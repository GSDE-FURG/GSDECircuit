//Converted to Combinational (Partial output: n80) , Module name: s1488_n80 , Timestamp: 2018-12-03T15:51:02.601892 
module s1488_n80 ( CLR, v7, v8, v2, v9, v1, v12, v11, v10, v6, v3, v5, v4, v0, n80 );
input CLR, v7, v8, v2, v9, v1, v12, v11, v10, v6, v3, v5, v4, v0;
output n80;
wire n267, n410, n416, n45, n403, n409, n415, n103, n79, n411, n63, n399, n402, n405, n408, n146, n154, n414, n413, n111, n236, n398, n401, n86, n400, n90, n109, n404, n406, n407, n82, n412, n230, n142, n397, n64, n72, n104, n68, n344, n61;
AOI21X1  g372(.A0(n416), .A1(n410), .B0(n267), .Y(n80));
INVX1    g222(.A(CLR), .Y(n267));
OAI21X1  g365(.A0(n409), .A1(n403), .B0(n45), .Y(n410));
AOI22X1  g371(.A0(n411), .A1(n79), .B0(n103), .B1(n415), .Y(n416));
INVX1    g000(.A(v7), .Y(n45));
AOI21X1  g358(.A0(n402), .A1(n399), .B0(n63), .Y(n403));
AOI21X1  g364(.A0(n408), .A1(n405), .B0(v8), .Y(n409));
OAI22X1  g370(.A0(n413), .A1(n414), .B0(n154), .B1(n146), .Y(n415));
INVX1    g058(.A(v2), .Y(n103));
AND2X1   g034(.A(v7), .B(v8), .Y(n79));
OAI22X1  g366(.A0(n236), .A1(n154), .B0(n111), .B1(n63), .Y(n411));
INVX1    g018(.A(v9), .Y(n63));
OR2X1    g354(.A(n398), .B(v1), .Y(n399));
AOI22X1  g357(.A0(n400), .A1(v12), .B0(n86), .B1(n401), .Y(n402));
NAND3X1  g360(.A(n404), .B(n109), .C(n90), .Y(n405));
OAI21X1  g363(.A0(n407), .A1(n406), .B0(v9), .Y(n408));
INVX1    g101(.A(n79), .Y(n146));
NAND2X1  g109(.A(n63), .B(v12), .Y(n154));
NAND3X1  g369(.A(n45), .B(v9), .C(n82), .Y(n414));
AOI21X1  g368(.A0(n230), .A1(n90), .B0(n412), .Y(n413));
OR2X1    g066(.A(v10), .B(v11), .Y(n111));
INVX1    g191(.A(n142), .Y(n236));
AOI21X1  g353(.A0(n64), .A1(v6), .B0(n397), .Y(n398));
OR2X1    g356(.A(n397), .B(n64), .Y(n401));
INVX1    g041(.A(v3), .Y(n86));
OAI21X1  g355(.A0(n72), .A1(v11), .B0(v10), .Y(n400));
AND2X1   g045(.A(v4), .B(v5), .Y(n90));
NOR2X1   g064(.A(n104), .B(v12), .Y(n109));
NOR3X1   g359(.A(v9), .B(n68), .C(v0), .Y(n404));
AOI21X1  g361(.A0(v10), .A1(n82), .B0(n104), .Y(n406));
AOI21X1  g362(.A0(n68), .A1(v6), .B0(n344), .Y(n407));
INVX1    g037(.A(v12), .Y(n82));
NOR2X1   g367(.A(v8), .B(v11), .Y(n412));
AND2X1   g185(.A(v8), .B(v11), .Y(n230));
NAND2X1  g097(.A(v10), .B(v11), .Y(n142));
NOR3X1   g352(.A(v8), .B(v11), .C(v12), .Y(n397));
AND2X1   g019(.A(v11), .B(v12), .Y(n64));
INVX1    g027(.A(v8), .Y(n72));
INVX1    g059(.A(v11), .Y(n104));
INVX1    g023(.A(v10), .Y(n68));
INVX1    g299(.A(n61), .Y(n344));
NOR2X1   g016(.A(v11), .B(v12), .Y(n61));

endmodule
