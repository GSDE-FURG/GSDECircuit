//Converted to Combinational (Partial output: n4250) , Module name: s38584_n4250 , Timestamp: 2018-12-03T15:51:17.159502 
module s38584_n4250 ( g35, g4917, g4922, g12, g16, g19, g28, g9, g7, g31, g6, g8, g2856, g2852, g4732, g5853, g3502, g46, g56, g57, g947, g1291, g53, g34, g54, g2999, g2912, g2917, g626, g772, g590, g1129, g1472, n4250 );
input g35, g4917, g4922, g12, g16, g19, g28, g9, g7, g31, g6, g8, g2856, g2852, g4732, g5853, g3502, g46, g56, g57, g947, g1291, g53, g34, g54, g2999, g2912, g2917, g626, g772, g590, g1129, g1472;
output n4250;
wire n8758, n6891_1, n6676, n5616, n5031, n5004, n5468, n5005, n4983, n5291, n5299_1, n5308_1, n5015, n5289_1, n5290, n5030, n5298, n5307, n5300, n5301, n5302, n4383, n5003, n5014, n5284_1, n5288, n5013, n5010, n4987, n5029, n5293, n5295, n5297, n5306, n5033, n5047_1, n5304, n4984_1, n4981, n5020, n5046, n5034, n5032_1, n4977, n4976, n5002_1, n4998, n4999, n5000, n5007_1, n5012_1, n5283, n5006, n5287, n4789, n4787, n5286, n5009, n4982, n5008, n5025, n5026, n5028, n5223, n5292, n5023, n5294_1, n5229, n5296, n5305, n5024, n5019, n5303_1, n4979_1, n4980, n4988_1, n5021, n4995, n5001, n4997_1, n5011, n5250_1, n5285, n5027_1, n5022_1, n4989, n4994, n4992_1, n4993, n4996;
MX2X1    g4112(.A(g4917), .B(n8758), .S0(g35), .Y(n4250));
MX2X1    g4111(.A(g4922), .B(n6676), .S0(n6891_1), .Y(n8758));
NOR3X1   g2249(.A(n5004), .B(n5031), .C(n5616), .Y(n6891_1));
INVX1    g1436(.A(n5468), .Y(n6676));
INVX1    g0976(.A(g12), .Y(n5616));
NAND3X1  g0411(.A(g19), .B(n5005), .C(g16), .Y(n5031));
NAND2X1  g0384(.A(n4983), .B(g28), .Y(n5004));
NOR3X1   g0828(.A(n5308_1), .B(n5299_1), .C(n5291), .Y(n5468));
INVX1    g0385(.A(g9), .Y(n5005));
NOR4X1   g0363(.A(g8), .B(g6), .C(g31), .D(g7), .Y(n4983));
AOI21X1  g0651(.A0(n5290), .A1(n5289_1), .B0(n5015), .Y(n5291));
NOR2X1   g0659(.A(n5298), .B(n5030), .Y(n5299_1));
NAND4X1  g0668(.A(n5302), .B(n5301), .C(n5300), .D(n5307), .Y(n5308_1));
OAI21X1  g0395(.A0(n5014), .A1(n5003), .B0(n4383), .Y(n5015));
NOR2X1   g0649(.A(n5288), .B(n5284_1), .Y(n5289_1));
AOI22X1  g0650(.A0(n5010), .A1(g2852), .B0(g2856), .B1(n5013), .Y(n5290));
OR2X1    g0410(.A(n5029), .B(n4987), .Y(n5030));
NOR3X1   g0658(.A(n5297), .B(n5295), .C(n5293), .Y(n5298));
AOI22X1  g0667(.A0(n5304), .A1(n5047_1), .B0(n5033), .B1(n5306), .Y(n5307));
NAND4X1  g0660(.A(n4981), .B(n4383), .C(g4732), .D(n4984_1), .Y(n5300));
AOI22X1  g0661(.A0(n5046), .A1(g3502), .B0(g5853), .B1(n5020), .Y(n5301));
AOI22X1  g0662(.A0(n5032_1), .A1(g4922), .B0(g46), .B1(n5034), .Y(n5302));
NOR4X1   g0358(.A(n4976), .B(g57), .C(g56), .D(n4977), .Y(n4383));
OR4X1    g0383(.A(n5000), .B(n4999), .C(n4998), .D(n5002_1), .Y(n5003));
OR4X1    g0394(.A(n5012_1), .B(n5010), .C(n5007_1), .D(n5013), .Y(n5014));
NOR3X1   g0644(.A(n5006), .B(n5004), .C(n5283), .Y(n5284_1));
OAI22X1  g0648(.A0(n5286), .A1(n4787), .B0(n4789), .B1(n5287), .Y(n5288));
NOR4X1   g0393(.A(n5008), .B(n4982), .C(n5005), .D(n5009), .Y(n5013));
NOR4X1   g0390(.A(n5008), .B(g28), .C(n5005), .D(n5009), .Y(n5010));
OR4X1    g0367(.A(n4976), .B(g57), .C(g56), .D(n4977), .Y(n4987));
NOR3X1   g0409(.A(n5028), .B(n5026), .C(n5025), .Y(n5029));
AOI21X1  g0653(.A0(n5292), .A1(g35), .B0(n5223), .Y(n5293));
AOI21X1  g0655(.A0(n5294_1), .A1(g35), .B0(n5023), .Y(n5295));
AOI21X1  g0657(.A0(n5296), .A1(g35), .B0(n5229), .Y(n5297));
NOR2X1   g0666(.A(g947), .B(n5305), .Y(n5306));
NOR3X1   g0413(.A(n5024), .B(n5004), .C(n4987), .Y(n5033));
NOR3X1   g0427(.A(n5006), .B(n5019), .C(n4987), .Y(n5047_1));
NOR2X1   g0664(.A(g1291), .B(n5303_1), .Y(n5304));
AND2X1   g0364(.A(n4983), .B(n4982), .Y(n4984_1));
NOR3X1   g0361(.A(n4980), .B(g9), .C(n4979_1), .Y(n4981));
NOR3X1   g0400(.A(n4988_1), .B(n5019), .C(n4987), .Y(n5020));
NOR3X1   g0426(.A(n5021), .B(n4988_1), .C(n4987), .Y(n5046));
NOR2X1   g0414(.A(n4383), .B(g53), .Y(n5034));
NOR3X1   g0412(.A(n5004), .B(n5031), .C(n4987), .Y(n5032_1));
OR2X1    g0357(.A(g34), .B(g53), .Y(n4977));
INVX1    g0356(.A(g54), .Y(n4976));
NOR3X1   g0382(.A(n5001), .B(n4995), .C(g28), .Y(n5002_1));
NOR3X1   g0378(.A(n4997_1), .B(n4995), .C(g28), .Y(n4998));
NOR3X1   g0379(.A(n4995), .B(n4988_1), .C(n4982), .Y(n4999));
NOR3X1   g0380(.A(n4997_1), .B(n4995), .C(n4982), .Y(n5000));
NOR2X1   g0387(.A(n5006), .B(n5004), .Y(n5007_1));
NOR2X1   g0392(.A(n5011), .B(n5006), .Y(n5012_1));
INVX1    g0643(.A(g2999), .Y(n5283));
NAND3X1  g0386(.A(n4980), .B(n5005), .C(g16), .Y(n5006));
NAND3X1  g0647(.A(n5285), .B(n5250_1), .C(g28), .Y(n5287));
INVX1    g0169(.A(g2912), .Y(n4789));
INVX1    g0167(.A(g2917), .Y(n4787));
NAND3X1  g0646(.A(n5285), .B(n5250_1), .C(n4982), .Y(n5286));
OR2X1    g0389(.A(g19), .B(g16), .Y(n5009));
INVX1    g0362(.A(g28), .Y(n4982));
OR4X1    g0388(.A(g8), .B(g6), .C(g31), .D(g7), .Y(n5008));
OAI21X1  g0405(.A0(n5024), .A1(n5021), .B0(n5023), .Y(n5025));
NOR4X1   g0406(.A(n5008), .B(g28), .C(g9), .D(n5009), .Y(n5026));
OAI21X1  g0408(.A0(n5024), .A1(n5019), .B0(n5027_1), .Y(n5028));
OR2X1    g0583(.A(n5024), .B(n5019), .Y(n5223));
INVX1    g0652(.A(g626), .Y(n5292));
NAND4X1  g0403(.A(n4989), .B(g28), .C(g31), .D(n5022_1), .Y(n5023));
INVX1    g0654(.A(g772), .Y(n5294_1));
OR2X1    g0589(.A(n5024), .B(n5021), .Y(n5229));
INVX1    g0656(.A(g590), .Y(n5296));
INVX1    g0665(.A(g1129), .Y(n5305));
NAND3X1  g0404(.A(g19), .B(n5005), .C(n4979_1), .Y(n5024));
NAND2X1  g0399(.A(n4983), .B(n4982), .Y(n5019));
INVX1    g0663(.A(g1472), .Y(n5303_1));
INVX1    g0359(.A(g16), .Y(n4979_1));
INVX1    g0360(.A(g19), .Y(n4980));
NAND3X1  g0368(.A(g19), .B(g9), .C(n4979_1), .Y(n4988_1));
NAND3X1  g0401(.A(n4989), .B(n4982), .C(g31), .Y(n5021));
OR4X1    g0375(.A(n4993), .B(n4992_1), .C(g31), .D(n4994), .Y(n4995));
NAND3X1  g0381(.A(n4980), .B(g9), .C(g16), .Y(n5001));
NAND2X1  g0377(.A(n4996), .B(g9), .Y(n4997_1));
NAND3X1  g0391(.A(n4989), .B(g28), .C(g31), .Y(n5011));
NOR4X1   g0610(.A(n4993), .B(n4992_1), .C(g31), .D(n4994), .Y(n5250_1));
NOR2X1   g0645(.A(n5009), .B(n5005), .Y(n5285));
NAND3X1  g0407(.A(n5022_1), .B(n4983), .C(g28), .Y(n5027_1));
NOR3X1   g0402(.A(g19), .B(g9), .C(g16), .Y(n5022_1));
NOR3X1   g0369(.A(g7), .B(g8), .C(g6), .Y(n4989));
INVX1    g0374(.A(g7), .Y(n4994));
INVX1    g0372(.A(g6), .Y(n4992_1));
INVX1    g0373(.A(g8), .Y(n4993));
NOR2X1   g0376(.A(g19), .B(g16), .Y(n4996));

endmodule
