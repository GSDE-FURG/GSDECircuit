// Benchmark "top" written by ABC on Mon Sep 21 04:05:09 2020

module top ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] ,
    \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] ;
  output \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F;
  wire new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n331_, new_n332_, new_n333_, new_n334_, new_n335_,
    new_n336_, new_n337_, new_n338_, new_n339_, new_n340_, new_n341_,
    new_n342_, new_n343_, new_n344_, new_n345_, new_n346_, new_n347_,
    new_n348_, new_n349_, new_n350_, new_n351_, new_n352_, new_n353_,
    new_n354_, new_n355_, new_n356_, new_n357_, new_n358_, new_n359_,
    new_n360_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n430_, new_n431_,
    new_n432_, new_n433_, new_n434_, new_n435_, new_n436_, new_n437_,
    new_n438_, new_n439_, new_n440_, new_n441_, new_n442_, new_n443_,
    new_n444_, new_n445_, new_n446_, new_n447_, new_n448_, new_n449_,
    new_n450_, new_n451_, new_n452_, new_n453_, new_n454_, new_n455_,
    new_n456_, new_n457_, new_n458_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n480_, new_n481_, new_n482_, new_n483_, new_n484_, new_n485_,
    new_n486_, new_n487_, new_n488_, new_n489_, new_n490_, new_n491_,
    new_n492_, new_n493_, new_n494_, new_n495_, new_n496_, new_n497_,
    new_n498_, new_n499_, new_n500_, new_n501_, new_n502_, new_n503_,
    new_n504_, new_n505_, new_n506_, new_n507_, new_n508_, new_n509_,
    new_n510_, new_n511_, new_n512_, new_n513_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n522_,
    new_n523_, new_n524_, new_n525_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n530_, new_n531_, new_n532_, new_n533_, new_n534_,
    new_n535_, new_n536_, new_n537_, new_n538_, new_n539_, new_n540_,
    new_n541_, new_n542_, new_n543_, new_n544_, new_n545_, new_n546_,
    new_n547_, new_n548_, new_n549_, new_n550_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n558_,
    new_n559_, new_n560_, new_n561_, new_n562_, new_n563_, new_n564_,
    new_n565_, new_n566_, new_n567_, new_n568_, new_n569_, new_n570_,
    new_n571_, new_n572_, new_n573_, new_n574_, new_n575_, new_n576_,
    new_n577_, new_n578_, new_n579_, new_n580_, new_n581_, new_n582_,
    new_n583_, new_n584_, new_n585_, new_n587_, new_n588_, new_n589_,
    new_n590_, new_n591_, new_n592_, new_n593_, new_n594_, new_n595_,
    new_n596_, new_n597_, new_n598_, new_n599_, new_n600_, new_n601_,
    new_n602_, new_n603_, new_n604_, new_n605_, new_n606_, new_n607_,
    new_n608_, new_n609_, new_n610_, new_n611_, new_n612_, new_n613_,
    new_n614_, new_n615_, new_n616_, new_n617_, new_n618_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n653_, new_n654_, new_n655_, new_n657_, new_n659_,
    new_n660_;
  INVX1    g000(.A(\A[12] ), .Y(new_n137_));
  INVX1    g001(.A(\A[22] ), .Y(new_n138_));
  INVX1    g002(.A(\A[24] ), .Y(new_n139_));
  INVX1    g003(.A(\A[26] ), .Y(new_n140_));
  INVX1    g004(.A(\A[32] ), .Y(new_n141_));
  INVX1    g005(.A(\A[34] ), .Y(new_n142_));
  INVX1    g006(.A(\A[36] ), .Y(new_n143_));
  INVX1    g007(.A(\A[42] ), .Y(new_n144_));
  INVX1    g008(.A(\A[44] ), .Y(new_n145_));
  INVX1    g009(.A(\A[46] ), .Y(new_n146_));
  INVX1    g010(.A(\A[52] ), .Y(new_n147_));
  INVX1    g011(.A(\A[54] ), .Y(new_n148_));
  INVX1    g012(.A(\A[56] ), .Y(new_n149_));
  INVX1    g013(.A(\A[62] ), .Y(new_n150_));
  INVX1    g014(.A(\A[64] ), .Y(new_n151_));
  INVX1    g015(.A(\A[66] ), .Y(new_n152_));
  INVX1    g016(.A(\A[72] ), .Y(new_n153_));
  INVX1    g017(.A(\A[74] ), .Y(new_n154_));
  INVX1    g018(.A(\A[76] ), .Y(new_n155_));
  INVX1    g019(.A(\A[82] ), .Y(new_n156_));
  INVX1    g020(.A(\A[84] ), .Y(new_n157_));
  INVX1    g021(.A(\A[86] ), .Y(new_n158_));
  INVX1    g022(.A(\A[88] ), .Y(new_n159_));
  INVX1    g023(.A(\A[90] ), .Y(new_n160_));
  INVX1    g024(.A(\A[92] ), .Y(new_n161_));
  INVX1    g025(.A(\A[94] ), .Y(new_n162_));
  INVX1    g026(.A(\A[96] ), .Y(new_n163_));
  INVX1    g027(.A(\A[98] ), .Y(new_n164_));
  INVX1    g028(.A(\A[102] ), .Y(new_n165_));
  INVX1    g029(.A(\A[106] ), .Y(new_n166_));
  INVX1    g030(.A(\A[108] ), .Y(new_n167_));
  INVX1    g031(.A(\A[120] ), .Y(new_n168_));
  INVX1    g032(.A(\A[126] ), .Y(new_n169_));
  NOR2X1   g033(.A(\A[127] ), .B(new_n169_), .Y(new_n170_));
  AOI21X1  g034(.A0(new_n169_), .A1(\A[125] ), .B0(\A[127] ), .Y(new_n171_));
  MX2X1    g035(.A(new_n170_), .B(new_n171_), .S0(\A[124] ), .Y(new_n172_));
  MX2X1    g036(.A(new_n171_), .B(new_n172_), .S0(\A[123] ), .Y(new_n173_));
  MX2X1    g037(.A(new_n172_), .B(new_n173_), .S0(\A[122] ), .Y(new_n174_));
  MX2X1    g038(.A(new_n173_), .B(new_n174_), .S0(\A[121] ), .Y(new_n175_));
  MX2X1    g039(.A(new_n175_), .B(new_n174_), .S0(new_n168_), .Y(new_n176_));
  MX2X1    g040(.A(new_n175_), .B(new_n176_), .S0(\A[119] ), .Y(new_n177_));
  MX2X1    g041(.A(new_n176_), .B(new_n177_), .S0(\A[118] ), .Y(new_n178_));
  MX2X1    g042(.A(new_n177_), .B(new_n178_), .S0(\A[117] ), .Y(new_n179_));
  MX2X1    g043(.A(new_n178_), .B(new_n179_), .S0(\A[116] ), .Y(new_n180_));
  MX2X1    g044(.A(new_n179_), .B(new_n180_), .S0(\A[115] ), .Y(new_n181_));
  MX2X1    g045(.A(new_n180_), .B(new_n181_), .S0(\A[114] ), .Y(new_n182_));
  MX2X1    g046(.A(new_n181_), .B(new_n182_), .S0(\A[113] ), .Y(new_n183_));
  MX2X1    g047(.A(new_n182_), .B(new_n183_), .S0(\A[112] ), .Y(new_n184_));
  MX2X1    g048(.A(new_n183_), .B(new_n184_), .S0(\A[111] ), .Y(new_n185_));
  MX2X1    g049(.A(new_n184_), .B(new_n185_), .S0(\A[110] ), .Y(new_n186_));
  INVX1    g050(.A(\A[109] ), .Y(new_n187_));
  MX2X1    g051(.A(new_n186_), .B(new_n185_), .S0(new_n187_), .Y(new_n188_));
  MX2X1    g052(.A(new_n188_), .B(new_n186_), .S0(new_n167_), .Y(new_n189_));
  INVX1    g053(.A(\A[107] ), .Y(new_n190_));
  MX2X1    g054(.A(new_n189_), .B(new_n188_), .S0(new_n190_), .Y(new_n191_));
  MX2X1    g055(.A(new_n191_), .B(new_n189_), .S0(new_n166_), .Y(new_n192_));
  MX2X1    g056(.A(new_n191_), .B(new_n192_), .S0(\A[105] ), .Y(new_n193_));
  MX2X1    g057(.A(new_n192_), .B(new_n193_), .S0(\A[104] ), .Y(new_n194_));
  INVX1    g058(.A(\A[103] ), .Y(new_n195_));
  MX2X1    g059(.A(new_n194_), .B(new_n193_), .S0(new_n195_), .Y(new_n196_));
  MX2X1    g060(.A(new_n196_), .B(new_n194_), .S0(new_n165_), .Y(new_n197_));
  MX2X1    g061(.A(new_n196_), .B(new_n197_), .S0(\A[101] ), .Y(new_n198_));
  MX2X1    g062(.A(new_n197_), .B(new_n198_), .S0(\A[100] ), .Y(new_n199_));
  INVX1    g063(.A(\A[99] ), .Y(new_n200_));
  MX2X1    g064(.A(new_n199_), .B(new_n198_), .S0(new_n200_), .Y(new_n201_));
  MX2X1    g065(.A(new_n201_), .B(new_n199_), .S0(new_n164_), .Y(new_n202_));
  INVX1    g066(.A(\A[97] ), .Y(new_n203_));
  MX2X1    g067(.A(new_n202_), .B(new_n201_), .S0(new_n203_), .Y(new_n204_));
  MX2X1    g068(.A(new_n204_), .B(new_n202_), .S0(new_n163_), .Y(new_n205_));
  INVX1    g069(.A(\A[95] ), .Y(new_n206_));
  MX2X1    g070(.A(new_n205_), .B(new_n204_), .S0(new_n206_), .Y(new_n207_));
  MX2X1    g071(.A(new_n207_), .B(new_n205_), .S0(new_n162_), .Y(new_n208_));
  INVX1    g072(.A(\A[93] ), .Y(new_n209_));
  MX2X1    g073(.A(new_n208_), .B(new_n207_), .S0(new_n209_), .Y(new_n210_));
  MX2X1    g074(.A(new_n210_), .B(new_n208_), .S0(new_n161_), .Y(new_n211_));
  INVX1    g075(.A(\A[91] ), .Y(new_n212_));
  MX2X1    g076(.A(new_n211_), .B(new_n210_), .S0(new_n212_), .Y(new_n213_));
  MX2X1    g077(.A(new_n213_), .B(new_n211_), .S0(new_n160_), .Y(new_n214_));
  INVX1    g078(.A(\A[89] ), .Y(new_n215_));
  MX2X1    g079(.A(new_n214_), .B(new_n213_), .S0(new_n215_), .Y(new_n216_));
  MX2X1    g080(.A(new_n216_), .B(new_n214_), .S0(new_n159_), .Y(new_n217_));
  INVX1    g081(.A(\A[87] ), .Y(new_n218_));
  MX2X1    g082(.A(new_n217_), .B(new_n216_), .S0(new_n218_), .Y(new_n219_));
  MX2X1    g083(.A(new_n219_), .B(new_n217_), .S0(new_n158_), .Y(new_n220_));
  INVX1    g084(.A(\A[85] ), .Y(new_n221_));
  MX2X1    g085(.A(new_n220_), .B(new_n219_), .S0(new_n221_), .Y(new_n222_));
  MX2X1    g086(.A(new_n222_), .B(new_n220_), .S0(new_n157_), .Y(new_n223_));
  INVX1    g087(.A(\A[83] ), .Y(new_n224_));
  MX2X1    g088(.A(new_n223_), .B(new_n222_), .S0(new_n224_), .Y(new_n225_));
  MX2X1    g089(.A(new_n225_), .B(new_n223_), .S0(new_n156_), .Y(new_n226_));
  MX2X1    g090(.A(new_n225_), .B(new_n226_), .S0(\A[81] ), .Y(new_n227_));
  MX2X1    g091(.A(new_n226_), .B(new_n227_), .S0(\A[80] ), .Y(new_n228_));
  MX2X1    g092(.A(new_n227_), .B(new_n228_), .S0(\A[79] ), .Y(new_n229_));
  MX2X1    g093(.A(new_n228_), .B(new_n229_), .S0(\A[78] ), .Y(new_n230_));
  INVX1    g094(.A(\A[77] ), .Y(new_n231_));
  MX2X1    g095(.A(new_n230_), .B(new_n229_), .S0(new_n231_), .Y(new_n232_));
  MX2X1    g096(.A(new_n232_), .B(new_n230_), .S0(new_n155_), .Y(new_n233_));
  INVX1    g097(.A(\A[75] ), .Y(new_n234_));
  MX2X1    g098(.A(new_n233_), .B(new_n232_), .S0(new_n234_), .Y(new_n235_));
  MX2X1    g099(.A(new_n235_), .B(new_n233_), .S0(new_n154_), .Y(new_n236_));
  INVX1    g100(.A(\A[73] ), .Y(new_n237_));
  MX2X1    g101(.A(new_n236_), .B(new_n235_), .S0(new_n237_), .Y(new_n238_));
  MX2X1    g102(.A(new_n238_), .B(new_n236_), .S0(new_n153_), .Y(new_n239_));
  MX2X1    g103(.A(new_n238_), .B(new_n239_), .S0(\A[71] ), .Y(new_n240_));
  MX2X1    g104(.A(new_n239_), .B(new_n240_), .S0(\A[70] ), .Y(new_n241_));
  MX2X1    g105(.A(new_n240_), .B(new_n241_), .S0(\A[69] ), .Y(new_n242_));
  MX2X1    g106(.A(new_n241_), .B(new_n242_), .S0(\A[68] ), .Y(new_n243_));
  INVX1    g107(.A(\A[67] ), .Y(new_n244_));
  MX2X1    g108(.A(new_n243_), .B(new_n242_), .S0(new_n244_), .Y(new_n245_));
  MX2X1    g109(.A(new_n245_), .B(new_n243_), .S0(new_n152_), .Y(new_n246_));
  INVX1    g110(.A(\A[65] ), .Y(new_n247_));
  MX2X1    g111(.A(new_n246_), .B(new_n245_), .S0(new_n247_), .Y(new_n248_));
  MX2X1    g112(.A(new_n248_), .B(new_n246_), .S0(new_n151_), .Y(new_n249_));
  INVX1    g113(.A(\A[63] ), .Y(new_n250_));
  MX2X1    g114(.A(new_n249_), .B(new_n248_), .S0(new_n250_), .Y(new_n251_));
  MX2X1    g115(.A(new_n251_), .B(new_n249_), .S0(new_n150_), .Y(new_n252_));
  MX2X1    g116(.A(new_n251_), .B(new_n252_), .S0(\A[61] ), .Y(new_n253_));
  MX2X1    g117(.A(new_n252_), .B(new_n253_), .S0(\A[60] ), .Y(new_n254_));
  MX2X1    g118(.A(new_n253_), .B(new_n254_), .S0(\A[59] ), .Y(new_n255_));
  MX2X1    g119(.A(new_n254_), .B(new_n255_), .S0(\A[58] ), .Y(new_n256_));
  INVX1    g120(.A(\A[57] ), .Y(new_n257_));
  MX2X1    g121(.A(new_n256_), .B(new_n255_), .S0(new_n257_), .Y(new_n258_));
  MX2X1    g122(.A(new_n258_), .B(new_n256_), .S0(new_n149_), .Y(new_n259_));
  INVX1    g123(.A(\A[55] ), .Y(new_n260_));
  MX2X1    g124(.A(new_n259_), .B(new_n258_), .S0(new_n260_), .Y(new_n261_));
  MX2X1    g125(.A(new_n261_), .B(new_n259_), .S0(new_n148_), .Y(new_n262_));
  INVX1    g126(.A(\A[53] ), .Y(new_n263_));
  MX2X1    g127(.A(new_n262_), .B(new_n261_), .S0(new_n263_), .Y(new_n264_));
  MX2X1    g128(.A(new_n264_), .B(new_n262_), .S0(new_n147_), .Y(new_n265_));
  MX2X1    g129(.A(new_n264_), .B(new_n265_), .S0(\A[51] ), .Y(new_n266_));
  MX2X1    g130(.A(new_n265_), .B(new_n266_), .S0(\A[50] ), .Y(new_n267_));
  MX2X1    g131(.A(new_n266_), .B(new_n267_), .S0(\A[49] ), .Y(new_n268_));
  MX2X1    g132(.A(new_n267_), .B(new_n268_), .S0(\A[48] ), .Y(new_n269_));
  INVX1    g133(.A(\A[47] ), .Y(new_n270_));
  MX2X1    g134(.A(new_n269_), .B(new_n268_), .S0(new_n270_), .Y(new_n271_));
  MX2X1    g135(.A(new_n271_), .B(new_n269_), .S0(new_n146_), .Y(new_n272_));
  INVX1    g136(.A(\A[45] ), .Y(new_n273_));
  MX2X1    g137(.A(new_n272_), .B(new_n271_), .S0(new_n273_), .Y(new_n274_));
  MX2X1    g138(.A(new_n274_), .B(new_n272_), .S0(new_n145_), .Y(new_n275_));
  INVX1    g139(.A(\A[43] ), .Y(new_n276_));
  MX2X1    g140(.A(new_n275_), .B(new_n274_), .S0(new_n276_), .Y(new_n277_));
  MX2X1    g141(.A(new_n277_), .B(new_n275_), .S0(new_n144_), .Y(new_n278_));
  MX2X1    g142(.A(new_n277_), .B(new_n278_), .S0(\A[41] ), .Y(new_n279_));
  MX2X1    g143(.A(new_n278_), .B(new_n279_), .S0(\A[40] ), .Y(new_n280_));
  MX2X1    g144(.A(new_n279_), .B(new_n280_), .S0(\A[39] ), .Y(new_n281_));
  MX2X1    g145(.A(new_n280_), .B(new_n281_), .S0(\A[38] ), .Y(new_n282_));
  INVX1    g146(.A(\A[37] ), .Y(new_n283_));
  MX2X1    g147(.A(new_n282_), .B(new_n281_), .S0(new_n283_), .Y(new_n284_));
  MX2X1    g148(.A(new_n284_), .B(new_n282_), .S0(new_n143_), .Y(new_n285_));
  INVX1    g149(.A(\A[35] ), .Y(new_n286_));
  MX2X1    g150(.A(new_n285_), .B(new_n284_), .S0(new_n286_), .Y(new_n287_));
  MX2X1    g151(.A(new_n287_), .B(new_n285_), .S0(new_n142_), .Y(new_n288_));
  INVX1    g152(.A(\A[33] ), .Y(new_n289_));
  MX2X1    g153(.A(new_n288_), .B(new_n287_), .S0(new_n289_), .Y(new_n290_));
  MX2X1    g154(.A(new_n290_), .B(new_n288_), .S0(new_n141_), .Y(new_n291_));
  MX2X1    g155(.A(new_n290_), .B(new_n291_), .S0(\A[31] ), .Y(new_n292_));
  MX2X1    g156(.A(new_n291_), .B(new_n292_), .S0(\A[30] ), .Y(new_n293_));
  MX2X1    g157(.A(new_n292_), .B(new_n293_), .S0(\A[29] ), .Y(new_n294_));
  MX2X1    g158(.A(new_n293_), .B(new_n294_), .S0(\A[28] ), .Y(new_n295_));
  INVX1    g159(.A(\A[27] ), .Y(new_n296_));
  MX2X1    g160(.A(new_n295_), .B(new_n294_), .S0(new_n296_), .Y(new_n297_));
  MX2X1    g161(.A(new_n297_), .B(new_n295_), .S0(new_n140_), .Y(new_n298_));
  INVX1    g162(.A(\A[25] ), .Y(new_n299_));
  MX2X1    g163(.A(new_n298_), .B(new_n297_), .S0(new_n299_), .Y(new_n300_));
  MX2X1    g164(.A(new_n300_), .B(new_n298_), .S0(new_n139_), .Y(new_n301_));
  INVX1    g165(.A(\A[23] ), .Y(new_n302_));
  MX2X1    g166(.A(new_n301_), .B(new_n300_), .S0(new_n302_), .Y(new_n303_));
  MX2X1    g167(.A(new_n303_), .B(new_n301_), .S0(new_n138_), .Y(new_n304_));
  MX2X1    g168(.A(new_n303_), .B(new_n304_), .S0(\A[21] ), .Y(new_n305_));
  MX2X1    g169(.A(new_n304_), .B(new_n305_), .S0(\A[20] ), .Y(new_n306_));
  MX2X1    g170(.A(new_n305_), .B(new_n306_), .S0(\A[19] ), .Y(new_n307_));
  MX2X1    g171(.A(new_n306_), .B(new_n307_), .S0(\A[18] ), .Y(new_n308_));
  MX2X1    g172(.A(new_n307_), .B(new_n308_), .S0(\A[17] ), .Y(new_n309_));
  MX2X1    g173(.A(new_n308_), .B(new_n309_), .S0(\A[16] ), .Y(new_n310_));
  MX2X1    g174(.A(new_n309_), .B(new_n310_), .S0(\A[15] ), .Y(new_n311_));
  MX2X1    g175(.A(new_n310_), .B(new_n311_), .S0(\A[14] ), .Y(new_n312_));
  INVX1    g176(.A(\A[13] ), .Y(new_n313_));
  MX2X1    g177(.A(new_n312_), .B(new_n311_), .S0(new_n313_), .Y(new_n314_));
  MX2X1    g178(.A(new_n314_), .B(new_n312_), .S0(new_n137_), .Y(new_n315_));
  MX2X1    g179(.A(new_n314_), .B(new_n315_), .S0(\A[11] ), .Y(new_n316_));
  MX2X1    g180(.A(new_n315_), .B(new_n316_), .S0(\A[10] ), .Y(new_n317_));
  MX2X1    g181(.A(new_n316_), .B(new_n317_), .S0(\A[9] ), .Y(new_n318_));
  MX2X1    g182(.A(new_n317_), .B(new_n318_), .S0(\A[8] ), .Y(new_n319_));
  MX2X1    g183(.A(new_n318_), .B(new_n319_), .S0(\A[7] ), .Y(new_n320_));
  MX2X1    g184(.A(new_n319_), .B(new_n320_), .S0(\A[6] ), .Y(new_n321_));
  MX2X1    g185(.A(new_n320_), .B(new_n321_), .S0(\A[5] ), .Y(new_n322_));
  MX2X1    g186(.A(new_n321_), .B(new_n322_), .S0(\A[4] ), .Y(new_n323_));
  INVX1    g187(.A(\A[3] ), .Y(new_n324_));
  OR2X1    g188(.A(new_n323_), .B(new_n324_), .Y(new_n325_));
  INVX1    g189(.A(\A[2] ), .Y(new_n326_));
  AND2X1   g190(.A(new_n326_), .B(\A[1] ), .Y(new_n327_));
  NOR2X1   g191(.A(new_n322_), .B(\A[3] ), .Y(new_n328_));
  NOR2X1   g192(.A(new_n327_), .B(new_n328_), .Y(new_n329_));
  AOI22X1  g193(.A0(new_n329_), .A1(new_n325_), .B0(new_n327_), .B1(new_n323_), .Y(\P[0] ));
  NOR2X1   g194(.A(\A[127] ), .B(\A[126] ), .Y(new_n331_));
  NOR2X1   g195(.A(\A[125] ), .B(\A[124] ), .Y(new_n332_));
  INVX1    g196(.A(new_n332_), .Y(new_n333_));
  NOR2X1   g197(.A(\A[123] ), .B(\A[122] ), .Y(new_n334_));
  OAI21X1  g198(.A0(new_n334_), .A1(new_n333_), .B0(new_n331_), .Y(new_n335_));
  INVX1    g199(.A(new_n331_), .Y(new_n336_));
  AOI21X1  g200(.A0(new_n334_), .A1(\A[121] ), .B0(new_n333_), .Y(new_n337_));
  OR2X1    g201(.A(new_n337_), .B(new_n336_), .Y(new_n338_));
  MX2X1    g202(.A(new_n335_), .B(new_n338_), .S0(new_n168_), .Y(new_n339_));
  NOR2X1   g203(.A(\A[119] ), .B(\A[118] ), .Y(new_n340_));
  MX2X1    g204(.A(new_n339_), .B(new_n335_), .S0(new_n340_), .Y(new_n341_));
  NOR2X1   g205(.A(\A[117] ), .B(\A[116] ), .Y(new_n342_));
  MX2X1    g206(.A(new_n341_), .B(new_n339_), .S0(new_n342_), .Y(new_n343_));
  NOR2X1   g207(.A(\A[115] ), .B(\A[114] ), .Y(new_n344_));
  MX2X1    g208(.A(new_n343_), .B(new_n341_), .S0(new_n344_), .Y(new_n345_));
  NOR2X1   g209(.A(\A[113] ), .B(\A[112] ), .Y(new_n346_));
  MX2X1    g210(.A(new_n345_), .B(new_n343_), .S0(new_n346_), .Y(new_n347_));
  OR2X1    g211(.A(\A[111] ), .B(\A[110] ), .Y(new_n348_));
  MX2X1    g212(.A(new_n345_), .B(new_n347_), .S0(new_n348_), .Y(new_n349_));
  OR2X1    g213(.A(\A[109] ), .B(\A[108] ), .Y(new_n350_));
  AND2X1   g214(.A(new_n350_), .B(new_n349_), .Y(new_n351_));
  INVX1    g215(.A(new_n351_), .Y(new_n352_));
  NAND3X1  g216(.A(new_n347_), .B(new_n187_), .C(new_n167_), .Y(new_n353_));
  AND2X1   g217(.A(new_n353_), .B(new_n352_), .Y(new_n354_));
  OR2X1    g218(.A(\A[107] ), .B(\A[106] ), .Y(new_n355_));
  AND2X1   g219(.A(new_n355_), .B(new_n354_), .Y(new_n356_));
  NOR2X1   g220(.A(new_n355_), .B(new_n349_), .Y(new_n357_));
  NOR2X1   g221(.A(\A[105] ), .B(\A[104] ), .Y(new_n358_));
  NOR3X1   g222(.A(new_n358_), .B(new_n357_), .C(new_n356_), .Y(new_n359_));
  NOR3X1   g223(.A(new_n354_), .B(\A[105] ), .C(\A[104] ), .Y(new_n360_));
  NOR2X1   g224(.A(new_n360_), .B(new_n359_), .Y(new_n361_));
  NOR2X1   g225(.A(\A[103] ), .B(\A[102] ), .Y(new_n362_));
  NOR3X1   g226(.A(new_n362_), .B(new_n360_), .C(new_n359_), .Y(new_n363_));
  AOI21X1  g227(.A0(new_n355_), .A1(new_n354_), .B0(new_n357_), .Y(new_n364_));
  NOR3X1   g228(.A(new_n364_), .B(\A[103] ), .C(\A[102] ), .Y(new_n365_));
  NOR2X1   g229(.A(new_n365_), .B(new_n363_), .Y(new_n366_));
  INVX1    g230(.A(new_n366_), .Y(new_n367_));
  OR2X1    g231(.A(\A[101] ), .B(\A[100] ), .Y(new_n368_));
  MX2X1    g232(.A(new_n361_), .B(new_n367_), .S0(new_n368_), .Y(new_n369_));
  OR2X1    g233(.A(\A[99] ), .B(\A[98] ), .Y(new_n370_));
  NOR2X1   g234(.A(new_n370_), .B(new_n366_), .Y(new_n371_));
  AOI21X1  g235(.A0(new_n370_), .A1(new_n369_), .B0(new_n371_), .Y(new_n372_));
  OR2X1    g236(.A(\A[97] ), .B(\A[96] ), .Y(new_n373_));
  NOR2X1   g237(.A(new_n373_), .B(new_n369_), .Y(new_n374_));
  AOI21X1  g238(.A0(new_n373_), .A1(new_n372_), .B0(new_n374_), .Y(new_n375_));
  OR2X1    g239(.A(\A[95] ), .B(\A[94] ), .Y(new_n376_));
  NOR2X1   g240(.A(new_n376_), .B(new_n372_), .Y(new_n377_));
  AOI21X1  g241(.A0(new_n376_), .A1(new_n375_), .B0(new_n377_), .Y(new_n378_));
  INVX1    g242(.A(new_n378_), .Y(new_n379_));
  OR2X1    g243(.A(\A[93] ), .B(\A[92] ), .Y(new_n380_));
  NOR2X1   g244(.A(new_n380_), .B(new_n375_), .Y(new_n381_));
  AOI21X1  g245(.A0(new_n380_), .A1(new_n378_), .B0(new_n381_), .Y(new_n382_));
  NOR2X1   g246(.A(\A[91] ), .B(\A[90] ), .Y(new_n383_));
  MX2X1    g247(.A(new_n382_), .B(new_n379_), .S0(new_n383_), .Y(new_n384_));
  AOI21X1  g248(.A0(new_n215_), .A1(new_n159_), .B0(new_n384_), .Y(new_n385_));
  NOR3X1   g249(.A(new_n382_), .B(\A[89] ), .C(\A[88] ), .Y(new_n386_));
  OR2X1    g250(.A(new_n386_), .B(new_n385_), .Y(new_n387_));
  INVX1    g251(.A(new_n387_), .Y(new_n388_));
  NOR2X1   g252(.A(\A[87] ), .B(\A[86] ), .Y(new_n389_));
  NAND3X1  g253(.A(new_n384_), .B(new_n218_), .C(new_n158_), .Y(new_n390_));
  OAI21X1  g254(.A0(new_n389_), .A1(new_n387_), .B0(new_n390_), .Y(new_n391_));
  NOR2X1   g255(.A(\A[85] ), .B(\A[84] ), .Y(new_n392_));
  MX2X1    g256(.A(new_n391_), .B(new_n388_), .S0(new_n392_), .Y(new_n393_));
  OAI21X1  g257(.A0(\A[83] ), .A1(\A[82] ), .B0(new_n393_), .Y(new_n394_));
  NAND3X1  g258(.A(new_n391_), .B(new_n224_), .C(new_n156_), .Y(new_n395_));
  AND2X1   g259(.A(new_n395_), .B(new_n394_), .Y(new_n396_));
  INVX1    g260(.A(new_n396_), .Y(new_n397_));
  OR2X1    g261(.A(\A[81] ), .B(\A[80] ), .Y(new_n398_));
  NOR2X1   g262(.A(new_n398_), .B(new_n393_), .Y(new_n399_));
  AOI21X1  g263(.A0(new_n398_), .A1(new_n396_), .B0(new_n399_), .Y(new_n400_));
  NOR2X1   g264(.A(\A[79] ), .B(\A[78] ), .Y(new_n401_));
  MX2X1    g265(.A(new_n400_), .B(new_n397_), .S0(new_n401_), .Y(new_n402_));
  INVX1    g266(.A(new_n402_), .Y(new_n403_));
  AOI21X1  g267(.A0(new_n231_), .A1(new_n155_), .B0(new_n402_), .Y(new_n404_));
  OR2X1    g268(.A(\A[77] ), .B(\A[76] ), .Y(new_n405_));
  NOR2X1   g269(.A(new_n405_), .B(new_n400_), .Y(new_n406_));
  OR2X1    g270(.A(new_n406_), .B(new_n404_), .Y(new_n407_));
  NOR2X1   g271(.A(\A[75] ), .B(\A[74] ), .Y(new_n408_));
  MX2X1    g272(.A(new_n407_), .B(new_n403_), .S0(new_n408_), .Y(new_n409_));
  OAI21X1  g273(.A0(\A[73] ), .A1(\A[72] ), .B0(new_n409_), .Y(new_n410_));
  NAND3X1  g274(.A(new_n407_), .B(new_n237_), .C(new_n153_), .Y(new_n411_));
  AND2X1   g275(.A(new_n411_), .B(new_n410_), .Y(new_n412_));
  INVX1    g276(.A(new_n412_), .Y(new_n413_));
  OR2X1    g277(.A(\A[71] ), .B(\A[70] ), .Y(new_n414_));
  NOR2X1   g278(.A(new_n414_), .B(new_n409_), .Y(new_n415_));
  AOI21X1  g279(.A0(new_n414_), .A1(new_n412_), .B0(new_n415_), .Y(new_n416_));
  NOR2X1   g280(.A(\A[69] ), .B(\A[68] ), .Y(new_n417_));
  MX2X1    g281(.A(new_n416_), .B(new_n413_), .S0(new_n417_), .Y(new_n418_));
  INVX1    g282(.A(new_n418_), .Y(new_n419_));
  AOI21X1  g283(.A0(new_n244_), .A1(new_n152_), .B0(new_n418_), .Y(new_n420_));
  NOR3X1   g284(.A(new_n416_), .B(\A[67] ), .C(\A[66] ), .Y(new_n421_));
  OR2X1    g285(.A(new_n421_), .B(new_n420_), .Y(new_n422_));
  NOR2X1   g286(.A(\A[65] ), .B(\A[64] ), .Y(new_n423_));
  MX2X1    g287(.A(new_n422_), .B(new_n419_), .S0(new_n423_), .Y(new_n424_));
  OAI21X1  g288(.A0(\A[63] ), .A1(\A[62] ), .B0(new_n424_), .Y(new_n425_));
  NAND3X1  g289(.A(new_n422_), .B(new_n250_), .C(new_n150_), .Y(new_n426_));
  AND2X1   g290(.A(new_n426_), .B(new_n425_), .Y(new_n427_));
  INVX1    g291(.A(new_n427_), .Y(new_n428_));
  OR2X1    g292(.A(\A[61] ), .B(\A[60] ), .Y(new_n429_));
  NOR2X1   g293(.A(new_n429_), .B(new_n424_), .Y(new_n430_));
  AOI21X1  g294(.A0(new_n429_), .A1(new_n427_), .B0(new_n430_), .Y(new_n431_));
  NOR2X1   g295(.A(\A[59] ), .B(\A[58] ), .Y(new_n432_));
  MX2X1    g296(.A(new_n431_), .B(new_n428_), .S0(new_n432_), .Y(new_n433_));
  INVX1    g297(.A(new_n433_), .Y(new_n434_));
  AOI21X1  g298(.A0(new_n257_), .A1(new_n149_), .B0(new_n433_), .Y(new_n435_));
  NOR3X1   g299(.A(new_n431_), .B(\A[57] ), .C(\A[56] ), .Y(new_n436_));
  OR2X1    g300(.A(new_n436_), .B(new_n435_), .Y(new_n437_));
  NOR2X1   g301(.A(\A[55] ), .B(\A[54] ), .Y(new_n438_));
  MX2X1    g302(.A(new_n437_), .B(new_n434_), .S0(new_n438_), .Y(new_n439_));
  OAI21X1  g303(.A0(\A[53] ), .A1(\A[52] ), .B0(new_n439_), .Y(new_n440_));
  NAND3X1  g304(.A(new_n437_), .B(new_n263_), .C(new_n147_), .Y(new_n441_));
  AND2X1   g305(.A(new_n441_), .B(new_n440_), .Y(new_n442_));
  INVX1    g306(.A(new_n442_), .Y(new_n443_));
  OR2X1    g307(.A(\A[51] ), .B(\A[50] ), .Y(new_n444_));
  NOR2X1   g308(.A(new_n444_), .B(new_n439_), .Y(new_n445_));
  AOI21X1  g309(.A0(new_n444_), .A1(new_n442_), .B0(new_n445_), .Y(new_n446_));
  NOR2X1   g310(.A(\A[49] ), .B(\A[48] ), .Y(new_n447_));
  MX2X1    g311(.A(new_n446_), .B(new_n443_), .S0(new_n447_), .Y(new_n448_));
  INVX1    g312(.A(new_n448_), .Y(new_n449_));
  AOI21X1  g313(.A0(new_n270_), .A1(new_n146_), .B0(new_n448_), .Y(new_n450_));
  NOR3X1   g314(.A(new_n446_), .B(\A[47] ), .C(\A[46] ), .Y(new_n451_));
  OR2X1    g315(.A(new_n451_), .B(new_n450_), .Y(new_n452_));
  NOR2X1   g316(.A(\A[45] ), .B(\A[44] ), .Y(new_n453_));
  MX2X1    g317(.A(new_n452_), .B(new_n449_), .S0(new_n453_), .Y(new_n454_));
  OAI21X1  g318(.A0(\A[43] ), .A1(\A[42] ), .B0(new_n454_), .Y(new_n455_));
  NAND3X1  g319(.A(new_n452_), .B(new_n276_), .C(new_n144_), .Y(new_n456_));
  AND2X1   g320(.A(new_n456_), .B(new_n455_), .Y(new_n457_));
  INVX1    g321(.A(new_n457_), .Y(new_n458_));
  OR2X1    g322(.A(\A[41] ), .B(\A[40] ), .Y(new_n459_));
  NOR2X1   g323(.A(new_n459_), .B(new_n454_), .Y(new_n460_));
  AOI21X1  g324(.A0(new_n459_), .A1(new_n457_), .B0(new_n460_), .Y(new_n461_));
  NOR2X1   g325(.A(\A[39] ), .B(\A[38] ), .Y(new_n462_));
  MX2X1    g326(.A(new_n461_), .B(new_n458_), .S0(new_n462_), .Y(new_n463_));
  INVX1    g327(.A(new_n463_), .Y(new_n464_));
  AOI21X1  g328(.A0(new_n283_), .A1(new_n143_), .B0(new_n463_), .Y(new_n465_));
  NOR3X1   g329(.A(new_n461_), .B(\A[37] ), .C(\A[36] ), .Y(new_n466_));
  OR2X1    g330(.A(new_n466_), .B(new_n465_), .Y(new_n467_));
  NOR2X1   g331(.A(\A[35] ), .B(\A[34] ), .Y(new_n468_));
  MX2X1    g332(.A(new_n467_), .B(new_n464_), .S0(new_n468_), .Y(new_n469_));
  OAI21X1  g333(.A0(\A[33] ), .A1(\A[32] ), .B0(new_n469_), .Y(new_n470_));
  NAND3X1  g334(.A(new_n467_), .B(new_n289_), .C(new_n141_), .Y(new_n471_));
  AND2X1   g335(.A(new_n471_), .B(new_n470_), .Y(new_n472_));
  INVX1    g336(.A(new_n472_), .Y(new_n473_));
  OR2X1    g337(.A(\A[31] ), .B(\A[30] ), .Y(new_n474_));
  NOR2X1   g338(.A(new_n474_), .B(new_n469_), .Y(new_n475_));
  AOI21X1  g339(.A0(new_n474_), .A1(new_n472_), .B0(new_n475_), .Y(new_n476_));
  NOR2X1   g340(.A(\A[29] ), .B(\A[28] ), .Y(new_n477_));
  MX2X1    g341(.A(new_n476_), .B(new_n473_), .S0(new_n477_), .Y(new_n478_));
  INVX1    g342(.A(new_n478_), .Y(new_n479_));
  AOI21X1  g343(.A0(new_n296_), .A1(new_n140_), .B0(new_n478_), .Y(new_n480_));
  NOR3X1   g344(.A(new_n476_), .B(\A[27] ), .C(\A[26] ), .Y(new_n481_));
  OR2X1    g345(.A(new_n481_), .B(new_n480_), .Y(new_n482_));
  NOR2X1   g346(.A(\A[25] ), .B(\A[24] ), .Y(new_n483_));
  MX2X1    g347(.A(new_n482_), .B(new_n479_), .S0(new_n483_), .Y(new_n484_));
  OAI21X1  g348(.A0(\A[23] ), .A1(\A[22] ), .B0(new_n484_), .Y(new_n485_));
  NAND3X1  g349(.A(new_n482_), .B(new_n302_), .C(new_n138_), .Y(new_n486_));
  AND2X1   g350(.A(new_n486_), .B(new_n485_), .Y(new_n487_));
  INVX1    g351(.A(new_n487_), .Y(new_n488_));
  OR2X1    g352(.A(\A[21] ), .B(\A[20] ), .Y(new_n489_));
  NOR2X1   g353(.A(new_n489_), .B(new_n484_), .Y(new_n490_));
  AOI21X1  g354(.A0(new_n489_), .A1(new_n487_), .B0(new_n490_), .Y(new_n491_));
  NOR2X1   g355(.A(\A[19] ), .B(\A[18] ), .Y(new_n492_));
  MX2X1    g356(.A(new_n491_), .B(new_n488_), .S0(new_n492_), .Y(new_n493_));
  NOR2X1   g357(.A(\A[17] ), .B(\A[16] ), .Y(new_n494_));
  NOR2X1   g358(.A(new_n494_), .B(new_n493_), .Y(new_n495_));
  NOR3X1   g359(.A(new_n491_), .B(\A[17] ), .C(\A[16] ), .Y(new_n496_));
  OR2X1    g360(.A(new_n496_), .B(new_n495_), .Y(new_n497_));
  INVX1    g361(.A(new_n497_), .Y(new_n498_));
  NOR2X1   g362(.A(\A[15] ), .B(\A[14] ), .Y(new_n499_));
  MX2X1    g363(.A(new_n498_), .B(new_n493_), .S0(new_n499_), .Y(new_n500_));
  NOR2X1   g364(.A(\A[13] ), .B(\A[12] ), .Y(new_n501_));
  MX2X1    g365(.A(new_n500_), .B(new_n498_), .S0(new_n501_), .Y(new_n502_));
  NOR2X1   g366(.A(\A[11] ), .B(\A[10] ), .Y(new_n503_));
  MX2X1    g367(.A(new_n502_), .B(new_n500_), .S0(new_n503_), .Y(new_n504_));
  NOR2X1   g368(.A(\A[9] ), .B(\A[8] ), .Y(new_n505_));
  MX2X1    g369(.A(new_n504_), .B(new_n502_), .S0(new_n505_), .Y(new_n506_));
  NOR2X1   g370(.A(\A[7] ), .B(\A[6] ), .Y(new_n507_));
  MX2X1    g371(.A(new_n506_), .B(new_n504_), .S0(new_n507_), .Y(new_n508_));
  NOR2X1   g372(.A(\A[5] ), .B(\A[4] ), .Y(new_n509_));
  OR2X1    g373(.A(new_n509_), .B(new_n508_), .Y(new_n510_));
  NOR2X1   g374(.A(\A[3] ), .B(\A[2] ), .Y(new_n511_));
  NOR3X1   g375(.A(new_n506_), .B(\A[5] ), .C(\A[4] ), .Y(new_n512_));
  NOR2X1   g376(.A(new_n511_), .B(new_n512_), .Y(new_n513_));
  AOI22X1  g377(.A0(new_n513_), .A1(new_n510_), .B0(new_n511_), .B1(new_n508_), .Y(\P[1] ));
  NOR4X1   g378(.A(\A[127] ), .B(\A[126] ), .C(\A[125] ), .D(\A[124] ), .Y(new_n515_));
  INVX1    g379(.A(new_n515_), .Y(new_n516_));
  NOR4X1   g380(.A(\A[123] ), .B(\A[122] ), .C(\A[121] ), .D(\A[120] ), .Y(new_n517_));
  NOR4X1   g381(.A(\A[119] ), .B(\A[118] ), .C(\A[117] ), .D(\A[116] ), .Y(new_n518_));
  INVX1    g382(.A(new_n518_), .Y(new_n519_));
  AOI21X1  g383(.A0(new_n519_), .A1(new_n517_), .B0(new_n516_), .Y(new_n520_));
  INVX1    g384(.A(new_n520_), .Y(new_n521_));
  NOR3X1   g385(.A(\A[114] ), .B(\A[113] ), .C(\A[112] ), .Y(new_n522_));
  INVX1    g386(.A(new_n517_), .Y(new_n523_));
  AOI21X1  g387(.A0(new_n518_), .A1(\A[115] ), .B0(new_n523_), .Y(new_n524_));
  AND2X1   g388(.A(new_n522_), .B(new_n515_), .Y(new_n525_));
  INVX1    g389(.A(new_n525_), .Y(new_n526_));
  OAI22X1  g390(.A0(new_n526_), .A1(new_n524_), .B0(new_n522_), .B1(new_n521_), .Y(new_n527_));
  NOR4X1   g391(.A(\A[111] ), .B(\A[110] ), .C(\A[109] ), .D(\A[108] ), .Y(new_n528_));
  MX2X1    g392(.A(new_n527_), .B(new_n520_), .S0(new_n528_), .Y(new_n529_));
  NOR4X1   g393(.A(\A[107] ), .B(\A[106] ), .C(\A[105] ), .D(\A[104] ), .Y(new_n530_));
  MX2X1    g394(.A(new_n529_), .B(new_n527_), .S0(new_n530_), .Y(new_n531_));
  NOR4X1   g395(.A(\A[103] ), .B(\A[102] ), .C(\A[101] ), .D(\A[100] ), .Y(new_n532_));
  MX2X1    g396(.A(new_n531_), .B(new_n529_), .S0(new_n532_), .Y(new_n533_));
  NOR4X1   g397(.A(\A[99] ), .B(\A[98] ), .C(\A[97] ), .D(\A[96] ), .Y(new_n534_));
  INVX1    g398(.A(new_n534_), .Y(new_n535_));
  MX2X1    g399(.A(new_n531_), .B(new_n533_), .S0(new_n535_), .Y(new_n536_));
  NOR4X1   g400(.A(\A[95] ), .B(\A[94] ), .C(\A[93] ), .D(\A[92] ), .Y(new_n537_));
  MX2X1    g401(.A(new_n536_), .B(new_n533_), .S0(new_n537_), .Y(new_n538_));
  NOR4X1   g402(.A(\A[91] ), .B(\A[90] ), .C(\A[89] ), .D(\A[88] ), .Y(new_n539_));
  MX2X1    g403(.A(new_n538_), .B(new_n536_), .S0(new_n539_), .Y(new_n540_));
  NOR4X1   g404(.A(\A[87] ), .B(\A[86] ), .C(\A[85] ), .D(\A[84] ), .Y(new_n541_));
  MX2X1    g405(.A(new_n540_), .B(new_n538_), .S0(new_n541_), .Y(new_n542_));
  NOR4X1   g406(.A(\A[83] ), .B(\A[82] ), .C(\A[81] ), .D(\A[80] ), .Y(new_n543_));
  MX2X1    g407(.A(new_n542_), .B(new_n540_), .S0(new_n543_), .Y(new_n544_));
  NOR4X1   g408(.A(\A[79] ), .B(\A[78] ), .C(\A[77] ), .D(\A[76] ), .Y(new_n545_));
  MX2X1    g409(.A(new_n544_), .B(new_n542_), .S0(new_n545_), .Y(new_n546_));
  NOR4X1   g410(.A(\A[75] ), .B(\A[74] ), .C(\A[73] ), .D(\A[72] ), .Y(new_n547_));
  MX2X1    g411(.A(new_n546_), .B(new_n544_), .S0(new_n547_), .Y(new_n548_));
  NOR4X1   g412(.A(\A[71] ), .B(\A[70] ), .C(\A[69] ), .D(\A[68] ), .Y(new_n549_));
  MX2X1    g413(.A(new_n548_), .B(new_n546_), .S0(new_n549_), .Y(new_n550_));
  NOR4X1   g414(.A(\A[67] ), .B(\A[66] ), .C(\A[65] ), .D(\A[64] ), .Y(new_n551_));
  MX2X1    g415(.A(new_n550_), .B(new_n548_), .S0(new_n551_), .Y(new_n552_));
  NOR4X1   g416(.A(\A[63] ), .B(\A[62] ), .C(\A[61] ), .D(\A[60] ), .Y(new_n553_));
  MX2X1    g417(.A(new_n552_), .B(new_n550_), .S0(new_n553_), .Y(new_n554_));
  NOR4X1   g418(.A(\A[59] ), .B(\A[58] ), .C(\A[57] ), .D(\A[56] ), .Y(new_n555_));
  MX2X1    g419(.A(new_n554_), .B(new_n552_), .S0(new_n555_), .Y(new_n556_));
  NOR4X1   g420(.A(\A[55] ), .B(\A[54] ), .C(\A[53] ), .D(\A[52] ), .Y(new_n557_));
  MX2X1    g421(.A(new_n556_), .B(new_n554_), .S0(new_n557_), .Y(new_n558_));
  NOR4X1   g422(.A(\A[51] ), .B(\A[50] ), .C(\A[49] ), .D(\A[48] ), .Y(new_n559_));
  MX2X1    g423(.A(new_n558_), .B(new_n556_), .S0(new_n559_), .Y(new_n560_));
  NOR4X1   g424(.A(\A[47] ), .B(\A[46] ), .C(\A[45] ), .D(\A[44] ), .Y(new_n561_));
  MX2X1    g425(.A(new_n560_), .B(new_n558_), .S0(new_n561_), .Y(new_n562_));
  NOR4X1   g426(.A(\A[43] ), .B(\A[42] ), .C(\A[41] ), .D(\A[40] ), .Y(new_n563_));
  MX2X1    g427(.A(new_n562_), .B(new_n560_), .S0(new_n563_), .Y(new_n564_));
  NOR4X1   g428(.A(\A[39] ), .B(\A[38] ), .C(\A[37] ), .D(\A[36] ), .Y(new_n565_));
  MX2X1    g429(.A(new_n564_), .B(new_n562_), .S0(new_n565_), .Y(new_n566_));
  NOR4X1   g430(.A(\A[35] ), .B(\A[34] ), .C(\A[33] ), .D(\A[32] ), .Y(new_n567_));
  MX2X1    g431(.A(new_n566_), .B(new_n564_), .S0(new_n567_), .Y(new_n568_));
  NOR4X1   g432(.A(\A[31] ), .B(\A[30] ), .C(\A[29] ), .D(\A[28] ), .Y(new_n569_));
  MX2X1    g433(.A(new_n568_), .B(new_n566_), .S0(new_n569_), .Y(new_n570_));
  NOR4X1   g434(.A(\A[27] ), .B(\A[26] ), .C(\A[25] ), .D(\A[24] ), .Y(new_n571_));
  MX2X1    g435(.A(new_n570_), .B(new_n568_), .S0(new_n571_), .Y(new_n572_));
  NOR4X1   g436(.A(\A[23] ), .B(\A[22] ), .C(\A[21] ), .D(\A[20] ), .Y(new_n573_));
  MX2X1    g437(.A(new_n572_), .B(new_n570_), .S0(new_n573_), .Y(new_n574_));
  NOR4X1   g438(.A(\A[19] ), .B(\A[18] ), .C(\A[17] ), .D(\A[16] ), .Y(new_n575_));
  MX2X1    g439(.A(new_n574_), .B(new_n572_), .S0(new_n575_), .Y(new_n576_));
  NOR4X1   g440(.A(\A[15] ), .B(\A[14] ), .C(\A[13] ), .D(\A[12] ), .Y(new_n577_));
  MX2X1    g441(.A(new_n576_), .B(new_n574_), .S0(new_n577_), .Y(new_n578_));
  NOR4X1   g442(.A(\A[11] ), .B(\A[10] ), .C(\A[9] ), .D(\A[8] ), .Y(new_n579_));
  INVX1    g443(.A(new_n579_), .Y(new_n580_));
  AND2X1   g444(.A(new_n580_), .B(new_n578_), .Y(new_n581_));
  NOR4X1   g445(.A(\A[7] ), .B(\A[6] ), .C(\A[5] ), .D(\A[4] ), .Y(new_n582_));
  INVX1    g446(.A(new_n582_), .Y(new_n583_));
  AND2X1   g447(.A(new_n579_), .B(new_n576_), .Y(new_n584_));
  OR2X1    g448(.A(new_n582_), .B(new_n584_), .Y(new_n585_));
  OAI22X1  g449(.A0(new_n585_), .A1(new_n581_), .B0(new_n583_), .B1(new_n578_), .Y(\P[2] ));
  AND2X1   g450(.A(new_n517_), .B(new_n515_), .Y(new_n587_));
  NAND3X1  g451(.A(new_n518_), .B(new_n346_), .C(new_n344_), .Y(new_n588_));
  AND2X1   g452(.A(new_n530_), .B(new_n528_), .Y(new_n589_));
  OR2X1    g453(.A(new_n589_), .B(new_n588_), .Y(new_n590_));
  AND2X1   g454(.A(new_n590_), .B(new_n587_), .Y(new_n591_));
  NOR4X1   g455(.A(new_n373_), .B(new_n370_), .C(new_n368_), .D(\A[102] ), .Y(new_n592_));
  INVX1    g456(.A(new_n592_), .Y(new_n593_));
  AOI21X1  g457(.A0(new_n589_), .A1(\A[103] ), .B0(new_n588_), .Y(new_n594_));
  INVX1    g458(.A(new_n594_), .Y(new_n595_));
  AND2X1   g459(.A(new_n592_), .B(new_n587_), .Y(new_n596_));
  AOI22X1  g460(.A0(new_n596_), .A1(new_n595_), .B0(new_n593_), .B1(new_n591_), .Y(new_n597_));
  INVX1    g461(.A(new_n597_), .Y(new_n598_));
  AND2X1   g462(.A(new_n539_), .B(new_n537_), .Y(new_n599_));
  MX2X1    g463(.A(new_n598_), .B(new_n591_), .S0(new_n599_), .Y(new_n600_));
  INVX1    g464(.A(new_n600_), .Y(new_n601_));
  AND2X1   g465(.A(new_n543_), .B(new_n541_), .Y(new_n602_));
  MX2X1    g466(.A(new_n601_), .B(new_n597_), .S0(new_n602_), .Y(new_n603_));
  INVX1    g467(.A(new_n603_), .Y(new_n604_));
  AND2X1   g468(.A(new_n547_), .B(new_n545_), .Y(new_n605_));
  MX2X1    g469(.A(new_n604_), .B(new_n600_), .S0(new_n605_), .Y(new_n606_));
  INVX1    g470(.A(new_n606_), .Y(new_n607_));
  AND2X1   g471(.A(new_n551_), .B(new_n549_), .Y(new_n608_));
  MX2X1    g472(.A(new_n607_), .B(new_n603_), .S0(new_n608_), .Y(new_n609_));
  INVX1    g473(.A(new_n609_), .Y(new_n610_));
  AND2X1   g474(.A(new_n555_), .B(new_n553_), .Y(new_n611_));
  MX2X1    g475(.A(new_n610_), .B(new_n606_), .S0(new_n611_), .Y(new_n612_));
  INVX1    g476(.A(new_n612_), .Y(new_n613_));
  AND2X1   g477(.A(new_n559_), .B(new_n557_), .Y(new_n614_));
  MX2X1    g478(.A(new_n613_), .B(new_n609_), .S0(new_n614_), .Y(new_n615_));
  INVX1    g479(.A(new_n615_), .Y(new_n616_));
  AND2X1   g480(.A(new_n563_), .B(new_n561_), .Y(new_n617_));
  MX2X1    g481(.A(new_n616_), .B(new_n612_), .S0(new_n617_), .Y(new_n618_));
  INVX1    g482(.A(new_n618_), .Y(new_n619_));
  AND2X1   g483(.A(new_n567_), .B(new_n565_), .Y(new_n620_));
  MX2X1    g484(.A(new_n619_), .B(new_n615_), .S0(new_n620_), .Y(new_n621_));
  AND2X1   g485(.A(new_n571_), .B(new_n569_), .Y(new_n622_));
  MX2X1    g486(.A(new_n621_), .B(new_n619_), .S0(new_n622_), .Y(new_n623_));
  AND2X1   g487(.A(new_n575_), .B(new_n573_), .Y(new_n624_));
  NOR2X1   g488(.A(new_n624_), .B(new_n623_), .Y(new_n625_));
  INVX1    g489(.A(new_n624_), .Y(new_n626_));
  NAND2X1  g490(.A(new_n579_), .B(new_n577_), .Y(new_n627_));
  OAI21X1  g491(.A0(new_n626_), .A1(new_n621_), .B0(new_n627_), .Y(new_n628_));
  NAND3X1  g492(.A(new_n623_), .B(new_n579_), .C(new_n577_), .Y(new_n629_));
  OAI21X1  g493(.A0(new_n628_), .A1(new_n625_), .B0(new_n629_), .Y(\P[3] ));
  INVX1    g494(.A(new_n587_), .Y(new_n631_));
  NAND4X1  g495(.A(new_n534_), .B(new_n532_), .C(new_n530_), .D(new_n528_), .Y(new_n632_));
  AOI21X1  g496(.A0(new_n602_), .A1(new_n599_), .B0(new_n632_), .Y(new_n633_));
  NOR3X1   g497(.A(new_n633_), .B(new_n588_), .C(new_n631_), .Y(new_n634_));
  INVX1    g498(.A(new_n547_), .Y(new_n635_));
  INVX1    g499(.A(new_n608_), .Y(new_n636_));
  NOR4X1   g500(.A(new_n636_), .B(new_n635_), .C(new_n405_), .D(\A[78] ), .Y(new_n637_));
  INVX1    g501(.A(new_n637_), .Y(new_n638_));
  AND2X1   g502(.A(new_n602_), .B(new_n599_), .Y(new_n639_));
  AOI21X1  g503(.A0(new_n639_), .A1(\A[79] ), .B0(new_n632_), .Y(new_n640_));
  NOR4X1   g504(.A(new_n640_), .B(new_n638_), .C(new_n588_), .D(new_n631_), .Y(new_n641_));
  AOI21X1  g505(.A0(new_n638_), .A1(new_n634_), .B0(new_n641_), .Y(new_n642_));
  INVX1    g506(.A(new_n642_), .Y(new_n643_));
  AND2X1   g507(.A(new_n614_), .B(new_n611_), .Y(new_n644_));
  MX2X1    g508(.A(new_n643_), .B(new_n634_), .S0(new_n644_), .Y(new_n645_));
  AND2X1   g509(.A(new_n624_), .B(new_n622_), .Y(new_n646_));
  INVX1    g510(.A(new_n646_), .Y(new_n647_));
  INVX1    g511(.A(new_n645_), .Y(new_n648_));
  AND2X1   g512(.A(new_n620_), .B(new_n617_), .Y(new_n649_));
  AOI21X1  g513(.A0(new_n649_), .A1(new_n643_), .B0(new_n646_), .Y(new_n650_));
  OAI21X1  g514(.A0(new_n649_), .A1(new_n648_), .B0(new_n650_), .Y(new_n651_));
  OAI21X1  g515(.A0(new_n647_), .A1(new_n645_), .B0(new_n651_), .Y(\P[4] ));
  NOR4X1   g516(.A(new_n632_), .B(new_n588_), .C(new_n523_), .D(new_n516_), .Y(new_n653_));
  NAND4X1  g517(.A(new_n608_), .B(new_n605_), .C(new_n602_), .D(new_n599_), .Y(new_n654_));
  AND2X1   g518(.A(new_n649_), .B(new_n644_), .Y(new_n655_));
  OAI21X1  g519(.A0(new_n655_), .A1(new_n654_), .B0(new_n653_), .Y(\P[5] ));
  NOR4X1   g520(.A(new_n654_), .B(new_n632_), .C(new_n588_), .D(new_n631_), .Y(new_n657_));
  INVX1    g521(.A(new_n657_), .Y(\P[6] ));
  OR4X1    g522(.A(\A[3] ), .B(\A[2] ), .C(\A[1] ), .D(\A[0] ), .Y(new_n659_));
  NOR3X1   g523(.A(new_n659_), .B(new_n627_), .C(new_n583_), .Y(new_n660_));
  NAND4X1  g524(.A(new_n660_), .B(new_n657_), .C(new_n655_), .D(new_n646_), .Y(F));
endmodule


