//Converted to Combinational (Partial output: n177) , Module name: s713_n177
module s713_n177 ( G5, G2, G75, G3, G77, G76, G64, G72, G65, G13, G9, G10, G22, G11, G66, G78, G24, G23, G71, G67, G4, G25, n177 );
input G5, G2, G75, G3, G77, G76, G64, G72, G65, G13, G9, G10, G22, G11, G66, G78, G24, G23, G71, G67, G4, G25;
output n177;
wire n216, n117, n215, n147_1, n126, n116, n115, G86BF, n214, n117_1, n133, n139, n143, n134, n140, n151, n213, n128, n132_1, n138, n141, n142_1, n125, n203, n127_1, n118, n124, n130, n131, n137_1, n135, n122_1, n172_1, n120, n123, n129, n136, n165, n119, n121;
OAI21X1  g102(.A0(n215), .A1(n117), .B0(n216), .Y(n177));
OAI21X1  g101(.A0(G5), .A1(n126), .B0(n147_1), .Y(n216));
AOI21X1  g030(.A0(G86BF), .A1(n115), .B0(n116), .Y(n117));
OAI21X1  g100(.A0(n133), .A1(n117_1), .B0(n214), .Y(n215));
INVX1    g032(.A(n139), .Y(n147_1));
INVX1    g011(.A(G2), .Y(n126));
INVX1    g001(.A(G75), .Y(n116));
INVX1    g000(.A(G3), .Y(n115));
OAI21X1  g029(.A0(n140), .A1(n134), .B0(n143), .Y(G86BF));
NOR2X1   g099(.A(n213), .B(n151), .Y(n214));
INVX1    g002(.A(G77), .Y(n117_1));
AOI21X1  g018(.A0(n132_1), .A1(n128), .B0(G3), .Y(n133));
OAI21X1  g024(.A0(n138), .A1(G3), .B0(G76), .Y(n139));
NOR2X1   g028(.A(n142_1), .B(n141), .Y(n143));
OAI21X1  g019(.A0(n133), .A1(n117_1), .B0(n125), .Y(n134));
NAND3X1  g025(.A(n139), .B(G64), .C(n126), .Y(n140));
INVX1    g036(.A(n125), .Y(n151));
NAND4X1  g098(.A(n138), .B(G72), .C(G5), .D(n203), .Y(n213));
OAI21X1  g013(.A0(n124), .A1(n118), .B0(n127_1), .Y(n128));
NOR2X1   g017(.A(n131), .B(n130), .Y(n132_1));
NOR4X1   g023(.A(n122_1), .B(G65), .C(n135), .D(n137_1), .Y(n138));
NOR4X1   g026(.A(G10), .B(G9), .C(G3), .D(G13), .Y(n141));
OAI21X1  g027(.A0(G11), .A1(G3), .B0(G22), .Y(n142_1));
OR2X1    g010(.A(n124), .B(n118), .Y(n125));
INVX1    g088(.A(n172_1), .Y(n203));
AND2X1   g012(.A(G66), .B(n126), .Y(n127_1));
INVX1    g003(.A(G78), .Y(n118));
AOI21X1  g009(.A0(n123), .A1(n120), .B0(G3), .Y(n124));
NOR4X1   g015(.A(G10), .B(n129), .C(G3), .D(G13), .Y(n130));
OAI21X1  g016(.A0(G11), .A1(G3), .B0(G24), .Y(n131));
NOR4X1   g022(.A(n136), .B(G9), .C(G3), .D(G13), .Y(n137_1));
INVX1    g020(.A(G23), .Y(n135));
NOR2X1   g007(.A(G11), .B(G3), .Y(n122_1));
NAND2X1  g057(.A(G71), .B(n165), .Y(n172_1));
NAND4X1  g005(.A(G10), .B(G9), .C(n115), .D(n119), .Y(n120));
NOR3X1   g008(.A(n122_1), .B(G67), .C(n121), .Y(n123));
INVX1    g014(.A(G9), .Y(n129));
INVX1    g021(.A(G10), .Y(n136));
INVX1    g050(.A(G4), .Y(n165));
INVX1    g004(.A(G13), .Y(n119));
INVX1    g006(.A(G25), .Y(n121));

endmodule
