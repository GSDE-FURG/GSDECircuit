//Converted to Combinational (Partial output: n1722) , Module name: s38417_n1722 , Timestamp: 2018-12-03T15:51:12.371353 
module s38417_n1722 ( g404, g405, g309, g403, g402, g181, g276, g401, g121, g169, g168, g170, g113, g109, g117, g97, g125, g157, g156, g158, g105, g101, g154, g153, g155, g172, g171, g173, g163, g162, g164, g138, g165, g135, g175, g174, g176, g160, g159, g161, g148, g147, g149, g145, g144, g146, g151, g150, g152, g130, g129, g131, g142, g141, g143, g133, g132, g134, n1722 );
input g404, g405, g309, g403, g402, g181, g276, g401, g121, g169, g168, g170, g113, g109, g117, g97, g125, g157, g156, g158, g105, g101, g154, g153, g155, g172, g171, g173, g163, g162, g164, g138, g165, g135, g175, g174, g176, g160, g159, g161, g148, g147, g149, g145, g144, g146, g151, g150, g152, g130, g129, g131, g142, g141, g143, g133, g132, g134;
output n1722;
wire n5923, n5920, n5569_1, n5437_1, n5454, n5468, n5567, n5568, n5436, n5425, n5428, n5432, n5453, n5441, n5445, n5449, n5467, n5455_1, n5459, n5463, n5545, n5548, n5547, n1741, n5435, n5393, n5424_1, n5426, n5427, n5387, n5431, n5452, n1759, n5440, n1768, n5444, n1750, n5448, n1795, n5466, n1732, n5450, n5451_1, n1777, n5458, n1786, n5462, n5433_1, n5434, n5391, n5392_1, n5422, n5423, n5382, n5385, n5384, n5383_1, n5386, n5429_1, n5430, n5438, n5439, n5442_1, n5443, n5446_1, n5447, n5464_1, n5465, n5456, n5457, n5460_1, n5461;
MX2X1    g0881(.A(g404), .B(n5920), .S0(n5923), .Y(n1722));
AND2X1   g0880(.A(g309), .B(g405), .Y(n5923));
NAND4X1  g0877(.A(n5468), .B(n5454), .C(n5437_1), .D(n5569_1), .Y(n5920));
NOR2X1   g0527(.A(n5568), .B(n5567), .Y(n5569_1));
NOR4X1   g0395(.A(n5432), .B(n5428), .C(n5425), .D(n5436), .Y(n5437_1));
NOR4X1   g0412(.A(n5449), .B(n5445), .C(n5441), .D(n5453), .Y(n5454));
NOR4X1   g0426(.A(n5463), .B(n5459), .C(n5455_1), .D(n5467), .Y(n5468));
NOR2X1   g0525(.A(g403), .B(n5545), .Y(n5567));
OAI22X1  g0526(.A0(g404), .A1(n5547), .B0(n5548), .B1(g402), .Y(n5568));
XOR2X1   g0394(.A(n5435), .B(n1741), .Y(n5436));
AND2X1   g0383(.A(n5424_1), .B(n5393), .Y(n5425));
OAI21X1  g0386(.A0(n5427), .A1(n5426), .B0(g181), .Y(n5428));
XOR2X1   g0390(.A(n5431), .B(n5387), .Y(n5432));
OAI21X1  g0411(.A0(n5424_1), .A1(n5393), .B0(n5452), .Y(n5453));
XOR2X1   g0399(.A(n5440), .B(n1759), .Y(n5441));
XOR2X1   g0403(.A(n5444), .B(n1768), .Y(n5445));
XOR2X1   g0407(.A(n5448), .B(n1750), .Y(n5449));
XOR2X1   g0425(.A(n5466), .B(n1795), .Y(n5467));
NOR3X1   g0413(.A(n5451_1), .B(n5450), .C(n1732), .Y(n5455_1));
XOR2X1   g0417(.A(n5458), .B(n1777), .Y(n5459));
XOR2X1   g0421(.A(n5462), .B(n1786), .Y(n5463));
INVX1    g0503(.A(g276), .Y(n5545));
INVX1    g0506(.A(g401), .Y(n5548));
INVX1    g0505(.A(g405), .Y(n5547));
INVX1    g0332(.A(g121), .Y(n1741));
NOR2X1   g0393(.A(n5434), .B(n5433_1), .Y(n5435));
NOR2X1   g0351(.A(n5392_1), .B(n5391), .Y(n5393));
OR2X1    g0382(.A(n5423), .B(n5422), .Y(n5424_1));
NOR2X1   g0384(.A(g169), .B(n5382), .Y(n5426));
OAI22X1  g0385(.A0(g170), .A1(n5384), .B0(n5385), .B1(g168), .Y(n5427));
NOR2X1   g0345(.A(n5386), .B(n5383_1), .Y(n5387));
NOR2X1   g0389(.A(n5430), .B(n5429_1), .Y(n5431));
OAI21X1  g0410(.A0(n5451_1), .A1(n5450), .B0(n1732), .Y(n5452));
INVX1    g0324(.A(g113), .Y(n1759));
NOR2X1   g0398(.A(n5439), .B(n5438), .Y(n5440));
INVX1    g0320(.A(g109), .Y(n1768));
NOR2X1   g0402(.A(n5443), .B(n5442_1), .Y(n5444));
INVX1    g0328(.A(g117), .Y(n1750));
NOR2X1   g0406(.A(n5447), .B(n5446_1), .Y(n5448));
INVX1    g0305(.A(g97), .Y(n1795));
NOR2X1   g0424(.A(n5465), .B(n5464_1), .Y(n5466));
INVX1    g0336(.A(g125), .Y(n1732));
NOR2X1   g0408(.A(g157), .B(n5382), .Y(n5450));
OAI22X1  g0409(.A0(g158), .A1(n5384), .B0(n5385), .B1(g156), .Y(n5451_1));
INVX1    g0316(.A(g105), .Y(n1777));
NOR2X1   g0416(.A(n5457), .B(n5456), .Y(n5458));
INVX1    g0312(.A(g101), .Y(n1786));
NOR2X1   g0420(.A(n5461), .B(n5460_1), .Y(n5462));
NOR2X1   g0391(.A(g154), .B(n5382), .Y(n5433_1));
OAI22X1  g0392(.A0(g155), .A1(n5384), .B0(n5385), .B1(g153), .Y(n5434));
NOR2X1   g0349(.A(g172), .B(n5382), .Y(n5391));
OAI22X1  g0350(.A0(g173), .A1(n5384), .B0(n5385), .B1(g171), .Y(n5392_1));
NOR2X1   g0380(.A(g163), .B(n5382), .Y(n5422));
OAI22X1  g0381(.A0(g164), .A1(n5384), .B0(n5385), .B1(g162), .Y(n5423));
INVX1    g0340(.A(g138), .Y(n5382));
INVX1    g0343(.A(g165), .Y(n5385));
INVX1    g0342(.A(g135), .Y(n5384));
NOR2X1   g0341(.A(g175), .B(n5382), .Y(n5383_1));
OAI22X1  g0344(.A0(g176), .A1(n5384), .B0(n5385), .B1(g174), .Y(n5386));
NOR2X1   g0387(.A(g160), .B(n5382), .Y(n5429_1));
OAI22X1  g0388(.A0(g161), .A1(n5384), .B0(n5385), .B1(g159), .Y(n5430));
NOR2X1   g0396(.A(g148), .B(n5382), .Y(n5438));
OAI22X1  g0397(.A0(g149), .A1(n5384), .B0(n5385), .B1(g147), .Y(n5439));
NOR2X1   g0400(.A(g145), .B(n5382), .Y(n5442_1));
OAI22X1  g0401(.A0(g146), .A1(n5384), .B0(n5385), .B1(g144), .Y(n5443));
NOR2X1   g0404(.A(g151), .B(n5382), .Y(n5446_1));
OAI22X1  g0405(.A0(g152), .A1(n5384), .B0(n5385), .B1(g150), .Y(n5447));
NOR2X1   g0422(.A(g130), .B(n5382), .Y(n5464_1));
OAI22X1  g0423(.A0(g131), .A1(n5384), .B0(n5385), .B1(g129), .Y(n5465));
NOR2X1   g0414(.A(g142), .B(n5382), .Y(n5456));
OAI22X1  g0415(.A0(g143), .A1(n5384), .B0(n5385), .B1(g141), .Y(n5457));
NOR2X1   g0418(.A(g133), .B(n5382), .Y(n5460_1));
OAI22X1  g0419(.A0(g134), .A1(n5384), .B0(n5385), .B1(g132), .Y(n5461));

endmodule
