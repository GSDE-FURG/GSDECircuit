//Converted to Combinational (Partial output: n1005) , Module name: s38584_n1005 , Timestamp: 2018-12-03T15:51:16.093154 
module s38584_n1005 ( g35, g6199, g12, g9, g19, g28, g7, g31, g8, g16, g56, g57, g53, g34, g54, g2844, g2907, g2902, g956, g1300, g4727, g3853, g4917, g45, g2848, g776, g632, g538, g595, g947, g1291, n1005 );
input g6, g35, g6199, g12, g9, g19, g28, g7, g31, g8, g16, g56, g57, g53, g34, g54, g2844, g2907, g2902, g956, g1300, g4727, g3853, g4917, g45, g2848, g776, g632, g538, g595, g947, g1291;
output n1005;
wire n6030, n6029, n3747, n5616, n5019, n4988_1, n5221_1, n5234, n5248, n4982, n4983, n4979_1, n4383, n5072, n5220, n5040, n5233, n5247, n5236_1, n5239, n5242, n4977, n4976, n5003, n5014, n5215, n5218, n5219, n4987, n5029, n5232, n5224, n5227, n5230, n5246_1, n5067, n5017_1, n5244, n5235, n5031, n5238, n5237, n4991, n5241_1, n5240, n5062, n5002_1, n4998, n4999, n5000, n5013, n5007_1, n5010, n5012_1, n5216_1, n5217, n5025, n5026, n5028, n5023, n5231_1, n5223, n5222, n5225, n5226_1, n5229, n5228, n5245, n5024, n5008, n4984_1, n5016, n5243, n5005, n5048, n4990, n5050, n4981, n4995, n5001, n4997_1, n5009, n5004, n5006, n5011, n4996, n5021, n5027_1, n5022_1, n4989, n4980, n4994, n4992_1, n4993;
AND2X1   g1391(.A(n6030), .B(g35), .Y(n1005));
MX2X1    g1390(.A(g6199), .B(n3747), .S0(n6029), .Y(n6030));
NOR3X1   g1389(.A(n4988_1), .B(n5019), .C(n5616), .Y(n6029));
NAND3X1  g0827(.A(n5248), .B(n5234), .C(n5221_1), .Y(n3747));
INVX1    g0976(.A(g12), .Y(n5616));
NAND2X1  g0399(.A(n4983), .B(n4982), .Y(n5019));
NAND3X1  g0368(.A(g19), .B(g9), .C(n4979_1), .Y(n4988_1));
NAND3X1  g0581(.A(n5220), .B(n5072), .C(n4383), .Y(n5221_1));
NAND2X1  g0594(.A(n5233), .B(n5040), .Y(n5234));
NOR4X1   g0608(.A(n5242), .B(n5239), .C(n5236_1), .D(n5247), .Y(n5248));
INVX1    g0362(.A(g28), .Y(n4982));
NOR4X1   g0363(.A(g8), .B(g6), .C(g31), .D(g7), .Y(n4983));
INVX1    g0359(.A(g16), .Y(n4979_1));
NOR4X1   g0358(.A(n4976), .B(g57), .C(g56), .D(n4977), .Y(n4383));
OR2X1    g0447(.A(n5014), .B(n5003), .Y(n5072));
NAND3X1  g0580(.A(n5219), .B(n5218), .C(n5215), .Y(n5220));
NOR2X1   g0420(.A(n5029), .B(n4987), .Y(n5040));
OR4X1    g0593(.A(n5230), .B(n5227), .C(n5224), .D(n5232), .Y(n5233));
OAI22X1  g0607(.A0(n5244), .A1(n5017_1), .B0(n5067), .B1(n5246_1), .Y(n5247));
NOR4X1   g0596(.A(n5031), .B(n4987), .C(n5235), .D(n5019), .Y(n5236_1));
OAI21X1  g0599(.A0(n4991), .A1(n5237), .B0(n5238), .Y(n5239));
OAI21X1  g0602(.A0(n5062), .A1(n5240), .B0(n5241_1), .Y(n5242));
OR2X1    g0357(.A(g34), .B(g53), .Y(n4977));
INVX1    g0356(.A(g54), .Y(n4976));
OR4X1    g0383(.A(n5000), .B(n4999), .C(n4998), .D(n5002_1), .Y(n5003));
OR4X1    g0394(.A(n5012_1), .B(n5010), .C(n5007_1), .D(n5013), .Y(n5014));
NAND2X1  g0575(.A(n5010), .B(g2844), .Y(n5215));
OR2X1    g0578(.A(n5217), .B(n5216_1), .Y(n5218));
AOI22X1  g0579(.A0(n4998), .A1(g2902), .B0(g2907), .B1(n5000), .Y(n5219));
OR4X1    g0367(.A(n4976), .B(g57), .C(g56), .D(n4977), .Y(n4987));
NOR3X1   g0409(.A(n5028), .B(n5026), .C(n5025), .Y(n5029));
AOI21X1  g0592(.A0(n5231_1), .A1(g35), .B0(n5023), .Y(n5232));
AOI21X1  g0584(.A0(n5222), .A1(g35), .B0(n5223), .Y(n5224));
NOR2X1   g0587(.A(n5226_1), .B(n5225), .Y(n5227));
AOI21X1  g0590(.A0(n5228), .A1(g35), .B0(n5229), .Y(n5230));
NAND2X1  g0606(.A(n5245), .B(g956), .Y(n5246_1));
OR4X1    g0444(.A(n5008), .B(n4987), .C(n4982), .D(n5024), .Y(n5067));
NAND3X1  g0397(.A(n5016), .B(n4984_1), .C(n4383), .Y(n5017_1));
NAND2X1  g0604(.A(g1300), .B(n5243), .Y(n5244));
INVX1    g0595(.A(g4727), .Y(n5235));
NAND3X1  g0411(.A(g19), .B(n5005), .C(g16), .Y(n5031));
NAND4X1  g0598(.A(n4984_1), .B(n4383), .C(g6199), .D(n5048), .Y(n5238));
INVX1    g0597(.A(g3853), .Y(n5237));
OR4X1    g0371(.A(n4988_1), .B(n4987), .C(g28), .D(n4990), .Y(n4991));
NAND4X1  g0601(.A(n4981), .B(n4383), .C(g4917), .D(n5050), .Y(n5241_1));
INVX1    g0600(.A(g45), .Y(n5240));
OR2X1    g0442(.A(n4383), .B(g53), .Y(n5062));
NOR3X1   g0382(.A(n5001), .B(n4995), .C(g28), .Y(n5002_1));
NOR3X1   g0378(.A(n4997_1), .B(n4995), .C(g28), .Y(n4998));
NOR3X1   g0379(.A(n4995), .B(n4988_1), .C(n4982), .Y(n4999));
NOR3X1   g0380(.A(n4997_1), .B(n4995), .C(n4982), .Y(n5000));
NOR4X1   g0393(.A(n5008), .B(n4982), .C(n5005), .D(n5009), .Y(n5013));
NOR2X1   g0387(.A(n5006), .B(n5004), .Y(n5007_1));
NOR4X1   g0390(.A(n5008), .B(g28), .C(n5005), .D(n5009), .Y(n5010));
NOR2X1   g0392(.A(n5011), .B(n5006), .Y(n5012_1));
INVX1    g0576(.A(g2848), .Y(n5216_1));
NAND4X1  g0577(.A(n4983), .B(g28), .C(g9), .D(n4996), .Y(n5217));
OAI21X1  g0405(.A0(n5024), .A1(n5021), .B0(n5023), .Y(n5025));
NOR4X1   g0406(.A(n5008), .B(g28), .C(g9), .D(n5009), .Y(n5026));
OAI21X1  g0408(.A0(n5024), .A1(n5019), .B0(n5027_1), .Y(n5028));
NAND4X1  g0403(.A(n4989), .B(g28), .C(g31), .D(n5022_1), .Y(n5023));
INVX1    g0591(.A(g776), .Y(n5231_1));
OR2X1    g0583(.A(n5024), .B(n5019), .Y(n5223));
INVX1    g0582(.A(g632), .Y(n5222));
INVX1    g0585(.A(g538), .Y(n5225));
NAND3X1  g0586(.A(n5022_1), .B(n4983), .C(n4982), .Y(n5226_1));
OR2X1    g0589(.A(n5024), .B(n5021), .Y(n5229));
INVX1    g0588(.A(g595), .Y(n5228));
INVX1    g0605(.A(g947), .Y(n5245));
NAND3X1  g0404(.A(g19), .B(n5005), .C(n4979_1), .Y(n5024));
OR4X1    g0388(.A(g8), .B(g6), .C(g31), .D(g7), .Y(n5008));
AND2X1   g0364(.A(n4983), .B(n4982), .Y(n4984_1));
NOR3X1   g0396(.A(g19), .B(g9), .C(n4979_1), .Y(n5016));
INVX1    g0603(.A(g1291), .Y(n5243));
INVX1    g0385(.A(g9), .Y(n5005));
NOR3X1   g0428(.A(n4980), .B(n5005), .C(g16), .Y(n5048));
NAND2X1  g0370(.A(n4989), .B(g31), .Y(n4990));
AND2X1   g0430(.A(n4983), .B(g28), .Y(n5050));
NOR3X1   g0361(.A(n4980), .B(g9), .C(n4979_1), .Y(n4981));
OR4X1    g0375(.A(n4993), .B(n4992_1), .C(g31), .D(n4994), .Y(n4995));
NAND3X1  g0381(.A(n4980), .B(g9), .C(g16), .Y(n5001));
NAND2X1  g0377(.A(n4996), .B(g9), .Y(n4997_1));
OR2X1    g0389(.A(g19), .B(g16), .Y(n5009));
NAND2X1  g0384(.A(n4983), .B(g28), .Y(n5004));
NAND3X1  g0386(.A(n4980), .B(n5005), .C(g16), .Y(n5006));
NAND3X1  g0391(.A(n4989), .B(g28), .C(g31), .Y(n5011));
NOR2X1   g0376(.A(g19), .B(g16), .Y(n4996));
NAND3X1  g0401(.A(n4989), .B(n4982), .C(g31), .Y(n5021));
NAND3X1  g0407(.A(n5022_1), .B(n4983), .C(g28), .Y(n5027_1));
NOR3X1   g0402(.A(g19), .B(g9), .C(g16), .Y(n5022_1));
NOR3X1   g0369(.A(g7), .B(g8), .C(g6), .Y(n4989));
INVX1    g0360(.A(g19), .Y(n4980));
INVX1    g0374(.A(g7), .Y(n4994));
INVX1    g0372(.A(g6), .Y(n4992_1));
INVX1    g0373(.A(g8), .Y(n4993));

endmodule
