// Benchmark "top" written by ABC on Mon Sep 21 03:43:56 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ;
  output \asquared[0] , \asquared[1] , \asquared[2] , \asquared[3] ,
    \asquared[4] , \asquared[5] , \asquared[6] , \asquared[7] ,
    \asquared[8] , \asquared[9] , \asquared[10] , \asquared[11] ,
    \asquared[12] , \asquared[13] , \asquared[14] , \asquared[15] ,
    \asquared[16] , \asquared[17] , \asquared[18] , \asquared[19] ,
    \asquared[20] , \asquared[21] , \asquared[22] , \asquared[23] ,
    \asquared[24] , \asquared[25] , \asquared[26] , \asquared[27] ,
    \asquared[28] , \asquared[29] , \asquared[30] , \asquared[31] ,
    \asquared[32] , \asquared[33] , \asquared[34] , \asquared[35] ,
    \asquared[36] , \asquared[37] , \asquared[38] , \asquared[39] ,
    \asquared[40] , \asquared[41] , \asquared[42] , \asquared[43] ,
    \asquared[44] , \asquared[45] , \asquared[46] , \asquared[47] ,
    \asquared[48] , \asquared[49] , \asquared[50] , \asquared[51] ,
    \asquared[52] , \asquared[53] , \asquared[54] , \asquared[55] ,
    \asquared[56] , \asquared[57] , \asquared[58] , \asquared[59] ,
    \asquared[60] , \asquared[61] , \asquared[62] , \asquared[63] ,
    \asquared[64] , \asquared[65] , \asquared[66] , \asquared[67] ,
    \asquared[68] , \asquared[69] , \asquared[70] , \asquared[71] ,
    \asquared[72] , \asquared[73] , \asquared[74] , \asquared[75] ,
    \asquared[76] , \asquared[77] , \asquared[78] , \asquared[79] ,
    \asquared[80] , \asquared[81] , \asquared[82] , \asquared[83] ,
    \asquared[84] , \asquared[85] , \asquared[86] , \asquared[87] ,
    \asquared[88] , \asquared[89] , \asquared[90] , \asquared[91] ,
    \asquared[92] , \asquared[93] , \asquared[94] , \asquared[95] ,
    \asquared[96] , \asquared[97] , \asquared[98] , \asquared[99] ,
    \asquared[100] , \asquared[101] , \asquared[102] , \asquared[103] ,
    \asquared[104] , \asquared[105] , \asquared[106] , \asquared[107] ,
    \asquared[108] , \asquared[109] , \asquared[110] , \asquared[111] ,
    \asquared[112] , \asquared[113] , \asquared[114] , \asquared[115] ,
    \asquared[116] , \asquared[117] , \asquared[118] , \asquared[119] ,
    \asquared[120] , \asquared[121] , \asquared[122] , \asquared[123] ,
    \asquared[124] , \asquared[125] , \asquared[126] , \asquared[127] ;
  wire new_n194_, new_n196_, new_n197_, new_n198_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n216_, new_n217_, new_n218_, new_n219_, new_n220_, new_n221_,
    new_n222_, new_n223_, new_n224_, new_n225_, new_n226_, new_n227_,
    new_n228_, new_n230_, new_n231_, new_n232_, new_n233_, new_n234_,
    new_n235_, new_n236_, new_n237_, new_n238_, new_n239_, new_n240_,
    new_n241_, new_n242_, new_n243_, new_n244_, new_n245_, new_n246_,
    new_n248_, new_n249_, new_n250_, new_n251_, new_n252_, new_n253_,
    new_n254_, new_n255_, new_n256_, new_n257_, new_n258_, new_n259_,
    new_n260_, new_n261_, new_n262_, new_n263_, new_n264_, new_n265_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n361_, new_n362_, new_n363_, new_n364_, new_n365_,
    new_n366_, new_n367_, new_n368_, new_n369_, new_n370_, new_n371_,
    new_n372_, new_n373_, new_n374_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n392_, new_n393_, new_n394_, new_n395_, new_n396_,
    new_n397_, new_n398_, new_n399_, new_n400_, new_n401_, new_n402_,
    new_n403_, new_n404_, new_n405_, new_n406_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n414_,
    new_n415_, new_n416_, new_n417_, new_n418_, new_n419_, new_n420_,
    new_n421_, new_n422_, new_n423_, new_n424_, new_n425_, new_n426_,
    new_n427_, new_n428_, new_n430_, new_n431_, new_n432_, new_n433_,
    new_n434_, new_n435_, new_n436_, new_n437_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n443_, new_n444_, new_n445_,
    new_n446_, new_n447_, new_n448_, new_n449_, new_n450_, new_n451_,
    new_n452_, new_n453_, new_n454_, new_n455_, new_n456_, new_n457_,
    new_n458_, new_n459_, new_n460_, new_n461_, new_n462_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n610_, new_n611_,
    new_n612_, new_n613_, new_n614_, new_n615_, new_n616_, new_n617_,
    new_n618_, new_n619_, new_n620_, new_n621_, new_n622_, new_n623_,
    new_n624_, new_n625_, new_n626_, new_n627_, new_n628_, new_n629_,
    new_n630_, new_n631_, new_n632_, new_n633_, new_n634_, new_n635_,
    new_n636_, new_n637_, new_n638_, new_n639_, new_n640_, new_n641_,
    new_n642_, new_n643_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n673_, new_n674_, new_n675_, new_n676_, new_n677_, new_n678_,
    new_n679_, new_n680_, new_n681_, new_n682_, new_n683_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n702_,
    new_n703_, new_n704_, new_n705_, new_n706_, new_n707_, new_n708_,
    new_n709_, new_n710_, new_n711_, new_n712_, new_n713_, new_n714_,
    new_n715_, new_n716_, new_n717_, new_n718_, new_n719_, new_n720_,
    new_n721_, new_n722_, new_n723_, new_n724_, new_n725_, new_n726_,
    new_n727_, new_n728_, new_n729_, new_n731_, new_n732_, new_n733_,
    new_n734_, new_n735_, new_n736_, new_n737_, new_n738_, new_n739_,
    new_n740_, new_n741_, new_n742_, new_n743_, new_n744_, new_n745_,
    new_n746_, new_n747_, new_n748_, new_n749_, new_n750_, new_n751_,
    new_n752_, new_n753_, new_n754_, new_n755_, new_n756_, new_n757_,
    new_n758_, new_n759_, new_n760_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n770_, new_n771_, new_n772_, new_n773_, new_n774_, new_n775_,
    new_n776_, new_n777_, new_n778_, new_n779_, new_n780_, new_n781_,
    new_n782_, new_n783_, new_n784_, new_n785_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n986_, new_n987_, new_n988_, new_n989_,
    new_n990_, new_n991_, new_n992_, new_n993_, new_n994_, new_n995_,
    new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_, new_n1001_,
    new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1062_,
    new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_, new_n1068_,
    new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_, new_n1074_,
    new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_, new_n1080_,
    new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_, new_n1086_,
    new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1098_,
    new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_, new_n1104_,
    new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_, new_n1110_,
    new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_, new_n1116_,
    new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_, new_n1122_,
    new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_, new_n1128_,
    new_n1129_, new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_,
    new_n1136_, new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_,
    new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_,
    new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_,
    new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_,
    new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_,
    new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_,
    new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_,
    new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_,
    new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_,
    new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_,
    new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_,
    new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_,
    new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_, new_n1566_,
    new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_, new_n1572_,
    new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_, new_n1578_,
    new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_, new_n1584_,
    new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_, new_n1590_,
    new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_, new_n1596_,
    new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_, new_n1602_,
    new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_, new_n1608_,
    new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_, new_n1614_,
    new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_, new_n1620_,
    new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_, new_n1626_,
    new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_, new_n1632_,
    new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_, new_n1638_,
    new_n1639_, new_n1640_, new_n1642_, new_n1643_, new_n1644_, new_n1645_,
    new_n1646_, new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_,
    new_n1652_, new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_,
    new_n1658_, new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_,
    new_n1664_, new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_,
    new_n1670_, new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_,
    new_n1676_, new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_,
    new_n1682_, new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_,
    new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_,
    new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_,
    new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_,
    new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_,
    new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_,
    new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_,
    new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_,
    new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_,
    new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_,
    new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2150_, new_n2151_, new_n2152_, new_n2153_, new_n2154_,
    new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_, new_n2160_,
    new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_, new_n2166_,
    new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_, new_n2172_,
    new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_, new_n2178_,
    new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_, new_n2184_,
    new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_, new_n2190_,
    new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_, new_n2196_,
    new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_, new_n2202_,
    new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_, new_n2208_,
    new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_, new_n2214_,
    new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_, new_n2220_,
    new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_, new_n2226_,
    new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_, new_n2232_,
    new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_, new_n2238_,
    new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_, new_n2244_,
    new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_, new_n2250_,
    new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_, new_n2256_,
    new_n2257_, new_n2258_, new_n2260_, new_n2261_, new_n2262_, new_n2263_,
    new_n2264_, new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_,
    new_n2270_, new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_,
    new_n2276_, new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_,
    new_n2282_, new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_,
    new_n2288_, new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_,
    new_n2294_, new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_,
    new_n2300_, new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_,
    new_n2306_, new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_,
    new_n2312_, new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_,
    new_n2318_, new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_,
    new_n2324_, new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_,
    new_n2330_, new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_,
    new_n2336_, new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_,
    new_n2342_, new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_,
    new_n2348_, new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_,
    new_n2354_, new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_,
    new_n2360_, new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_,
    new_n2366_, new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_,
    new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_,
    new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_,
    new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_,
    new_n2427_, new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_,
    new_n2433_, new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_,
    new_n2439_, new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_,
    new_n2445_, new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_,
    new_n2451_, new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_,
    new_n2457_, new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_,
    new_n2463_, new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_,
    new_n2469_, new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_,
    new_n2475_, new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_,
    new_n2481_, new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_,
    new_n2487_, new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_,
    new_n2493_, new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_,
    new_n2499_, new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_,
    new_n2505_, new_n2506_, new_n2507_, new_n2509_, new_n2510_, new_n2511_,
    new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_,
    new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_,
    new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_,
    new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_,
    new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_,
    new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_,
    new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_,
    new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_,
    new_n2620_, new_n2621_, new_n2622_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_, new_n2880_,
    new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_, new_n2886_,
    new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_, new_n2892_,
    new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_, new_n2898_,
    new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_, new_n2904_,
    new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_, new_n2910_,
    new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_, new_n2916_,
    new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_, new_n2922_,
    new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_, new_n2928_,
    new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_, new_n2934_,
    new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_, new_n2940_,
    new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_, new_n2946_,
    new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_, new_n2952_,
    new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_, new_n2958_,
    new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_, new_n2964_,
    new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_, new_n2970_,
    new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_, new_n2976_,
    new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_, new_n2982_,
    new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_, new_n2988_,
    new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_, new_n2994_,
    new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n3000_, new_n3001_,
    new_n3002_, new_n3003_, new_n3004_, new_n3005_, new_n3006_, new_n3007_,
    new_n3008_, new_n3009_, new_n3010_, new_n3011_, new_n3012_, new_n3013_,
    new_n3014_, new_n3015_, new_n3016_, new_n3017_, new_n3018_, new_n3019_,
    new_n3020_, new_n3021_, new_n3022_, new_n3023_, new_n3024_, new_n3025_,
    new_n3026_, new_n3027_, new_n3028_, new_n3029_, new_n3030_, new_n3031_,
    new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_, new_n3037_,
    new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_, new_n3043_,
    new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_, new_n3049_,
    new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_, new_n3055_,
    new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_, new_n3061_,
    new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_, new_n3067_,
    new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_, new_n3073_,
    new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_, new_n3079_,
    new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_, new_n3085_,
    new_n3086_, new_n3087_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_,
    new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_,
    new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_,
    new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_,
    new_n3128_, new_n3129_, new_n3130_, new_n3131_, new_n3132_, new_n3133_,
    new_n3134_, new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_,
    new_n3183_, new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_,
    new_n3189_, new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_,
    new_n3195_, new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_,
    new_n3201_, new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_,
    new_n3207_, new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_,
    new_n3213_, new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_,
    new_n3219_, new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_,
    new_n3225_, new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_,
    new_n3231_, new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_,
    new_n3237_, new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_,
    new_n3243_, new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_,
    new_n3249_, new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_,
    new_n3255_, new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_,
    new_n3261_, new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_,
    new_n3267_, new_n3268_, new_n3269_, new_n3270_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3412_,
    new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_,
    new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_,
    new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_,
    new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_,
    new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_,
    new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_,
    new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_,
    new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_,
    new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_,
    new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_,
    new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_,
    new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_,
    new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_,
    new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_,
    new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_,
    new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_,
    new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_,
    new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_,
    new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_,
    new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_,
    new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_,
    new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_,
    new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3698_, new_n3699_, new_n3700_, new_n3701_, new_n3702_,
    new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_, new_n3708_,
    new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_, new_n3714_,
    new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_, new_n3720_,
    new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_, new_n3726_,
    new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_, new_n3732_,
    new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_, new_n3738_,
    new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_, new_n3744_,
    new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_, new_n3750_,
    new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_, new_n3756_,
    new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_, new_n3762_,
    new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_, new_n3768_,
    new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_, new_n3774_,
    new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_, new_n3780_,
    new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_, new_n3786_,
    new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_, new_n3792_,
    new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_, new_n3798_,
    new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_, new_n3804_,
    new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_, new_n3810_,
    new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_, new_n3816_,
    new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_, new_n3822_,
    new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_, new_n3828_,
    new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_, new_n3834_,
    new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_, new_n3840_,
    new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_, new_n3846_,
    new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_, new_n3852_,
    new_n3854_, new_n3855_, new_n3856_, new_n3857_, new_n3858_, new_n3859_,
    new_n3860_, new_n3861_, new_n3862_, new_n3863_, new_n3864_, new_n3865_,
    new_n3866_, new_n3867_, new_n3868_, new_n3869_, new_n3870_, new_n3871_,
    new_n3872_, new_n3873_, new_n3874_, new_n3875_, new_n3876_, new_n3877_,
    new_n3878_, new_n3879_, new_n3880_, new_n3881_, new_n3882_, new_n3883_,
    new_n3884_, new_n3885_, new_n3886_, new_n3887_, new_n3888_, new_n3889_,
    new_n3890_, new_n3891_, new_n3892_, new_n3893_, new_n3894_, new_n3895_,
    new_n3896_, new_n3897_, new_n3898_, new_n3899_, new_n3900_, new_n3901_,
    new_n3902_, new_n3903_, new_n3904_, new_n3905_, new_n3906_, new_n3907_,
    new_n3908_, new_n3909_, new_n3910_, new_n3911_, new_n3912_, new_n3913_,
    new_n3914_, new_n3915_, new_n3916_, new_n3917_, new_n3918_, new_n3919_,
    new_n3920_, new_n3921_, new_n3922_, new_n3923_, new_n3924_, new_n3925_,
    new_n3926_, new_n3927_, new_n3928_, new_n3929_, new_n3930_, new_n3931_,
    new_n3932_, new_n3933_, new_n3934_, new_n3935_, new_n3936_, new_n3937_,
    new_n3938_, new_n3939_, new_n3940_, new_n3941_, new_n3942_, new_n3943_,
    new_n3944_, new_n3945_, new_n3946_, new_n3947_, new_n3948_, new_n3949_,
    new_n3950_, new_n3951_, new_n3952_, new_n3953_, new_n3954_, new_n3955_,
    new_n3956_, new_n3957_, new_n3958_, new_n3959_, new_n3960_, new_n3961_,
    new_n3962_, new_n3963_, new_n3964_, new_n3965_, new_n3966_, new_n3967_,
    new_n3968_, new_n3969_, new_n3970_, new_n3971_, new_n3972_, new_n3973_,
    new_n3974_, new_n3975_, new_n3976_, new_n3977_, new_n3978_, new_n3979_,
    new_n3980_, new_n3981_, new_n3982_, new_n3983_, new_n3984_, new_n3985_,
    new_n3986_, new_n3987_, new_n3988_, new_n3989_, new_n3990_, new_n3991_,
    new_n3992_, new_n3993_, new_n3994_, new_n3995_, new_n3996_, new_n3997_,
    new_n3998_, new_n3999_, new_n4000_, new_n4002_, new_n4003_, new_n4004_,
    new_n4005_, new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_,
    new_n4011_, new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_,
    new_n4017_, new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_,
    new_n4023_, new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_,
    new_n4029_, new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_,
    new_n4035_, new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_,
    new_n4041_, new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_,
    new_n4047_, new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_,
    new_n4053_, new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_,
    new_n4059_, new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_,
    new_n4065_, new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_,
    new_n4071_, new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_,
    new_n4077_, new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_,
    new_n4083_, new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_,
    new_n4089_, new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_,
    new_n4095_, new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_,
    new_n4101_, new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_,
    new_n4107_, new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_,
    new_n4113_, new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_,
    new_n4119_, new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_,
    new_n4125_, new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_,
    new_n4131_, new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_,
    new_n4137_, new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_,
    new_n4143_, new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_,
    new_n4149_, new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_,
    new_n4155_, new_n4156_, new_n4157_, new_n4158_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4311_, new_n4312_,
    new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_,
    new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_,
    new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_,
    new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_,
    new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_,
    new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_,
    new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_,
    new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_,
    new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_,
    new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_,
    new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_,
    new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_,
    new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_,
    new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_,
    new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_,
    new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_,
    new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_,
    new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_,
    new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_,
    new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_,
    new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_,
    new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_,
    new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_,
    new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_,
    new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_,
    new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_, new_n4626_,
    new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_, new_n4632_,
    new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_, new_n4638_,
    new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_, new_n4644_,
    new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_, new_n4650_,
    new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_, new_n4656_,
    new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_, new_n4662_,
    new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_, new_n4668_,
    new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_, new_n4674_,
    new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_, new_n4680_,
    new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_, new_n4686_,
    new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_, new_n4692_,
    new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_, new_n4698_,
    new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_, new_n4704_,
    new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_, new_n4710_,
    new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_, new_n4716_,
    new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_, new_n4722_,
    new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_, new_n4728_,
    new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_, new_n4734_,
    new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_, new_n4740_,
    new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_, new_n4746_,
    new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_, new_n4752_,
    new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_, new_n4758_,
    new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_, new_n4764_,
    new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_, new_n4770_,
    new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_, new_n4776_,
    new_n4777_, new_n4778_, new_n4779_, new_n4781_, new_n4782_, new_n4783_,
    new_n4784_, new_n4785_, new_n4786_, new_n4787_, new_n4788_, new_n4789_,
    new_n4790_, new_n4791_, new_n4792_, new_n4793_, new_n4794_, new_n4795_,
    new_n4796_, new_n4797_, new_n4798_, new_n4799_, new_n4800_, new_n4801_,
    new_n4802_, new_n4803_, new_n4804_, new_n4805_, new_n4806_, new_n4807_,
    new_n4808_, new_n4809_, new_n4810_, new_n4811_, new_n4812_, new_n4813_,
    new_n4814_, new_n4815_, new_n4816_, new_n4817_, new_n4818_, new_n4819_,
    new_n4820_, new_n4821_, new_n4822_, new_n4823_, new_n4824_, new_n4825_,
    new_n4826_, new_n4827_, new_n4828_, new_n4829_, new_n4830_, new_n4831_,
    new_n4832_, new_n4833_, new_n4834_, new_n4835_, new_n4836_, new_n4837_,
    new_n4838_, new_n4839_, new_n4840_, new_n4841_, new_n4842_, new_n4843_,
    new_n4844_, new_n4845_, new_n4846_, new_n4847_, new_n4848_, new_n4849_,
    new_n4850_, new_n4851_, new_n4852_, new_n4853_, new_n4854_, new_n4855_,
    new_n4856_, new_n4857_, new_n4858_, new_n4859_, new_n4860_, new_n4861_,
    new_n4862_, new_n4863_, new_n4864_, new_n4865_, new_n4866_, new_n4867_,
    new_n4868_, new_n4869_, new_n4870_, new_n4871_, new_n4872_, new_n4873_,
    new_n4874_, new_n4875_, new_n4876_, new_n4877_, new_n4878_, new_n4879_,
    new_n4880_, new_n4881_, new_n4882_, new_n4883_, new_n4884_, new_n4885_,
    new_n4886_, new_n4887_, new_n4888_, new_n4889_, new_n4890_, new_n4891_,
    new_n4892_, new_n4893_, new_n4894_, new_n4895_, new_n4896_, new_n4897_,
    new_n4898_, new_n4899_, new_n4900_, new_n4901_, new_n4902_, new_n4903_,
    new_n4904_, new_n4905_, new_n4906_, new_n4907_, new_n4908_, new_n4909_,
    new_n4910_, new_n4911_, new_n4912_, new_n4913_, new_n4914_, new_n4915_,
    new_n4916_, new_n4917_, new_n4918_, new_n4919_, new_n4920_, new_n4921_,
    new_n4922_, new_n4923_, new_n4924_, new_n4925_, new_n4926_, new_n4927_,
    new_n4928_, new_n4929_, new_n4930_, new_n4931_, new_n4932_, new_n4933_,
    new_n4934_, new_n4935_, new_n4936_, new_n4937_, new_n4938_, new_n4939_,
    new_n4941_, new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_,
    new_n4947_, new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_,
    new_n4953_, new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_,
    new_n4959_, new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_,
    new_n4965_, new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_,
    new_n4971_, new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_,
    new_n4977_, new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_,
    new_n4983_, new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_,
    new_n4989_, new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_,
    new_n4995_, new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_,
    new_n5001_, new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_,
    new_n5007_, new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_,
    new_n5013_, new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_,
    new_n5019_, new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_,
    new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_,
    new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_,
    new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_,
    new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_,
    new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_,
    new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_,
    new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_,
    new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_,
    new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_,
    new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_,
    new_n5085_, new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_,
    new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_,
    new_n5097_, new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_,
    new_n5103_, new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_,
    new_n5109_, new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_,
    new_n5115_, new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_,
    new_n5121_, new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_,
    new_n5127_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_,
    new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_,
    new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_,
    new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_,
    new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_,
    new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_,
    new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_,
    new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_,
    new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_,
    new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_,
    new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_,
    new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_,
    new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_,
    new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_,
    new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_,
    new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_,
    new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_,
    new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_,
    new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_,
    new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_,
    new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_,
    new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_,
    new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_,
    new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_,
    new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_,
    new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_,
    new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_,
    new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_,
    new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_,
    new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_,
    new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_,
    new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_,
    new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_,
    new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_,
    new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_,
    new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_,
    new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_,
    new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_,
    new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_,
    new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5676_,
    new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_, new_n5682_,
    new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_, new_n5688_,
    new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_, new_n5694_,
    new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_, new_n5700_,
    new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_, new_n5706_,
    new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_, new_n5712_,
    new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_, new_n5778_,
    new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_,
    new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_,
    new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_,
    new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_,
    new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_,
    new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_,
    new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_, new_n5820_,
    new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_, new_n5826_,
    new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_, new_n5832_,
    new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_, new_n5838_,
    new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_, new_n5844_,
    new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_, new_n5850_,
    new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_, new_n5856_,
    new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_, new_n5862_,
    new_n5864_, new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_,
    new_n5870_, new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_,
    new_n5876_, new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_,
    new_n5882_, new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_,
    new_n5888_, new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_,
    new_n5894_, new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_,
    new_n5900_, new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_,
    new_n5906_, new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_,
    new_n5912_, new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_,
    new_n5918_, new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_,
    new_n5924_, new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_,
    new_n5930_, new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_,
    new_n5936_, new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_,
    new_n5942_, new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_,
    new_n5948_, new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_,
    new_n5954_, new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_,
    new_n5960_, new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_,
    new_n5966_, new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_,
    new_n5972_, new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_,
    new_n5978_, new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_,
    new_n5984_, new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_,
    new_n5990_, new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_,
    new_n5996_, new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_,
    new_n6002_, new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_,
    new_n6008_, new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_,
    new_n6014_, new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_,
    new_n6020_, new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_,
    new_n6026_, new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_,
    new_n6032_, new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_,
    new_n6038_, new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_,
    new_n6044_, new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_,
    new_n6050_, new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_,
    new_n6056_, new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_,
    new_n6062_, new_n6063_, new_n6064_, new_n6066_, new_n6067_, new_n6068_,
    new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_,
    new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_,
    new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_,
    new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_,
    new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_,
    new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_,
    new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_,
    new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_,
    new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_,
    new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_,
    new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_,
    new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_,
    new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_,
    new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_,
    new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_,
    new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_,
    new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_,
    new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_,
    new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_,
    new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_,
    new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_,
    new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_,
    new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_,
    new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_,
    new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_,
    new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_,
    new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_,
    new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_,
    new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_,
    new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_,
    new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_,
    new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_,
    new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_,
    new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_,
    new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_,
    new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_,
    new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_,
    new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_,
    new_n6316_, new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_,
    new_n6322_, new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_,
    new_n6328_, new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_,
    new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_,
    new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_,
    new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_,
    new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_,
    new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_,
    new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_,
    new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_,
    new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_,
    new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_,
    new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_,
    new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_,
    new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_,
    new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_,
    new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_,
    new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_,
    new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_,
    new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_,
    new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_,
    new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_,
    new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_,
    new_n6454_, new_n6455_, new_n6456_, new_n6458_, new_n6459_, new_n6460_,
    new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_,
    new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_,
    new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_,
    new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_,
    new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_,
    new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_,
    new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_,
    new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_,
    new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_,
    new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_,
    new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_,
    new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_,
    new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_,
    new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_,
    new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_,
    new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_,
    new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_,
    new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_,
    new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_,
    new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_,
    new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_,
    new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_,
    new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_,
    new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_,
    new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_,
    new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_,
    new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_,
    new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_,
    new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_,
    new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_,
    new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_,
    new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_,
    new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_,
    new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_,
    new_n6828_, new_n6829_, new_n6831_, new_n6832_, new_n6833_, new_n6834_,
    new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_,
    new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_,
    new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_,
    new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_,
    new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_,
    new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_,
    new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_,
    new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_,
    new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_,
    new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_,
    new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_,
    new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_,
    new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_,
    new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_,
    new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_,
    new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_,
    new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_,
    new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_,
    new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_,
    new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_,
    new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_,
    new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_,
    new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_,
    new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_,
    new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_,
    new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_,
    new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_,
    new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_,
    new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_,
    new_n7009_, new_n7010_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7208_,
    new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_,
    new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_,
    new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_,
    new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_,
    new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_,
    new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_,
    new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_,
    new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_,
    new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_,
    new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_,
    new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_,
    new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_,
    new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_,
    new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_,
    new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_,
    new_n7299_, new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_,
    new_n7305_, new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_,
    new_n7311_, new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_,
    new_n7317_, new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_,
    new_n7323_, new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_,
    new_n7329_, new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_,
    new_n7335_, new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_,
    new_n7341_, new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_,
    new_n7347_, new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_,
    new_n7353_, new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_,
    new_n7359_, new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_,
    new_n7365_, new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_,
    new_n7371_, new_n7372_, new_n7373_, new_n7374_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7546_,
    new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_,
    new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_,
    new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_,
    new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_,
    new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_,
    new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_,
    new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_,
    new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_,
    new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_,
    new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_,
    new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_,
    new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_,
    new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_,
    new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_,
    new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_,
    new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_,
    new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_,
    new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_,
    new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_,
    new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_,
    new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_,
    new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_,
    new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_,
    new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_,
    new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_,
    new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_,
    new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_,
    new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_,
    new_n7727_, new_n7728_, new_n7730_, new_n7731_, new_n7732_, new_n7733_,
    new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_,
    new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_,
    new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_,
    new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_,
    new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_,
    new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_,
    new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_,
    new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_,
    new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_,
    new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_,
    new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_,
    new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_,
    new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_,
    new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_,
    new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_,
    new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_,
    new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_,
    new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_,
    new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_,
    new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_,
    new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_,
    new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_,
    new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_,
    new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_, new_n7890_,
    new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_, new_n7896_,
    new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_, new_n7902_,
    new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_, new_n7908_,
    new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_, new_n7914_,
    new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_, new_n7920_,
    new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_, new_n7926_,
    new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_, new_n7932_,
    new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_, new_n7938_,
    new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_, new_n7944_,
    new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_, new_n7950_,
    new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_, new_n7956_,
    new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_, new_n7962_,
    new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_, new_n7968_,
    new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_, new_n7974_,
    new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_, new_n7980_,
    new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_, new_n7986_,
    new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_, new_n7992_,
    new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_, new_n7998_,
    new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_, new_n8004_,
    new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_, new_n8010_,
    new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_, new_n8016_,
    new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_, new_n8022_,
    new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_, new_n8028_,
    new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_, new_n8034_,
    new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_, new_n8040_,
    new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_, new_n8046_,
    new_n8047_, new_n8048_, new_n8049_, new_n8051_, new_n8052_, new_n8053_,
    new_n8054_, new_n8055_, new_n8056_, new_n8057_, new_n8058_, new_n8059_,
    new_n8060_, new_n8061_, new_n8062_, new_n8063_, new_n8064_, new_n8065_,
    new_n8066_, new_n8067_, new_n8068_, new_n8069_, new_n8070_, new_n8071_,
    new_n8072_, new_n8073_, new_n8074_, new_n8075_, new_n8076_, new_n8077_,
    new_n8078_, new_n8079_, new_n8080_, new_n8081_, new_n8082_, new_n8083_,
    new_n8084_, new_n8085_, new_n8086_, new_n8087_, new_n8088_, new_n8089_,
    new_n8090_, new_n8091_, new_n8092_, new_n8093_, new_n8094_, new_n8095_,
    new_n8096_, new_n8097_, new_n8098_, new_n8099_, new_n8100_, new_n8101_,
    new_n8102_, new_n8103_, new_n8104_, new_n8105_, new_n8106_, new_n8107_,
    new_n8108_, new_n8109_, new_n8110_, new_n8111_, new_n8112_, new_n8113_,
    new_n8114_, new_n8115_, new_n8116_, new_n8117_, new_n8118_, new_n8119_,
    new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_, new_n8125_,
    new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_, new_n8131_,
    new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_, new_n8137_,
    new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_, new_n8143_,
    new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_, new_n8149_,
    new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_, new_n8155_,
    new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_, new_n8161_,
    new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_, new_n8167_,
    new_n8168_, new_n8169_, new_n8170_, new_n8171_, new_n8172_, new_n8173_,
    new_n8174_, new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_,
    new_n8180_, new_n8181_, new_n8182_, new_n8183_, new_n8184_, new_n8185_,
    new_n8186_, new_n8187_, new_n8188_, new_n8189_, new_n8190_, new_n8191_,
    new_n8192_, new_n8193_, new_n8194_, new_n8195_, new_n8196_, new_n8197_,
    new_n8198_, new_n8199_, new_n8200_, new_n8201_, new_n8202_, new_n8203_,
    new_n8204_, new_n8205_, new_n8206_, new_n8207_, new_n8208_, new_n8209_,
    new_n8210_, new_n8211_, new_n8212_, new_n8213_, new_n8214_, new_n8216_,
    new_n8217_, new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_,
    new_n8223_, new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_,
    new_n8229_, new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_,
    new_n8235_, new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_,
    new_n8241_, new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8246_,
    new_n8247_, new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_,
    new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_,
    new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_,
    new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_,
    new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_,
    new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_,
    new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_,
    new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_,
    new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_,
    new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_,
    new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_,
    new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_,
    new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_,
    new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_,
    new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_,
    new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_,
    new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_,
    new_n8349_, new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_,
    new_n8355_, new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_,
    new_n8361_, new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_,
    new_n8367_, new_n8368_, new_n8369_, new_n8370_, new_n8372_, new_n8373_,
    new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_,
    new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_,
    new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_,
    new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_,
    new_n8398_, new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_,
    new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_,
    new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_,
    new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_,
    new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_,
    new_n8428_, new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_,
    new_n8434_, new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_,
    new_n8440_, new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_,
    new_n8446_, new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_,
    new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_,
    new_n8458_, new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_,
    new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_,
    new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_,
    new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_,
    new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_,
    new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_,
    new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_,
    new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_,
    new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_,
    new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_,
    new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_,
    new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8529_, new_n8530_,
    new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_,
    new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_,
    new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_,
    new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_,
    new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_,
    new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_,
    new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_,
    new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_,
    new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_,
    new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_,
    new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_,
    new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_,
    new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_,
    new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_,
    new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_,
    new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_,
    new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_,
    new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_,
    new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_,
    new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_,
    new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_,
    new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_,
    new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_,
    new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_,
    new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_,
    new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_,
    new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_,
    new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_,
    new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_,
    new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_,
    new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_,
    new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_,
    new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_,
    new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_,
    new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_,
    new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_,
    new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_,
    new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_,
    new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_,
    new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_,
    new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_,
    new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_,
    new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_,
    new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_,
    new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_,
    new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_,
    new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_,
    new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_,
    new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_,
    new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_,
    new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_,
    new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_,
    new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_,
    new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_,
    new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_,
    new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_,
    new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_,
    new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_,
    new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_,
    new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_,
    new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_,
    new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_,
    new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_,
    new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_,
    new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_,
    new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_,
    new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_,
    new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_,
    new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_,
    new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_,
    new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9110_,
    new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_,
    new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_,
    new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_,
    new_n9141_, new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_,
    new_n9147_, new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_,
    new_n9153_, new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_,
    new_n9159_, new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_,
    new_n9165_, new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_,
    new_n9171_, new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_,
    new_n9177_, new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_,
    new_n9183_, new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_,
    new_n9189_, new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_,
    new_n9195_, new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_,
    new_n9201_, new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_,
    new_n9207_, new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_,
    new_n9213_, new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_,
    new_n9219_, new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_,
    new_n9225_, new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_,
    new_n9231_, new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_,
    new_n9237_, new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_,
    new_n9243_, new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_,
    new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9382_,
    new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_,
    new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_,
    new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_,
    new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_,
    new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_,
    new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_,
    new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_,
    new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_,
    new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_,
    new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_,
    new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_,
    new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_,
    new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_,
    new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_,
    new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_,
    new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_,
    new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_,
    new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_,
    new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_,
    new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_,
    new_n9509_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9646_, new_n9647_, new_n9648_,
    new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_, new_n9654_,
    new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_, new_n9660_,
    new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_, new_n9666_,
    new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_,
    new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_, new_n9678_,
    new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_, new_n9684_,
    new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_, new_n9690_,
    new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_,
    new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_,
    new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_,
    new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_,
    new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_,
    new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_,
    new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_,
    new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_,
    new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_,
    new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_,
    new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_,
    new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_,
    new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_,
    new_n9769_, new_n9771_, new_n9772_, new_n9773_, new_n9774_, new_n9775_,
    new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_, new_n9781_,
    new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_, new_n9787_,
    new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_, new_n9793_,
    new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_, new_n9799_,
    new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_, new_n9805_,
    new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_, new_n9811_,
    new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_, new_n9817_,
    new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_, new_n9823_,
    new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_, new_n9829_,
    new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_, new_n9835_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_,
    new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_,
    new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_,
    new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_,
    new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_,
    new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_,
    new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_,
    new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_,
    new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_,
    new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_,
    new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_,
    new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_,
    new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_,
    new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_,
    new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_,
    new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_,
    new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_,
    new_n9999_, new_n10000_, new_n10001_, new_n10002_, new_n10003_,
    new_n10004_, new_n10005_, new_n10006_, new_n10007_, new_n10008_,
    new_n10009_, new_n10010_, new_n10011_, new_n10012_, new_n10013_,
    new_n10014_, new_n10015_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10242_, new_n10243_, new_n10244_, new_n10245_, new_n10246_,
    new_n10247_, new_n10248_, new_n10249_, new_n10250_, new_n10251_,
    new_n10252_, new_n10253_, new_n10254_, new_n10255_, new_n10256_,
    new_n10257_, new_n10258_, new_n10259_, new_n10260_, new_n10261_,
    new_n10262_, new_n10263_, new_n10264_, new_n10265_, new_n10266_,
    new_n10267_, new_n10268_, new_n10269_, new_n10270_, new_n10271_,
    new_n10272_, new_n10273_, new_n10274_, new_n10275_, new_n10276_,
    new_n10277_, new_n10278_, new_n10279_, new_n10280_, new_n10281_,
    new_n10282_, new_n10283_, new_n10284_, new_n10285_, new_n10286_,
    new_n10287_, new_n10288_, new_n10289_, new_n10290_, new_n10291_,
    new_n10292_, new_n10293_, new_n10294_, new_n10295_, new_n10296_,
    new_n10297_, new_n10298_, new_n10299_, new_n10300_, new_n10301_,
    new_n10302_, new_n10303_, new_n10304_, new_n10305_, new_n10306_,
    new_n10307_, new_n10308_, new_n10309_, new_n10310_, new_n10311_,
    new_n10312_, new_n10313_, new_n10314_, new_n10315_, new_n10316_,
    new_n10317_, new_n10318_, new_n10319_, new_n10320_, new_n10321_,
    new_n10322_, new_n10323_, new_n10324_, new_n10325_, new_n10326_,
    new_n10327_, new_n10328_, new_n10329_, new_n10330_, new_n10331_,
    new_n10332_, new_n10333_, new_n10334_, new_n10335_, new_n10336_,
    new_n10337_, new_n10338_, new_n10339_, new_n10340_, new_n10341_,
    new_n10342_, new_n10343_, new_n10344_, new_n10345_, new_n10346_,
    new_n10347_, new_n10348_, new_n10349_, new_n10350_, new_n10351_,
    new_n10353_, new_n10354_, new_n10355_, new_n10356_, new_n10357_,
    new_n10358_, new_n10359_, new_n10360_, new_n10361_, new_n10362_,
    new_n10363_, new_n10364_, new_n10365_, new_n10366_, new_n10367_,
    new_n10368_, new_n10369_, new_n10370_, new_n10371_, new_n10372_,
    new_n10373_, new_n10374_, new_n10375_, new_n10376_, new_n10377_,
    new_n10378_, new_n10379_, new_n10380_, new_n10381_, new_n10382_,
    new_n10383_, new_n10384_, new_n10385_, new_n10386_, new_n10387_,
    new_n10388_, new_n10389_, new_n10390_, new_n10391_, new_n10392_,
    new_n10393_, new_n10394_, new_n10395_, new_n10396_, new_n10397_,
    new_n10398_, new_n10399_, new_n10400_, new_n10401_, new_n10402_,
    new_n10403_, new_n10404_, new_n10405_, new_n10406_, new_n10407_,
    new_n10408_, new_n10409_, new_n10410_, new_n10411_, new_n10412_,
    new_n10413_, new_n10414_, new_n10415_, new_n10416_, new_n10417_,
    new_n10418_, new_n10419_, new_n10420_, new_n10421_, new_n10422_,
    new_n10423_, new_n10424_, new_n10425_, new_n10426_, new_n10427_,
    new_n10428_, new_n10429_, new_n10430_, new_n10431_, new_n10432_,
    new_n10433_, new_n10434_, new_n10435_, new_n10436_, new_n10437_,
    new_n10438_, new_n10439_, new_n10440_, new_n10441_, new_n10442_,
    new_n10443_, new_n10444_, new_n10445_, new_n10446_, new_n10447_,
    new_n10448_, new_n10449_, new_n10450_, new_n10451_, new_n10452_,
    new_n10453_, new_n10454_, new_n10455_, new_n10456_, new_n10457_,
    new_n10458_, new_n10459_, new_n10460_, new_n10461_, new_n10462_,
    new_n10463_, new_n10464_, new_n10465_, new_n10466_, new_n10467_,
    new_n10468_, new_n10469_, new_n10471_, new_n10472_, new_n10473_,
    new_n10474_, new_n10475_, new_n10476_, new_n10477_, new_n10478_,
    new_n10479_, new_n10480_, new_n10481_, new_n10482_, new_n10483_,
    new_n10484_, new_n10485_, new_n10486_, new_n10487_, new_n10488_,
    new_n10489_, new_n10490_, new_n10491_, new_n10492_, new_n10493_,
    new_n10494_, new_n10495_, new_n10496_, new_n10497_, new_n10498_,
    new_n10499_, new_n10500_, new_n10501_, new_n10502_, new_n10503_,
    new_n10504_, new_n10505_, new_n10506_, new_n10507_, new_n10508_,
    new_n10509_, new_n10510_, new_n10511_, new_n10512_, new_n10513_,
    new_n10514_, new_n10515_, new_n10516_, new_n10517_, new_n10518_,
    new_n10519_, new_n10520_, new_n10521_, new_n10522_, new_n10523_,
    new_n10524_, new_n10525_, new_n10526_, new_n10527_, new_n10528_,
    new_n10529_, new_n10530_, new_n10531_, new_n10532_, new_n10533_,
    new_n10534_, new_n10535_, new_n10536_, new_n10537_, new_n10538_,
    new_n10539_, new_n10540_, new_n10541_, new_n10542_, new_n10543_,
    new_n10544_, new_n10545_, new_n10546_, new_n10547_, new_n10548_,
    new_n10549_, new_n10550_, new_n10551_, new_n10552_, new_n10553_,
    new_n10554_, new_n10555_, new_n10556_, new_n10557_, new_n10558_,
    new_n10559_, new_n10560_, new_n10561_, new_n10562_, new_n10563_,
    new_n10564_, new_n10565_, new_n10566_, new_n10567_, new_n10568_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10776_,
    new_n10777_, new_n10778_, new_n10779_, new_n10780_, new_n10781_,
    new_n10782_, new_n10783_, new_n10784_, new_n10785_, new_n10786_,
    new_n10787_, new_n10788_, new_n10789_, new_n10790_, new_n10791_,
    new_n10792_, new_n10793_, new_n10794_, new_n10795_, new_n10796_,
    new_n10797_, new_n10798_, new_n10799_, new_n10800_, new_n10801_,
    new_n10802_, new_n10803_, new_n10804_, new_n10805_, new_n10806_,
    new_n10807_, new_n10808_, new_n10809_, new_n10810_, new_n10811_,
    new_n10812_, new_n10813_, new_n10814_, new_n10815_, new_n10816_,
    new_n10817_, new_n10818_, new_n10819_, new_n10820_, new_n10821_,
    new_n10822_, new_n10823_, new_n10824_, new_n10825_, new_n10826_,
    new_n10827_, new_n10828_, new_n10829_, new_n10830_, new_n10831_,
    new_n10832_, new_n10833_, new_n10834_, new_n10835_, new_n10836_,
    new_n10837_, new_n10838_, new_n10839_, new_n10840_, new_n10841_,
    new_n10842_, new_n10843_, new_n10844_, new_n10845_, new_n10846_,
    new_n10847_, new_n10848_, new_n10849_, new_n10850_, new_n10851_,
    new_n10852_, new_n10853_, new_n10854_, new_n10855_, new_n10856_,
    new_n10857_, new_n10858_, new_n10859_, new_n10860_, new_n10861_,
    new_n10862_, new_n10863_, new_n10864_, new_n10865_, new_n10866_,
    new_n10868_, new_n10869_, new_n10870_, new_n10871_, new_n10872_,
    new_n10873_, new_n10874_, new_n10875_, new_n10876_, new_n10877_,
    new_n10878_, new_n10879_, new_n10880_, new_n10881_, new_n10882_,
    new_n10883_, new_n10884_, new_n10885_, new_n10886_, new_n10887_,
    new_n10888_, new_n10889_, new_n10890_, new_n10891_, new_n10892_,
    new_n10893_, new_n10894_, new_n10895_, new_n10896_, new_n10897_,
    new_n10898_, new_n10899_, new_n10900_, new_n10901_, new_n10902_,
    new_n10903_, new_n10904_, new_n10905_, new_n10906_, new_n10907_,
    new_n10908_, new_n10909_, new_n10910_, new_n10911_, new_n10912_,
    new_n10913_, new_n10914_, new_n10915_, new_n10916_, new_n10917_,
    new_n10918_, new_n10919_, new_n10920_, new_n10921_, new_n10922_,
    new_n10923_, new_n10924_, new_n10925_, new_n10926_, new_n10927_,
    new_n10928_, new_n10929_, new_n10930_, new_n10931_, new_n10932_,
    new_n10933_, new_n10934_, new_n10935_, new_n10936_, new_n10937_,
    new_n10938_, new_n10939_, new_n10940_, new_n10941_, new_n10942_,
    new_n10943_, new_n10944_, new_n10945_, new_n10946_, new_n10947_,
    new_n10948_, new_n10949_, new_n10950_, new_n10951_, new_n10952_,
    new_n10953_, new_n10954_, new_n10955_, new_n10956_, new_n10957_,
    new_n10959_, new_n10960_, new_n10961_, new_n10962_, new_n10963_,
    new_n10964_, new_n10965_, new_n10966_, new_n10967_, new_n10968_,
    new_n10969_, new_n10970_, new_n10971_, new_n10972_, new_n10973_,
    new_n10974_, new_n10975_, new_n10976_, new_n10977_, new_n10978_,
    new_n10979_, new_n10980_, new_n10981_, new_n10982_, new_n10983_,
    new_n10984_, new_n10985_, new_n10986_, new_n10987_, new_n10988_,
    new_n10989_, new_n10990_, new_n10991_, new_n10992_, new_n10993_,
    new_n10994_, new_n10995_, new_n10996_, new_n10997_, new_n10998_,
    new_n10999_, new_n11000_, new_n11001_, new_n11002_, new_n11003_,
    new_n11004_, new_n11005_, new_n11006_, new_n11007_, new_n11008_,
    new_n11009_, new_n11010_, new_n11011_, new_n11012_, new_n11013_,
    new_n11014_, new_n11015_, new_n11016_, new_n11017_, new_n11018_,
    new_n11019_, new_n11020_, new_n11021_, new_n11022_, new_n11023_,
    new_n11024_, new_n11025_, new_n11026_, new_n11027_, new_n11028_,
    new_n11029_, new_n11030_, new_n11031_, new_n11032_, new_n11033_,
    new_n11034_, new_n11035_, new_n11036_, new_n11037_, new_n11038_,
    new_n11039_, new_n11040_, new_n11041_, new_n11042_, new_n11043_,
    new_n11044_, new_n11045_, new_n11046_, new_n11047_, new_n11048_,
    new_n11049_, new_n11050_, new_n11051_, new_n11052_, new_n11053_,
    new_n11054_, new_n11055_, new_n11056_, new_n11057_, new_n11058_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11073_, new_n11074_,
    new_n11075_, new_n11076_, new_n11077_, new_n11078_, new_n11079_,
    new_n11080_, new_n11081_, new_n11082_, new_n11083_, new_n11084_,
    new_n11085_, new_n11086_, new_n11087_, new_n11088_, new_n11089_,
    new_n11090_, new_n11091_, new_n11092_, new_n11093_, new_n11094_,
    new_n11095_, new_n11096_, new_n11097_, new_n11098_, new_n11099_,
    new_n11100_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11106_, new_n11107_, new_n11108_, new_n11109_,
    new_n11110_, new_n11111_, new_n11112_, new_n11113_, new_n11114_,
    new_n11115_, new_n11116_, new_n11117_, new_n11118_, new_n11119_,
    new_n11120_, new_n11121_, new_n11122_, new_n11123_, new_n11124_,
    new_n11125_, new_n11126_, new_n11127_, new_n11128_, new_n11129_,
    new_n11130_, new_n11131_, new_n11132_, new_n11133_, new_n11134_,
    new_n11135_, new_n11136_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11231_,
    new_n11232_, new_n11233_, new_n11234_, new_n11235_, new_n11236_,
    new_n11237_, new_n11238_, new_n11239_, new_n11240_, new_n11241_,
    new_n11242_, new_n11243_, new_n11244_, new_n11245_, new_n11246_,
    new_n11247_, new_n11248_, new_n11249_, new_n11250_, new_n11251_,
    new_n11252_, new_n11253_, new_n11254_, new_n11255_, new_n11256_,
    new_n11257_, new_n11258_, new_n11259_, new_n11260_, new_n11261_,
    new_n11262_, new_n11263_, new_n11264_, new_n11265_, new_n11266_,
    new_n11267_, new_n11268_, new_n11269_, new_n11270_, new_n11271_,
    new_n11272_, new_n11273_, new_n11274_, new_n11275_, new_n11276_,
    new_n11277_, new_n11278_, new_n11279_, new_n11280_, new_n11281_,
    new_n11282_, new_n11283_, new_n11284_, new_n11285_, new_n11286_,
    new_n11287_, new_n11288_, new_n11289_, new_n11290_, new_n11291_,
    new_n11292_, new_n11293_, new_n11294_, new_n11295_, new_n11296_,
    new_n11297_, new_n11298_, new_n11299_, new_n11300_, new_n11301_,
    new_n11302_, new_n11303_, new_n11304_, new_n11305_, new_n11306_,
    new_n11307_, new_n11308_, new_n11309_, new_n11310_, new_n11311_,
    new_n11312_, new_n11313_, new_n11314_, new_n11315_, new_n11316_,
    new_n11317_, new_n11319_, new_n11320_, new_n11321_, new_n11322_,
    new_n11323_, new_n11324_, new_n11325_, new_n11326_, new_n11327_,
    new_n11328_, new_n11329_, new_n11330_, new_n11331_, new_n11332_,
    new_n11333_, new_n11334_, new_n11335_, new_n11336_, new_n11337_,
    new_n11338_, new_n11339_, new_n11340_, new_n11341_, new_n11342_,
    new_n11343_, new_n11344_, new_n11345_, new_n11346_, new_n11347_,
    new_n11348_, new_n11349_, new_n11350_, new_n11351_, new_n11352_,
    new_n11353_, new_n11354_, new_n11355_, new_n11356_, new_n11357_,
    new_n11358_, new_n11359_, new_n11360_, new_n11361_, new_n11362_,
    new_n11363_, new_n11364_, new_n11365_, new_n11366_, new_n11367_,
    new_n11368_, new_n11369_, new_n11370_, new_n11371_, new_n11372_,
    new_n11373_, new_n11374_, new_n11375_, new_n11376_, new_n11377_,
    new_n11378_, new_n11379_, new_n11380_, new_n11381_, new_n11382_,
    new_n11383_, new_n11384_, new_n11385_, new_n11386_, new_n11387_,
    new_n11388_, new_n11389_, new_n11390_, new_n11391_, new_n11392_,
    new_n11393_, new_n11394_, new_n11396_, new_n11397_, new_n11398_,
    new_n11399_, new_n11400_, new_n11401_, new_n11402_, new_n11403_,
    new_n11404_, new_n11405_, new_n11406_, new_n11407_, new_n11408_,
    new_n11409_, new_n11410_, new_n11411_, new_n11412_, new_n11413_,
    new_n11414_, new_n11415_, new_n11416_, new_n11417_, new_n11418_,
    new_n11419_, new_n11420_, new_n11421_, new_n11422_, new_n11423_,
    new_n11424_, new_n11425_, new_n11426_, new_n11427_, new_n11428_,
    new_n11429_, new_n11430_, new_n11431_, new_n11432_, new_n11433_,
    new_n11434_, new_n11435_, new_n11436_, new_n11437_, new_n11438_,
    new_n11439_, new_n11440_, new_n11441_, new_n11442_, new_n11443_,
    new_n11444_, new_n11445_, new_n11446_, new_n11447_, new_n11448_,
    new_n11449_, new_n11450_, new_n11451_, new_n11452_, new_n11453_,
    new_n11454_, new_n11455_, new_n11456_, new_n11457_, new_n11458_,
    new_n11459_, new_n11460_, new_n11461_, new_n11462_, new_n11463_,
    new_n11464_, new_n11465_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11528_, new_n11529_,
    new_n11530_, new_n11531_, new_n11532_, new_n11533_, new_n11534_,
    new_n11535_, new_n11536_, new_n11537_, new_n11538_, new_n11539_,
    new_n11540_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11607_, new_n11608_, new_n11609_, new_n11610_, new_n11611_,
    new_n11612_, new_n11613_, new_n11614_, new_n11615_, new_n11616_,
    new_n11617_, new_n11618_, new_n11619_, new_n11620_, new_n11621_,
    new_n11622_, new_n11623_, new_n11624_, new_n11625_, new_n11626_,
    new_n11627_, new_n11628_, new_n11629_, new_n11630_, new_n11631_,
    new_n11632_, new_n11633_, new_n11634_, new_n11635_, new_n11636_,
    new_n11637_, new_n11638_, new_n11639_, new_n11640_, new_n11641_,
    new_n11642_, new_n11643_, new_n11644_, new_n11645_, new_n11646_,
    new_n11647_, new_n11648_, new_n11649_, new_n11650_, new_n11651_,
    new_n11652_, new_n11653_, new_n11654_, new_n11655_, new_n11656_,
    new_n11657_, new_n11658_, new_n11659_, new_n11660_, new_n11661_,
    new_n11662_, new_n11663_, new_n11664_, new_n11665_, new_n11666_,
    new_n11668_, new_n11669_, new_n11670_, new_n11671_, new_n11672_,
    new_n11673_, new_n11674_, new_n11675_, new_n11676_, new_n11677_,
    new_n11678_, new_n11679_, new_n11680_, new_n11681_, new_n11682_,
    new_n11683_, new_n11684_, new_n11685_, new_n11686_, new_n11687_,
    new_n11688_, new_n11689_, new_n11690_, new_n11691_, new_n11692_,
    new_n11693_, new_n11694_, new_n11695_, new_n11696_, new_n11697_,
    new_n11698_, new_n11699_, new_n11700_, new_n11701_, new_n11702_,
    new_n11703_, new_n11704_, new_n11705_, new_n11706_, new_n11707_,
    new_n11708_, new_n11709_, new_n11710_, new_n11711_, new_n11712_,
    new_n11713_, new_n11714_, new_n11715_, new_n11716_, new_n11717_,
    new_n11718_, new_n11719_, new_n11720_, new_n11721_, new_n11722_,
    new_n11723_, new_n11724_, new_n11725_, new_n11726_, new_n11727_,
    new_n11728_, new_n11729_, new_n11730_, new_n11731_, new_n11733_,
    new_n11734_, new_n11735_, new_n11736_, new_n11737_, new_n11738_,
    new_n11739_, new_n11740_, new_n11741_, new_n11742_, new_n11743_,
    new_n11744_, new_n11745_, new_n11746_, new_n11747_, new_n11748_,
    new_n11749_, new_n11750_, new_n11751_, new_n11752_, new_n11753_,
    new_n11754_, new_n11755_, new_n11756_, new_n11757_, new_n11758_,
    new_n11759_, new_n11760_, new_n11761_, new_n11762_, new_n11763_,
    new_n11764_, new_n11765_, new_n11766_, new_n11767_, new_n11768_,
    new_n11769_, new_n11770_, new_n11771_, new_n11772_, new_n11773_,
    new_n11774_, new_n11775_, new_n11776_, new_n11777_, new_n11778_,
    new_n11779_, new_n11780_, new_n11781_, new_n11782_, new_n11783_,
    new_n11784_, new_n11785_, new_n11786_, new_n11787_, new_n11788_,
    new_n11789_, new_n11790_, new_n11791_, new_n11792_, new_n11793_,
    new_n11794_, new_n11795_, new_n11797_, new_n11798_, new_n11799_,
    new_n11800_, new_n11801_, new_n11802_, new_n11803_, new_n11804_,
    new_n11805_, new_n11806_, new_n11807_, new_n11808_, new_n11809_,
    new_n11810_, new_n11811_, new_n11812_, new_n11813_, new_n11814_,
    new_n11815_, new_n11816_, new_n11817_, new_n11818_, new_n11819_,
    new_n11820_, new_n11821_, new_n11822_, new_n11823_, new_n11824_,
    new_n11825_, new_n11826_, new_n11827_, new_n11828_, new_n11829_,
    new_n11830_, new_n11831_, new_n11832_, new_n11833_, new_n11834_,
    new_n11835_, new_n11836_, new_n11837_, new_n11838_, new_n11839_,
    new_n11840_, new_n11841_, new_n11842_, new_n11843_, new_n11844_,
    new_n11845_, new_n11846_, new_n11847_, new_n11848_, new_n11849_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11906_,
    new_n11907_, new_n11908_, new_n11909_, new_n11910_, new_n11911_,
    new_n11912_, new_n11913_, new_n11914_, new_n11915_, new_n11916_,
    new_n11917_, new_n11918_, new_n11919_, new_n11920_, new_n11921_,
    new_n11922_, new_n11923_, new_n11924_, new_n11925_, new_n11926_,
    new_n11927_, new_n11928_, new_n11929_, new_n11930_, new_n11931_,
    new_n11932_, new_n11933_, new_n11934_, new_n11935_, new_n11936_,
    new_n11937_, new_n11938_, new_n11939_, new_n11940_, new_n11941_,
    new_n11942_, new_n11943_, new_n11944_, new_n11945_, new_n11946_,
    new_n11947_, new_n11948_, new_n11949_, new_n11950_, new_n11951_,
    new_n11952_, new_n11953_, new_n11954_, new_n11956_, new_n11957_,
    new_n11958_, new_n11959_, new_n11960_, new_n11961_, new_n11962_,
    new_n11963_, new_n11964_, new_n11965_, new_n11966_, new_n11967_,
    new_n11968_, new_n11969_, new_n11970_, new_n11971_, new_n11972_,
    new_n11973_, new_n11974_, new_n11975_, new_n11976_, new_n11977_,
    new_n11978_, new_n11979_, new_n11980_, new_n11981_, new_n11982_,
    new_n11983_, new_n11984_, new_n11985_, new_n11986_, new_n11987_,
    new_n11988_, new_n11989_, new_n11990_, new_n11991_, new_n11992_,
    new_n11993_, new_n11994_, new_n11995_, new_n11996_, new_n11997_,
    new_n11998_, new_n11999_, new_n12000_, new_n12001_, new_n12002_,
    new_n12003_, new_n12004_, new_n12005_, new_n12006_, new_n12007_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12056_, new_n12057_, new_n12058_, new_n12059_,
    new_n12060_, new_n12061_, new_n12062_, new_n12063_, new_n12064_,
    new_n12065_, new_n12066_, new_n12067_, new_n12068_, new_n12069_,
    new_n12070_, new_n12071_, new_n12072_, new_n12073_, new_n12074_,
    new_n12075_, new_n12076_, new_n12077_, new_n12078_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12084_,
    new_n12085_, new_n12086_, new_n12087_, new_n12088_, new_n12089_,
    new_n12090_, new_n12091_, new_n12092_, new_n12093_, new_n12094_,
    new_n12095_, new_n12096_, new_n12097_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12138_, new_n12139_, new_n12140_, new_n12141_,
    new_n12142_, new_n12143_, new_n12144_, new_n12145_, new_n12146_,
    new_n12147_, new_n12148_, new_n12149_, new_n12150_, new_n12151_,
    new_n12152_, new_n12153_, new_n12154_, new_n12155_, new_n12156_,
    new_n12157_, new_n12158_, new_n12159_, new_n12160_, new_n12161_,
    new_n12162_, new_n12163_, new_n12164_, new_n12165_, new_n12166_,
    new_n12167_, new_n12168_, new_n12169_, new_n12170_, new_n12171_,
    new_n12172_, new_n12173_, new_n12174_, new_n12175_, new_n12176_,
    new_n12177_, new_n12178_, new_n12179_, new_n12180_, new_n12182_,
    new_n12183_, new_n12184_, new_n12185_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12248_, new_n12249_,
    new_n12250_, new_n12251_, new_n12252_, new_n12253_, new_n12254_,
    new_n12255_, new_n12256_, new_n12257_, new_n12258_, new_n12259_,
    new_n12260_, new_n12261_, new_n12262_, new_n12263_, new_n12264_,
    new_n12265_, new_n12266_, new_n12267_, new_n12268_, new_n12269_,
    new_n12270_, new_n12271_, new_n12272_, new_n12273_, new_n12274_,
    new_n12275_, new_n12276_, new_n12277_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12304_, new_n12305_, new_n12306_,
    new_n12307_, new_n12308_, new_n12309_, new_n12310_, new_n12311_,
    new_n12312_, new_n12313_, new_n12314_, new_n12315_, new_n12316_,
    new_n12317_, new_n12318_, new_n12319_, new_n12320_, new_n12321_,
    new_n12322_, new_n12323_, new_n12324_, new_n12325_, new_n12326_,
    new_n12328_, new_n12329_, new_n12330_, new_n12331_, new_n12332_,
    new_n12333_, new_n12334_, new_n12335_, new_n12336_, new_n12337_,
    new_n12338_, new_n12339_, new_n12340_, new_n12341_, new_n12342_,
    new_n12343_, new_n12344_, new_n12345_, new_n12346_, new_n12348_,
    new_n12349_, new_n12350_, new_n12351_, new_n12352_, new_n12353_,
    new_n12354_, new_n12355_, new_n12356_, new_n12357_, new_n12358_,
    new_n12359_, new_n12360_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12380_,
    new_n12381_, new_n12382_, new_n12383_, new_n12385_, new_n12386_,
    new_n12387_, new_n12388_, new_n12389_, new_n12390_, new_n12391_,
    new_n12393_, new_n12394_, new_n12395_;
  INVX1    g00000(.A(\a[0] ), .Y(new_n194_));
  AND2X1   g00001(.A(\a[1] ), .B(new_n194_), .Y(\asquared[2] ));
  NAND2X1  g00002(.A(\a[1] ), .B(\a[0] ), .Y(new_n196_));
  AND2X1   g00003(.A(\a[2] ), .B(\a[0] ), .Y(new_n197_));
  INVX1    g00004(.A(new_n197_), .Y(new_n198_));
  XOR2X1   g00005(.A(new_n198_), .B(new_n196_), .Y(\asquared[3] ));
  INVX1    g00006(.A(\a[2] ), .Y(new_n200_));
  NOR3X1   g00007(.A(new_n196_), .B(new_n200_), .C(new_n194_), .Y(new_n201_));
  INVX1    g00008(.A(\a[1] ), .Y(new_n202_));
  AND2X1   g00009(.A(\a[2] ), .B(new_n202_), .Y(new_n203_));
  AND2X1   g00010(.A(\a[3] ), .B(\a[0] ), .Y(new_n204_));
  XOR2X1   g00011(.A(new_n204_), .B(new_n203_), .Y(new_n205_));
  XOR2X1   g00012(.A(new_n205_), .B(new_n201_), .Y(\asquared[4] ));
  NAND2X1  g00013(.A(\a[2] ), .B(\a[1] ), .Y(new_n207_));
  NAND4X1  g00014(.A(\a[4] ), .B(\a[3] ), .C(\a[1] ), .D(\a[0] ), .Y(new_n208_));
  AND2X1   g00015(.A(\a[3] ), .B(\a[1] ), .Y(new_n209_));
  AND2X1   g00016(.A(\a[4] ), .B(\a[0] ), .Y(new_n210_));
  OAI21X1  g00017(.A0(new_n210_), .A1(new_n209_), .B0(new_n208_), .Y(new_n211_));
  XOR2X1   g00018(.A(new_n211_), .B(new_n207_), .Y(new_n212_));
  NAND3X1  g00019(.A(\a[3] ), .B(\a[2] ), .C(\a[0] ), .Y(new_n213_));
  INVX1    g00020(.A(new_n213_), .Y(new_n214_));
  XOR2X1   g00021(.A(new_n214_), .B(new_n212_), .Y(\asquared[5] ));
  AOI22X1  g00022(.A0(\a[5] ), .A1(\a[0] ), .B0(\a[4] ), .B1(\a[1] ), .Y(new_n216_));
  NAND2X1  g00023(.A(\a[4] ), .B(\a[3] ), .Y(new_n217_));
  AND2X1   g00024(.A(\a[5] ), .B(\a[4] ), .Y(new_n218_));
  NOR4X1   g00025(.A(new_n218_), .B(new_n216_), .C(new_n217_), .D(new_n196_), .Y(new_n219_));
  NAND2X1  g00026(.A(\a[5] ), .B(\a[4] ), .Y(new_n220_));
  OAI22X1  g00027(.A0(new_n220_), .A1(new_n196_), .B0(new_n216_), .B1(new_n208_), .Y(new_n221_));
  OAI22X1  g00028(.A0(new_n221_), .A1(new_n216_), .B0(new_n219_), .B1(new_n208_), .Y(new_n222_));
  INVX1    g00029(.A(\a[3] ), .Y(new_n223_));
  OR2X1    g00030(.A(new_n223_), .B(\a[2] ), .Y(new_n224_));
  XOR2X1   g00031(.A(new_n224_), .B(new_n222_), .Y(new_n225_));
  NOR2X1   g00032(.A(new_n211_), .B(new_n207_), .Y(new_n226_));
  AOI21X1  g00033(.A0(new_n211_), .A1(new_n207_), .B0(new_n213_), .Y(new_n227_));
  NOR2X1   g00034(.A(new_n227_), .B(new_n226_), .Y(new_n228_));
  XOR2X1   g00035(.A(new_n228_), .B(new_n225_), .Y(\asquared[6] ));
  INVX1    g00036(.A(\a[6] ), .Y(new_n230_));
  AND2X1   g00037(.A(\a[3] ), .B(\a[2] ), .Y(new_n231_));
  AND2X1   g00038(.A(\a[6] ), .B(\a[0] ), .Y(new_n232_));
  OAI22X1  g00039(.A0(new_n232_), .A1(new_n231_), .B0(new_n213_), .B1(new_n230_), .Y(new_n233_));
  AND2X1   g00040(.A(\a[5] ), .B(\a[1] ), .Y(new_n234_));
  AND2X1   g00041(.A(\a[4] ), .B(\a[2] ), .Y(new_n235_));
  OAI22X1  g00042(.A0(new_n235_), .A1(new_n234_), .B0(new_n220_), .B1(new_n207_), .Y(new_n236_));
  XOR2X1   g00043(.A(new_n236_), .B(new_n233_), .Y(new_n237_));
  AND2X1   g00044(.A(new_n237_), .B(new_n221_), .Y(new_n238_));
  INVX1    g00045(.A(new_n238_), .Y(new_n239_));
  AND2X1   g00046(.A(\a[3] ), .B(new_n200_), .Y(new_n240_));
  NAND2X1  g00047(.A(new_n240_), .B(new_n222_), .Y(new_n241_));
  OAI22X1  g00048(.A0(new_n227_), .A1(new_n226_), .B0(new_n240_), .B1(new_n222_), .Y(new_n242_));
  NAND2X1  g00049(.A(new_n242_), .B(new_n241_), .Y(new_n243_));
  OR2X1    g00050(.A(new_n237_), .B(new_n221_), .Y(new_n244_));
  AOI21X1  g00051(.A0(new_n239_), .A1(new_n244_), .B0(new_n243_), .Y(new_n245_));
  AND2X1   g00052(.A(new_n244_), .B(new_n243_), .Y(new_n246_));
  AOI21X1  g00053(.A0(new_n246_), .A1(new_n239_), .B0(new_n245_), .Y(\asquared[7] ));
  AND2X1   g00054(.A(\a[7] ), .B(\a[0] ), .Y(new_n248_));
  NAND2X1  g00055(.A(\a[3] ), .B(\a[2] ), .Y(new_n249_));
  NAND4X1  g00056(.A(\a[7] ), .B(\a[4] ), .C(\a[3] ), .D(\a[0] ), .Y(new_n250_));
  NAND4X1  g00057(.A(\a[7] ), .B(\a[5] ), .C(\a[2] ), .D(\a[0] ), .Y(new_n251_));
  NAND2X1  g00058(.A(new_n251_), .B(new_n250_), .Y(new_n252_));
  OAI21X1  g00059(.A0(new_n220_), .A1(new_n249_), .B0(new_n252_), .Y(new_n253_));
  AOI21X1  g00060(.A0(new_n218_), .A1(new_n231_), .B0(new_n252_), .Y(new_n254_));
  INVX1    g00061(.A(\a[5] ), .Y(new_n255_));
  OAI21X1  g00062(.A0(new_n255_), .A1(new_n200_), .B0(new_n217_), .Y(new_n256_));
  AOI22X1  g00063(.A0(new_n256_), .A1(new_n254_), .B0(new_n253_), .B1(new_n248_), .Y(new_n257_));
  OAI22X1  g00064(.A0(new_n236_), .A1(new_n233_), .B0(new_n213_), .B1(new_n230_), .Y(new_n258_));
  NOR2X1   g00065(.A(new_n220_), .B(new_n207_), .Y(new_n259_));
  AND2X1   g00066(.A(\a[6] ), .B(\a[1] ), .Y(new_n260_));
  XOR2X1   g00067(.A(new_n260_), .B(\a[4] ), .Y(new_n261_));
  MX2X1    g00068(.A(new_n261_), .B(new_n260_), .S0(new_n259_), .Y(new_n262_));
  XOR2X1   g00069(.A(new_n262_), .B(new_n258_), .Y(new_n263_));
  XOR2X1   g00070(.A(new_n263_), .B(new_n257_), .Y(new_n264_));
  AOI21X1  g00071(.A0(new_n244_), .A1(new_n243_), .B0(new_n238_), .Y(new_n265_));
  XOR2X1   g00072(.A(new_n265_), .B(new_n264_), .Y(\asquared[8] ));
  NOR3X1   g00073(.A(new_n260_), .B(new_n220_), .C(new_n207_), .Y(new_n267_));
  AND2X1   g00074(.A(new_n262_), .B(new_n258_), .Y(new_n268_));
  OR2X1    g00075(.A(new_n268_), .B(new_n267_), .Y(new_n269_));
  OAI21X1  g00076(.A0(new_n220_), .A1(new_n249_), .B0(new_n253_), .Y(new_n270_));
  AND2X1   g00077(.A(\a[7] ), .B(\a[1] ), .Y(new_n271_));
  AND2X1   g00078(.A(\a[5] ), .B(\a[3] ), .Y(new_n272_));
  XOR2X1   g00079(.A(new_n272_), .B(new_n271_), .Y(new_n273_));
  XOR2X1   g00080(.A(new_n273_), .B(new_n270_), .Y(new_n274_));
  NAND3X1  g00081(.A(\a[6] ), .B(\a[4] ), .C(\a[1] ), .Y(new_n275_));
  AOI22X1  g00082(.A0(\a[8] ), .A1(\a[0] ), .B0(\a[6] ), .B1(\a[2] ), .Y(new_n276_));
  AND2X1   g00083(.A(\a[8] ), .B(\a[6] ), .Y(new_n277_));
  AND2X1   g00084(.A(new_n277_), .B(new_n197_), .Y(new_n278_));
  NOR3X1   g00085(.A(new_n278_), .B(new_n276_), .C(new_n275_), .Y(new_n279_));
  INVX1    g00086(.A(new_n277_), .Y(new_n280_));
  OAI22X1  g00087(.A0(new_n280_), .A1(new_n198_), .B0(new_n276_), .B1(new_n275_), .Y(new_n281_));
  OAI22X1  g00088(.A0(new_n281_), .A1(new_n276_), .B0(new_n279_), .B1(new_n275_), .Y(new_n282_));
  XOR2X1   g00089(.A(new_n282_), .B(new_n274_), .Y(new_n283_));
  XOR2X1   g00090(.A(new_n283_), .B(new_n269_), .Y(new_n284_));
  NOR2X1   g00091(.A(new_n262_), .B(new_n258_), .Y(new_n285_));
  OR2X1    g00092(.A(new_n285_), .B(new_n268_), .Y(new_n286_));
  AND2X1   g00093(.A(new_n286_), .B(new_n257_), .Y(new_n287_));
  OR2X1    g00094(.A(new_n286_), .B(new_n257_), .Y(new_n288_));
  OAI21X1  g00095(.A0(new_n265_), .A1(new_n287_), .B0(new_n288_), .Y(new_n289_));
  XOR2X1   g00096(.A(new_n289_), .B(new_n284_), .Y(\asquared[9] ));
  AND2X1   g00097(.A(new_n273_), .B(new_n270_), .Y(new_n291_));
  AOI21X1  g00098(.A0(new_n282_), .A1(new_n274_), .B0(new_n291_), .Y(new_n292_));
  INVX1    g00099(.A(new_n281_), .Y(new_n293_));
  INVX1    g00100(.A(new_n217_), .Y(new_n294_));
  AND2X1   g00101(.A(\a[6] ), .B(\a[5] ), .Y(new_n295_));
  NAND4X1  g00102(.A(\a[7] ), .B(\a[5] ), .C(\a[4] ), .D(\a[2] ), .Y(new_n296_));
  NAND4X1  g00103(.A(\a[7] ), .B(\a[6] ), .C(\a[3] ), .D(\a[2] ), .Y(new_n297_));
  AOI22X1  g00104(.A0(new_n297_), .A1(new_n296_), .B0(new_n295_), .B1(new_n294_), .Y(new_n298_));
  NAND4X1  g00105(.A(\a[6] ), .B(\a[5] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n299_));
  NAND3X1  g00106(.A(new_n297_), .B(new_n296_), .C(new_n299_), .Y(new_n300_));
  AOI22X1  g00107(.A0(\a[6] ), .A1(\a[3] ), .B0(\a[5] ), .B1(\a[4] ), .Y(new_n301_));
  NAND2X1  g00108(.A(\a[7] ), .B(\a[2] ), .Y(new_n302_));
  OAI22X1  g00109(.A0(new_n302_), .A1(new_n298_), .B0(new_n301_), .B1(new_n300_), .Y(new_n303_));
  AND2X1   g00110(.A(new_n303_), .B(new_n293_), .Y(new_n304_));
  XOR2X1   g00111(.A(new_n303_), .B(new_n293_), .Y(new_n305_));
  NAND4X1  g00112(.A(\a[7] ), .B(\a[5] ), .C(\a[3] ), .D(\a[1] ), .Y(new_n306_));
  AND2X1   g00113(.A(\a[9] ), .B(\a[0] ), .Y(new_n307_));
  XOR2X1   g00114(.A(new_n307_), .B(new_n306_), .Y(new_n308_));
  INVX1    g00115(.A(new_n308_), .Y(new_n309_));
  NAND3X1  g00116(.A(\a[8] ), .B(\a[5] ), .C(\a[1] ), .Y(new_n310_));
  AND2X1   g00117(.A(\a[8] ), .B(\a[1] ), .Y(new_n311_));
  OAI21X1  g00118(.A0(new_n311_), .A1(\a[5] ), .B0(new_n310_), .Y(new_n312_));
  XOR2X1   g00119(.A(new_n312_), .B(new_n309_), .Y(new_n313_));
  OAI21X1  g00120(.A0(new_n303_), .A1(new_n293_), .B0(new_n313_), .Y(new_n314_));
  OAI22X1  g00121(.A0(new_n314_), .A1(new_n304_), .B0(new_n313_), .B1(new_n305_), .Y(new_n315_));
  XOR2X1   g00122(.A(new_n315_), .B(new_n292_), .Y(new_n316_));
  OR2X1    g00123(.A(new_n283_), .B(new_n269_), .Y(new_n317_));
  AND2X1   g00124(.A(new_n283_), .B(new_n269_), .Y(new_n318_));
  AOI21X1  g00125(.A0(new_n289_), .A1(new_n317_), .B0(new_n318_), .Y(new_n319_));
  INVX1    g00126(.A(new_n319_), .Y(new_n320_));
  XOR2X1   g00127(.A(new_n320_), .B(new_n316_), .Y(\asquared[10] ));
  NOR2X1   g00128(.A(new_n313_), .B(new_n305_), .Y(new_n322_));
  AOI21X1  g00129(.A0(new_n303_), .A1(new_n281_), .B0(new_n322_), .Y(new_n323_));
  AND2X1   g00130(.A(\a[10] ), .B(\a[8] ), .Y(new_n324_));
  AND2X1   g00131(.A(\a[8] ), .B(\a[7] ), .Y(new_n325_));
  AOI22X1  g00132(.A0(new_n325_), .A1(new_n231_), .B0(new_n324_), .B1(new_n197_), .Y(new_n326_));
  NAND4X1  g00133(.A(\a[10] ), .B(\a[7] ), .C(\a[3] ), .D(\a[0] ), .Y(new_n327_));
  INVX1    g00134(.A(new_n327_), .Y(new_n328_));
  OR2X1    g00135(.A(new_n328_), .B(new_n326_), .Y(new_n329_));
  NAND3X1  g00136(.A(new_n329_), .B(\a[8] ), .C(\a[2] ), .Y(new_n330_));
  NAND2X1  g00137(.A(new_n327_), .B(new_n326_), .Y(new_n331_));
  AOI22X1  g00138(.A0(\a[10] ), .A1(\a[0] ), .B0(\a[7] ), .B1(\a[3] ), .Y(new_n332_));
  OR2X1    g00139(.A(new_n332_), .B(new_n331_), .Y(new_n333_));
  AND2X1   g00140(.A(new_n333_), .B(new_n330_), .Y(new_n334_));
  OR2X1    g00141(.A(new_n312_), .B(new_n308_), .Y(new_n335_));
  NAND3X1  g00142(.A(new_n307_), .B(new_n272_), .C(new_n271_), .Y(new_n336_));
  AND2X1   g00143(.A(new_n336_), .B(new_n335_), .Y(new_n337_));
  XOR2X1   g00144(.A(new_n337_), .B(new_n334_), .Y(new_n338_));
  NAND4X1  g00145(.A(\a[9] ), .B(\a[6] ), .C(\a[4] ), .D(\a[1] ), .Y(new_n339_));
  INVX1    g00146(.A(\a[4] ), .Y(new_n340_));
  INVX1    g00147(.A(\a[9] ), .Y(new_n341_));
  OAI22X1  g00148(.A0(new_n341_), .A1(new_n202_), .B0(new_n230_), .B1(new_n340_), .Y(new_n342_));
  NAND3X1  g00149(.A(new_n342_), .B(new_n339_), .C(new_n310_), .Y(new_n343_));
  NAND2X1  g00150(.A(new_n342_), .B(new_n339_), .Y(new_n344_));
  XOR2X1   g00151(.A(new_n344_), .B(new_n310_), .Y(new_n345_));
  AOI21X1  g00152(.A0(new_n342_), .A1(new_n339_), .B0(new_n310_), .Y(new_n346_));
  NOR2X1   g00153(.A(new_n346_), .B(new_n300_), .Y(new_n347_));
  AOI22X1  g00154(.A0(new_n347_), .A1(new_n343_), .B0(new_n345_), .B1(new_n300_), .Y(new_n348_));
  NAND2X1  g00155(.A(new_n348_), .B(new_n338_), .Y(new_n349_));
  OR2X1    g00156(.A(new_n348_), .B(new_n338_), .Y(new_n350_));
  NAND2X1  g00157(.A(new_n350_), .B(new_n349_), .Y(new_n351_));
  NOR2X1   g00158(.A(new_n351_), .B(new_n323_), .Y(new_n352_));
  INVX1    g00159(.A(new_n352_), .Y(new_n353_));
  OR2X1    g00160(.A(new_n315_), .B(new_n292_), .Y(new_n354_));
  AND2X1   g00161(.A(new_n315_), .B(new_n292_), .Y(new_n355_));
  OAI21X1  g00162(.A0(new_n319_), .A1(new_n355_), .B0(new_n354_), .Y(new_n356_));
  NAND2X1  g00163(.A(new_n351_), .B(new_n323_), .Y(new_n357_));
  AOI21X1  g00164(.A0(new_n353_), .A1(new_n357_), .B0(new_n356_), .Y(new_n358_));
  AND2X1   g00165(.A(new_n357_), .B(new_n356_), .Y(new_n359_));
  AOI21X1  g00166(.A0(new_n359_), .A1(new_n353_), .B0(new_n358_), .Y(\asquared[11] ));
  OAI21X1  g00167(.A0(new_n337_), .A1(new_n334_), .B0(new_n349_), .Y(new_n361_));
  NAND2X1  g00168(.A(\a[10] ), .B(\a[1] ), .Y(new_n362_));
  AOI22X1  g00169(.A0(new_n362_), .A1(new_n230_), .B0(new_n260_), .B1(\a[10] ), .Y(new_n363_));
  XOR2X1   g00170(.A(new_n363_), .B(new_n331_), .Y(new_n364_));
  AOI22X1  g00171(.A0(\a[9] ), .A1(\a[2] ), .B0(\a[8] ), .B1(\a[3] ), .Y(new_n365_));
  NAND2X1  g00172(.A(\a[9] ), .B(\a[8] ), .Y(new_n366_));
  NOR2X1   g00173(.A(new_n366_), .B(new_n249_), .Y(new_n367_));
  NOR3X1   g00174(.A(new_n365_), .B(new_n367_), .C(new_n339_), .Y(new_n368_));
  OAI22X1  g00175(.A0(new_n365_), .A1(new_n339_), .B0(new_n366_), .B1(new_n249_), .Y(new_n369_));
  OAI22X1  g00176(.A0(new_n369_), .A1(new_n365_), .B0(new_n368_), .B1(new_n339_), .Y(new_n370_));
  XOR2X1   g00177(.A(new_n370_), .B(new_n364_), .Y(new_n371_));
  NAND2X1  g00178(.A(new_n345_), .B(new_n300_), .Y(new_n372_));
  OAI21X1  g00179(.A0(new_n344_), .A1(new_n310_), .B0(new_n372_), .Y(new_n373_));
  AOI22X1  g00180(.A0(\a[7] ), .A1(\a[4] ), .B0(\a[6] ), .B1(\a[5] ), .Y(new_n374_));
  AND2X1   g00181(.A(\a[7] ), .B(\a[6] ), .Y(new_n375_));
  INVX1    g00182(.A(new_n375_), .Y(new_n376_));
  AND2X1   g00183(.A(\a[11] ), .B(\a[0] ), .Y(new_n377_));
  INVX1    g00184(.A(new_n377_), .Y(new_n378_));
  OAI22X1  g00185(.A0(new_n378_), .A1(new_n374_), .B0(new_n376_), .B1(new_n220_), .Y(new_n379_));
  AND2X1   g00186(.A(new_n375_), .B(new_n218_), .Y(new_n380_));
  OAI21X1  g00187(.A0(new_n380_), .A1(new_n374_), .B0(new_n377_), .Y(new_n381_));
  OAI21X1  g00188(.A0(new_n379_), .A1(new_n374_), .B0(new_n381_), .Y(new_n382_));
  INVX1    g00189(.A(new_n382_), .Y(new_n383_));
  OR2X1    g00190(.A(new_n383_), .B(new_n373_), .Y(new_n384_));
  XOR2X1   g00191(.A(new_n382_), .B(new_n373_), .Y(new_n385_));
  AOI21X1  g00192(.A0(new_n383_), .A1(new_n373_), .B0(new_n371_), .Y(new_n386_));
  AOI22X1  g00193(.A0(new_n386_), .A1(new_n384_), .B0(new_n385_), .B1(new_n371_), .Y(new_n387_));
  XOR2X1   g00194(.A(new_n387_), .B(new_n361_), .Y(new_n388_));
  AOI21X1  g00195(.A0(new_n357_), .A1(new_n356_), .B0(new_n352_), .Y(new_n389_));
  INVX1    g00196(.A(new_n389_), .Y(new_n390_));
  XOR2X1   g00197(.A(new_n390_), .B(new_n388_), .Y(\asquared[12] ));
  AND2X1   g00198(.A(new_n382_), .B(new_n373_), .Y(new_n392_));
  AND2X1   g00199(.A(new_n385_), .B(new_n371_), .Y(new_n393_));
  OR2X1    g00200(.A(new_n393_), .B(new_n392_), .Y(new_n394_));
  XOR2X1   g00201(.A(new_n379_), .B(new_n369_), .Y(new_n395_));
  AND2X1   g00202(.A(\a[12] ), .B(\a[10] ), .Y(new_n396_));
  NAND4X1  g00203(.A(\a[12] ), .B(\a[9] ), .C(\a[3] ), .D(\a[0] ), .Y(new_n397_));
  NAND4X1  g00204(.A(\a[10] ), .B(\a[9] ), .C(\a[3] ), .D(\a[2] ), .Y(new_n398_));
  AOI22X1  g00205(.A0(new_n398_), .A1(new_n397_), .B0(new_n396_), .B1(new_n197_), .Y(new_n399_));
  NOR3X1   g00206(.A(new_n399_), .B(new_n341_), .C(new_n223_), .Y(new_n400_));
  AOI21X1  g00207(.A0(new_n396_), .A1(new_n197_), .B0(new_n399_), .Y(new_n401_));
  AOI22X1  g00208(.A0(\a[12] ), .A1(\a[0] ), .B0(\a[10] ), .B1(\a[2] ), .Y(new_n402_));
  INVX1    g00209(.A(new_n402_), .Y(new_n403_));
  AOI21X1  g00210(.A0(new_n403_), .A1(new_n401_), .B0(new_n400_), .Y(new_n404_));
  XOR2X1   g00211(.A(new_n404_), .B(new_n395_), .Y(new_n405_));
  AND2X1   g00212(.A(new_n363_), .B(new_n331_), .Y(new_n406_));
  AOI21X1  g00213(.A0(new_n370_), .A1(new_n364_), .B0(new_n406_), .Y(new_n407_));
  AOI22X1  g00214(.A0(new_n260_), .A1(\a[10] ), .B0(\a[8] ), .B1(\a[4] ), .Y(new_n408_));
  AND2X1   g00215(.A(\a[11] ), .B(\a[5] ), .Y(new_n409_));
  AND2X1   g00216(.A(new_n409_), .B(new_n271_), .Y(new_n410_));
  AOI22X1  g00217(.A0(\a[11] ), .A1(\a[1] ), .B0(\a[7] ), .B1(\a[5] ), .Y(new_n411_));
  OR2X1    g00218(.A(new_n411_), .B(new_n410_), .Y(new_n412_));
  INVX1    g00219(.A(\a[8] ), .Y(new_n413_));
  NAND3X1  g00220(.A(\a[10] ), .B(\a[6] ), .C(\a[1] ), .Y(new_n414_));
  NOR3X1   g00221(.A(new_n414_), .B(new_n413_), .C(new_n340_), .Y(new_n415_));
  NOR4X1   g00222(.A(new_n411_), .B(new_n410_), .C(new_n415_), .D(new_n408_), .Y(new_n416_));
  OR2X1    g00223(.A(new_n416_), .B(new_n415_), .Y(new_n417_));
  OAI22X1  g00224(.A0(new_n417_), .A1(new_n408_), .B0(new_n416_), .B1(new_n412_), .Y(new_n418_));
  XOR2X1   g00225(.A(new_n418_), .B(new_n407_), .Y(new_n419_));
  XOR2X1   g00226(.A(new_n419_), .B(new_n405_), .Y(new_n420_));
  AND2X1   g00227(.A(new_n420_), .B(new_n394_), .Y(new_n421_));
  INVX1    g00228(.A(new_n421_), .Y(new_n422_));
  NOR2X1   g00229(.A(new_n387_), .B(new_n361_), .Y(new_n423_));
  NAND2X1  g00230(.A(new_n387_), .B(new_n361_), .Y(new_n424_));
  OAI21X1  g00231(.A0(new_n389_), .A1(new_n423_), .B0(new_n424_), .Y(new_n425_));
  OR2X1    g00232(.A(new_n420_), .B(new_n394_), .Y(new_n426_));
  AOI21X1  g00233(.A0(new_n422_), .A1(new_n426_), .B0(new_n425_), .Y(new_n427_));
  AND2X1   g00234(.A(new_n426_), .B(new_n425_), .Y(new_n428_));
  AOI21X1  g00235(.A0(new_n428_), .A1(new_n422_), .B0(new_n427_), .Y(\asquared[13] ));
  AND2X1   g00236(.A(\a[13] ), .B(\a[9] ), .Y(new_n430_));
  NAND4X1  g00237(.A(\a[10] ), .B(\a[9] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n431_));
  NAND4X1  g00238(.A(\a[13] ), .B(\a[10] ), .C(\a[3] ), .D(\a[0] ), .Y(new_n432_));
  AOI22X1  g00239(.A0(new_n432_), .A1(new_n431_), .B0(new_n430_), .B1(new_n210_), .Y(new_n433_));
  NAND2X1  g00240(.A(\a[10] ), .B(\a[3] ), .Y(new_n434_));
  NAND4X1  g00241(.A(\a[13] ), .B(\a[9] ), .C(\a[4] ), .D(\a[0] ), .Y(new_n435_));
  NAND3X1  g00242(.A(new_n432_), .B(new_n431_), .C(new_n435_), .Y(new_n436_));
  AOI22X1  g00243(.A0(\a[13] ), .A1(\a[0] ), .B0(\a[9] ), .B1(\a[4] ), .Y(new_n437_));
  OAI22X1  g00244(.A0(new_n437_), .A1(new_n436_), .B0(new_n434_), .B1(new_n433_), .Y(new_n438_));
  XOR2X1   g00245(.A(new_n438_), .B(new_n417_), .Y(new_n439_));
  NAND2X1  g00246(.A(\a[11] ), .B(\a[2] ), .Y(new_n440_));
  AOI22X1  g00247(.A0(\a[8] ), .A1(\a[5] ), .B0(\a[7] ), .B1(\a[6] ), .Y(new_n441_));
  AND2X1   g00248(.A(new_n325_), .B(new_n295_), .Y(new_n442_));
  NOR3X1   g00249(.A(new_n441_), .B(new_n442_), .C(new_n440_), .Y(new_n443_));
  INVX1    g00250(.A(new_n295_), .Y(new_n444_));
  INVX1    g00251(.A(new_n325_), .Y(new_n445_));
  OAI22X1  g00252(.A0(new_n441_), .A1(new_n440_), .B0(new_n445_), .B1(new_n444_), .Y(new_n446_));
  OAI22X1  g00253(.A0(new_n446_), .A1(new_n441_), .B0(new_n443_), .B1(new_n440_), .Y(new_n447_));
  XOR2X1   g00254(.A(new_n447_), .B(new_n439_), .Y(new_n448_));
  NAND2X1  g00255(.A(new_n379_), .B(new_n369_), .Y(new_n449_));
  AND2X1   g00256(.A(new_n403_), .B(new_n401_), .Y(new_n450_));
  OAI21X1  g00257(.A0(new_n450_), .A1(new_n400_), .B0(new_n395_), .Y(new_n451_));
  AND2X1   g00258(.A(new_n451_), .B(new_n449_), .Y(new_n452_));
  INVX1    g00259(.A(\a[12] ), .Y(new_n453_));
  NAND3X1  g00260(.A(new_n409_), .B(new_n271_), .C(new_n453_), .Y(new_n454_));
  AOI21X1  g00261(.A0(\a[12] ), .A1(\a[1] ), .B0(\a[7] ), .Y(new_n455_));
  AOI21X1  g00262(.A0(new_n271_), .A1(\a[12] ), .B0(new_n455_), .Y(new_n456_));
  OAI21X1  g00263(.A0(new_n456_), .A1(new_n410_), .B0(new_n454_), .Y(new_n457_));
  INVX1    g00264(.A(new_n457_), .Y(new_n458_));
  XOR2X1   g00265(.A(new_n458_), .B(new_n401_), .Y(new_n459_));
  XOR2X1   g00266(.A(new_n459_), .B(new_n452_), .Y(new_n460_));
  AND2X1   g00267(.A(new_n370_), .B(new_n364_), .Y(new_n461_));
  OAI21X1  g00268(.A0(new_n461_), .A1(new_n406_), .B0(new_n418_), .Y(new_n462_));
  OAI21X1  g00269(.A0(new_n419_), .A1(new_n405_), .B0(new_n462_), .Y(new_n463_));
  XOR2X1   g00270(.A(new_n463_), .B(new_n460_), .Y(new_n464_));
  NOR2X1   g00271(.A(new_n464_), .B(new_n448_), .Y(new_n465_));
  NAND2X1  g00272(.A(new_n464_), .B(new_n448_), .Y(new_n466_));
  INVX1    g00273(.A(new_n466_), .Y(new_n467_));
  OR2X1    g00274(.A(new_n467_), .B(new_n465_), .Y(new_n468_));
  AOI21X1  g00275(.A0(new_n426_), .A1(new_n425_), .B0(new_n421_), .Y(new_n469_));
  XOR2X1   g00276(.A(new_n469_), .B(new_n468_), .Y(\asquared[14] ));
  AOI21X1  g00277(.A0(new_n451_), .A1(new_n449_), .B0(new_n459_), .Y(new_n471_));
  AOI21X1  g00278(.A0(new_n463_), .A1(new_n460_), .B0(new_n471_), .Y(new_n472_));
  AND2X1   g00279(.A(\a[13] ), .B(\a[1] ), .Y(new_n473_));
  XOR2X1   g00280(.A(new_n473_), .B(new_n277_), .Y(new_n474_));
  INVX1    g00281(.A(new_n474_), .Y(new_n475_));
  XOR2X1   g00282(.A(new_n475_), .B(new_n446_), .Y(new_n476_));
  XOR2X1   g00283(.A(new_n476_), .B(new_n436_), .Y(new_n477_));
  INVX1    g00284(.A(new_n477_), .Y(new_n478_));
  AND2X1   g00285(.A(new_n438_), .B(new_n417_), .Y(new_n479_));
  AOI21X1  g00286(.A0(new_n447_), .A1(new_n439_), .B0(new_n479_), .Y(new_n480_));
  XOR2X1   g00287(.A(new_n480_), .B(new_n478_), .Y(new_n481_));
  AND2X1   g00288(.A(\a[12] ), .B(\a[11] ), .Y(new_n482_));
  AND2X1   g00289(.A(new_n482_), .B(new_n231_), .Y(new_n483_));
  NAND4X1  g00290(.A(\a[14] ), .B(\a[11] ), .C(\a[3] ), .D(\a[0] ), .Y(new_n484_));
  NAND4X1  g00291(.A(\a[14] ), .B(\a[12] ), .C(\a[2] ), .D(\a[0] ), .Y(new_n485_));
  AOI22X1  g00292(.A0(new_n485_), .A1(new_n484_), .B0(new_n482_), .B1(new_n231_), .Y(new_n486_));
  NOR2X1   g00293(.A(new_n486_), .B(new_n483_), .Y(new_n487_));
  INVX1    g00294(.A(\a[11] ), .Y(new_n488_));
  OAI22X1  g00295(.A0(new_n453_), .A1(new_n200_), .B0(new_n488_), .B1(new_n223_), .Y(new_n489_));
  INVX1    g00296(.A(\a[14] ), .Y(new_n490_));
  NOR3X1   g00297(.A(new_n486_), .B(new_n490_), .C(new_n194_), .Y(new_n491_));
  AOI21X1  g00298(.A0(new_n489_), .A1(new_n487_), .B0(new_n491_), .Y(new_n492_));
  NAND3X1  g00299(.A(\a[12] ), .B(\a[7] ), .C(\a[1] ), .Y(new_n493_));
  AOI22X1  g00300(.A0(\a[10] ), .A1(\a[4] ), .B0(\a[9] ), .B1(\a[5] ), .Y(new_n494_));
  INVX1    g00301(.A(new_n494_), .Y(new_n495_));
  NAND4X1  g00302(.A(\a[10] ), .B(\a[9] ), .C(\a[5] ), .D(\a[4] ), .Y(new_n496_));
  AOI21X1  g00303(.A0(new_n496_), .A1(new_n495_), .B0(new_n493_), .Y(new_n497_));
  OAI21X1  g00304(.A0(new_n494_), .A1(new_n493_), .B0(new_n496_), .Y(new_n498_));
  NOR2X1   g00305(.A(new_n498_), .B(new_n494_), .Y(new_n499_));
  NOR2X1   g00306(.A(new_n499_), .B(new_n497_), .Y(new_n500_));
  XOR2X1   g00307(.A(new_n500_), .B(new_n492_), .Y(new_n501_));
  OAI21X1  g00308(.A0(new_n457_), .A1(new_n401_), .B0(new_n454_), .Y(new_n502_));
  XOR2X1   g00309(.A(new_n502_), .B(new_n501_), .Y(new_n503_));
  XOR2X1   g00310(.A(new_n503_), .B(new_n481_), .Y(new_n504_));
  NOR2X1   g00311(.A(new_n504_), .B(new_n472_), .Y(new_n505_));
  INVX1    g00312(.A(new_n505_), .Y(new_n506_));
  OAI21X1  g00313(.A0(new_n469_), .A1(new_n465_), .B0(new_n466_), .Y(new_n507_));
  NAND2X1  g00314(.A(new_n504_), .B(new_n472_), .Y(new_n508_));
  AOI21X1  g00315(.A0(new_n508_), .A1(new_n506_), .B0(new_n507_), .Y(new_n509_));
  AND2X1   g00316(.A(new_n508_), .B(new_n507_), .Y(new_n510_));
  AOI21X1  g00317(.A0(new_n510_), .A1(new_n506_), .B0(new_n509_), .Y(\asquared[15] ));
  AOI21X1  g00318(.A0(new_n508_), .A1(new_n507_), .B0(new_n505_), .Y(new_n512_));
  NAND2X1  g00319(.A(new_n480_), .B(new_n477_), .Y(new_n513_));
  NOR2X1   g00320(.A(new_n480_), .B(new_n477_), .Y(new_n514_));
  AOI21X1  g00321(.A0(new_n503_), .A1(new_n513_), .B0(new_n514_), .Y(new_n515_));
  NAND4X1  g00322(.A(\a[13] ), .B(\a[8] ), .C(\a[6] ), .D(\a[1] ), .Y(new_n516_));
  NAND2X1  g00323(.A(\a[11] ), .B(\a[4] ), .Y(new_n517_));
  NAND2X1  g00324(.A(new_n517_), .B(new_n516_), .Y(new_n518_));
  AND2X1   g00325(.A(\a[14] ), .B(\a[1] ), .Y(new_n519_));
  XOR2X1   g00326(.A(new_n519_), .B(\a[8] ), .Y(new_n520_));
  XOR2X1   g00327(.A(new_n517_), .B(new_n516_), .Y(new_n521_));
  NAND2X1  g00328(.A(new_n521_), .B(new_n520_), .Y(new_n522_));
  NOR2X1   g00329(.A(new_n517_), .B(new_n516_), .Y(new_n523_));
  AOI21X1  g00330(.A0(new_n520_), .A1(new_n518_), .B0(new_n523_), .Y(new_n524_));
  AOI22X1  g00331(.A0(new_n524_), .A1(new_n518_), .B0(new_n522_), .B1(new_n520_), .Y(new_n525_));
  AOI22X1  g00332(.A0(\a[9] ), .A1(\a[6] ), .B0(\a[8] ), .B1(\a[7] ), .Y(new_n526_));
  INVX1    g00333(.A(new_n526_), .Y(new_n527_));
  AND2X1   g00334(.A(\a[13] ), .B(\a[2] ), .Y(new_n528_));
  INVX1    g00335(.A(new_n528_), .Y(new_n529_));
  NAND4X1  g00336(.A(\a[9] ), .B(\a[8] ), .C(\a[7] ), .D(\a[6] ), .Y(new_n530_));
  AOI21X1  g00337(.A0(new_n527_), .A1(new_n530_), .B0(new_n529_), .Y(new_n531_));
  INVX1    g00338(.A(\a[7] ), .Y(new_n532_));
  NOR4X1   g00339(.A(new_n341_), .B(new_n413_), .C(new_n532_), .D(new_n230_), .Y(new_n533_));
  AOI21X1  g00340(.A0(new_n527_), .A1(new_n528_), .B0(new_n533_), .Y(new_n534_));
  AOI21X1  g00341(.A0(new_n534_), .A1(new_n527_), .B0(new_n531_), .Y(new_n535_));
  XOR2X1   g00342(.A(new_n535_), .B(new_n525_), .Y(new_n536_));
  INVX1    g00343(.A(new_n436_), .Y(new_n537_));
  NAND2X1  g00344(.A(new_n474_), .B(new_n446_), .Y(new_n538_));
  OAI21X1  g00345(.A0(new_n476_), .A1(new_n537_), .B0(new_n538_), .Y(new_n539_));
  XOR2X1   g00346(.A(new_n539_), .B(new_n536_), .Y(new_n540_));
  XOR2X1   g00347(.A(new_n498_), .B(new_n487_), .Y(new_n541_));
  AND2X1   g00348(.A(\a[10] ), .B(\a[5] ), .Y(new_n542_));
  INVX1    g00349(.A(new_n396_), .Y(new_n543_));
  NAND2X1  g00350(.A(\a[15] ), .B(\a[10] ), .Y(new_n544_));
  OAI22X1  g00351(.A0(new_n544_), .A1(new_n194_), .B0(new_n543_), .B1(new_n223_), .Y(new_n545_));
  NAND4X1  g00352(.A(\a[15] ), .B(\a[12] ), .C(\a[3] ), .D(\a[0] ), .Y(new_n546_));
  NAND3X1  g00353(.A(new_n546_), .B(new_n545_), .C(\a[5] ), .Y(new_n547_));
  AND2X1   g00354(.A(new_n547_), .B(new_n546_), .Y(new_n548_));
  INVX1    g00355(.A(\a[15] ), .Y(new_n549_));
  OAI22X1  g00356(.A0(new_n549_), .A1(new_n194_), .B0(new_n453_), .B1(new_n223_), .Y(new_n550_));
  AOI22X1  g00357(.A0(new_n550_), .A1(new_n548_), .B0(new_n547_), .B1(new_n542_), .Y(new_n551_));
  XOR2X1   g00358(.A(new_n551_), .B(new_n541_), .Y(new_n552_));
  NAND2X1  g00359(.A(new_n502_), .B(new_n501_), .Y(new_n553_));
  OAI21X1  g00360(.A0(new_n500_), .A1(new_n492_), .B0(new_n553_), .Y(new_n554_));
  XOR2X1   g00361(.A(new_n554_), .B(new_n552_), .Y(new_n555_));
  XOR2X1   g00362(.A(new_n555_), .B(new_n540_), .Y(new_n556_));
  XOR2X1   g00363(.A(new_n556_), .B(new_n515_), .Y(new_n557_));
  XOR2X1   g00364(.A(new_n557_), .B(new_n512_), .Y(\asquared[16] ));
  AND2X1   g00365(.A(new_n554_), .B(new_n552_), .Y(new_n559_));
  AOI21X1  g00366(.A0(new_n555_), .A1(new_n540_), .B0(new_n559_), .Y(new_n560_));
  OAI21X1  g00367(.A0(new_n517_), .A1(new_n516_), .B0(new_n522_), .Y(new_n561_));
  XOR2X1   g00368(.A(new_n548_), .B(new_n561_), .Y(new_n562_));
  AND2X1   g00369(.A(\a[10] ), .B(\a[0] ), .Y(new_n563_));
  AND2X1   g00370(.A(\a[16] ), .B(\a[6] ), .Y(new_n564_));
  NAND4X1  g00371(.A(\a[11] ), .B(\a[10] ), .C(\a[6] ), .D(\a[5] ), .Y(new_n565_));
  NAND4X1  g00372(.A(\a[16] ), .B(\a[11] ), .C(\a[5] ), .D(\a[0] ), .Y(new_n566_));
  AOI22X1  g00373(.A0(new_n566_), .A1(new_n565_), .B0(new_n564_), .B1(new_n563_), .Y(new_n567_));
  NOR3X1   g00374(.A(new_n567_), .B(new_n488_), .C(new_n255_), .Y(new_n568_));
  AOI21X1  g00375(.A0(new_n564_), .A1(new_n563_), .B0(new_n567_), .Y(new_n569_));
  INVX1    g00376(.A(\a[10] ), .Y(new_n570_));
  INVX1    g00377(.A(\a[16] ), .Y(new_n571_));
  OAI22X1  g00378(.A0(new_n571_), .A1(new_n194_), .B0(new_n570_), .B1(new_n230_), .Y(new_n572_));
  AOI21X1  g00379(.A0(new_n572_), .A1(new_n569_), .B0(new_n568_), .Y(new_n573_));
  XOR2X1   g00380(.A(new_n573_), .B(new_n562_), .Y(new_n574_));
  INVX1    g00381(.A(new_n574_), .Y(new_n575_));
  NOR2X1   g00382(.A(new_n535_), .B(new_n525_), .Y(new_n576_));
  AOI21X1  g00383(.A0(new_n539_), .A1(new_n536_), .B0(new_n576_), .Y(new_n577_));
  XOR2X1   g00384(.A(new_n577_), .B(new_n575_), .Y(new_n578_));
  OAI21X1  g00385(.A0(new_n486_), .A1(new_n483_), .B0(new_n498_), .Y(new_n579_));
  OAI21X1  g00386(.A0(new_n551_), .A1(new_n541_), .B0(new_n579_), .Y(new_n580_));
  AND2X1   g00387(.A(\a[12] ), .B(\a[4] ), .Y(new_n581_));
  AND2X1   g00388(.A(\a[14] ), .B(\a[13] ), .Y(new_n582_));
  INVX1    g00389(.A(new_n582_), .Y(new_n583_));
  INVX1    g00390(.A(new_n235_), .Y(new_n584_));
  NAND2X1  g00391(.A(\a[14] ), .B(\a[12] ), .Y(new_n585_));
  AND2X1   g00392(.A(\a[13] ), .B(\a[12] ), .Y(new_n586_));
  INVX1    g00393(.A(new_n586_), .Y(new_n587_));
  OAI22X1  g00394(.A0(new_n587_), .A1(new_n217_), .B0(new_n585_), .B1(new_n584_), .Y(new_n588_));
  OAI21X1  g00395(.A0(new_n583_), .A1(new_n249_), .B0(new_n588_), .Y(new_n589_));
  AOI21X1  g00396(.A0(new_n582_), .A1(new_n231_), .B0(new_n588_), .Y(new_n590_));
  INVX1    g00397(.A(\a[13] ), .Y(new_n591_));
  OAI22X1  g00398(.A0(new_n490_), .A1(new_n200_), .B0(new_n591_), .B1(new_n223_), .Y(new_n592_));
  AOI22X1  g00399(.A0(new_n592_), .A1(new_n590_), .B0(new_n589_), .B1(new_n581_), .Y(new_n593_));
  XOR2X1   g00400(.A(new_n593_), .B(new_n580_), .Y(new_n594_));
  NAND3X1  g00401(.A(\a[14] ), .B(\a[8] ), .C(\a[1] ), .Y(new_n595_));
  AND2X1   g00402(.A(\a[9] ), .B(\a[7] ), .Y(new_n596_));
  AND2X1   g00403(.A(\a[15] ), .B(\a[1] ), .Y(new_n597_));
  XOR2X1   g00404(.A(new_n597_), .B(new_n596_), .Y(new_n598_));
  XOR2X1   g00405(.A(new_n598_), .B(new_n595_), .Y(new_n599_));
  XOR2X1   g00406(.A(new_n599_), .B(new_n534_), .Y(new_n600_));
  XOR2X1   g00407(.A(new_n600_), .B(new_n594_), .Y(new_n601_));
  XOR2X1   g00408(.A(new_n601_), .B(new_n578_), .Y(new_n602_));
  XOR2X1   g00409(.A(new_n602_), .B(new_n560_), .Y(new_n603_));
  INVX1    g00410(.A(new_n540_), .Y(new_n604_));
  XOR2X1   g00411(.A(new_n555_), .B(new_n604_), .Y(new_n605_));
  OR2X1    g00412(.A(new_n605_), .B(new_n515_), .Y(new_n606_));
  AND2X1   g00413(.A(new_n605_), .B(new_n515_), .Y(new_n607_));
  OAI21X1  g00414(.A0(new_n607_), .A1(new_n512_), .B0(new_n606_), .Y(new_n608_));
  XOR2X1   g00415(.A(new_n608_), .B(new_n603_), .Y(\asquared[17] ));
  AND2X1   g00416(.A(new_n577_), .B(new_n575_), .Y(new_n610_));
  OR2X1    g00417(.A(new_n577_), .B(new_n575_), .Y(new_n611_));
  OAI21X1  g00418(.A0(new_n601_), .A1(new_n610_), .B0(new_n611_), .Y(new_n612_));
  AND2X1   g00419(.A(new_n597_), .B(new_n596_), .Y(new_n613_));
  INVX1    g00420(.A(new_n613_), .Y(new_n614_));
  AOI22X1  g00421(.A0(\a[17] ), .A1(\a[0] ), .B0(\a[12] ), .B1(\a[5] ), .Y(new_n615_));
  INVX1    g00422(.A(\a[17] ), .Y(new_n616_));
  NOR4X1   g00423(.A(new_n616_), .B(new_n453_), .C(new_n255_), .D(new_n194_), .Y(new_n617_));
  NOR3X1   g00424(.A(new_n617_), .B(new_n615_), .C(new_n614_), .Y(new_n618_));
  NOR2X1   g00425(.A(new_n618_), .B(new_n617_), .Y(new_n619_));
  INVX1    g00426(.A(new_n619_), .Y(new_n620_));
  OAI22X1  g00427(.A0(new_n620_), .A1(new_n615_), .B0(new_n618_), .B1(new_n614_), .Y(new_n621_));
  AOI22X1  g00428(.A0(\a[10] ), .A1(\a[7] ), .B0(\a[9] ), .B1(\a[8] ), .Y(new_n622_));
  INVX1    g00429(.A(new_n622_), .Y(new_n623_));
  NAND2X1  g00430(.A(\a[14] ), .B(\a[3] ), .Y(new_n624_));
  NAND4X1  g00431(.A(\a[10] ), .B(\a[9] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n625_));
  AOI21X1  g00432(.A0(new_n623_), .A1(new_n625_), .B0(new_n624_), .Y(new_n626_));
  OR2X1    g00433(.A(new_n622_), .B(new_n624_), .Y(new_n627_));
  AND2X1   g00434(.A(new_n627_), .B(new_n625_), .Y(new_n628_));
  AOI21X1  g00435(.A0(new_n628_), .A1(new_n623_), .B0(new_n626_), .Y(new_n629_));
  XOR2X1   g00436(.A(new_n629_), .B(new_n621_), .Y(new_n630_));
  INVX1    g00437(.A(new_n630_), .Y(new_n631_));
  AND2X1   g00438(.A(\a[11] ), .B(\a[6] ), .Y(new_n632_));
  NAND2X1  g00439(.A(\a[15] ), .B(\a[11] ), .Y(new_n633_));
  AND2X1   g00440(.A(\a[13] ), .B(\a[11] ), .Y(new_n634_));
  INVX1    g00441(.A(new_n634_), .Y(new_n635_));
  OAI22X1  g00442(.A0(new_n635_), .A1(new_n340_), .B0(new_n633_), .B1(new_n200_), .Y(new_n636_));
  NAND4X1  g00443(.A(\a[15] ), .B(\a[13] ), .C(\a[4] ), .D(\a[2] ), .Y(new_n637_));
  NAND3X1  g00444(.A(new_n637_), .B(new_n636_), .C(\a[6] ), .Y(new_n638_));
  AND2X1   g00445(.A(\a[15] ), .B(\a[13] ), .Y(new_n639_));
  AOI22X1  g00446(.A0(new_n639_), .A1(new_n235_), .B0(new_n636_), .B1(\a[6] ), .Y(new_n640_));
  OAI22X1  g00447(.A0(new_n549_), .A1(new_n200_), .B0(new_n591_), .B1(new_n340_), .Y(new_n641_));
  AOI22X1  g00448(.A0(new_n641_), .A1(new_n640_), .B0(new_n638_), .B1(new_n632_), .Y(new_n642_));
  XOR2X1   g00449(.A(new_n642_), .B(new_n631_), .Y(new_n643_));
  OR2X1    g00450(.A(new_n551_), .B(new_n541_), .Y(new_n644_));
  AOI21X1  g00451(.A0(new_n644_), .A1(new_n579_), .B0(new_n593_), .Y(new_n645_));
  INVX1    g00452(.A(new_n600_), .Y(new_n646_));
  NOR2X1   g00453(.A(new_n646_), .B(new_n594_), .Y(new_n647_));
  NOR2X1   g00454(.A(new_n647_), .B(new_n645_), .Y(new_n648_));
  XOR2X1   g00455(.A(new_n648_), .B(new_n643_), .Y(new_n649_));
  NAND3X1  g00456(.A(new_n598_), .B(new_n519_), .C(\a[8] ), .Y(new_n650_));
  OAI21X1  g00457(.A0(new_n599_), .A1(new_n534_), .B0(new_n650_), .Y(new_n651_));
  INVX1    g00458(.A(new_n651_), .Y(new_n652_));
  OR2X1    g00459(.A(new_n548_), .B(new_n524_), .Y(new_n653_));
  OAI21X1  g00460(.A0(new_n573_), .A1(new_n562_), .B0(new_n653_), .Y(new_n654_));
  XOR2X1   g00461(.A(new_n654_), .B(new_n652_), .Y(new_n655_));
  AOI21X1  g00462(.A0(\a[16] ), .A1(\a[1] ), .B0(\a[9] ), .Y(new_n656_));
  AND2X1   g00463(.A(\a[16] ), .B(\a[9] ), .Y(new_n657_));
  AOI21X1  g00464(.A0(new_n657_), .A1(\a[1] ), .B0(new_n656_), .Y(new_n658_));
  XOR2X1   g00465(.A(new_n658_), .B(new_n590_), .Y(new_n659_));
  INVX1    g00466(.A(new_n659_), .Y(new_n660_));
  XOR2X1   g00467(.A(new_n660_), .B(new_n569_), .Y(new_n661_));
  XOR2X1   g00468(.A(new_n661_), .B(new_n655_), .Y(new_n662_));
  XOR2X1   g00469(.A(new_n662_), .B(new_n649_), .Y(new_n663_));
  NAND2X1  g00470(.A(new_n663_), .B(new_n612_), .Y(new_n664_));
  INVX1    g00471(.A(new_n664_), .Y(new_n665_));
  NOR2X1   g00472(.A(new_n663_), .B(new_n612_), .Y(new_n666_));
  OR2X1    g00473(.A(new_n666_), .B(new_n665_), .Y(new_n667_));
  NOR2X1   g00474(.A(new_n602_), .B(new_n560_), .Y(new_n668_));
  AND2X1   g00475(.A(new_n602_), .B(new_n560_), .Y(new_n669_));
  INVX1    g00476(.A(new_n669_), .Y(new_n670_));
  AOI21X1  g00477(.A0(new_n608_), .A1(new_n670_), .B0(new_n668_), .Y(new_n671_));
  XOR2X1   g00478(.A(new_n671_), .B(new_n667_), .Y(\asquared[18] ));
  NOR2X1   g00479(.A(new_n648_), .B(new_n643_), .Y(new_n673_));
  AOI21X1  g00480(.A0(new_n662_), .A1(new_n649_), .B0(new_n673_), .Y(new_n674_));
  INVX1    g00481(.A(\a[18] ), .Y(new_n675_));
  NOR4X1   g00482(.A(new_n675_), .B(new_n591_), .C(new_n255_), .D(new_n194_), .Y(new_n676_));
  AND2X1   g00483(.A(\a[18] ), .B(\a[7] ), .Y(new_n677_));
  NAND2X1  g00484(.A(\a[7] ), .B(\a[5] ), .Y(new_n678_));
  NOR3X1   g00485(.A(new_n678_), .B(new_n591_), .C(new_n488_), .Y(new_n679_));
  AOI21X1  g00486(.A0(new_n677_), .A1(new_n377_), .B0(new_n679_), .Y(new_n680_));
  NOR2X1   g00487(.A(new_n680_), .B(new_n676_), .Y(new_n681_));
  INVX1    g00488(.A(new_n676_), .Y(new_n682_));
  AND2X1   g00489(.A(new_n680_), .B(new_n682_), .Y(new_n683_));
  INVX1    g00490(.A(new_n683_), .Y(new_n684_));
  AOI22X1  g00491(.A0(\a[18] ), .A1(\a[0] ), .B0(\a[13] ), .B1(\a[5] ), .Y(new_n685_));
  NAND2X1  g00492(.A(\a[11] ), .B(\a[7] ), .Y(new_n686_));
  OAI22X1  g00493(.A0(new_n686_), .A1(new_n681_), .B0(new_n685_), .B1(new_n684_), .Y(new_n687_));
  NAND2X1  g00494(.A(\a[14] ), .B(\a[4] ), .Y(new_n688_));
  AND2X1   g00495(.A(\a[16] ), .B(\a[15] ), .Y(new_n689_));
  AND2X1   g00496(.A(\a[16] ), .B(\a[14] ), .Y(new_n690_));
  AND2X1   g00497(.A(\a[15] ), .B(\a[14] ), .Y(new_n691_));
  AOI22X1  g00498(.A0(new_n691_), .A1(new_n294_), .B0(new_n690_), .B1(new_n235_), .Y(new_n692_));
  AOI21X1  g00499(.A0(new_n689_), .A1(new_n231_), .B0(new_n692_), .Y(new_n693_));
  AOI21X1  g00500(.A0(new_n689_), .A1(new_n231_), .B0(new_n693_), .Y(new_n694_));
  INVX1    g00501(.A(new_n694_), .Y(new_n695_));
  AOI22X1  g00502(.A0(\a[16] ), .A1(\a[2] ), .B0(\a[15] ), .B1(\a[3] ), .Y(new_n696_));
  OAI22X1  g00503(.A0(new_n696_), .A1(new_n695_), .B0(new_n693_), .B1(new_n688_), .Y(new_n697_));
  XOR2X1   g00504(.A(new_n697_), .B(new_n687_), .Y(new_n698_));
  INVX1    g00505(.A(new_n324_), .Y(new_n699_));
  AND2X1   g00506(.A(\a[17] ), .B(\a[1] ), .Y(new_n700_));
  XOR2X1   g00507(.A(new_n700_), .B(new_n699_), .Y(new_n701_));
  AOI22X1  g00508(.A0(new_n657_), .A1(\a[1] ), .B0(\a[12] ), .B1(\a[6] ), .Y(new_n702_));
  NAND4X1  g00509(.A(new_n657_), .B(\a[12] ), .C(\a[6] ), .D(\a[1] ), .Y(new_n703_));
  INVX1    g00510(.A(new_n703_), .Y(new_n704_));
  NOR3X1   g00511(.A(new_n704_), .B(new_n702_), .C(new_n701_), .Y(new_n705_));
  OAI21X1  g00512(.A0(new_n702_), .A1(new_n701_), .B0(new_n703_), .Y(new_n706_));
  OAI22X1  g00513(.A0(new_n706_), .A1(new_n702_), .B0(new_n705_), .B1(new_n701_), .Y(new_n707_));
  XOR2X1   g00514(.A(new_n707_), .B(new_n698_), .Y(new_n708_));
  NOR2X1   g00515(.A(new_n661_), .B(new_n655_), .Y(new_n709_));
  AOI21X1  g00516(.A0(new_n654_), .A1(new_n651_), .B0(new_n709_), .Y(new_n710_));
  XOR2X1   g00517(.A(new_n710_), .B(new_n708_), .Y(new_n711_));
  XOR2X1   g00518(.A(new_n640_), .B(new_n628_), .Y(new_n712_));
  XOR2X1   g00519(.A(new_n712_), .B(new_n620_), .Y(new_n713_));
  AND2X1   g00520(.A(new_n582_), .B(new_n231_), .Y(new_n714_));
  OAI21X1  g00521(.A0(new_n588_), .A1(new_n714_), .B0(new_n658_), .Y(new_n715_));
  OAI21X1  g00522(.A0(new_n659_), .A1(new_n569_), .B0(new_n715_), .Y(new_n716_));
  INVX1    g00523(.A(new_n621_), .Y(new_n717_));
  OR2X1    g00524(.A(new_n642_), .B(new_n630_), .Y(new_n718_));
  OAI21X1  g00525(.A0(new_n629_), .A1(new_n717_), .B0(new_n718_), .Y(new_n719_));
  XOR2X1   g00526(.A(new_n719_), .B(new_n716_), .Y(new_n720_));
  XOR2X1   g00527(.A(new_n720_), .B(new_n713_), .Y(new_n721_));
  XOR2X1   g00528(.A(new_n721_), .B(new_n711_), .Y(new_n722_));
  NOR2X1   g00529(.A(new_n722_), .B(new_n674_), .Y(new_n723_));
  INVX1    g00530(.A(new_n723_), .Y(new_n724_));
  OAI21X1  g00531(.A0(new_n671_), .A1(new_n666_), .B0(new_n664_), .Y(new_n725_));
  AND2X1   g00532(.A(new_n722_), .B(new_n674_), .Y(new_n726_));
  INVX1    g00533(.A(new_n726_), .Y(new_n727_));
  AOI21X1  g00534(.A0(new_n727_), .A1(new_n724_), .B0(new_n725_), .Y(new_n728_));
  AND2X1   g00535(.A(new_n727_), .B(new_n725_), .Y(new_n729_));
  AOI21X1  g00536(.A0(new_n729_), .A1(new_n724_), .B0(new_n728_), .Y(\asquared[19] ));
  XOR2X1   g00537(.A(new_n706_), .B(new_n683_), .Y(new_n731_));
  AND2X1   g00538(.A(\a[16] ), .B(\a[3] ), .Y(new_n732_));
  AOI22X1  g00539(.A0(\a[11] ), .A1(\a[8] ), .B0(\a[10] ), .B1(\a[9] ), .Y(new_n733_));
  INVX1    g00540(.A(new_n733_), .Y(new_n734_));
  NAND2X1  g00541(.A(\a[10] ), .B(\a[9] ), .Y(new_n735_));
  NOR3X1   g00542(.A(new_n735_), .B(new_n488_), .C(new_n413_), .Y(new_n736_));
  OR4X1    g00543(.A(new_n733_), .B(new_n736_), .C(new_n571_), .D(new_n223_), .Y(new_n737_));
  AOI21X1  g00544(.A0(new_n734_), .A1(new_n732_), .B0(new_n736_), .Y(new_n738_));
  AOI22X1  g00545(.A0(new_n738_), .A1(new_n734_), .B0(new_n737_), .B1(new_n732_), .Y(new_n739_));
  XOR2X1   g00546(.A(new_n739_), .B(new_n731_), .Y(new_n740_));
  AND2X1   g00547(.A(new_n697_), .B(new_n687_), .Y(new_n741_));
  AOI21X1  g00548(.A0(new_n707_), .A1(new_n698_), .B0(new_n741_), .Y(new_n742_));
  AND2X1   g00549(.A(new_n700_), .B(new_n324_), .Y(new_n743_));
  NAND4X1  g00550(.A(new_n324_), .B(new_n675_), .C(\a[17] ), .D(\a[1] ), .Y(new_n744_));
  AND2X1   g00551(.A(\a[18] ), .B(\a[1] ), .Y(new_n745_));
  XOR2X1   g00552(.A(new_n745_), .B(\a[10] ), .Y(new_n746_));
  OAI21X1  g00553(.A0(new_n746_), .A1(new_n743_), .B0(new_n744_), .Y(new_n747_));
  XOR2X1   g00554(.A(new_n747_), .B(new_n695_), .Y(new_n748_));
  XOR2X1   g00555(.A(new_n748_), .B(new_n742_), .Y(new_n749_));
  XOR2X1   g00556(.A(new_n749_), .B(new_n740_), .Y(new_n750_));
  INVX1    g00557(.A(new_n750_), .Y(new_n751_));
  INVX1    g00558(.A(\a[19] ), .Y(new_n752_));
  AND2X1   g00559(.A(\a[17] ), .B(\a[15] ), .Y(new_n753_));
  AND2X1   g00560(.A(new_n753_), .B(new_n235_), .Y(new_n754_));
  AOI22X1  g00561(.A0(new_n210_), .A1(\a[15] ), .B0(new_n197_), .B1(\a[17] ), .Y(new_n755_));
  NOR3X1   g00562(.A(new_n755_), .B(new_n754_), .C(new_n752_), .Y(new_n756_));
  NOR2X1   g00563(.A(new_n756_), .B(new_n754_), .Y(new_n757_));
  INVX1    g00564(.A(new_n757_), .Y(new_n758_));
  AOI22X1  g00565(.A0(\a[17] ), .A1(\a[2] ), .B0(\a[15] ), .B1(\a[4] ), .Y(new_n759_));
  AND2X1   g00566(.A(\a[19] ), .B(\a[0] ), .Y(new_n760_));
  INVX1    g00567(.A(new_n760_), .Y(new_n761_));
  OAI22X1  g00568(.A0(new_n761_), .A1(new_n756_), .B0(new_n759_), .B1(new_n758_), .Y(new_n762_));
  OAI22X1  g00569(.A0(new_n583_), .A1(new_n444_), .B0(new_n585_), .B1(new_n678_), .Y(new_n763_));
  OAI21X1  g00570(.A0(new_n587_), .A1(new_n376_), .B0(new_n763_), .Y(new_n764_));
  AND2X1   g00571(.A(\a[14] ), .B(\a[5] ), .Y(new_n765_));
  AOI21X1  g00572(.A0(new_n586_), .A1(new_n375_), .B0(new_n763_), .Y(new_n766_));
  OAI22X1  g00573(.A0(new_n591_), .A1(new_n230_), .B0(new_n453_), .B1(new_n532_), .Y(new_n767_));
  AOI22X1  g00574(.A0(new_n767_), .A1(new_n766_), .B0(new_n765_), .B1(new_n764_), .Y(new_n768_));
  XOR2X1   g00575(.A(new_n768_), .B(new_n762_), .Y(new_n769_));
  INVX1    g00576(.A(new_n769_), .Y(new_n770_));
  NOR2X1   g00577(.A(new_n640_), .B(new_n628_), .Y(new_n771_));
  AOI21X1  g00578(.A0(new_n712_), .A1(new_n620_), .B0(new_n771_), .Y(new_n772_));
  XOR2X1   g00579(.A(new_n772_), .B(new_n770_), .Y(new_n773_));
  AND2X1   g00580(.A(new_n719_), .B(new_n716_), .Y(new_n774_));
  AOI21X1  g00581(.A0(new_n720_), .A1(new_n713_), .B0(new_n774_), .Y(new_n775_));
  XOR2X1   g00582(.A(new_n775_), .B(new_n773_), .Y(new_n776_));
  XOR2X1   g00583(.A(new_n776_), .B(new_n751_), .Y(new_n777_));
  INVX1    g00584(.A(new_n708_), .Y(new_n778_));
  NOR2X1   g00585(.A(new_n710_), .B(new_n778_), .Y(new_n779_));
  INVX1    g00586(.A(new_n711_), .Y(new_n780_));
  AOI21X1  g00587(.A0(new_n721_), .A1(new_n780_), .B0(new_n779_), .Y(new_n781_));
  AND2X1   g00588(.A(new_n781_), .B(new_n777_), .Y(new_n782_));
  NOR2X1   g00589(.A(new_n781_), .B(new_n777_), .Y(new_n783_));
  OR2X1    g00590(.A(new_n783_), .B(new_n782_), .Y(new_n784_));
  AOI21X1  g00591(.A0(new_n727_), .A1(new_n725_), .B0(new_n723_), .Y(new_n785_));
  XOR2X1   g00592(.A(new_n785_), .B(new_n784_), .Y(\asquared[20] ));
  INVX1    g00593(.A(new_n783_), .Y(new_n787_));
  OAI21X1  g00594(.A0(new_n785_), .A1(new_n782_), .B0(new_n787_), .Y(new_n788_));
  NOR2X1   g00595(.A(new_n775_), .B(new_n773_), .Y(new_n789_));
  AOI21X1  g00596(.A0(new_n776_), .A1(new_n750_), .B0(new_n789_), .Y(new_n790_));
  OAI21X1  g00597(.A0(new_n747_), .A1(new_n694_), .B0(new_n744_), .Y(new_n791_));
  AND2X1   g00598(.A(\a[17] ), .B(\a[16] ), .Y(new_n792_));
  INVX1    g00599(.A(new_n792_), .Y(new_n793_));
  AND2X1   g00600(.A(\a[18] ), .B(\a[16] ), .Y(new_n794_));
  INVX1    g00601(.A(new_n794_), .Y(new_n795_));
  AND2X1   g00602(.A(\a[18] ), .B(\a[17] ), .Y(new_n796_));
  INVX1    g00603(.A(new_n796_), .Y(new_n797_));
  OAI22X1  g00604(.A0(new_n797_), .A1(new_n249_), .B0(new_n795_), .B1(new_n584_), .Y(new_n798_));
  OAI21X1  g00605(.A0(new_n793_), .A1(new_n217_), .B0(new_n798_), .Y(new_n799_));
  AND2X1   g00606(.A(\a[18] ), .B(\a[2] ), .Y(new_n800_));
  AOI21X1  g00607(.A0(new_n792_), .A1(new_n294_), .B0(new_n798_), .Y(new_n801_));
  OAI22X1  g00608(.A0(new_n616_), .A1(new_n223_), .B0(new_n571_), .B1(new_n340_), .Y(new_n802_));
  AOI22X1  g00609(.A0(new_n802_), .A1(new_n801_), .B0(new_n800_), .B1(new_n799_), .Y(new_n803_));
  XOR2X1   g00610(.A(new_n803_), .B(new_n791_), .Y(new_n804_));
  NOR2X1   g00611(.A(new_n739_), .B(new_n731_), .Y(new_n805_));
  AOI21X1  g00612(.A0(new_n706_), .A1(new_n684_), .B0(new_n805_), .Y(new_n806_));
  XOR2X1   g00613(.A(new_n806_), .B(new_n804_), .Y(new_n807_));
  INVX1    g00614(.A(new_n807_), .Y(new_n808_));
  NOR2X1   g00615(.A(new_n748_), .B(new_n742_), .Y(new_n809_));
  AOI21X1  g00616(.A0(new_n749_), .A1(new_n740_), .B0(new_n809_), .Y(new_n810_));
  XOR2X1   g00617(.A(new_n810_), .B(new_n808_), .Y(new_n811_));
  INVX1    g00618(.A(new_n811_), .Y(new_n812_));
  AND2X1   g00619(.A(\a[11] ), .B(\a[9] ), .Y(new_n813_));
  AND2X1   g00620(.A(\a[19] ), .B(\a[1] ), .Y(new_n814_));
  XOR2X1   g00621(.A(new_n814_), .B(new_n813_), .Y(new_n815_));
  XOR2X1   g00622(.A(new_n815_), .B(new_n738_), .Y(new_n816_));
  XOR2X1   g00623(.A(new_n816_), .B(new_n758_), .Y(new_n817_));
  INVX1    g00624(.A(new_n817_), .Y(new_n818_));
  INVX1    g00625(.A(new_n762_), .Y(new_n819_));
  OR2X1    g00626(.A(new_n768_), .B(new_n819_), .Y(new_n820_));
  OR2X1    g00627(.A(new_n772_), .B(new_n769_), .Y(new_n821_));
  AND2X1   g00628(.A(new_n821_), .B(new_n820_), .Y(new_n822_));
  XOR2X1   g00629(.A(new_n822_), .B(new_n818_), .Y(new_n823_));
  AND2X1   g00630(.A(new_n745_), .B(\a[10] ), .Y(new_n824_));
  AND2X1   g00631(.A(\a[20] ), .B(\a[0] ), .Y(new_n825_));
  AND2X1   g00632(.A(\a[13] ), .B(\a[7] ), .Y(new_n826_));
  XOR2X1   g00633(.A(new_n826_), .B(new_n825_), .Y(new_n827_));
  XOR2X1   g00634(.A(new_n827_), .B(new_n824_), .Y(new_n828_));
  INVX1    g00635(.A(new_n828_), .Y(new_n829_));
  XOR2X1   g00636(.A(new_n829_), .B(new_n766_), .Y(new_n830_));
  NAND4X1  g00637(.A(\a[14] ), .B(\a[12] ), .C(\a[8] ), .D(\a[6] ), .Y(new_n831_));
  NAND4X1  g00638(.A(\a[15] ), .B(\a[12] ), .C(\a[8] ), .D(\a[5] ), .Y(new_n832_));
  AOI22X1  g00639(.A0(new_n832_), .A1(new_n831_), .B0(new_n691_), .B1(new_n295_), .Y(new_n833_));
  NOR3X1   g00640(.A(new_n833_), .B(new_n453_), .C(new_n413_), .Y(new_n834_));
  AOI21X1  g00641(.A0(new_n691_), .A1(new_n295_), .B0(new_n833_), .Y(new_n835_));
  OAI22X1  g00642(.A0(new_n549_), .A1(new_n255_), .B0(new_n490_), .B1(new_n230_), .Y(new_n836_));
  AOI21X1  g00643(.A0(new_n836_), .A1(new_n835_), .B0(new_n834_), .Y(new_n837_));
  XOR2X1   g00644(.A(new_n837_), .B(new_n830_), .Y(new_n838_));
  XOR2X1   g00645(.A(new_n838_), .B(new_n823_), .Y(new_n839_));
  XOR2X1   g00646(.A(new_n839_), .B(new_n812_), .Y(new_n840_));
  XOR2X1   g00647(.A(new_n840_), .B(new_n790_), .Y(new_n841_));
  XOR2X1   g00648(.A(new_n841_), .B(new_n788_), .Y(\asquared[21] ));
  NOR2X1   g00649(.A(new_n810_), .B(new_n808_), .Y(new_n843_));
  AOI21X1  g00650(.A0(new_n839_), .A1(new_n811_), .B0(new_n843_), .Y(new_n844_));
  XOR2X1   g00651(.A(new_n835_), .B(new_n801_), .Y(new_n845_));
  AND2X1   g00652(.A(new_n826_), .B(new_n825_), .Y(new_n846_));
  AOI21X1  g00653(.A0(new_n827_), .A1(new_n824_), .B0(new_n846_), .Y(new_n847_));
  INVX1    g00654(.A(new_n847_), .Y(new_n848_));
  XOR2X1   g00655(.A(new_n848_), .B(new_n845_), .Y(new_n849_));
  INVX1    g00656(.A(new_n849_), .Y(new_n850_));
  INVX1    g00657(.A(new_n791_), .Y(new_n851_));
  OR2X1    g00658(.A(new_n803_), .B(new_n851_), .Y(new_n852_));
  OAI21X1  g00659(.A0(new_n806_), .A1(new_n804_), .B0(new_n852_), .Y(new_n853_));
  XOR2X1   g00660(.A(new_n853_), .B(new_n850_), .Y(new_n854_));
  AND2X1   g00661(.A(\a[19] ), .B(\a[18] ), .Y(new_n855_));
  AND2X1   g00662(.A(new_n855_), .B(new_n231_), .Y(new_n856_));
  AND2X1   g00663(.A(\a[16] ), .B(\a[2] ), .Y(new_n857_));
  AOI22X1  g00664(.A0(new_n794_), .A1(\a[3] ), .B0(new_n857_), .B1(\a[19] ), .Y(new_n858_));
  NOR3X1   g00665(.A(new_n858_), .B(new_n856_), .C(new_n255_), .Y(new_n859_));
  NOR2X1   g00666(.A(new_n859_), .B(new_n856_), .Y(new_n860_));
  INVX1    g00667(.A(new_n860_), .Y(new_n861_));
  AOI22X1  g00668(.A0(\a[19] ), .A1(\a[2] ), .B0(\a[18] ), .B1(\a[3] ), .Y(new_n862_));
  AND2X1   g00669(.A(\a[16] ), .B(\a[5] ), .Y(new_n863_));
  INVX1    g00670(.A(new_n863_), .Y(new_n864_));
  OAI22X1  g00671(.A0(new_n864_), .A1(new_n859_), .B0(new_n862_), .B1(new_n861_), .Y(new_n865_));
  INVX1    g00672(.A(new_n639_), .Y(new_n866_));
  INVX1    g00673(.A(new_n691_), .Y(new_n867_));
  OAI22X1  g00674(.A0(new_n867_), .A1(new_n376_), .B0(new_n866_), .B1(new_n280_), .Y(new_n868_));
  OAI21X1  g00675(.A0(new_n583_), .A1(new_n445_), .B0(new_n868_), .Y(new_n869_));
  AND2X1   g00676(.A(\a[15] ), .B(\a[6] ), .Y(new_n870_));
  AOI21X1  g00677(.A0(new_n582_), .A1(new_n325_), .B0(new_n868_), .Y(new_n871_));
  OAI22X1  g00678(.A0(new_n490_), .A1(new_n532_), .B0(new_n591_), .B1(new_n413_), .Y(new_n872_));
  AOI22X1  g00679(.A0(new_n872_), .A1(new_n871_), .B0(new_n870_), .B1(new_n869_), .Y(new_n873_));
  XOR2X1   g00680(.A(new_n873_), .B(new_n865_), .Y(new_n874_));
  INVX1    g00681(.A(new_n874_), .Y(new_n875_));
  AND2X1   g00682(.A(\a[17] ), .B(\a[4] ), .Y(new_n876_));
  AOI22X1  g00683(.A0(\a[12] ), .A1(\a[9] ), .B0(\a[11] ), .B1(\a[10] ), .Y(new_n877_));
  INVX1    g00684(.A(new_n877_), .Y(new_n878_));
  NAND4X1  g00685(.A(\a[12] ), .B(\a[11] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n879_));
  NAND3X1  g00686(.A(new_n878_), .B(new_n879_), .C(new_n876_), .Y(new_n880_));
  INVX1    g00687(.A(new_n735_), .Y(new_n881_));
  AOI22X1  g00688(.A0(new_n878_), .A1(new_n876_), .B0(new_n482_), .B1(new_n881_), .Y(new_n882_));
  AOI22X1  g00689(.A0(new_n882_), .A1(new_n878_), .B0(new_n880_), .B1(new_n876_), .Y(new_n883_));
  XOR2X1   g00690(.A(new_n883_), .B(new_n875_), .Y(new_n884_));
  XOR2X1   g00691(.A(new_n884_), .B(new_n854_), .Y(new_n885_));
  INVX1    g00692(.A(new_n815_), .Y(new_n886_));
  NOR2X1   g00693(.A(new_n886_), .B(new_n738_), .Y(new_n887_));
  NOR2X1   g00694(.A(new_n816_), .B(new_n757_), .Y(new_n888_));
  NOR2X1   g00695(.A(new_n888_), .B(new_n887_), .Y(new_n889_));
  AND2X1   g00696(.A(new_n814_), .B(new_n813_), .Y(new_n890_));
  AND2X1   g00697(.A(\a[21] ), .B(\a[0] ), .Y(new_n891_));
  XOR2X1   g00698(.A(new_n891_), .B(new_n890_), .Y(new_n892_));
  INVX1    g00699(.A(new_n892_), .Y(new_n893_));
  AND2X1   g00700(.A(\a[20] ), .B(\a[1] ), .Y(new_n894_));
  XOR2X1   g00701(.A(new_n894_), .B(new_n488_), .Y(new_n895_));
  XOR2X1   g00702(.A(new_n895_), .B(new_n893_), .Y(new_n896_));
  XOR2X1   g00703(.A(new_n896_), .B(new_n889_), .Y(new_n897_));
  OR2X1    g00704(.A(new_n829_), .B(new_n766_), .Y(new_n898_));
  AND2X1   g00705(.A(new_n829_), .B(new_n766_), .Y(new_n899_));
  OAI21X1  g00706(.A0(new_n837_), .A1(new_n899_), .B0(new_n898_), .Y(new_n900_));
  XOR2X1   g00707(.A(new_n900_), .B(new_n897_), .Y(new_n901_));
  OR2X1    g00708(.A(new_n822_), .B(new_n817_), .Y(new_n902_));
  OR2X1    g00709(.A(new_n838_), .B(new_n823_), .Y(new_n903_));
  AND2X1   g00710(.A(new_n903_), .B(new_n902_), .Y(new_n904_));
  XOR2X1   g00711(.A(new_n904_), .B(new_n901_), .Y(new_n905_));
  XOR2X1   g00712(.A(new_n905_), .B(new_n885_), .Y(new_n906_));
  XOR2X1   g00713(.A(new_n906_), .B(new_n844_), .Y(new_n907_));
  NOR2X1   g00714(.A(new_n840_), .B(new_n790_), .Y(new_n908_));
  AND2X1   g00715(.A(new_n840_), .B(new_n790_), .Y(new_n909_));
  INVX1    g00716(.A(new_n909_), .Y(new_n910_));
  AOI21X1  g00717(.A0(new_n910_), .A1(new_n788_), .B0(new_n908_), .Y(new_n911_));
  XOR2X1   g00718(.A(new_n911_), .B(new_n907_), .Y(\asquared[22] ));
  NAND2X1  g00719(.A(new_n905_), .B(new_n885_), .Y(new_n913_));
  OAI21X1  g00720(.A0(new_n904_), .A1(new_n901_), .B0(new_n913_), .Y(new_n914_));
  XOR2X1   g00721(.A(new_n871_), .B(new_n860_), .Y(new_n915_));
  INVX1    g00722(.A(new_n915_), .Y(new_n916_));
  NOR2X1   g00723(.A(new_n895_), .B(new_n893_), .Y(new_n917_));
  AOI21X1  g00724(.A0(new_n891_), .A1(new_n890_), .B0(new_n917_), .Y(new_n918_));
  XOR2X1   g00725(.A(new_n918_), .B(new_n916_), .Y(new_n919_));
  INVX1    g00726(.A(new_n889_), .Y(new_n920_));
  OR2X1    g00727(.A(new_n896_), .B(new_n920_), .Y(new_n921_));
  AND2X1   g00728(.A(new_n896_), .B(new_n920_), .Y(new_n922_));
  AOI21X1  g00729(.A0(new_n900_), .A1(new_n921_), .B0(new_n922_), .Y(new_n923_));
  XOR2X1   g00730(.A(new_n923_), .B(new_n919_), .Y(new_n924_));
  AOI22X1  g00731(.A0(\a[15] ), .A1(\a[7] ), .B0(\a[14] ), .B1(\a[8] ), .Y(new_n925_));
  AND2X1   g00732(.A(\a[22] ), .B(\a[0] ), .Y(new_n926_));
  INVX1    g00733(.A(new_n926_), .Y(new_n927_));
  AND2X1   g00734(.A(new_n691_), .B(new_n325_), .Y(new_n928_));
  NOR3X1   g00735(.A(new_n927_), .B(new_n928_), .C(new_n925_), .Y(new_n929_));
  INVX1    g00736(.A(new_n925_), .Y(new_n930_));
  AOI21X1  g00737(.A0(new_n926_), .A1(new_n930_), .B0(new_n928_), .Y(new_n931_));
  INVX1    g00738(.A(new_n931_), .Y(new_n932_));
  OAI22X1  g00739(.A0(new_n932_), .A1(new_n925_), .B0(new_n929_), .B1(new_n927_), .Y(new_n933_));
  INVX1    g00740(.A(\a[20] ), .Y(new_n934_));
  NOR4X1   g00741(.A(new_n934_), .B(new_n571_), .C(new_n230_), .D(new_n200_), .Y(new_n935_));
  AOI22X1  g00742(.A0(\a[20] ), .A1(\a[2] ), .B0(\a[16] ), .B1(\a[6] ), .Y(new_n936_));
  OR4X1    g00743(.A(new_n936_), .B(new_n935_), .C(new_n591_), .D(new_n341_), .Y(new_n937_));
  NOR3X1   g00744(.A(new_n936_), .B(new_n935_), .C(new_n430_), .Y(new_n938_));
  AOI21X1  g00745(.A0(new_n937_), .A1(new_n430_), .B0(new_n938_), .Y(new_n939_));
  XOR2X1   g00746(.A(new_n939_), .B(new_n933_), .Y(new_n940_));
  INVX1    g00747(.A(new_n940_), .Y(new_n941_));
  AND2X1   g00748(.A(\a[19] ), .B(\a[3] ), .Y(new_n942_));
  INVX1    g00749(.A(new_n942_), .Y(new_n943_));
  NAND4X1  g00750(.A(\a[19] ), .B(\a[18] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n944_));
  NAND4X1  g00751(.A(\a[19] ), .B(\a[17] ), .C(\a[5] ), .D(\a[3] ), .Y(new_n945_));
  AOI22X1  g00752(.A0(new_n945_), .A1(new_n944_), .B0(new_n796_), .B1(new_n218_), .Y(new_n946_));
  NOR2X1   g00753(.A(new_n946_), .B(new_n943_), .Y(new_n947_));
  AOI21X1  g00754(.A0(new_n796_), .A1(new_n218_), .B0(new_n946_), .Y(new_n948_));
  OAI22X1  g00755(.A0(new_n675_), .A1(new_n340_), .B0(new_n616_), .B1(new_n255_), .Y(new_n949_));
  AOI21X1  g00756(.A0(new_n949_), .A1(new_n948_), .B0(new_n947_), .Y(new_n950_));
  XOR2X1   g00757(.A(new_n950_), .B(new_n941_), .Y(new_n951_));
  XOR2X1   g00758(.A(new_n951_), .B(new_n924_), .Y(new_n952_));
  NAND2X1  g00759(.A(new_n853_), .B(new_n849_), .Y(new_n953_));
  OAI21X1  g00760(.A0(new_n884_), .A1(new_n854_), .B0(new_n953_), .Y(new_n954_));
  INVX1    g00761(.A(new_n865_), .Y(new_n955_));
  NOR2X1   g00762(.A(new_n873_), .B(new_n955_), .Y(new_n956_));
  NOR2X1   g00763(.A(new_n883_), .B(new_n874_), .Y(new_n957_));
  NOR2X1   g00764(.A(new_n957_), .B(new_n956_), .Y(new_n958_));
  NOR2X1   g00765(.A(new_n835_), .B(new_n801_), .Y(new_n959_));
  AOI21X1  g00766(.A0(new_n848_), .A1(new_n845_), .B0(new_n959_), .Y(new_n960_));
  INVX1    g00767(.A(new_n882_), .Y(new_n961_));
  AND2X1   g00768(.A(new_n894_), .B(\a[11] ), .Y(new_n962_));
  AND2X1   g00769(.A(\a[21] ), .B(\a[1] ), .Y(new_n963_));
  XOR2X1   g00770(.A(new_n963_), .B(new_n396_), .Y(new_n964_));
  XOR2X1   g00771(.A(new_n964_), .B(new_n962_), .Y(new_n965_));
  XOR2X1   g00772(.A(new_n965_), .B(new_n961_), .Y(new_n966_));
  XOR2X1   g00773(.A(new_n966_), .B(new_n960_), .Y(new_n967_));
  XOR2X1   g00774(.A(new_n967_), .B(new_n958_), .Y(new_n968_));
  INVX1    g00775(.A(new_n968_), .Y(new_n969_));
  OR2X1    g00776(.A(new_n969_), .B(new_n954_), .Y(new_n970_));
  XOR2X1   g00777(.A(new_n968_), .B(new_n954_), .Y(new_n971_));
  AOI21X1  g00778(.A0(new_n969_), .A1(new_n954_), .B0(new_n952_), .Y(new_n972_));
  AOI22X1  g00779(.A0(new_n972_), .A1(new_n970_), .B0(new_n971_), .B1(new_n952_), .Y(new_n973_));
  AND2X1   g00780(.A(new_n973_), .B(new_n914_), .Y(new_n974_));
  INVX1    g00781(.A(new_n974_), .Y(new_n975_));
  INVX1    g00782(.A(new_n844_), .Y(new_n976_));
  AND2X1   g00783(.A(new_n906_), .B(new_n976_), .Y(new_n977_));
  INVX1    g00784(.A(new_n977_), .Y(new_n978_));
  NOR2X1   g00785(.A(new_n906_), .B(new_n976_), .Y(new_n979_));
  OAI21X1  g00786(.A0(new_n911_), .A1(new_n979_), .B0(new_n978_), .Y(new_n980_));
  NOR2X1   g00787(.A(new_n973_), .B(new_n914_), .Y(new_n981_));
  INVX1    g00788(.A(new_n981_), .Y(new_n982_));
  AOI21X1  g00789(.A0(new_n982_), .A1(new_n975_), .B0(new_n980_), .Y(new_n983_));
  AND2X1   g00790(.A(new_n982_), .B(new_n980_), .Y(new_n984_));
  AOI21X1  g00791(.A0(new_n984_), .A1(new_n975_), .B0(new_n983_), .Y(\asquared[23] ));
  AND2X1   g00792(.A(new_n968_), .B(new_n954_), .Y(new_n986_));
  AOI21X1  g00793(.A0(new_n971_), .A1(new_n952_), .B0(new_n986_), .Y(new_n987_));
  INVX1    g00794(.A(new_n966_), .Y(new_n988_));
  NOR2X1   g00795(.A(new_n988_), .B(new_n960_), .Y(new_n989_));
  INVX1    g00796(.A(new_n989_), .Y(new_n990_));
  OAI21X1  g00797(.A0(new_n967_), .A1(new_n958_), .B0(new_n990_), .Y(new_n991_));
  AND2X1   g00798(.A(\a[20] ), .B(\a[18] ), .Y(new_n992_));
  NAND4X1  g00799(.A(\a[20] ), .B(\a[17] ), .C(\a[6] ), .D(\a[3] ), .Y(new_n993_));
  NAND4X1  g00800(.A(\a[18] ), .B(\a[17] ), .C(\a[6] ), .D(\a[5] ), .Y(new_n994_));
  AOI22X1  g00801(.A0(new_n994_), .A1(new_n993_), .B0(new_n992_), .B1(new_n272_), .Y(new_n995_));
  AOI21X1  g00802(.A0(new_n992_), .A1(new_n272_), .B0(new_n995_), .Y(new_n996_));
  OAI22X1  g00803(.A0(new_n934_), .A1(new_n223_), .B0(new_n675_), .B1(new_n255_), .Y(new_n997_));
  NOR3X1   g00804(.A(new_n995_), .B(new_n616_), .C(new_n230_), .Y(new_n998_));
  AOI21X1  g00805(.A0(new_n997_), .A1(new_n996_), .B0(new_n998_), .Y(new_n999_));
  AOI22X1  g00806(.A0(\a[13] ), .A1(\a[10] ), .B0(\a[12] ), .B1(\a[11] ), .Y(new_n1000_));
  AND2X1   g00807(.A(\a[19] ), .B(\a[4] ), .Y(new_n1001_));
  AND2X1   g00808(.A(\a[11] ), .B(\a[10] ), .Y(new_n1002_));
  AND2X1   g00809(.A(new_n586_), .B(new_n1002_), .Y(new_n1003_));
  OAI21X1  g00810(.A0(new_n1000_), .A1(new_n1003_), .B0(new_n1001_), .Y(new_n1004_));
  INVX1    g00811(.A(new_n1000_), .Y(new_n1005_));
  AOI21X1  g00812(.A0(new_n1005_), .A1(new_n1001_), .B0(new_n1003_), .Y(new_n1006_));
  INVX1    g00813(.A(new_n1006_), .Y(new_n1007_));
  OAI21X1  g00814(.A0(new_n1007_), .A1(new_n1000_), .B0(new_n1004_), .Y(new_n1008_));
  XOR2X1   g00815(.A(new_n1008_), .B(new_n999_), .Y(new_n1009_));
  AND2X1   g00816(.A(new_n964_), .B(new_n962_), .Y(new_n1010_));
  AOI21X1  g00817(.A0(new_n965_), .A1(new_n961_), .B0(new_n1010_), .Y(new_n1011_));
  XOR2X1   g00818(.A(new_n1011_), .B(new_n1009_), .Y(new_n1012_));
  AOI22X1  g00819(.A0(\a[23] ), .A1(\a[0] ), .B0(\a[21] ), .B1(\a[2] ), .Y(new_n1013_));
  INVX1    g00820(.A(new_n1013_), .Y(new_n1014_));
  AND2X1   g00821(.A(new_n963_), .B(new_n396_), .Y(new_n1015_));
  AND2X1   g00822(.A(\a[23] ), .B(\a[21] ), .Y(new_n1016_));
  AND2X1   g00823(.A(new_n1016_), .B(new_n197_), .Y(new_n1017_));
  AOI21X1  g00824(.A0(new_n1014_), .A1(new_n1015_), .B0(new_n1017_), .Y(new_n1018_));
  NAND2X1  g00825(.A(new_n1018_), .B(new_n1014_), .Y(new_n1019_));
  OAI21X1  g00826(.A0(new_n1017_), .A1(new_n1013_), .B0(new_n1015_), .Y(new_n1020_));
  AND2X1   g00827(.A(new_n1020_), .B(new_n1019_), .Y(new_n1021_));
  XOR2X1   g00828(.A(new_n1021_), .B(new_n932_), .Y(new_n1022_));
  INVX1    g00829(.A(new_n596_), .Y(new_n1023_));
  INVX1    g00830(.A(new_n689_), .Y(new_n1024_));
  INVX1    g00831(.A(new_n690_), .Y(new_n1025_));
  OAI22X1  g00832(.A0(new_n1025_), .A1(new_n1023_), .B0(new_n1024_), .B1(new_n445_), .Y(new_n1026_));
  OAI21X1  g00833(.A0(new_n867_), .A1(new_n366_), .B0(new_n1026_), .Y(new_n1027_));
  AND2X1   g00834(.A(\a[16] ), .B(\a[7] ), .Y(new_n1028_));
  OAI22X1  g00835(.A0(new_n549_), .A1(new_n413_), .B0(new_n490_), .B1(new_n341_), .Y(new_n1029_));
  INVX1    g00836(.A(new_n366_), .Y(new_n1030_));
  AOI21X1  g00837(.A0(new_n691_), .A1(new_n1030_), .B0(new_n1026_), .Y(new_n1031_));
  AOI22X1  g00838(.A0(new_n1031_), .A1(new_n1029_), .B0(new_n1028_), .B1(new_n1027_), .Y(new_n1032_));
  XOR2X1   g00839(.A(new_n1032_), .B(new_n1022_), .Y(new_n1033_));
  XOR2X1   g00840(.A(new_n1033_), .B(new_n1012_), .Y(new_n1034_));
  XOR2X1   g00841(.A(new_n1034_), .B(new_n991_), .Y(new_n1035_));
  INVX1    g00842(.A(new_n1035_), .Y(new_n1036_));
  INVX1    g00843(.A(new_n919_), .Y(new_n1037_));
  OR2X1    g00844(.A(new_n923_), .B(new_n1037_), .Y(new_n1038_));
  OAI21X1  g00845(.A0(new_n951_), .A1(new_n924_), .B0(new_n1038_), .Y(new_n1039_));
  OR2X1    g00846(.A(new_n871_), .B(new_n860_), .Y(new_n1040_));
  OAI21X1  g00847(.A0(new_n918_), .A1(new_n916_), .B0(new_n1040_), .Y(new_n1041_));
  INVX1    g00848(.A(new_n933_), .Y(new_n1042_));
  OR2X1    g00849(.A(new_n950_), .B(new_n940_), .Y(new_n1043_));
  OAI21X1  g00850(.A0(new_n939_), .A1(new_n1042_), .B0(new_n1043_), .Y(new_n1044_));
  XOR2X1   g00851(.A(new_n1044_), .B(new_n1041_), .Y(new_n1045_));
  NOR3X1   g00852(.A(new_n936_), .B(new_n591_), .C(new_n341_), .Y(new_n1046_));
  NOR2X1   g00853(.A(new_n1046_), .B(new_n935_), .Y(new_n1047_));
  INVX1    g00854(.A(new_n1047_), .Y(new_n1048_));
  INVX1    g00855(.A(new_n948_), .Y(new_n1049_));
  AND2X1   g00856(.A(\a[22] ), .B(\a[1] ), .Y(new_n1050_));
  XOR2X1   g00857(.A(new_n1050_), .B(\a[12] ), .Y(new_n1051_));
  XOR2X1   g00858(.A(new_n1051_), .B(new_n1049_), .Y(new_n1052_));
  XOR2X1   g00859(.A(new_n1052_), .B(new_n1048_), .Y(new_n1053_));
  XOR2X1   g00860(.A(new_n1053_), .B(new_n1045_), .Y(new_n1054_));
  XOR2X1   g00861(.A(new_n1054_), .B(new_n1039_), .Y(new_n1055_));
  XOR2X1   g00862(.A(new_n1055_), .B(new_n1036_), .Y(new_n1056_));
  AND2X1   g00863(.A(new_n1056_), .B(new_n987_), .Y(new_n1057_));
  NOR2X1   g00864(.A(new_n1056_), .B(new_n987_), .Y(new_n1058_));
  OR2X1    g00865(.A(new_n1058_), .B(new_n1057_), .Y(new_n1059_));
  AOI21X1  g00866(.A0(new_n982_), .A1(new_n980_), .B0(new_n974_), .Y(new_n1060_));
  XOR2X1   g00867(.A(new_n1060_), .B(new_n1059_), .Y(\asquared[24] ));
  AND2X1   g00868(.A(new_n1054_), .B(new_n1039_), .Y(new_n1062_));
  AOI21X1  g00869(.A0(new_n1055_), .A1(new_n1035_), .B0(new_n1062_), .Y(new_n1063_));
  INVX1    g00870(.A(new_n1063_), .Y(new_n1064_));
  AND2X1   g00871(.A(new_n1033_), .B(new_n1012_), .Y(new_n1065_));
  AND2X1   g00872(.A(new_n1034_), .B(new_n991_), .Y(new_n1066_));
  OR2X1    g00873(.A(new_n1066_), .B(new_n1065_), .Y(new_n1067_));
  XOR2X1   g00874(.A(new_n1006_), .B(new_n996_), .Y(new_n1068_));
  XOR2X1   g00875(.A(new_n1068_), .B(new_n1031_), .Y(new_n1069_));
  AND2X1   g00876(.A(new_n997_), .B(new_n996_), .Y(new_n1070_));
  OAI21X1  g00877(.A0(new_n998_), .A1(new_n1070_), .B0(new_n1008_), .Y(new_n1071_));
  OAI21X1  g00878(.A0(new_n1011_), .A1(new_n1009_), .B0(new_n1071_), .Y(new_n1072_));
  OR2X1    g00879(.A(new_n1021_), .B(new_n931_), .Y(new_n1073_));
  OAI21X1  g00880(.A0(new_n1032_), .A1(new_n1022_), .B0(new_n1073_), .Y(new_n1074_));
  INVX1    g00881(.A(new_n1074_), .Y(new_n1075_));
  XOR2X1   g00882(.A(new_n1075_), .B(new_n1072_), .Y(new_n1076_));
  XOR2X1   g00883(.A(new_n1076_), .B(new_n1069_), .Y(new_n1077_));
  XOR2X1   g00884(.A(new_n1077_), .B(new_n1067_), .Y(new_n1078_));
  NAND3X1  g00885(.A(\a[22] ), .B(\a[12] ), .C(\a[1] ), .Y(new_n1079_));
  AND2X1   g00886(.A(\a[24] ), .B(\a[0] ), .Y(new_n1080_));
  XOR2X1   g00887(.A(new_n1080_), .B(new_n1079_), .Y(new_n1081_));
  AND2X1   g00888(.A(\a[23] ), .B(\a[1] ), .Y(new_n1082_));
  XOR2X1   g00889(.A(new_n1082_), .B(new_n635_), .Y(new_n1083_));
  XOR2X1   g00890(.A(new_n1083_), .B(new_n1081_), .Y(new_n1084_));
  NAND2X1  g00891(.A(\a[17] ), .B(\a[7] ), .Y(new_n1085_));
  INVX1    g00892(.A(\a[22] ), .Y(new_n1086_));
  NOR4X1   g00893(.A(new_n1086_), .B(new_n675_), .C(new_n230_), .D(new_n200_), .Y(new_n1087_));
  NAND4X1  g00894(.A(\a[18] ), .B(\a[17] ), .C(\a[7] ), .D(\a[6] ), .Y(new_n1088_));
  NAND4X1  g00895(.A(\a[22] ), .B(\a[17] ), .C(\a[7] ), .D(\a[2] ), .Y(new_n1089_));
  AOI21X1  g00896(.A0(new_n1089_), .A1(new_n1088_), .B0(new_n1087_), .Y(new_n1090_));
  OR2X1    g00897(.A(new_n1090_), .B(new_n1087_), .Y(new_n1091_));
  AOI22X1  g00898(.A0(\a[22] ), .A1(\a[2] ), .B0(\a[18] ), .B1(\a[6] ), .Y(new_n1092_));
  OAI22X1  g00899(.A0(new_n1092_), .A1(new_n1091_), .B0(new_n1090_), .B1(new_n1085_), .Y(new_n1093_));
  XOR2X1   g00900(.A(new_n1093_), .B(new_n1084_), .Y(new_n1094_));
  AND2X1   g00901(.A(new_n1051_), .B(new_n1049_), .Y(new_n1095_));
  AOI21X1  g00902(.A0(new_n1052_), .A1(new_n1048_), .B0(new_n1095_), .Y(new_n1096_));
  XOR2X1   g00903(.A(new_n1096_), .B(new_n1094_), .Y(new_n1097_));
  INVX1    g00904(.A(\a[21] ), .Y(new_n1098_));
  AND2X1   g00905(.A(\a[20] ), .B(\a[19] ), .Y(new_n1099_));
  NAND4X1  g00906(.A(\a[21] ), .B(\a[19] ), .C(\a[5] ), .D(\a[3] ), .Y(new_n1100_));
  NAND4X1  g00907(.A(\a[21] ), .B(\a[20] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n1101_));
  AOI22X1  g00908(.A0(new_n1101_), .A1(new_n1100_), .B0(new_n1099_), .B1(new_n218_), .Y(new_n1102_));
  NOR3X1   g00909(.A(new_n1102_), .B(new_n1098_), .C(new_n223_), .Y(new_n1103_));
  AOI21X1  g00910(.A0(new_n1099_), .A1(new_n218_), .B0(new_n1102_), .Y(new_n1104_));
  AOI22X1  g00911(.A0(\a[20] ), .A1(\a[4] ), .B0(\a[19] ), .B1(\a[5] ), .Y(new_n1105_));
  INVX1    g00912(.A(new_n1105_), .Y(new_n1106_));
  AOI21X1  g00913(.A0(new_n1106_), .A1(new_n1104_), .B0(new_n1103_), .Y(new_n1107_));
  XOR2X1   g00914(.A(new_n1107_), .B(new_n1018_), .Y(new_n1108_));
  INVX1    g00915(.A(new_n1108_), .Y(new_n1109_));
  AND2X1   g00916(.A(\a[16] ), .B(\a[8] ), .Y(new_n1110_));
  OAI22X1  g00917(.A0(new_n1025_), .A1(new_n699_), .B0(new_n1024_), .B1(new_n366_), .Y(new_n1111_));
  OAI21X1  g00918(.A0(new_n867_), .A1(new_n735_), .B0(new_n1111_), .Y(new_n1112_));
  AOI21X1  g00919(.A0(new_n691_), .A1(new_n881_), .B0(new_n1111_), .Y(new_n1113_));
  OAI22X1  g00920(.A0(new_n549_), .A1(new_n341_), .B0(new_n490_), .B1(new_n570_), .Y(new_n1114_));
  AOI22X1  g00921(.A0(new_n1114_), .A1(new_n1113_), .B0(new_n1112_), .B1(new_n1110_), .Y(new_n1115_));
  XOR2X1   g00922(.A(new_n1115_), .B(new_n1109_), .Y(new_n1116_));
  XOR2X1   g00923(.A(new_n1116_), .B(new_n1097_), .Y(new_n1117_));
  AND2X1   g00924(.A(new_n1044_), .B(new_n1041_), .Y(new_n1118_));
  AOI21X1  g00925(.A0(new_n1053_), .A1(new_n1045_), .B0(new_n1118_), .Y(new_n1119_));
  XOR2X1   g00926(.A(new_n1119_), .B(new_n1117_), .Y(new_n1120_));
  XOR2X1   g00927(.A(new_n1120_), .B(new_n1078_), .Y(new_n1121_));
  AND2X1   g00928(.A(new_n1121_), .B(new_n1064_), .Y(new_n1122_));
  INVX1    g00929(.A(new_n1122_), .Y(new_n1123_));
  INVX1    g00930(.A(new_n1058_), .Y(new_n1124_));
  OAI21X1  g00931(.A0(new_n1060_), .A1(new_n1057_), .B0(new_n1124_), .Y(new_n1125_));
  NOR2X1   g00932(.A(new_n1121_), .B(new_n1064_), .Y(new_n1126_));
  INVX1    g00933(.A(new_n1126_), .Y(new_n1127_));
  AOI21X1  g00934(.A0(new_n1127_), .A1(new_n1123_), .B0(new_n1125_), .Y(new_n1128_));
  AND2X1   g00935(.A(new_n1127_), .B(new_n1125_), .Y(new_n1129_));
  AOI21X1  g00936(.A0(new_n1129_), .A1(new_n1123_), .B0(new_n1128_), .Y(\asquared[25] ));
  AND2X1   g00937(.A(new_n1077_), .B(new_n1067_), .Y(new_n1131_));
  AND2X1   g00938(.A(new_n1120_), .B(new_n1078_), .Y(new_n1132_));
  AOI22X1  g00939(.A0(\a[25] ), .A1(\a[0] ), .B0(\a[23] ), .B1(\a[2] ), .Y(new_n1133_));
  AND2X1   g00940(.A(\a[25] ), .B(\a[23] ), .Y(new_n1134_));
  AND2X1   g00941(.A(new_n1134_), .B(new_n197_), .Y(new_n1135_));
  NOR3X1   g00942(.A(new_n1135_), .B(new_n1133_), .C(new_n544_), .Y(new_n1136_));
  INVX1    g00943(.A(new_n544_), .Y(new_n1137_));
  INVX1    g00944(.A(new_n1133_), .Y(new_n1138_));
  AOI21X1  g00945(.A0(new_n1138_), .A1(new_n1137_), .B0(new_n1135_), .Y(new_n1139_));
  INVX1    g00946(.A(new_n1139_), .Y(new_n1140_));
  OAI22X1  g00947(.A0(new_n1140_), .A1(new_n1133_), .B0(new_n1136_), .B1(new_n544_), .Y(new_n1141_));
  OAI22X1  g00948(.A0(new_n797_), .A1(new_n445_), .B0(new_n795_), .B1(new_n1023_), .Y(new_n1142_));
  OAI21X1  g00949(.A0(new_n793_), .A1(new_n366_), .B0(new_n1142_), .Y(new_n1143_));
  AOI21X1  g00950(.A0(new_n792_), .A1(new_n1030_), .B0(new_n1142_), .Y(new_n1144_));
  OAI22X1  g00951(.A0(new_n616_), .A1(new_n413_), .B0(new_n571_), .B1(new_n341_), .Y(new_n1145_));
  AOI22X1  g00952(.A0(new_n1145_), .A1(new_n1144_), .B0(new_n1143_), .B1(new_n677_), .Y(new_n1146_));
  XOR2X1   g00953(.A(new_n1146_), .B(new_n1141_), .Y(new_n1147_));
  AND2X1   g00954(.A(\a[21] ), .B(\a[19] ), .Y(new_n1148_));
  INVX1    g00955(.A(new_n1148_), .Y(new_n1149_));
  OAI22X1  g00956(.A0(new_n1149_), .A1(new_n340_), .B0(new_n943_), .B1(new_n1086_), .Y(new_n1150_));
  NAND4X1  g00957(.A(\a[22] ), .B(\a[21] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n1151_));
  NAND3X1  g00958(.A(new_n1151_), .B(new_n1150_), .C(\a[6] ), .Y(new_n1152_));
  AND2X1   g00959(.A(\a[19] ), .B(\a[6] ), .Y(new_n1153_));
  AND2X1   g00960(.A(\a[22] ), .B(\a[21] ), .Y(new_n1154_));
  AOI22X1  g00961(.A0(new_n1154_), .A1(new_n294_), .B0(new_n1150_), .B1(\a[6] ), .Y(new_n1155_));
  OAI22X1  g00962(.A0(new_n1086_), .A1(new_n223_), .B0(new_n1098_), .B1(new_n340_), .Y(new_n1156_));
  AOI22X1  g00963(.A0(new_n1156_), .A1(new_n1155_), .B0(new_n1153_), .B1(new_n1152_), .Y(new_n1157_));
  XOR2X1   g00964(.A(new_n1157_), .B(new_n1147_), .Y(new_n1158_));
  NAND2X1  g00965(.A(new_n1074_), .B(new_n1072_), .Y(new_n1159_));
  OAI21X1  g00966(.A0(new_n1076_), .A1(new_n1069_), .B0(new_n1159_), .Y(new_n1160_));
  XOR2X1   g00967(.A(new_n1160_), .B(new_n1158_), .Y(new_n1161_));
  AND2X1   g00968(.A(new_n1082_), .B(new_n634_), .Y(new_n1162_));
  AND2X1   g00969(.A(\a[24] ), .B(\a[1] ), .Y(new_n1163_));
  XOR2X1   g00970(.A(new_n1163_), .B(\a[13] ), .Y(new_n1164_));
  XOR2X1   g00971(.A(new_n1164_), .B(new_n1162_), .Y(new_n1165_));
  INVX1    g00972(.A(new_n1165_), .Y(new_n1166_));
  XOR2X1   g00973(.A(new_n1166_), .B(new_n1104_), .Y(new_n1167_));
  INVX1    g00974(.A(new_n1031_), .Y(new_n1168_));
  NOR2X1   g00975(.A(new_n1006_), .B(new_n996_), .Y(new_n1169_));
  AOI21X1  g00976(.A0(new_n1068_), .A1(new_n1168_), .B0(new_n1169_), .Y(new_n1170_));
  AND2X1   g00977(.A(\a[20] ), .B(\a[5] ), .Y(new_n1171_));
  INVX1    g00978(.A(new_n1171_), .Y(new_n1172_));
  AOI22X1  g00979(.A0(\a[14] ), .A1(\a[11] ), .B0(\a[13] ), .B1(\a[12] ), .Y(new_n1173_));
  NOR4X1   g00980(.A(new_n490_), .B(new_n591_), .C(new_n453_), .D(new_n488_), .Y(new_n1174_));
  NOR3X1   g00981(.A(new_n1173_), .B(new_n1174_), .C(new_n1172_), .Y(new_n1175_));
  INVX1    g00982(.A(new_n1173_), .Y(new_n1176_));
  AOI21X1  g00983(.A0(new_n1176_), .A1(new_n1171_), .B0(new_n1174_), .Y(new_n1177_));
  INVX1    g00984(.A(new_n1177_), .Y(new_n1178_));
  OAI22X1  g00985(.A0(new_n1178_), .A1(new_n1173_), .B0(new_n1175_), .B1(new_n1172_), .Y(new_n1179_));
  XOR2X1   g00986(.A(new_n1179_), .B(new_n1170_), .Y(new_n1180_));
  XOR2X1   g00987(.A(new_n1180_), .B(new_n1167_), .Y(new_n1181_));
  XOR2X1   g00988(.A(new_n1181_), .B(new_n1161_), .Y(new_n1182_));
  INVX1    g00989(.A(new_n1113_), .Y(new_n1183_));
  XOR2X1   g00990(.A(new_n1183_), .B(new_n1091_), .Y(new_n1184_));
  INVX1    g00991(.A(\a[24] ), .Y(new_n1185_));
  NOR3X1   g00992(.A(new_n1079_), .B(new_n1185_), .C(new_n194_), .Y(new_n1186_));
  NOR2X1   g00993(.A(new_n1083_), .B(new_n1081_), .Y(new_n1187_));
  NOR2X1   g00994(.A(new_n1187_), .B(new_n1186_), .Y(new_n1188_));
  INVX1    g00995(.A(new_n1188_), .Y(new_n1189_));
  XOR2X1   g00996(.A(new_n1189_), .B(new_n1184_), .Y(new_n1190_));
  INVX1    g00997(.A(new_n1190_), .Y(new_n1191_));
  OR2X1    g00998(.A(new_n1107_), .B(new_n1018_), .Y(new_n1192_));
  OAI21X1  g00999(.A0(new_n1115_), .A1(new_n1109_), .B0(new_n1192_), .Y(new_n1193_));
  XOR2X1   g01000(.A(new_n1193_), .B(new_n1191_), .Y(new_n1194_));
  AND2X1   g01001(.A(new_n1093_), .B(new_n1084_), .Y(new_n1195_));
  INVX1    g01002(.A(new_n1195_), .Y(new_n1196_));
  INVX1    g01003(.A(new_n1094_), .Y(new_n1197_));
  OAI21X1  g01004(.A0(new_n1096_), .A1(new_n1197_), .B0(new_n1196_), .Y(new_n1198_));
  INVX1    g01005(.A(new_n1198_), .Y(new_n1199_));
  XOR2X1   g01006(.A(new_n1199_), .B(new_n1194_), .Y(new_n1200_));
  INVX1    g01007(.A(new_n1200_), .Y(new_n1201_));
  INVX1    g01008(.A(new_n1116_), .Y(new_n1202_));
  OR2X1    g01009(.A(new_n1202_), .B(new_n1097_), .Y(new_n1203_));
  OAI21X1  g01010(.A0(new_n1119_), .A1(new_n1117_), .B0(new_n1203_), .Y(new_n1204_));
  XOR2X1   g01011(.A(new_n1204_), .B(new_n1201_), .Y(new_n1205_));
  XOR2X1   g01012(.A(new_n1205_), .B(new_n1182_), .Y(new_n1206_));
  NOR3X1   g01013(.A(new_n1206_), .B(new_n1132_), .C(new_n1131_), .Y(new_n1207_));
  OR2X1    g01014(.A(new_n1132_), .B(new_n1131_), .Y(new_n1208_));
  AND2X1   g01015(.A(new_n1206_), .B(new_n1208_), .Y(new_n1209_));
  OR2X1    g01016(.A(new_n1209_), .B(new_n1207_), .Y(new_n1210_));
  AOI21X1  g01017(.A0(new_n1127_), .A1(new_n1125_), .B0(new_n1122_), .Y(new_n1211_));
  XOR2X1   g01018(.A(new_n1211_), .B(new_n1210_), .Y(\asquared[26] ));
  NAND2X1  g01019(.A(new_n1204_), .B(new_n1200_), .Y(new_n1213_));
  OAI21X1  g01020(.A0(new_n1205_), .A1(new_n1182_), .B0(new_n1213_), .Y(new_n1214_));
  AOI22X1  g01021(.A0(\a[23] ), .A1(\a[3] ), .B0(\a[19] ), .B1(\a[7] ), .Y(new_n1215_));
  INVX1    g01022(.A(\a[23] ), .Y(new_n1216_));
  NOR4X1   g01023(.A(new_n1216_), .B(new_n752_), .C(new_n532_), .D(new_n223_), .Y(new_n1217_));
  NOR3X1   g01024(.A(new_n302_), .B(new_n1185_), .C(new_n752_), .Y(new_n1218_));
  AND2X1   g01025(.A(\a[24] ), .B(\a[23] ), .Y(new_n1219_));
  AOI21X1  g01026(.A0(new_n1219_), .A1(new_n231_), .B0(new_n1218_), .Y(new_n1220_));
  NOR2X1   g01027(.A(new_n1220_), .B(new_n1217_), .Y(new_n1221_));
  NOR2X1   g01028(.A(new_n1221_), .B(new_n1217_), .Y(new_n1222_));
  INVX1    g01029(.A(new_n1222_), .Y(new_n1223_));
  NAND2X1  g01030(.A(\a[24] ), .B(\a[2] ), .Y(new_n1224_));
  OAI22X1  g01031(.A0(new_n1224_), .A1(new_n1221_), .B0(new_n1223_), .B1(new_n1215_), .Y(new_n1225_));
  AND2X1   g01032(.A(\a[17] ), .B(\a[9] ), .Y(new_n1226_));
  INVX1    g01033(.A(new_n1226_), .Y(new_n1227_));
  NAND4X1  g01034(.A(\a[17] ), .B(\a[15] ), .C(\a[11] ), .D(\a[9] ), .Y(new_n1228_));
  NAND4X1  g01035(.A(\a[17] ), .B(\a[16] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n1229_));
  AOI22X1  g01036(.A0(new_n1229_), .A1(new_n1228_), .B0(new_n689_), .B1(new_n1002_), .Y(new_n1230_));
  NAND4X1  g01037(.A(\a[16] ), .B(\a[15] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n1231_));
  NAND3X1  g01038(.A(new_n1229_), .B(new_n1228_), .C(new_n1231_), .Y(new_n1232_));
  AOI22X1  g01039(.A0(\a[16] ), .A1(\a[10] ), .B0(\a[15] ), .B1(\a[11] ), .Y(new_n1233_));
  OAI22X1  g01040(.A0(new_n1233_), .A1(new_n1232_), .B0(new_n1230_), .B1(new_n1227_), .Y(new_n1234_));
  XOR2X1   g01041(.A(new_n1234_), .B(new_n1225_), .Y(new_n1235_));
  AND2X1   g01042(.A(\a[21] ), .B(\a[20] ), .Y(new_n1236_));
  NAND4X1  g01043(.A(\a[22] ), .B(\a[20] ), .C(\a[6] ), .D(\a[4] ), .Y(new_n1237_));
  NAND4X1  g01044(.A(\a[22] ), .B(\a[21] ), .C(\a[5] ), .D(\a[4] ), .Y(new_n1238_));
  AOI22X1  g01045(.A0(new_n1238_), .A1(new_n1237_), .B0(new_n1236_), .B1(new_n295_), .Y(new_n1239_));
  AND2X1   g01046(.A(\a[22] ), .B(\a[4] ), .Y(new_n1240_));
  INVX1    g01047(.A(new_n1240_), .Y(new_n1241_));
  AOI21X1  g01048(.A0(new_n1236_), .A1(new_n295_), .B0(new_n1239_), .Y(new_n1242_));
  INVX1    g01049(.A(new_n1242_), .Y(new_n1243_));
  AOI22X1  g01050(.A0(\a[21] ), .A1(\a[5] ), .B0(\a[20] ), .B1(\a[6] ), .Y(new_n1244_));
  OAI22X1  g01051(.A0(new_n1244_), .A1(new_n1243_), .B0(new_n1241_), .B1(new_n1239_), .Y(new_n1245_));
  XOR2X1   g01052(.A(new_n1245_), .B(new_n1235_), .Y(new_n1246_));
  AND2X1   g01053(.A(new_n1193_), .B(new_n1190_), .Y(new_n1247_));
  INVX1    g01054(.A(new_n1247_), .Y(new_n1248_));
  OAI21X1  g01055(.A0(new_n1199_), .A1(new_n1194_), .B0(new_n1248_), .Y(new_n1249_));
  INVX1    g01056(.A(new_n1249_), .Y(new_n1250_));
  XOR2X1   g01057(.A(new_n1250_), .B(new_n1246_), .Y(new_n1251_));
  AND2X1   g01058(.A(new_n1183_), .B(new_n1091_), .Y(new_n1252_));
  AOI21X1  g01059(.A0(new_n1189_), .A1(new_n1184_), .B0(new_n1252_), .Y(new_n1253_));
  NAND2X1  g01060(.A(new_n1164_), .B(new_n1162_), .Y(new_n1254_));
  OR2X1    g01061(.A(new_n1166_), .B(new_n1104_), .Y(new_n1255_));
  AND2X1   g01062(.A(new_n1255_), .B(new_n1254_), .Y(new_n1256_));
  INVX1    g01063(.A(new_n1256_), .Y(new_n1257_));
  XOR2X1   g01064(.A(new_n1257_), .B(new_n1253_), .Y(new_n1258_));
  XOR2X1   g01065(.A(new_n1144_), .B(new_n1140_), .Y(new_n1259_));
  AND2X1   g01066(.A(new_n1163_), .B(\a[13] ), .Y(new_n1260_));
  INVX1    g01067(.A(new_n1260_), .Y(new_n1261_));
  AOI22X1  g01068(.A0(\a[26] ), .A1(\a[0] ), .B0(\a[18] ), .B1(\a[8] ), .Y(new_n1262_));
  INVX1    g01069(.A(\a[26] ), .Y(new_n1263_));
  NOR4X1   g01070(.A(new_n1263_), .B(new_n675_), .C(new_n413_), .D(new_n194_), .Y(new_n1264_));
  NOR3X1   g01071(.A(new_n1262_), .B(new_n1264_), .C(new_n1261_), .Y(new_n1265_));
  NOR2X1   g01072(.A(new_n1265_), .B(new_n1264_), .Y(new_n1266_));
  INVX1    g01073(.A(new_n1266_), .Y(new_n1267_));
  OAI22X1  g01074(.A0(new_n1267_), .A1(new_n1262_), .B0(new_n1265_), .B1(new_n1261_), .Y(new_n1268_));
  XOR2X1   g01075(.A(new_n1268_), .B(new_n1259_), .Y(new_n1269_));
  XOR2X1   g01076(.A(new_n1269_), .B(new_n1258_), .Y(new_n1270_));
  XOR2X1   g01077(.A(new_n1270_), .B(new_n1251_), .Y(new_n1271_));
  NAND2X1  g01078(.A(new_n1160_), .B(new_n1158_), .Y(new_n1272_));
  INVX1    g01079(.A(new_n1161_), .Y(new_n1273_));
  OAI21X1  g01080(.A0(new_n1181_), .A1(new_n1273_), .B0(new_n1272_), .Y(new_n1274_));
  INVX1    g01081(.A(new_n1167_), .Y(new_n1275_));
  INVX1    g01082(.A(new_n1179_), .Y(new_n1276_));
  OR2X1    g01083(.A(new_n1276_), .B(new_n1170_), .Y(new_n1277_));
  OAI21X1  g01084(.A0(new_n1180_), .A1(new_n1275_), .B0(new_n1277_), .Y(new_n1278_));
  INVX1    g01085(.A(new_n1141_), .Y(new_n1279_));
  OR2X1    g01086(.A(new_n1146_), .B(new_n1279_), .Y(new_n1280_));
  OAI21X1  g01087(.A0(new_n1157_), .A1(new_n1147_), .B0(new_n1280_), .Y(new_n1281_));
  INVX1    g01088(.A(new_n585_), .Y(new_n1282_));
  AND2X1   g01089(.A(\a[25] ), .B(\a[1] ), .Y(new_n1283_));
  XOR2X1   g01090(.A(new_n1283_), .B(new_n1282_), .Y(new_n1284_));
  XOR2X1   g01091(.A(new_n1284_), .B(new_n1177_), .Y(new_n1285_));
  OR2X1    g01092(.A(new_n1285_), .B(new_n1155_), .Y(new_n1286_));
  OR2X1    g01093(.A(new_n1284_), .B(new_n1177_), .Y(new_n1287_));
  NAND2X1  g01094(.A(new_n1284_), .B(new_n1177_), .Y(new_n1288_));
  NAND3X1  g01095(.A(new_n1288_), .B(new_n1287_), .C(new_n1155_), .Y(new_n1289_));
  AND2X1   g01096(.A(new_n1289_), .B(new_n1286_), .Y(new_n1290_));
  XOR2X1   g01097(.A(new_n1290_), .B(new_n1281_), .Y(new_n1291_));
  XOR2X1   g01098(.A(new_n1291_), .B(new_n1278_), .Y(new_n1292_));
  XOR2X1   g01099(.A(new_n1292_), .B(new_n1274_), .Y(new_n1293_));
  XOR2X1   g01100(.A(new_n1293_), .B(new_n1271_), .Y(new_n1294_));
  INVX1    g01101(.A(new_n1294_), .Y(new_n1295_));
  XOR2X1   g01102(.A(new_n1295_), .B(new_n1214_), .Y(new_n1296_));
  INVX1    g01103(.A(new_n1209_), .Y(new_n1297_));
  OAI21X1  g01104(.A0(new_n1211_), .A1(new_n1207_), .B0(new_n1297_), .Y(new_n1298_));
  XOR2X1   g01105(.A(new_n1298_), .B(new_n1296_), .Y(\asquared[27] ));
  INVX1    g01106(.A(new_n1271_), .Y(new_n1300_));
  AND2X1   g01107(.A(new_n1292_), .B(new_n1274_), .Y(new_n1301_));
  AOI21X1  g01108(.A0(new_n1293_), .A1(new_n1300_), .B0(new_n1301_), .Y(new_n1302_));
  AND2X1   g01109(.A(new_n1249_), .B(new_n1246_), .Y(new_n1303_));
  XOR2X1   g01110(.A(new_n1249_), .B(new_n1246_), .Y(new_n1304_));
  AOI21X1  g01111(.A0(new_n1270_), .A1(new_n1304_), .B0(new_n1303_), .Y(new_n1305_));
  INVX1    g01112(.A(new_n1305_), .Y(new_n1306_));
  NOR4X1   g01113(.A(new_n1216_), .B(new_n1098_), .C(new_n230_), .D(new_n340_), .Y(new_n1307_));
  NOR4X1   g01114(.A(new_n1185_), .B(new_n1098_), .C(new_n230_), .D(new_n223_), .Y(new_n1308_));
  AOI21X1  g01115(.A0(new_n1219_), .A1(new_n294_), .B0(new_n1308_), .Y(new_n1309_));
  OR2X1    g01116(.A(new_n1309_), .B(new_n1307_), .Y(new_n1310_));
  NOR3X1   g01117(.A(new_n217_), .B(new_n1185_), .C(new_n1216_), .Y(new_n1311_));
  NOR3X1   g01118(.A(new_n1311_), .B(new_n1308_), .C(new_n1307_), .Y(new_n1312_));
  OAI22X1  g01119(.A0(new_n1216_), .A1(new_n340_), .B0(new_n1098_), .B1(new_n230_), .Y(new_n1313_));
  AND2X1   g01120(.A(\a[24] ), .B(\a[3] ), .Y(new_n1314_));
  AOI22X1  g01121(.A0(new_n1314_), .A1(new_n1310_), .B0(new_n1313_), .B1(new_n1312_), .Y(new_n1315_));
  AND2X1   g01122(.A(\a[22] ), .B(\a[5] ), .Y(new_n1316_));
  INVX1    g01123(.A(new_n1316_), .Y(new_n1317_));
  AOI22X1  g01124(.A0(\a[15] ), .A1(\a[12] ), .B0(\a[14] ), .B1(\a[13] ), .Y(new_n1318_));
  AND2X1   g01125(.A(new_n691_), .B(new_n586_), .Y(new_n1319_));
  NOR3X1   g01126(.A(new_n1318_), .B(new_n1319_), .C(new_n1317_), .Y(new_n1320_));
  INVX1    g01127(.A(new_n1318_), .Y(new_n1321_));
  AOI21X1  g01128(.A0(new_n1321_), .A1(new_n1316_), .B0(new_n1319_), .Y(new_n1322_));
  INVX1    g01129(.A(new_n1322_), .Y(new_n1323_));
  OAI22X1  g01130(.A0(new_n1323_), .A1(new_n1318_), .B0(new_n1320_), .B1(new_n1317_), .Y(new_n1324_));
  XOR2X1   g01131(.A(new_n1324_), .B(new_n1315_), .Y(new_n1325_));
  INVX1    g01132(.A(\a[25] ), .Y(new_n1326_));
  NOR3X1   g01133(.A(new_n585_), .B(new_n1326_), .C(new_n202_), .Y(new_n1327_));
  AND2X1   g01134(.A(\a[27] ), .B(\a[0] ), .Y(new_n1328_));
  XOR2X1   g01135(.A(new_n1328_), .B(new_n1327_), .Y(new_n1329_));
  INVX1    g01136(.A(new_n1329_), .Y(new_n1330_));
  AND2X1   g01137(.A(new_n519_), .B(\a[26] ), .Y(new_n1331_));
  INVX1    g01138(.A(new_n1331_), .Y(new_n1332_));
  AND2X1   g01139(.A(\a[26] ), .B(\a[1] ), .Y(new_n1333_));
  OAI21X1  g01140(.A0(new_n1333_), .A1(\a[14] ), .B0(new_n1332_), .Y(new_n1334_));
  XOR2X1   g01141(.A(new_n1334_), .B(new_n1330_), .Y(new_n1335_));
  XOR2X1   g01142(.A(new_n1335_), .B(new_n1325_), .Y(new_n1336_));
  XOR2X1   g01143(.A(new_n1243_), .B(new_n1232_), .Y(new_n1337_));
  XOR2X1   g01144(.A(new_n1337_), .B(new_n1223_), .Y(new_n1338_));
  INVX1    g01145(.A(new_n1338_), .Y(new_n1339_));
  OR2X1    g01146(.A(new_n1256_), .B(new_n1253_), .Y(new_n1340_));
  OAI21X1  g01147(.A0(new_n1269_), .A1(new_n1258_), .B0(new_n1340_), .Y(new_n1341_));
  XOR2X1   g01148(.A(new_n1341_), .B(new_n1339_), .Y(new_n1342_));
  XOR2X1   g01149(.A(new_n1342_), .B(new_n1336_), .Y(new_n1343_));
  XOR2X1   g01150(.A(new_n1343_), .B(new_n1306_), .Y(new_n1344_));
  AND2X1   g01151(.A(\a[16] ), .B(\a[11] ), .Y(new_n1345_));
  NOR3X1   g01152(.A(new_n302_), .B(new_n1326_), .C(new_n934_), .Y(new_n1346_));
  AOI22X1  g01153(.A0(\a[25] ), .A1(\a[2] ), .B0(\a[20] ), .B1(\a[7] ), .Y(new_n1347_));
  NOR2X1   g01154(.A(new_n1347_), .B(new_n1346_), .Y(new_n1348_));
  XOR2X1   g01155(.A(new_n1348_), .B(new_n1345_), .Y(new_n1349_));
  XOR2X1   g01156(.A(new_n1349_), .B(new_n1267_), .Y(new_n1350_));
  NAND4X1  g01157(.A(\a[19] ), .B(\a[17] ), .C(\a[10] ), .D(\a[8] ), .Y(new_n1351_));
  NAND4X1  g01158(.A(\a[19] ), .B(\a[18] ), .C(\a[9] ), .D(\a[8] ), .Y(new_n1352_));
  AOI22X1  g01159(.A0(new_n1352_), .A1(new_n1351_), .B0(new_n796_), .B1(new_n881_), .Y(new_n1353_));
  NOR3X1   g01160(.A(new_n1353_), .B(new_n752_), .C(new_n413_), .Y(new_n1354_));
  AOI21X1  g01161(.A0(new_n796_), .A1(new_n881_), .B0(new_n1353_), .Y(new_n1355_));
  OAI22X1  g01162(.A0(new_n675_), .A1(new_n341_), .B0(new_n616_), .B1(new_n570_), .Y(new_n1356_));
  AOI21X1  g01163(.A0(new_n1356_), .A1(new_n1355_), .B0(new_n1354_), .Y(new_n1357_));
  XOR2X1   g01164(.A(new_n1357_), .B(new_n1350_), .Y(new_n1358_));
  AND2X1   g01165(.A(new_n1290_), .B(new_n1281_), .Y(new_n1359_));
  AOI21X1  g01166(.A0(new_n1291_), .A1(new_n1278_), .B0(new_n1359_), .Y(new_n1360_));
  XOR2X1   g01167(.A(new_n1360_), .B(new_n1358_), .Y(new_n1361_));
  OAI21X1  g01168(.A0(new_n1175_), .A1(new_n1174_), .B0(new_n1284_), .Y(new_n1362_));
  AND2X1   g01169(.A(new_n1286_), .B(new_n1362_), .Y(new_n1363_));
  NAND2X1  g01170(.A(new_n1144_), .B(new_n1139_), .Y(new_n1364_));
  NOR2X1   g01171(.A(new_n1144_), .B(new_n1139_), .Y(new_n1365_));
  AOI21X1  g01172(.A0(new_n1268_), .A1(new_n1364_), .B0(new_n1365_), .Y(new_n1366_));
  XOR2X1   g01173(.A(new_n1366_), .B(new_n1363_), .Y(new_n1367_));
  AND2X1   g01174(.A(new_n1234_), .B(new_n1225_), .Y(new_n1368_));
  AND2X1   g01175(.A(new_n1245_), .B(new_n1235_), .Y(new_n1369_));
  OR2X1    g01176(.A(new_n1369_), .B(new_n1368_), .Y(new_n1370_));
  XOR2X1   g01177(.A(new_n1370_), .B(new_n1367_), .Y(new_n1371_));
  XOR2X1   g01178(.A(new_n1371_), .B(new_n1361_), .Y(new_n1372_));
  XOR2X1   g01179(.A(new_n1372_), .B(new_n1344_), .Y(new_n1373_));
  XOR2X1   g01180(.A(new_n1373_), .B(new_n1302_), .Y(new_n1374_));
  AND2X1   g01181(.A(new_n1295_), .B(new_n1214_), .Y(new_n1375_));
  NOR2X1   g01182(.A(new_n1295_), .B(new_n1214_), .Y(new_n1376_));
  INVX1    g01183(.A(new_n1376_), .Y(new_n1377_));
  AOI21X1  g01184(.A0(new_n1298_), .A1(new_n1377_), .B0(new_n1375_), .Y(new_n1378_));
  XOR2X1   g01185(.A(new_n1378_), .B(new_n1374_), .Y(\asquared[28] ));
  NAND2X1  g01186(.A(new_n1341_), .B(new_n1338_), .Y(new_n1380_));
  OAI21X1  g01187(.A0(new_n1342_), .A1(new_n1336_), .B0(new_n1380_), .Y(new_n1381_));
  AND2X1   g01188(.A(\a[20] ), .B(\a[8] ), .Y(new_n1382_));
  NOR3X1   g01189(.A(new_n217_), .B(new_n1326_), .C(new_n1185_), .Y(new_n1383_));
  AOI22X1  g01190(.A0(\a[25] ), .A1(\a[3] ), .B0(\a[24] ), .B1(\a[4] ), .Y(new_n1384_));
  OAI21X1  g01191(.A0(new_n1384_), .A1(new_n1383_), .B0(new_n1382_), .Y(new_n1385_));
  INVX1    g01192(.A(new_n1384_), .Y(new_n1386_));
  AOI21X1  g01193(.A0(new_n1386_), .A1(new_n1382_), .B0(new_n1383_), .Y(new_n1387_));
  NAND2X1  g01194(.A(new_n1387_), .B(new_n1386_), .Y(new_n1388_));
  AND2X1   g01195(.A(new_n1388_), .B(new_n1385_), .Y(new_n1389_));
  NOR2X1   g01196(.A(new_n1334_), .B(new_n1330_), .Y(new_n1390_));
  AOI21X1  g01197(.A0(new_n1328_), .A1(new_n1327_), .B0(new_n1390_), .Y(new_n1391_));
  XOR2X1   g01198(.A(new_n1391_), .B(new_n1389_), .Y(new_n1392_));
  INVX1    g01199(.A(new_n1392_), .Y(new_n1393_));
  AND2X1   g01200(.A(\a[23] ), .B(\a[22] ), .Y(new_n1394_));
  INVX1    g01201(.A(new_n1394_), .Y(new_n1395_));
  INVX1    g01202(.A(new_n1016_), .Y(new_n1396_));
  INVX1    g01203(.A(new_n1154_), .Y(new_n1397_));
  OAI22X1  g01204(.A0(new_n1397_), .A1(new_n376_), .B0(new_n1396_), .B1(new_n678_), .Y(new_n1398_));
  OAI21X1  g01205(.A0(new_n1395_), .A1(new_n444_), .B0(new_n1398_), .Y(new_n1399_));
  AND2X1   g01206(.A(\a[21] ), .B(\a[7] ), .Y(new_n1400_));
  AOI21X1  g01207(.A0(new_n1394_), .A1(new_n295_), .B0(new_n1398_), .Y(new_n1401_));
  OAI22X1  g01208(.A0(new_n1216_), .A1(new_n255_), .B0(new_n1086_), .B1(new_n230_), .Y(new_n1402_));
  AOI22X1  g01209(.A0(new_n1402_), .A1(new_n1401_), .B0(new_n1400_), .B1(new_n1399_), .Y(new_n1403_));
  XOR2X1   g01210(.A(new_n1403_), .B(new_n1393_), .Y(new_n1404_));
  XOR2X1   g01211(.A(new_n1404_), .B(new_n1381_), .Y(new_n1405_));
  INVX1    g01212(.A(new_n1324_), .Y(new_n1406_));
  OR2X1    g01213(.A(new_n1406_), .B(new_n1315_), .Y(new_n1407_));
  INVX1    g01214(.A(new_n1335_), .Y(new_n1408_));
  OAI21X1  g01215(.A0(new_n1408_), .A1(new_n1325_), .B0(new_n1407_), .Y(new_n1409_));
  OAI21X1  g01216(.A0(new_n1265_), .A1(new_n1264_), .B0(new_n1349_), .Y(new_n1410_));
  NOR3X1   g01217(.A(new_n1349_), .B(new_n1265_), .C(new_n1264_), .Y(new_n1411_));
  OAI21X1  g01218(.A0(new_n1357_), .A1(new_n1411_), .B0(new_n1410_), .Y(new_n1412_));
  AND2X1   g01219(.A(\a[27] ), .B(\a[1] ), .Y(new_n1413_));
  XOR2X1   g01220(.A(new_n1413_), .B(new_n639_), .Y(new_n1414_));
  XOR2X1   g01221(.A(new_n1414_), .B(new_n1332_), .Y(new_n1415_));
  XOR2X1   g01222(.A(new_n1415_), .B(new_n1322_), .Y(new_n1416_));
  XOR2X1   g01223(.A(new_n1416_), .B(new_n1412_), .Y(new_n1417_));
  XOR2X1   g01224(.A(new_n1417_), .B(new_n1409_), .Y(new_n1418_));
  XOR2X1   g01225(.A(new_n1418_), .B(new_n1405_), .Y(new_n1419_));
  AND2X1   g01226(.A(new_n1343_), .B(new_n1306_), .Y(new_n1420_));
  AND2X1   g01227(.A(new_n1372_), .B(new_n1344_), .Y(new_n1421_));
  OR2X1    g01228(.A(new_n1421_), .B(new_n1420_), .Y(new_n1422_));
  NAND2X1  g01229(.A(new_n1371_), .B(new_n1361_), .Y(new_n1423_));
  OAI21X1  g01230(.A0(new_n1360_), .A1(new_n1358_), .B0(new_n1423_), .Y(new_n1424_));
  XOR2X1   g01231(.A(new_n1355_), .B(new_n1312_), .Y(new_n1425_));
  AOI21X1  g01232(.A0(new_n1348_), .A1(new_n1345_), .B0(new_n1346_), .Y(new_n1426_));
  XOR2X1   g01233(.A(new_n1426_), .B(new_n1425_), .Y(new_n1427_));
  NOR2X1   g01234(.A(new_n1366_), .B(new_n1363_), .Y(new_n1428_));
  AOI21X1  g01235(.A0(new_n1370_), .A1(new_n1367_), .B0(new_n1428_), .Y(new_n1429_));
  XOR2X1   g01236(.A(new_n1429_), .B(new_n1427_), .Y(new_n1430_));
  INVX1    g01237(.A(\a[28] ), .Y(new_n1431_));
  NOR4X1   g01238(.A(new_n1431_), .B(new_n571_), .C(new_n453_), .D(new_n194_), .Y(new_n1432_));
  AND2X1   g01239(.A(\a[17] ), .B(\a[0] ), .Y(new_n1433_));
  AND2X1   g01240(.A(\a[28] ), .B(\a[11] ), .Y(new_n1434_));
  AOI22X1  g01241(.A0(new_n1434_), .A1(new_n1433_), .B0(new_n792_), .B1(new_n482_), .Y(new_n1435_));
  OR2X1    g01242(.A(new_n1435_), .B(new_n1432_), .Y(new_n1436_));
  INVX1    g01243(.A(new_n1432_), .Y(new_n1437_));
  AND2X1   g01244(.A(new_n1435_), .B(new_n1437_), .Y(new_n1438_));
  OAI22X1  g01245(.A0(new_n1431_), .A1(new_n194_), .B0(new_n571_), .B1(new_n453_), .Y(new_n1439_));
  AND2X1   g01246(.A(\a[17] ), .B(\a[11] ), .Y(new_n1440_));
  AOI22X1  g01247(.A0(new_n1440_), .A1(new_n1436_), .B0(new_n1439_), .B1(new_n1438_), .Y(new_n1441_));
  AND2X1   g01248(.A(\a[26] ), .B(\a[2] ), .Y(new_n1442_));
  INVX1    g01249(.A(new_n1442_), .Y(new_n1443_));
  AOI22X1  g01250(.A0(\a[19] ), .A1(\a[9] ), .B0(\a[18] ), .B1(\a[10] ), .Y(new_n1444_));
  NOR3X1   g01251(.A(new_n735_), .B(new_n752_), .C(new_n675_), .Y(new_n1445_));
  NOR3X1   g01252(.A(new_n1444_), .B(new_n1445_), .C(new_n1443_), .Y(new_n1446_));
  INVX1    g01253(.A(new_n1444_), .Y(new_n1447_));
  AOI21X1  g01254(.A0(new_n1447_), .A1(new_n1442_), .B0(new_n1445_), .Y(new_n1448_));
  INVX1    g01255(.A(new_n1448_), .Y(new_n1449_));
  OAI22X1  g01256(.A0(new_n1449_), .A1(new_n1444_), .B0(new_n1446_), .B1(new_n1443_), .Y(new_n1450_));
  XOR2X1   g01257(.A(new_n1450_), .B(new_n1441_), .Y(new_n1451_));
  AND2X1   g01258(.A(new_n1243_), .B(new_n1232_), .Y(new_n1452_));
  AOI21X1  g01259(.A0(new_n1337_), .A1(new_n1223_), .B0(new_n1452_), .Y(new_n1453_));
  XOR2X1   g01260(.A(new_n1453_), .B(new_n1451_), .Y(new_n1454_));
  XOR2X1   g01261(.A(new_n1454_), .B(new_n1430_), .Y(new_n1455_));
  XOR2X1   g01262(.A(new_n1455_), .B(new_n1424_), .Y(new_n1456_));
  XOR2X1   g01263(.A(new_n1456_), .B(new_n1422_), .Y(new_n1457_));
  XOR2X1   g01264(.A(new_n1457_), .B(new_n1419_), .Y(new_n1458_));
  INVX1    g01265(.A(new_n1373_), .Y(new_n1459_));
  NOR2X1   g01266(.A(new_n1459_), .B(new_n1302_), .Y(new_n1460_));
  INVX1    g01267(.A(new_n1460_), .Y(new_n1461_));
  AND2X1   g01268(.A(new_n1459_), .B(new_n1302_), .Y(new_n1462_));
  OAI21X1  g01269(.A0(new_n1378_), .A1(new_n1462_), .B0(new_n1461_), .Y(new_n1463_));
  XOR2X1   g01270(.A(new_n1463_), .B(new_n1458_), .Y(\asquared[29] ));
  AND2X1   g01271(.A(new_n1455_), .B(new_n1424_), .Y(new_n1465_));
  AOI21X1  g01272(.A0(new_n1456_), .A1(new_n1422_), .B0(new_n1465_), .Y(new_n1466_));
  NOR2X1   g01273(.A(new_n1429_), .B(new_n1427_), .Y(new_n1467_));
  AOI21X1  g01274(.A0(new_n1454_), .A1(new_n1430_), .B0(new_n1467_), .Y(new_n1468_));
  AND2X1   g01275(.A(new_n1416_), .B(new_n1412_), .Y(new_n1469_));
  AOI21X1  g01276(.A0(new_n1417_), .A1(new_n1409_), .B0(new_n1469_), .Y(new_n1470_));
  XOR2X1   g01277(.A(new_n1470_), .B(new_n1468_), .Y(new_n1471_));
  INVX1    g01278(.A(new_n1450_), .Y(new_n1472_));
  OR2X1    g01279(.A(new_n1472_), .B(new_n1441_), .Y(new_n1473_));
  OAI21X1  g01280(.A0(new_n1453_), .A1(new_n1451_), .B0(new_n1473_), .Y(new_n1474_));
  OR2X1    g01281(.A(new_n1391_), .B(new_n1389_), .Y(new_n1475_));
  OAI21X1  g01282(.A0(new_n1403_), .A1(new_n1393_), .B0(new_n1475_), .Y(new_n1476_));
  XOR2X1   g01283(.A(new_n1476_), .B(new_n1474_), .Y(new_n1477_));
  XOR2X1   g01284(.A(new_n1449_), .B(new_n1438_), .Y(new_n1478_));
  AND2X1   g01285(.A(new_n1413_), .B(new_n639_), .Y(new_n1479_));
  AOI22X1  g01286(.A0(\a[29] ), .A1(\a[0] ), .B0(\a[27] ), .B1(\a[2] ), .Y(new_n1480_));
  INVX1    g01287(.A(new_n1480_), .Y(new_n1481_));
  NAND4X1  g01288(.A(\a[29] ), .B(\a[27] ), .C(\a[2] ), .D(\a[0] ), .Y(new_n1482_));
  NAND3X1  g01289(.A(new_n1482_), .B(new_n1481_), .C(new_n1479_), .Y(new_n1483_));
  AND2X1   g01290(.A(\a[29] ), .B(\a[27] ), .Y(new_n1484_));
  AOI22X1  g01291(.A0(new_n1484_), .A1(new_n197_), .B0(new_n1481_), .B1(new_n1479_), .Y(new_n1485_));
  AOI22X1  g01292(.A0(new_n1485_), .A1(new_n1481_), .B0(new_n1483_), .B1(new_n1479_), .Y(new_n1486_));
  XOR2X1   g01293(.A(new_n1486_), .B(new_n1478_), .Y(new_n1487_));
  XOR2X1   g01294(.A(new_n1487_), .B(new_n1477_), .Y(new_n1488_));
  XOR2X1   g01295(.A(new_n1488_), .B(new_n1471_), .Y(new_n1489_));
  AND2X1   g01296(.A(new_n1404_), .B(new_n1381_), .Y(new_n1490_));
  AOI21X1  g01297(.A0(new_n1418_), .A1(new_n1405_), .B0(new_n1490_), .Y(new_n1491_));
  AND2X1   g01298(.A(new_n1414_), .B(new_n1331_), .Y(new_n1492_));
  INVX1    g01299(.A(new_n1492_), .Y(new_n1493_));
  OR2X1    g01300(.A(new_n1415_), .B(new_n1322_), .Y(new_n1494_));
  AND2X1   g01301(.A(new_n1494_), .B(new_n1493_), .Y(new_n1495_));
  INVX1    g01302(.A(new_n1495_), .Y(new_n1496_));
  AND2X1   g01303(.A(\a[23] ), .B(\a[6] ), .Y(new_n1497_));
  NOR4X1   g01304(.A(new_n571_), .B(new_n549_), .C(new_n490_), .D(new_n591_), .Y(new_n1498_));
  AOI22X1  g01305(.A0(\a[16] ), .A1(\a[13] ), .B0(\a[15] ), .B1(\a[14] ), .Y(new_n1499_));
  OR4X1    g01306(.A(new_n1499_), .B(new_n1498_), .C(new_n1216_), .D(new_n230_), .Y(new_n1500_));
  NOR3X1   g01307(.A(new_n1499_), .B(new_n1498_), .C(new_n1497_), .Y(new_n1501_));
  AOI21X1  g01308(.A0(new_n1500_), .A1(new_n1497_), .B0(new_n1501_), .Y(new_n1502_));
  XOR2X1   g01309(.A(new_n1502_), .B(new_n1496_), .Y(new_n1503_));
  NOR2X1   g01310(.A(new_n1355_), .B(new_n1312_), .Y(new_n1504_));
  INVX1    g01311(.A(new_n1426_), .Y(new_n1505_));
  AOI21X1  g01312(.A0(new_n1505_), .A1(new_n1425_), .B0(new_n1504_), .Y(new_n1506_));
  XOR2X1   g01313(.A(new_n1506_), .B(new_n1503_), .Y(new_n1507_));
  AOI22X1  g01314(.A0(\a[26] ), .A1(\a[3] ), .B0(\a[21] ), .B1(\a[8] ), .Y(new_n1508_));
  AND2X1   g01315(.A(\a[17] ), .B(\a[12] ), .Y(new_n1509_));
  INVX1    g01316(.A(new_n1509_), .Y(new_n1510_));
  NOR4X1   g01317(.A(new_n1263_), .B(new_n1098_), .C(new_n413_), .D(new_n223_), .Y(new_n1511_));
  NOR3X1   g01318(.A(new_n1510_), .B(new_n1511_), .C(new_n1508_), .Y(new_n1512_));
  INVX1    g01319(.A(new_n1508_), .Y(new_n1513_));
  AOI21X1  g01320(.A0(new_n1509_), .A1(new_n1513_), .B0(new_n1511_), .Y(new_n1514_));
  INVX1    g01321(.A(new_n1514_), .Y(new_n1515_));
  OAI22X1  g01322(.A0(new_n1515_), .A1(new_n1508_), .B0(new_n1512_), .B1(new_n1510_), .Y(new_n1516_));
  INVX1    g01323(.A(new_n1002_), .Y(new_n1517_));
  INVX1    g01324(.A(new_n855_), .Y(new_n1518_));
  INVX1    g01325(.A(new_n813_), .Y(new_n1519_));
  INVX1    g01326(.A(new_n992_), .Y(new_n1520_));
  INVX1    g01327(.A(new_n1099_), .Y(new_n1521_));
  OAI22X1  g01328(.A0(new_n1521_), .A1(new_n735_), .B0(new_n1520_), .B1(new_n1519_), .Y(new_n1522_));
  OAI21X1  g01329(.A0(new_n1518_), .A1(new_n1517_), .B0(new_n1522_), .Y(new_n1523_));
  AND2X1   g01330(.A(\a[20] ), .B(\a[9] ), .Y(new_n1524_));
  AOI21X1  g01331(.A0(new_n855_), .A1(new_n1002_), .B0(new_n1522_), .Y(new_n1525_));
  OAI22X1  g01332(.A0(new_n752_), .A1(new_n570_), .B0(new_n675_), .B1(new_n488_), .Y(new_n1526_));
  AOI22X1  g01333(.A0(new_n1526_), .A1(new_n1525_), .B0(new_n1524_), .B1(new_n1523_), .Y(new_n1527_));
  XOR2X1   g01334(.A(new_n1527_), .B(new_n1516_), .Y(new_n1528_));
  AND2X1   g01335(.A(\a[25] ), .B(\a[4] ), .Y(new_n1529_));
  AND2X1   g01336(.A(\a[24] ), .B(\a[22] ), .Y(new_n1530_));
  INVX1    g01337(.A(new_n1530_), .Y(new_n1531_));
  AND2X1   g01338(.A(\a[25] ), .B(\a[24] ), .Y(new_n1532_));
  AND2X1   g01339(.A(new_n1532_), .B(new_n218_), .Y(new_n1533_));
  NOR4X1   g01340(.A(new_n1326_), .B(new_n1086_), .C(new_n532_), .D(new_n340_), .Y(new_n1534_));
  OAI22X1  g01341(.A0(new_n1534_), .A1(new_n1533_), .B0(new_n1531_), .B1(new_n678_), .Y(new_n1535_));
  OAI21X1  g01342(.A0(new_n1531_), .A1(new_n678_), .B0(new_n1535_), .Y(new_n1536_));
  INVX1    g01343(.A(new_n1536_), .Y(new_n1537_));
  OAI22X1  g01344(.A0(new_n1185_), .A1(new_n255_), .B0(new_n1086_), .B1(new_n532_), .Y(new_n1538_));
  AOI22X1  g01345(.A0(new_n1538_), .A1(new_n1537_), .B0(new_n1535_), .B1(new_n1529_), .Y(new_n1539_));
  XOR2X1   g01346(.A(new_n1539_), .B(new_n1528_), .Y(new_n1540_));
  INVX1    g01347(.A(new_n1401_), .Y(new_n1541_));
  NAND3X1  g01348(.A(\a[28] ), .B(\a[15] ), .C(\a[1] ), .Y(new_n1542_));
  AND2X1   g01349(.A(\a[28] ), .B(\a[1] ), .Y(new_n1543_));
  OAI21X1  g01350(.A0(new_n1543_), .A1(\a[15] ), .B0(new_n1542_), .Y(new_n1544_));
  XOR2X1   g01351(.A(new_n1544_), .B(new_n1541_), .Y(new_n1545_));
  XOR2X1   g01352(.A(new_n1545_), .B(new_n1387_), .Y(new_n1546_));
  XOR2X1   g01353(.A(new_n1546_), .B(new_n1540_), .Y(new_n1547_));
  XOR2X1   g01354(.A(new_n1547_), .B(new_n1507_), .Y(new_n1548_));
  NAND2X1  g01355(.A(new_n1548_), .B(new_n1491_), .Y(new_n1549_));
  INVX1    g01356(.A(new_n1491_), .Y(new_n1550_));
  XOR2X1   g01357(.A(new_n1548_), .B(new_n1550_), .Y(new_n1551_));
  NAND2X1  g01358(.A(new_n1548_), .B(new_n1550_), .Y(new_n1552_));
  AOI21X1  g01359(.A0(new_n1552_), .A1(new_n1550_), .B0(new_n1489_), .Y(new_n1553_));
  AOI22X1  g01360(.A0(new_n1553_), .A1(new_n1549_), .B0(new_n1551_), .B1(new_n1489_), .Y(new_n1554_));
  XOR2X1   g01361(.A(new_n1554_), .B(new_n1466_), .Y(new_n1555_));
  NOR2X1   g01362(.A(new_n1457_), .B(new_n1419_), .Y(new_n1556_));
  INVX1    g01363(.A(new_n1556_), .Y(new_n1557_));
  AND2X1   g01364(.A(new_n1457_), .B(new_n1419_), .Y(new_n1558_));
  AOI21X1  g01365(.A0(new_n1463_), .A1(new_n1557_), .B0(new_n1558_), .Y(new_n1559_));
  XOR2X1   g01366(.A(new_n1559_), .B(new_n1555_), .Y(\asquared[30] ));
  AND2X1   g01367(.A(new_n1548_), .B(new_n1550_), .Y(new_n1561_));
  AOI21X1  g01368(.A0(new_n1551_), .A1(new_n1489_), .B0(new_n1561_), .Y(new_n1562_));
  INVX1    g01369(.A(new_n1562_), .Y(new_n1563_));
  AND2X1   g01370(.A(\a[30] ), .B(\a[0] ), .Y(new_n1564_));
  XOR2X1   g01371(.A(new_n1564_), .B(new_n1542_), .Y(new_n1565_));
  NAND2X1  g01372(.A(\a[29] ), .B(\a[1] ), .Y(new_n1566_));
  XOR2X1   g01373(.A(new_n1566_), .B(new_n690_), .Y(new_n1567_));
  XOR2X1   g01374(.A(new_n1567_), .B(new_n1565_), .Y(new_n1568_));
  OR2X1    g01375(.A(new_n1544_), .B(new_n1401_), .Y(new_n1569_));
  OAI21X1  g01376(.A0(new_n1545_), .A1(new_n1387_), .B0(new_n1569_), .Y(new_n1570_));
  XOR2X1   g01377(.A(new_n1570_), .B(new_n1568_), .Y(new_n1571_));
  INVX1    g01378(.A(new_n1571_), .Y(new_n1572_));
  OR2X1    g01379(.A(new_n1448_), .B(new_n1438_), .Y(new_n1573_));
  OAI21X1  g01380(.A0(new_n1486_), .A1(new_n1478_), .B0(new_n1573_), .Y(new_n1574_));
  XOR2X1   g01381(.A(new_n1574_), .B(new_n1572_), .Y(new_n1575_));
  AND2X1   g01382(.A(new_n1546_), .B(new_n1540_), .Y(new_n1576_));
  AOI21X1  g01383(.A0(new_n1547_), .A1(new_n1507_), .B0(new_n1576_), .Y(new_n1577_));
  XOR2X1   g01384(.A(new_n1577_), .B(new_n1575_), .Y(new_n1578_));
  NOR3X1   g01385(.A(new_n1499_), .B(new_n1216_), .C(new_n230_), .Y(new_n1579_));
  NOR2X1   g01386(.A(new_n1579_), .B(new_n1498_), .Y(new_n1580_));
  XOR2X1   g01387(.A(new_n1536_), .B(new_n1580_), .Y(new_n1581_));
  AND2X1   g01388(.A(\a[17] ), .B(\a[13] ), .Y(new_n1582_));
  NOR4X1   g01389(.A(new_n1431_), .B(new_n1098_), .C(new_n341_), .D(new_n200_), .Y(new_n1583_));
  AOI22X1  g01390(.A0(\a[28] ), .A1(\a[2] ), .B0(\a[21] ), .B1(\a[9] ), .Y(new_n1584_));
  OR4X1    g01391(.A(new_n1584_), .B(new_n1583_), .C(new_n616_), .D(new_n591_), .Y(new_n1585_));
  NOR3X1   g01392(.A(new_n1584_), .B(new_n1583_), .C(new_n1582_), .Y(new_n1586_));
  AOI21X1  g01393(.A0(new_n1585_), .A1(new_n1582_), .B0(new_n1586_), .Y(new_n1587_));
  XOR2X1   g01394(.A(new_n1587_), .B(new_n1581_), .Y(new_n1588_));
  INVX1    g01395(.A(new_n1516_), .Y(new_n1589_));
  OR2X1    g01396(.A(new_n1527_), .B(new_n1589_), .Y(new_n1590_));
  OAI21X1  g01397(.A0(new_n1539_), .A1(new_n1528_), .B0(new_n1590_), .Y(new_n1591_));
  XOR2X1   g01398(.A(new_n1591_), .B(new_n1588_), .Y(new_n1592_));
  INVX1    g01399(.A(new_n1485_), .Y(new_n1593_));
  XOR2X1   g01400(.A(new_n1525_), .B(new_n1514_), .Y(new_n1594_));
  XOR2X1   g01401(.A(new_n1594_), .B(new_n1593_), .Y(new_n1595_));
  XOR2X1   g01402(.A(new_n1595_), .B(new_n1592_), .Y(new_n1596_));
  XOR2X1   g01403(.A(new_n1596_), .B(new_n1578_), .Y(new_n1597_));
  NAND2X1  g01404(.A(new_n1488_), .B(new_n1471_), .Y(new_n1598_));
  OAI21X1  g01405(.A0(new_n1470_), .A1(new_n1468_), .B0(new_n1598_), .Y(new_n1599_));
  NOR4X1   g01406(.A(new_n1263_), .B(new_n1086_), .C(new_n413_), .D(new_n340_), .Y(new_n1600_));
  NAND4X1  g01407(.A(\a[27] ), .B(\a[26] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n1601_));
  NAND4X1  g01408(.A(\a[27] ), .B(\a[22] ), .C(\a[8] ), .D(\a[3] ), .Y(new_n1602_));
  AOI21X1  g01409(.A0(new_n1602_), .A1(new_n1601_), .B0(new_n1600_), .Y(new_n1603_));
  OR2X1    g01410(.A(new_n1603_), .B(new_n1600_), .Y(new_n1604_));
  AOI22X1  g01411(.A0(\a[26] ), .A1(\a[4] ), .B0(\a[22] ), .B1(\a[8] ), .Y(new_n1605_));
  NAND2X1  g01412(.A(\a[27] ), .B(\a[3] ), .Y(new_n1606_));
  OAI22X1  g01413(.A0(new_n1606_), .A1(new_n1603_), .B0(new_n1605_), .B1(new_n1604_), .Y(new_n1607_));
  NAND4X1  g01414(.A(\a[25] ), .B(\a[23] ), .C(\a[7] ), .D(\a[5] ), .Y(new_n1608_));
  NAND4X1  g01415(.A(\a[25] ), .B(\a[24] ), .C(\a[6] ), .D(\a[5] ), .Y(new_n1609_));
  AOI22X1  g01416(.A0(new_n1609_), .A1(new_n1608_), .B0(new_n1219_), .B1(new_n375_), .Y(new_n1610_));
  NAND2X1  g01417(.A(\a[25] ), .B(\a[5] ), .Y(new_n1611_));
  AOI21X1  g01418(.A0(new_n1219_), .A1(new_n375_), .B0(new_n1610_), .Y(new_n1612_));
  INVX1    g01419(.A(new_n1612_), .Y(new_n1613_));
  AOI22X1  g01420(.A0(\a[24] ), .A1(\a[6] ), .B0(\a[23] ), .B1(\a[7] ), .Y(new_n1614_));
  OAI22X1  g01421(.A0(new_n1614_), .A1(new_n1613_), .B0(new_n1611_), .B1(new_n1610_), .Y(new_n1615_));
  XOR2X1   g01422(.A(new_n1615_), .B(new_n1607_), .Y(new_n1616_));
  AOI22X1  g01423(.A0(new_n1099_), .A1(new_n1002_), .B0(new_n992_), .B1(new_n396_), .Y(new_n1617_));
  AOI21X1  g01424(.A0(new_n855_), .A1(new_n482_), .B0(new_n1617_), .Y(new_n1618_));
  AND2X1   g01425(.A(\a[20] ), .B(\a[10] ), .Y(new_n1619_));
  INVX1    g01426(.A(new_n1619_), .Y(new_n1620_));
  AOI22X1  g01427(.A0(\a[19] ), .A1(\a[11] ), .B0(\a[18] ), .B1(\a[12] ), .Y(new_n1621_));
  OAI22X1  g01428(.A0(new_n1521_), .A1(new_n1517_), .B0(new_n1520_), .B1(new_n543_), .Y(new_n1622_));
  AOI21X1  g01429(.A0(new_n855_), .A1(new_n482_), .B0(new_n1622_), .Y(new_n1623_));
  INVX1    g01430(.A(new_n1623_), .Y(new_n1624_));
  OAI22X1  g01431(.A0(new_n1624_), .A1(new_n1621_), .B0(new_n1620_), .B1(new_n1618_), .Y(new_n1625_));
  XOR2X1   g01432(.A(new_n1625_), .B(new_n1616_), .Y(new_n1626_));
  INVX1    g01433(.A(new_n1626_), .Y(new_n1627_));
  OR2X1    g01434(.A(new_n1502_), .B(new_n1495_), .Y(new_n1628_));
  OAI21X1  g01435(.A0(new_n1506_), .A1(new_n1503_), .B0(new_n1628_), .Y(new_n1629_));
  XOR2X1   g01436(.A(new_n1629_), .B(new_n1627_), .Y(new_n1630_));
  AND2X1   g01437(.A(new_n1476_), .B(new_n1474_), .Y(new_n1631_));
  AOI21X1  g01438(.A0(new_n1487_), .A1(new_n1477_), .B0(new_n1631_), .Y(new_n1632_));
  XOR2X1   g01439(.A(new_n1632_), .B(new_n1630_), .Y(new_n1633_));
  XOR2X1   g01440(.A(new_n1633_), .B(new_n1599_), .Y(new_n1634_));
  XOR2X1   g01441(.A(new_n1634_), .B(new_n1597_), .Y(new_n1635_));
  XOR2X1   g01442(.A(new_n1635_), .B(new_n1563_), .Y(new_n1636_));
  INVX1    g01443(.A(new_n1466_), .Y(new_n1637_));
  NAND2X1  g01444(.A(new_n1554_), .B(new_n1637_), .Y(new_n1638_));
  NOR2X1   g01445(.A(new_n1554_), .B(new_n1637_), .Y(new_n1639_));
  OAI21X1  g01446(.A0(new_n1559_), .A1(new_n1639_), .B0(new_n1638_), .Y(new_n1640_));
  XOR2X1   g01447(.A(new_n1640_), .B(new_n1636_), .Y(\asquared[31] ));
  AND2X1   g01448(.A(new_n1633_), .B(new_n1599_), .Y(new_n1642_));
  AOI21X1  g01449(.A0(new_n1634_), .A1(new_n1597_), .B0(new_n1642_), .Y(new_n1643_));
  NOR2X1   g01450(.A(new_n1577_), .B(new_n1575_), .Y(new_n1644_));
  AOI21X1  g01451(.A0(new_n1596_), .A1(new_n1578_), .B0(new_n1644_), .Y(new_n1645_));
  INVX1    g01452(.A(new_n1645_), .Y(new_n1646_));
  AND2X1   g01453(.A(new_n1591_), .B(new_n1588_), .Y(new_n1647_));
  AND2X1   g01454(.A(new_n1595_), .B(new_n1592_), .Y(new_n1648_));
  OR2X1    g01455(.A(new_n1648_), .B(new_n1647_), .Y(new_n1649_));
  AND2X1   g01456(.A(\a[26] ), .B(\a[24] ), .Y(new_n1650_));
  INVX1    g01457(.A(new_n1650_), .Y(new_n1651_));
  INVX1    g01458(.A(new_n1219_), .Y(new_n1652_));
  NAND4X1  g01459(.A(\a[26] ), .B(\a[23] ), .C(\a[8] ), .D(\a[5] ), .Y(new_n1653_));
  OAI21X1  g01460(.A0(new_n1652_), .A1(new_n445_), .B0(new_n1653_), .Y(new_n1654_));
  OAI21X1  g01461(.A0(new_n1651_), .A1(new_n678_), .B0(new_n1654_), .Y(new_n1655_));
  NOR3X1   g01462(.A(new_n678_), .B(new_n1263_), .C(new_n1185_), .Y(new_n1656_));
  NOR2X1   g01463(.A(new_n1654_), .B(new_n1656_), .Y(new_n1657_));
  OAI22X1  g01464(.A0(new_n1263_), .A1(new_n255_), .B0(new_n1185_), .B1(new_n532_), .Y(new_n1658_));
  AND2X1   g01465(.A(\a[23] ), .B(\a[8] ), .Y(new_n1659_));
  AOI22X1  g01466(.A0(new_n1659_), .A1(new_n1655_), .B0(new_n1658_), .B1(new_n1657_), .Y(new_n1660_));
  AND2X1   g01467(.A(\a[25] ), .B(\a[6] ), .Y(new_n1661_));
  INVX1    g01468(.A(new_n1661_), .Y(new_n1662_));
  AOI22X1  g01469(.A0(\a[17] ), .A1(\a[14] ), .B0(\a[16] ), .B1(\a[15] ), .Y(new_n1663_));
  AND2X1   g01470(.A(new_n792_), .B(new_n691_), .Y(new_n1664_));
  NOR3X1   g01471(.A(new_n1663_), .B(new_n1664_), .C(new_n1662_), .Y(new_n1665_));
  INVX1    g01472(.A(new_n1663_), .Y(new_n1666_));
  AOI21X1  g01473(.A0(new_n1666_), .A1(new_n1661_), .B0(new_n1664_), .Y(new_n1667_));
  INVX1    g01474(.A(new_n1667_), .Y(new_n1668_));
  OAI22X1  g01475(.A0(new_n1668_), .A1(new_n1663_), .B0(new_n1665_), .B1(new_n1662_), .Y(new_n1669_));
  XOR2X1   g01476(.A(new_n1669_), .B(new_n1660_), .Y(new_n1670_));
  AND2X1   g01477(.A(\a[28] ), .B(\a[27] ), .Y(new_n1671_));
  INVX1    g01478(.A(new_n1671_), .Y(new_n1672_));
  INVX1    g01479(.A(new_n1484_), .Y(new_n1673_));
  AND2X1   g01480(.A(\a[29] ), .B(\a[28] ), .Y(new_n1674_));
  INVX1    g01481(.A(new_n1674_), .Y(new_n1675_));
  OAI22X1  g01482(.A0(new_n1675_), .A1(new_n249_), .B0(new_n1673_), .B1(new_n584_), .Y(new_n1676_));
  OAI21X1  g01483(.A0(new_n1672_), .A1(new_n217_), .B0(new_n1676_), .Y(new_n1677_));
  AND2X1   g01484(.A(\a[29] ), .B(\a[2] ), .Y(new_n1678_));
  INVX1    g01485(.A(\a[27] ), .Y(new_n1679_));
  OAI22X1  g01486(.A0(new_n1431_), .A1(new_n223_), .B0(new_n1679_), .B1(new_n340_), .Y(new_n1680_));
  AOI21X1  g01487(.A0(new_n1671_), .A1(new_n294_), .B0(new_n1676_), .Y(new_n1681_));
  AOI22X1  g01488(.A0(new_n1681_), .A1(new_n1680_), .B0(new_n1678_), .B1(new_n1677_), .Y(new_n1682_));
  XOR2X1   g01489(.A(new_n1682_), .B(new_n1670_), .Y(new_n1683_));
  INVX1    g01490(.A(\a[30] ), .Y(new_n1684_));
  NOR3X1   g01491(.A(new_n1542_), .B(new_n1684_), .C(new_n194_), .Y(new_n1685_));
  NOR2X1   g01492(.A(new_n1567_), .B(new_n1565_), .Y(new_n1686_));
  NOR2X1   g01493(.A(new_n1686_), .B(new_n1685_), .Y(new_n1687_));
  NAND4X1  g01494(.A(\a[20] ), .B(\a[18] ), .C(\a[13] ), .D(\a[11] ), .Y(new_n1688_));
  NAND4X1  g01495(.A(\a[20] ), .B(\a[19] ), .C(\a[12] ), .D(\a[11] ), .Y(new_n1689_));
  AOI22X1  g01496(.A0(new_n1689_), .A1(new_n1688_), .B0(new_n855_), .B1(new_n586_), .Y(new_n1690_));
  NAND2X1  g01497(.A(\a[20] ), .B(\a[11] ), .Y(new_n1691_));
  NAND4X1  g01498(.A(\a[19] ), .B(\a[18] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n1692_));
  NAND3X1  g01499(.A(new_n1689_), .B(new_n1688_), .C(new_n1692_), .Y(new_n1693_));
  AOI22X1  g01500(.A0(\a[19] ), .A1(\a[12] ), .B0(\a[18] ), .B1(\a[13] ), .Y(new_n1694_));
  OAI22X1  g01501(.A0(new_n1694_), .A1(new_n1693_), .B0(new_n1691_), .B1(new_n1690_), .Y(new_n1695_));
  NAND2X1  g01502(.A(new_n1695_), .B(new_n1687_), .Y(new_n1696_));
  NAND2X1  g01503(.A(\a[31] ), .B(\a[22] ), .Y(new_n1697_));
  NOR3X1   g01504(.A(new_n1697_), .B(new_n341_), .C(new_n194_), .Y(new_n1698_));
  AND2X1   g01505(.A(\a[31] ), .B(\a[10] ), .Y(new_n1699_));
  AOI22X1  g01506(.A0(new_n1699_), .A1(new_n891_), .B0(new_n1154_), .B1(new_n881_), .Y(new_n1700_));
  OR2X1    g01507(.A(new_n1700_), .B(new_n1698_), .Y(new_n1701_));
  INVX1    g01508(.A(new_n1698_), .Y(new_n1702_));
  AND2X1   g01509(.A(new_n1700_), .B(new_n1702_), .Y(new_n1703_));
  INVX1    g01510(.A(\a[31] ), .Y(new_n1704_));
  OAI22X1  g01511(.A0(new_n1704_), .A1(new_n194_), .B0(new_n1086_), .B1(new_n341_), .Y(new_n1705_));
  AND2X1   g01512(.A(\a[21] ), .B(\a[10] ), .Y(new_n1706_));
  AOI22X1  g01513(.A0(new_n1706_), .A1(new_n1701_), .B0(new_n1705_), .B1(new_n1703_), .Y(new_n1707_));
  OR2X1    g01514(.A(new_n1695_), .B(new_n1687_), .Y(new_n1708_));
  AOI21X1  g01515(.A0(new_n1696_), .A1(new_n1708_), .B0(new_n1707_), .Y(new_n1709_));
  AND2X1   g01516(.A(new_n1708_), .B(new_n1707_), .Y(new_n1710_));
  AOI21X1  g01517(.A0(new_n1710_), .A1(new_n1696_), .B0(new_n1709_), .Y(new_n1711_));
  XOR2X1   g01518(.A(new_n1711_), .B(new_n1683_), .Y(new_n1712_));
  XOR2X1   g01519(.A(new_n1712_), .B(new_n1649_), .Y(new_n1713_));
  XOR2X1   g01520(.A(new_n1713_), .B(new_n1646_), .Y(new_n1714_));
  NAND2X1  g01521(.A(new_n1629_), .B(new_n1626_), .Y(new_n1715_));
  OAI21X1  g01522(.A0(new_n1632_), .A1(new_n1630_), .B0(new_n1715_), .Y(new_n1716_));
  INVX1    g01523(.A(new_n1580_), .Y(new_n1717_));
  NOR2X1   g01524(.A(new_n1587_), .B(new_n1581_), .Y(new_n1718_));
  AOI21X1  g01525(.A0(new_n1536_), .A1(new_n1717_), .B0(new_n1718_), .Y(new_n1719_));
  NOR2X1   g01526(.A(new_n1525_), .B(new_n1514_), .Y(new_n1720_));
  AOI21X1  g01527(.A0(new_n1594_), .A1(new_n1593_), .B0(new_n1720_), .Y(new_n1721_));
  XOR2X1   g01528(.A(new_n1721_), .B(new_n1719_), .Y(new_n1722_));
  NAND4X1  g01529(.A(\a[29] ), .B(\a[16] ), .C(\a[14] ), .D(\a[1] ), .Y(new_n1723_));
  AND2X1   g01530(.A(\a[30] ), .B(\a[1] ), .Y(new_n1724_));
  XOR2X1   g01531(.A(new_n1724_), .B(\a[16] ), .Y(new_n1725_));
  XOR2X1   g01532(.A(new_n1725_), .B(new_n1723_), .Y(new_n1726_));
  XOR2X1   g01533(.A(new_n1726_), .B(new_n1612_), .Y(new_n1727_));
  XOR2X1   g01534(.A(new_n1727_), .B(new_n1722_), .Y(new_n1728_));
  XOR2X1   g01535(.A(new_n1728_), .B(new_n1716_), .Y(new_n1729_));
  NOR3X1   g01536(.A(new_n1584_), .B(new_n616_), .C(new_n591_), .Y(new_n1730_));
  NOR2X1   g01537(.A(new_n1730_), .B(new_n1583_), .Y(new_n1731_));
  INVX1    g01538(.A(new_n1731_), .Y(new_n1732_));
  XOR2X1   g01539(.A(new_n1604_), .B(new_n1732_), .Y(new_n1733_));
  XOR2X1   g01540(.A(new_n1733_), .B(new_n1623_), .Y(new_n1734_));
  AND2X1   g01541(.A(new_n1615_), .B(new_n1607_), .Y(new_n1735_));
  AOI21X1  g01542(.A0(new_n1625_), .A1(new_n1616_), .B0(new_n1735_), .Y(new_n1736_));
  XOR2X1   g01543(.A(new_n1736_), .B(new_n1734_), .Y(new_n1737_));
  AND2X1   g01544(.A(new_n1570_), .B(new_n1568_), .Y(new_n1738_));
  AND2X1   g01545(.A(new_n1574_), .B(new_n1571_), .Y(new_n1739_));
  OR2X1    g01546(.A(new_n1739_), .B(new_n1738_), .Y(new_n1740_));
  XOR2X1   g01547(.A(new_n1740_), .B(new_n1737_), .Y(new_n1741_));
  XOR2X1   g01548(.A(new_n1741_), .B(new_n1729_), .Y(new_n1742_));
  XOR2X1   g01549(.A(new_n1742_), .B(new_n1714_), .Y(new_n1743_));
  XOR2X1   g01550(.A(new_n1743_), .B(new_n1643_), .Y(new_n1744_));
  AND2X1   g01551(.A(new_n1635_), .B(new_n1563_), .Y(new_n1745_));
  OR2X1    g01552(.A(new_n1635_), .B(new_n1563_), .Y(new_n1746_));
  AOI21X1  g01553(.A0(new_n1640_), .A1(new_n1746_), .B0(new_n1745_), .Y(new_n1747_));
  XOR2X1   g01554(.A(new_n1747_), .B(new_n1744_), .Y(\asquared[32] ));
  INVX1    g01555(.A(new_n1743_), .Y(new_n1749_));
  OR2X1    g01556(.A(new_n1749_), .B(new_n1643_), .Y(new_n1750_));
  AND2X1   g01557(.A(new_n1749_), .B(new_n1643_), .Y(new_n1751_));
  OAI21X1  g01558(.A0(new_n1747_), .A1(new_n1751_), .B0(new_n1750_), .Y(new_n1752_));
  AND2X1   g01559(.A(new_n1713_), .B(new_n1646_), .Y(new_n1753_));
  AND2X1   g01560(.A(new_n1742_), .B(new_n1714_), .Y(new_n1754_));
  OR2X1    g01561(.A(new_n1754_), .B(new_n1753_), .Y(new_n1755_));
  AND2X1   g01562(.A(new_n1728_), .B(new_n1716_), .Y(new_n1756_));
  AND2X1   g01563(.A(new_n1741_), .B(new_n1729_), .Y(new_n1757_));
  OR2X1    g01564(.A(new_n1757_), .B(new_n1756_), .Y(new_n1758_));
  NOR2X1   g01565(.A(new_n1736_), .B(new_n1734_), .Y(new_n1759_));
  AOI21X1  g01566(.A0(new_n1740_), .A1(new_n1737_), .B0(new_n1759_), .Y(new_n1760_));
  AOI22X1  g01567(.A0(\a[28] ), .A1(\a[4] ), .B0(\a[27] ), .B1(\a[5] ), .Y(new_n1761_));
  AND2X1   g01568(.A(\a[23] ), .B(\a[9] ), .Y(new_n1762_));
  INVX1    g01569(.A(new_n1762_), .Y(new_n1763_));
  AND2X1   g01570(.A(new_n1671_), .B(new_n218_), .Y(new_n1764_));
  NOR3X1   g01571(.A(new_n1763_), .B(new_n1764_), .C(new_n1761_), .Y(new_n1765_));
  INVX1    g01572(.A(new_n1761_), .Y(new_n1766_));
  AOI21X1  g01573(.A0(new_n1762_), .A1(new_n1766_), .B0(new_n1764_), .Y(new_n1767_));
  INVX1    g01574(.A(new_n1767_), .Y(new_n1768_));
  OAI22X1  g01575(.A0(new_n1768_), .A1(new_n1761_), .B0(new_n1765_), .B1(new_n1763_), .Y(new_n1769_));
  AND2X1   g01576(.A(\a[26] ), .B(\a[25] ), .Y(new_n1770_));
  INVX1    g01577(.A(new_n1770_), .Y(new_n1771_));
  INVX1    g01578(.A(new_n1532_), .Y(new_n1772_));
  OAI22X1  g01579(.A0(new_n1651_), .A1(new_n280_), .B0(new_n1772_), .B1(new_n445_), .Y(new_n1773_));
  OAI21X1  g01580(.A0(new_n1771_), .A1(new_n376_), .B0(new_n1773_), .Y(new_n1774_));
  AND2X1   g01581(.A(\a[24] ), .B(\a[8] ), .Y(new_n1775_));
  AOI21X1  g01582(.A0(new_n1770_), .A1(new_n375_), .B0(new_n1773_), .Y(new_n1776_));
  OAI22X1  g01583(.A0(new_n1263_), .A1(new_n230_), .B0(new_n1326_), .B1(new_n532_), .Y(new_n1777_));
  AOI22X1  g01584(.A0(new_n1777_), .A1(new_n1776_), .B0(new_n1775_), .B1(new_n1774_), .Y(new_n1778_));
  XOR2X1   g01585(.A(new_n1778_), .B(new_n1769_), .Y(new_n1779_));
  INVX1    g01586(.A(new_n1779_), .Y(new_n1780_));
  OR4X1    g01587(.A(new_n1724_), .B(new_n1566_), .C(new_n571_), .D(new_n490_), .Y(new_n1781_));
  OAI21X1  g01588(.A0(new_n1726_), .A1(new_n1612_), .B0(new_n1781_), .Y(new_n1782_));
  XOR2X1   g01589(.A(new_n1782_), .B(new_n1780_), .Y(new_n1783_));
  AOI22X1  g01590(.A0(\a[32] ), .A1(\a[0] ), .B0(\a[30] ), .B1(\a[2] ), .Y(new_n1784_));
  INVX1    g01591(.A(new_n1784_), .Y(new_n1785_));
  AND2X1   g01592(.A(new_n1724_), .B(\a[16] ), .Y(new_n1786_));
  AND2X1   g01593(.A(\a[32] ), .B(\a[30] ), .Y(new_n1787_));
  AND2X1   g01594(.A(new_n1787_), .B(new_n197_), .Y(new_n1788_));
  AOI21X1  g01595(.A0(new_n1785_), .A1(new_n1786_), .B0(new_n1788_), .Y(new_n1789_));
  NAND2X1  g01596(.A(new_n1789_), .B(new_n1785_), .Y(new_n1790_));
  OAI21X1  g01597(.A0(new_n1788_), .A1(new_n1784_), .B0(new_n1786_), .Y(new_n1791_));
  AND2X1   g01598(.A(new_n1791_), .B(new_n1790_), .Y(new_n1792_));
  INVX1    g01599(.A(new_n482_), .Y(new_n1793_));
  INVX1    g01600(.A(new_n1236_), .Y(new_n1794_));
  OAI22X1  g01601(.A0(new_n1794_), .A1(new_n1793_), .B0(new_n1149_), .B1(new_n635_), .Y(new_n1795_));
  OAI21X1  g01602(.A0(new_n1521_), .A1(new_n587_), .B0(new_n1795_), .Y(new_n1796_));
  AND2X1   g01603(.A(\a[21] ), .B(\a[11] ), .Y(new_n1797_));
  AOI21X1  g01604(.A0(new_n1099_), .A1(new_n586_), .B0(new_n1795_), .Y(new_n1798_));
  OAI22X1  g01605(.A0(new_n934_), .A1(new_n453_), .B0(new_n752_), .B1(new_n591_), .Y(new_n1799_));
  AOI22X1  g01606(.A0(new_n1799_), .A1(new_n1798_), .B0(new_n1797_), .B1(new_n1796_), .Y(new_n1800_));
  XOR2X1   g01607(.A(new_n1800_), .B(new_n1792_), .Y(new_n1801_));
  AND2X1   g01608(.A(\a[18] ), .B(\a[14] ), .Y(new_n1802_));
  INVX1    g01609(.A(\a[29] ), .Y(new_n1803_));
  NOR4X1   g01610(.A(new_n1803_), .B(new_n1086_), .C(new_n570_), .D(new_n223_), .Y(new_n1804_));
  AOI22X1  g01611(.A0(\a[29] ), .A1(\a[3] ), .B0(\a[22] ), .B1(\a[10] ), .Y(new_n1805_));
  OR4X1    g01612(.A(new_n1805_), .B(new_n1804_), .C(new_n675_), .D(new_n490_), .Y(new_n1806_));
  NOR3X1   g01613(.A(new_n1805_), .B(new_n1804_), .C(new_n1802_), .Y(new_n1807_));
  AOI21X1  g01614(.A0(new_n1806_), .A1(new_n1802_), .B0(new_n1807_), .Y(new_n1808_));
  XOR2X1   g01615(.A(new_n1808_), .B(new_n1801_), .Y(new_n1809_));
  XOR2X1   g01616(.A(new_n1809_), .B(new_n1783_), .Y(new_n1810_));
  XOR2X1   g01617(.A(new_n1810_), .B(new_n1760_), .Y(new_n1811_));
  XOR2X1   g01618(.A(new_n1811_), .B(new_n1758_), .Y(new_n1812_));
  NOR2X1   g01619(.A(new_n1721_), .B(new_n1719_), .Y(new_n1813_));
  AOI21X1  g01620(.A0(new_n1727_), .A1(new_n1722_), .B0(new_n1813_), .Y(new_n1814_));
  INVX1    g01621(.A(new_n1681_), .Y(new_n1815_));
  INVX1    g01622(.A(new_n1703_), .Y(new_n1816_));
  XOR2X1   g01623(.A(new_n1693_), .B(new_n1816_), .Y(new_n1817_));
  XOR2X1   g01624(.A(new_n1817_), .B(new_n1815_), .Y(new_n1818_));
  AND2X1   g01625(.A(\a[31] ), .B(\a[1] ), .Y(new_n1819_));
  XOR2X1   g01626(.A(new_n1819_), .B(new_n753_), .Y(new_n1820_));
  INVX1    g01627(.A(new_n1820_), .Y(new_n1821_));
  XOR2X1   g01628(.A(new_n1821_), .B(new_n1667_), .Y(new_n1822_));
  INVX1    g01629(.A(new_n1822_), .Y(new_n1823_));
  XOR2X1   g01630(.A(new_n1823_), .B(new_n1657_), .Y(new_n1824_));
  INVX1    g01631(.A(new_n1824_), .Y(new_n1825_));
  XOR2X1   g01632(.A(new_n1825_), .B(new_n1818_), .Y(new_n1826_));
  XOR2X1   g01633(.A(new_n1826_), .B(new_n1814_), .Y(new_n1827_));
  INVX1    g01634(.A(new_n1687_), .Y(new_n1828_));
  AOI21X1  g01635(.A0(new_n1695_), .A1(new_n1828_), .B0(new_n1709_), .Y(new_n1829_));
  AND2X1   g01636(.A(new_n1604_), .B(new_n1732_), .Y(new_n1830_));
  AOI21X1  g01637(.A0(new_n1733_), .A1(new_n1624_), .B0(new_n1830_), .Y(new_n1831_));
  XOR2X1   g01638(.A(new_n1831_), .B(new_n1829_), .Y(new_n1832_));
  INVX1    g01639(.A(new_n1832_), .Y(new_n1833_));
  INVX1    g01640(.A(new_n1669_), .Y(new_n1834_));
  OR2X1    g01641(.A(new_n1834_), .B(new_n1660_), .Y(new_n1835_));
  OAI21X1  g01642(.A0(new_n1682_), .A1(new_n1670_), .B0(new_n1835_), .Y(new_n1836_));
  XOR2X1   g01643(.A(new_n1836_), .B(new_n1833_), .Y(new_n1837_));
  AND2X1   g01644(.A(new_n1711_), .B(new_n1683_), .Y(new_n1838_));
  AOI21X1  g01645(.A0(new_n1712_), .A1(new_n1649_), .B0(new_n1838_), .Y(new_n1839_));
  XOR2X1   g01646(.A(new_n1839_), .B(new_n1837_), .Y(new_n1840_));
  XOR2X1   g01647(.A(new_n1840_), .B(new_n1827_), .Y(new_n1841_));
  XOR2X1   g01648(.A(new_n1841_), .B(new_n1812_), .Y(new_n1842_));
  XOR2X1   g01649(.A(new_n1842_), .B(new_n1755_), .Y(new_n1843_));
  XOR2X1   g01650(.A(new_n1843_), .B(new_n1752_), .Y(\asquared[33] ));
  NOR3X1   g01651(.A(new_n1805_), .B(new_n675_), .C(new_n490_), .Y(new_n1845_));
  NOR2X1   g01652(.A(new_n1845_), .B(new_n1804_), .Y(new_n1846_));
  INVX1    g01653(.A(new_n1846_), .Y(new_n1847_));
  XOR2X1   g01654(.A(new_n1798_), .B(new_n1789_), .Y(new_n1848_));
  XOR2X1   g01655(.A(new_n1848_), .B(new_n1847_), .Y(new_n1849_));
  XOR2X1   g01656(.A(new_n1776_), .B(new_n1767_), .Y(new_n1850_));
  INVX1    g01657(.A(\a[33] ), .Y(new_n1851_));
  NOR4X1   g01658(.A(new_n1851_), .B(new_n1086_), .C(new_n488_), .D(new_n194_), .Y(new_n1852_));
  NAND4X1  g01659(.A(\a[31] ), .B(\a[22] ), .C(\a[11] ), .D(\a[2] ), .Y(new_n1853_));
  NAND4X1  g01660(.A(\a[33] ), .B(\a[31] ), .C(\a[2] ), .D(\a[0] ), .Y(new_n1854_));
  AOI21X1  g01661(.A0(new_n1854_), .A1(new_n1853_), .B0(new_n1852_), .Y(new_n1855_));
  NAND2X1  g01662(.A(\a[31] ), .B(\a[2] ), .Y(new_n1856_));
  OR2X1    g01663(.A(new_n1855_), .B(new_n1852_), .Y(new_n1857_));
  AOI22X1  g01664(.A0(\a[33] ), .A1(\a[0] ), .B0(\a[22] ), .B1(\a[11] ), .Y(new_n1858_));
  OAI22X1  g01665(.A0(new_n1858_), .A1(new_n1857_), .B0(new_n1856_), .B1(new_n1855_), .Y(new_n1859_));
  XOR2X1   g01666(.A(new_n1859_), .B(new_n1850_), .Y(new_n1860_));
  XOR2X1   g01667(.A(new_n1860_), .B(new_n1849_), .Y(new_n1861_));
  NOR4X1   g01668(.A(new_n1803_), .B(new_n1185_), .C(new_n341_), .D(new_n340_), .Y(new_n1862_));
  NAND4X1  g01669(.A(\a[30] ), .B(\a[29] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n1863_));
  NAND4X1  g01670(.A(\a[30] ), .B(\a[24] ), .C(\a[9] ), .D(\a[3] ), .Y(new_n1864_));
  AOI21X1  g01671(.A0(new_n1864_), .A1(new_n1863_), .B0(new_n1862_), .Y(new_n1865_));
  OR2X1    g01672(.A(new_n1865_), .B(new_n1862_), .Y(new_n1866_));
  AOI22X1  g01673(.A0(\a[29] ), .A1(\a[4] ), .B0(\a[24] ), .B1(\a[9] ), .Y(new_n1867_));
  NAND2X1  g01674(.A(\a[30] ), .B(\a[3] ), .Y(new_n1868_));
  OAI22X1  g01675(.A0(new_n1868_), .A1(new_n1865_), .B0(new_n1867_), .B1(new_n1866_), .Y(new_n1869_));
  NAND2X1  g01676(.A(\a[28] ), .B(\a[5] ), .Y(new_n1870_));
  AND2X1   g01677(.A(\a[27] ), .B(\a[25] ), .Y(new_n1871_));
  NAND4X1  g01678(.A(\a[28] ), .B(\a[27] ), .C(\a[6] ), .D(\a[5] ), .Y(new_n1872_));
  NAND4X1  g01679(.A(\a[28] ), .B(\a[25] ), .C(\a[8] ), .D(\a[5] ), .Y(new_n1873_));
  AOI22X1  g01680(.A0(new_n1873_), .A1(new_n1872_), .B0(new_n1871_), .B1(new_n277_), .Y(new_n1874_));
  AOI22X1  g01681(.A0(\a[27] ), .A1(\a[6] ), .B0(\a[25] ), .B1(\a[8] ), .Y(new_n1875_));
  AOI21X1  g01682(.A0(new_n1871_), .A1(new_n277_), .B0(new_n1874_), .Y(new_n1876_));
  INVX1    g01683(.A(new_n1876_), .Y(new_n1877_));
  OAI22X1  g01684(.A0(new_n1877_), .A1(new_n1875_), .B0(new_n1874_), .B1(new_n1870_), .Y(new_n1878_));
  XOR2X1   g01685(.A(new_n1878_), .B(new_n1869_), .Y(new_n1879_));
  AND2X1   g01686(.A(\a[26] ), .B(\a[7] ), .Y(new_n1880_));
  INVX1    g01687(.A(new_n1880_), .Y(new_n1881_));
  AOI22X1  g01688(.A0(\a[18] ), .A1(\a[15] ), .B0(\a[17] ), .B1(\a[16] ), .Y(new_n1882_));
  AND2X1   g01689(.A(new_n796_), .B(new_n689_), .Y(new_n1883_));
  NOR3X1   g01690(.A(new_n1882_), .B(new_n1883_), .C(new_n1881_), .Y(new_n1884_));
  NOR2X1   g01691(.A(new_n1884_), .B(new_n1883_), .Y(new_n1885_));
  INVX1    g01692(.A(new_n1885_), .Y(new_n1886_));
  OAI22X1  g01693(.A0(new_n1886_), .A1(new_n1882_), .B0(new_n1884_), .B1(new_n1881_), .Y(new_n1887_));
  XOR2X1   g01694(.A(new_n1887_), .B(new_n1879_), .Y(new_n1888_));
  INVX1    g01695(.A(new_n1888_), .Y(new_n1889_));
  XOR2X1   g01696(.A(new_n1889_), .B(new_n1861_), .Y(new_n1890_));
  AND2X1   g01697(.A(new_n1693_), .B(new_n1816_), .Y(new_n1891_));
  AOI21X1  g01698(.A0(new_n1817_), .A1(new_n1815_), .B0(new_n1891_), .Y(new_n1892_));
  INVX1    g01699(.A(new_n1892_), .Y(new_n1893_));
  OR2X1    g01700(.A(new_n1800_), .B(new_n1792_), .Y(new_n1894_));
  INVX1    g01701(.A(new_n1801_), .Y(new_n1895_));
  OAI21X1  g01702(.A0(new_n1808_), .A1(new_n1895_), .B0(new_n1894_), .Y(new_n1896_));
  XOR2X1   g01703(.A(new_n1896_), .B(new_n1893_), .Y(new_n1897_));
  INVX1    g01704(.A(new_n1769_), .Y(new_n1898_));
  NAND2X1  g01705(.A(new_n1782_), .B(new_n1780_), .Y(new_n1899_));
  OAI21X1  g01706(.A0(new_n1778_), .A1(new_n1898_), .B0(new_n1899_), .Y(new_n1900_));
  XOR2X1   g01707(.A(new_n1900_), .B(new_n1897_), .Y(new_n1901_));
  XOR2X1   g01708(.A(new_n1808_), .B(new_n1895_), .Y(new_n1902_));
  AND2X1   g01709(.A(new_n1902_), .B(new_n1783_), .Y(new_n1903_));
  INVX1    g01710(.A(new_n1903_), .Y(new_n1904_));
  OAI21X1  g01711(.A0(new_n1810_), .A1(new_n1760_), .B0(new_n1904_), .Y(new_n1905_));
  INVX1    g01712(.A(new_n1905_), .Y(new_n1906_));
  XOR2X1   g01713(.A(new_n1906_), .B(new_n1901_), .Y(new_n1907_));
  XOR2X1   g01714(.A(new_n1907_), .B(new_n1890_), .Y(new_n1908_));
  AOI22X1  g01715(.A0(new_n1819_), .A1(new_n753_), .B0(\a[23] ), .B1(\a[10] ), .Y(new_n1909_));
  INVX1    g01716(.A(new_n1909_), .Y(new_n1910_));
  NAND4X1  g01717(.A(new_n1819_), .B(new_n753_), .C(\a[23] ), .D(\a[10] ), .Y(new_n1911_));
  INVX1    g01718(.A(new_n1911_), .Y(new_n1912_));
  AND2X1   g01719(.A(\a[32] ), .B(\a[1] ), .Y(new_n1913_));
  XOR2X1   g01720(.A(new_n1913_), .B(new_n616_), .Y(new_n1914_));
  INVX1    g01721(.A(new_n1914_), .Y(new_n1915_));
  AOI21X1  g01722(.A0(new_n1915_), .A1(new_n1910_), .B0(new_n1912_), .Y(new_n1916_));
  AOI21X1  g01723(.A0(new_n1911_), .A1(new_n1910_), .B0(new_n1914_), .Y(new_n1917_));
  AOI21X1  g01724(.A0(new_n1916_), .A1(new_n1910_), .B0(new_n1917_), .Y(new_n1918_));
  OAI22X1  g01725(.A0(new_n1794_), .A1(new_n587_), .B0(new_n1149_), .B1(new_n585_), .Y(new_n1919_));
  OAI21X1  g01726(.A0(new_n1521_), .A1(new_n583_), .B0(new_n1919_), .Y(new_n1920_));
  AND2X1   g01727(.A(\a[21] ), .B(\a[12] ), .Y(new_n1921_));
  AOI21X1  g01728(.A0(new_n1099_), .A1(new_n582_), .B0(new_n1919_), .Y(new_n1922_));
  OAI22X1  g01729(.A0(new_n934_), .A1(new_n591_), .B0(new_n752_), .B1(new_n490_), .Y(new_n1923_));
  AOI22X1  g01730(.A0(new_n1923_), .A1(new_n1922_), .B0(new_n1921_), .B1(new_n1920_), .Y(new_n1924_));
  XOR2X1   g01731(.A(new_n1924_), .B(new_n1918_), .Y(new_n1925_));
  OR2X1    g01732(.A(new_n1821_), .B(new_n1667_), .Y(new_n1926_));
  OAI21X1  g01733(.A0(new_n1823_), .A1(new_n1657_), .B0(new_n1926_), .Y(new_n1927_));
  XOR2X1   g01734(.A(new_n1927_), .B(new_n1925_), .Y(new_n1928_));
  NOR2X1   g01735(.A(new_n1831_), .B(new_n1829_), .Y(new_n1929_));
  AOI21X1  g01736(.A0(new_n1836_), .A1(new_n1832_), .B0(new_n1929_), .Y(new_n1930_));
  XOR2X1   g01737(.A(new_n1930_), .B(new_n1928_), .Y(new_n1931_));
  NOR2X1   g01738(.A(new_n1826_), .B(new_n1814_), .Y(new_n1932_));
  AOI21X1  g01739(.A0(new_n1824_), .A1(new_n1818_), .B0(new_n1932_), .Y(new_n1933_));
  XOR2X1   g01740(.A(new_n1933_), .B(new_n1931_), .Y(new_n1934_));
  NAND2X1  g01741(.A(new_n1840_), .B(new_n1827_), .Y(new_n1935_));
  OAI21X1  g01742(.A0(new_n1839_), .A1(new_n1837_), .B0(new_n1935_), .Y(new_n1936_));
  XOR2X1   g01743(.A(new_n1936_), .B(new_n1934_), .Y(new_n1937_));
  XOR2X1   g01744(.A(new_n1937_), .B(new_n1908_), .Y(new_n1938_));
  AND2X1   g01745(.A(new_n1811_), .B(new_n1758_), .Y(new_n1939_));
  AOI21X1  g01746(.A0(new_n1841_), .A1(new_n1812_), .B0(new_n1939_), .Y(new_n1940_));
  XOR2X1   g01747(.A(new_n1940_), .B(new_n1938_), .Y(new_n1941_));
  AND2X1   g01748(.A(new_n1842_), .B(new_n1755_), .Y(new_n1942_));
  OR2X1    g01749(.A(new_n1842_), .B(new_n1755_), .Y(new_n1943_));
  AOI21X1  g01750(.A0(new_n1943_), .A1(new_n1752_), .B0(new_n1942_), .Y(new_n1944_));
  XOR2X1   g01751(.A(new_n1944_), .B(new_n1941_), .Y(\asquared[34] ));
  AND2X1   g01752(.A(new_n1936_), .B(new_n1934_), .Y(new_n1946_));
  AND2X1   g01753(.A(new_n1937_), .B(new_n1908_), .Y(new_n1947_));
  OR2X1    g01754(.A(new_n1947_), .B(new_n1946_), .Y(new_n1948_));
  XOR2X1   g01755(.A(new_n1866_), .B(new_n1857_), .Y(new_n1949_));
  XOR2X1   g01756(.A(new_n1949_), .B(new_n1876_), .Y(new_n1950_));
  AND2X1   g01757(.A(new_n1878_), .B(new_n1869_), .Y(new_n1951_));
  AOI21X1  g01758(.A0(new_n1887_), .A1(new_n1879_), .B0(new_n1951_), .Y(new_n1952_));
  AND2X1   g01759(.A(new_n1913_), .B(\a[17] ), .Y(new_n1953_));
  AND2X1   g01760(.A(\a[33] ), .B(\a[1] ), .Y(new_n1954_));
  XOR2X1   g01761(.A(new_n1954_), .B(new_n794_), .Y(new_n1955_));
  XOR2X1   g01762(.A(new_n1955_), .B(new_n1953_), .Y(new_n1956_));
  XOR2X1   g01763(.A(new_n1956_), .B(new_n1886_), .Y(new_n1957_));
  INVX1    g01764(.A(new_n1957_), .Y(new_n1958_));
  XOR2X1   g01765(.A(new_n1958_), .B(new_n1952_), .Y(new_n1959_));
  INVX1    g01766(.A(new_n1959_), .Y(new_n1960_));
  XOR2X1   g01767(.A(new_n1960_), .B(new_n1950_), .Y(new_n1961_));
  XOR2X1   g01768(.A(new_n1922_), .B(new_n1916_), .Y(new_n1962_));
  AND2X1   g01769(.A(\a[32] ), .B(\a[2] ), .Y(new_n1963_));
  INVX1    g01770(.A(new_n1963_), .Y(new_n1964_));
  AOI22X1  g01771(.A0(\a[23] ), .A1(\a[11] ), .B0(\a[22] ), .B1(\a[12] ), .Y(new_n1965_));
  AND2X1   g01772(.A(new_n1394_), .B(new_n482_), .Y(new_n1966_));
  NOR3X1   g01773(.A(new_n1965_), .B(new_n1966_), .C(new_n1964_), .Y(new_n1967_));
  NOR2X1   g01774(.A(new_n1967_), .B(new_n1966_), .Y(new_n1968_));
  INVX1    g01775(.A(new_n1968_), .Y(new_n1969_));
  OAI22X1  g01776(.A0(new_n1969_), .A1(new_n1965_), .B0(new_n1967_), .B1(new_n1964_), .Y(new_n1970_));
  XOR2X1   g01777(.A(new_n1970_), .B(new_n1962_), .Y(new_n1971_));
  INVX1    g01778(.A(new_n1971_), .Y(new_n1972_));
  NAND2X1  g01779(.A(new_n1927_), .B(new_n1925_), .Y(new_n1973_));
  OAI21X1  g01780(.A0(new_n1924_), .A1(new_n1918_), .B0(new_n1973_), .Y(new_n1974_));
  XOR2X1   g01781(.A(new_n1974_), .B(new_n1972_), .Y(new_n1975_));
  NOR4X1   g01782(.A(new_n1803_), .B(new_n1326_), .C(new_n341_), .D(new_n255_), .Y(new_n1976_));
  NAND4X1  g01783(.A(\a[29] ), .B(\a[24] ), .C(\a[10] ), .D(\a[5] ), .Y(new_n1977_));
  NAND4X1  g01784(.A(\a[25] ), .B(\a[24] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n1978_));
  AOI21X1  g01785(.A0(new_n1978_), .A1(new_n1977_), .B0(new_n1976_), .Y(new_n1979_));
  NAND2X1  g01786(.A(new_n1978_), .B(new_n1977_), .Y(new_n1980_));
  NOR2X1   g01787(.A(new_n1980_), .B(new_n1976_), .Y(new_n1981_));
  INVX1    g01788(.A(new_n1981_), .Y(new_n1982_));
  AOI22X1  g01789(.A0(\a[29] ), .A1(\a[5] ), .B0(\a[25] ), .B1(\a[9] ), .Y(new_n1983_));
  NAND2X1  g01790(.A(\a[24] ), .B(\a[10] ), .Y(new_n1984_));
  OAI22X1  g01791(.A0(new_n1984_), .A1(new_n1979_), .B0(new_n1983_), .B1(new_n1982_), .Y(new_n1985_));
  NAND4X1  g01792(.A(\a[21] ), .B(\a[19] ), .C(\a[15] ), .D(\a[13] ), .Y(new_n1986_));
  NAND4X1  g01793(.A(\a[21] ), .B(\a[20] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n1987_));
  AOI22X1  g01794(.A0(new_n1987_), .A1(new_n1986_), .B0(new_n1099_), .B1(new_n691_), .Y(new_n1988_));
  NAND2X1  g01795(.A(\a[21] ), .B(\a[13] ), .Y(new_n1989_));
  NAND4X1  g01796(.A(\a[20] ), .B(\a[19] ), .C(\a[15] ), .D(\a[14] ), .Y(new_n1990_));
  NAND3X1  g01797(.A(new_n1987_), .B(new_n1986_), .C(new_n1990_), .Y(new_n1991_));
  AOI22X1  g01798(.A0(\a[20] ), .A1(\a[14] ), .B0(\a[19] ), .B1(\a[15] ), .Y(new_n1992_));
  OAI22X1  g01799(.A0(new_n1992_), .A1(new_n1991_), .B0(new_n1989_), .B1(new_n1988_), .Y(new_n1993_));
  XOR2X1   g01800(.A(new_n1993_), .B(new_n1985_), .Y(new_n1994_));
  AND2X1   g01801(.A(\a[27] ), .B(\a[26] ), .Y(new_n1995_));
  AND2X1   g01802(.A(\a[28] ), .B(\a[26] ), .Y(new_n1996_));
  AOI22X1  g01803(.A0(new_n1996_), .A1(new_n277_), .B0(new_n1671_), .B1(new_n375_), .Y(new_n1997_));
  AOI21X1  g01804(.A0(new_n1995_), .A1(new_n325_), .B0(new_n1997_), .Y(new_n1998_));
  AND2X1   g01805(.A(\a[28] ), .B(\a[6] ), .Y(new_n1999_));
  INVX1    g01806(.A(new_n1999_), .Y(new_n2000_));
  AOI21X1  g01807(.A0(new_n1995_), .A1(new_n325_), .B0(new_n1998_), .Y(new_n2001_));
  INVX1    g01808(.A(new_n2001_), .Y(new_n2002_));
  AOI22X1  g01809(.A0(\a[27] ), .A1(\a[7] ), .B0(\a[26] ), .B1(\a[8] ), .Y(new_n2003_));
  OAI22X1  g01810(.A0(new_n2003_), .A1(new_n2002_), .B0(new_n2000_), .B1(new_n1998_), .Y(new_n2004_));
  INVX1    g01811(.A(new_n2004_), .Y(new_n2005_));
  XOR2X1   g01812(.A(new_n2005_), .B(new_n1994_), .Y(new_n2006_));
  AND2X1   g01813(.A(new_n2006_), .B(new_n1975_), .Y(new_n2007_));
  OAI21X1  g01814(.A0(new_n2006_), .A1(new_n1975_), .B0(new_n1961_), .Y(new_n2008_));
  XOR2X1   g01815(.A(new_n2006_), .B(new_n1975_), .Y(new_n2009_));
  OAI22X1  g01816(.A0(new_n2009_), .A1(new_n1961_), .B0(new_n2008_), .B1(new_n2007_), .Y(new_n2010_));
  INVX1    g01817(.A(new_n1928_), .Y(new_n2011_));
  OR2X1    g01818(.A(new_n1930_), .B(new_n2011_), .Y(new_n2012_));
  OAI21X1  g01819(.A0(new_n1933_), .A1(new_n1931_), .B0(new_n2012_), .Y(new_n2013_));
  XOR2X1   g01820(.A(new_n2013_), .B(new_n2010_), .Y(new_n2014_));
  AND2X1   g01821(.A(new_n1905_), .B(new_n1901_), .Y(new_n2015_));
  NOR2X1   g01822(.A(new_n1907_), .B(new_n1890_), .Y(new_n2016_));
  NOR2X1   g01823(.A(new_n2016_), .B(new_n2015_), .Y(new_n2017_));
  AND2X1   g01824(.A(new_n1860_), .B(new_n1849_), .Y(new_n2018_));
  AOI21X1  g01825(.A0(new_n1888_), .A1(new_n1861_), .B0(new_n2018_), .Y(new_n2019_));
  AND2X1   g01826(.A(new_n1896_), .B(new_n1893_), .Y(new_n2020_));
  AOI21X1  g01827(.A0(new_n1900_), .A1(new_n1897_), .B0(new_n2020_), .Y(new_n2021_));
  XOR2X1   g01828(.A(new_n2021_), .B(new_n2019_), .Y(new_n2022_));
  NAND2X1  g01829(.A(new_n1859_), .B(new_n1850_), .Y(new_n2023_));
  OAI21X1  g01830(.A0(new_n1776_), .A1(new_n1767_), .B0(new_n2023_), .Y(new_n2024_));
  NOR2X1   g01831(.A(new_n1798_), .B(new_n1789_), .Y(new_n2025_));
  AOI21X1  g01832(.A0(new_n1848_), .A1(new_n1847_), .B0(new_n2025_), .Y(new_n2026_));
  AOI22X1  g01833(.A0(new_n210_), .A1(\a[30] ), .B0(new_n204_), .B1(\a[31] ), .Y(new_n2027_));
  INVX1    g01834(.A(\a[34] ), .Y(new_n2028_));
  NOR3X1   g01835(.A(new_n217_), .B(new_n1704_), .C(new_n1684_), .Y(new_n2029_));
  OR2X1    g01836(.A(new_n2029_), .B(new_n2028_), .Y(new_n2030_));
  AOI22X1  g01837(.A0(\a[31] ), .A1(\a[3] ), .B0(\a[30] ), .B1(\a[4] ), .Y(new_n2031_));
  OAI22X1  g01838(.A0(new_n2031_), .A1(new_n2029_), .B0(new_n2028_), .B1(new_n194_), .Y(new_n2032_));
  OAI21X1  g01839(.A0(new_n2030_), .A1(new_n2027_), .B0(new_n2032_), .Y(new_n2033_));
  XOR2X1   g01840(.A(new_n2033_), .B(new_n2026_), .Y(new_n2034_));
  XOR2X1   g01841(.A(new_n2034_), .B(new_n2024_), .Y(new_n2035_));
  XOR2X1   g01842(.A(new_n2035_), .B(new_n2022_), .Y(new_n2036_));
  XOR2X1   g01843(.A(new_n2036_), .B(new_n2017_), .Y(new_n2037_));
  XOR2X1   g01844(.A(new_n2037_), .B(new_n2014_), .Y(new_n2038_));
  AND2X1   g01845(.A(new_n2038_), .B(new_n1948_), .Y(new_n2039_));
  INVX1    g01846(.A(new_n2039_), .Y(new_n2040_));
  INVX1    g01847(.A(new_n1938_), .Y(new_n2041_));
  AND2X1   g01848(.A(new_n1940_), .B(new_n2041_), .Y(new_n2042_));
  OR2X1    g01849(.A(new_n1940_), .B(new_n2041_), .Y(new_n2043_));
  OAI21X1  g01850(.A0(new_n1944_), .A1(new_n2042_), .B0(new_n2043_), .Y(new_n2044_));
  NOR2X1   g01851(.A(new_n2038_), .B(new_n1948_), .Y(new_n2045_));
  INVX1    g01852(.A(new_n2045_), .Y(new_n2046_));
  AOI21X1  g01853(.A0(new_n2046_), .A1(new_n2040_), .B0(new_n2044_), .Y(new_n2047_));
  AND2X1   g01854(.A(new_n2046_), .B(new_n2044_), .Y(new_n2048_));
  AOI21X1  g01855(.A0(new_n2048_), .A1(new_n2040_), .B0(new_n2047_), .Y(\asquared[35] ));
  AOI21X1  g01856(.A0(new_n2046_), .A1(new_n2044_), .B0(new_n2039_), .Y(new_n2050_));
  OAI21X1  g01857(.A0(new_n2016_), .A1(new_n2015_), .B0(new_n2036_), .Y(new_n2051_));
  OAI21X1  g01858(.A0(new_n2037_), .A1(new_n2014_), .B0(new_n2051_), .Y(new_n2052_));
  NOR2X1   g01859(.A(new_n2008_), .B(new_n2007_), .Y(new_n2053_));
  INVX1    g01860(.A(new_n2010_), .Y(new_n2054_));
  AOI21X1  g01861(.A0(new_n2013_), .A1(new_n2054_), .B0(new_n2053_), .Y(new_n2055_));
  AND2X1   g01862(.A(new_n1866_), .B(new_n1857_), .Y(new_n2056_));
  AOI21X1  g01863(.A0(new_n1949_), .A1(new_n1877_), .B0(new_n2056_), .Y(new_n2057_));
  AND2X1   g01864(.A(new_n1955_), .B(new_n1953_), .Y(new_n2058_));
  AOI21X1  g01865(.A0(new_n1956_), .A1(new_n1886_), .B0(new_n2058_), .Y(new_n2059_));
  XOR2X1   g01866(.A(new_n2059_), .B(new_n2057_), .Y(new_n2060_));
  INVX1    g01867(.A(new_n2060_), .Y(new_n2061_));
  NOR2X1   g01868(.A(new_n1922_), .B(new_n1916_), .Y(new_n2062_));
  AOI21X1  g01869(.A0(new_n1970_), .A1(new_n1962_), .B0(new_n2062_), .Y(new_n2063_));
  XOR2X1   g01870(.A(new_n2063_), .B(new_n2061_), .Y(new_n2064_));
  OR2X1    g01871(.A(new_n1958_), .B(new_n1952_), .Y(new_n2065_));
  OAI21X1  g01872(.A0(new_n1960_), .A1(new_n1950_), .B0(new_n2065_), .Y(new_n2066_));
  XOR2X1   g01873(.A(new_n2066_), .B(new_n2064_), .Y(new_n2067_));
  NAND2X1  g01874(.A(new_n1974_), .B(new_n1971_), .Y(new_n2068_));
  OAI21X1  g01875(.A0(new_n2006_), .A1(new_n1975_), .B0(new_n2068_), .Y(new_n2069_));
  XOR2X1   g01876(.A(new_n2069_), .B(new_n2067_), .Y(new_n2070_));
  XOR2X1   g01877(.A(new_n2070_), .B(new_n2055_), .Y(new_n2071_));
  NOR2X1   g01878(.A(new_n2021_), .B(new_n2019_), .Y(new_n2072_));
  AOI21X1  g01879(.A0(new_n2035_), .A1(new_n2022_), .B0(new_n2072_), .Y(new_n2073_));
  XOR2X1   g01880(.A(new_n1991_), .B(new_n1969_), .Y(new_n2074_));
  AND2X1   g01881(.A(\a[31] ), .B(\a[30] ), .Y(new_n2075_));
  INVX1    g01882(.A(new_n2075_), .Y(new_n2076_));
  OAI22X1  g01883(.A0(new_n2076_), .A1(new_n217_), .B0(new_n2027_), .B1(new_n2028_), .Y(new_n2077_));
  XOR2X1   g01884(.A(new_n2077_), .B(new_n2074_), .Y(new_n2078_));
  AND2X1   g01885(.A(new_n1993_), .B(new_n1985_), .Y(new_n2079_));
  AOI21X1  g01886(.A0(new_n2004_), .A1(new_n1994_), .B0(new_n2079_), .Y(new_n2080_));
  AOI21X1  g01887(.A0(\a[34] ), .A1(\a[1] ), .B0(\a[18] ), .Y(new_n2081_));
  AOI21X1  g01888(.A0(new_n745_), .A1(\a[34] ), .B0(new_n2081_), .Y(new_n2082_));
  XOR2X1   g01889(.A(new_n2082_), .B(new_n2002_), .Y(new_n2083_));
  XOR2X1   g01890(.A(new_n2083_), .B(new_n1981_), .Y(new_n2084_));
  XOR2X1   g01891(.A(new_n2084_), .B(new_n2080_), .Y(new_n2085_));
  XOR2X1   g01892(.A(new_n2085_), .B(new_n2078_), .Y(new_n2086_));
  INVX1    g01893(.A(new_n2086_), .Y(new_n2087_));
  XOR2X1   g01894(.A(new_n2087_), .B(new_n2073_), .Y(new_n2088_));
  INVX1    g01895(.A(new_n2088_), .Y(new_n2089_));
  NAND4X1  g01896(.A(\a[30] ), .B(\a[27] ), .C(\a[8] ), .D(\a[5] ), .Y(new_n2090_));
  NAND4X1  g01897(.A(\a[30] ), .B(\a[29] ), .C(\a[6] ), .D(\a[5] ), .Y(new_n2091_));
  AOI22X1  g01898(.A0(new_n2091_), .A1(new_n2090_), .B0(new_n1484_), .B1(new_n277_), .Y(new_n2092_));
  AOI21X1  g01899(.A0(new_n1484_), .A1(new_n277_), .B0(new_n2092_), .Y(new_n2093_));
  OAI22X1  g01900(.A0(new_n1803_), .A1(new_n230_), .B0(new_n1679_), .B1(new_n413_), .Y(new_n2094_));
  NOR3X1   g01901(.A(new_n2092_), .B(new_n1684_), .C(new_n255_), .Y(new_n2095_));
  AOI21X1  g01902(.A0(new_n2094_), .A1(new_n2093_), .B0(new_n2095_), .Y(new_n2096_));
  AND2X1   g01903(.A(\a[28] ), .B(\a[7] ), .Y(new_n2097_));
  INVX1    g01904(.A(new_n2097_), .Y(new_n2098_));
  AOI22X1  g01905(.A0(\a[19] ), .A1(\a[16] ), .B0(\a[18] ), .B1(\a[17] ), .Y(new_n2099_));
  NOR4X1   g01906(.A(new_n752_), .B(new_n675_), .C(new_n616_), .D(new_n571_), .Y(new_n2100_));
  NOR3X1   g01907(.A(new_n2099_), .B(new_n2100_), .C(new_n2098_), .Y(new_n2101_));
  NOR2X1   g01908(.A(new_n2101_), .B(new_n2100_), .Y(new_n2102_));
  INVX1    g01909(.A(new_n2102_), .Y(new_n2103_));
  OAI22X1  g01910(.A0(new_n2103_), .A1(new_n2099_), .B0(new_n2101_), .B1(new_n2098_), .Y(new_n2104_));
  XOR2X1   g01911(.A(new_n2104_), .B(new_n2096_), .Y(new_n2105_));
  AND2X1   g01912(.A(\a[31] ), .B(\a[4] ), .Y(new_n2106_));
  AOI22X1  g01913(.A0(\a[26] ), .A1(\a[9] ), .B0(\a[25] ), .B1(\a[10] ), .Y(new_n2107_));
  INVX1    g01914(.A(new_n2107_), .Y(new_n2108_));
  NAND4X1  g01915(.A(\a[26] ), .B(\a[25] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n2109_));
  NAND3X1  g01916(.A(new_n2108_), .B(new_n2109_), .C(new_n2106_), .Y(new_n2110_));
  AOI22X1  g01917(.A0(new_n2108_), .A1(new_n2106_), .B0(new_n1770_), .B1(new_n881_), .Y(new_n2111_));
  AOI22X1  g01918(.A0(new_n2111_), .A1(new_n2108_), .B0(new_n2110_), .B1(new_n2106_), .Y(new_n2112_));
  XOR2X1   g01919(.A(new_n2112_), .B(new_n2105_), .Y(new_n2113_));
  NOR2X1   g01920(.A(new_n2033_), .B(new_n2026_), .Y(new_n2114_));
  AOI21X1  g01921(.A0(new_n2034_), .A1(new_n2024_), .B0(new_n2114_), .Y(new_n2115_));
  XOR2X1   g01922(.A(new_n2115_), .B(new_n2113_), .Y(new_n2116_));
  AOI22X1  g01923(.A0(\a[35] ), .A1(\a[0] ), .B0(\a[33] ), .B1(\a[2] ), .Y(new_n2117_));
  INVX1    g01924(.A(new_n2117_), .Y(new_n2118_));
  AND2X1   g01925(.A(new_n1954_), .B(new_n794_), .Y(new_n2119_));
  AND2X1   g01926(.A(\a[35] ), .B(\a[33] ), .Y(new_n2120_));
  AND2X1   g01927(.A(new_n2120_), .B(new_n197_), .Y(new_n2121_));
  AOI21X1  g01928(.A0(new_n2118_), .A1(new_n2119_), .B0(new_n2121_), .Y(new_n2122_));
  NAND2X1  g01929(.A(new_n2122_), .B(new_n2118_), .Y(new_n2123_));
  OAI21X1  g01930(.A0(new_n2121_), .A1(new_n2117_), .B0(new_n2119_), .Y(new_n2124_));
  AND2X1   g01931(.A(new_n2124_), .B(new_n2123_), .Y(new_n2125_));
  AND2X1   g01932(.A(\a[32] ), .B(\a[3] ), .Y(new_n2126_));
  AOI22X1  g01933(.A0(\a[24] ), .A1(\a[11] ), .B0(\a[23] ), .B1(\a[12] ), .Y(new_n2127_));
  INVX1    g01934(.A(new_n2127_), .Y(new_n2128_));
  NAND4X1  g01935(.A(\a[24] ), .B(\a[23] ), .C(\a[12] ), .D(\a[11] ), .Y(new_n2129_));
  NAND3X1  g01936(.A(new_n2128_), .B(new_n2129_), .C(new_n2126_), .Y(new_n2130_));
  AOI22X1  g01937(.A0(new_n2128_), .A1(new_n2126_), .B0(new_n1219_), .B1(new_n482_), .Y(new_n2131_));
  AOI22X1  g01938(.A0(new_n2131_), .A1(new_n2128_), .B0(new_n2130_), .B1(new_n2126_), .Y(new_n2132_));
  XOR2X1   g01939(.A(new_n2132_), .B(new_n2125_), .Y(new_n2133_));
  AND2X1   g01940(.A(\a[22] ), .B(\a[20] ), .Y(new_n2134_));
  INVX1    g01941(.A(new_n2134_), .Y(new_n2135_));
  OAI22X1  g01942(.A0(new_n2135_), .A1(new_n866_), .B0(new_n1397_), .B1(new_n583_), .Y(new_n2136_));
  OAI21X1  g01943(.A0(new_n1794_), .A1(new_n867_), .B0(new_n2136_), .Y(new_n2137_));
  AND2X1   g01944(.A(\a[22] ), .B(\a[13] ), .Y(new_n2138_));
  AOI21X1  g01945(.A0(new_n1236_), .A1(new_n691_), .B0(new_n2136_), .Y(new_n2139_));
  OAI22X1  g01946(.A0(new_n1098_), .A1(new_n490_), .B0(new_n934_), .B1(new_n549_), .Y(new_n2140_));
  AOI22X1  g01947(.A0(new_n2140_), .A1(new_n2139_), .B0(new_n2138_), .B1(new_n2137_), .Y(new_n2141_));
  XOR2X1   g01948(.A(new_n2141_), .B(new_n2133_), .Y(new_n2142_));
  XOR2X1   g01949(.A(new_n2142_), .B(new_n2116_), .Y(new_n2143_));
  XOR2X1   g01950(.A(new_n2143_), .B(new_n2089_), .Y(new_n2144_));
  XOR2X1   g01951(.A(new_n2144_), .B(new_n2071_), .Y(new_n2145_));
  NOR2X1   g01952(.A(new_n2145_), .B(new_n2052_), .Y(new_n2146_));
  AND2X1   g01953(.A(new_n2145_), .B(new_n2052_), .Y(new_n2147_));
  OR2X1    g01954(.A(new_n2147_), .B(new_n2146_), .Y(new_n2148_));
  XOR2X1   g01955(.A(new_n2148_), .B(new_n2050_), .Y(\asquared[36] ));
  INVX1    g01956(.A(new_n2070_), .Y(new_n2150_));
  NOR2X1   g01957(.A(new_n2150_), .B(new_n2055_), .Y(new_n2151_));
  NOR2X1   g01958(.A(new_n2144_), .B(new_n2071_), .Y(new_n2152_));
  NOR2X1   g01959(.A(new_n2152_), .B(new_n2151_), .Y(new_n2153_));
  INVX1    g01960(.A(new_n2153_), .Y(new_n2154_));
  NOR2X1   g01961(.A(new_n2087_), .B(new_n2073_), .Y(new_n2155_));
  AOI21X1  g01962(.A0(new_n2143_), .A1(new_n2088_), .B0(new_n2155_), .Y(new_n2156_));
  AND2X1   g01963(.A(new_n1991_), .B(new_n1969_), .Y(new_n2157_));
  AOI21X1  g01964(.A0(new_n2077_), .A1(new_n2074_), .B0(new_n2157_), .Y(new_n2158_));
  AND2X1   g01965(.A(new_n2082_), .B(new_n2002_), .Y(new_n2159_));
  AOI21X1  g01966(.A0(new_n2083_), .A1(new_n1982_), .B0(new_n2159_), .Y(new_n2160_));
  XOR2X1   g01967(.A(new_n2160_), .B(new_n2158_), .Y(new_n2161_));
  INVX1    g01968(.A(new_n2161_), .Y(new_n2162_));
  OR2X1    g01969(.A(new_n2132_), .B(new_n2125_), .Y(new_n2163_));
  INVX1    g01970(.A(new_n2133_), .Y(new_n2164_));
  OAI21X1  g01971(.A0(new_n2141_), .A1(new_n2164_), .B0(new_n2163_), .Y(new_n2165_));
  XOR2X1   g01972(.A(new_n2165_), .B(new_n2162_), .Y(new_n2166_));
  NOR2X1   g01973(.A(new_n2084_), .B(new_n2080_), .Y(new_n2167_));
  AOI21X1  g01974(.A0(new_n2085_), .A1(new_n2078_), .B0(new_n2167_), .Y(new_n2168_));
  XOR2X1   g01975(.A(new_n2168_), .B(new_n2166_), .Y(new_n2169_));
  INVX1    g01976(.A(new_n2169_), .Y(new_n2170_));
  AND2X1   g01977(.A(new_n2034_), .B(new_n2024_), .Y(new_n2171_));
  OAI21X1  g01978(.A0(new_n2171_), .A1(new_n2114_), .B0(new_n2113_), .Y(new_n2172_));
  OR2X1    g01979(.A(new_n2142_), .B(new_n2116_), .Y(new_n2173_));
  AND2X1   g01980(.A(new_n2173_), .B(new_n2172_), .Y(new_n2174_));
  XOR2X1   g01981(.A(new_n2174_), .B(new_n2170_), .Y(new_n2175_));
  XOR2X1   g01982(.A(new_n2175_), .B(new_n2156_), .Y(new_n2176_));
  AOI22X1  g01983(.A0(\a[24] ), .A1(\a[12] ), .B0(\a[23] ), .B1(\a[13] ), .Y(new_n2177_));
  AND2X1   g01984(.A(\a[34] ), .B(\a[2] ), .Y(new_n2178_));
  INVX1    g01985(.A(new_n2178_), .Y(new_n2179_));
  AND2X1   g01986(.A(new_n1219_), .B(new_n586_), .Y(new_n2180_));
  NOR3X1   g01987(.A(new_n2179_), .B(new_n2180_), .C(new_n2177_), .Y(new_n2181_));
  INVX1    g01988(.A(new_n2177_), .Y(new_n2182_));
  AOI21X1  g01989(.A0(new_n2178_), .A1(new_n2182_), .B0(new_n2180_), .Y(new_n2183_));
  INVX1    g01990(.A(new_n2183_), .Y(new_n2184_));
  OAI22X1  g01991(.A0(new_n2184_), .A1(new_n2177_), .B0(new_n2181_), .B1(new_n2179_), .Y(new_n2185_));
  NOR4X1   g01992(.A(new_n1704_), .B(new_n1679_), .C(new_n341_), .D(new_n255_), .Y(new_n2186_));
  AND2X1   g01993(.A(\a[26] ), .B(\a[5] ), .Y(new_n2187_));
  AOI22X1  g01994(.A0(new_n1699_), .A1(new_n2187_), .B0(new_n1995_), .B1(new_n881_), .Y(new_n2188_));
  OR2X1    g01995(.A(new_n2188_), .B(new_n2186_), .Y(new_n2189_));
  AND2X1   g01996(.A(\a[26] ), .B(\a[10] ), .Y(new_n2190_));
  INVX1    g01997(.A(new_n2186_), .Y(new_n2191_));
  AND2X1   g01998(.A(new_n2188_), .B(new_n2191_), .Y(new_n2192_));
  OAI22X1  g01999(.A0(new_n1704_), .A1(new_n255_), .B0(new_n1679_), .B1(new_n341_), .Y(new_n2193_));
  AOI22X1  g02000(.A0(new_n2193_), .A1(new_n2192_), .B0(new_n2190_), .B1(new_n2189_), .Y(new_n2194_));
  XOR2X1   g02001(.A(new_n2194_), .B(new_n2185_), .Y(new_n2195_));
  AND2X1   g02002(.A(\a[30] ), .B(\a[29] ), .Y(new_n2196_));
  INVX1    g02003(.A(new_n2196_), .Y(new_n2197_));
  AND2X1   g02004(.A(\a[30] ), .B(\a[28] ), .Y(new_n2198_));
  INVX1    g02005(.A(new_n2198_), .Y(new_n2199_));
  OAI22X1  g02006(.A0(new_n2199_), .A1(new_n280_), .B0(new_n2197_), .B1(new_n376_), .Y(new_n2200_));
  OAI21X1  g02007(.A0(new_n1675_), .A1(new_n445_), .B0(new_n2200_), .Y(new_n2201_));
  AND2X1   g02008(.A(\a[30] ), .B(\a[6] ), .Y(new_n2202_));
  AOI21X1  g02009(.A0(new_n1674_), .A1(new_n325_), .B0(new_n2200_), .Y(new_n2203_));
  OAI22X1  g02010(.A0(new_n1803_), .A1(new_n532_), .B0(new_n1431_), .B1(new_n413_), .Y(new_n2204_));
  AOI22X1  g02011(.A0(new_n2204_), .A1(new_n2203_), .B0(new_n2202_), .B1(new_n2201_), .Y(new_n2205_));
  XOR2X1   g02012(.A(new_n2205_), .B(new_n2195_), .Y(new_n2206_));
  OR2X1    g02013(.A(new_n2059_), .B(new_n2057_), .Y(new_n2207_));
  OAI21X1  g02014(.A0(new_n2063_), .A1(new_n2061_), .B0(new_n2207_), .Y(new_n2208_));
  NAND3X1  g02015(.A(\a[34] ), .B(\a[18] ), .C(\a[1] ), .Y(new_n2209_));
  NAND2X1  g02016(.A(\a[36] ), .B(\a[0] ), .Y(new_n2210_));
  XOR2X1   g02017(.A(new_n2210_), .B(new_n2209_), .Y(new_n2211_));
  AND2X1   g02018(.A(\a[35] ), .B(\a[1] ), .Y(new_n2212_));
  AND2X1   g02019(.A(\a[19] ), .B(\a[17] ), .Y(new_n2213_));
  INVX1    g02020(.A(new_n2213_), .Y(new_n2214_));
  XOR2X1   g02021(.A(new_n2214_), .B(new_n2212_), .Y(new_n2215_));
  XOR2X1   g02022(.A(new_n2215_), .B(new_n2211_), .Y(new_n2216_));
  AND2X1   g02023(.A(\a[33] ), .B(\a[3] ), .Y(new_n2217_));
  INVX1    g02024(.A(new_n2217_), .Y(new_n2218_));
  INVX1    g02025(.A(\a[32] ), .Y(new_n2219_));
  NOR4X1   g02026(.A(new_n2219_), .B(new_n1326_), .C(new_n488_), .D(new_n340_), .Y(new_n2220_));
  NAND4X1  g02027(.A(\a[33] ), .B(\a[32] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n2221_));
  NAND4X1  g02028(.A(\a[33] ), .B(\a[25] ), .C(\a[11] ), .D(\a[3] ), .Y(new_n2222_));
  AOI21X1  g02029(.A0(new_n2222_), .A1(new_n2221_), .B0(new_n2220_), .Y(new_n2223_));
  OR2X1    g02030(.A(new_n2223_), .B(new_n2220_), .Y(new_n2224_));
  AOI22X1  g02031(.A0(\a[32] ), .A1(\a[4] ), .B0(\a[25] ), .B1(\a[11] ), .Y(new_n2225_));
  OAI22X1  g02032(.A0(new_n2225_), .A1(new_n2224_), .B0(new_n2223_), .B1(new_n2218_), .Y(new_n2226_));
  NAND4X1  g02033(.A(\a[22] ), .B(\a[20] ), .C(\a[16] ), .D(\a[14] ), .Y(new_n2227_));
  NAND4X1  g02034(.A(\a[22] ), .B(\a[21] ), .C(\a[15] ), .D(\a[14] ), .Y(new_n2228_));
  AOI22X1  g02035(.A0(new_n2228_), .A1(new_n2227_), .B0(new_n1236_), .B1(new_n689_), .Y(new_n2229_));
  NAND2X1  g02036(.A(\a[22] ), .B(\a[14] ), .Y(new_n2230_));
  NAND4X1  g02037(.A(\a[21] ), .B(\a[20] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n2231_));
  NAND3X1  g02038(.A(new_n2228_), .B(new_n2227_), .C(new_n2231_), .Y(new_n2232_));
  AOI22X1  g02039(.A0(\a[21] ), .A1(\a[15] ), .B0(\a[20] ), .B1(\a[16] ), .Y(new_n2233_));
  OAI22X1  g02040(.A0(new_n2233_), .A1(new_n2232_), .B0(new_n2230_), .B1(new_n2229_), .Y(new_n2234_));
  XOR2X1   g02041(.A(new_n2234_), .B(new_n2226_), .Y(new_n2235_));
  XOR2X1   g02042(.A(new_n2235_), .B(new_n2216_), .Y(new_n2236_));
  XOR2X1   g02043(.A(new_n2236_), .B(new_n2208_), .Y(new_n2237_));
  XOR2X1   g02044(.A(new_n2237_), .B(new_n2206_), .Y(new_n2238_));
  AND2X1   g02045(.A(new_n2066_), .B(new_n2064_), .Y(new_n2239_));
  AOI21X1  g02046(.A0(new_n2069_), .A1(new_n2067_), .B0(new_n2239_), .Y(new_n2240_));
  XOR2X1   g02047(.A(new_n2111_), .B(new_n2093_), .Y(new_n2241_));
  XOR2X1   g02048(.A(new_n2241_), .B(new_n2103_), .Y(new_n2242_));
  INVX1    g02049(.A(new_n2122_), .Y(new_n2243_));
  XOR2X1   g02050(.A(new_n2139_), .B(new_n2131_), .Y(new_n2244_));
  XOR2X1   g02051(.A(new_n2244_), .B(new_n2243_), .Y(new_n2245_));
  AND2X1   g02052(.A(new_n2094_), .B(new_n2093_), .Y(new_n2246_));
  OAI21X1  g02053(.A0(new_n2095_), .A1(new_n2246_), .B0(new_n2104_), .Y(new_n2247_));
  OAI21X1  g02054(.A0(new_n2112_), .A1(new_n2105_), .B0(new_n2247_), .Y(new_n2248_));
  XOR2X1   g02055(.A(new_n2248_), .B(new_n2245_), .Y(new_n2249_));
  XOR2X1   g02056(.A(new_n2249_), .B(new_n2242_), .Y(new_n2250_));
  AND2X1   g02057(.A(new_n2250_), .B(new_n2240_), .Y(new_n2251_));
  XOR2X1   g02058(.A(new_n2250_), .B(new_n2240_), .Y(new_n2252_));
  OAI21X1  g02059(.A0(new_n2250_), .A1(new_n2240_), .B0(new_n2238_), .Y(new_n2253_));
  OAI22X1  g02060(.A0(new_n2253_), .A1(new_n2251_), .B0(new_n2252_), .B1(new_n2238_), .Y(new_n2254_));
  XOR2X1   g02061(.A(new_n2254_), .B(new_n2176_), .Y(new_n2255_));
  XOR2X1   g02062(.A(new_n2255_), .B(new_n2154_), .Y(new_n2256_));
  INVX1    g02063(.A(new_n2147_), .Y(new_n2257_));
  OAI21X1  g02064(.A0(new_n2146_), .A1(new_n2050_), .B0(new_n2257_), .Y(new_n2258_));
  XOR2X1   g02065(.A(new_n2258_), .B(new_n2256_), .Y(\asquared[37] ));
  INVX1    g02066(.A(new_n2175_), .Y(new_n2260_));
  OR2X1    g02067(.A(new_n2260_), .B(new_n2156_), .Y(new_n2261_));
  OAI21X1  g02068(.A0(new_n2254_), .A1(new_n2176_), .B0(new_n2261_), .Y(new_n2262_));
  INVX1    g02069(.A(new_n2250_), .Y(new_n2263_));
  NOR2X1   g02070(.A(new_n2263_), .B(new_n2240_), .Y(new_n2264_));
  NOR2X1   g02071(.A(new_n2252_), .B(new_n2238_), .Y(new_n2265_));
  NOR2X1   g02072(.A(new_n2265_), .B(new_n2264_), .Y(new_n2266_));
  INVX1    g02073(.A(new_n2206_), .Y(new_n2267_));
  INVX1    g02074(.A(new_n2236_), .Y(new_n2268_));
  NAND2X1  g02075(.A(new_n2268_), .B(new_n2208_), .Y(new_n2269_));
  OAI21X1  g02076(.A0(new_n2237_), .A1(new_n2267_), .B0(new_n2269_), .Y(new_n2270_));
  AND2X1   g02077(.A(new_n2248_), .B(new_n2245_), .Y(new_n2271_));
  AND2X1   g02078(.A(new_n2249_), .B(new_n2242_), .Y(new_n2272_));
  OR2X1    g02079(.A(new_n2272_), .B(new_n2271_), .Y(new_n2273_));
  INVX1    g02080(.A(new_n2185_), .Y(new_n2274_));
  OR2X1    g02081(.A(new_n2194_), .B(new_n2274_), .Y(new_n2275_));
  OAI21X1  g02082(.A0(new_n2205_), .A1(new_n2195_), .B0(new_n2275_), .Y(new_n2276_));
  NOR2X1   g02083(.A(new_n2111_), .B(new_n2093_), .Y(new_n2277_));
  AOI21X1  g02084(.A0(new_n2241_), .A1(new_n2103_), .B0(new_n2277_), .Y(new_n2278_));
  NAND4X1  g02085(.A(\a[35] ), .B(\a[19] ), .C(\a[17] ), .D(\a[1] ), .Y(new_n2279_));
  AOI21X1  g02086(.A0(\a[36] ), .A1(\a[1] ), .B0(\a[19] ), .Y(new_n2280_));
  AOI21X1  g02087(.A0(new_n814_), .A1(\a[36] ), .B0(new_n2280_), .Y(new_n2281_));
  AND2X1   g02088(.A(new_n2281_), .B(new_n2279_), .Y(new_n2282_));
  XOR2X1   g02089(.A(new_n2281_), .B(new_n2279_), .Y(new_n2283_));
  AND2X1   g02090(.A(new_n814_), .B(\a[36] ), .Y(new_n2284_));
  NOR3X1   g02091(.A(new_n2280_), .B(new_n2284_), .C(new_n2279_), .Y(new_n2285_));
  OAI21X1  g02092(.A0(new_n2285_), .A1(new_n2279_), .B0(new_n2203_), .Y(new_n2286_));
  OAI22X1  g02093(.A0(new_n2286_), .A1(new_n2282_), .B0(new_n2283_), .B1(new_n2203_), .Y(new_n2287_));
  XOR2X1   g02094(.A(new_n2287_), .B(new_n2278_), .Y(new_n2288_));
  XOR2X1   g02095(.A(new_n2288_), .B(new_n2276_), .Y(new_n2289_));
  XOR2X1   g02096(.A(new_n2289_), .B(new_n2273_), .Y(new_n2290_));
  XOR2X1   g02097(.A(new_n2290_), .B(new_n2270_), .Y(new_n2291_));
  NAND2X1  g02098(.A(new_n2291_), .B(new_n2266_), .Y(new_n2292_));
  NOR2X1   g02099(.A(new_n2168_), .B(new_n2166_), .Y(new_n2293_));
  INVX1    g02100(.A(new_n2293_), .Y(new_n2294_));
  OAI21X1  g02101(.A0(new_n2174_), .A1(new_n2170_), .B0(new_n2294_), .Y(new_n2295_));
  INVX1    g02102(.A(new_n2295_), .Y(new_n2296_));
  INVX1    g02103(.A(new_n2192_), .Y(new_n2297_));
  INVX1    g02104(.A(new_n2215_), .Y(new_n2298_));
  NAND2X1  g02105(.A(new_n2298_), .B(new_n2211_), .Y(new_n2299_));
  OAI21X1  g02106(.A0(new_n2210_), .A1(new_n2209_), .B0(new_n2299_), .Y(new_n2300_));
  XOR2X1   g02107(.A(new_n2300_), .B(new_n2297_), .Y(new_n2301_));
  OAI22X1  g02108(.A0(new_n1531_), .A1(new_n866_), .B0(new_n1652_), .B1(new_n583_), .Y(new_n2302_));
  OAI21X1  g02109(.A0(new_n1395_), .A1(new_n867_), .B0(new_n2302_), .Y(new_n2303_));
  AND2X1   g02110(.A(\a[24] ), .B(\a[13] ), .Y(new_n2304_));
  OAI22X1  g02111(.A0(new_n1216_), .A1(new_n490_), .B0(new_n1086_), .B1(new_n549_), .Y(new_n2305_));
  AOI21X1  g02112(.A0(new_n1394_), .A1(new_n691_), .B0(new_n2302_), .Y(new_n2306_));
  AOI22X1  g02113(.A0(new_n2306_), .A1(new_n2305_), .B0(new_n2304_), .B1(new_n2303_), .Y(new_n2307_));
  XOR2X1   g02114(.A(new_n2307_), .B(new_n2301_), .Y(new_n2308_));
  XOR2X1   g02115(.A(new_n2232_), .B(new_n2224_), .Y(new_n2309_));
  XOR2X1   g02116(.A(new_n2309_), .B(new_n2183_), .Y(new_n2310_));
  INVX1    g02117(.A(new_n2216_), .Y(new_n2311_));
  AND2X1   g02118(.A(new_n2234_), .B(new_n2226_), .Y(new_n2312_));
  AOI21X1  g02119(.A0(new_n2235_), .A1(new_n2311_), .B0(new_n2312_), .Y(new_n2313_));
  XOR2X1   g02120(.A(new_n2313_), .B(new_n2310_), .Y(new_n2314_));
  XOR2X1   g02121(.A(new_n2314_), .B(new_n2308_), .Y(new_n2315_));
  XOR2X1   g02122(.A(new_n2315_), .B(new_n2296_), .Y(new_n2316_));
  NOR4X1   g02123(.A(new_n2219_), .B(new_n1679_), .C(new_n570_), .D(new_n255_), .Y(new_n2317_));
  AND2X1   g02124(.A(\a[32] ), .B(\a[26] ), .Y(new_n2318_));
  AOI22X1  g02125(.A0(new_n2318_), .A1(new_n409_), .B0(new_n1995_), .B1(new_n1002_), .Y(new_n2319_));
  OR2X1    g02126(.A(new_n2319_), .B(new_n2317_), .Y(new_n2320_));
  INVX1    g02127(.A(new_n2317_), .Y(new_n2321_));
  AND2X1   g02128(.A(new_n2319_), .B(new_n2321_), .Y(new_n2322_));
  OAI22X1  g02129(.A0(new_n2219_), .A1(new_n255_), .B0(new_n1679_), .B1(new_n570_), .Y(new_n2323_));
  AND2X1   g02130(.A(\a[26] ), .B(\a[11] ), .Y(new_n2324_));
  AOI22X1  g02131(.A0(new_n2324_), .A1(new_n2320_), .B0(new_n2323_), .B1(new_n2322_), .Y(new_n2325_));
  AND2X1   g02132(.A(\a[29] ), .B(\a[8] ), .Y(new_n2326_));
  INVX1    g02133(.A(new_n2326_), .Y(new_n2327_));
  AOI22X1  g02134(.A0(\a[20] ), .A1(\a[17] ), .B0(\a[19] ), .B1(\a[18] ), .Y(new_n2328_));
  AND2X1   g02135(.A(new_n1099_), .B(new_n796_), .Y(new_n2329_));
  NOR3X1   g02136(.A(new_n2328_), .B(new_n2329_), .C(new_n2327_), .Y(new_n2330_));
  INVX1    g02137(.A(new_n2328_), .Y(new_n2331_));
  AOI21X1  g02138(.A0(new_n2331_), .A1(new_n2326_), .B0(new_n2329_), .Y(new_n2332_));
  INVX1    g02139(.A(new_n2332_), .Y(new_n2333_));
  OAI22X1  g02140(.A0(new_n2333_), .A1(new_n2328_), .B0(new_n2330_), .B1(new_n2327_), .Y(new_n2334_));
  XOR2X1   g02141(.A(new_n2334_), .B(new_n2325_), .Y(new_n2335_));
  NOR2X1   g02142(.A(new_n2139_), .B(new_n2131_), .Y(new_n2336_));
  AOI21X1  g02143(.A0(new_n2244_), .A1(new_n2243_), .B0(new_n2336_), .Y(new_n2337_));
  XOR2X1   g02144(.A(new_n2337_), .B(new_n2335_), .Y(new_n2338_));
  NOR2X1   g02145(.A(new_n2160_), .B(new_n2158_), .Y(new_n2339_));
  AOI21X1  g02146(.A0(new_n2165_), .A1(new_n2161_), .B0(new_n2339_), .Y(new_n2340_));
  XOR2X1   g02147(.A(new_n2340_), .B(new_n2338_), .Y(new_n2341_));
  INVX1    g02148(.A(new_n210_), .Y(new_n2342_));
  NAND2X1  g02149(.A(\a[12] ), .B(\a[0] ), .Y(new_n2343_));
  OAI22X1  g02150(.A0(new_n2343_), .A1(new_n1326_), .B0(new_n2342_), .B1(new_n1851_), .Y(new_n2344_));
  INVX1    g02151(.A(\a[37] ), .Y(new_n2345_));
  AND2X1   g02152(.A(\a[33] ), .B(\a[25] ), .Y(new_n2346_));
  AOI21X1  g02153(.A0(new_n2346_), .A1(new_n581_), .B0(new_n2345_), .Y(new_n2347_));
  AND2X1   g02154(.A(new_n2347_), .B(new_n2344_), .Y(new_n2348_));
  AND2X1   g02155(.A(new_n2346_), .B(new_n581_), .Y(new_n2349_));
  AOI21X1  g02156(.A0(new_n2344_), .A1(\a[37] ), .B0(new_n2349_), .Y(new_n2350_));
  INVX1    g02157(.A(new_n2350_), .Y(new_n2351_));
  AOI22X1  g02158(.A0(\a[33] ), .A1(\a[4] ), .B0(\a[25] ), .B1(\a[12] ), .Y(new_n2352_));
  AND2X1   g02159(.A(\a[37] ), .B(\a[0] ), .Y(new_n2353_));
  INVX1    g02160(.A(new_n2353_), .Y(new_n2354_));
  OAI22X1  g02161(.A0(new_n2354_), .A1(new_n2348_), .B0(new_n2352_), .B1(new_n2351_), .Y(new_n2355_));
  AND2X1   g02162(.A(\a[21] ), .B(\a[16] ), .Y(new_n2356_));
  AOI22X1  g02163(.A0(\a[35] ), .A1(\a[2] ), .B0(\a[34] ), .B1(\a[3] ), .Y(new_n2357_));
  INVX1    g02164(.A(new_n2357_), .Y(new_n2358_));
  NAND4X1  g02165(.A(\a[35] ), .B(\a[34] ), .C(\a[3] ), .D(\a[2] ), .Y(new_n2359_));
  NAND3X1  g02166(.A(new_n2358_), .B(new_n2359_), .C(new_n2356_), .Y(new_n2360_));
  AND2X1   g02167(.A(\a[35] ), .B(\a[34] ), .Y(new_n2361_));
  AOI22X1  g02168(.A0(new_n2358_), .A1(new_n2356_), .B0(new_n2361_), .B1(new_n231_), .Y(new_n2362_));
  AOI22X1  g02169(.A0(new_n2362_), .A1(new_n2358_), .B0(new_n2360_), .B1(new_n2356_), .Y(new_n2363_));
  XOR2X1   g02170(.A(new_n2363_), .B(new_n2355_), .Y(new_n2364_));
  INVX1    g02171(.A(new_n2364_), .Y(new_n2365_));
  NAND4X1  g02172(.A(\a[30] ), .B(\a[28] ), .C(\a[9] ), .D(\a[7] ), .Y(new_n2366_));
  NAND4X1  g02173(.A(\a[31] ), .B(\a[28] ), .C(\a[9] ), .D(\a[6] ), .Y(new_n2367_));
  AOI22X1  g02174(.A0(new_n2367_), .A1(new_n2366_), .B0(new_n2075_), .B1(new_n375_), .Y(new_n2368_));
  NOR3X1   g02175(.A(new_n2368_), .B(new_n1431_), .C(new_n341_), .Y(new_n2369_));
  AOI21X1  g02176(.A0(new_n2075_), .A1(new_n375_), .B0(new_n2368_), .Y(new_n2370_));
  OAI22X1  g02177(.A0(new_n1704_), .A1(new_n230_), .B0(new_n1684_), .B1(new_n532_), .Y(new_n2371_));
  AOI21X1  g02178(.A0(new_n2371_), .A1(new_n2370_), .B0(new_n2369_), .Y(new_n2372_));
  XOR2X1   g02179(.A(new_n2372_), .B(new_n2365_), .Y(new_n2373_));
  XOR2X1   g02180(.A(new_n2373_), .B(new_n2341_), .Y(new_n2374_));
  XOR2X1   g02181(.A(new_n2374_), .B(new_n2316_), .Y(new_n2375_));
  INVX1    g02182(.A(new_n2375_), .Y(new_n2376_));
  XOR2X1   g02183(.A(new_n2291_), .B(new_n2266_), .Y(new_n2377_));
  NOR2X1   g02184(.A(new_n2377_), .B(new_n2376_), .Y(new_n2378_));
  NOR2X1   g02185(.A(new_n2291_), .B(new_n2266_), .Y(new_n2379_));
  NOR2X1   g02186(.A(new_n2379_), .B(new_n2375_), .Y(new_n2380_));
  AOI21X1  g02187(.A0(new_n2380_), .A1(new_n2292_), .B0(new_n2378_), .Y(new_n2381_));
  AND2X1   g02188(.A(new_n2381_), .B(new_n2262_), .Y(new_n2382_));
  NOR2X1   g02189(.A(new_n2381_), .B(new_n2262_), .Y(new_n2383_));
  OR2X1    g02190(.A(new_n2383_), .B(new_n2382_), .Y(new_n2384_));
  NOR3X1   g02191(.A(new_n2255_), .B(new_n2152_), .C(new_n2151_), .Y(new_n2385_));
  INVX1    g02192(.A(new_n2385_), .Y(new_n2386_));
  AND2X1   g02193(.A(new_n2255_), .B(new_n2154_), .Y(new_n2387_));
  AOI21X1  g02194(.A0(new_n2258_), .A1(new_n2386_), .B0(new_n2387_), .Y(new_n2388_));
  XOR2X1   g02195(.A(new_n2388_), .B(new_n2384_), .Y(\asquared[38] ));
  INVX1    g02196(.A(new_n2266_), .Y(new_n2390_));
  AOI21X1  g02197(.A0(new_n2291_), .A1(new_n2390_), .B0(new_n2378_), .Y(new_n2391_));
  INVX1    g02198(.A(new_n2338_), .Y(new_n2392_));
  NOR2X1   g02199(.A(new_n2340_), .B(new_n2392_), .Y(new_n2393_));
  NOR2X1   g02200(.A(new_n2373_), .B(new_n2341_), .Y(new_n2394_));
  NOR2X1   g02201(.A(new_n2394_), .B(new_n2393_), .Y(new_n2395_));
  INVX1    g02202(.A(new_n2308_), .Y(new_n2396_));
  NOR2X1   g02203(.A(new_n2313_), .B(new_n2310_), .Y(new_n2397_));
  AOI21X1  g02204(.A0(new_n2314_), .A1(new_n2396_), .B0(new_n2397_), .Y(new_n2398_));
  XOR2X1   g02205(.A(new_n2398_), .B(new_n2395_), .Y(new_n2399_));
  XOR2X1   g02206(.A(new_n2362_), .B(new_n2350_), .Y(new_n2400_));
  INVX1    g02207(.A(new_n2400_), .Y(new_n2401_));
  XOR2X1   g02208(.A(new_n2401_), .B(new_n2306_), .Y(new_n2402_));
  INVX1    g02209(.A(new_n2402_), .Y(new_n2403_));
  INVX1    g02210(.A(new_n2334_), .Y(new_n2404_));
  OR2X1    g02211(.A(new_n2404_), .B(new_n2325_), .Y(new_n2405_));
  OAI21X1  g02212(.A0(new_n2337_), .A1(new_n2335_), .B0(new_n2405_), .Y(new_n2406_));
  XOR2X1   g02213(.A(new_n2406_), .B(new_n2403_), .Y(new_n2407_));
  AND2X1   g02214(.A(\a[33] ), .B(\a[5] ), .Y(new_n2408_));
  INVX1    g02215(.A(new_n2408_), .Y(new_n2409_));
  AND2X1   g02216(.A(\a[32] ), .B(\a[6] ), .Y(new_n2410_));
  AND2X1   g02217(.A(\a[28] ), .B(\a[10] ), .Y(new_n2411_));
  NAND4X1  g02218(.A(\a[33] ), .B(\a[32] ), .C(\a[6] ), .D(\a[5] ), .Y(new_n2412_));
  NAND4X1  g02219(.A(\a[33] ), .B(\a[28] ), .C(\a[10] ), .D(\a[5] ), .Y(new_n2413_));
  AOI22X1  g02220(.A0(new_n2413_), .A1(new_n2412_), .B0(new_n2411_), .B1(new_n2410_), .Y(new_n2414_));
  AND2X1   g02221(.A(new_n2411_), .B(new_n2410_), .Y(new_n2415_));
  NOR2X1   g02222(.A(new_n2414_), .B(new_n2415_), .Y(new_n2416_));
  OAI21X1  g02223(.A0(new_n2411_), .A1(new_n2410_), .B0(new_n2416_), .Y(new_n2417_));
  OAI21X1  g02224(.A0(new_n2414_), .A1(new_n2409_), .B0(new_n2417_), .Y(new_n2418_));
  NAND4X1  g02225(.A(\a[23] ), .B(\a[22] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n2419_));
  NAND4X1  g02226(.A(\a[23] ), .B(\a[21] ), .C(\a[17] ), .D(\a[15] ), .Y(new_n2420_));
  AOI22X1  g02227(.A0(new_n2420_), .A1(new_n2419_), .B0(new_n1154_), .B1(new_n792_), .Y(new_n2421_));
  NAND2X1  g02228(.A(\a[23] ), .B(\a[15] ), .Y(new_n2422_));
  AOI22X1  g02229(.A0(\a[22] ), .A1(\a[16] ), .B0(\a[21] ), .B1(\a[17] ), .Y(new_n2423_));
  AOI21X1  g02230(.A0(new_n1154_), .A1(new_n792_), .B0(new_n2421_), .Y(new_n2424_));
  INVX1    g02231(.A(new_n2424_), .Y(new_n2425_));
  OAI22X1  g02232(.A0(new_n2425_), .A1(new_n2423_), .B0(new_n2422_), .B1(new_n2421_), .Y(new_n2426_));
  XOR2X1   g02233(.A(new_n2426_), .B(new_n2418_), .Y(new_n2427_));
  NAND4X1  g02234(.A(\a[31] ), .B(\a[30] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n2428_));
  AND2X1   g02235(.A(\a[31] ), .B(\a[29] ), .Y(new_n2429_));
  INVX1    g02236(.A(new_n2429_), .Y(new_n2430_));
  OAI22X1  g02237(.A0(new_n2430_), .A1(new_n1023_), .B0(new_n2197_), .B1(new_n366_), .Y(new_n2431_));
  AND2X1   g02238(.A(new_n2431_), .B(new_n2428_), .Y(new_n2432_));
  AND2X1   g02239(.A(\a[29] ), .B(\a[9] ), .Y(new_n2433_));
  INVX1    g02240(.A(new_n2433_), .Y(new_n2434_));
  AOI21X1  g02241(.A0(new_n2075_), .A1(new_n325_), .B0(new_n2431_), .Y(new_n2435_));
  INVX1    g02242(.A(new_n2435_), .Y(new_n2436_));
  AOI22X1  g02243(.A0(\a[31] ), .A1(\a[7] ), .B0(\a[30] ), .B1(\a[8] ), .Y(new_n2437_));
  OAI22X1  g02244(.A0(new_n2437_), .A1(new_n2436_), .B0(new_n2434_), .B1(new_n2432_), .Y(new_n2438_));
  INVX1    g02245(.A(new_n2438_), .Y(new_n2439_));
  XOR2X1   g02246(.A(new_n2439_), .B(new_n2427_), .Y(new_n2440_));
  XOR2X1   g02247(.A(new_n2440_), .B(new_n2407_), .Y(new_n2441_));
  XOR2X1   g02248(.A(new_n2441_), .B(new_n2399_), .Y(new_n2442_));
  INVX1    g02249(.A(new_n2442_), .Y(new_n2443_));
  NOR2X1   g02250(.A(new_n2315_), .B(new_n2296_), .Y(new_n2444_));
  AOI21X1  g02251(.A0(new_n2374_), .A1(new_n2316_), .B0(new_n2444_), .Y(new_n2445_));
  XOR2X1   g02252(.A(new_n2445_), .B(new_n2443_), .Y(new_n2446_));
  AND2X1   g02253(.A(new_n2289_), .B(new_n2273_), .Y(new_n2447_));
  AND2X1   g02254(.A(new_n2290_), .B(new_n2270_), .Y(new_n2448_));
  OR2X1    g02255(.A(new_n2448_), .B(new_n2447_), .Y(new_n2449_));
  NOR2X1   g02256(.A(new_n2300_), .B(new_n2297_), .Y(new_n2450_));
  NAND2X1  g02257(.A(new_n2300_), .B(new_n2297_), .Y(new_n2451_));
  OAI21X1  g02258(.A0(new_n2307_), .A1(new_n2450_), .B0(new_n2451_), .Y(new_n2452_));
  INVX1    g02259(.A(new_n2355_), .Y(new_n2453_));
  OR2X1    g02260(.A(new_n2363_), .B(new_n2453_), .Y(new_n2454_));
  OAI21X1  g02261(.A0(new_n2372_), .A1(new_n2364_), .B0(new_n2454_), .Y(new_n2455_));
  XOR2X1   g02262(.A(new_n2455_), .B(new_n2452_), .Y(new_n2456_));
  AND2X1   g02263(.A(\a[37] ), .B(\a[1] ), .Y(new_n2457_));
  XOR2X1   g02264(.A(new_n2457_), .B(new_n992_), .Y(new_n2458_));
  XOR2X1   g02265(.A(new_n2458_), .B(new_n2332_), .Y(new_n2459_));
  XOR2X1   g02266(.A(new_n2459_), .B(new_n2370_), .Y(new_n2460_));
  XOR2X1   g02267(.A(new_n2460_), .B(new_n2456_), .Y(new_n2461_));
  XOR2X1   g02268(.A(new_n2461_), .B(new_n2449_), .Y(new_n2462_));
  NOR2X1   g02269(.A(new_n2283_), .B(new_n2203_), .Y(new_n2463_));
  NOR2X1   g02270(.A(new_n2463_), .B(new_n2285_), .Y(new_n2464_));
  INVX1    g02271(.A(new_n2464_), .Y(new_n2465_));
  NOR3X1   g02272(.A(new_n517_), .B(new_n2028_), .C(new_n1679_), .Y(new_n2466_));
  AND2X1   g02273(.A(\a[26] ), .B(\a[4] ), .Y(new_n2467_));
  AND2X1   g02274(.A(\a[34] ), .B(\a[12] ), .Y(new_n2468_));
  AOI22X1  g02275(.A0(new_n2468_), .A1(new_n2467_), .B0(new_n1995_), .B1(new_n482_), .Y(new_n2469_));
  OR2X1    g02276(.A(new_n2469_), .B(new_n2466_), .Y(new_n2470_));
  AND2X1   g02277(.A(\a[26] ), .B(\a[12] ), .Y(new_n2471_));
  INVX1    g02278(.A(new_n2466_), .Y(new_n2472_));
  AND2X1   g02279(.A(new_n2469_), .B(new_n2472_), .Y(new_n2473_));
  OAI22X1  g02280(.A0(new_n2028_), .A1(new_n340_), .B0(new_n1679_), .B1(new_n488_), .Y(new_n2474_));
  AOI22X1  g02281(.A0(new_n2474_), .A1(new_n2473_), .B0(new_n2471_), .B1(new_n2470_), .Y(new_n2475_));
  XOR2X1   g02282(.A(new_n2475_), .B(new_n2465_), .Y(new_n2476_));
  AND2X1   g02283(.A(new_n2232_), .B(new_n2224_), .Y(new_n2477_));
  AOI21X1  g02284(.A0(new_n2309_), .A1(new_n2184_), .B0(new_n2477_), .Y(new_n2478_));
  XOR2X1   g02285(.A(new_n2478_), .B(new_n2476_), .Y(new_n2479_));
  NOR2X1   g02286(.A(new_n2287_), .B(new_n2278_), .Y(new_n2480_));
  AOI21X1  g02287(.A0(new_n2288_), .A1(new_n2276_), .B0(new_n2480_), .Y(new_n2481_));
  AOI22X1  g02288(.A0(\a[38] ), .A1(\a[0] ), .B0(\a[36] ), .B1(\a[2] ), .Y(new_n2482_));
  INVX1    g02289(.A(new_n2482_), .Y(new_n2483_));
  AND2X1   g02290(.A(\a[38] ), .B(\a[36] ), .Y(new_n2484_));
  AND2X1   g02291(.A(new_n2484_), .B(new_n197_), .Y(new_n2485_));
  AOI21X1  g02292(.A0(new_n2483_), .A1(new_n2284_), .B0(new_n2485_), .Y(new_n2486_));
  INVX1    g02293(.A(new_n2486_), .Y(new_n2487_));
  OAI21X1  g02294(.A0(new_n2485_), .A1(new_n2482_), .B0(new_n2284_), .Y(new_n2488_));
  OAI21X1  g02295(.A0(new_n2487_), .A1(new_n2482_), .B0(new_n2488_), .Y(new_n2489_));
  XOR2X1   g02296(.A(new_n2489_), .B(new_n2322_), .Y(new_n2490_));
  INVX1    g02297(.A(new_n2490_), .Y(new_n2491_));
  AND2X1   g02298(.A(\a[35] ), .B(\a[3] ), .Y(new_n2492_));
  AOI22X1  g02299(.A0(\a[25] ), .A1(\a[13] ), .B0(\a[24] ), .B1(\a[14] ), .Y(new_n2493_));
  INVX1    g02300(.A(new_n2493_), .Y(new_n2494_));
  NAND4X1  g02301(.A(\a[25] ), .B(\a[24] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n2495_));
  NAND3X1  g02302(.A(new_n2494_), .B(new_n2495_), .C(new_n2492_), .Y(new_n2496_));
  AOI22X1  g02303(.A0(new_n2494_), .A1(new_n2492_), .B0(new_n1532_), .B1(new_n582_), .Y(new_n2497_));
  AOI22X1  g02304(.A0(new_n2497_), .A1(new_n2494_), .B0(new_n2496_), .B1(new_n2492_), .Y(new_n2498_));
  XOR2X1   g02305(.A(new_n2498_), .B(new_n2491_), .Y(new_n2499_));
  XOR2X1   g02306(.A(new_n2499_), .B(new_n2481_), .Y(new_n2500_));
  XOR2X1   g02307(.A(new_n2500_), .B(new_n2479_), .Y(new_n2501_));
  XOR2X1   g02308(.A(new_n2501_), .B(new_n2462_), .Y(new_n2502_));
  XOR2X1   g02309(.A(new_n2502_), .B(new_n2446_), .Y(new_n2503_));
  INVX1    g02310(.A(new_n2503_), .Y(new_n2504_));
  XOR2X1   g02311(.A(new_n2504_), .B(new_n2391_), .Y(new_n2505_));
  INVX1    g02312(.A(new_n2382_), .Y(new_n2506_));
  OAI21X1  g02313(.A0(new_n2388_), .A1(new_n2383_), .B0(new_n2506_), .Y(new_n2507_));
  XOR2X1   g02314(.A(new_n2507_), .B(new_n2505_), .Y(\asquared[39] ));
  NOR2X1   g02315(.A(new_n2445_), .B(new_n2443_), .Y(new_n2509_));
  AOI21X1  g02316(.A0(new_n2502_), .A1(new_n2446_), .B0(new_n2509_), .Y(new_n2510_));
  AND2X1   g02317(.A(new_n2461_), .B(new_n2449_), .Y(new_n2511_));
  AOI21X1  g02318(.A0(new_n2501_), .A1(new_n2462_), .B0(new_n2511_), .Y(new_n2512_));
  INVX1    g02319(.A(new_n2512_), .Y(new_n2513_));
  NOR2X1   g02320(.A(new_n2499_), .B(new_n2481_), .Y(new_n2514_));
  AOI21X1  g02321(.A0(new_n2500_), .A1(new_n2479_), .B0(new_n2514_), .Y(new_n2515_));
  NAND4X1  g02322(.A(\a[37] ), .B(\a[20] ), .C(\a[18] ), .D(\a[1] ), .Y(new_n2516_));
  AND2X1   g02323(.A(\a[39] ), .B(\a[0] ), .Y(new_n2517_));
  XOR2X1   g02324(.A(new_n2517_), .B(new_n2516_), .Y(new_n2518_));
  INVX1    g02325(.A(\a[38] ), .Y(new_n2519_));
  OAI21X1  g02326(.A0(new_n2519_), .A1(new_n202_), .B0(\a[20] ), .Y(new_n2520_));
  NAND3X1  g02327(.A(\a[38] ), .B(new_n934_), .C(\a[1] ), .Y(new_n2521_));
  AND2X1   g02328(.A(new_n2521_), .B(new_n2520_), .Y(new_n2522_));
  XOR2X1   g02329(.A(new_n2522_), .B(new_n2518_), .Y(new_n2523_));
  OAI21X1  g02330(.A0(new_n2330_), .A1(new_n2329_), .B0(new_n2458_), .Y(new_n2524_));
  OAI21X1  g02331(.A0(new_n2459_), .A1(new_n2370_), .B0(new_n2524_), .Y(new_n2525_));
  XOR2X1   g02332(.A(new_n2525_), .B(new_n2523_), .Y(new_n2526_));
  OR2X1    g02333(.A(new_n2362_), .B(new_n2350_), .Y(new_n2527_));
  OAI21X1  g02334(.A0(new_n2401_), .A1(new_n2306_), .B0(new_n2527_), .Y(new_n2528_));
  XOR2X1   g02335(.A(new_n2528_), .B(new_n2526_), .Y(new_n2529_));
  INVX1    g02336(.A(new_n2529_), .Y(new_n2530_));
  XOR2X1   g02337(.A(new_n2497_), .B(new_n2486_), .Y(new_n2531_));
  XOR2X1   g02338(.A(new_n2531_), .B(new_n2424_), .Y(new_n2532_));
  AND2X1   g02339(.A(new_n2426_), .B(new_n2418_), .Y(new_n2533_));
  AOI21X1  g02340(.A0(new_n2438_), .A1(new_n2427_), .B0(new_n2533_), .Y(new_n2534_));
  INVX1    g02341(.A(new_n2534_), .Y(new_n2535_));
  INVX1    g02342(.A(new_n2322_), .Y(new_n2536_));
  NOR2X1   g02343(.A(new_n2498_), .B(new_n2490_), .Y(new_n2537_));
  AOI21X1  g02344(.A0(new_n2489_), .A1(new_n2536_), .B0(new_n2537_), .Y(new_n2538_));
  XOR2X1   g02345(.A(new_n2538_), .B(new_n2535_), .Y(new_n2539_));
  XOR2X1   g02346(.A(new_n2539_), .B(new_n2532_), .Y(new_n2540_));
  XOR2X1   g02347(.A(new_n2540_), .B(new_n2530_), .Y(new_n2541_));
  XOR2X1   g02348(.A(new_n2541_), .B(new_n2515_), .Y(new_n2542_));
  XOR2X1   g02349(.A(new_n2542_), .B(new_n2513_), .Y(new_n2543_));
  INVX1    g02350(.A(new_n2543_), .Y(new_n2544_));
  NOR2X1   g02351(.A(new_n2398_), .B(new_n2395_), .Y(new_n2545_));
  AOI21X1  g02352(.A0(new_n2441_), .A1(new_n2399_), .B0(new_n2545_), .Y(new_n2546_));
  INVX1    g02353(.A(new_n2416_), .Y(new_n2547_));
  XOR2X1   g02354(.A(new_n2473_), .B(new_n2435_), .Y(new_n2548_));
  XOR2X1   g02355(.A(new_n2548_), .B(new_n2547_), .Y(new_n2549_));
  INVX1    g02356(.A(new_n2549_), .Y(new_n2550_));
  OR2X1    g02357(.A(new_n2475_), .B(new_n2464_), .Y(new_n2551_));
  OAI21X1  g02358(.A0(new_n2478_), .A1(new_n2476_), .B0(new_n2551_), .Y(new_n2552_));
  XOR2X1   g02359(.A(new_n2552_), .B(new_n2550_), .Y(new_n2553_));
  AOI22X1  g02360(.A0(\a[35] ), .A1(\a[4] ), .B0(\a[27] ), .B1(\a[12] ), .Y(new_n2554_));
  AND2X1   g02361(.A(\a[22] ), .B(\a[17] ), .Y(new_n2555_));
  INVX1    g02362(.A(new_n2555_), .Y(new_n2556_));
  INVX1    g02363(.A(\a[35] ), .Y(new_n2557_));
  NOR4X1   g02364(.A(new_n2557_), .B(new_n1679_), .C(new_n453_), .D(new_n340_), .Y(new_n2558_));
  NOR3X1   g02365(.A(new_n2556_), .B(new_n2558_), .C(new_n2554_), .Y(new_n2559_));
  NOR2X1   g02366(.A(new_n2559_), .B(new_n2558_), .Y(new_n2560_));
  INVX1    g02367(.A(new_n2560_), .Y(new_n2561_));
  OAI22X1  g02368(.A0(new_n2561_), .A1(new_n2554_), .B0(new_n2559_), .B1(new_n2556_), .Y(new_n2562_));
  AND2X1   g02369(.A(\a[31] ), .B(\a[8] ), .Y(new_n2563_));
  AOI22X1  g02370(.A0(\a[21] ), .A1(\a[18] ), .B0(\a[20] ), .B1(\a[19] ), .Y(new_n2564_));
  INVX1    g02371(.A(new_n2564_), .Y(new_n2565_));
  NAND4X1  g02372(.A(\a[21] ), .B(\a[20] ), .C(\a[19] ), .D(\a[18] ), .Y(new_n2566_));
  NAND3X1  g02373(.A(new_n2565_), .B(new_n2566_), .C(new_n2563_), .Y(new_n2567_));
  AOI22X1  g02374(.A0(new_n2565_), .A1(new_n2563_), .B0(new_n1236_), .B1(new_n855_), .Y(new_n2568_));
  AOI22X1  g02375(.A0(new_n2568_), .A1(new_n2565_), .B0(new_n2567_), .B1(new_n2563_), .Y(new_n2569_));
  XOR2X1   g02376(.A(new_n2569_), .B(new_n2562_), .Y(new_n2570_));
  INVX1    g02377(.A(new_n2570_), .Y(new_n2571_));
  NOR4X1   g02378(.A(new_n2028_), .B(new_n1803_), .C(new_n570_), .D(new_n255_), .Y(new_n2572_));
  AND2X1   g02379(.A(\a[34] ), .B(\a[5] ), .Y(new_n2573_));
  AOI22X1  g02380(.A0(new_n2573_), .A1(new_n1434_), .B0(new_n1674_), .B1(new_n1002_), .Y(new_n2574_));
  OR2X1    g02381(.A(new_n2574_), .B(new_n2572_), .Y(new_n2575_));
  INVX1    g02382(.A(new_n2572_), .Y(new_n2576_));
  AND2X1   g02383(.A(new_n2574_), .B(new_n2576_), .Y(new_n2577_));
  OAI22X1  g02384(.A0(new_n2028_), .A1(new_n255_), .B0(new_n1803_), .B1(new_n570_), .Y(new_n2578_));
  AOI22X1  g02385(.A0(new_n2578_), .A1(new_n2577_), .B0(new_n2575_), .B1(new_n1434_), .Y(new_n2579_));
  XOR2X1   g02386(.A(new_n2579_), .B(new_n2571_), .Y(new_n2580_));
  XOR2X1   g02387(.A(new_n2580_), .B(new_n2553_), .Y(new_n2581_));
  XOR2X1   g02388(.A(new_n2581_), .B(new_n2546_), .Y(new_n2582_));
  INVX1    g02389(.A(\a[36] ), .Y(new_n2583_));
  NOR4X1   g02390(.A(new_n2583_), .B(new_n1263_), .C(new_n591_), .D(new_n223_), .Y(new_n2584_));
  NAND4X1  g02391(.A(\a[37] ), .B(\a[36] ), .C(\a[3] ), .D(\a[2] ), .Y(new_n2585_));
  NAND4X1  g02392(.A(\a[37] ), .B(\a[26] ), .C(\a[13] ), .D(\a[2] ), .Y(new_n2586_));
  AOI21X1  g02393(.A0(new_n2586_), .A1(new_n2585_), .B0(new_n2584_), .Y(new_n2587_));
  OR2X1    g02394(.A(new_n2587_), .B(new_n2584_), .Y(new_n2588_));
  AOI22X1  g02395(.A0(\a[36] ), .A1(\a[3] ), .B0(\a[26] ), .B1(\a[13] ), .Y(new_n2589_));
  NAND2X1  g02396(.A(\a[37] ), .B(\a[2] ), .Y(new_n2590_));
  OAI22X1  g02397(.A0(new_n2590_), .A1(new_n2587_), .B0(new_n2589_), .B1(new_n2588_), .Y(new_n2591_));
  AOI22X1  g02398(.A0(new_n1532_), .A1(new_n691_), .B0(new_n1134_), .B1(new_n690_), .Y(new_n2592_));
  AOI21X1  g02399(.A0(new_n1219_), .A1(new_n689_), .B0(new_n2592_), .Y(new_n2593_));
  NAND2X1  g02400(.A(\a[25] ), .B(\a[14] ), .Y(new_n2594_));
  OAI21X1  g02401(.A0(new_n1652_), .A1(new_n1024_), .B0(new_n2592_), .Y(new_n2595_));
  AOI22X1  g02402(.A0(\a[24] ), .A1(\a[15] ), .B0(\a[23] ), .B1(\a[16] ), .Y(new_n2596_));
  OAI22X1  g02403(.A0(new_n2596_), .A1(new_n2595_), .B0(new_n2594_), .B1(new_n2593_), .Y(new_n2597_));
  XOR2X1   g02404(.A(new_n2597_), .B(new_n2591_), .Y(new_n2598_));
  AND2X1   g02405(.A(\a[33] ), .B(\a[6] ), .Y(new_n2599_));
  INVX1    g02406(.A(new_n2599_), .Y(new_n2600_));
  NAND4X1  g02407(.A(\a[33] ), .B(\a[32] ), .C(\a[7] ), .D(\a[6] ), .Y(new_n2601_));
  NAND4X1  g02408(.A(\a[33] ), .B(\a[30] ), .C(\a[9] ), .D(\a[6] ), .Y(new_n2602_));
  AOI22X1  g02409(.A0(new_n2602_), .A1(new_n2601_), .B0(new_n1787_), .B1(new_n596_), .Y(new_n2603_));
  AOI21X1  g02410(.A0(new_n1787_), .A1(new_n596_), .B0(new_n2603_), .Y(new_n2604_));
  INVX1    g02411(.A(new_n2604_), .Y(new_n2605_));
  AOI22X1  g02412(.A0(\a[32] ), .A1(\a[7] ), .B0(\a[30] ), .B1(\a[9] ), .Y(new_n2606_));
  OAI22X1  g02413(.A0(new_n2606_), .A1(new_n2605_), .B0(new_n2603_), .B1(new_n2600_), .Y(new_n2607_));
  INVX1    g02414(.A(new_n2607_), .Y(new_n2608_));
  XOR2X1   g02415(.A(new_n2608_), .B(new_n2598_), .Y(new_n2609_));
  AND2X1   g02416(.A(new_n2455_), .B(new_n2452_), .Y(new_n2610_));
  AOI21X1  g02417(.A0(new_n2460_), .A1(new_n2456_), .B0(new_n2610_), .Y(new_n2611_));
  XOR2X1   g02418(.A(new_n2611_), .B(new_n2609_), .Y(new_n2612_));
  NAND2X1  g02419(.A(new_n2406_), .B(new_n2402_), .Y(new_n2613_));
  OAI21X1  g02420(.A0(new_n2440_), .A1(new_n2407_), .B0(new_n2613_), .Y(new_n2614_));
  XOR2X1   g02421(.A(new_n2614_), .B(new_n2612_), .Y(new_n2615_));
  XOR2X1   g02422(.A(new_n2615_), .B(new_n2582_), .Y(new_n2616_));
  XOR2X1   g02423(.A(new_n2616_), .B(new_n2544_), .Y(new_n2617_));
  XOR2X1   g02424(.A(new_n2617_), .B(new_n2510_), .Y(new_n2618_));
  NOR2X1   g02425(.A(new_n2504_), .B(new_n2391_), .Y(new_n2619_));
  AND2X1   g02426(.A(new_n2504_), .B(new_n2391_), .Y(new_n2620_));
  INVX1    g02427(.A(new_n2620_), .Y(new_n2621_));
  AOI21X1  g02428(.A0(new_n2507_), .A1(new_n2621_), .B0(new_n2619_), .Y(new_n2622_));
  XOR2X1   g02429(.A(new_n2622_), .B(new_n2618_), .Y(\asquared[40] ));
  NAND2X1  g02430(.A(new_n2542_), .B(new_n2513_), .Y(new_n2624_));
  OAI21X1  g02431(.A0(new_n2616_), .A1(new_n2544_), .B0(new_n2624_), .Y(new_n2625_));
  NOR2X1   g02432(.A(new_n2611_), .B(new_n2609_), .Y(new_n2626_));
  AOI21X1  g02433(.A0(new_n2614_), .A1(new_n2612_), .B0(new_n2626_), .Y(new_n2627_));
  NAND2X1  g02434(.A(new_n2552_), .B(new_n2549_), .Y(new_n2628_));
  OAI21X1  g02435(.A0(new_n2580_), .A1(new_n2553_), .B0(new_n2628_), .Y(new_n2629_));
  INVX1    g02436(.A(new_n2577_), .Y(new_n2630_));
  XOR2X1   g02437(.A(new_n2588_), .B(new_n2630_), .Y(new_n2631_));
  XOR2X1   g02438(.A(new_n2631_), .B(new_n2561_), .Y(new_n2632_));
  INVX1    g02439(.A(new_n2562_), .Y(new_n2633_));
  OR2X1    g02440(.A(new_n2579_), .B(new_n2570_), .Y(new_n2634_));
  OAI21X1  g02441(.A0(new_n2569_), .A1(new_n2633_), .B0(new_n2634_), .Y(new_n2635_));
  AND2X1   g02442(.A(new_n2597_), .B(new_n2591_), .Y(new_n2636_));
  AND2X1   g02443(.A(new_n2607_), .B(new_n2598_), .Y(new_n2637_));
  OR2X1    g02444(.A(new_n2637_), .B(new_n2636_), .Y(new_n2638_));
  XOR2X1   g02445(.A(new_n2638_), .B(new_n2635_), .Y(new_n2639_));
  XOR2X1   g02446(.A(new_n2639_), .B(new_n2632_), .Y(new_n2640_));
  XOR2X1   g02447(.A(new_n2640_), .B(new_n2629_), .Y(new_n2641_));
  INVX1    g02448(.A(new_n2641_), .Y(new_n2642_));
  XOR2X1   g02449(.A(new_n2642_), .B(new_n2627_), .Y(new_n2643_));
  INVX1    g02450(.A(new_n2546_), .Y(new_n2644_));
  AND2X1   g02451(.A(new_n2581_), .B(new_n2644_), .Y(new_n2645_));
  INVX1    g02452(.A(new_n2582_), .Y(new_n2646_));
  AOI21X1  g02453(.A0(new_n2615_), .A1(new_n2646_), .B0(new_n2645_), .Y(new_n2647_));
  OR2X1    g02454(.A(new_n2647_), .B(new_n2643_), .Y(new_n2648_));
  INVX1    g02455(.A(new_n2643_), .Y(new_n2649_));
  XOR2X1   g02456(.A(new_n2647_), .B(new_n2649_), .Y(new_n2650_));
  XOR2X1   g02457(.A(new_n2605_), .B(new_n2595_), .Y(new_n2651_));
  INVX1    g02458(.A(\a[39] ), .Y(new_n2652_));
  NOR3X1   g02459(.A(new_n2516_), .B(new_n2652_), .C(new_n194_), .Y(new_n2653_));
  AOI21X1  g02460(.A0(new_n2521_), .A1(new_n2520_), .B0(new_n2518_), .Y(new_n2654_));
  NOR2X1   g02461(.A(new_n2654_), .B(new_n2653_), .Y(new_n2655_));
  XOR2X1   g02462(.A(new_n2655_), .B(new_n2651_), .Y(new_n2656_));
  AND2X1   g02463(.A(new_n2525_), .B(new_n2523_), .Y(new_n2657_));
  AOI21X1  g02464(.A0(new_n2528_), .A1(new_n2526_), .B0(new_n2657_), .Y(new_n2658_));
  XOR2X1   g02465(.A(new_n2658_), .B(new_n2656_), .Y(new_n2659_));
  AND2X1   g02466(.A(\a[22] ), .B(\a[18] ), .Y(new_n2660_));
  INVX1    g02467(.A(new_n2660_), .Y(new_n2661_));
  AOI22X1  g02468(.A0(\a[40] ), .A1(\a[0] ), .B0(\a[38] ), .B1(\a[2] ), .Y(new_n2662_));
  AND2X1   g02469(.A(\a[40] ), .B(\a[38] ), .Y(new_n2663_));
  AND2X1   g02470(.A(new_n2663_), .B(new_n197_), .Y(new_n2664_));
  NOR3X1   g02471(.A(new_n2664_), .B(new_n2662_), .C(new_n2661_), .Y(new_n2665_));
  INVX1    g02472(.A(new_n2662_), .Y(new_n2666_));
  AOI21X1  g02473(.A0(new_n2666_), .A1(new_n2660_), .B0(new_n2664_), .Y(new_n2667_));
  INVX1    g02474(.A(new_n2667_), .Y(new_n2668_));
  OAI22X1  g02475(.A0(new_n2668_), .A1(new_n2662_), .B0(new_n2665_), .B1(new_n2661_), .Y(new_n2669_));
  AND2X1   g02476(.A(\a[33] ), .B(\a[7] ), .Y(new_n2670_));
  AND2X1   g02477(.A(\a[32] ), .B(\a[31] ), .Y(new_n2671_));
  INVX1    g02478(.A(new_n2671_), .Y(new_n2672_));
  NAND2X1  g02479(.A(\a[33] ), .B(\a[31] ), .Y(new_n2673_));
  AND2X1   g02480(.A(\a[33] ), .B(\a[32] ), .Y(new_n2674_));
  INVX1    g02481(.A(new_n2674_), .Y(new_n2675_));
  OAI22X1  g02482(.A0(new_n2675_), .A1(new_n445_), .B0(new_n2673_), .B1(new_n1023_), .Y(new_n2676_));
  OAI21X1  g02483(.A0(new_n2672_), .A1(new_n366_), .B0(new_n2676_), .Y(new_n2677_));
  AOI21X1  g02484(.A0(new_n2671_), .A1(new_n1030_), .B0(new_n2676_), .Y(new_n2678_));
  OAI22X1  g02485(.A0(new_n2219_), .A1(new_n413_), .B0(new_n1704_), .B1(new_n341_), .Y(new_n2679_));
  AOI22X1  g02486(.A0(new_n2679_), .A1(new_n2678_), .B0(new_n2677_), .B1(new_n2670_), .Y(new_n2680_));
  XOR2X1   g02487(.A(new_n2680_), .B(new_n2669_), .Y(new_n2681_));
  AND2X1   g02488(.A(\a[36] ), .B(\a[35] ), .Y(new_n2682_));
  NOR4X1   g02489(.A(new_n2583_), .B(new_n1431_), .C(new_n453_), .D(new_n340_), .Y(new_n2683_));
  AOI21X1  g02490(.A0(new_n2682_), .A1(new_n218_), .B0(new_n2683_), .Y(new_n2684_));
  NOR4X1   g02491(.A(new_n2557_), .B(new_n1431_), .C(new_n453_), .D(new_n255_), .Y(new_n2685_));
  OR2X1    g02492(.A(new_n2685_), .B(new_n2684_), .Y(new_n2686_));
  AND2X1   g02493(.A(\a[36] ), .B(\a[4] ), .Y(new_n2687_));
  AND2X1   g02494(.A(new_n2682_), .B(new_n218_), .Y(new_n2688_));
  NOR3X1   g02495(.A(new_n2685_), .B(new_n2683_), .C(new_n2688_), .Y(new_n2689_));
  OAI22X1  g02496(.A0(new_n2557_), .A1(new_n255_), .B0(new_n1431_), .B1(new_n453_), .Y(new_n2690_));
  AOI22X1  g02497(.A0(new_n2690_), .A1(new_n2689_), .B0(new_n2687_), .B1(new_n2686_), .Y(new_n2691_));
  XOR2X1   g02498(.A(new_n2691_), .B(new_n2681_), .Y(new_n2692_));
  XOR2X1   g02499(.A(new_n2692_), .B(new_n2659_), .Y(new_n2693_));
  NAND2X1  g02500(.A(new_n2540_), .B(new_n2529_), .Y(new_n2694_));
  OAI21X1  g02501(.A0(new_n2541_), .A1(new_n2515_), .B0(new_n2694_), .Y(new_n2695_));
  XOR2X1   g02502(.A(new_n2695_), .B(new_n2693_), .Y(new_n2696_));
  AOI22X1  g02503(.A0(\a[27] ), .A1(\a[13] ), .B0(\a[26] ), .B1(\a[14] ), .Y(new_n2697_));
  AND2X1   g02504(.A(\a[37] ), .B(\a[3] ), .Y(new_n2698_));
  INVX1    g02505(.A(new_n2698_), .Y(new_n2699_));
  AND2X1   g02506(.A(new_n1995_), .B(new_n582_), .Y(new_n2700_));
  NOR3X1   g02507(.A(new_n2699_), .B(new_n2700_), .C(new_n2697_), .Y(new_n2701_));
  NOR2X1   g02508(.A(new_n2701_), .B(new_n2700_), .Y(new_n2702_));
  INVX1    g02509(.A(new_n2702_), .Y(new_n2703_));
  OAI22X1  g02510(.A0(new_n2703_), .A1(new_n2697_), .B0(new_n2701_), .B1(new_n2699_), .Y(new_n2704_));
  INVX1    g02511(.A(new_n753_), .Y(new_n2705_));
  INVX1    g02512(.A(new_n1134_), .Y(new_n2706_));
  OAI22X1  g02513(.A0(new_n1772_), .A1(new_n1024_), .B0(new_n2706_), .B1(new_n2705_), .Y(new_n2707_));
  OAI21X1  g02514(.A0(new_n1652_), .A1(new_n793_), .B0(new_n2707_), .Y(new_n2708_));
  AND2X1   g02515(.A(\a[25] ), .B(\a[15] ), .Y(new_n2709_));
  AOI21X1  g02516(.A0(new_n1219_), .A1(new_n792_), .B0(new_n2707_), .Y(new_n2710_));
  OAI22X1  g02517(.A0(new_n1185_), .A1(new_n571_), .B0(new_n1216_), .B1(new_n616_), .Y(new_n2711_));
  AOI22X1  g02518(.A0(new_n2711_), .A1(new_n2710_), .B0(new_n2709_), .B1(new_n2708_), .Y(new_n2712_));
  XOR2X1   g02519(.A(new_n2712_), .B(new_n2704_), .Y(new_n2713_));
  NOR4X1   g02520(.A(new_n2028_), .B(new_n1684_), .C(new_n570_), .D(new_n230_), .Y(new_n2714_));
  AND2X1   g02521(.A(new_n2196_), .B(new_n1002_), .Y(new_n2715_));
  NOR4X1   g02522(.A(new_n2028_), .B(new_n1803_), .C(new_n488_), .D(new_n230_), .Y(new_n2716_));
  NOR2X1   g02523(.A(new_n2716_), .B(new_n2715_), .Y(new_n2717_));
  NOR2X1   g02524(.A(new_n2717_), .B(new_n2714_), .Y(new_n2718_));
  NOR3X1   g02525(.A(new_n2718_), .B(new_n1803_), .C(new_n488_), .Y(new_n2719_));
  NOR3X1   g02526(.A(new_n2716_), .B(new_n2715_), .C(new_n2714_), .Y(new_n2720_));
  OAI22X1  g02527(.A0(new_n2028_), .A1(new_n230_), .B0(new_n1684_), .B1(new_n570_), .Y(new_n2721_));
  AOI21X1  g02528(.A0(new_n2721_), .A1(new_n2720_), .B0(new_n2719_), .Y(new_n2722_));
  XOR2X1   g02529(.A(new_n2722_), .B(new_n2713_), .Y(new_n2723_));
  OR2X1    g02530(.A(new_n2538_), .B(new_n2534_), .Y(new_n2724_));
  OAI21X1  g02531(.A0(new_n2539_), .A1(new_n2532_), .B0(new_n2724_), .Y(new_n2725_));
  XOR2X1   g02532(.A(new_n2725_), .B(new_n2723_), .Y(new_n2726_));
  NOR2X1   g02533(.A(new_n2473_), .B(new_n2435_), .Y(new_n2727_));
  AOI21X1  g02534(.A0(new_n2548_), .A1(new_n2547_), .B0(new_n2727_), .Y(new_n2728_));
  NOR2X1   g02535(.A(new_n2497_), .B(new_n2486_), .Y(new_n2729_));
  AOI21X1  g02536(.A0(new_n2531_), .A1(new_n2425_), .B0(new_n2729_), .Y(new_n2730_));
  XOR2X1   g02537(.A(new_n2730_), .B(new_n2728_), .Y(new_n2731_));
  INVX1    g02538(.A(new_n2568_), .Y(new_n2732_));
  AND2X1   g02539(.A(new_n894_), .B(\a[38] ), .Y(new_n2733_));
  AND2X1   g02540(.A(\a[39] ), .B(\a[1] ), .Y(new_n2734_));
  XOR2X1   g02541(.A(new_n2734_), .B(new_n1148_), .Y(new_n2735_));
  XOR2X1   g02542(.A(new_n2735_), .B(new_n2733_), .Y(new_n2736_));
  XOR2X1   g02543(.A(new_n2736_), .B(new_n2732_), .Y(new_n2737_));
  XOR2X1   g02544(.A(new_n2737_), .B(new_n2731_), .Y(new_n2738_));
  XOR2X1   g02545(.A(new_n2738_), .B(new_n2726_), .Y(new_n2739_));
  XOR2X1   g02546(.A(new_n2739_), .B(new_n2696_), .Y(new_n2740_));
  AOI21X1  g02547(.A0(new_n2647_), .A1(new_n2643_), .B0(new_n2740_), .Y(new_n2741_));
  AOI22X1  g02548(.A0(new_n2741_), .A1(new_n2648_), .B0(new_n2740_), .B1(new_n2650_), .Y(new_n2742_));
  AND2X1   g02549(.A(new_n2742_), .B(new_n2625_), .Y(new_n2743_));
  INVX1    g02550(.A(new_n2743_), .Y(new_n2744_));
  INVX1    g02551(.A(new_n2617_), .Y(new_n2745_));
  NOR2X1   g02552(.A(new_n2745_), .B(new_n2510_), .Y(new_n2746_));
  INVX1    g02553(.A(new_n2746_), .Y(new_n2747_));
  AND2X1   g02554(.A(new_n2745_), .B(new_n2510_), .Y(new_n2748_));
  OAI21X1  g02555(.A0(new_n2622_), .A1(new_n2748_), .B0(new_n2747_), .Y(new_n2749_));
  NOR2X1   g02556(.A(new_n2742_), .B(new_n2625_), .Y(new_n2750_));
  INVX1    g02557(.A(new_n2750_), .Y(new_n2751_));
  AOI21X1  g02558(.A0(new_n2751_), .A1(new_n2744_), .B0(new_n2749_), .Y(new_n2752_));
  AND2X1   g02559(.A(new_n2751_), .B(new_n2749_), .Y(new_n2753_));
  AOI21X1  g02560(.A0(new_n2753_), .A1(new_n2744_), .B0(new_n2752_), .Y(\asquared[41] ));
  NAND2X1  g02561(.A(new_n2740_), .B(new_n2650_), .Y(new_n2755_));
  OAI21X1  g02562(.A0(new_n2647_), .A1(new_n2649_), .B0(new_n2755_), .Y(new_n2756_));
  AND2X1   g02563(.A(new_n2725_), .B(new_n2723_), .Y(new_n2757_));
  AOI21X1  g02564(.A0(new_n2738_), .A1(new_n2726_), .B0(new_n2757_), .Y(new_n2758_));
  NOR2X1   g02565(.A(new_n2658_), .B(new_n2656_), .Y(new_n2759_));
  AOI21X1  g02566(.A0(new_n2692_), .A1(new_n2659_), .B0(new_n2759_), .Y(new_n2760_));
  XOR2X1   g02567(.A(new_n2710_), .B(new_n2667_), .Y(new_n2761_));
  XOR2X1   g02568(.A(new_n2761_), .B(new_n2703_), .Y(new_n2762_));
  INVX1    g02569(.A(new_n2669_), .Y(new_n2763_));
  OR2X1    g02570(.A(new_n2680_), .B(new_n2763_), .Y(new_n2764_));
  OAI21X1  g02571(.A0(new_n2691_), .A1(new_n2681_), .B0(new_n2764_), .Y(new_n2765_));
  XOR2X1   g02572(.A(new_n2765_), .B(new_n2762_), .Y(new_n2766_));
  INVX1    g02573(.A(new_n2766_), .Y(new_n2767_));
  AOI21X1  g02574(.A0(\a[40] ), .A1(\a[1] ), .B0(\a[21] ), .Y(new_n2768_));
  AOI21X1  g02575(.A0(new_n963_), .A1(\a[40] ), .B0(new_n2768_), .Y(new_n2769_));
  XOR2X1   g02576(.A(new_n2769_), .B(new_n2678_), .Y(new_n2770_));
  XOR2X1   g02577(.A(new_n2770_), .B(new_n2720_), .Y(new_n2771_));
  XOR2X1   g02578(.A(new_n2771_), .B(new_n2767_), .Y(new_n2772_));
  XOR2X1   g02579(.A(new_n2772_), .B(new_n2760_), .Y(new_n2773_));
  XOR2X1   g02580(.A(new_n2773_), .B(new_n2758_), .Y(new_n2774_));
  AND2X1   g02581(.A(new_n2695_), .B(new_n2693_), .Y(new_n2775_));
  AOI21X1  g02582(.A0(new_n2739_), .A1(new_n2696_), .B0(new_n2775_), .Y(new_n2776_));
  XOR2X1   g02583(.A(new_n2776_), .B(new_n2774_), .Y(new_n2777_));
  OAI22X1  g02584(.A0(new_n2557_), .A1(new_n230_), .B0(new_n1684_), .B1(new_n488_), .Y(new_n2778_));
  AND2X1   g02585(.A(\a[35] ), .B(\a[30] ), .Y(new_n2779_));
  AND2X1   g02586(.A(new_n2779_), .B(new_n632_), .Y(new_n2780_));
  NAND4X1  g02587(.A(\a[36] ), .B(\a[35] ), .C(\a[6] ), .D(\a[5] ), .Y(new_n2781_));
  NAND4X1  g02588(.A(\a[36] ), .B(\a[30] ), .C(\a[11] ), .D(\a[5] ), .Y(new_n2782_));
  AOI22X1  g02589(.A0(new_n2782_), .A1(new_n2781_), .B0(new_n2779_), .B1(new_n632_), .Y(new_n2783_));
  NOR2X1   g02590(.A(new_n2783_), .B(new_n2780_), .Y(new_n2784_));
  NOR3X1   g02591(.A(new_n2783_), .B(new_n2583_), .C(new_n255_), .Y(new_n2785_));
  AOI21X1  g02592(.A0(new_n2784_), .A1(new_n2778_), .B0(new_n2785_), .Y(new_n2786_));
  AND2X1   g02593(.A(\a[33] ), .B(\a[8] ), .Y(new_n2787_));
  INVX1    g02594(.A(new_n2787_), .Y(new_n2788_));
  AOI22X1  g02595(.A0(\a[22] ), .A1(\a[19] ), .B0(\a[21] ), .B1(\a[20] ), .Y(new_n2789_));
  NOR4X1   g02596(.A(new_n1086_), .B(new_n1098_), .C(new_n934_), .D(new_n752_), .Y(new_n2790_));
  NOR3X1   g02597(.A(new_n2789_), .B(new_n2790_), .C(new_n2788_), .Y(new_n2791_));
  NOR2X1   g02598(.A(new_n2791_), .B(new_n2790_), .Y(new_n2792_));
  INVX1    g02599(.A(new_n2792_), .Y(new_n2793_));
  OAI22X1  g02600(.A0(new_n2793_), .A1(new_n2789_), .B0(new_n2791_), .B1(new_n2788_), .Y(new_n2794_));
  XOR2X1   g02601(.A(new_n2794_), .B(new_n2786_), .Y(new_n2795_));
  AND2X1   g02602(.A(new_n2735_), .B(new_n2733_), .Y(new_n2796_));
  AOI21X1  g02603(.A0(new_n2736_), .A1(new_n2732_), .B0(new_n2796_), .Y(new_n2797_));
  XOR2X1   g02604(.A(new_n2797_), .B(new_n2795_), .Y(new_n2798_));
  NOR2X1   g02605(.A(new_n2730_), .B(new_n2728_), .Y(new_n2799_));
  AOI21X1  g02606(.A0(new_n2737_), .A1(new_n2731_), .B0(new_n2799_), .Y(new_n2800_));
  XOR2X1   g02607(.A(new_n2800_), .B(new_n2798_), .Y(new_n2801_));
  NOR4X1   g02608(.A(new_n2345_), .B(new_n1803_), .C(new_n453_), .D(new_n340_), .Y(new_n2802_));
  NAND4X1  g02609(.A(\a[37] ), .B(\a[27] ), .C(\a[14] ), .D(\a[4] ), .Y(new_n2803_));
  NAND4X1  g02610(.A(\a[29] ), .B(\a[27] ), .C(\a[14] ), .D(\a[12] ), .Y(new_n2804_));
  AOI21X1  g02611(.A0(new_n2804_), .A1(new_n2803_), .B0(new_n2802_), .Y(new_n2805_));
  OR2X1    g02612(.A(new_n2805_), .B(new_n2802_), .Y(new_n2806_));
  AOI22X1  g02613(.A0(\a[37] ), .A1(\a[4] ), .B0(\a[29] ), .B1(\a[12] ), .Y(new_n2807_));
  NAND2X1  g02614(.A(\a[27] ), .B(\a[14] ), .Y(new_n2808_));
  OAI22X1  g02615(.A0(new_n2808_), .A1(new_n2805_), .B0(new_n2807_), .B1(new_n2806_), .Y(new_n2809_));
  NAND4X1  g02616(.A(\a[25] ), .B(\a[23] ), .C(\a[18] ), .D(\a[16] ), .Y(new_n2810_));
  NAND4X1  g02617(.A(\a[25] ), .B(\a[24] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n2811_));
  AOI22X1  g02618(.A0(new_n2811_), .A1(new_n2810_), .B0(new_n1219_), .B1(new_n796_), .Y(new_n2812_));
  NAND2X1  g02619(.A(\a[25] ), .B(\a[16] ), .Y(new_n2813_));
  NAND4X1  g02620(.A(\a[24] ), .B(\a[23] ), .C(\a[18] ), .D(\a[17] ), .Y(new_n2814_));
  NAND3X1  g02621(.A(new_n2811_), .B(new_n2810_), .C(new_n2814_), .Y(new_n2815_));
  AOI22X1  g02622(.A0(\a[24] ), .A1(\a[17] ), .B0(\a[23] ), .B1(\a[18] ), .Y(new_n2816_));
  OAI22X1  g02623(.A0(new_n2816_), .A1(new_n2815_), .B0(new_n2813_), .B1(new_n2812_), .Y(new_n2817_));
  XOR2X1   g02624(.A(new_n2817_), .B(new_n2809_), .Y(new_n2818_));
  INVX1    g02625(.A(new_n1699_), .Y(new_n2819_));
  AND2X1   g02626(.A(\a[34] ), .B(\a[32] ), .Y(new_n2820_));
  NAND4X1  g02627(.A(\a[32] ), .B(\a[31] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n2821_));
  NAND4X1  g02628(.A(\a[34] ), .B(\a[31] ), .C(\a[10] ), .D(\a[7] ), .Y(new_n2822_));
  AOI22X1  g02629(.A0(new_n2822_), .A1(new_n2821_), .B0(new_n2820_), .B1(new_n596_), .Y(new_n2823_));
  AOI21X1  g02630(.A0(new_n2820_), .A1(new_n596_), .B0(new_n2823_), .Y(new_n2824_));
  INVX1    g02631(.A(new_n2824_), .Y(new_n2825_));
  AOI22X1  g02632(.A0(\a[34] ), .A1(\a[7] ), .B0(\a[32] ), .B1(\a[9] ), .Y(new_n2826_));
  OAI22X1  g02633(.A0(new_n2826_), .A1(new_n2825_), .B0(new_n2823_), .B1(new_n2819_), .Y(new_n2827_));
  INVX1    g02634(.A(new_n2827_), .Y(new_n2828_));
  XOR2X1   g02635(.A(new_n2828_), .B(new_n2818_), .Y(new_n2829_));
  XOR2X1   g02636(.A(new_n2829_), .B(new_n2801_), .Y(new_n2830_));
  NAND2X1  g02637(.A(new_n2640_), .B(new_n2629_), .Y(new_n2831_));
  OAI21X1  g02638(.A0(new_n2642_), .A1(new_n2627_), .B0(new_n2831_), .Y(new_n2832_));
  AND2X1   g02639(.A(new_n2830_), .B(new_n2832_), .Y(new_n2833_));
  INVX1    g02640(.A(new_n2833_), .Y(new_n2834_));
  NAND2X1  g02641(.A(new_n2834_), .B(new_n2830_), .Y(new_n2835_));
  AND2X1   g02642(.A(new_n2605_), .B(new_n2595_), .Y(new_n2836_));
  INVX1    g02643(.A(new_n2655_), .Y(new_n2837_));
  AOI21X1  g02644(.A0(new_n2837_), .A1(new_n2651_), .B0(new_n2836_), .Y(new_n2838_));
  AND2X1   g02645(.A(new_n2588_), .B(new_n2630_), .Y(new_n2839_));
  AOI21X1  g02646(.A0(new_n2631_), .A1(new_n2561_), .B0(new_n2839_), .Y(new_n2840_));
  XOR2X1   g02647(.A(new_n2840_), .B(new_n2838_), .Y(new_n2841_));
  INVX1    g02648(.A(new_n2704_), .Y(new_n2842_));
  OR2X1    g02649(.A(new_n2712_), .B(new_n2842_), .Y(new_n2843_));
  OAI21X1  g02650(.A0(new_n2722_), .A1(new_n2713_), .B0(new_n2843_), .Y(new_n2844_));
  XOR2X1   g02651(.A(new_n2844_), .B(new_n2841_), .Y(new_n2845_));
  AND2X1   g02652(.A(new_n2734_), .B(new_n1148_), .Y(new_n2846_));
  AND2X1   g02653(.A(\a[41] ), .B(\a[39] ), .Y(new_n2847_));
  AOI22X1  g02654(.A0(\a[41] ), .A1(\a[0] ), .B0(\a[39] ), .B1(\a[2] ), .Y(new_n2848_));
  AOI21X1  g02655(.A0(new_n2847_), .A1(new_n197_), .B0(new_n2848_), .Y(new_n2849_));
  XOR2X1   g02656(.A(new_n2849_), .B(new_n2846_), .Y(new_n2850_));
  INVX1    g02657(.A(new_n2850_), .Y(new_n2851_));
  XOR2X1   g02658(.A(new_n2851_), .B(new_n2689_), .Y(new_n2852_));
  AND2X1   g02659(.A(\a[38] ), .B(\a[3] ), .Y(new_n2853_));
  AOI22X1  g02660(.A0(\a[28] ), .A1(\a[13] ), .B0(\a[26] ), .B1(\a[15] ), .Y(new_n2854_));
  INVX1    g02661(.A(new_n2854_), .Y(new_n2855_));
  NAND4X1  g02662(.A(\a[28] ), .B(\a[26] ), .C(\a[15] ), .D(\a[13] ), .Y(new_n2856_));
  NAND3X1  g02663(.A(new_n2855_), .B(new_n2856_), .C(new_n2853_), .Y(new_n2857_));
  AOI22X1  g02664(.A0(new_n2855_), .A1(new_n2853_), .B0(new_n1996_), .B1(new_n639_), .Y(new_n2858_));
  AOI22X1  g02665(.A0(new_n2858_), .A1(new_n2855_), .B0(new_n2857_), .B1(new_n2853_), .Y(new_n2859_));
  XOR2X1   g02666(.A(new_n2859_), .B(new_n2852_), .Y(new_n2860_));
  AND2X1   g02667(.A(new_n2638_), .B(new_n2635_), .Y(new_n2861_));
  AOI21X1  g02668(.A0(new_n2639_), .A1(new_n2632_), .B0(new_n2861_), .Y(new_n2862_));
  XOR2X1   g02669(.A(new_n2862_), .B(new_n2860_), .Y(new_n2863_));
  XOR2X1   g02670(.A(new_n2863_), .B(new_n2845_), .Y(new_n2864_));
  XOR2X1   g02671(.A(new_n2830_), .B(new_n2832_), .Y(new_n2865_));
  AND2X1   g02672(.A(new_n2865_), .B(new_n2864_), .Y(new_n2866_));
  AOI21X1  g02673(.A0(new_n2834_), .A1(new_n2832_), .B0(new_n2864_), .Y(new_n2867_));
  AOI21X1  g02674(.A0(new_n2867_), .A1(new_n2835_), .B0(new_n2866_), .Y(new_n2868_));
  XOR2X1   g02675(.A(new_n2868_), .B(new_n2777_), .Y(new_n2869_));
  NOR2X1   g02676(.A(new_n2869_), .B(new_n2756_), .Y(new_n2870_));
  AND2X1   g02677(.A(new_n2869_), .B(new_n2756_), .Y(new_n2871_));
  OR2X1    g02678(.A(new_n2871_), .B(new_n2870_), .Y(new_n2872_));
  AOI21X1  g02679(.A0(new_n2751_), .A1(new_n2749_), .B0(new_n2743_), .Y(new_n2873_));
  XOR2X1   g02680(.A(new_n2873_), .B(new_n2872_), .Y(\asquared[42] ));
  NAND2X1  g02681(.A(new_n2869_), .B(new_n2756_), .Y(new_n2875_));
  OAI21X1  g02682(.A0(new_n2873_), .A1(new_n2870_), .B0(new_n2875_), .Y(new_n2876_));
  NOR2X1   g02683(.A(new_n2776_), .B(new_n2774_), .Y(new_n2877_));
  AOI21X1  g02684(.A0(new_n2868_), .A1(new_n2777_), .B0(new_n2877_), .Y(new_n2878_));
  OR2X1    g02685(.A(new_n2866_), .B(new_n2833_), .Y(new_n2879_));
  NOR2X1   g02686(.A(new_n2862_), .B(new_n2860_), .Y(new_n2880_));
  AOI21X1  g02687(.A0(new_n2863_), .A1(new_n2845_), .B0(new_n2880_), .Y(new_n2881_));
  NOR2X1   g02688(.A(new_n2710_), .B(new_n2667_), .Y(new_n2882_));
  AOI21X1  g02689(.A0(new_n2761_), .A1(new_n2703_), .B0(new_n2882_), .Y(new_n2883_));
  NOR2X1   g02690(.A(new_n2851_), .B(new_n2689_), .Y(new_n2884_));
  INVX1    g02691(.A(new_n2884_), .Y(new_n2885_));
  INVX1    g02692(.A(new_n2852_), .Y(new_n2886_));
  OAI21X1  g02693(.A0(new_n2859_), .A1(new_n2886_), .B0(new_n2885_), .Y(new_n2887_));
  INVX1    g02694(.A(new_n2887_), .Y(new_n2888_));
  XOR2X1   g02695(.A(new_n2888_), .B(new_n2883_), .Y(new_n2889_));
  AND2X1   g02696(.A(new_n2817_), .B(new_n2809_), .Y(new_n2890_));
  AND2X1   g02697(.A(new_n2827_), .B(new_n2818_), .Y(new_n2891_));
  OR2X1    g02698(.A(new_n2891_), .B(new_n2890_), .Y(new_n2892_));
  XOR2X1   g02699(.A(new_n2892_), .B(new_n2889_), .Y(new_n2893_));
  INVX1    g02700(.A(new_n2893_), .Y(new_n2894_));
  AND2X1   g02701(.A(new_n2737_), .B(new_n2731_), .Y(new_n2895_));
  OAI21X1  g02702(.A0(new_n2895_), .A1(new_n2799_), .B0(new_n2798_), .Y(new_n2896_));
  OAI21X1  g02703(.A0(new_n2829_), .A1(new_n2801_), .B0(new_n2896_), .Y(new_n2897_));
  XOR2X1   g02704(.A(new_n2897_), .B(new_n2894_), .Y(new_n2898_));
  XOR2X1   g02705(.A(new_n2898_), .B(new_n2881_), .Y(new_n2899_));
  XOR2X1   g02706(.A(new_n2899_), .B(new_n2879_), .Y(new_n2900_));
  INVX1    g02707(.A(new_n2758_), .Y(new_n2901_));
  NOR2X1   g02708(.A(new_n2772_), .B(new_n2760_), .Y(new_n2902_));
  AOI21X1  g02709(.A0(new_n2773_), .A1(new_n2901_), .B0(new_n2902_), .Y(new_n2903_));
  NOR2X1   g02710(.A(new_n2840_), .B(new_n2838_), .Y(new_n2904_));
  AOI21X1  g02711(.A0(new_n2844_), .A1(new_n2841_), .B0(new_n2904_), .Y(new_n2905_));
  NOR4X1   g02712(.A(new_n2557_), .B(new_n1704_), .C(new_n488_), .D(new_n532_), .Y(new_n2906_));
  AND2X1   g02713(.A(\a[36] ), .B(\a[31] ), .Y(new_n2907_));
  AOI22X1  g02714(.A0(new_n2907_), .A1(new_n632_), .B0(new_n2682_), .B1(new_n375_), .Y(new_n2908_));
  AND2X1   g02715(.A(\a[36] ), .B(\a[6] ), .Y(new_n2909_));
  OAI21X1  g02716(.A0(new_n2908_), .A1(new_n2906_), .B0(new_n2909_), .Y(new_n2910_));
  INVX1    g02717(.A(new_n2906_), .Y(new_n2911_));
  AND2X1   g02718(.A(new_n2908_), .B(new_n2911_), .Y(new_n2912_));
  INVX1    g02719(.A(new_n2912_), .Y(new_n2913_));
  AOI22X1  g02720(.A0(\a[35] ), .A1(\a[7] ), .B0(\a[31] ), .B1(\a[11] ), .Y(new_n2914_));
  OAI21X1  g02721(.A0(new_n2914_), .A1(new_n2913_), .B0(new_n2910_), .Y(new_n2915_));
  XOR2X1   g02722(.A(new_n2915_), .B(new_n2824_), .Y(new_n2916_));
  AND2X1   g02723(.A(\a[32] ), .B(\a[10] ), .Y(new_n2917_));
  AND2X1   g02724(.A(\a[34] ), .B(\a[33] ), .Y(new_n2918_));
  INVX1    g02725(.A(new_n2918_), .Y(new_n2919_));
  INVX1    g02726(.A(new_n2820_), .Y(new_n2920_));
  OAI22X1  g02727(.A0(new_n2920_), .A1(new_n699_), .B0(new_n2675_), .B1(new_n735_), .Y(new_n2921_));
  OAI21X1  g02728(.A0(new_n2919_), .A1(new_n366_), .B0(new_n2921_), .Y(new_n2922_));
  AOI21X1  g02729(.A0(new_n2918_), .A1(new_n1030_), .B0(new_n2921_), .Y(new_n2923_));
  OAI22X1  g02730(.A0(new_n2028_), .A1(new_n413_), .B0(new_n1851_), .B1(new_n341_), .Y(new_n2924_));
  AOI22X1  g02731(.A0(new_n2924_), .A1(new_n2923_), .B0(new_n2922_), .B1(new_n2917_), .Y(new_n2925_));
  XOR2X1   g02732(.A(new_n2925_), .B(new_n2916_), .Y(new_n2926_));
  XOR2X1   g02733(.A(new_n2926_), .B(new_n2905_), .Y(new_n2927_));
  NOR4X1   g02734(.A(new_n2652_), .B(new_n1263_), .C(new_n571_), .D(new_n223_), .Y(new_n2928_));
  NAND4X1  g02735(.A(\a[40] ), .B(\a[26] ), .C(\a[16] ), .D(\a[2] ), .Y(new_n2929_));
  NAND4X1  g02736(.A(\a[40] ), .B(\a[39] ), .C(\a[3] ), .D(\a[2] ), .Y(new_n2930_));
  AOI21X1  g02737(.A0(new_n2930_), .A1(new_n2929_), .B0(new_n2928_), .Y(new_n2931_));
  OR2X1    g02738(.A(new_n2931_), .B(new_n2928_), .Y(new_n2932_));
  AOI22X1  g02739(.A0(\a[39] ), .A1(\a[3] ), .B0(\a[26] ), .B1(\a[16] ), .Y(new_n2933_));
  NAND2X1  g02740(.A(\a[40] ), .B(\a[2] ), .Y(new_n2934_));
  OAI22X1  g02741(.A0(new_n2934_), .A1(new_n2931_), .B0(new_n2933_), .B1(new_n2932_), .Y(new_n2935_));
  NAND4X1  g02742(.A(\a[25] ), .B(\a[23] ), .C(\a[19] ), .D(\a[17] ), .Y(new_n2936_));
  NAND4X1  g02743(.A(\a[25] ), .B(\a[24] ), .C(\a[18] ), .D(\a[17] ), .Y(new_n2937_));
  AOI22X1  g02744(.A0(new_n2937_), .A1(new_n2936_), .B0(new_n1219_), .B1(new_n855_), .Y(new_n2938_));
  NAND2X1  g02745(.A(\a[25] ), .B(\a[17] ), .Y(new_n2939_));
  AOI22X1  g02746(.A0(\a[24] ), .A1(\a[18] ), .B0(\a[23] ), .B1(\a[19] ), .Y(new_n2940_));
  AOI21X1  g02747(.A0(new_n1219_), .A1(new_n855_), .B0(new_n2938_), .Y(new_n2941_));
  INVX1    g02748(.A(new_n2941_), .Y(new_n2942_));
  OAI22X1  g02749(.A0(new_n2942_), .A1(new_n2940_), .B0(new_n2939_), .B1(new_n2938_), .Y(new_n2943_));
  XOR2X1   g02750(.A(new_n2943_), .B(new_n2935_), .Y(new_n2944_));
  NOR4X1   g02751(.A(new_n2519_), .B(new_n1431_), .C(new_n490_), .D(new_n340_), .Y(new_n2945_));
  NOR4X1   g02752(.A(new_n2519_), .B(new_n1679_), .C(new_n549_), .D(new_n340_), .Y(new_n2946_));
  AOI21X1  g02753(.A0(new_n1671_), .A1(new_n691_), .B0(new_n2946_), .Y(new_n2947_));
  AND2X1   g02754(.A(\a[27] ), .B(\a[15] ), .Y(new_n2948_));
  OAI21X1  g02755(.A0(new_n2947_), .A1(new_n2945_), .B0(new_n2948_), .Y(new_n2949_));
  NOR2X1   g02756(.A(new_n2947_), .B(new_n2945_), .Y(new_n2950_));
  NOR2X1   g02757(.A(new_n2950_), .B(new_n2945_), .Y(new_n2951_));
  INVX1    g02758(.A(new_n2951_), .Y(new_n2952_));
  AOI22X1  g02759(.A0(\a[38] ), .A1(\a[4] ), .B0(\a[28] ), .B1(\a[14] ), .Y(new_n2953_));
  OAI21X1  g02760(.A0(new_n2953_), .A1(new_n2952_), .B0(new_n2949_), .Y(new_n2954_));
  INVX1    g02761(.A(new_n2954_), .Y(new_n2955_));
  XOR2X1   g02762(.A(new_n2955_), .B(new_n2944_), .Y(new_n2956_));
  XOR2X1   g02763(.A(new_n2956_), .B(new_n2927_), .Y(new_n2957_));
  XOR2X1   g02764(.A(new_n2957_), .B(new_n2903_), .Y(new_n2958_));
  NAND3X1  g02765(.A(\a[40] ), .B(\a[21] ), .C(\a[1] ), .Y(new_n2959_));
  AND2X1   g02766(.A(\a[42] ), .B(\a[0] ), .Y(new_n2960_));
  XOR2X1   g02767(.A(new_n2960_), .B(new_n2959_), .Y(new_n2961_));
  AND2X1   g02768(.A(\a[41] ), .B(\a[1] ), .Y(new_n2962_));
  XOR2X1   g02769(.A(new_n2962_), .B(new_n2135_), .Y(new_n2963_));
  XOR2X1   g02770(.A(new_n2963_), .B(new_n2961_), .Y(new_n2964_));
  NOR4X1   g02771(.A(new_n2345_), .B(new_n1684_), .C(new_n453_), .D(new_n255_), .Y(new_n2965_));
  NAND4X1  g02772(.A(\a[30] ), .B(\a[29] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n2966_));
  NAND4X1  g02773(.A(\a[37] ), .B(\a[29] ), .C(\a[13] ), .D(\a[5] ), .Y(new_n2967_));
  AOI21X1  g02774(.A0(new_n2967_), .A1(new_n2966_), .B0(new_n2965_), .Y(new_n2968_));
  NAND2X1  g02775(.A(\a[29] ), .B(\a[13] ), .Y(new_n2969_));
  OR2X1    g02776(.A(new_n2968_), .B(new_n2965_), .Y(new_n2970_));
  AOI22X1  g02777(.A0(\a[37] ), .A1(\a[5] ), .B0(\a[30] ), .B1(\a[12] ), .Y(new_n2971_));
  OAI22X1  g02778(.A0(new_n2971_), .A1(new_n2970_), .B0(new_n2969_), .B1(new_n2968_), .Y(new_n2972_));
  XOR2X1   g02779(.A(new_n2972_), .B(new_n2964_), .Y(new_n2973_));
  NOR3X1   g02780(.A(new_n366_), .B(new_n2219_), .C(new_n1704_), .Y(new_n2974_));
  OAI21X1  g02781(.A0(new_n2676_), .A1(new_n2974_), .B0(new_n2769_), .Y(new_n2975_));
  OAI21X1  g02782(.A0(new_n2770_), .A1(new_n2720_), .B0(new_n2975_), .Y(new_n2976_));
  XOR2X1   g02783(.A(new_n2976_), .B(new_n2973_), .Y(new_n2977_));
  INVX1    g02784(.A(new_n2977_), .Y(new_n2978_));
  AND2X1   g02785(.A(new_n2765_), .B(new_n2762_), .Y(new_n2979_));
  AOI21X1  g02786(.A0(new_n2771_), .A1(new_n2766_), .B0(new_n2979_), .Y(new_n2980_));
  XOR2X1   g02787(.A(new_n2980_), .B(new_n2978_), .Y(new_n2981_));
  INVX1    g02788(.A(new_n2784_), .Y(new_n2982_));
  XOR2X1   g02789(.A(new_n2806_), .B(new_n2793_), .Y(new_n2983_));
  XOR2X1   g02790(.A(new_n2983_), .B(new_n2982_), .Y(new_n2984_));
  INVX1    g02791(.A(new_n2984_), .Y(new_n2985_));
  AND2X1   g02792(.A(new_n2784_), .B(new_n2778_), .Y(new_n2986_));
  OAI21X1  g02793(.A0(new_n2785_), .A1(new_n2986_), .B0(new_n2794_), .Y(new_n2987_));
  OAI21X1  g02794(.A0(new_n2797_), .A1(new_n2795_), .B0(new_n2987_), .Y(new_n2988_));
  XOR2X1   g02795(.A(new_n2988_), .B(new_n2985_), .Y(new_n2989_));
  INVX1    g02796(.A(new_n2858_), .Y(new_n2990_));
  XOR2X1   g02797(.A(new_n2815_), .B(new_n2990_), .Y(new_n2991_));
  AOI22X1  g02798(.A0(new_n2849_), .A1(new_n2846_), .B0(new_n2847_), .B1(new_n197_), .Y(new_n2992_));
  XOR2X1   g02799(.A(new_n2992_), .B(new_n2991_), .Y(new_n2993_));
  XOR2X1   g02800(.A(new_n2993_), .B(new_n2989_), .Y(new_n2994_));
  XOR2X1   g02801(.A(new_n2994_), .B(new_n2981_), .Y(new_n2995_));
  XOR2X1   g02802(.A(new_n2995_), .B(new_n2958_), .Y(new_n2996_));
  XOR2X1   g02803(.A(new_n2996_), .B(new_n2900_), .Y(new_n2997_));
  XOR2X1   g02804(.A(new_n2997_), .B(new_n2878_), .Y(new_n2998_));
  XOR2X1   g02805(.A(new_n2998_), .B(new_n2876_), .Y(\asquared[43] ));
  AND2X1   g02806(.A(new_n2899_), .B(new_n2879_), .Y(new_n3000_));
  INVX1    g02807(.A(new_n2996_), .Y(new_n3001_));
  AOI21X1  g02808(.A0(new_n3001_), .A1(new_n2900_), .B0(new_n3000_), .Y(new_n3002_));
  INVX1    g02809(.A(new_n2903_), .Y(new_n3003_));
  AND2X1   g02810(.A(new_n2957_), .B(new_n3003_), .Y(new_n3004_));
  INVX1    g02811(.A(new_n2995_), .Y(new_n3005_));
  NOR2X1   g02812(.A(new_n3005_), .B(new_n2958_), .Y(new_n3006_));
  NOR2X1   g02813(.A(new_n3006_), .B(new_n3004_), .Y(new_n3007_));
  NAND2X1  g02814(.A(new_n2994_), .B(new_n2981_), .Y(new_n3008_));
  OAI21X1  g02815(.A0(new_n2980_), .A1(new_n2978_), .B0(new_n3008_), .Y(new_n3009_));
  INVX1    g02816(.A(new_n2926_), .Y(new_n3010_));
  OR2X1    g02817(.A(new_n3010_), .B(new_n2905_), .Y(new_n3011_));
  OAI21X1  g02818(.A0(new_n2956_), .A1(new_n2927_), .B0(new_n3011_), .Y(new_n3012_));
  AND2X1   g02819(.A(new_n2943_), .B(new_n2935_), .Y(new_n3013_));
  AND2X1   g02820(.A(new_n2954_), .B(new_n2944_), .Y(new_n3014_));
  OR2X1    g02821(.A(new_n3014_), .B(new_n3013_), .Y(new_n3015_));
  NAND2X1  g02822(.A(new_n2915_), .B(new_n2825_), .Y(new_n3016_));
  OAI21X1  g02823(.A0(new_n2925_), .A1(new_n2916_), .B0(new_n3016_), .Y(new_n3017_));
  AND2X1   g02824(.A(new_n2962_), .B(new_n2134_), .Y(new_n3018_));
  AOI21X1  g02825(.A0(\a[42] ), .A1(\a[1] ), .B0(\a[22] ), .Y(new_n3019_));
  AOI21X1  g02826(.A0(new_n1050_), .A1(\a[42] ), .B0(new_n3019_), .Y(new_n3020_));
  XOR2X1   g02827(.A(new_n3020_), .B(new_n3018_), .Y(new_n3021_));
  INVX1    g02828(.A(new_n3021_), .Y(new_n3022_));
  XOR2X1   g02829(.A(new_n3022_), .B(new_n2923_), .Y(new_n3023_));
  INVX1    g02830(.A(new_n3023_), .Y(new_n3024_));
  OR2X1    g02831(.A(new_n3024_), .B(new_n3017_), .Y(new_n3025_));
  XOR2X1   g02832(.A(new_n3023_), .B(new_n3017_), .Y(new_n3026_));
  AOI21X1  g02833(.A0(new_n3024_), .A1(new_n3017_), .B0(new_n3015_), .Y(new_n3027_));
  AOI22X1  g02834(.A0(new_n3027_), .A1(new_n3025_), .B0(new_n3026_), .B1(new_n3015_), .Y(new_n3028_));
  XOR2X1   g02835(.A(new_n3028_), .B(new_n3012_), .Y(new_n3029_));
  XOR2X1   g02836(.A(new_n3029_), .B(new_n3009_), .Y(new_n3030_));
  XOR2X1   g02837(.A(new_n3030_), .B(new_n3007_), .Y(new_n3031_));
  NAND2X1  g02838(.A(new_n2897_), .B(new_n2893_), .Y(new_n3032_));
  OAI21X1  g02839(.A0(new_n2898_), .A1(new_n2881_), .B0(new_n3032_), .Y(new_n3033_));
  NOR2X1   g02840(.A(new_n2888_), .B(new_n2883_), .Y(new_n3034_));
  AOI21X1  g02841(.A0(new_n2892_), .A1(new_n2889_), .B0(new_n3034_), .Y(new_n3035_));
  INVX1    g02842(.A(\a[40] ), .Y(new_n3036_));
  INVX1    g02843(.A(\a[43] ), .Y(new_n3037_));
  NOR4X1   g02844(.A(new_n3037_), .B(new_n3036_), .C(new_n223_), .D(new_n194_), .Y(new_n3038_));
  NAND4X1  g02845(.A(\a[40] ), .B(\a[39] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n3039_));
  NAND4X1  g02846(.A(\a[43] ), .B(\a[39] ), .C(\a[4] ), .D(\a[0] ), .Y(new_n3040_));
  AOI21X1  g02847(.A0(new_n3040_), .A1(new_n3039_), .B0(new_n3038_), .Y(new_n3041_));
  OR2X1    g02848(.A(new_n3041_), .B(new_n3038_), .Y(new_n3042_));
  AOI22X1  g02849(.A0(\a[43] ), .A1(\a[0] ), .B0(\a[40] ), .B1(\a[3] ), .Y(new_n3043_));
  NAND2X1  g02850(.A(\a[39] ), .B(\a[4] ), .Y(new_n3044_));
  OAI22X1  g02851(.A0(new_n3044_), .A1(new_n3041_), .B0(new_n3043_), .B1(new_n3042_), .Y(new_n3045_));
  AOI22X1  g02852(.A0(new_n1674_), .A1(new_n691_), .B0(new_n1484_), .B1(new_n690_), .Y(new_n3046_));
  AOI21X1  g02853(.A0(new_n1671_), .A1(new_n689_), .B0(new_n3046_), .Y(new_n3047_));
  NAND2X1  g02854(.A(\a[29] ), .B(\a[14] ), .Y(new_n3048_));
  OAI21X1  g02855(.A0(new_n1672_), .A1(new_n1024_), .B0(new_n3046_), .Y(new_n3049_));
  AOI22X1  g02856(.A0(\a[28] ), .A1(\a[15] ), .B0(\a[27] ), .B1(\a[16] ), .Y(new_n3050_));
  OAI22X1  g02857(.A0(new_n3050_), .A1(new_n3049_), .B0(new_n3048_), .B1(new_n3047_), .Y(new_n3051_));
  XOR2X1   g02858(.A(new_n3051_), .B(new_n3045_), .Y(new_n3052_));
  AOI22X1  g02859(.A0(new_n2213_), .A1(new_n1650_), .B0(new_n1770_), .B1(new_n796_), .Y(new_n3053_));
  AOI21X1  g02860(.A0(new_n1532_), .A1(new_n855_), .B0(new_n3053_), .Y(new_n3054_));
  AND2X1   g02861(.A(\a[26] ), .B(\a[17] ), .Y(new_n3055_));
  INVX1    g02862(.A(new_n3055_), .Y(new_n3056_));
  AOI22X1  g02863(.A0(\a[25] ), .A1(\a[18] ), .B0(\a[24] ), .B1(\a[19] ), .Y(new_n3057_));
  AOI21X1  g02864(.A0(new_n1532_), .A1(new_n855_), .B0(new_n3054_), .Y(new_n3058_));
  INVX1    g02865(.A(new_n3058_), .Y(new_n3059_));
  OAI22X1  g02866(.A0(new_n3059_), .A1(new_n3057_), .B0(new_n3056_), .B1(new_n3054_), .Y(new_n3060_));
  INVX1    g02867(.A(new_n3060_), .Y(new_n3061_));
  XOR2X1   g02868(.A(new_n3061_), .B(new_n3052_), .Y(new_n3062_));
  NAND4X1  g02869(.A(\a[36] ), .B(\a[35] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n3063_));
  NAND4X1  g02870(.A(\a[36] ), .B(\a[33] ), .C(\a[10] ), .D(\a[7] ), .Y(new_n3064_));
  AOI22X1  g02871(.A0(new_n3064_), .A1(new_n3063_), .B0(new_n2120_), .B1(new_n324_), .Y(new_n3065_));
  AOI21X1  g02872(.A0(new_n2120_), .A1(new_n324_), .B0(new_n3065_), .Y(new_n3066_));
  OAI22X1  g02873(.A0(new_n2557_), .A1(new_n413_), .B0(new_n1851_), .B1(new_n570_), .Y(new_n3067_));
  NOR3X1   g02874(.A(new_n3065_), .B(new_n2583_), .C(new_n532_), .Y(new_n3068_));
  AOI21X1  g02875(.A0(new_n3067_), .A1(new_n3066_), .B0(new_n3068_), .Y(new_n3069_));
  AND2X1   g02876(.A(\a[34] ), .B(\a[9] ), .Y(new_n3070_));
  INVX1    g02877(.A(new_n3070_), .Y(new_n3071_));
  AOI22X1  g02878(.A0(\a[23] ), .A1(\a[20] ), .B0(\a[22] ), .B1(\a[21] ), .Y(new_n3072_));
  AND2X1   g02879(.A(new_n1394_), .B(new_n1236_), .Y(new_n3073_));
  NOR3X1   g02880(.A(new_n3072_), .B(new_n3073_), .C(new_n3071_), .Y(new_n3074_));
  INVX1    g02881(.A(new_n3072_), .Y(new_n3075_));
  AOI21X1  g02882(.A0(new_n3075_), .A1(new_n3070_), .B0(new_n3073_), .Y(new_n3076_));
  INVX1    g02883(.A(new_n3076_), .Y(new_n3077_));
  OAI22X1  g02884(.A0(new_n3077_), .A1(new_n3072_), .B0(new_n3074_), .B1(new_n3071_), .Y(new_n3078_));
  XOR2X1   g02885(.A(new_n3078_), .B(new_n3069_), .Y(new_n3079_));
  AND2X1   g02886(.A(\a[41] ), .B(\a[2] ), .Y(new_n3080_));
  INVX1    g02887(.A(\a[41] ), .Y(new_n3081_));
  NOR4X1   g02888(.A(new_n2519_), .B(new_n1684_), .C(new_n591_), .D(new_n255_), .Y(new_n3082_));
  AOI22X1  g02889(.A0(\a[38] ), .A1(\a[5] ), .B0(\a[30] ), .B1(\a[13] ), .Y(new_n3083_));
  OR4X1    g02890(.A(new_n3083_), .B(new_n3082_), .C(new_n3081_), .D(new_n200_), .Y(new_n3084_));
  NOR3X1   g02891(.A(new_n3083_), .B(new_n3082_), .C(new_n3080_), .Y(new_n3085_));
  AOI21X1  g02892(.A0(new_n3084_), .A1(new_n3080_), .B0(new_n3085_), .Y(new_n3086_));
  XOR2X1   g02893(.A(new_n3086_), .B(new_n3079_), .Y(new_n3087_));
  XOR2X1   g02894(.A(new_n3087_), .B(new_n3062_), .Y(new_n3088_));
  XOR2X1   g02895(.A(new_n3088_), .B(new_n3035_), .Y(new_n3089_));
  XOR2X1   g02896(.A(new_n3089_), .B(new_n3033_), .Y(new_n3090_));
  AND2X1   g02897(.A(new_n2972_), .B(new_n2964_), .Y(new_n3091_));
  AOI21X1  g02898(.A0(new_n2976_), .A1(new_n2973_), .B0(new_n3091_), .Y(new_n3092_));
  XOR2X1   g02899(.A(new_n2951_), .B(new_n2912_), .Y(new_n3093_));
  XOR2X1   g02900(.A(new_n3093_), .B(new_n2941_), .Y(new_n3094_));
  XOR2X1   g02901(.A(new_n2970_), .B(new_n2932_), .Y(new_n3095_));
  INVX1    g02902(.A(\a[42] ), .Y(new_n3096_));
  NOR3X1   g02903(.A(new_n2959_), .B(new_n3096_), .C(new_n194_), .Y(new_n3097_));
  NOR2X1   g02904(.A(new_n2963_), .B(new_n2961_), .Y(new_n3098_));
  NOR2X1   g02905(.A(new_n3098_), .B(new_n3097_), .Y(new_n3099_));
  INVX1    g02906(.A(new_n3099_), .Y(new_n3100_));
  XOR2X1   g02907(.A(new_n3100_), .B(new_n3095_), .Y(new_n3101_));
  INVX1    g02908(.A(new_n3101_), .Y(new_n3102_));
  XOR2X1   g02909(.A(new_n3102_), .B(new_n3094_), .Y(new_n3103_));
  XOR2X1   g02910(.A(new_n3103_), .B(new_n3092_), .Y(new_n3104_));
  AND2X1   g02911(.A(new_n2806_), .B(new_n2793_), .Y(new_n3105_));
  AOI21X1  g02912(.A0(new_n2983_), .A1(new_n2982_), .B0(new_n3105_), .Y(new_n3106_));
  NOR4X1   g02913(.A(new_n2345_), .B(new_n1704_), .C(new_n453_), .D(new_n230_), .Y(new_n3107_));
  AOI21X1  g02914(.A0(new_n2671_), .A1(new_n482_), .B0(new_n3107_), .Y(new_n3108_));
  NAND2X1  g02915(.A(\a[37] ), .B(\a[6] ), .Y(new_n3109_));
  NOR3X1   g02916(.A(new_n3109_), .B(new_n2219_), .C(new_n488_), .Y(new_n3110_));
  AND2X1   g02917(.A(\a[31] ), .B(\a[12] ), .Y(new_n3111_));
  OAI21X1  g02918(.A0(new_n3110_), .A1(new_n3108_), .B0(new_n3111_), .Y(new_n3112_));
  AND2X1   g02919(.A(new_n2671_), .B(new_n482_), .Y(new_n3113_));
  NOR3X1   g02920(.A(new_n3110_), .B(new_n3107_), .C(new_n3113_), .Y(new_n3114_));
  INVX1    g02921(.A(new_n3114_), .Y(new_n3115_));
  AOI22X1  g02922(.A0(\a[37] ), .A1(\a[6] ), .B0(\a[32] ), .B1(\a[11] ), .Y(new_n3116_));
  OAI21X1  g02923(.A0(new_n3116_), .A1(new_n3115_), .B0(new_n3112_), .Y(new_n3117_));
  XOR2X1   g02924(.A(new_n3117_), .B(new_n3106_), .Y(new_n3118_));
  AND2X1   g02925(.A(new_n2815_), .B(new_n2990_), .Y(new_n3119_));
  INVX1    g02926(.A(new_n2992_), .Y(new_n3120_));
  AOI21X1  g02927(.A0(new_n3120_), .A1(new_n2991_), .B0(new_n3119_), .Y(new_n3121_));
  XOR2X1   g02928(.A(new_n3121_), .B(new_n3118_), .Y(new_n3122_));
  NOR2X1   g02929(.A(new_n2993_), .B(new_n2989_), .Y(new_n3123_));
  AOI21X1  g02930(.A0(new_n2988_), .A1(new_n2984_), .B0(new_n3123_), .Y(new_n3124_));
  XOR2X1   g02931(.A(new_n3124_), .B(new_n3122_), .Y(new_n3125_));
  XOR2X1   g02932(.A(new_n3125_), .B(new_n3104_), .Y(new_n3126_));
  XOR2X1   g02933(.A(new_n3126_), .B(new_n3090_), .Y(new_n3127_));
  INVX1    g02934(.A(new_n3127_), .Y(new_n3128_));
  NOR2X1   g02935(.A(new_n3128_), .B(new_n3031_), .Y(new_n3129_));
  OAI21X1  g02936(.A0(new_n3006_), .A1(new_n3004_), .B0(new_n3030_), .Y(new_n3130_));
  OAI21X1  g02937(.A0(new_n3030_), .A1(new_n3007_), .B0(new_n3128_), .Y(new_n3131_));
  AOI21X1  g02938(.A0(new_n3130_), .A1(new_n3030_), .B0(new_n3131_), .Y(new_n3132_));
  NOR2X1   g02939(.A(new_n3132_), .B(new_n3129_), .Y(new_n3133_));
  XOR2X1   g02940(.A(new_n3133_), .B(new_n3002_), .Y(new_n3134_));
  NOR2X1   g02941(.A(new_n2997_), .B(new_n2878_), .Y(new_n3135_));
  AND2X1   g02942(.A(new_n2997_), .B(new_n2878_), .Y(new_n3136_));
  INVX1    g02943(.A(new_n3136_), .Y(new_n3137_));
  AOI21X1  g02944(.A0(new_n3137_), .A1(new_n2876_), .B0(new_n3135_), .Y(new_n3138_));
  XOR2X1   g02945(.A(new_n3138_), .B(new_n3134_), .Y(\asquared[44] ));
  OAI21X1  g02946(.A0(new_n3128_), .A1(new_n3031_), .B0(new_n3130_), .Y(new_n3140_));
  AND2X1   g02947(.A(new_n3028_), .B(new_n3012_), .Y(new_n3141_));
  AOI21X1  g02948(.A0(new_n3029_), .A1(new_n3009_), .B0(new_n3141_), .Y(new_n3142_));
  AND2X1   g02949(.A(new_n3023_), .B(new_n3017_), .Y(new_n3143_));
  AOI21X1  g02950(.A0(new_n3026_), .A1(new_n3015_), .B0(new_n3143_), .Y(new_n3144_));
  AOI22X1  g02951(.A0(\a[29] ), .A1(\a[15] ), .B0(\a[27] ), .B1(\a[17] ), .Y(new_n3145_));
  AND2X1   g02952(.A(\a[41] ), .B(\a[3] ), .Y(new_n3146_));
  INVX1    g02953(.A(new_n3146_), .Y(new_n3147_));
  AND2X1   g02954(.A(new_n1484_), .B(new_n753_), .Y(new_n3148_));
  NOR3X1   g02955(.A(new_n3147_), .B(new_n3148_), .C(new_n3145_), .Y(new_n3149_));
  NOR2X1   g02956(.A(new_n3149_), .B(new_n3148_), .Y(new_n3150_));
  INVX1    g02957(.A(new_n3150_), .Y(new_n3151_));
  OAI22X1  g02958(.A0(new_n3151_), .A1(new_n3145_), .B0(new_n3149_), .B1(new_n3147_), .Y(new_n3152_));
  AND2X1   g02959(.A(\a[26] ), .B(\a[18] ), .Y(new_n3153_));
  OAI22X1  g02960(.A0(new_n1771_), .A1(new_n1518_), .B0(new_n1651_), .B1(new_n1520_), .Y(new_n3154_));
  OAI21X1  g02961(.A0(new_n1772_), .A1(new_n1521_), .B0(new_n3154_), .Y(new_n3155_));
  OAI22X1  g02962(.A0(new_n1326_), .A1(new_n752_), .B0(new_n1185_), .B1(new_n934_), .Y(new_n3156_));
  AOI21X1  g02963(.A0(new_n1532_), .A1(new_n1099_), .B0(new_n3154_), .Y(new_n3157_));
  AOI22X1  g02964(.A0(new_n3157_), .A1(new_n3156_), .B0(new_n3155_), .B1(new_n3153_), .Y(new_n3158_));
  XOR2X1   g02965(.A(new_n3158_), .B(new_n3152_), .Y(new_n3159_));
  AND2X1   g02966(.A(\a[38] ), .B(\a[6] ), .Y(new_n3160_));
  AND2X1   g02967(.A(\a[37] ), .B(\a[11] ), .Y(new_n3161_));
  AND2X1   g02968(.A(new_n3161_), .B(new_n2670_), .Y(new_n3162_));
  AND2X1   g02969(.A(\a[38] ), .B(\a[33] ), .Y(new_n3163_));
  AND2X1   g02970(.A(\a[38] ), .B(\a[37] ), .Y(new_n3164_));
  AOI22X1  g02971(.A0(new_n3164_), .A1(new_n375_), .B0(new_n3163_), .B1(new_n632_), .Y(new_n3165_));
  OR2X1    g02972(.A(new_n3165_), .B(new_n3162_), .Y(new_n3166_));
  INVX1    g02973(.A(new_n3162_), .Y(new_n3167_));
  AND2X1   g02974(.A(new_n3165_), .B(new_n3167_), .Y(new_n3168_));
  OAI22X1  g02975(.A0(new_n2345_), .A1(new_n532_), .B0(new_n1851_), .B1(new_n488_), .Y(new_n3169_));
  AOI22X1  g02976(.A0(new_n3169_), .A1(new_n3168_), .B0(new_n3166_), .B1(new_n3160_), .Y(new_n3170_));
  XOR2X1   g02977(.A(new_n3170_), .B(new_n3159_), .Y(new_n3171_));
  INVX1    g02978(.A(new_n3171_), .Y(new_n3172_));
  NOR4X1   g02979(.A(new_n3036_), .B(new_n1684_), .C(new_n490_), .D(new_n340_), .Y(new_n3173_));
  NAND4X1  g02980(.A(\a[40] ), .B(\a[28] ), .C(\a[16] ), .D(\a[4] ), .Y(new_n3174_));
  NAND4X1  g02981(.A(\a[30] ), .B(\a[28] ), .C(\a[16] ), .D(\a[14] ), .Y(new_n3175_));
  AOI21X1  g02982(.A0(new_n3175_), .A1(new_n3174_), .B0(new_n3173_), .Y(new_n3176_));
  OR2X1    g02983(.A(new_n3176_), .B(new_n3173_), .Y(new_n3177_));
  AOI22X1  g02984(.A0(\a[40] ), .A1(\a[4] ), .B0(\a[30] ), .B1(\a[14] ), .Y(new_n3178_));
  NAND2X1  g02985(.A(\a[28] ), .B(\a[16] ), .Y(new_n3179_));
  OAI22X1  g02986(.A0(new_n3179_), .A1(new_n3176_), .B0(new_n3178_), .B1(new_n3177_), .Y(new_n3180_));
  NAND2X1  g02987(.A(\a[36] ), .B(\a[8] ), .Y(new_n3181_));
  NAND4X1  g02988(.A(\a[36] ), .B(\a[34] ), .C(\a[10] ), .D(\a[8] ), .Y(new_n3182_));
  NAND4X1  g02989(.A(\a[36] ), .B(\a[35] ), .C(\a[9] ), .D(\a[8] ), .Y(new_n3183_));
  AOI22X1  g02990(.A0(new_n3183_), .A1(new_n3182_), .B0(new_n2361_), .B1(new_n881_), .Y(new_n3184_));
  AOI21X1  g02991(.A0(new_n2361_), .A1(new_n881_), .B0(new_n3184_), .Y(new_n3185_));
  INVX1    g02992(.A(new_n3185_), .Y(new_n3186_));
  AOI22X1  g02993(.A0(\a[35] ), .A1(\a[9] ), .B0(\a[34] ), .B1(\a[10] ), .Y(new_n3187_));
  OAI22X1  g02994(.A0(new_n3187_), .A1(new_n3186_), .B0(new_n3184_), .B1(new_n3181_), .Y(new_n3188_));
  XOR2X1   g02995(.A(new_n3188_), .B(new_n3180_), .Y(new_n3189_));
  AND2X1   g02996(.A(\a[39] ), .B(\a[5] ), .Y(new_n3190_));
  INVX1    g02997(.A(new_n3190_), .Y(new_n3191_));
  AOI22X1  g02998(.A0(\a[32] ), .A1(\a[12] ), .B0(\a[31] ), .B1(\a[13] ), .Y(new_n3192_));
  AND2X1   g02999(.A(new_n2671_), .B(new_n586_), .Y(new_n3193_));
  NOR3X1   g03000(.A(new_n3192_), .B(new_n3193_), .C(new_n3191_), .Y(new_n3194_));
  NOR2X1   g03001(.A(new_n3194_), .B(new_n3193_), .Y(new_n3195_));
  INVX1    g03002(.A(new_n3195_), .Y(new_n3196_));
  OAI22X1  g03003(.A0(new_n3196_), .A1(new_n3192_), .B0(new_n3194_), .B1(new_n3191_), .Y(new_n3197_));
  INVX1    g03004(.A(new_n3197_), .Y(new_n3198_));
  XOR2X1   g03005(.A(new_n3198_), .B(new_n3189_), .Y(new_n3199_));
  XOR2X1   g03006(.A(new_n3199_), .B(new_n3172_), .Y(new_n3200_));
  INVX1    g03007(.A(new_n3200_), .Y(new_n3201_));
  XOR2X1   g03008(.A(new_n3201_), .B(new_n3144_), .Y(new_n3202_));
  INVX1    g03009(.A(new_n3202_), .Y(new_n3203_));
  XOR2X1   g03010(.A(new_n3203_), .B(new_n3142_), .Y(new_n3204_));
  XOR2X1   g03011(.A(new_n3115_), .B(new_n3049_), .Y(new_n3205_));
  AOI22X1  g03012(.A0(\a[44] ), .A1(\a[0] ), .B0(\a[42] ), .B1(\a[2] ), .Y(new_n3206_));
  AND2X1   g03013(.A(new_n1050_), .B(\a[42] ), .Y(new_n3207_));
  AND2X1   g03014(.A(\a[44] ), .B(\a[42] ), .Y(new_n3208_));
  AND2X1   g03015(.A(new_n3208_), .B(new_n197_), .Y(new_n3209_));
  OAI21X1  g03016(.A0(new_n3209_), .A1(new_n3206_), .B0(new_n3207_), .Y(new_n3210_));
  INVX1    g03017(.A(new_n3207_), .Y(new_n3211_));
  INVX1    g03018(.A(new_n3208_), .Y(new_n3212_));
  OAI22X1  g03019(.A0(new_n3212_), .A1(new_n198_), .B0(new_n3206_), .B1(new_n3211_), .Y(new_n3213_));
  OAI21X1  g03020(.A0(new_n3213_), .A1(new_n3206_), .B0(new_n3210_), .Y(new_n3214_));
  XOR2X1   g03021(.A(new_n3214_), .B(new_n3205_), .Y(new_n3215_));
  AND2X1   g03022(.A(\a[43] ), .B(\a[1] ), .Y(new_n3216_));
  XOR2X1   g03023(.A(new_n3216_), .B(new_n1016_), .Y(new_n3217_));
  XOR2X1   g03024(.A(new_n3217_), .B(new_n3076_), .Y(new_n3218_));
  XOR2X1   g03025(.A(new_n3218_), .B(new_n3066_), .Y(new_n3219_));
  XOR2X1   g03026(.A(new_n3219_), .B(new_n3215_), .Y(new_n3220_));
  INVX1    g03027(.A(new_n3117_), .Y(new_n3221_));
  OR2X1    g03028(.A(new_n3221_), .B(new_n3106_), .Y(new_n3222_));
  OAI21X1  g03029(.A0(new_n3121_), .A1(new_n3118_), .B0(new_n3222_), .Y(new_n3223_));
  XOR2X1   g03030(.A(new_n3223_), .B(new_n3220_), .Y(new_n3224_));
  AND2X1   g03031(.A(new_n3102_), .B(new_n3094_), .Y(new_n3225_));
  OR2X1    g03032(.A(new_n3102_), .B(new_n3094_), .Y(new_n3226_));
  OAI21X1  g03033(.A0(new_n3225_), .A1(new_n3092_), .B0(new_n3226_), .Y(new_n3227_));
  AND2X1   g03034(.A(new_n2970_), .B(new_n2932_), .Y(new_n3228_));
  AOI21X1  g03035(.A0(new_n3100_), .A1(new_n3095_), .B0(new_n3228_), .Y(new_n3229_));
  AND2X1   g03036(.A(new_n3020_), .B(new_n3018_), .Y(new_n3230_));
  NOR2X1   g03037(.A(new_n3022_), .B(new_n2923_), .Y(new_n3231_));
  NOR2X1   g03038(.A(new_n3231_), .B(new_n3230_), .Y(new_n3232_));
  INVX1    g03039(.A(new_n3232_), .Y(new_n3233_));
  XOR2X1   g03040(.A(new_n3233_), .B(new_n3229_), .Y(new_n3234_));
  NOR2X1   g03041(.A(new_n2951_), .B(new_n2912_), .Y(new_n3235_));
  AOI21X1  g03042(.A0(new_n3093_), .A1(new_n2942_), .B0(new_n3235_), .Y(new_n3236_));
  XOR2X1   g03043(.A(new_n3236_), .B(new_n3234_), .Y(new_n3237_));
  XOR2X1   g03044(.A(new_n3237_), .B(new_n3227_), .Y(new_n3238_));
  XOR2X1   g03045(.A(new_n3238_), .B(new_n3224_), .Y(new_n3239_));
  XOR2X1   g03046(.A(new_n3239_), .B(new_n3204_), .Y(new_n3240_));
  AND2X1   g03047(.A(new_n3089_), .B(new_n3033_), .Y(new_n3241_));
  AOI21X1  g03048(.A0(new_n3126_), .A1(new_n3090_), .B0(new_n3241_), .Y(new_n3242_));
  INVX1    g03049(.A(new_n3124_), .Y(new_n3243_));
  NOR2X1   g03050(.A(new_n3125_), .B(new_n3104_), .Y(new_n3244_));
  AOI21X1  g03051(.A0(new_n3243_), .A1(new_n3122_), .B0(new_n3244_), .Y(new_n3245_));
  XOR2X1   g03052(.A(new_n3060_), .B(new_n3052_), .Y(new_n3246_));
  NAND2X1  g03053(.A(new_n3087_), .B(new_n3246_), .Y(new_n3247_));
  OAI21X1  g03054(.A0(new_n3088_), .A1(new_n3035_), .B0(new_n3247_), .Y(new_n3248_));
  NOR3X1   g03055(.A(new_n3083_), .B(new_n3081_), .C(new_n200_), .Y(new_n3249_));
  NOR2X1   g03056(.A(new_n3249_), .B(new_n3082_), .Y(new_n3250_));
  INVX1    g03057(.A(new_n3250_), .Y(new_n3251_));
  XOR2X1   g03058(.A(new_n3251_), .B(new_n3042_), .Y(new_n3252_));
  XOR2X1   g03059(.A(new_n3252_), .B(new_n3059_), .Y(new_n3253_));
  AND2X1   g03060(.A(new_n3067_), .B(new_n3066_), .Y(new_n3254_));
  OAI21X1  g03061(.A0(new_n3068_), .A1(new_n3254_), .B0(new_n3078_), .Y(new_n3255_));
  OAI21X1  g03062(.A0(new_n3086_), .A1(new_n3079_), .B0(new_n3255_), .Y(new_n3256_));
  AND2X1   g03063(.A(new_n3051_), .B(new_n3045_), .Y(new_n3257_));
  AND2X1   g03064(.A(new_n3060_), .B(new_n3052_), .Y(new_n3258_));
  OR2X1    g03065(.A(new_n3258_), .B(new_n3257_), .Y(new_n3259_));
  XOR2X1   g03066(.A(new_n3259_), .B(new_n3256_), .Y(new_n3260_));
  XOR2X1   g03067(.A(new_n3260_), .B(new_n3253_), .Y(new_n3261_));
  XOR2X1   g03068(.A(new_n3261_), .B(new_n3248_), .Y(new_n3262_));
  XOR2X1   g03069(.A(new_n3262_), .B(new_n3245_), .Y(new_n3263_));
  XOR2X1   g03070(.A(new_n3263_), .B(new_n3242_), .Y(new_n3264_));
  XOR2X1   g03071(.A(new_n3264_), .B(new_n3240_), .Y(new_n3265_));
  XOR2X1   g03072(.A(new_n3265_), .B(new_n3140_), .Y(new_n3266_));
  INVX1    g03073(.A(new_n3002_), .Y(new_n3267_));
  NAND2X1  g03074(.A(new_n3133_), .B(new_n3267_), .Y(new_n3268_));
  NOR2X1   g03075(.A(new_n3133_), .B(new_n3267_), .Y(new_n3269_));
  OAI21X1  g03076(.A0(new_n3138_), .A1(new_n3269_), .B0(new_n3268_), .Y(new_n3270_));
  XOR2X1   g03077(.A(new_n3270_), .B(new_n3266_), .Y(\asquared[45] ));
  OR2X1    g03078(.A(new_n3199_), .B(new_n3172_), .Y(new_n3272_));
  OAI21X1  g03079(.A0(new_n3201_), .A1(new_n3144_), .B0(new_n3272_), .Y(new_n3273_));
  AND2X1   g03080(.A(new_n3237_), .B(new_n3227_), .Y(new_n3274_));
  AOI21X1  g03081(.A0(new_n3238_), .A1(new_n3224_), .B0(new_n3274_), .Y(new_n3275_));
  XOR2X1   g03082(.A(new_n3275_), .B(new_n3273_), .Y(new_n3276_));
  INVX1    g03083(.A(new_n3157_), .Y(new_n3277_));
  XOR2X1   g03084(.A(new_n3213_), .B(new_n3151_), .Y(new_n3278_));
  XOR2X1   g03085(.A(new_n3278_), .B(new_n3277_), .Y(new_n3279_));
  INVX1    g03086(.A(new_n3279_), .Y(new_n3280_));
  OR2X1    g03087(.A(new_n3232_), .B(new_n3229_), .Y(new_n3281_));
  OAI21X1  g03088(.A0(new_n3236_), .A1(new_n3234_), .B0(new_n3281_), .Y(new_n3282_));
  XOR2X1   g03089(.A(new_n3282_), .B(new_n3280_), .Y(new_n3283_));
  AOI22X1  g03090(.A0(\a[39] ), .A1(\a[6] ), .B0(\a[34] ), .B1(\a[11] ), .Y(new_n3284_));
  AND2X1   g03091(.A(\a[39] ), .B(\a[34] ), .Y(new_n3285_));
  NAND4X1  g03092(.A(\a[39] ), .B(\a[33] ), .C(\a[12] ), .D(\a[6] ), .Y(new_n3286_));
  NAND4X1  g03093(.A(\a[34] ), .B(\a[33] ), .C(\a[12] ), .D(\a[11] ), .Y(new_n3287_));
  AOI22X1  g03094(.A0(new_n3287_), .A1(new_n3286_), .B0(new_n3285_), .B1(new_n632_), .Y(new_n3288_));
  AOI21X1  g03095(.A0(new_n3285_), .A1(new_n632_), .B0(new_n3288_), .Y(new_n3289_));
  INVX1    g03096(.A(new_n3289_), .Y(new_n3290_));
  NAND2X1  g03097(.A(\a[33] ), .B(\a[12] ), .Y(new_n3291_));
  OAI22X1  g03098(.A0(new_n3291_), .A1(new_n3288_), .B0(new_n3290_), .B1(new_n3284_), .Y(new_n3292_));
  NAND4X1  g03099(.A(\a[30] ), .B(\a[28] ), .C(\a[17] ), .D(\a[15] ), .Y(new_n3293_));
  NAND4X1  g03100(.A(\a[30] ), .B(\a[29] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n3294_));
  AOI22X1  g03101(.A0(new_n3294_), .A1(new_n3293_), .B0(new_n1674_), .B1(new_n792_), .Y(new_n3295_));
  NAND2X1  g03102(.A(\a[30] ), .B(\a[15] ), .Y(new_n3296_));
  NAND4X1  g03103(.A(\a[29] ), .B(\a[28] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n3297_));
  NAND3X1  g03104(.A(new_n3294_), .B(new_n3293_), .C(new_n3297_), .Y(new_n3298_));
  AOI22X1  g03105(.A0(\a[29] ), .A1(\a[16] ), .B0(\a[28] ), .B1(\a[17] ), .Y(new_n3299_));
  OAI22X1  g03106(.A0(new_n3299_), .A1(new_n3298_), .B0(new_n3296_), .B1(new_n3295_), .Y(new_n3300_));
  XOR2X1   g03107(.A(new_n3300_), .B(new_n3292_), .Y(new_n3301_));
  AND2X1   g03108(.A(new_n1082_), .B(\a[44] ), .Y(new_n3302_));
  INVX1    g03109(.A(new_n3302_), .Y(new_n3303_));
  AND2X1   g03110(.A(\a[44] ), .B(\a[1] ), .Y(new_n3304_));
  OAI21X1  g03111(.A0(new_n3304_), .A1(\a[23] ), .B0(new_n3303_), .Y(new_n3305_));
  AOI22X1  g03112(.A0(new_n3216_), .A1(new_n1016_), .B0(\a[42] ), .B1(\a[3] ), .Y(new_n3306_));
  NAND4X1  g03113(.A(new_n3216_), .B(new_n1016_), .C(\a[42] ), .D(\a[3] ), .Y(new_n3307_));
  INVX1    g03114(.A(new_n3307_), .Y(new_n3308_));
  NOR3X1   g03115(.A(new_n3308_), .B(new_n3306_), .C(new_n3305_), .Y(new_n3309_));
  NOR2X1   g03116(.A(new_n3309_), .B(new_n3308_), .Y(new_n3310_));
  INVX1    g03117(.A(new_n3310_), .Y(new_n3311_));
  OAI22X1  g03118(.A0(new_n3311_), .A1(new_n3306_), .B0(new_n3309_), .B1(new_n3305_), .Y(new_n3312_));
  INVX1    g03119(.A(new_n3312_), .Y(new_n3313_));
  XOR2X1   g03120(.A(new_n3313_), .B(new_n3301_), .Y(new_n3314_));
  XOR2X1   g03121(.A(new_n3314_), .B(new_n3283_), .Y(new_n3315_));
  XOR2X1   g03122(.A(new_n3315_), .B(new_n3276_), .Y(new_n3316_));
  NOR2X1   g03123(.A(new_n3203_), .B(new_n3142_), .Y(new_n3317_));
  AOI21X1  g03124(.A0(new_n3239_), .A1(new_n3204_), .B0(new_n3317_), .Y(new_n3318_));
  XOR2X1   g03125(.A(new_n3318_), .B(new_n3316_), .Y(new_n3319_));
  AND2X1   g03126(.A(\a[43] ), .B(\a[41] ), .Y(new_n3320_));
  NAND4X1  g03127(.A(\a[45] ), .B(\a[41] ), .C(\a[4] ), .D(\a[0] ), .Y(new_n3321_));
  NAND4X1  g03128(.A(\a[45] ), .B(\a[43] ), .C(\a[2] ), .D(\a[0] ), .Y(new_n3322_));
  AOI22X1  g03129(.A0(new_n3322_), .A1(new_n3321_), .B0(new_n3320_), .B1(new_n235_), .Y(new_n3323_));
  NAND4X1  g03130(.A(\a[43] ), .B(\a[41] ), .C(\a[4] ), .D(\a[2] ), .Y(new_n3324_));
  NAND3X1  g03131(.A(new_n3322_), .B(new_n3321_), .C(new_n3324_), .Y(new_n3325_));
  AOI22X1  g03132(.A0(\a[43] ), .A1(\a[2] ), .B0(\a[41] ), .B1(\a[4] ), .Y(new_n3326_));
  NAND2X1  g03133(.A(\a[45] ), .B(\a[0] ), .Y(new_n3327_));
  OAI22X1  g03134(.A0(new_n3327_), .A1(new_n3323_), .B0(new_n3326_), .B1(new_n3325_), .Y(new_n3328_));
  NAND2X1  g03135(.A(\a[38] ), .B(\a[7] ), .Y(new_n3329_));
  AND2X1   g03136(.A(\a[37] ), .B(\a[36] ), .Y(new_n3330_));
  NAND4X1  g03137(.A(\a[38] ), .B(\a[36] ), .C(\a[9] ), .D(\a[7] ), .Y(new_n3331_));
  NAND4X1  g03138(.A(\a[38] ), .B(\a[37] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n3332_));
  AOI22X1  g03139(.A0(new_n3332_), .A1(new_n3331_), .B0(new_n3330_), .B1(new_n1030_), .Y(new_n3333_));
  AOI22X1  g03140(.A0(\a[37] ), .A1(\a[8] ), .B0(\a[36] ), .B1(\a[9] ), .Y(new_n3334_));
  AOI21X1  g03141(.A0(new_n3330_), .A1(new_n1030_), .B0(new_n3333_), .Y(new_n3335_));
  INVX1    g03142(.A(new_n3335_), .Y(new_n3336_));
  OAI22X1  g03143(.A0(new_n3336_), .A1(new_n3334_), .B0(new_n3333_), .B1(new_n3329_), .Y(new_n3337_));
  XOR2X1   g03144(.A(new_n3337_), .B(new_n3328_), .Y(new_n3338_));
  AOI22X1  g03145(.A0(\a[24] ), .A1(\a[21] ), .B0(\a[23] ), .B1(\a[22] ), .Y(new_n3339_));
  AND2X1   g03146(.A(\a[35] ), .B(\a[10] ), .Y(new_n3340_));
  AND2X1   g03147(.A(new_n1219_), .B(new_n1154_), .Y(new_n3341_));
  OAI21X1  g03148(.A0(new_n3339_), .A1(new_n3341_), .B0(new_n3340_), .Y(new_n3342_));
  INVX1    g03149(.A(new_n3339_), .Y(new_n3343_));
  AOI21X1  g03150(.A0(new_n3343_), .A1(new_n3340_), .B0(new_n3341_), .Y(new_n3344_));
  INVX1    g03151(.A(new_n3344_), .Y(new_n3345_));
  OAI21X1  g03152(.A0(new_n3345_), .A1(new_n3339_), .B0(new_n3342_), .Y(new_n3346_));
  XOR2X1   g03153(.A(new_n3346_), .B(new_n3338_), .Y(new_n3347_));
  INVX1    g03154(.A(new_n3347_), .Y(new_n3348_));
  NOR4X1   g03155(.A(new_n3036_), .B(new_n2219_), .C(new_n591_), .D(new_n255_), .Y(new_n3349_));
  AND2X1   g03156(.A(\a[31] ), .B(\a[5] ), .Y(new_n3350_));
  AND2X1   g03157(.A(\a[40] ), .B(\a[14] ), .Y(new_n3351_));
  AOI22X1  g03158(.A0(new_n3351_), .A1(new_n3350_), .B0(new_n2671_), .B1(new_n582_), .Y(new_n3352_));
  OR2X1    g03159(.A(new_n3352_), .B(new_n3349_), .Y(new_n3353_));
  INVX1    g03160(.A(new_n3349_), .Y(new_n3354_));
  AND2X1   g03161(.A(new_n3352_), .B(new_n3354_), .Y(new_n3355_));
  OAI22X1  g03162(.A0(new_n3036_), .A1(new_n255_), .B0(new_n2219_), .B1(new_n591_), .Y(new_n3356_));
  AND2X1   g03163(.A(\a[31] ), .B(\a[14] ), .Y(new_n3357_));
  AOI22X1  g03164(.A0(new_n3357_), .A1(new_n3353_), .B0(new_n3356_), .B1(new_n3355_), .Y(new_n3358_));
  NAND4X1  g03165(.A(\a[27] ), .B(\a[25] ), .C(\a[20] ), .D(\a[18] ), .Y(new_n3359_));
  NAND4X1  g03166(.A(\a[27] ), .B(\a[26] ), .C(\a[19] ), .D(\a[18] ), .Y(new_n3360_));
  AOI22X1  g03167(.A0(new_n3360_), .A1(new_n3359_), .B0(new_n1770_), .B1(new_n1099_), .Y(new_n3361_));
  NAND2X1  g03168(.A(\a[27] ), .B(\a[18] ), .Y(new_n3362_));
  NAND4X1  g03169(.A(\a[26] ), .B(\a[25] ), .C(\a[20] ), .D(\a[19] ), .Y(new_n3363_));
  NAND3X1  g03170(.A(new_n3360_), .B(new_n3359_), .C(new_n3363_), .Y(new_n3364_));
  AOI22X1  g03171(.A0(\a[26] ), .A1(\a[19] ), .B0(\a[25] ), .B1(\a[20] ), .Y(new_n3365_));
  OAI22X1  g03172(.A0(new_n3365_), .A1(new_n3364_), .B0(new_n3362_), .B1(new_n3361_), .Y(new_n3366_));
  XOR2X1   g03173(.A(new_n3366_), .B(new_n3185_), .Y(new_n3367_));
  XOR2X1   g03174(.A(new_n3367_), .B(new_n3358_), .Y(new_n3368_));
  XOR2X1   g03175(.A(new_n3368_), .B(new_n3348_), .Y(new_n3369_));
  AND2X1   g03176(.A(new_n3259_), .B(new_n3256_), .Y(new_n3370_));
  AOI21X1  g03177(.A0(new_n3260_), .A1(new_n3253_), .B0(new_n3370_), .Y(new_n3371_));
  XOR2X1   g03178(.A(new_n3371_), .B(new_n3369_), .Y(new_n3372_));
  NAND2X1  g03179(.A(new_n3261_), .B(new_n3248_), .Y(new_n3373_));
  NOR2X1   g03180(.A(new_n3261_), .B(new_n3248_), .Y(new_n3374_));
  OAI21X1  g03181(.A0(new_n3374_), .A1(new_n3245_), .B0(new_n3373_), .Y(new_n3375_));
  XOR2X1   g03182(.A(new_n3375_), .B(new_n3372_), .Y(new_n3376_));
  NAND2X1  g03183(.A(new_n3115_), .B(new_n3049_), .Y(new_n3377_));
  NAND2X1  g03184(.A(new_n3214_), .B(new_n3205_), .Y(new_n3378_));
  AND2X1   g03185(.A(new_n3378_), .B(new_n3377_), .Y(new_n3379_));
  AND2X1   g03186(.A(new_n3251_), .B(new_n3042_), .Y(new_n3380_));
  AOI21X1  g03187(.A0(new_n3252_), .A1(new_n3059_), .B0(new_n3380_), .Y(new_n3381_));
  XOR2X1   g03188(.A(new_n3381_), .B(new_n3379_), .Y(new_n3382_));
  INVX1    g03189(.A(new_n3382_), .Y(new_n3383_));
  OAI21X1  g03190(.A0(new_n3074_), .A1(new_n3073_), .B0(new_n3217_), .Y(new_n3384_));
  OAI21X1  g03191(.A0(new_n3218_), .A1(new_n3066_), .B0(new_n3384_), .Y(new_n3385_));
  XOR2X1   g03192(.A(new_n3385_), .B(new_n3383_), .Y(new_n3386_));
  AND2X1   g03193(.A(new_n3219_), .B(new_n3215_), .Y(new_n3387_));
  AOI21X1  g03194(.A0(new_n3223_), .A1(new_n3220_), .B0(new_n3387_), .Y(new_n3388_));
  XOR2X1   g03195(.A(new_n3388_), .B(new_n3386_), .Y(new_n3389_));
  INVX1    g03196(.A(new_n3168_), .Y(new_n3390_));
  XOR2X1   g03197(.A(new_n3177_), .B(new_n3390_), .Y(new_n3391_));
  XOR2X1   g03198(.A(new_n3391_), .B(new_n3196_), .Y(new_n3392_));
  AND2X1   g03199(.A(new_n3188_), .B(new_n3180_), .Y(new_n3393_));
  AND2X1   g03200(.A(new_n3197_), .B(new_n3189_), .Y(new_n3394_));
  OR2X1    g03201(.A(new_n3394_), .B(new_n3393_), .Y(new_n3395_));
  INVX1    g03202(.A(new_n3152_), .Y(new_n3396_));
  OR2X1    g03203(.A(new_n3158_), .B(new_n3396_), .Y(new_n3397_));
  OAI21X1  g03204(.A0(new_n3170_), .A1(new_n3159_), .B0(new_n3397_), .Y(new_n3398_));
  XOR2X1   g03205(.A(new_n3398_), .B(new_n3395_), .Y(new_n3399_));
  XOR2X1   g03206(.A(new_n3399_), .B(new_n3392_), .Y(new_n3400_));
  XOR2X1   g03207(.A(new_n3400_), .B(new_n3389_), .Y(new_n3401_));
  XOR2X1   g03208(.A(new_n3401_), .B(new_n3376_), .Y(new_n3402_));
  XOR2X1   g03209(.A(new_n3402_), .B(new_n3319_), .Y(new_n3403_));
  NOR2X1   g03210(.A(new_n3263_), .B(new_n3242_), .Y(new_n3404_));
  AOI21X1  g03211(.A0(new_n3264_), .A1(new_n3240_), .B0(new_n3404_), .Y(new_n3405_));
  XOR2X1   g03212(.A(new_n3405_), .B(new_n3403_), .Y(new_n3406_));
  AND2X1   g03213(.A(new_n3265_), .B(new_n3140_), .Y(new_n3407_));
  NOR2X1   g03214(.A(new_n3265_), .B(new_n3140_), .Y(new_n3408_));
  INVX1    g03215(.A(new_n3408_), .Y(new_n3409_));
  AOI21X1  g03216(.A0(new_n3270_), .A1(new_n3409_), .B0(new_n3407_), .Y(new_n3410_));
  XOR2X1   g03217(.A(new_n3410_), .B(new_n3406_), .Y(\asquared[46] ));
  NOR2X1   g03218(.A(new_n3318_), .B(new_n3316_), .Y(new_n3412_));
  AOI21X1  g03219(.A0(new_n3402_), .A1(new_n3319_), .B0(new_n3412_), .Y(new_n3413_));
  INVX1    g03220(.A(new_n3413_), .Y(new_n3414_));
  AND2X1   g03221(.A(new_n3375_), .B(new_n3372_), .Y(new_n3415_));
  AND2X1   g03222(.A(new_n3401_), .B(new_n3376_), .Y(new_n3416_));
  OR2X1    g03223(.A(new_n3416_), .B(new_n3415_), .Y(new_n3417_));
  NAND2X1  g03224(.A(new_n3400_), .B(new_n3389_), .Y(new_n3418_));
  OAI21X1  g03225(.A0(new_n3388_), .A1(new_n3386_), .B0(new_n3418_), .Y(new_n3419_));
  NAND2X1  g03226(.A(new_n3368_), .B(new_n3347_), .Y(new_n3420_));
  OAI21X1  g03227(.A0(new_n3371_), .A1(new_n3369_), .B0(new_n3420_), .Y(new_n3421_));
  XOR2X1   g03228(.A(new_n3421_), .B(new_n3419_), .Y(new_n3422_));
  AOI22X1  g03229(.A0(\a[41] ), .A1(\a[5] ), .B0(\a[31] ), .B1(\a[15] ), .Y(new_n3423_));
  AND2X1   g03230(.A(\a[44] ), .B(\a[2] ), .Y(new_n3424_));
  INVX1    g03231(.A(new_n3424_), .Y(new_n3425_));
  NOR4X1   g03232(.A(new_n3081_), .B(new_n1704_), .C(new_n549_), .D(new_n255_), .Y(new_n3426_));
  NOR3X1   g03233(.A(new_n3425_), .B(new_n3426_), .C(new_n3423_), .Y(new_n3427_));
  INVX1    g03234(.A(new_n3423_), .Y(new_n3428_));
  AOI21X1  g03235(.A0(new_n3424_), .A1(new_n3428_), .B0(new_n3426_), .Y(new_n3429_));
  INVX1    g03236(.A(new_n3429_), .Y(new_n3430_));
  OAI22X1  g03237(.A0(new_n3430_), .A1(new_n3423_), .B0(new_n3427_), .B1(new_n3425_), .Y(new_n3431_));
  AOI22X1  g03238(.A0(new_n3351_), .A1(new_n2410_), .B0(new_n2674_), .B1(new_n582_), .Y(new_n3432_));
  NOR4X1   g03239(.A(new_n3036_), .B(new_n1851_), .C(new_n591_), .D(new_n230_), .Y(new_n3433_));
  OR2X1    g03240(.A(new_n3433_), .B(new_n3432_), .Y(new_n3434_));
  AND2X1   g03241(.A(\a[32] ), .B(\a[14] ), .Y(new_n3435_));
  INVX1    g03242(.A(new_n3433_), .Y(new_n3436_));
  AND2X1   g03243(.A(new_n3436_), .B(new_n3432_), .Y(new_n3437_));
  OAI22X1  g03244(.A0(new_n3036_), .A1(new_n230_), .B0(new_n1851_), .B1(new_n591_), .Y(new_n3438_));
  AOI22X1  g03245(.A0(new_n3438_), .A1(new_n3437_), .B0(new_n3435_), .B1(new_n3434_), .Y(new_n3439_));
  XOR2X1   g03246(.A(new_n3439_), .B(new_n3431_), .Y(new_n3440_));
  AND2X1   g03247(.A(new_n3177_), .B(new_n3390_), .Y(new_n3441_));
  AOI21X1  g03248(.A0(new_n3391_), .A1(new_n3196_), .B0(new_n3441_), .Y(new_n3442_));
  XOR2X1   g03249(.A(new_n3442_), .B(new_n3440_), .Y(new_n3443_));
  XOR2X1   g03250(.A(new_n3364_), .B(new_n3298_), .Y(new_n3444_));
  XOR2X1   g03251(.A(new_n3444_), .B(new_n3289_), .Y(new_n3445_));
  AOI21X1  g03252(.A0(new_n3378_), .A1(new_n3377_), .B0(new_n3381_), .Y(new_n3446_));
  AOI21X1  g03253(.A0(new_n3385_), .A1(new_n3382_), .B0(new_n3446_), .Y(new_n3447_));
  XOR2X1   g03254(.A(new_n3447_), .B(new_n3445_), .Y(new_n3448_));
  XOR2X1   g03255(.A(new_n3448_), .B(new_n3443_), .Y(new_n3449_));
  XOR2X1   g03256(.A(new_n3449_), .B(new_n3422_), .Y(new_n3450_));
  XOR2X1   g03257(.A(new_n3450_), .B(new_n3417_), .Y(new_n3451_));
  XOR2X1   g03258(.A(new_n3451_), .B(new_n3414_), .Y(new_n3452_));
  INVX1    g03259(.A(new_n3276_), .Y(new_n3453_));
  OR2X1    g03260(.A(new_n3201_), .B(new_n3144_), .Y(new_n3454_));
  AOI21X1  g03261(.A0(new_n3454_), .A1(new_n3272_), .B0(new_n3275_), .Y(new_n3455_));
  AOI21X1  g03262(.A0(new_n3315_), .A1(new_n3453_), .B0(new_n3455_), .Y(new_n3456_));
  AND2X1   g03263(.A(new_n3398_), .B(new_n3395_), .Y(new_n3457_));
  AOI21X1  g03264(.A0(new_n3399_), .A1(new_n3392_), .B0(new_n3457_), .Y(new_n3458_));
  AOI22X1  g03265(.A0(\a[46] ), .A1(\a[0] ), .B0(\a[42] ), .B1(\a[4] ), .Y(new_n3459_));
  INVX1    g03266(.A(\a[46] ), .Y(new_n3460_));
  NOR4X1   g03267(.A(new_n3460_), .B(new_n3096_), .C(new_n340_), .D(new_n194_), .Y(new_n3461_));
  AND2X1   g03268(.A(\a[43] ), .B(\a[42] ), .Y(new_n3462_));
  NOR4X1   g03269(.A(new_n3460_), .B(new_n3037_), .C(new_n223_), .D(new_n194_), .Y(new_n3463_));
  AOI21X1  g03270(.A0(new_n3462_), .A1(new_n294_), .B0(new_n3463_), .Y(new_n3464_));
  NOR2X1   g03271(.A(new_n3464_), .B(new_n3461_), .Y(new_n3465_));
  NOR2X1   g03272(.A(new_n3465_), .B(new_n3461_), .Y(new_n3466_));
  INVX1    g03273(.A(new_n3466_), .Y(new_n3467_));
  NAND2X1  g03274(.A(\a[43] ), .B(\a[3] ), .Y(new_n3468_));
  OAI22X1  g03275(.A0(new_n3468_), .A1(new_n3465_), .B0(new_n3467_), .B1(new_n3459_), .Y(new_n3469_));
  NAND4X1  g03276(.A(\a[37] ), .B(\a[35] ), .C(\a[11] ), .D(\a[9] ), .Y(new_n3470_));
  NAND4X1  g03277(.A(\a[37] ), .B(\a[36] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n3471_));
  AOI22X1  g03278(.A0(new_n3471_), .A1(new_n3470_), .B0(new_n2682_), .B1(new_n1002_), .Y(new_n3472_));
  NAND2X1  g03279(.A(\a[37] ), .B(\a[9] ), .Y(new_n3473_));
  AOI21X1  g03280(.A0(new_n2682_), .A1(new_n1002_), .B0(new_n3472_), .Y(new_n3474_));
  INVX1    g03281(.A(new_n3474_), .Y(new_n3475_));
  AOI22X1  g03282(.A0(\a[36] ), .A1(\a[10] ), .B0(\a[35] ), .B1(\a[11] ), .Y(new_n3476_));
  OAI22X1  g03283(.A0(new_n3476_), .A1(new_n3475_), .B0(new_n3473_), .B1(new_n3472_), .Y(new_n3477_));
  XOR2X1   g03284(.A(new_n3477_), .B(new_n3469_), .Y(new_n3478_));
  AOI22X1  g03285(.A0(new_n1871_), .A1(new_n1148_), .B0(new_n1995_), .B1(new_n1099_), .Y(new_n3479_));
  AOI21X1  g03286(.A0(new_n1770_), .A1(new_n1236_), .B0(new_n3479_), .Y(new_n3480_));
  AND2X1   g03287(.A(\a[27] ), .B(\a[19] ), .Y(new_n3481_));
  INVX1    g03288(.A(new_n3481_), .Y(new_n3482_));
  INVX1    g03289(.A(new_n1995_), .Y(new_n3483_));
  INVX1    g03290(.A(new_n1871_), .Y(new_n3484_));
  OAI22X1  g03291(.A0(new_n3484_), .A1(new_n1149_), .B0(new_n3483_), .B1(new_n1521_), .Y(new_n3485_));
  AOI21X1  g03292(.A0(new_n1770_), .A1(new_n1236_), .B0(new_n3485_), .Y(new_n3486_));
  INVX1    g03293(.A(new_n3486_), .Y(new_n3487_));
  AOI22X1  g03294(.A0(\a[26] ), .A1(\a[20] ), .B0(\a[25] ), .B1(\a[21] ), .Y(new_n3488_));
  OAI22X1  g03295(.A0(new_n3488_), .A1(new_n3487_), .B0(new_n3482_), .B1(new_n3480_), .Y(new_n3489_));
  INVX1    g03296(.A(new_n3489_), .Y(new_n3490_));
  XOR2X1   g03297(.A(new_n3490_), .B(new_n3478_), .Y(new_n3491_));
  NAND4X1  g03298(.A(\a[30] ), .B(\a[28] ), .C(\a[18] ), .D(\a[16] ), .Y(new_n3492_));
  NAND4X1  g03299(.A(\a[30] ), .B(\a[29] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n3493_));
  AOI22X1  g03300(.A0(new_n3493_), .A1(new_n3492_), .B0(new_n1674_), .B1(new_n796_), .Y(new_n3494_));
  AND2X1   g03301(.A(\a[30] ), .B(\a[16] ), .Y(new_n3495_));
  INVX1    g03302(.A(new_n3495_), .Y(new_n3496_));
  AOI21X1  g03303(.A0(new_n1674_), .A1(new_n796_), .B0(new_n3494_), .Y(new_n3497_));
  INVX1    g03304(.A(new_n3497_), .Y(new_n3498_));
  AOI22X1  g03305(.A0(\a[29] ), .A1(\a[17] ), .B0(\a[28] ), .B1(\a[18] ), .Y(new_n3499_));
  OAI22X1  g03306(.A0(new_n3499_), .A1(new_n3498_), .B0(new_n3496_), .B1(new_n3494_), .Y(new_n3500_));
  XOR2X1   g03307(.A(new_n3500_), .B(new_n3310_), .Y(new_n3501_));
  AOI22X1  g03308(.A0(\a[39] ), .A1(\a[7] ), .B0(\a[38] ), .B1(\a[8] ), .Y(new_n3502_));
  AND2X1   g03309(.A(\a[39] ), .B(\a[38] ), .Y(new_n3503_));
  AND2X1   g03310(.A(new_n3503_), .B(new_n325_), .Y(new_n3504_));
  OAI21X1  g03311(.A0(new_n3502_), .A1(new_n3504_), .B0(new_n2468_), .Y(new_n3505_));
  INVX1    g03312(.A(new_n3502_), .Y(new_n3506_));
  AOI21X1  g03313(.A0(new_n3506_), .A1(new_n2468_), .B0(new_n3504_), .Y(new_n3507_));
  INVX1    g03314(.A(new_n3507_), .Y(new_n3508_));
  OAI21X1  g03315(.A0(new_n3508_), .A1(new_n3502_), .B0(new_n3505_), .Y(new_n3509_));
  INVX1    g03316(.A(new_n3509_), .Y(new_n3510_));
  XOR2X1   g03317(.A(new_n3510_), .B(new_n3501_), .Y(new_n3511_));
  XOR2X1   g03318(.A(new_n3511_), .B(new_n3491_), .Y(new_n3512_));
  INVX1    g03319(.A(new_n3512_), .Y(new_n3513_));
  XOR2X1   g03320(.A(new_n3513_), .B(new_n3458_), .Y(new_n3514_));
  XOR2X1   g03321(.A(new_n3514_), .B(new_n3456_), .Y(new_n3515_));
  NOR2X1   g03322(.A(new_n3367_), .B(new_n3358_), .Y(new_n3516_));
  AOI21X1  g03323(.A0(new_n3366_), .A1(new_n3186_), .B0(new_n3516_), .Y(new_n3517_));
  AND2X1   g03324(.A(new_n3337_), .B(new_n3328_), .Y(new_n3518_));
  AOI21X1  g03325(.A0(new_n3346_), .A1(new_n3338_), .B0(new_n3518_), .Y(new_n3519_));
  XOR2X1   g03326(.A(new_n3519_), .B(new_n3517_), .Y(new_n3520_));
  AND2X1   g03327(.A(new_n3300_), .B(new_n3292_), .Y(new_n3521_));
  AOI21X1  g03328(.A0(new_n3312_), .A1(new_n3301_), .B0(new_n3521_), .Y(new_n3522_));
  XOR2X1   g03329(.A(new_n3522_), .B(new_n3520_), .Y(new_n3523_));
  NAND2X1  g03330(.A(new_n3282_), .B(new_n3279_), .Y(new_n3524_));
  OAI21X1  g03331(.A0(new_n3314_), .A1(new_n3283_), .B0(new_n3524_), .Y(new_n3525_));
  INVX1    g03332(.A(new_n3355_), .Y(new_n3526_));
  XOR2X1   g03333(.A(new_n3526_), .B(new_n3325_), .Y(new_n3527_));
  XOR2X1   g03334(.A(new_n3527_), .B(new_n3335_), .Y(new_n3528_));
  AND2X1   g03335(.A(new_n3213_), .B(new_n3151_), .Y(new_n3529_));
  AOI21X1  g03336(.A0(new_n3278_), .A1(new_n3277_), .B0(new_n3529_), .Y(new_n3530_));
  AND2X1   g03337(.A(\a[45] ), .B(\a[1] ), .Y(new_n3531_));
  XOR2X1   g03338(.A(new_n3531_), .B(new_n1530_), .Y(new_n3532_));
  XOR2X1   g03339(.A(new_n3532_), .B(new_n3303_), .Y(new_n3533_));
  XOR2X1   g03340(.A(new_n3533_), .B(new_n3344_), .Y(new_n3534_));
  INVX1    g03341(.A(new_n3534_), .Y(new_n3535_));
  XOR2X1   g03342(.A(new_n3535_), .B(new_n3530_), .Y(new_n3536_));
  INVX1    g03343(.A(new_n3536_), .Y(new_n3537_));
  XOR2X1   g03344(.A(new_n3537_), .B(new_n3528_), .Y(new_n3538_));
  INVX1    g03345(.A(new_n3538_), .Y(new_n3539_));
  XOR2X1   g03346(.A(new_n3539_), .B(new_n3525_), .Y(new_n3540_));
  XOR2X1   g03347(.A(new_n3540_), .B(new_n3523_), .Y(new_n3541_));
  XOR2X1   g03348(.A(new_n3541_), .B(new_n3515_), .Y(new_n3542_));
  XOR2X1   g03349(.A(new_n3542_), .B(new_n3452_), .Y(new_n3543_));
  INVX1    g03350(.A(new_n3403_), .Y(new_n3544_));
  NOR2X1   g03351(.A(new_n3405_), .B(new_n3544_), .Y(new_n3545_));
  INVX1    g03352(.A(new_n3545_), .Y(new_n3546_));
  AND2X1   g03353(.A(new_n3405_), .B(new_n3544_), .Y(new_n3547_));
  OAI21X1  g03354(.A0(new_n3410_), .A1(new_n3547_), .B0(new_n3546_), .Y(new_n3548_));
  XOR2X1   g03355(.A(new_n3548_), .B(new_n3543_), .Y(\asquared[47] ));
  AND2X1   g03356(.A(new_n3450_), .B(new_n3417_), .Y(new_n3550_));
  AOI21X1  g03357(.A0(new_n3451_), .A1(new_n3414_), .B0(new_n3550_), .Y(new_n3551_));
  NOR2X1   g03358(.A(new_n3514_), .B(new_n3456_), .Y(new_n3552_));
  AOI21X1  g03359(.A0(new_n3541_), .A1(new_n3515_), .B0(new_n3552_), .Y(new_n3553_));
  AOI22X1  g03360(.A0(\a[47] ), .A1(\a[0] ), .B0(\a[45] ), .B1(\a[2] ), .Y(new_n3554_));
  INVX1    g03361(.A(new_n3554_), .Y(new_n3555_));
  AND2X1   g03362(.A(new_n3531_), .B(new_n1530_), .Y(new_n3556_));
  AND2X1   g03363(.A(\a[47] ), .B(\a[45] ), .Y(new_n3557_));
  AND2X1   g03364(.A(new_n3557_), .B(new_n197_), .Y(new_n3558_));
  AOI21X1  g03365(.A0(new_n3555_), .A1(new_n3556_), .B0(new_n3558_), .Y(new_n3559_));
  NAND2X1  g03366(.A(new_n3559_), .B(new_n3555_), .Y(new_n3560_));
  OAI21X1  g03367(.A0(new_n3558_), .A1(new_n3554_), .B0(new_n3556_), .Y(new_n3561_));
  AND2X1   g03368(.A(new_n3561_), .B(new_n3560_), .Y(new_n3562_));
  OAI22X1  g03369(.A0(new_n2430_), .A1(new_n795_), .B0(new_n2076_), .B1(new_n793_), .Y(new_n3563_));
  OAI21X1  g03370(.A0(new_n2197_), .A1(new_n797_), .B0(new_n3563_), .Y(new_n3564_));
  AND2X1   g03371(.A(\a[31] ), .B(\a[16] ), .Y(new_n3565_));
  AOI21X1  g03372(.A0(new_n2196_), .A1(new_n796_), .B0(new_n3563_), .Y(new_n3566_));
  OAI22X1  g03373(.A0(new_n1684_), .A1(new_n616_), .B0(new_n1803_), .B1(new_n675_), .Y(new_n3567_));
  AOI22X1  g03374(.A0(new_n3567_), .A1(new_n3566_), .B0(new_n3565_), .B1(new_n3564_), .Y(new_n3568_));
  XOR2X1   g03375(.A(new_n3568_), .B(new_n3562_), .Y(new_n3569_));
  INVX1    g03376(.A(new_n1996_), .Y(new_n3570_));
  OAI22X1  g03377(.A0(new_n3570_), .A1(new_n1149_), .B0(new_n1672_), .B1(new_n1521_), .Y(new_n3571_));
  OAI21X1  g03378(.A0(new_n3483_), .A1(new_n1794_), .B0(new_n3571_), .Y(new_n3572_));
  AND2X1   g03379(.A(\a[28] ), .B(\a[19] ), .Y(new_n3573_));
  AOI21X1  g03380(.A0(new_n1995_), .A1(new_n1236_), .B0(new_n3571_), .Y(new_n3574_));
  OAI22X1  g03381(.A0(new_n1679_), .A1(new_n934_), .B0(new_n1263_), .B1(new_n1098_), .Y(new_n3575_));
  AOI22X1  g03382(.A0(new_n3575_), .A1(new_n3574_), .B0(new_n3573_), .B1(new_n3572_), .Y(new_n3576_));
  XOR2X1   g03383(.A(new_n3576_), .B(new_n3569_), .Y(new_n3577_));
  XOR2X1   g03384(.A(new_n3497_), .B(new_n3437_), .Y(new_n3578_));
  INVX1    g03385(.A(new_n3578_), .Y(new_n3579_));
  NOR4X1   g03386(.A(new_n3037_), .B(new_n2219_), .C(new_n549_), .D(new_n340_), .Y(new_n3580_));
  NAND4X1  g03387(.A(\a[44] ), .B(\a[43] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n3581_));
  NAND4X1  g03388(.A(\a[44] ), .B(\a[32] ), .C(\a[15] ), .D(\a[3] ), .Y(new_n3582_));
  AOI21X1  g03389(.A0(new_n3582_), .A1(new_n3581_), .B0(new_n3580_), .Y(new_n3583_));
  NAND2X1  g03390(.A(\a[44] ), .B(\a[3] ), .Y(new_n3584_));
  OR2X1    g03391(.A(new_n3583_), .B(new_n3580_), .Y(new_n3585_));
  AOI22X1  g03392(.A0(\a[43] ), .A1(\a[4] ), .B0(\a[32] ), .B1(\a[15] ), .Y(new_n3586_));
  OAI22X1  g03393(.A0(new_n3586_), .A1(new_n3585_), .B0(new_n3584_), .B1(new_n3583_), .Y(new_n3587_));
  XOR2X1   g03394(.A(new_n3587_), .B(new_n3579_), .Y(new_n3588_));
  NAND4X1  g03395(.A(\a[39] ), .B(\a[38] ), .C(\a[9] ), .D(\a[8] ), .Y(new_n3589_));
  NAND4X1  g03396(.A(\a[39] ), .B(\a[36] ), .C(\a[11] ), .D(\a[8] ), .Y(new_n3590_));
  AOI22X1  g03397(.A0(new_n3590_), .A1(new_n3589_), .B0(new_n2484_), .B1(new_n813_), .Y(new_n3591_));
  AOI21X1  g03398(.A0(new_n2484_), .A1(new_n813_), .B0(new_n3591_), .Y(new_n3592_));
  OAI22X1  g03399(.A0(new_n2519_), .A1(new_n341_), .B0(new_n2583_), .B1(new_n488_), .Y(new_n3593_));
  NOR3X1   g03400(.A(new_n3591_), .B(new_n2652_), .C(new_n413_), .Y(new_n3594_));
  AOI21X1  g03401(.A0(new_n3593_), .A1(new_n3592_), .B0(new_n3594_), .Y(new_n3595_));
  AND2X1   g03402(.A(\a[37] ), .B(\a[10] ), .Y(new_n3596_));
  INVX1    g03403(.A(new_n3596_), .Y(new_n3597_));
  AOI22X1  g03404(.A0(\a[25] ), .A1(\a[22] ), .B0(\a[24] ), .B1(\a[23] ), .Y(new_n3598_));
  AND2X1   g03405(.A(new_n1394_), .B(new_n1532_), .Y(new_n3599_));
  NOR3X1   g03406(.A(new_n3598_), .B(new_n3599_), .C(new_n3597_), .Y(new_n3600_));
  INVX1    g03407(.A(new_n3598_), .Y(new_n3601_));
  AOI21X1  g03408(.A0(new_n3601_), .A1(new_n3596_), .B0(new_n3599_), .Y(new_n3602_));
  INVX1    g03409(.A(new_n3602_), .Y(new_n3603_));
  OAI22X1  g03410(.A0(new_n3603_), .A1(new_n3598_), .B0(new_n3600_), .B1(new_n3597_), .Y(new_n3604_));
  XOR2X1   g03411(.A(new_n3604_), .B(new_n3595_), .Y(new_n3605_));
  NOR4X1   g03412(.A(new_n3081_), .B(new_n1851_), .C(new_n490_), .D(new_n230_), .Y(new_n3606_));
  AND2X1   g03413(.A(\a[42] ), .B(\a[41] ), .Y(new_n3607_));
  AND2X1   g03414(.A(\a[42] ), .B(\a[14] ), .Y(new_n3608_));
  AOI22X1  g03415(.A0(new_n3608_), .A1(new_n2408_), .B0(new_n3607_), .B1(new_n295_), .Y(new_n3609_));
  OR2X1    g03416(.A(new_n3609_), .B(new_n3606_), .Y(new_n3610_));
  AND2X1   g03417(.A(\a[42] ), .B(\a[5] ), .Y(new_n3611_));
  OAI22X1  g03418(.A0(new_n3081_), .A1(new_n230_), .B0(new_n1851_), .B1(new_n490_), .Y(new_n3612_));
  INVX1    g03419(.A(new_n3606_), .Y(new_n3613_));
  AND2X1   g03420(.A(new_n3609_), .B(new_n3613_), .Y(new_n3614_));
  AOI22X1  g03421(.A0(new_n3614_), .A1(new_n3612_), .B0(new_n3611_), .B1(new_n3610_), .Y(new_n3615_));
  XOR2X1   g03422(.A(new_n3615_), .B(new_n3605_), .Y(new_n3616_));
  XOR2X1   g03423(.A(new_n3616_), .B(new_n3588_), .Y(new_n3617_));
  XOR2X1   g03424(.A(new_n3617_), .B(new_n3577_), .Y(new_n3618_));
  NOR2X1   g03425(.A(new_n3510_), .B(new_n3501_), .Y(new_n3619_));
  AOI21X1  g03426(.A0(new_n3500_), .A1(new_n3311_), .B0(new_n3619_), .Y(new_n3620_));
  INVX1    g03427(.A(new_n3620_), .Y(new_n3621_));
  AND2X1   g03428(.A(new_n3526_), .B(new_n3325_), .Y(new_n3622_));
  AOI21X1  g03429(.A0(new_n3527_), .A1(new_n3336_), .B0(new_n3622_), .Y(new_n3623_));
  XOR2X1   g03430(.A(new_n3623_), .B(new_n3621_), .Y(new_n3624_));
  OAI21X1  g03431(.A0(new_n3460_), .A1(new_n202_), .B0(new_n1185_), .Y(new_n3625_));
  NAND3X1  g03432(.A(\a[46] ), .B(\a[24] ), .C(\a[1] ), .Y(new_n3626_));
  AND2X1   g03433(.A(new_n3626_), .B(new_n3625_), .Y(new_n3627_));
  XOR2X1   g03434(.A(new_n3627_), .B(new_n3474_), .Y(new_n3628_));
  XOR2X1   g03435(.A(new_n3628_), .B(new_n3508_), .Y(new_n3629_));
  XOR2X1   g03436(.A(new_n3629_), .B(new_n3624_), .Y(new_n3630_));
  AND2X1   g03437(.A(new_n3618_), .B(new_n3630_), .Y(new_n3631_));
  INVX1    g03438(.A(new_n3631_), .Y(new_n3632_));
  NAND2X1  g03439(.A(new_n3632_), .B(new_n3618_), .Y(new_n3633_));
  NOR2X1   g03440(.A(new_n3533_), .B(new_n3344_), .Y(new_n3634_));
  AOI21X1  g03441(.A0(new_n3532_), .A1(new_n3302_), .B0(new_n3634_), .Y(new_n3635_));
  NOR4X1   g03442(.A(new_n3036_), .B(new_n2557_), .C(new_n453_), .D(new_n532_), .Y(new_n3636_));
  AND2X1   g03443(.A(\a[40] ), .B(\a[34] ), .Y(new_n3637_));
  AOI22X1  g03444(.A0(new_n3637_), .A1(new_n826_), .B0(new_n2361_), .B1(new_n586_), .Y(new_n3638_));
  NOR2X1   g03445(.A(new_n3638_), .B(new_n3636_), .Y(new_n3639_));
  NOR3X1   g03446(.A(new_n3639_), .B(new_n2028_), .C(new_n591_), .Y(new_n3640_));
  NOR2X1   g03447(.A(new_n3639_), .B(new_n3636_), .Y(new_n3641_));
  OAI22X1  g03448(.A0(new_n3036_), .A1(new_n532_), .B0(new_n2557_), .B1(new_n453_), .Y(new_n3642_));
  AOI21X1  g03449(.A0(new_n3642_), .A1(new_n3641_), .B0(new_n3640_), .Y(new_n3643_));
  XOR2X1   g03450(.A(new_n3643_), .B(new_n3635_), .Y(new_n3644_));
  INVX1    g03451(.A(new_n3644_), .Y(new_n3645_));
  AND2X1   g03452(.A(new_n3364_), .B(new_n3298_), .Y(new_n3646_));
  AOI21X1  g03453(.A0(new_n3444_), .A1(new_n3290_), .B0(new_n3646_), .Y(new_n3647_));
  XOR2X1   g03454(.A(new_n3647_), .B(new_n3645_), .Y(new_n3648_));
  INVX1    g03455(.A(new_n3648_), .Y(new_n3649_));
  OR2X1    g03456(.A(new_n3535_), .B(new_n3530_), .Y(new_n3650_));
  OAI21X1  g03457(.A0(new_n3537_), .A1(new_n3528_), .B0(new_n3650_), .Y(new_n3651_));
  XOR2X1   g03458(.A(new_n3651_), .B(new_n3649_), .Y(new_n3652_));
  OR2X1    g03459(.A(new_n3519_), .B(new_n3517_), .Y(new_n3653_));
  AND2X1   g03460(.A(new_n3312_), .B(new_n3301_), .Y(new_n3654_));
  OAI21X1  g03461(.A0(new_n3654_), .A1(new_n3521_), .B0(new_n3520_), .Y(new_n3655_));
  AND2X1   g03462(.A(new_n3655_), .B(new_n3653_), .Y(new_n3656_));
  XOR2X1   g03463(.A(new_n3656_), .B(new_n3652_), .Y(new_n3657_));
  XOR2X1   g03464(.A(new_n3618_), .B(new_n3630_), .Y(new_n3658_));
  AND2X1   g03465(.A(new_n3658_), .B(new_n3657_), .Y(new_n3659_));
  AOI21X1  g03466(.A0(new_n3632_), .A1(new_n3630_), .B0(new_n3657_), .Y(new_n3660_));
  AOI21X1  g03467(.A0(new_n3660_), .A1(new_n3633_), .B0(new_n3659_), .Y(new_n3661_));
  NAND2X1  g03468(.A(new_n3661_), .B(new_n3553_), .Y(new_n3662_));
  AND2X1   g03469(.A(new_n3421_), .B(new_n3419_), .Y(new_n3663_));
  AOI21X1  g03470(.A0(new_n3449_), .A1(new_n3422_), .B0(new_n3663_), .Y(new_n3664_));
  INVX1    g03471(.A(new_n3664_), .Y(new_n3665_));
  NAND2X1  g03472(.A(new_n3538_), .B(new_n3525_), .Y(new_n3666_));
  OAI21X1  g03473(.A0(new_n3540_), .A1(new_n3523_), .B0(new_n3666_), .Y(new_n3667_));
  XOR2X1   g03474(.A(new_n3667_), .B(new_n3665_), .Y(new_n3668_));
  XOR2X1   g03475(.A(new_n3486_), .B(new_n3429_), .Y(new_n3669_));
  XOR2X1   g03476(.A(new_n3669_), .B(new_n3467_), .Y(new_n3670_));
  INVX1    g03477(.A(new_n3670_), .Y(new_n3671_));
  AND2X1   g03478(.A(new_n3477_), .B(new_n3469_), .Y(new_n3672_));
  AOI21X1  g03479(.A0(new_n3489_), .A1(new_n3478_), .B0(new_n3672_), .Y(new_n3673_));
  XOR2X1   g03480(.A(new_n3673_), .B(new_n3671_), .Y(new_n3674_));
  INVX1    g03481(.A(new_n3431_), .Y(new_n3675_));
  OR2X1    g03482(.A(new_n3439_), .B(new_n3675_), .Y(new_n3676_));
  OAI21X1  g03483(.A0(new_n3442_), .A1(new_n3440_), .B0(new_n3676_), .Y(new_n3677_));
  XOR2X1   g03484(.A(new_n3677_), .B(new_n3674_), .Y(new_n3678_));
  INVX1    g03485(.A(new_n3511_), .Y(new_n3679_));
  OR2X1    g03486(.A(new_n3679_), .B(new_n3491_), .Y(new_n3680_));
  OAI21X1  g03487(.A0(new_n3512_), .A1(new_n3458_), .B0(new_n3680_), .Y(new_n3681_));
  NOR2X1   g03488(.A(new_n3447_), .B(new_n3445_), .Y(new_n3682_));
  AOI21X1  g03489(.A0(new_n3448_), .A1(new_n3443_), .B0(new_n3682_), .Y(new_n3683_));
  XOR2X1   g03490(.A(new_n3683_), .B(new_n3681_), .Y(new_n3684_));
  XOR2X1   g03491(.A(new_n3684_), .B(new_n3678_), .Y(new_n3685_));
  XOR2X1   g03492(.A(new_n3685_), .B(new_n3668_), .Y(new_n3686_));
  XOR2X1   g03493(.A(new_n3661_), .B(new_n3553_), .Y(new_n3687_));
  NOR2X1   g03494(.A(new_n3687_), .B(new_n3686_), .Y(new_n3688_));
  OR2X1    g03495(.A(new_n3661_), .B(new_n3553_), .Y(new_n3689_));
  AND2X1   g03496(.A(new_n3689_), .B(new_n3686_), .Y(new_n3690_));
  AOI21X1  g03497(.A0(new_n3690_), .A1(new_n3662_), .B0(new_n3688_), .Y(new_n3691_));
  XOR2X1   g03498(.A(new_n3691_), .B(new_n3551_), .Y(new_n3692_));
  NOR2X1   g03499(.A(new_n3542_), .B(new_n3452_), .Y(new_n3693_));
  INVX1    g03500(.A(new_n3693_), .Y(new_n3694_));
  AND2X1   g03501(.A(new_n3542_), .B(new_n3452_), .Y(new_n3695_));
  AOI21X1  g03502(.A0(new_n3548_), .A1(new_n3694_), .B0(new_n3695_), .Y(new_n3696_));
  XOR2X1   g03503(.A(new_n3696_), .B(new_n3692_), .Y(\asquared[48] ));
  AND2X1   g03504(.A(new_n3541_), .B(new_n3515_), .Y(new_n3698_));
  OAI21X1  g03505(.A0(new_n3698_), .A1(new_n3552_), .B0(new_n3661_), .Y(new_n3699_));
  OAI21X1  g03506(.A0(new_n3687_), .A1(new_n3686_), .B0(new_n3699_), .Y(new_n3700_));
  NOR2X1   g03507(.A(new_n3667_), .B(new_n3665_), .Y(new_n3701_));
  NAND2X1  g03508(.A(new_n3667_), .B(new_n3665_), .Y(new_n3702_));
  OAI21X1  g03509(.A0(new_n3685_), .A1(new_n3701_), .B0(new_n3702_), .Y(new_n3703_));
  INVX1    g03510(.A(new_n3678_), .Y(new_n3704_));
  INVX1    g03511(.A(new_n3683_), .Y(new_n3705_));
  NAND2X1  g03512(.A(new_n3705_), .B(new_n3681_), .Y(new_n3706_));
  OAI21X1  g03513(.A0(new_n3684_), .A1(new_n3704_), .B0(new_n3706_), .Y(new_n3707_));
  NAND2X1  g03514(.A(new_n3651_), .B(new_n3648_), .Y(new_n3708_));
  OAI21X1  g03515(.A0(new_n3656_), .A1(new_n3652_), .B0(new_n3708_), .Y(new_n3709_));
  NOR4X1   g03516(.A(new_n3096_), .B(new_n2557_), .C(new_n591_), .D(new_n230_), .Y(new_n3710_));
  NAND4X1  g03517(.A(\a[35] ), .B(\a[34] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n3711_));
  NAND4X1  g03518(.A(\a[42] ), .B(\a[34] ), .C(\a[14] ), .D(\a[6] ), .Y(new_n3712_));
  AOI21X1  g03519(.A0(new_n3712_), .A1(new_n3711_), .B0(new_n3710_), .Y(new_n3713_));
  OR2X1    g03520(.A(new_n3713_), .B(new_n3710_), .Y(new_n3714_));
  AOI22X1  g03521(.A0(\a[42] ), .A1(\a[6] ), .B0(\a[35] ), .B1(\a[13] ), .Y(new_n3715_));
  NAND2X1  g03522(.A(\a[34] ), .B(\a[14] ), .Y(new_n3716_));
  OAI22X1  g03523(.A0(new_n3716_), .A1(new_n3713_), .B0(new_n3715_), .B1(new_n3714_), .Y(new_n3717_));
  AND2X1   g03524(.A(\a[41] ), .B(\a[7] ), .Y(new_n3718_));
  INVX1    g03525(.A(new_n3718_), .Y(new_n3719_));
  NOR3X1   g03526(.A(new_n3181_), .B(new_n3036_), .C(new_n453_), .Y(new_n3720_));
  NAND4X1  g03527(.A(\a[41] ), .B(\a[40] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n3721_));
  NAND4X1  g03528(.A(\a[41] ), .B(\a[36] ), .C(\a[12] ), .D(\a[7] ), .Y(new_n3722_));
  AOI21X1  g03529(.A0(new_n3722_), .A1(new_n3721_), .B0(new_n3720_), .Y(new_n3723_));
  AOI22X1  g03530(.A0(\a[40] ), .A1(\a[8] ), .B0(\a[36] ), .B1(\a[12] ), .Y(new_n3724_));
  OR2X1    g03531(.A(new_n3723_), .B(new_n3720_), .Y(new_n3725_));
  OAI22X1  g03532(.A0(new_n3725_), .A1(new_n3724_), .B0(new_n3723_), .B1(new_n3719_), .Y(new_n3726_));
  XOR2X1   g03533(.A(new_n3726_), .B(new_n3717_), .Y(new_n3727_));
  NAND4X1  g03534(.A(\a[38] ), .B(\a[37] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n3728_));
  INVX1    g03535(.A(new_n3503_), .Y(new_n3729_));
  AND2X1   g03536(.A(\a[39] ), .B(\a[37] ), .Y(new_n3730_));
  INVX1    g03537(.A(new_n3730_), .Y(new_n3731_));
  OAI22X1  g03538(.A0(new_n3731_), .A1(new_n1519_), .B0(new_n3729_), .B1(new_n735_), .Y(new_n3732_));
  AND2X1   g03539(.A(new_n3732_), .B(new_n3728_), .Y(new_n3733_));
  NOR3X1   g03540(.A(new_n3733_), .B(new_n2652_), .C(new_n341_), .Y(new_n3734_));
  AOI21X1  g03541(.A0(new_n3164_), .A1(new_n1002_), .B0(new_n3732_), .Y(new_n3735_));
  AOI22X1  g03542(.A0(\a[38] ), .A1(\a[10] ), .B0(\a[37] ), .B1(\a[11] ), .Y(new_n3736_));
  INVX1    g03543(.A(new_n3736_), .Y(new_n3737_));
  AOI21X1  g03544(.A0(new_n3737_), .A1(new_n3735_), .B0(new_n3734_), .Y(new_n3738_));
  XOR2X1   g03545(.A(new_n3738_), .B(new_n3727_), .Y(new_n3739_));
  OR2X1    g03546(.A(new_n3643_), .B(new_n3635_), .Y(new_n3740_));
  OAI21X1  g03547(.A0(new_n3647_), .A1(new_n3645_), .B0(new_n3740_), .Y(new_n3741_));
  XOR2X1   g03548(.A(new_n3741_), .B(new_n3739_), .Y(new_n3742_));
  AND2X1   g03549(.A(\a[15] ), .B(\a[5] ), .Y(new_n3743_));
  AND2X1   g03550(.A(\a[43] ), .B(\a[33] ), .Y(new_n3744_));
  NAND4X1  g03551(.A(\a[44] ), .B(\a[33] ), .C(\a[15] ), .D(\a[4] ), .Y(new_n3745_));
  NAND4X1  g03552(.A(\a[44] ), .B(\a[43] ), .C(\a[5] ), .D(\a[4] ), .Y(new_n3746_));
  AOI22X1  g03553(.A0(new_n3746_), .A1(new_n3745_), .B0(new_n3744_), .B1(new_n3743_), .Y(new_n3747_));
  NAND4X1  g03554(.A(\a[43] ), .B(\a[33] ), .C(\a[15] ), .D(\a[5] ), .Y(new_n3748_));
  NAND3X1  g03555(.A(new_n3746_), .B(new_n3745_), .C(new_n3748_), .Y(new_n3749_));
  AOI22X1  g03556(.A0(\a[43] ), .A1(\a[5] ), .B0(\a[33] ), .B1(\a[15] ), .Y(new_n3750_));
  NAND2X1  g03557(.A(\a[44] ), .B(\a[4] ), .Y(new_n3751_));
  OAI22X1  g03558(.A0(new_n3751_), .A1(new_n3747_), .B0(new_n3750_), .B1(new_n3749_), .Y(new_n3752_));
  AOI22X1  g03559(.A0(new_n1996_), .A1(new_n2134_), .B0(new_n1671_), .B1(new_n1236_), .Y(new_n3753_));
  AOI21X1  g03560(.A0(new_n1995_), .A1(new_n1154_), .B0(new_n3753_), .Y(new_n3754_));
  NAND2X1  g03561(.A(\a[28] ), .B(\a[20] ), .Y(new_n3755_));
  AOI22X1  g03562(.A0(\a[27] ), .A1(\a[21] ), .B0(\a[26] ), .B1(\a[22] ), .Y(new_n3756_));
  AOI21X1  g03563(.A0(new_n1995_), .A1(new_n1154_), .B0(new_n3754_), .Y(new_n3757_));
  INVX1    g03564(.A(new_n3757_), .Y(new_n3758_));
  OAI22X1  g03565(.A0(new_n3758_), .A1(new_n3756_), .B0(new_n3755_), .B1(new_n3754_), .Y(new_n3759_));
  XOR2X1   g03566(.A(new_n3759_), .B(new_n3752_), .Y(new_n3760_));
  AOI22X1  g03567(.A0(new_n2429_), .A1(new_n2213_), .B0(new_n2075_), .B1(new_n796_), .Y(new_n3761_));
  AOI21X1  g03568(.A0(new_n2196_), .A1(new_n855_), .B0(new_n3761_), .Y(new_n3762_));
  AND2X1   g03569(.A(\a[31] ), .B(\a[17] ), .Y(new_n3763_));
  INVX1    g03570(.A(new_n3763_), .Y(new_n3764_));
  AOI21X1  g03571(.A0(new_n2196_), .A1(new_n855_), .B0(new_n3762_), .Y(new_n3765_));
  INVX1    g03572(.A(new_n3765_), .Y(new_n3766_));
  AOI22X1  g03573(.A0(\a[30] ), .A1(\a[18] ), .B0(\a[29] ), .B1(\a[19] ), .Y(new_n3767_));
  OAI22X1  g03574(.A0(new_n3767_), .A1(new_n3766_), .B0(new_n3764_), .B1(new_n3762_), .Y(new_n3768_));
  INVX1    g03575(.A(new_n3768_), .Y(new_n3769_));
  XOR2X1   g03576(.A(new_n3769_), .B(new_n3760_), .Y(new_n3770_));
  XOR2X1   g03577(.A(new_n3770_), .B(new_n3742_), .Y(new_n3771_));
  XOR2X1   g03578(.A(new_n3771_), .B(new_n3709_), .Y(new_n3772_));
  XOR2X1   g03579(.A(new_n3772_), .B(new_n3707_), .Y(new_n3773_));
  XOR2X1   g03580(.A(new_n3773_), .B(new_n3703_), .Y(new_n3774_));
  AOI21X1  g03581(.A0(new_n3658_), .A1(new_n3657_), .B0(new_n3631_), .Y(new_n3775_));
  NOR2X1   g03582(.A(new_n3673_), .B(new_n3671_), .Y(new_n3776_));
  AOI21X1  g03583(.A0(new_n3677_), .A1(new_n3674_), .B0(new_n3776_), .Y(new_n3777_));
  NOR2X1   g03584(.A(new_n3623_), .B(new_n3620_), .Y(new_n3778_));
  INVX1    g03585(.A(new_n3778_), .Y(new_n3779_));
  OAI21X1  g03586(.A0(new_n3629_), .A1(new_n3624_), .B0(new_n3779_), .Y(new_n3780_));
  XOR2X1   g03587(.A(new_n3780_), .B(new_n3777_), .Y(new_n3781_));
  AND2X1   g03588(.A(\a[48] ), .B(\a[0] ), .Y(new_n3782_));
  XOR2X1   g03589(.A(new_n3782_), .B(new_n3626_), .Y(new_n3783_));
  AND2X1   g03590(.A(\a[47] ), .B(\a[1] ), .Y(new_n3784_));
  XOR2X1   g03591(.A(new_n3784_), .B(new_n2706_), .Y(new_n3785_));
  XOR2X1   g03592(.A(new_n3785_), .B(new_n3783_), .Y(new_n3786_));
  INVX1    g03593(.A(new_n3786_), .Y(new_n3787_));
  NOR2X1   g03594(.A(new_n3486_), .B(new_n3429_), .Y(new_n3788_));
  AOI21X1  g03595(.A0(new_n3669_), .A1(new_n3467_), .B0(new_n3788_), .Y(new_n3789_));
  XOR2X1   g03596(.A(new_n3789_), .B(new_n3787_), .Y(new_n3790_));
  INVX1    g03597(.A(new_n3790_), .Y(new_n3791_));
  NAND2X1  g03598(.A(new_n3587_), .B(new_n3578_), .Y(new_n3792_));
  OAI21X1  g03599(.A0(new_n3497_), .A1(new_n3437_), .B0(new_n3792_), .Y(new_n3793_));
  XOR2X1   g03600(.A(new_n3793_), .B(new_n3791_), .Y(new_n3794_));
  XOR2X1   g03601(.A(new_n3794_), .B(new_n3781_), .Y(new_n3795_));
  NAND2X1  g03602(.A(new_n3795_), .B(new_n3775_), .Y(new_n3796_));
  INVX1    g03603(.A(new_n3775_), .Y(new_n3797_));
  XOR2X1   g03604(.A(new_n3795_), .B(new_n3797_), .Y(new_n3798_));
  INVX1    g03605(.A(new_n3614_), .Y(new_n3799_));
  XOR2X1   g03606(.A(new_n3592_), .B(new_n3574_), .Y(new_n3800_));
  XOR2X1   g03607(.A(new_n3800_), .B(new_n3799_), .Y(new_n3801_));
  INVX1    g03608(.A(new_n3801_), .Y(new_n3802_));
  AND2X1   g03609(.A(new_n3593_), .B(new_n3592_), .Y(new_n3803_));
  OAI21X1  g03610(.A0(new_n3594_), .A1(new_n3803_), .B0(new_n3604_), .Y(new_n3804_));
  OAI21X1  g03611(.A0(new_n3615_), .A1(new_n3605_), .B0(new_n3804_), .Y(new_n3805_));
  XOR2X1   g03612(.A(new_n3805_), .B(new_n3802_), .Y(new_n3806_));
  XOR2X1   g03613(.A(new_n3603_), .B(new_n3641_), .Y(new_n3807_));
  AND2X1   g03614(.A(\a[46] ), .B(\a[32] ), .Y(new_n3808_));
  AND2X1   g03615(.A(\a[46] ), .B(\a[45] ), .Y(new_n3809_));
  AOI22X1  g03616(.A0(new_n3809_), .A1(new_n231_), .B0(new_n3808_), .B1(new_n857_), .Y(new_n3810_));
  INVX1    g03617(.A(\a[45] ), .Y(new_n3811_));
  NOR4X1   g03618(.A(new_n3811_), .B(new_n2219_), .C(new_n571_), .D(new_n223_), .Y(new_n3812_));
  AND2X1   g03619(.A(\a[46] ), .B(\a[2] ), .Y(new_n3813_));
  OAI21X1  g03620(.A0(new_n3812_), .A1(new_n3810_), .B0(new_n3813_), .Y(new_n3814_));
  INVX1    g03621(.A(new_n3812_), .Y(new_n3815_));
  AND2X1   g03622(.A(new_n3815_), .B(new_n3810_), .Y(new_n3816_));
  INVX1    g03623(.A(new_n3816_), .Y(new_n3817_));
  AOI22X1  g03624(.A0(\a[45] ), .A1(\a[3] ), .B0(\a[32] ), .B1(\a[16] ), .Y(new_n3818_));
  OAI21X1  g03625(.A0(new_n3818_), .A1(new_n3817_), .B0(new_n3814_), .Y(new_n3819_));
  XOR2X1   g03626(.A(new_n3819_), .B(new_n3807_), .Y(new_n3820_));
  XOR2X1   g03627(.A(new_n3820_), .B(new_n3806_), .Y(new_n3821_));
  INVX1    g03628(.A(new_n3616_), .Y(new_n3822_));
  OR2X1    g03629(.A(new_n3617_), .B(new_n3577_), .Y(new_n3823_));
  OAI21X1  g03630(.A0(new_n3822_), .A1(new_n3588_), .B0(new_n3823_), .Y(new_n3824_));
  XOR2X1   g03631(.A(new_n3824_), .B(new_n3821_), .Y(new_n3825_));
  INVX1    g03632(.A(new_n3559_), .Y(new_n3826_));
  INVX1    g03633(.A(new_n3566_), .Y(new_n3827_));
  XOR2X1   g03634(.A(new_n3585_), .B(new_n3827_), .Y(new_n3828_));
  XOR2X1   g03635(.A(new_n3828_), .B(new_n3826_), .Y(new_n3829_));
  NAND2X1  g03636(.A(new_n3627_), .B(new_n3475_), .Y(new_n3830_));
  OAI21X1  g03637(.A0(new_n3628_), .A1(new_n3507_), .B0(new_n3830_), .Y(new_n3831_));
  OR2X1    g03638(.A(new_n3568_), .B(new_n3562_), .Y(new_n3832_));
  INVX1    g03639(.A(new_n3569_), .Y(new_n3833_));
  OAI21X1  g03640(.A0(new_n3576_), .A1(new_n3833_), .B0(new_n3832_), .Y(new_n3834_));
  XOR2X1   g03641(.A(new_n3834_), .B(new_n3831_), .Y(new_n3835_));
  XOR2X1   g03642(.A(new_n3835_), .B(new_n3829_), .Y(new_n3836_));
  XOR2X1   g03643(.A(new_n3836_), .B(new_n3825_), .Y(new_n3837_));
  NOR2X1   g03644(.A(new_n3795_), .B(new_n3775_), .Y(new_n3838_));
  NOR2X1   g03645(.A(new_n3837_), .B(new_n3838_), .Y(new_n3839_));
  AOI22X1  g03646(.A0(new_n3839_), .A1(new_n3796_), .B0(new_n3837_), .B1(new_n3798_), .Y(new_n3840_));
  XOR2X1   g03647(.A(new_n3840_), .B(new_n3774_), .Y(new_n3841_));
  AND2X1   g03648(.A(new_n3841_), .B(new_n3700_), .Y(new_n3842_));
  INVX1    g03649(.A(new_n3842_), .Y(new_n3843_));
  INVX1    g03650(.A(new_n3551_), .Y(new_n3844_));
  AND2X1   g03651(.A(new_n3691_), .B(new_n3844_), .Y(new_n3845_));
  INVX1    g03652(.A(new_n3845_), .Y(new_n3846_));
  NOR2X1   g03653(.A(new_n3691_), .B(new_n3844_), .Y(new_n3847_));
  OAI21X1  g03654(.A0(new_n3696_), .A1(new_n3847_), .B0(new_n3846_), .Y(new_n3848_));
  NOR2X1   g03655(.A(new_n3841_), .B(new_n3700_), .Y(new_n3849_));
  INVX1    g03656(.A(new_n3849_), .Y(new_n3850_));
  AOI21X1  g03657(.A0(new_n3843_), .A1(new_n3850_), .B0(new_n3848_), .Y(new_n3851_));
  AND2X1   g03658(.A(new_n3850_), .B(new_n3848_), .Y(new_n3852_));
  AOI21X1  g03659(.A0(new_n3852_), .A1(new_n3843_), .B0(new_n3851_), .Y(\asquared[49] ));
  AND2X1   g03660(.A(new_n3795_), .B(new_n3797_), .Y(new_n3854_));
  AOI21X1  g03661(.A0(new_n3837_), .A1(new_n3798_), .B0(new_n3854_), .Y(new_n3855_));
  AND2X1   g03662(.A(new_n3824_), .B(new_n3821_), .Y(new_n3856_));
  AOI21X1  g03663(.A0(new_n3836_), .A1(new_n3825_), .B0(new_n3856_), .Y(new_n3857_));
  INVX1    g03664(.A(new_n3857_), .Y(new_n3858_));
  AND2X1   g03665(.A(new_n3677_), .B(new_n3674_), .Y(new_n3859_));
  OAI21X1  g03666(.A0(new_n3859_), .A1(new_n3776_), .B0(new_n3780_), .Y(new_n3860_));
  OAI21X1  g03667(.A0(new_n3794_), .A1(new_n3781_), .B0(new_n3860_), .Y(new_n3861_));
  AOI22X1  g03668(.A0(\a[42] ), .A1(\a[7] ), .B0(\a[41] ), .B1(\a[8] ), .Y(new_n3862_));
  AND2X1   g03669(.A(\a[36] ), .B(\a[13] ), .Y(new_n3863_));
  INVX1    g03670(.A(new_n3863_), .Y(new_n3864_));
  AND2X1   g03671(.A(new_n3607_), .B(new_n325_), .Y(new_n3865_));
  NOR3X1   g03672(.A(new_n3864_), .B(new_n3865_), .C(new_n3862_), .Y(new_n3866_));
  NOR2X1   g03673(.A(new_n3866_), .B(new_n3865_), .Y(new_n3867_));
  INVX1    g03674(.A(new_n3867_), .Y(new_n3868_));
  OAI22X1  g03675(.A0(new_n3868_), .A1(new_n3862_), .B0(new_n3866_), .B1(new_n3864_), .Y(new_n3869_));
  AND2X1   g03676(.A(\a[38] ), .B(\a[11] ), .Y(new_n3870_));
  AOI22X1  g03677(.A0(\a[26] ), .A1(\a[23] ), .B0(\a[25] ), .B1(\a[24] ), .Y(new_n3871_));
  INVX1    g03678(.A(new_n3871_), .Y(new_n3872_));
  NAND2X1  g03679(.A(\a[26] ), .B(\a[23] ), .Y(new_n3873_));
  NOR3X1   g03680(.A(new_n3873_), .B(new_n1326_), .C(new_n1185_), .Y(new_n3874_));
  OR4X1    g03681(.A(new_n3871_), .B(new_n3874_), .C(new_n2519_), .D(new_n488_), .Y(new_n3875_));
  AOI21X1  g03682(.A0(new_n3872_), .A1(new_n3870_), .B0(new_n3874_), .Y(new_n3876_));
  AOI22X1  g03683(.A0(new_n3876_), .A1(new_n3872_), .B0(new_n3875_), .B1(new_n3870_), .Y(new_n3877_));
  XOR2X1   g03684(.A(new_n3877_), .B(new_n3869_), .Y(new_n3878_));
  INVX1    g03685(.A(new_n3878_), .Y(new_n3879_));
  NOR4X1   g03686(.A(new_n3037_), .B(new_n2557_), .C(new_n490_), .D(new_n230_), .Y(new_n3880_));
  NOR4X1   g03687(.A(new_n3037_), .B(new_n2028_), .C(new_n549_), .D(new_n230_), .Y(new_n3881_));
  AOI21X1  g03688(.A0(new_n2361_), .A1(new_n691_), .B0(new_n3881_), .Y(new_n3882_));
  OR2X1    g03689(.A(new_n3882_), .B(new_n3880_), .Y(new_n3883_));
  AND2X1   g03690(.A(\a[34] ), .B(\a[15] ), .Y(new_n3884_));
  OAI22X1  g03691(.A0(new_n3037_), .A1(new_n230_), .B0(new_n2557_), .B1(new_n490_), .Y(new_n3885_));
  AND2X1   g03692(.A(new_n2361_), .B(new_n691_), .Y(new_n3886_));
  NOR3X1   g03693(.A(new_n3886_), .B(new_n3881_), .C(new_n3880_), .Y(new_n3887_));
  AOI22X1  g03694(.A0(new_n3887_), .A1(new_n3885_), .B0(new_n3884_), .B1(new_n3883_), .Y(new_n3888_));
  XOR2X1   g03695(.A(new_n3888_), .B(new_n3879_), .Y(new_n3889_));
  AOI22X1  g03696(.A0(\a[47] ), .A1(\a[2] ), .B0(\a[46] ), .B1(\a[3] ), .Y(new_n3890_));
  AND2X1   g03697(.A(\a[27] ), .B(\a[22] ), .Y(new_n3891_));
  INVX1    g03698(.A(new_n3891_), .Y(new_n3892_));
  AND2X1   g03699(.A(\a[47] ), .B(\a[46] ), .Y(new_n3893_));
  AND2X1   g03700(.A(new_n3893_), .B(new_n231_), .Y(new_n3894_));
  NOR3X1   g03701(.A(new_n3892_), .B(new_n3894_), .C(new_n3890_), .Y(new_n3895_));
  NOR2X1   g03702(.A(new_n3895_), .B(new_n3894_), .Y(new_n3896_));
  INVX1    g03703(.A(new_n3896_), .Y(new_n3897_));
  OAI22X1  g03704(.A0(new_n3897_), .A1(new_n3890_), .B0(new_n3895_), .B1(new_n3892_), .Y(new_n3898_));
  OAI22X1  g03705(.A0(new_n2199_), .A1(new_n1149_), .B0(new_n2197_), .B1(new_n1521_), .Y(new_n3899_));
  OAI21X1  g03706(.A0(new_n1675_), .A1(new_n1794_), .B0(new_n3899_), .Y(new_n3900_));
  AND2X1   g03707(.A(\a[30] ), .B(\a[19] ), .Y(new_n3901_));
  AOI21X1  g03708(.A0(new_n1674_), .A1(new_n1236_), .B0(new_n3899_), .Y(new_n3902_));
  OAI22X1  g03709(.A0(new_n1803_), .A1(new_n934_), .B0(new_n1431_), .B1(new_n1098_), .Y(new_n3903_));
  AOI22X1  g03710(.A0(new_n3903_), .A1(new_n3902_), .B0(new_n3901_), .B1(new_n3900_), .Y(new_n3904_));
  XOR2X1   g03711(.A(new_n3904_), .B(new_n3898_), .Y(new_n3905_));
  NAND4X1  g03712(.A(\a[40] ), .B(\a[39] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n3906_));
  NAND4X1  g03713(.A(\a[40] ), .B(\a[37] ), .C(\a[12] ), .D(\a[9] ), .Y(new_n3907_));
  AOI22X1  g03714(.A0(new_n3907_), .A1(new_n3906_), .B0(new_n3730_), .B1(new_n396_), .Y(new_n3908_));
  NOR3X1   g03715(.A(new_n3908_), .B(new_n3036_), .C(new_n341_), .Y(new_n3909_));
  AOI21X1  g03716(.A0(new_n3730_), .A1(new_n396_), .B0(new_n3908_), .Y(new_n3910_));
  OAI22X1  g03717(.A0(new_n2652_), .A1(new_n570_), .B0(new_n2345_), .B1(new_n453_), .Y(new_n3911_));
  AOI21X1  g03718(.A0(new_n3911_), .A1(new_n3910_), .B0(new_n3909_), .Y(new_n3912_));
  XOR2X1   g03719(.A(new_n3912_), .B(new_n3905_), .Y(new_n3913_));
  INVX1    g03720(.A(new_n3913_), .Y(new_n3914_));
  INVX1    g03721(.A(\a[49] ), .Y(new_n3915_));
  AND2X1   g03722(.A(\a[5] ), .B(\a[0] ), .Y(new_n3916_));
  AOI22X1  g03723(.A0(new_n3916_), .A1(\a[44] ), .B0(new_n210_), .B1(\a[45] ), .Y(new_n3917_));
  AND2X1   g03724(.A(\a[45] ), .B(\a[44] ), .Y(new_n3918_));
  AND2X1   g03725(.A(new_n3918_), .B(new_n218_), .Y(new_n3919_));
  NOR3X1   g03726(.A(new_n3919_), .B(new_n3917_), .C(new_n3915_), .Y(new_n3920_));
  NOR3X1   g03727(.A(new_n3920_), .B(new_n3915_), .C(new_n194_), .Y(new_n3921_));
  NOR2X1   g03728(.A(new_n3920_), .B(new_n3919_), .Y(new_n3922_));
  AOI22X1  g03729(.A0(\a[45] ), .A1(\a[4] ), .B0(\a[44] ), .B1(\a[5] ), .Y(new_n3923_));
  INVX1    g03730(.A(new_n3923_), .Y(new_n3924_));
  AOI21X1  g03731(.A0(new_n3924_), .A1(new_n3922_), .B0(new_n3921_), .Y(new_n3925_));
  INVX1    g03732(.A(\a[48] ), .Y(new_n3926_));
  NOR3X1   g03733(.A(new_n3626_), .B(new_n3926_), .C(new_n194_), .Y(new_n3927_));
  NOR2X1   g03734(.A(new_n3785_), .B(new_n3783_), .Y(new_n3928_));
  NOR2X1   g03735(.A(new_n3928_), .B(new_n3927_), .Y(new_n3929_));
  INVX1    g03736(.A(new_n3929_), .Y(new_n3930_));
  XOR2X1   g03737(.A(new_n3930_), .B(new_n3925_), .Y(new_n3931_));
  OAI22X1  g03738(.A0(new_n2675_), .A1(new_n793_), .B0(new_n2673_), .B1(new_n795_), .Y(new_n3932_));
  OAI21X1  g03739(.A0(new_n2672_), .A1(new_n797_), .B0(new_n3932_), .Y(new_n3933_));
  AND2X1   g03740(.A(\a[33] ), .B(\a[16] ), .Y(new_n3934_));
  AOI21X1  g03741(.A0(new_n2671_), .A1(new_n796_), .B0(new_n3932_), .Y(new_n3935_));
  OAI22X1  g03742(.A0(new_n2219_), .A1(new_n616_), .B0(new_n1704_), .B1(new_n675_), .Y(new_n3936_));
  AOI22X1  g03743(.A0(new_n3936_), .A1(new_n3935_), .B0(new_n3934_), .B1(new_n3933_), .Y(new_n3937_));
  XOR2X1   g03744(.A(new_n3937_), .B(new_n3931_), .Y(new_n3938_));
  XOR2X1   g03745(.A(new_n3938_), .B(new_n3914_), .Y(new_n3939_));
  XOR2X1   g03746(.A(new_n3939_), .B(new_n3889_), .Y(new_n3940_));
  XOR2X1   g03747(.A(new_n3940_), .B(new_n3861_), .Y(new_n3941_));
  XOR2X1   g03748(.A(new_n3941_), .B(new_n3858_), .Y(new_n3942_));
  XOR2X1   g03749(.A(new_n3942_), .B(new_n3855_), .Y(new_n3943_));
  AND2X1   g03750(.A(new_n3771_), .B(new_n3709_), .Y(new_n3944_));
  AOI21X1  g03751(.A0(new_n3772_), .A1(new_n3707_), .B0(new_n3944_), .Y(new_n3945_));
  NOR2X1   g03752(.A(new_n3592_), .B(new_n3574_), .Y(new_n3946_));
  AOI21X1  g03753(.A0(new_n3800_), .A1(new_n3799_), .B0(new_n3946_), .Y(new_n3947_));
  OR4X1    g03754(.A(new_n3600_), .B(new_n3599_), .C(new_n3639_), .D(new_n3636_), .Y(new_n3948_));
  NOR2X1   g03755(.A(new_n3602_), .B(new_n3641_), .Y(new_n3949_));
  AOI21X1  g03756(.A0(new_n3819_), .A1(new_n3948_), .B0(new_n3949_), .Y(new_n3950_));
  XOR2X1   g03757(.A(new_n3950_), .B(new_n3947_), .Y(new_n3951_));
  AND2X1   g03758(.A(new_n3585_), .B(new_n3827_), .Y(new_n3952_));
  AOI21X1  g03759(.A0(new_n3828_), .A1(new_n3826_), .B0(new_n3952_), .Y(new_n3953_));
  XOR2X1   g03760(.A(new_n3953_), .B(new_n3951_), .Y(new_n3954_));
  NAND2X1  g03761(.A(new_n3805_), .B(new_n3801_), .Y(new_n3955_));
  OAI21X1  g03762(.A0(new_n3820_), .A1(new_n3806_), .B0(new_n3955_), .Y(new_n3956_));
  AND2X1   g03763(.A(new_n3834_), .B(new_n3831_), .Y(new_n3957_));
  AOI21X1  g03764(.A0(new_n3835_), .A1(new_n3829_), .B0(new_n3957_), .Y(new_n3958_));
  XOR2X1   g03765(.A(new_n3958_), .B(new_n3956_), .Y(new_n3959_));
  XOR2X1   g03766(.A(new_n3959_), .B(new_n3954_), .Y(new_n3960_));
  AND2X1   g03767(.A(new_n3960_), .B(new_n3945_), .Y(new_n3961_));
  XOR2X1   g03768(.A(new_n3960_), .B(new_n3945_), .Y(new_n3962_));
  XOR2X1   g03769(.A(new_n3766_), .B(new_n3714_), .Y(new_n3963_));
  XOR2X1   g03770(.A(new_n3963_), .B(new_n3725_), .Y(new_n3964_));
  AND2X1   g03771(.A(new_n3759_), .B(new_n3752_), .Y(new_n3965_));
  AOI21X1  g03772(.A0(new_n3768_), .A1(new_n3760_), .B0(new_n3965_), .Y(new_n3966_));
  INVX1    g03773(.A(new_n3966_), .Y(new_n3967_));
  XOR2X1   g03774(.A(new_n3967_), .B(new_n3964_), .Y(new_n3968_));
  INVX1    g03775(.A(new_n3968_), .Y(new_n3969_));
  NOR2X1   g03776(.A(new_n3789_), .B(new_n3787_), .Y(new_n3970_));
  AOI21X1  g03777(.A0(new_n3793_), .A1(new_n3790_), .B0(new_n3970_), .Y(new_n3971_));
  XOR2X1   g03778(.A(new_n3971_), .B(new_n3969_), .Y(new_n3972_));
  INVX1    g03779(.A(new_n3739_), .Y(new_n3973_));
  NAND2X1  g03780(.A(new_n3741_), .B(new_n3973_), .Y(new_n3974_));
  OAI21X1  g03781(.A0(new_n3770_), .A1(new_n3742_), .B0(new_n3974_), .Y(new_n3975_));
  XOR2X1   g03782(.A(new_n3975_), .B(new_n3972_), .Y(new_n3976_));
  XOR2X1   g03783(.A(new_n3817_), .B(new_n3749_), .Y(new_n3977_));
  XOR2X1   g03784(.A(new_n3977_), .B(new_n3757_), .Y(new_n3978_));
  AND2X1   g03785(.A(new_n3726_), .B(new_n3717_), .Y(new_n3979_));
  INVX1    g03786(.A(new_n3738_), .Y(new_n3980_));
  AOI21X1  g03787(.A0(new_n3980_), .A1(new_n3727_), .B0(new_n3979_), .Y(new_n3981_));
  AND2X1   g03788(.A(new_n3784_), .B(new_n1134_), .Y(new_n3982_));
  AOI21X1  g03789(.A0(\a[48] ), .A1(\a[1] ), .B0(\a[25] ), .Y(new_n3983_));
  AOI21X1  g03790(.A0(new_n1283_), .A1(\a[48] ), .B0(new_n3983_), .Y(new_n3984_));
  XOR2X1   g03791(.A(new_n3984_), .B(new_n3982_), .Y(new_n3985_));
  INVX1    g03792(.A(new_n3985_), .Y(new_n3986_));
  XOR2X1   g03793(.A(new_n3986_), .B(new_n3735_), .Y(new_n3987_));
  INVX1    g03794(.A(new_n3987_), .Y(new_n3988_));
  XOR2X1   g03795(.A(new_n3988_), .B(new_n3981_), .Y(new_n3989_));
  INVX1    g03796(.A(new_n3989_), .Y(new_n3990_));
  XOR2X1   g03797(.A(new_n3990_), .B(new_n3978_), .Y(new_n3991_));
  INVX1    g03798(.A(new_n3991_), .Y(new_n3992_));
  XOR2X1   g03799(.A(new_n3992_), .B(new_n3976_), .Y(new_n3993_));
  OAI21X1  g03800(.A0(new_n3960_), .A1(new_n3945_), .B0(new_n3993_), .Y(new_n3994_));
  OAI22X1  g03801(.A0(new_n3994_), .A1(new_n3961_), .B0(new_n3993_), .B1(new_n3962_), .Y(new_n3995_));
  XOR2X1   g03802(.A(new_n3995_), .B(new_n3943_), .Y(new_n3996_));
  AND2X1   g03803(.A(new_n3773_), .B(new_n3703_), .Y(new_n3997_));
  AOI21X1  g03804(.A0(new_n3840_), .A1(new_n3774_), .B0(new_n3997_), .Y(new_n3998_));
  XOR2X1   g03805(.A(new_n3998_), .B(new_n3996_), .Y(new_n3999_));
  AOI21X1  g03806(.A0(new_n3850_), .A1(new_n3848_), .B0(new_n3842_), .Y(new_n4000_));
  XOR2X1   g03807(.A(new_n4000_), .B(new_n3999_), .Y(\asquared[50] ));
  INVX1    g03808(.A(new_n3942_), .Y(new_n4002_));
  OR2X1    g03809(.A(new_n4002_), .B(new_n3855_), .Y(new_n4003_));
  OAI21X1  g03810(.A0(new_n3995_), .A1(new_n3943_), .B0(new_n4003_), .Y(new_n4004_));
  INVX1    g03811(.A(new_n3960_), .Y(new_n4005_));
  NOR2X1   g03812(.A(new_n4005_), .B(new_n3945_), .Y(new_n4006_));
  NOR2X1   g03813(.A(new_n3993_), .B(new_n3962_), .Y(new_n4007_));
  OR2X1    g03814(.A(new_n4007_), .B(new_n4006_), .Y(new_n4008_));
  NAND2X1  g03815(.A(\a[45] ), .B(\a[35] ), .Y(new_n4009_));
  NOR3X1   g03816(.A(new_n4009_), .B(new_n549_), .C(new_n255_), .Y(new_n4010_));
  NAND4X1  g03817(.A(\a[45] ), .B(\a[34] ), .C(\a[16] ), .D(\a[5] ), .Y(new_n4011_));
  NAND4X1  g03818(.A(\a[35] ), .B(\a[34] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n4012_));
  AOI21X1  g03819(.A0(new_n4012_), .A1(new_n4011_), .B0(new_n4010_), .Y(new_n4013_));
  OR2X1    g03820(.A(new_n4013_), .B(new_n4010_), .Y(new_n4014_));
  AOI22X1  g03821(.A0(\a[45] ), .A1(\a[5] ), .B0(\a[35] ), .B1(\a[15] ), .Y(new_n4015_));
  NAND2X1  g03822(.A(\a[34] ), .B(\a[16] ), .Y(new_n4016_));
  OAI22X1  g03823(.A0(new_n4016_), .A1(new_n4013_), .B0(new_n4015_), .B1(new_n4014_), .Y(new_n4017_));
  AND2X1   g03824(.A(\a[32] ), .B(\a[28] ), .Y(new_n4018_));
  AOI22X1  g03825(.A0(new_n4018_), .A1(new_n2660_), .B0(new_n1671_), .B1(new_n1394_), .Y(new_n4019_));
  NOR4X1   g03826(.A(new_n2219_), .B(new_n1679_), .C(new_n1216_), .D(new_n675_), .Y(new_n4020_));
  NOR2X1   g03827(.A(new_n4020_), .B(new_n4019_), .Y(new_n4021_));
  NAND2X1  g03828(.A(\a[28] ), .B(\a[22] ), .Y(new_n4022_));
  AOI22X1  g03829(.A0(\a[32] ), .A1(\a[18] ), .B0(\a[27] ), .B1(\a[23] ), .Y(new_n4023_));
  INVX1    g03830(.A(new_n4020_), .Y(new_n4024_));
  AND2X1   g03831(.A(new_n4024_), .B(new_n4019_), .Y(new_n4025_));
  INVX1    g03832(.A(new_n4025_), .Y(new_n4026_));
  OAI22X1  g03833(.A0(new_n4026_), .A1(new_n4023_), .B0(new_n4022_), .B1(new_n4021_), .Y(new_n4027_));
  XOR2X1   g03834(.A(new_n4027_), .B(new_n4017_), .Y(new_n4028_));
  NAND2X1  g03835(.A(new_n3984_), .B(new_n3982_), .Y(new_n4029_));
  OAI21X1  g03836(.A0(new_n3986_), .A1(new_n3735_), .B0(new_n4029_), .Y(new_n4030_));
  XOR2X1   g03837(.A(new_n4030_), .B(new_n4028_), .Y(new_n4031_));
  AOI22X1  g03838(.A0(\a[50] ), .A1(\a[0] ), .B0(\a[48] ), .B1(\a[2] ), .Y(new_n4032_));
  INVX1    g03839(.A(new_n4032_), .Y(new_n4033_));
  AND2X1   g03840(.A(new_n1283_), .B(\a[48] ), .Y(new_n4034_));
  AND2X1   g03841(.A(\a[50] ), .B(\a[48] ), .Y(new_n4035_));
  AND2X1   g03842(.A(new_n4035_), .B(new_n197_), .Y(new_n4036_));
  AOI21X1  g03843(.A0(new_n4033_), .A1(new_n4034_), .B0(new_n4036_), .Y(new_n4037_));
  NAND2X1  g03844(.A(new_n4037_), .B(new_n4033_), .Y(new_n4038_));
  OAI21X1  g03845(.A0(new_n4036_), .A1(new_n4032_), .B0(new_n4034_), .Y(new_n4039_));
  AND2X1   g03846(.A(new_n4039_), .B(new_n4038_), .Y(new_n4040_));
  INVX1    g03847(.A(\a[47] ), .Y(new_n4041_));
  NOR4X1   g03848(.A(new_n3460_), .B(new_n1851_), .C(new_n616_), .D(new_n340_), .Y(new_n4042_));
  NAND4X1  g03849(.A(\a[47] ), .B(\a[46] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n4043_));
  NAND4X1  g03850(.A(\a[47] ), .B(\a[33] ), .C(\a[17] ), .D(\a[3] ), .Y(new_n4044_));
  AOI21X1  g03851(.A0(new_n4044_), .A1(new_n4043_), .B0(new_n4042_), .Y(new_n4045_));
  NOR3X1   g03852(.A(new_n4045_), .B(new_n4041_), .C(new_n223_), .Y(new_n4046_));
  NOR2X1   g03853(.A(new_n4045_), .B(new_n4042_), .Y(new_n4047_));
  OAI22X1  g03854(.A0(new_n3460_), .A1(new_n340_), .B0(new_n1851_), .B1(new_n616_), .Y(new_n4048_));
  AOI21X1  g03855(.A0(new_n4048_), .A1(new_n4047_), .B0(new_n4046_), .Y(new_n4049_));
  XOR2X1   g03856(.A(new_n4049_), .B(new_n4040_), .Y(new_n4050_));
  OAI22X1  g03857(.A0(new_n2430_), .A1(new_n1149_), .B0(new_n2076_), .B1(new_n1521_), .Y(new_n4051_));
  OAI21X1  g03858(.A0(new_n2197_), .A1(new_n1794_), .B0(new_n4051_), .Y(new_n4052_));
  AND2X1   g03859(.A(\a[31] ), .B(\a[19] ), .Y(new_n4053_));
  AOI21X1  g03860(.A0(new_n2196_), .A1(new_n1236_), .B0(new_n4051_), .Y(new_n4054_));
  OAI22X1  g03861(.A0(new_n1684_), .A1(new_n934_), .B0(new_n1803_), .B1(new_n1098_), .Y(new_n4055_));
  AOI22X1  g03862(.A0(new_n4055_), .A1(new_n4054_), .B0(new_n4053_), .B1(new_n4052_), .Y(new_n4056_));
  XOR2X1   g03863(.A(new_n4056_), .B(new_n4050_), .Y(new_n4057_));
  INVX1    g03864(.A(new_n4057_), .Y(new_n4058_));
  NOR4X1   g03865(.A(new_n3037_), .B(new_n2583_), .C(new_n490_), .D(new_n532_), .Y(new_n4059_));
  NAND4X1  g03866(.A(\a[44] ), .B(\a[43] ), .C(\a[7] ), .D(\a[6] ), .Y(new_n4060_));
  NAND4X1  g03867(.A(\a[44] ), .B(\a[36] ), .C(\a[14] ), .D(\a[6] ), .Y(new_n4061_));
  AOI21X1  g03868(.A0(new_n4061_), .A1(new_n4060_), .B0(new_n4059_), .Y(new_n4062_));
  OR2X1    g03869(.A(new_n4062_), .B(new_n4059_), .Y(new_n4063_));
  AOI22X1  g03870(.A0(\a[43] ), .A1(\a[7] ), .B0(\a[36] ), .B1(\a[14] ), .Y(new_n4064_));
  NAND2X1  g03871(.A(\a[44] ), .B(\a[6] ), .Y(new_n4065_));
  OAI22X1  g03872(.A0(new_n4065_), .A1(new_n4062_), .B0(new_n4064_), .B1(new_n4063_), .Y(new_n4066_));
  AND2X1   g03873(.A(\a[41] ), .B(\a[37] ), .Y(new_n4067_));
  NAND4X1  g03874(.A(\a[42] ), .B(\a[41] ), .C(\a[9] ), .D(\a[8] ), .Y(new_n4068_));
  NAND4X1  g03875(.A(\a[42] ), .B(\a[37] ), .C(\a[13] ), .D(\a[8] ), .Y(new_n4069_));
  AOI22X1  g03876(.A0(new_n4069_), .A1(new_n4068_), .B0(new_n4067_), .B1(new_n430_), .Y(new_n4070_));
  NAND2X1  g03877(.A(\a[42] ), .B(\a[8] ), .Y(new_n4071_));
  NAND4X1  g03878(.A(\a[41] ), .B(\a[37] ), .C(\a[13] ), .D(\a[9] ), .Y(new_n4072_));
  NAND3X1  g03879(.A(new_n4069_), .B(new_n4068_), .C(new_n4072_), .Y(new_n4073_));
  AOI22X1  g03880(.A0(\a[41] ), .A1(\a[9] ), .B0(\a[37] ), .B1(\a[13] ), .Y(new_n4074_));
  OAI22X1  g03881(.A0(new_n4074_), .A1(new_n4073_), .B0(new_n4071_), .B1(new_n4070_), .Y(new_n4075_));
  XOR2X1   g03882(.A(new_n4075_), .B(new_n4066_), .Y(new_n4076_));
  AND2X1   g03883(.A(\a[40] ), .B(\a[39] ), .Y(new_n4077_));
  AOI22X1  g03884(.A0(new_n3503_), .A1(new_n482_), .B0(new_n2663_), .B1(new_n396_), .Y(new_n4078_));
  AOI21X1  g03885(.A0(new_n4077_), .A1(new_n1002_), .B0(new_n4078_), .Y(new_n4079_));
  AND2X1   g03886(.A(\a[38] ), .B(\a[12] ), .Y(new_n4080_));
  INVX1    g03887(.A(new_n4080_), .Y(new_n4081_));
  AOI21X1  g03888(.A0(new_n4077_), .A1(new_n1002_), .B0(new_n4079_), .Y(new_n4082_));
  INVX1    g03889(.A(new_n4082_), .Y(new_n4083_));
  AOI22X1  g03890(.A0(\a[40] ), .A1(\a[10] ), .B0(\a[39] ), .B1(\a[11] ), .Y(new_n4084_));
  OAI22X1  g03891(.A0(new_n4084_), .A1(new_n4083_), .B0(new_n4081_), .B1(new_n4079_), .Y(new_n4085_));
  XOR2X1   g03892(.A(new_n4085_), .B(new_n4076_), .Y(new_n4086_));
  XOR2X1   g03893(.A(new_n4086_), .B(new_n4058_), .Y(new_n4087_));
  XOR2X1   g03894(.A(new_n4087_), .B(new_n4031_), .Y(new_n4088_));
  AND2X1   g03895(.A(new_n3835_), .B(new_n3829_), .Y(new_n4089_));
  OAI21X1  g03896(.A0(new_n4089_), .A1(new_n3957_), .B0(new_n3956_), .Y(new_n4090_));
  OAI21X1  g03897(.A0(new_n3959_), .A1(new_n3954_), .B0(new_n4090_), .Y(new_n4091_));
  AND2X1   g03898(.A(new_n4088_), .B(new_n4091_), .Y(new_n4092_));
  INVX1    g03899(.A(new_n4092_), .Y(new_n4093_));
  NAND2X1  g03900(.A(new_n4093_), .B(new_n4088_), .Y(new_n4094_));
  NAND2X1  g03901(.A(new_n3975_), .B(new_n3972_), .Y(new_n4095_));
  NOR2X1   g03902(.A(new_n3975_), .B(new_n3972_), .Y(new_n4096_));
  OAI21X1  g03903(.A0(new_n3992_), .A1(new_n4096_), .B0(new_n4095_), .Y(new_n4097_));
  XOR2X1   g03904(.A(new_n4088_), .B(new_n4091_), .Y(new_n4098_));
  AND2X1   g03905(.A(new_n4098_), .B(new_n4097_), .Y(new_n4099_));
  AOI21X1  g03906(.A0(new_n4093_), .A1(new_n4091_), .B0(new_n4097_), .Y(new_n4100_));
  AOI21X1  g03907(.A0(new_n4100_), .A1(new_n4094_), .B0(new_n4099_), .Y(new_n4101_));
  XOR2X1   g03908(.A(new_n4101_), .B(new_n4008_), .Y(new_n4102_));
  NAND2X1  g03909(.A(new_n3940_), .B(new_n3861_), .Y(new_n4103_));
  NOR2X1   g03910(.A(new_n3940_), .B(new_n3861_), .Y(new_n4104_));
  OAI21X1  g03911(.A0(new_n4104_), .A1(new_n3857_), .B0(new_n4103_), .Y(new_n4105_));
  NAND2X1  g03912(.A(new_n3967_), .B(new_n3964_), .Y(new_n4106_));
  OAI21X1  g03913(.A0(new_n3971_), .A1(new_n3969_), .B0(new_n4106_), .Y(new_n4107_));
  OR2X1    g03914(.A(new_n3988_), .B(new_n3981_), .Y(new_n4108_));
  OAI21X1  g03915(.A0(new_n3990_), .A1(new_n3978_), .B0(new_n4108_), .Y(new_n4109_));
  XOR2X1   g03916(.A(new_n4109_), .B(new_n4107_), .Y(new_n4110_));
  AND2X1   g03917(.A(new_n3766_), .B(new_n3714_), .Y(new_n4111_));
  AOI21X1  g03918(.A0(new_n3963_), .A1(new_n3725_), .B0(new_n4111_), .Y(new_n4112_));
  AND2X1   g03919(.A(new_n3817_), .B(new_n3749_), .Y(new_n4113_));
  AOI21X1  g03920(.A0(new_n3977_), .A1(new_n3758_), .B0(new_n4113_), .Y(new_n4114_));
  XOR2X1   g03921(.A(new_n4114_), .B(new_n4112_), .Y(new_n4115_));
  XOR2X1   g03922(.A(new_n3922_), .B(new_n3897_), .Y(new_n4116_));
  XOR2X1   g03923(.A(new_n4116_), .B(new_n3887_), .Y(new_n4117_));
  XOR2X1   g03924(.A(new_n4117_), .B(new_n4115_), .Y(new_n4118_));
  XOR2X1   g03925(.A(new_n4118_), .B(new_n4110_), .Y(new_n4119_));
  XOR2X1   g03926(.A(new_n4119_), .B(new_n4105_), .Y(new_n4120_));
  INVX1    g03927(.A(new_n3898_), .Y(new_n4121_));
  OR2X1    g03928(.A(new_n3904_), .B(new_n4121_), .Y(new_n4122_));
  OAI21X1  g03929(.A0(new_n3912_), .A1(new_n3905_), .B0(new_n4122_), .Y(new_n4123_));
  OR2X1    g03930(.A(new_n3929_), .B(new_n3925_), .Y(new_n4124_));
  OAI21X1  g03931(.A0(new_n3937_), .A1(new_n3931_), .B0(new_n4124_), .Y(new_n4125_));
  XOR2X1   g03932(.A(new_n4125_), .B(new_n4123_), .Y(new_n4126_));
  AND2X1   g03933(.A(\a[49] ), .B(\a[1] ), .Y(new_n4127_));
  XOR2X1   g03934(.A(new_n4127_), .B(new_n1650_), .Y(new_n4128_));
  XOR2X1   g03935(.A(new_n4128_), .B(new_n3876_), .Y(new_n4129_));
  XOR2X1   g03936(.A(new_n4129_), .B(new_n3910_), .Y(new_n4130_));
  XOR2X1   g03937(.A(new_n4130_), .B(new_n4126_), .Y(new_n4131_));
  XOR2X1   g03938(.A(new_n3935_), .B(new_n3902_), .Y(new_n4132_));
  XOR2X1   g03939(.A(new_n4132_), .B(new_n3868_), .Y(new_n4133_));
  INVX1    g03940(.A(new_n3869_), .Y(new_n4134_));
  OR2X1    g03941(.A(new_n3888_), .B(new_n3878_), .Y(new_n4135_));
  OAI21X1  g03942(.A0(new_n3877_), .A1(new_n4134_), .B0(new_n4135_), .Y(new_n4136_));
  XOR2X1   g03943(.A(new_n4136_), .B(new_n4133_), .Y(new_n4137_));
  INVX1    g03944(.A(new_n4137_), .Y(new_n4138_));
  AND2X1   g03945(.A(new_n3950_), .B(new_n3947_), .Y(new_n4139_));
  OR2X1    g03946(.A(new_n3950_), .B(new_n3947_), .Y(new_n4140_));
  OAI21X1  g03947(.A0(new_n3953_), .A1(new_n4139_), .B0(new_n4140_), .Y(new_n4141_));
  XOR2X1   g03948(.A(new_n4141_), .B(new_n4138_), .Y(new_n4142_));
  NOR2X1   g03949(.A(new_n3939_), .B(new_n3889_), .Y(new_n4143_));
  AOI21X1  g03950(.A0(new_n3938_), .A1(new_n3913_), .B0(new_n4143_), .Y(new_n4144_));
  XOR2X1   g03951(.A(new_n4144_), .B(new_n4142_), .Y(new_n4145_));
  XOR2X1   g03952(.A(new_n4145_), .B(new_n4131_), .Y(new_n4146_));
  XOR2X1   g03953(.A(new_n4146_), .B(new_n4120_), .Y(new_n4147_));
  XOR2X1   g03954(.A(new_n4147_), .B(new_n4102_), .Y(new_n4148_));
  AND2X1   g03955(.A(new_n4148_), .B(new_n4004_), .Y(new_n4149_));
  INVX1    g03956(.A(new_n4149_), .Y(new_n4150_));
  AND2X1   g03957(.A(new_n3840_), .B(new_n3774_), .Y(new_n4151_));
  NOR3X1   g03958(.A(new_n3996_), .B(new_n4151_), .C(new_n3997_), .Y(new_n4152_));
  OAI21X1  g03959(.A0(new_n4151_), .A1(new_n3997_), .B0(new_n3996_), .Y(new_n4153_));
  OAI21X1  g03960(.A0(new_n4000_), .A1(new_n4152_), .B0(new_n4153_), .Y(new_n4154_));
  NOR2X1   g03961(.A(new_n4148_), .B(new_n4004_), .Y(new_n4155_));
  INVX1    g03962(.A(new_n4155_), .Y(new_n4156_));
  AOI21X1  g03963(.A0(new_n4150_), .A1(new_n4156_), .B0(new_n4154_), .Y(new_n4157_));
  AND2X1   g03964(.A(new_n4156_), .B(new_n4154_), .Y(new_n4158_));
  AOI21X1  g03965(.A0(new_n4158_), .A1(new_n4150_), .B0(new_n4157_), .Y(\asquared[51] ));
  AOI21X1  g03966(.A0(new_n4156_), .A1(new_n4154_), .B0(new_n4149_), .Y(new_n4160_));
  AND2X1   g03967(.A(new_n4101_), .B(new_n4008_), .Y(new_n4161_));
  AND2X1   g03968(.A(new_n4147_), .B(new_n4102_), .Y(new_n4162_));
  OR2X1    g03969(.A(new_n4162_), .B(new_n4161_), .Y(new_n4163_));
  AND2X1   g03970(.A(new_n4119_), .B(new_n4105_), .Y(new_n4164_));
  AND2X1   g03971(.A(new_n4146_), .B(new_n4120_), .Y(new_n4165_));
  OR2X1    g03972(.A(new_n4165_), .B(new_n4164_), .Y(new_n4166_));
  NAND2X1  g03973(.A(new_n4145_), .B(new_n4131_), .Y(new_n4167_));
  OAI21X1  g03974(.A0(new_n4144_), .A1(new_n4142_), .B0(new_n4167_), .Y(new_n4168_));
  AND2X1   g03975(.A(new_n4109_), .B(new_n4107_), .Y(new_n4169_));
  AOI21X1  g03976(.A0(new_n4118_), .A1(new_n4110_), .B0(new_n4169_), .Y(new_n4170_));
  NAND4X1  g03977(.A(\a[49] ), .B(\a[26] ), .C(\a[24] ), .D(\a[1] ), .Y(new_n4171_));
  AND2X1   g03978(.A(\a[51] ), .B(\a[0] ), .Y(new_n4172_));
  XOR2X1   g03979(.A(new_n4172_), .B(new_n4171_), .Y(new_n4173_));
  AND2X1   g03980(.A(\a[50] ), .B(\a[1] ), .Y(new_n4174_));
  XOR2X1   g03981(.A(new_n4174_), .B(new_n1263_), .Y(new_n4175_));
  XOR2X1   g03982(.A(new_n4175_), .B(new_n4173_), .Y(new_n4176_));
  AND2X1   g03983(.A(\a[34] ), .B(\a[17] ), .Y(new_n4177_));
  AOI22X1  g03984(.A0(\a[32] ), .A1(\a[19] ), .B0(\a[31] ), .B1(\a[20] ), .Y(new_n4178_));
  INVX1    g03985(.A(new_n4178_), .Y(new_n4179_));
  NAND4X1  g03986(.A(\a[32] ), .B(\a[31] ), .C(\a[20] ), .D(\a[19] ), .Y(new_n4180_));
  NAND3X1  g03987(.A(new_n4180_), .B(new_n4179_), .C(new_n4177_), .Y(new_n4181_));
  AOI22X1  g03988(.A0(new_n4179_), .A1(new_n4177_), .B0(new_n2671_), .B1(new_n1099_), .Y(new_n4182_));
  AOI22X1  g03989(.A0(new_n4182_), .A1(new_n4179_), .B0(new_n4181_), .B1(new_n4177_), .Y(new_n4183_));
  XOR2X1   g03990(.A(new_n4183_), .B(new_n4176_), .Y(new_n4184_));
  NOR2X1   g03991(.A(new_n3935_), .B(new_n3902_), .Y(new_n4185_));
  AOI21X1  g03992(.A0(new_n4132_), .A1(new_n3868_), .B0(new_n4185_), .Y(new_n4186_));
  XOR2X1   g03993(.A(new_n4186_), .B(new_n4184_), .Y(new_n4187_));
  NOR4X1   g03994(.A(new_n3460_), .B(new_n2557_), .C(new_n571_), .D(new_n255_), .Y(new_n4188_));
  NAND4X1  g03995(.A(\a[46] ), .B(\a[33] ), .C(\a[18] ), .D(\a[5] ), .Y(new_n4189_));
  NAND4X1  g03996(.A(\a[35] ), .B(\a[33] ), .C(\a[18] ), .D(\a[16] ), .Y(new_n4190_));
  AOI21X1  g03997(.A0(new_n4190_), .A1(new_n4189_), .B0(new_n4188_), .Y(new_n4191_));
  OR2X1    g03998(.A(new_n4191_), .B(new_n4188_), .Y(new_n4192_));
  AOI22X1  g03999(.A0(\a[46] ), .A1(\a[5] ), .B0(\a[35] ), .B1(\a[16] ), .Y(new_n4193_));
  NAND2X1  g04000(.A(\a[33] ), .B(\a[18] ), .Y(new_n4194_));
  OAI22X1  g04001(.A0(new_n4194_), .A1(new_n4191_), .B0(new_n4193_), .B1(new_n4192_), .Y(new_n4195_));
  NAND4X1  g04002(.A(\a[30] ), .B(\a[28] ), .C(\a[23] ), .D(\a[21] ), .Y(new_n4196_));
  NAND4X1  g04003(.A(\a[30] ), .B(\a[29] ), .C(\a[22] ), .D(\a[21] ), .Y(new_n4197_));
  AOI22X1  g04004(.A0(new_n4197_), .A1(new_n4196_), .B0(new_n1674_), .B1(new_n1394_), .Y(new_n4198_));
  NAND2X1  g04005(.A(\a[30] ), .B(\a[21] ), .Y(new_n4199_));
  AOI22X1  g04006(.A0(\a[29] ), .A1(\a[22] ), .B0(\a[28] ), .B1(\a[23] ), .Y(new_n4200_));
  AOI21X1  g04007(.A0(new_n1674_), .A1(new_n1394_), .B0(new_n4198_), .Y(new_n4201_));
  INVX1    g04008(.A(new_n4201_), .Y(new_n4202_));
  OAI22X1  g04009(.A0(new_n4202_), .A1(new_n4200_), .B0(new_n4199_), .B1(new_n4198_), .Y(new_n4203_));
  XOR2X1   g04010(.A(new_n4203_), .B(new_n4195_), .Y(new_n4204_));
  AND2X1   g04011(.A(\a[36] ), .B(\a[15] ), .Y(new_n4205_));
  INVX1    g04012(.A(new_n4205_), .Y(new_n4206_));
  NOR4X1   g04013(.A(new_n3811_), .B(new_n2345_), .C(new_n490_), .D(new_n230_), .Y(new_n4207_));
  INVX1    g04014(.A(new_n4207_), .Y(new_n4208_));
  NOR4X1   g04015(.A(new_n3811_), .B(new_n2583_), .C(new_n549_), .D(new_n230_), .Y(new_n4209_));
  AND2X1   g04016(.A(new_n3330_), .B(new_n691_), .Y(new_n4210_));
  OR2X1    g04017(.A(new_n4210_), .B(new_n4209_), .Y(new_n4211_));
  AND2X1   g04018(.A(new_n4211_), .B(new_n4208_), .Y(new_n4212_));
  AOI22X1  g04019(.A0(\a[45] ), .A1(\a[6] ), .B0(\a[37] ), .B1(\a[14] ), .Y(new_n4213_));
  NOR3X1   g04020(.A(new_n4210_), .B(new_n4209_), .C(new_n4207_), .Y(new_n4214_));
  INVX1    g04021(.A(new_n4214_), .Y(new_n4215_));
  OAI22X1  g04022(.A0(new_n4215_), .A1(new_n4213_), .B0(new_n4212_), .B1(new_n4206_), .Y(new_n4216_));
  INVX1    g04023(.A(new_n4216_), .Y(new_n4217_));
  XOR2X1   g04024(.A(new_n4217_), .B(new_n4204_), .Y(new_n4218_));
  NOR4X1   g04025(.A(new_n3037_), .B(new_n2519_), .C(new_n591_), .D(new_n413_), .Y(new_n4219_));
  NAND4X1  g04026(.A(\a[44] ), .B(\a[43] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n4220_));
  NAND4X1  g04027(.A(\a[44] ), .B(\a[38] ), .C(\a[13] ), .D(\a[7] ), .Y(new_n4221_));
  AOI21X1  g04028(.A0(new_n4221_), .A1(new_n4220_), .B0(new_n4219_), .Y(new_n4222_));
  OR2X1    g04029(.A(new_n4222_), .B(new_n4219_), .Y(new_n4223_));
  AOI22X1  g04030(.A0(\a[43] ), .A1(\a[8] ), .B0(\a[38] ), .B1(\a[13] ), .Y(new_n4224_));
  NAND2X1  g04031(.A(\a[44] ), .B(\a[7] ), .Y(new_n4225_));
  OAI22X1  g04032(.A0(new_n4225_), .A1(new_n4222_), .B0(new_n4224_), .B1(new_n4223_), .Y(new_n4226_));
  AND2X1   g04033(.A(\a[42] ), .B(\a[9] ), .Y(new_n4227_));
  INVX1    g04034(.A(new_n4227_), .Y(new_n4228_));
  NAND4X1  g04035(.A(\a[42] ), .B(\a[39] ), .C(\a[12] ), .D(\a[9] ), .Y(new_n4229_));
  NAND4X1  g04036(.A(\a[42] ), .B(\a[41] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n4230_));
  AOI22X1  g04037(.A0(new_n4230_), .A1(new_n4229_), .B0(new_n2847_), .B1(new_n396_), .Y(new_n4231_));
  AOI21X1  g04038(.A0(new_n2847_), .A1(new_n396_), .B0(new_n4231_), .Y(new_n4232_));
  INVX1    g04039(.A(new_n4232_), .Y(new_n4233_));
  AOI22X1  g04040(.A0(\a[41] ), .A1(\a[10] ), .B0(\a[39] ), .B1(\a[12] ), .Y(new_n4234_));
  OAI22X1  g04041(.A0(new_n4234_), .A1(new_n4233_), .B0(new_n4231_), .B1(new_n4228_), .Y(new_n4235_));
  XOR2X1   g04042(.A(new_n4235_), .B(new_n4226_), .Y(new_n4236_));
  AND2X1   g04043(.A(\a[40] ), .B(\a[11] ), .Y(new_n4237_));
  INVX1    g04044(.A(new_n4237_), .Y(new_n4238_));
  AOI22X1  g04045(.A0(\a[27] ), .A1(\a[24] ), .B0(\a[26] ), .B1(\a[25] ), .Y(new_n4239_));
  AND2X1   g04046(.A(new_n1995_), .B(new_n1532_), .Y(new_n4240_));
  NOR3X1   g04047(.A(new_n4239_), .B(new_n4240_), .C(new_n4238_), .Y(new_n4241_));
  NOR2X1   g04048(.A(new_n4241_), .B(new_n4240_), .Y(new_n4242_));
  INVX1    g04049(.A(new_n4242_), .Y(new_n4243_));
  OAI22X1  g04050(.A0(new_n4243_), .A1(new_n4239_), .B0(new_n4241_), .B1(new_n4238_), .Y(new_n4244_));
  XOR2X1   g04051(.A(new_n4244_), .B(new_n4236_), .Y(new_n4245_));
  XOR2X1   g04052(.A(new_n4245_), .B(new_n4218_), .Y(new_n4246_));
  XOR2X1   g04053(.A(new_n4246_), .B(new_n4187_), .Y(new_n4247_));
  XOR2X1   g04054(.A(new_n4247_), .B(new_n4170_), .Y(new_n4248_));
  XOR2X1   g04055(.A(new_n4248_), .B(new_n4168_), .Y(new_n4249_));
  XOR2X1   g04056(.A(new_n4249_), .B(new_n4166_), .Y(new_n4250_));
  OR2X1    g04057(.A(new_n4099_), .B(new_n4092_), .Y(new_n4251_));
  AND2X1   g04058(.A(new_n4136_), .B(new_n4133_), .Y(new_n4252_));
  AOI21X1  g04059(.A0(new_n4141_), .A1(new_n4137_), .B0(new_n4252_), .Y(new_n4253_));
  AND2X1   g04060(.A(new_n4125_), .B(new_n4123_), .Y(new_n4254_));
  AOI21X1  g04061(.A0(new_n4130_), .A1(new_n4126_), .B0(new_n4254_), .Y(new_n4255_));
  XOR2X1   g04062(.A(new_n4255_), .B(new_n4253_), .Y(new_n4256_));
  OAI22X1  g04063(.A0(new_n3920_), .A1(new_n3919_), .B0(new_n3895_), .B1(new_n3894_), .Y(new_n4257_));
  OAI21X1  g04064(.A0(new_n4116_), .A1(new_n3887_), .B0(new_n4257_), .Y(new_n4258_));
  NOR3X1   g04065(.A(new_n3871_), .B(new_n2519_), .C(new_n488_), .Y(new_n4259_));
  OAI21X1  g04066(.A0(new_n4259_), .A1(new_n3874_), .B0(new_n4128_), .Y(new_n4260_));
  OAI21X1  g04067(.A0(new_n4129_), .A1(new_n3910_), .B0(new_n4260_), .Y(new_n4261_));
  XOR2X1   g04068(.A(new_n4261_), .B(new_n4258_), .Y(new_n4262_));
  OR2X1    g04069(.A(new_n4049_), .B(new_n4040_), .Y(new_n4263_));
  INVX1    g04070(.A(new_n4050_), .Y(new_n4264_));
  OAI21X1  g04071(.A0(new_n4056_), .A1(new_n4264_), .B0(new_n4263_), .Y(new_n4265_));
  XOR2X1   g04072(.A(new_n4265_), .B(new_n4262_), .Y(new_n4266_));
  XOR2X1   g04073(.A(new_n4266_), .B(new_n4256_), .Y(new_n4267_));
  XOR2X1   g04074(.A(new_n4267_), .B(new_n4251_), .Y(new_n4268_));
  AND2X1   g04075(.A(new_n4086_), .B(new_n4058_), .Y(new_n4269_));
  AOI21X1  g04076(.A0(new_n4087_), .A1(new_n4031_), .B0(new_n4269_), .Y(new_n4270_));
  XOR2X1   g04077(.A(new_n4083_), .B(new_n4014_), .Y(new_n4271_));
  AND2X1   g04078(.A(\a[48] ), .B(\a[47] ), .Y(new_n4272_));
  AND2X1   g04079(.A(\a[49] ), .B(\a[47] ), .Y(new_n4273_));
  AND2X1   g04080(.A(\a[49] ), .B(\a[48] ), .Y(new_n4274_));
  AOI22X1  g04081(.A0(new_n4274_), .A1(new_n231_), .B0(new_n4273_), .B1(new_n235_), .Y(new_n4275_));
  AOI21X1  g04082(.A0(new_n4272_), .A1(new_n294_), .B0(new_n4275_), .Y(new_n4276_));
  AND2X1   g04083(.A(\a[49] ), .B(\a[2] ), .Y(new_n4277_));
  INVX1    g04084(.A(new_n4277_), .Y(new_n4278_));
  INVX1    g04085(.A(new_n4273_), .Y(new_n4279_));
  INVX1    g04086(.A(new_n4274_), .Y(new_n4280_));
  OAI22X1  g04087(.A0(new_n4280_), .A1(new_n249_), .B0(new_n4279_), .B1(new_n584_), .Y(new_n4281_));
  AOI21X1  g04088(.A0(new_n4272_), .A1(new_n294_), .B0(new_n4281_), .Y(new_n4282_));
  INVX1    g04089(.A(new_n4282_), .Y(new_n4283_));
  AOI22X1  g04090(.A0(\a[48] ), .A1(\a[3] ), .B0(\a[47] ), .B1(\a[4] ), .Y(new_n4284_));
  OAI22X1  g04091(.A0(new_n4284_), .A1(new_n4283_), .B0(new_n4278_), .B1(new_n4276_), .Y(new_n4285_));
  XOR2X1   g04092(.A(new_n4285_), .B(new_n4271_), .Y(new_n4286_));
  INVX1    g04093(.A(new_n4286_), .Y(new_n4287_));
  AND2X1   g04094(.A(new_n4027_), .B(new_n4017_), .Y(new_n4288_));
  AOI21X1  g04095(.A0(new_n4030_), .A1(new_n4028_), .B0(new_n4288_), .Y(new_n4289_));
  XOR2X1   g04096(.A(new_n4289_), .B(new_n4287_), .Y(new_n4290_));
  NOR2X1   g04097(.A(new_n4114_), .B(new_n4112_), .Y(new_n4291_));
  AOI21X1  g04098(.A0(new_n4117_), .A1(new_n4115_), .B0(new_n4291_), .Y(new_n4292_));
  XOR2X1   g04099(.A(new_n4292_), .B(new_n4290_), .Y(new_n4293_));
  XOR2X1   g04100(.A(new_n4293_), .B(new_n4270_), .Y(new_n4294_));
  XOR2X1   g04101(.A(new_n4073_), .B(new_n4063_), .Y(new_n4295_));
  XOR2X1   g04102(.A(new_n4295_), .B(new_n4025_), .Y(new_n4296_));
  AND2X1   g04103(.A(new_n4075_), .B(new_n4066_), .Y(new_n4297_));
  AOI21X1  g04104(.A0(new_n4085_), .A1(new_n4076_), .B0(new_n4297_), .Y(new_n4298_));
  XOR2X1   g04105(.A(new_n4298_), .B(new_n4296_), .Y(new_n4299_));
  INVX1    g04106(.A(new_n4037_), .Y(new_n4300_));
  XOR2X1   g04107(.A(new_n4054_), .B(new_n4047_), .Y(new_n4301_));
  XOR2X1   g04108(.A(new_n4301_), .B(new_n4300_), .Y(new_n4302_));
  XOR2X1   g04109(.A(new_n4302_), .B(new_n4299_), .Y(new_n4303_));
  XOR2X1   g04110(.A(new_n4303_), .B(new_n4294_), .Y(new_n4304_));
  XOR2X1   g04111(.A(new_n4304_), .B(new_n4268_), .Y(new_n4305_));
  XOR2X1   g04112(.A(new_n4305_), .B(new_n4250_), .Y(new_n4306_));
  AND2X1   g04113(.A(new_n4306_), .B(new_n4163_), .Y(new_n4307_));
  NOR2X1   g04114(.A(new_n4306_), .B(new_n4163_), .Y(new_n4308_));
  OR2X1    g04115(.A(new_n4308_), .B(new_n4307_), .Y(new_n4309_));
  XOR2X1   g04116(.A(new_n4309_), .B(new_n4160_), .Y(\asquared[52] ));
  AND2X1   g04117(.A(new_n4249_), .B(new_n4166_), .Y(new_n4311_));
  AOI21X1  g04118(.A0(new_n4305_), .A1(new_n4250_), .B0(new_n4311_), .Y(new_n4312_));
  NOR2X1   g04119(.A(new_n4247_), .B(new_n4170_), .Y(new_n4313_));
  AOI21X1  g04120(.A0(new_n4248_), .A1(new_n4168_), .B0(new_n4313_), .Y(new_n4314_));
  INVX1    g04121(.A(new_n4314_), .Y(new_n4315_));
  NOR2X1   g04122(.A(new_n4054_), .B(new_n4047_), .Y(new_n4316_));
  AOI21X1  g04123(.A0(new_n4301_), .A1(new_n4300_), .B0(new_n4316_), .Y(new_n4317_));
  AND2X1   g04124(.A(\a[33] ), .B(\a[19] ), .Y(new_n4318_));
  INVX1    g04125(.A(new_n4318_), .Y(new_n4319_));
  AOI22X1  g04126(.A0(\a[50] ), .A1(\a[2] ), .B0(\a[49] ), .B1(\a[3] ), .Y(new_n4320_));
  AND2X1   g04127(.A(\a[50] ), .B(\a[49] ), .Y(new_n4321_));
  AND2X1   g04128(.A(new_n4321_), .B(new_n231_), .Y(new_n4322_));
  NOR3X1   g04129(.A(new_n4320_), .B(new_n4322_), .C(new_n4319_), .Y(new_n4323_));
  INVX1    g04130(.A(new_n4320_), .Y(new_n4324_));
  AOI21X1  g04131(.A0(new_n4324_), .A1(new_n4318_), .B0(new_n4322_), .Y(new_n4325_));
  INVX1    g04132(.A(new_n4325_), .Y(new_n4326_));
  OAI22X1  g04133(.A0(new_n4326_), .A1(new_n4320_), .B0(new_n4323_), .B1(new_n4319_), .Y(new_n4327_));
  XOR2X1   g04134(.A(new_n4327_), .B(new_n4317_), .Y(new_n4328_));
  AND2X1   g04135(.A(new_n4073_), .B(new_n4063_), .Y(new_n4329_));
  AOI21X1  g04136(.A0(new_n4295_), .A1(new_n4026_), .B0(new_n4329_), .Y(new_n4330_));
  XOR2X1   g04137(.A(new_n4330_), .B(new_n4328_), .Y(new_n4331_));
  AND2X1   g04138(.A(new_n4289_), .B(new_n4287_), .Y(new_n4332_));
  OR2X1    g04139(.A(new_n4289_), .B(new_n4287_), .Y(new_n4333_));
  OAI21X1  g04140(.A0(new_n4292_), .A1(new_n4332_), .B0(new_n4333_), .Y(new_n4334_));
  XOR2X1   g04141(.A(new_n4334_), .B(new_n4331_), .Y(new_n4335_));
  AND2X1   g04142(.A(new_n4235_), .B(new_n4226_), .Y(new_n4336_));
  AOI21X1  g04143(.A0(new_n4244_), .A1(new_n4236_), .B0(new_n4336_), .Y(new_n4337_));
  AND2X1   g04144(.A(new_n4083_), .B(new_n4014_), .Y(new_n4338_));
  AOI21X1  g04145(.A0(new_n4285_), .A1(new_n4271_), .B0(new_n4338_), .Y(new_n4339_));
  AND2X1   g04146(.A(new_n4174_), .B(\a[26] ), .Y(new_n4340_));
  AND2X1   g04147(.A(\a[51] ), .B(\a[1] ), .Y(new_n4341_));
  XOR2X1   g04148(.A(new_n4341_), .B(new_n1871_), .Y(new_n4342_));
  XOR2X1   g04149(.A(new_n4342_), .B(new_n4340_), .Y(new_n4343_));
  XOR2X1   g04150(.A(new_n4343_), .B(new_n4243_), .Y(new_n4344_));
  XOR2X1   g04151(.A(new_n4344_), .B(new_n4339_), .Y(new_n4345_));
  XOR2X1   g04152(.A(new_n4345_), .B(new_n4337_), .Y(new_n4346_));
  XOR2X1   g04153(.A(new_n4346_), .B(new_n4335_), .Y(new_n4347_));
  XOR2X1   g04154(.A(new_n4347_), .B(new_n4315_), .Y(new_n4348_));
  INVX1    g04155(.A(\a[51] ), .Y(new_n4349_));
  NOR3X1   g04156(.A(new_n4171_), .B(new_n4349_), .C(new_n194_), .Y(new_n4350_));
  NOR2X1   g04157(.A(new_n4175_), .B(new_n4173_), .Y(new_n4351_));
  NOR2X1   g04158(.A(new_n4351_), .B(new_n4350_), .Y(new_n4352_));
  XOR2X1   g04159(.A(new_n4352_), .B(new_n4232_), .Y(new_n4353_));
  INVX1    g04160(.A(\a[52] ), .Y(new_n4354_));
  AOI22X1  g04161(.A0(new_n1433_), .A1(\a[35] ), .B0(new_n210_), .B1(\a[48] ), .Y(new_n4355_));
  NOR4X1   g04162(.A(new_n3926_), .B(new_n2557_), .C(new_n616_), .D(new_n340_), .Y(new_n4356_));
  NOR3X1   g04163(.A(new_n4356_), .B(new_n4355_), .C(new_n4354_), .Y(new_n4357_));
  NOR3X1   g04164(.A(new_n4357_), .B(new_n4354_), .C(new_n194_), .Y(new_n4358_));
  NOR2X1   g04165(.A(new_n4357_), .B(new_n4356_), .Y(new_n4359_));
  AOI22X1  g04166(.A0(\a[48] ), .A1(\a[4] ), .B0(\a[35] ), .B1(\a[17] ), .Y(new_n4360_));
  INVX1    g04167(.A(new_n4360_), .Y(new_n4361_));
  AOI21X1  g04168(.A0(new_n4361_), .A1(new_n4359_), .B0(new_n4358_), .Y(new_n4362_));
  XOR2X1   g04169(.A(new_n4362_), .B(new_n4353_), .Y(new_n4363_));
  INVX1    g04170(.A(new_n4363_), .Y(new_n4364_));
  INVX1    g04171(.A(new_n4176_), .Y(new_n4365_));
  OR2X1    g04172(.A(new_n4183_), .B(new_n4365_), .Y(new_n4366_));
  OAI21X1  g04173(.A0(new_n4186_), .A1(new_n4184_), .B0(new_n4366_), .Y(new_n4367_));
  XOR2X1   g04174(.A(new_n4367_), .B(new_n4364_), .Y(new_n4368_));
  INVX1    g04175(.A(new_n4368_), .Y(new_n4369_));
  AND2X1   g04176(.A(new_n4261_), .B(new_n4258_), .Y(new_n4370_));
  AOI21X1  g04177(.A0(new_n4265_), .A1(new_n4262_), .B0(new_n4370_), .Y(new_n4371_));
  XOR2X1   g04178(.A(new_n4371_), .B(new_n4369_), .Y(new_n4372_));
  XOR2X1   g04179(.A(new_n4216_), .B(new_n4204_), .Y(new_n4373_));
  INVX1    g04180(.A(new_n4187_), .Y(new_n4374_));
  NOR2X1   g04181(.A(new_n4246_), .B(new_n4374_), .Y(new_n4375_));
  AOI21X1  g04182(.A0(new_n4245_), .A1(new_n4373_), .B0(new_n4375_), .Y(new_n4376_));
  XOR2X1   g04183(.A(new_n4223_), .B(new_n4192_), .Y(new_n4377_));
  XOR2X1   g04184(.A(new_n4377_), .B(new_n4202_), .Y(new_n4378_));
  XOR2X1   g04185(.A(new_n4282_), .B(new_n4182_), .Y(new_n4379_));
  XOR2X1   g04186(.A(new_n4379_), .B(new_n4215_), .Y(new_n4380_));
  INVX1    g04187(.A(new_n4380_), .Y(new_n4381_));
  AND2X1   g04188(.A(new_n4203_), .B(new_n4195_), .Y(new_n4382_));
  AOI21X1  g04189(.A0(new_n4216_), .A1(new_n4204_), .B0(new_n4382_), .Y(new_n4383_));
  XOR2X1   g04190(.A(new_n4383_), .B(new_n4381_), .Y(new_n4384_));
  XOR2X1   g04191(.A(new_n4384_), .B(new_n4378_), .Y(new_n4385_));
  XOR2X1   g04192(.A(new_n4385_), .B(new_n4376_), .Y(new_n4386_));
  XOR2X1   g04193(.A(new_n4386_), .B(new_n4372_), .Y(new_n4387_));
  XOR2X1   g04194(.A(new_n4387_), .B(new_n4348_), .Y(new_n4388_));
  NOR2X1   g04195(.A(new_n4293_), .B(new_n4270_), .Y(new_n4389_));
  AOI21X1  g04196(.A0(new_n4303_), .A1(new_n4294_), .B0(new_n4389_), .Y(new_n4390_));
  NOR2X1   g04197(.A(new_n4255_), .B(new_n4253_), .Y(new_n4391_));
  AOI21X1  g04198(.A0(new_n4266_), .A1(new_n4256_), .B0(new_n4391_), .Y(new_n4392_));
  NOR2X1   g04199(.A(new_n4298_), .B(new_n4296_), .Y(new_n4393_));
  AOI21X1  g04200(.A0(new_n4302_), .A1(new_n4299_), .B0(new_n4393_), .Y(new_n4394_));
  NAND2X1  g04201(.A(\a[47] ), .B(\a[5] ), .Y(new_n4395_));
  NOR4X1   g04202(.A(new_n3460_), .B(new_n2583_), .C(new_n571_), .D(new_n230_), .Y(new_n4396_));
  NAND4X1  g04203(.A(\a[47] ), .B(\a[46] ), .C(\a[6] ), .D(\a[5] ), .Y(new_n4397_));
  NAND4X1  g04204(.A(\a[47] ), .B(\a[36] ), .C(\a[16] ), .D(\a[5] ), .Y(new_n4398_));
  AOI21X1  g04205(.A0(new_n4398_), .A1(new_n4397_), .B0(new_n4396_), .Y(new_n4399_));
  OR2X1    g04206(.A(new_n4399_), .B(new_n4396_), .Y(new_n4400_));
  AOI22X1  g04207(.A0(\a[46] ), .A1(\a[6] ), .B0(\a[36] ), .B1(\a[16] ), .Y(new_n4401_));
  OAI22X1  g04208(.A0(new_n4401_), .A1(new_n4400_), .B0(new_n4399_), .B1(new_n4395_), .Y(new_n4402_));
  NAND2X1  g04209(.A(\a[42] ), .B(\a[10] ), .Y(new_n4403_));
  AND2X1   g04210(.A(\a[41] ), .B(\a[40] ), .Y(new_n4404_));
  NAND4X1  g04211(.A(\a[42] ), .B(\a[40] ), .C(\a[12] ), .D(\a[10] ), .Y(new_n4405_));
  NAND4X1  g04212(.A(\a[42] ), .B(\a[41] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n4406_));
  AOI22X1  g04213(.A0(new_n4406_), .A1(new_n4405_), .B0(new_n4404_), .B1(new_n482_), .Y(new_n4407_));
  NAND4X1  g04214(.A(\a[41] ), .B(\a[40] ), .C(\a[12] ), .D(\a[11] ), .Y(new_n4408_));
  NAND3X1  g04215(.A(new_n4406_), .B(new_n4405_), .C(new_n4408_), .Y(new_n4409_));
  AOI22X1  g04216(.A0(\a[41] ), .A1(\a[11] ), .B0(\a[40] ), .B1(\a[12] ), .Y(new_n4410_));
  OAI22X1  g04217(.A0(new_n4410_), .A1(new_n4409_), .B0(new_n4407_), .B1(new_n4403_), .Y(new_n4411_));
  XOR2X1   g04218(.A(new_n4411_), .B(new_n4402_), .Y(new_n4412_));
  AND2X1   g04219(.A(\a[37] ), .B(\a[15] ), .Y(new_n4413_));
  INVX1    g04220(.A(new_n4413_), .Y(new_n4414_));
  AOI22X1  g04221(.A0(\a[45] ), .A1(\a[7] ), .B0(\a[44] ), .B1(\a[8] ), .Y(new_n4415_));
  AND2X1   g04222(.A(new_n3918_), .B(new_n325_), .Y(new_n4416_));
  NOR3X1   g04223(.A(new_n4415_), .B(new_n4416_), .C(new_n4414_), .Y(new_n4417_));
  NOR2X1   g04224(.A(new_n4417_), .B(new_n4416_), .Y(new_n4418_));
  INVX1    g04225(.A(new_n4418_), .Y(new_n4419_));
  OAI22X1  g04226(.A0(new_n4419_), .A1(new_n4415_), .B0(new_n4417_), .B1(new_n4414_), .Y(new_n4420_));
  XOR2X1   g04227(.A(new_n4420_), .B(new_n4412_), .Y(new_n4421_));
  INVX1    g04228(.A(new_n4421_), .Y(new_n4422_));
  NAND4X1  g04229(.A(\a[34] ), .B(\a[31] ), .C(\a[21] ), .D(\a[18] ), .Y(new_n4423_));
  NAND4X1  g04230(.A(\a[34] ), .B(\a[32] ), .C(\a[20] ), .D(\a[18] ), .Y(new_n4424_));
  AOI22X1  g04231(.A0(new_n4424_), .A1(new_n4423_), .B0(new_n2671_), .B1(new_n1236_), .Y(new_n4425_));
  NAND4X1  g04232(.A(\a[32] ), .B(\a[31] ), .C(\a[21] ), .D(\a[20] ), .Y(new_n4426_));
  NAND3X1  g04233(.A(new_n4424_), .B(new_n4423_), .C(new_n4426_), .Y(new_n4427_));
  AOI22X1  g04234(.A0(\a[32] ), .A1(\a[20] ), .B0(\a[31] ), .B1(\a[21] ), .Y(new_n4428_));
  NAND2X1  g04235(.A(\a[34] ), .B(\a[18] ), .Y(new_n4429_));
  OAI22X1  g04236(.A0(new_n4429_), .A1(new_n4425_), .B0(new_n4428_), .B1(new_n4427_), .Y(new_n4430_));
  NAND4X1  g04237(.A(\a[30] ), .B(\a[28] ), .C(\a[24] ), .D(\a[22] ), .Y(new_n4431_));
  NAND4X1  g04238(.A(\a[30] ), .B(\a[29] ), .C(\a[23] ), .D(\a[22] ), .Y(new_n4432_));
  AOI22X1  g04239(.A0(new_n4432_), .A1(new_n4431_), .B0(new_n1674_), .B1(new_n1219_), .Y(new_n4433_));
  NAND2X1  g04240(.A(\a[30] ), .B(\a[22] ), .Y(new_n4434_));
  AOI22X1  g04241(.A0(\a[29] ), .A1(\a[23] ), .B0(\a[28] ), .B1(\a[24] ), .Y(new_n4435_));
  AOI21X1  g04242(.A0(new_n1674_), .A1(new_n1219_), .B0(new_n4433_), .Y(new_n4436_));
  INVX1    g04243(.A(new_n4436_), .Y(new_n4437_));
  OAI22X1  g04244(.A0(new_n4437_), .A1(new_n4435_), .B0(new_n4434_), .B1(new_n4433_), .Y(new_n4438_));
  XOR2X1   g04245(.A(new_n4438_), .B(new_n4430_), .Y(new_n4439_));
  AND2X1   g04246(.A(\a[38] ), .B(\a[14] ), .Y(new_n4440_));
  NOR4X1   g04247(.A(new_n3037_), .B(new_n2652_), .C(new_n591_), .D(new_n341_), .Y(new_n4441_));
  AND2X1   g04248(.A(\a[43] ), .B(\a[9] ), .Y(new_n4442_));
  AOI22X1  g04249(.A0(new_n4442_), .A1(new_n4440_), .B0(new_n3503_), .B1(new_n582_), .Y(new_n4443_));
  OAI21X1  g04250(.A0(new_n4443_), .A1(new_n4441_), .B0(new_n4440_), .Y(new_n4444_));
  INVX1    g04251(.A(new_n4441_), .Y(new_n4445_));
  AND2X1   g04252(.A(new_n4443_), .B(new_n4445_), .Y(new_n4446_));
  AND2X1   g04253(.A(\a[39] ), .B(\a[13] ), .Y(new_n4447_));
  OAI21X1  g04254(.A0(new_n4447_), .A1(new_n4442_), .B0(new_n4446_), .Y(new_n4448_));
  AND2X1   g04255(.A(new_n4448_), .B(new_n4444_), .Y(new_n4449_));
  XOR2X1   g04256(.A(new_n4449_), .B(new_n4439_), .Y(new_n4450_));
  XOR2X1   g04257(.A(new_n4450_), .B(new_n4422_), .Y(new_n4451_));
  INVX1    g04258(.A(new_n4451_), .Y(new_n4452_));
  XOR2X1   g04259(.A(new_n4452_), .B(new_n4394_), .Y(new_n4453_));
  INVX1    g04260(.A(new_n4453_), .Y(new_n4454_));
  XOR2X1   g04261(.A(new_n4454_), .B(new_n4392_), .Y(new_n4455_));
  XOR2X1   g04262(.A(new_n4455_), .B(new_n4390_), .Y(new_n4456_));
  AND2X1   g04263(.A(new_n4267_), .B(new_n4251_), .Y(new_n4457_));
  AOI21X1  g04264(.A0(new_n4304_), .A1(new_n4268_), .B0(new_n4457_), .Y(new_n4458_));
  XOR2X1   g04265(.A(new_n4458_), .B(new_n4456_), .Y(new_n4459_));
  XOR2X1   g04266(.A(new_n4459_), .B(new_n4388_), .Y(new_n4460_));
  NOR2X1   g04267(.A(new_n4460_), .B(new_n4312_), .Y(new_n4461_));
  INVX1    g04268(.A(new_n4461_), .Y(new_n4462_));
  INVX1    g04269(.A(new_n4307_), .Y(new_n4463_));
  OAI21X1  g04270(.A0(new_n4308_), .A1(new_n4160_), .B0(new_n4463_), .Y(new_n4464_));
  AND2X1   g04271(.A(new_n4460_), .B(new_n4312_), .Y(new_n4465_));
  INVX1    g04272(.A(new_n4465_), .Y(new_n4466_));
  AOI21X1  g04273(.A0(new_n4462_), .A1(new_n4466_), .B0(new_n4464_), .Y(new_n4467_));
  AND2X1   g04274(.A(new_n4466_), .B(new_n4464_), .Y(new_n4468_));
  AOI21X1  g04275(.A0(new_n4468_), .A1(new_n4462_), .B0(new_n4467_), .Y(\asquared[53] ));
  AOI21X1  g04276(.A0(new_n4466_), .A1(new_n4464_), .B0(new_n4461_), .Y(new_n4470_));
  OR2X1    g04277(.A(new_n4458_), .B(new_n4456_), .Y(new_n4471_));
  AND2X1   g04278(.A(new_n4458_), .B(new_n4456_), .Y(new_n4472_));
  OAI21X1  g04279(.A0(new_n4472_), .A1(new_n4388_), .B0(new_n4471_), .Y(new_n4473_));
  NOR2X1   g04280(.A(new_n4347_), .B(new_n4315_), .Y(new_n4474_));
  NAND2X1  g04281(.A(new_n4347_), .B(new_n4315_), .Y(new_n4475_));
  OAI21X1  g04282(.A0(new_n4387_), .A1(new_n4474_), .B0(new_n4475_), .Y(new_n4476_));
  INVX1    g04283(.A(new_n4372_), .Y(new_n4477_));
  AND2X1   g04284(.A(new_n4245_), .B(new_n4373_), .Y(new_n4478_));
  OAI21X1  g04285(.A0(new_n4478_), .A1(new_n4375_), .B0(new_n4385_), .Y(new_n4479_));
  OAI21X1  g04286(.A0(new_n4386_), .A1(new_n4477_), .B0(new_n4479_), .Y(new_n4480_));
  AOI22X1  g04287(.A0(\a[51] ), .A1(\a[2] ), .B0(\a[50] ), .B1(\a[3] ), .Y(new_n4481_));
  INVX1    g04288(.A(new_n4481_), .Y(new_n4482_));
  AND2X1   g04289(.A(new_n4341_), .B(new_n1871_), .Y(new_n4483_));
  AND2X1   g04290(.A(\a[51] ), .B(\a[50] ), .Y(new_n4484_));
  AND2X1   g04291(.A(new_n4484_), .B(new_n231_), .Y(new_n4485_));
  AOI21X1  g04292(.A0(new_n4482_), .A1(new_n4483_), .B0(new_n4485_), .Y(new_n4486_));
  NAND2X1  g04293(.A(new_n4486_), .B(new_n4482_), .Y(new_n4487_));
  OAI21X1  g04294(.A0(new_n4485_), .A1(new_n4481_), .B0(new_n4483_), .Y(new_n4488_));
  AND2X1   g04295(.A(new_n4488_), .B(new_n4487_), .Y(new_n4489_));
  AND2X1   g04296(.A(\a[49] ), .B(\a[4] ), .Y(new_n4490_));
  AOI22X1  g04297(.A0(\a[36] ), .A1(\a[17] ), .B0(\a[35] ), .B1(\a[18] ), .Y(new_n4491_));
  INVX1    g04298(.A(new_n4491_), .Y(new_n4492_));
  NAND4X1  g04299(.A(\a[36] ), .B(\a[35] ), .C(\a[18] ), .D(\a[17] ), .Y(new_n4493_));
  NAND3X1  g04300(.A(new_n4492_), .B(new_n4493_), .C(new_n4490_), .Y(new_n4494_));
  AOI22X1  g04301(.A0(new_n4492_), .A1(new_n4490_), .B0(new_n2682_), .B1(new_n796_), .Y(new_n4495_));
  AOI22X1  g04302(.A0(new_n4495_), .A1(new_n4492_), .B0(new_n4494_), .B1(new_n4490_), .Y(new_n4496_));
  XOR2X1   g04303(.A(new_n4496_), .B(new_n4489_), .Y(new_n4497_));
  OAI22X1  g04304(.A0(new_n2919_), .A1(new_n1521_), .B0(new_n2920_), .B1(new_n1149_), .Y(new_n4498_));
  OAI21X1  g04305(.A0(new_n2675_), .A1(new_n1794_), .B0(new_n4498_), .Y(new_n4499_));
  AND2X1   g04306(.A(\a[34] ), .B(\a[19] ), .Y(new_n4500_));
  AOI21X1  g04307(.A0(new_n2674_), .A1(new_n1236_), .B0(new_n4498_), .Y(new_n4501_));
  OAI22X1  g04308(.A0(new_n1851_), .A1(new_n934_), .B0(new_n2219_), .B1(new_n1098_), .Y(new_n4502_));
  AOI22X1  g04309(.A0(new_n4502_), .A1(new_n4501_), .B0(new_n4500_), .B1(new_n4499_), .Y(new_n4503_));
  XOR2X1   g04310(.A(new_n4503_), .B(new_n4497_), .Y(new_n4504_));
  INVX1    g04311(.A(new_n4327_), .Y(new_n4505_));
  OR2X1    g04312(.A(new_n4505_), .B(new_n4317_), .Y(new_n4506_));
  OAI21X1  g04313(.A0(new_n4330_), .A1(new_n4328_), .B0(new_n4506_), .Y(new_n4507_));
  XOR2X1   g04314(.A(new_n4507_), .B(new_n4504_), .Y(new_n4508_));
  NAND2X1  g04315(.A(\a[47] ), .B(\a[6] ), .Y(new_n4509_));
  NOR4X1   g04316(.A(new_n3460_), .B(new_n2519_), .C(new_n549_), .D(new_n532_), .Y(new_n4510_));
  NAND4X1  g04317(.A(\a[47] ), .B(\a[46] ), .C(\a[7] ), .D(\a[6] ), .Y(new_n4511_));
  NAND4X1  g04318(.A(\a[47] ), .B(\a[38] ), .C(\a[15] ), .D(\a[6] ), .Y(new_n4512_));
  AOI21X1  g04319(.A0(new_n4512_), .A1(new_n4511_), .B0(new_n4510_), .Y(new_n4513_));
  OR2X1    g04320(.A(new_n4513_), .B(new_n4510_), .Y(new_n4514_));
  AOI22X1  g04321(.A0(\a[46] ), .A1(\a[7] ), .B0(\a[38] ), .B1(\a[15] ), .Y(new_n4515_));
  OAI22X1  g04322(.A0(new_n4515_), .A1(new_n4514_), .B0(new_n4513_), .B1(new_n4509_), .Y(new_n4516_));
  NAND2X1  g04323(.A(\a[45] ), .B(\a[8] ), .Y(new_n4517_));
  NAND2X1  g04324(.A(\a[44] ), .B(\a[14] ), .Y(new_n4518_));
  NOR3X1   g04325(.A(new_n4518_), .B(new_n2652_), .C(new_n341_), .Y(new_n4519_));
  NAND4X1  g04326(.A(\a[45] ), .B(\a[44] ), .C(\a[9] ), .D(\a[8] ), .Y(new_n4520_));
  NAND4X1  g04327(.A(\a[45] ), .B(\a[39] ), .C(\a[14] ), .D(\a[8] ), .Y(new_n4521_));
  AOI21X1  g04328(.A0(new_n4521_), .A1(new_n4520_), .B0(new_n4519_), .Y(new_n4522_));
  OR2X1    g04329(.A(new_n4522_), .B(new_n4519_), .Y(new_n4523_));
  AOI22X1  g04330(.A0(\a[44] ), .A1(\a[9] ), .B0(\a[39] ), .B1(\a[14] ), .Y(new_n4524_));
  OAI22X1  g04331(.A0(new_n4524_), .A1(new_n4523_), .B0(new_n4522_), .B1(new_n4517_), .Y(new_n4525_));
  XOR2X1   g04332(.A(new_n4525_), .B(new_n4516_), .Y(new_n4526_));
  AND2X1   g04333(.A(\a[53] ), .B(\a[0] ), .Y(new_n4527_));
  INVX1    g04334(.A(new_n4527_), .Y(new_n4528_));
  AOI22X1  g04335(.A0(\a[48] ), .A1(\a[5] ), .B0(\a[37] ), .B1(\a[16] ), .Y(new_n4529_));
  NOR4X1   g04336(.A(new_n3926_), .B(new_n2345_), .C(new_n571_), .D(new_n255_), .Y(new_n4530_));
  NOR3X1   g04337(.A(new_n4529_), .B(new_n4530_), .C(new_n4528_), .Y(new_n4531_));
  NOR2X1   g04338(.A(new_n4531_), .B(new_n4530_), .Y(new_n4532_));
  INVX1    g04339(.A(new_n4532_), .Y(new_n4533_));
  OAI22X1  g04340(.A0(new_n4533_), .A1(new_n4529_), .B0(new_n4531_), .B1(new_n4528_), .Y(new_n4534_));
  INVX1    g04341(.A(new_n4534_), .Y(new_n4535_));
  XOR2X1   g04342(.A(new_n4535_), .B(new_n4526_), .Y(new_n4536_));
  XOR2X1   g04343(.A(new_n4536_), .B(new_n4508_), .Y(new_n4537_));
  AOI22X1  g04344(.A0(\a[43] ), .A1(\a[10] ), .B0(\a[41] ), .B1(\a[12] ), .Y(new_n4538_));
  NAND4X1  g04345(.A(\a[43] ), .B(\a[40] ), .C(\a[13] ), .D(\a[10] ), .Y(new_n4539_));
  NAND4X1  g04346(.A(\a[41] ), .B(\a[40] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n4540_));
  AOI22X1  g04347(.A0(new_n4540_), .A1(new_n4539_), .B0(new_n3320_), .B1(new_n396_), .Y(new_n4541_));
  AOI21X1  g04348(.A0(new_n3320_), .A1(new_n396_), .B0(new_n4541_), .Y(new_n4542_));
  INVX1    g04349(.A(new_n4542_), .Y(new_n4543_));
  NAND2X1  g04350(.A(\a[40] ), .B(\a[13] ), .Y(new_n4544_));
  OAI22X1  g04351(.A0(new_n4544_), .A1(new_n4541_), .B0(new_n4543_), .B1(new_n4538_), .Y(new_n4545_));
  NAND4X1  g04352(.A(\a[31] ), .B(\a[29] ), .C(\a[24] ), .D(\a[22] ), .Y(new_n4546_));
  NAND4X1  g04353(.A(\a[31] ), .B(\a[30] ), .C(\a[23] ), .D(\a[22] ), .Y(new_n4547_));
  AOI22X1  g04354(.A0(new_n4547_), .A1(new_n4546_), .B0(new_n2196_), .B1(new_n1219_), .Y(new_n4548_));
  AOI22X1  g04355(.A0(\a[30] ), .A1(\a[23] ), .B0(\a[29] ), .B1(\a[24] ), .Y(new_n4549_));
  AOI21X1  g04356(.A0(new_n2196_), .A1(new_n1219_), .B0(new_n4548_), .Y(new_n4550_));
  INVX1    g04357(.A(new_n4550_), .Y(new_n4551_));
  OAI22X1  g04358(.A0(new_n4551_), .A1(new_n4549_), .B0(new_n4548_), .B1(new_n1697_), .Y(new_n4552_));
  XOR2X1   g04359(.A(new_n4552_), .B(new_n4545_), .Y(new_n4553_));
  NAND2X1  g04360(.A(\a[42] ), .B(\a[11] ), .Y(new_n4554_));
  AOI22X1  g04361(.A0(\a[28] ), .A1(\a[25] ), .B0(\a[27] ), .B1(\a[26] ), .Y(new_n4555_));
  AND2X1   g04362(.A(new_n1770_), .B(new_n1671_), .Y(new_n4556_));
  NOR3X1   g04363(.A(new_n4555_), .B(new_n4556_), .C(new_n4554_), .Y(new_n4557_));
  OAI22X1  g04364(.A0(new_n4555_), .A1(new_n4554_), .B0(new_n1771_), .B1(new_n1672_), .Y(new_n4558_));
  OAI22X1  g04365(.A0(new_n4558_), .A1(new_n4555_), .B0(new_n4557_), .B1(new_n4554_), .Y(new_n4559_));
  XOR2X1   g04366(.A(new_n4559_), .B(new_n4553_), .Y(new_n4560_));
  INVX1    g04367(.A(new_n4344_), .Y(new_n4561_));
  OR2X1    g04368(.A(new_n4561_), .B(new_n4339_), .Y(new_n4562_));
  OAI21X1  g04369(.A0(new_n4345_), .A1(new_n4337_), .B0(new_n4562_), .Y(new_n4563_));
  XOR2X1   g04370(.A(new_n4563_), .B(new_n4560_), .Y(new_n4564_));
  NAND2X1  g04371(.A(new_n4384_), .B(new_n4378_), .Y(new_n4565_));
  OAI21X1  g04372(.A0(new_n4383_), .A1(new_n4381_), .B0(new_n4565_), .Y(new_n4566_));
  XOR2X1   g04373(.A(new_n4566_), .B(new_n4564_), .Y(new_n4567_));
  XOR2X1   g04374(.A(new_n4567_), .B(new_n4537_), .Y(new_n4568_));
  XOR2X1   g04375(.A(new_n4568_), .B(new_n4480_), .Y(new_n4569_));
  XOR2X1   g04376(.A(new_n4569_), .B(new_n4476_), .Y(new_n4570_));
  XOR2X1   g04377(.A(new_n4359_), .B(new_n4325_), .Y(new_n4571_));
  XOR2X1   g04378(.A(new_n4571_), .B(new_n4437_), .Y(new_n4572_));
  AND2X1   g04379(.A(new_n4438_), .B(new_n4430_), .Y(new_n4573_));
  INVX1    g04380(.A(new_n4449_), .Y(new_n4574_));
  AOI21X1  g04381(.A0(new_n4574_), .A1(new_n4439_), .B0(new_n4573_), .Y(new_n4575_));
  NOR2X1   g04382(.A(new_n4352_), .B(new_n4232_), .Y(new_n4576_));
  INVX1    g04383(.A(new_n4362_), .Y(new_n4577_));
  AOI21X1  g04384(.A0(new_n4577_), .A1(new_n4353_), .B0(new_n4576_), .Y(new_n4578_));
  XOR2X1   g04385(.A(new_n4578_), .B(new_n4575_), .Y(new_n4579_));
  XOR2X1   g04386(.A(new_n4579_), .B(new_n4572_), .Y(new_n4580_));
  XOR2X1   g04387(.A(new_n4427_), .B(new_n4400_), .Y(new_n4581_));
  XOR2X1   g04388(.A(new_n4581_), .B(new_n4419_), .Y(new_n4582_));
  AND2X1   g04389(.A(new_n4411_), .B(new_n4402_), .Y(new_n4583_));
  AOI21X1  g04390(.A0(new_n4420_), .A1(new_n4412_), .B0(new_n4583_), .Y(new_n4584_));
  AOI21X1  g04391(.A0(\a[52] ), .A1(\a[1] ), .B0(\a[27] ), .Y(new_n4585_));
  AOI21X1  g04392(.A0(new_n1413_), .A1(\a[52] ), .B0(new_n4585_), .Y(new_n4586_));
  XOR2X1   g04393(.A(new_n4586_), .B(new_n4409_), .Y(new_n4587_));
  INVX1    g04394(.A(new_n4587_), .Y(new_n4588_));
  XOR2X1   g04395(.A(new_n4588_), .B(new_n4446_), .Y(new_n4589_));
  XOR2X1   g04396(.A(new_n4589_), .B(new_n4584_), .Y(new_n4590_));
  XOR2X1   g04397(.A(new_n4590_), .B(new_n4582_), .Y(new_n4591_));
  XOR2X1   g04398(.A(new_n4591_), .B(new_n4580_), .Y(new_n4592_));
  AND2X1   g04399(.A(new_n4334_), .B(new_n4331_), .Y(new_n4593_));
  AOI21X1  g04400(.A0(new_n4346_), .A1(new_n4335_), .B0(new_n4593_), .Y(new_n4594_));
  XOR2X1   g04401(.A(new_n4594_), .B(new_n4592_), .Y(new_n4595_));
  OR2X1    g04402(.A(new_n4450_), .B(new_n4422_), .Y(new_n4596_));
  OAI21X1  g04403(.A0(new_n4452_), .A1(new_n4394_), .B0(new_n4596_), .Y(new_n4597_));
  AND2X1   g04404(.A(new_n4223_), .B(new_n4192_), .Y(new_n4598_));
  AOI21X1  g04405(.A0(new_n4377_), .A1(new_n4202_), .B0(new_n4598_), .Y(new_n4599_));
  AND2X1   g04406(.A(new_n4342_), .B(new_n4340_), .Y(new_n4600_));
  AOI21X1  g04407(.A0(new_n4343_), .A1(new_n4243_), .B0(new_n4600_), .Y(new_n4601_));
  INVX1    g04408(.A(new_n4601_), .Y(new_n4602_));
  XOR2X1   g04409(.A(new_n4602_), .B(new_n4599_), .Y(new_n4603_));
  NOR2X1   g04410(.A(new_n4282_), .B(new_n4182_), .Y(new_n4604_));
  AOI21X1  g04411(.A0(new_n4379_), .A1(new_n4215_), .B0(new_n4604_), .Y(new_n4605_));
  XOR2X1   g04412(.A(new_n4605_), .B(new_n4603_), .Y(new_n4606_));
  NAND2X1  g04413(.A(new_n4367_), .B(new_n4364_), .Y(new_n4607_));
  OAI21X1  g04414(.A0(new_n4371_), .A1(new_n4369_), .B0(new_n4607_), .Y(new_n4608_));
  XOR2X1   g04415(.A(new_n4608_), .B(new_n4606_), .Y(new_n4609_));
  XOR2X1   g04416(.A(new_n4609_), .B(new_n4597_), .Y(new_n4610_));
  OR2X1    g04417(.A(new_n4454_), .B(new_n4392_), .Y(new_n4611_));
  AND2X1   g04418(.A(new_n4454_), .B(new_n4392_), .Y(new_n4612_));
  OAI21X1  g04419(.A0(new_n4612_), .A1(new_n4390_), .B0(new_n4611_), .Y(new_n4613_));
  XOR2X1   g04420(.A(new_n4613_), .B(new_n4610_), .Y(new_n4614_));
  XOR2X1   g04421(.A(new_n4614_), .B(new_n4595_), .Y(new_n4615_));
  XOR2X1   g04422(.A(new_n4615_), .B(new_n4570_), .Y(new_n4616_));
  AND2X1   g04423(.A(new_n4616_), .B(new_n4473_), .Y(new_n4617_));
  NOR2X1   g04424(.A(new_n4616_), .B(new_n4473_), .Y(new_n4618_));
  OR2X1    g04425(.A(new_n4618_), .B(new_n4617_), .Y(new_n4619_));
  XOR2X1   g04426(.A(new_n4619_), .B(new_n4470_), .Y(\asquared[54] ));
  AND2X1   g04427(.A(new_n4569_), .B(new_n4476_), .Y(new_n4621_));
  AND2X1   g04428(.A(new_n4615_), .B(new_n4570_), .Y(new_n4622_));
  OR2X1    g04429(.A(new_n4622_), .B(new_n4621_), .Y(new_n4623_));
  INVX1    g04430(.A(new_n4591_), .Y(new_n4624_));
  NOR2X1   g04431(.A(new_n4594_), .B(new_n4592_), .Y(new_n4625_));
  AOI21X1  g04432(.A0(new_n4624_), .A1(new_n4580_), .B0(new_n4625_), .Y(new_n4626_));
  AND2X1   g04433(.A(new_n4608_), .B(new_n4606_), .Y(new_n4627_));
  AOI21X1  g04434(.A0(new_n4609_), .A1(new_n4597_), .B0(new_n4627_), .Y(new_n4628_));
  XOR2X1   g04435(.A(new_n4628_), .B(new_n4626_), .Y(new_n4629_));
  INVX1    g04436(.A(new_n4582_), .Y(new_n4630_));
  INVX1    g04437(.A(new_n4589_), .Y(new_n4631_));
  OR2X1    g04438(.A(new_n4631_), .B(new_n4584_), .Y(new_n4632_));
  OAI21X1  g04439(.A0(new_n4590_), .A1(new_n4630_), .B0(new_n4632_), .Y(new_n4633_));
  NOR2X1   g04440(.A(new_n4578_), .B(new_n4575_), .Y(new_n4634_));
  AOI21X1  g04441(.A0(new_n4579_), .A1(new_n4572_), .B0(new_n4634_), .Y(new_n4635_));
  NAND3X1  g04442(.A(\a[52] ), .B(\a[27] ), .C(\a[1] ), .Y(new_n4636_));
  AND2X1   g04443(.A(\a[54] ), .B(\a[0] ), .Y(new_n4637_));
  XOR2X1   g04444(.A(new_n4637_), .B(new_n4636_), .Y(new_n4638_));
  NAND2X1  g04445(.A(\a[53] ), .B(\a[1] ), .Y(new_n4639_));
  XOR2X1   g04446(.A(new_n4639_), .B(new_n1996_), .Y(new_n4640_));
  XOR2X1   g04447(.A(new_n4640_), .B(new_n4638_), .Y(new_n4641_));
  NAND4X1  g04448(.A(\a[35] ), .B(\a[32] ), .C(\a[22] ), .D(\a[19] ), .Y(new_n4642_));
  NAND4X1  g04449(.A(\a[35] ), .B(\a[33] ), .C(\a[21] ), .D(\a[19] ), .Y(new_n4643_));
  AOI22X1  g04450(.A0(new_n4643_), .A1(new_n4642_), .B0(new_n2674_), .B1(new_n1154_), .Y(new_n4644_));
  NAND4X1  g04451(.A(\a[33] ), .B(\a[32] ), .C(\a[22] ), .D(\a[21] ), .Y(new_n4645_));
  NAND3X1  g04452(.A(new_n4643_), .B(new_n4642_), .C(new_n4645_), .Y(new_n4646_));
  AOI22X1  g04453(.A0(\a[33] ), .A1(\a[21] ), .B0(\a[32] ), .B1(\a[22] ), .Y(new_n4647_));
  NAND2X1  g04454(.A(\a[35] ), .B(\a[19] ), .Y(new_n4648_));
  OAI22X1  g04455(.A0(new_n4648_), .A1(new_n4644_), .B0(new_n4647_), .B1(new_n4646_), .Y(new_n4649_));
  NAND4X1  g04456(.A(\a[31] ), .B(\a[29] ), .C(\a[25] ), .D(\a[23] ), .Y(new_n4650_));
  NAND4X1  g04457(.A(\a[31] ), .B(\a[30] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n4651_));
  AOI22X1  g04458(.A0(new_n4651_), .A1(new_n4650_), .B0(new_n2196_), .B1(new_n1532_), .Y(new_n4652_));
  NAND2X1  g04459(.A(\a[31] ), .B(\a[23] ), .Y(new_n4653_));
  NAND4X1  g04460(.A(\a[30] ), .B(\a[29] ), .C(\a[25] ), .D(\a[24] ), .Y(new_n4654_));
  NAND3X1  g04461(.A(new_n4651_), .B(new_n4650_), .C(new_n4654_), .Y(new_n4655_));
  AOI22X1  g04462(.A0(\a[30] ), .A1(\a[24] ), .B0(\a[29] ), .B1(\a[25] ), .Y(new_n4656_));
  OAI22X1  g04463(.A0(new_n4656_), .A1(new_n4655_), .B0(new_n4653_), .B1(new_n4652_), .Y(new_n4657_));
  XOR2X1   g04464(.A(new_n4657_), .B(new_n4649_), .Y(new_n4658_));
  XOR2X1   g04465(.A(new_n4658_), .B(new_n4641_), .Y(new_n4659_));
  XOR2X1   g04466(.A(new_n4659_), .B(new_n4635_), .Y(new_n4660_));
  XOR2X1   g04467(.A(new_n4660_), .B(new_n4633_), .Y(new_n4661_));
  XOR2X1   g04468(.A(new_n4661_), .B(new_n4629_), .Y(new_n4662_));
  AND2X1   g04469(.A(new_n4613_), .B(new_n4610_), .Y(new_n4663_));
  AOI21X1  g04470(.A0(new_n4614_), .A1(new_n4595_), .B0(new_n4663_), .Y(new_n4664_));
  XOR2X1   g04471(.A(new_n4664_), .B(new_n4662_), .Y(new_n4665_));
  AND2X1   g04472(.A(new_n4567_), .B(new_n4537_), .Y(new_n4666_));
  AOI21X1  g04473(.A0(new_n4568_), .A1(new_n4480_), .B0(new_n4666_), .Y(new_n4667_));
  INVX1    g04474(.A(new_n4667_), .Y(new_n4668_));
  AND2X1   g04475(.A(new_n4427_), .B(new_n4400_), .Y(new_n4669_));
  AOI21X1  g04476(.A0(new_n4581_), .A1(new_n4419_), .B0(new_n4669_), .Y(new_n4670_));
  NOR2X1   g04477(.A(new_n4359_), .B(new_n4325_), .Y(new_n4671_));
  AOI21X1  g04478(.A0(new_n4571_), .A1(new_n4437_), .B0(new_n4671_), .Y(new_n4672_));
  XOR2X1   g04479(.A(new_n4672_), .B(new_n4670_), .Y(new_n4673_));
  AND2X1   g04480(.A(new_n4586_), .B(new_n4409_), .Y(new_n4674_));
  INVX1    g04481(.A(new_n4674_), .Y(new_n4675_));
  OAI21X1  g04482(.A0(new_n4588_), .A1(new_n4446_), .B0(new_n4675_), .Y(new_n4676_));
  INVX1    g04483(.A(new_n4676_), .Y(new_n4677_));
  XOR2X1   g04484(.A(new_n4677_), .B(new_n4673_), .Y(new_n4678_));
  INVX1    g04485(.A(new_n4504_), .Y(new_n4679_));
  NOR2X1   g04486(.A(new_n4536_), .B(new_n4508_), .Y(new_n4680_));
  AOI21X1  g04487(.A0(new_n4507_), .A1(new_n4679_), .B0(new_n4680_), .Y(new_n4681_));
  XOR2X1   g04488(.A(new_n4681_), .B(new_n4678_), .Y(new_n4682_));
  XOR2X1   g04489(.A(new_n4533_), .B(new_n4514_), .Y(new_n4683_));
  XOR2X1   g04490(.A(new_n4683_), .B(new_n4558_), .Y(new_n4684_));
  XOR2X1   g04491(.A(new_n4501_), .B(new_n4495_), .Y(new_n4685_));
  XOR2X1   g04492(.A(new_n4685_), .B(new_n4550_), .Y(new_n4686_));
  AND2X1   g04493(.A(new_n4525_), .B(new_n4516_), .Y(new_n4687_));
  AOI21X1  g04494(.A0(new_n4534_), .A1(new_n4526_), .B0(new_n4687_), .Y(new_n4688_));
  XOR2X1   g04495(.A(new_n4688_), .B(new_n4686_), .Y(new_n4689_));
  XOR2X1   g04496(.A(new_n4689_), .B(new_n4684_), .Y(new_n4690_));
  XOR2X1   g04497(.A(new_n4690_), .B(new_n4682_), .Y(new_n4691_));
  XOR2X1   g04498(.A(new_n4691_), .B(new_n4668_), .Y(new_n4692_));
  AOI22X1  g04499(.A0(\a[49] ), .A1(\a[5] ), .B0(\a[36] ), .B1(\a[18] ), .Y(new_n4693_));
  NOR4X1   g04500(.A(new_n3915_), .B(new_n2583_), .C(new_n675_), .D(new_n255_), .Y(new_n4694_));
  AND2X1   g04501(.A(\a[36] ), .B(\a[34] ), .Y(new_n4695_));
  AND2X1   g04502(.A(\a[49] ), .B(\a[20] ), .Y(new_n4696_));
  AOI22X1  g04503(.A0(new_n4696_), .A1(new_n2573_), .B0(new_n4695_), .B1(new_n992_), .Y(new_n4697_));
  NOR2X1   g04504(.A(new_n4697_), .B(new_n4694_), .Y(new_n4698_));
  INVX1    g04505(.A(new_n4694_), .Y(new_n4699_));
  AND2X1   g04506(.A(new_n4697_), .B(new_n4699_), .Y(new_n4700_));
  INVX1    g04507(.A(new_n4700_), .Y(new_n4701_));
  NAND2X1  g04508(.A(\a[34] ), .B(\a[20] ), .Y(new_n4702_));
  OAI22X1  g04509(.A0(new_n4702_), .A1(new_n4698_), .B0(new_n4701_), .B1(new_n4693_), .Y(new_n4703_));
  NAND4X1  g04510(.A(\a[43] ), .B(\a[41] ), .C(\a[13] ), .D(\a[11] ), .Y(new_n4704_));
  NAND4X1  g04511(.A(\a[42] ), .B(\a[41] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n4705_));
  AOI22X1  g04512(.A0(new_n4705_), .A1(new_n4704_), .B0(new_n3462_), .B1(new_n482_), .Y(new_n4706_));
  NAND2X1  g04513(.A(\a[41] ), .B(\a[13] ), .Y(new_n4707_));
  AOI21X1  g04514(.A0(new_n3462_), .A1(new_n482_), .B0(new_n4706_), .Y(new_n4708_));
  INVX1    g04515(.A(new_n4708_), .Y(new_n4709_));
  AOI22X1  g04516(.A0(\a[43] ), .A1(\a[11] ), .B0(\a[42] ), .B1(\a[12] ), .Y(new_n4710_));
  OAI22X1  g04517(.A0(new_n4710_), .A1(new_n4709_), .B0(new_n4707_), .B1(new_n4706_), .Y(new_n4711_));
  XOR2X1   g04518(.A(new_n4711_), .B(new_n4703_), .Y(new_n4712_));
  AND2X1   g04519(.A(\a[48] ), .B(\a[38] ), .Y(new_n4713_));
  NAND4X1  g04520(.A(\a[48] ), .B(\a[37] ), .C(\a[17] ), .D(\a[6] ), .Y(new_n4714_));
  NAND4X1  g04521(.A(\a[38] ), .B(\a[37] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n4715_));
  AOI22X1  g04522(.A0(new_n4715_), .A1(new_n4714_), .B0(new_n4713_), .B1(new_n564_), .Y(new_n4716_));
  AND2X1   g04523(.A(\a[37] ), .B(\a[17] ), .Y(new_n4717_));
  INVX1    g04524(.A(new_n4717_), .Y(new_n4718_));
  AOI22X1  g04525(.A0(\a[48] ), .A1(\a[6] ), .B0(\a[38] ), .B1(\a[16] ), .Y(new_n4719_));
  AOI21X1  g04526(.A0(new_n4713_), .A1(new_n564_), .B0(new_n4716_), .Y(new_n4720_));
  INVX1    g04527(.A(new_n4720_), .Y(new_n4721_));
  OAI22X1  g04528(.A0(new_n4721_), .A1(new_n4719_), .B0(new_n4718_), .B1(new_n4716_), .Y(new_n4722_));
  XOR2X1   g04529(.A(new_n4722_), .B(new_n4712_), .Y(new_n4723_));
  INVX1    g04530(.A(new_n4723_), .Y(new_n4724_));
  OR2X1    g04531(.A(new_n4601_), .B(new_n4599_), .Y(new_n4725_));
  OAI21X1  g04532(.A0(new_n4605_), .A1(new_n4603_), .B0(new_n4725_), .Y(new_n4726_));
  XOR2X1   g04533(.A(new_n4726_), .B(new_n4724_), .Y(new_n4727_));
  NAND4X1  g04534(.A(\a[52] ), .B(\a[50] ), .C(\a[4] ), .D(\a[2] ), .Y(new_n4728_));
  NAND4X1  g04535(.A(\a[52] ), .B(\a[51] ), .C(\a[3] ), .D(\a[2] ), .Y(new_n4729_));
  AOI22X1  g04536(.A0(new_n4729_), .A1(new_n4728_), .B0(new_n4484_), .B1(new_n294_), .Y(new_n4730_));
  NAND4X1  g04537(.A(\a[51] ), .B(\a[50] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n4731_));
  NAND3X1  g04538(.A(new_n4729_), .B(new_n4728_), .C(new_n4731_), .Y(new_n4732_));
  AOI22X1  g04539(.A0(\a[51] ), .A1(\a[3] ), .B0(\a[50] ), .B1(\a[4] ), .Y(new_n4733_));
  NAND2X1  g04540(.A(\a[52] ), .B(\a[2] ), .Y(new_n4734_));
  OAI22X1  g04541(.A0(new_n4734_), .A1(new_n4730_), .B0(new_n4733_), .B1(new_n4732_), .Y(new_n4735_));
  AND2X1   g04542(.A(\a[47] ), .B(\a[7] ), .Y(new_n4736_));
  AND2X1   g04543(.A(\a[39] ), .B(\a[15] ), .Y(new_n4737_));
  AOI22X1  g04544(.A0(new_n4737_), .A1(new_n4736_), .B0(new_n3893_), .B1(new_n325_), .Y(new_n4738_));
  NOR4X1   g04545(.A(new_n3460_), .B(new_n2652_), .C(new_n549_), .D(new_n413_), .Y(new_n4739_));
  OAI21X1  g04546(.A0(new_n4739_), .A1(new_n4738_), .B0(new_n4736_), .Y(new_n4740_));
  INVX1    g04547(.A(new_n4739_), .Y(new_n4741_));
  AND2X1   g04548(.A(new_n4741_), .B(new_n4738_), .Y(new_n4742_));
  INVX1    g04549(.A(new_n4742_), .Y(new_n4743_));
  AOI22X1  g04550(.A0(\a[46] ), .A1(\a[8] ), .B0(\a[39] ), .B1(\a[15] ), .Y(new_n4744_));
  OAI21X1  g04551(.A0(new_n4744_), .A1(new_n4743_), .B0(new_n4740_), .Y(new_n4745_));
  XOR2X1   g04552(.A(new_n4745_), .B(new_n4735_), .Y(new_n4746_));
  AND2X1   g04553(.A(\a[45] ), .B(\a[9] ), .Y(new_n4747_));
  NOR3X1   g04554(.A(new_n4518_), .B(new_n3036_), .C(new_n570_), .Y(new_n4748_));
  AOI22X1  g04555(.A0(new_n4747_), .A1(new_n3351_), .B0(new_n3918_), .B1(new_n881_), .Y(new_n4749_));
  OAI21X1  g04556(.A0(new_n4749_), .A1(new_n4748_), .B0(new_n4747_), .Y(new_n4750_));
  INVX1    g04557(.A(new_n4748_), .Y(new_n4751_));
  AND2X1   g04558(.A(new_n4749_), .B(new_n4751_), .Y(new_n4752_));
  INVX1    g04559(.A(new_n4752_), .Y(new_n4753_));
  AOI22X1  g04560(.A0(\a[44] ), .A1(\a[10] ), .B0(\a[40] ), .B1(\a[14] ), .Y(new_n4754_));
  OAI21X1  g04561(.A0(new_n4754_), .A1(new_n4753_), .B0(new_n4750_), .Y(new_n4755_));
  INVX1    g04562(.A(new_n4755_), .Y(new_n4756_));
  XOR2X1   g04563(.A(new_n4756_), .B(new_n4746_), .Y(new_n4757_));
  XOR2X1   g04564(.A(new_n4757_), .B(new_n4727_), .Y(new_n4758_));
  AND2X1   g04565(.A(new_n4563_), .B(new_n4560_), .Y(new_n4759_));
  AOI21X1  g04566(.A0(new_n4566_), .A1(new_n4564_), .B0(new_n4759_), .Y(new_n4760_));
  INVX1    g04567(.A(new_n4486_), .Y(new_n4761_));
  XOR2X1   g04568(.A(new_n4523_), .B(new_n4761_), .Y(new_n4762_));
  XOR2X1   g04569(.A(new_n4762_), .B(new_n4543_), .Y(new_n4763_));
  INVX1    g04570(.A(new_n4763_), .Y(new_n4764_));
  AND2X1   g04571(.A(new_n4552_), .B(new_n4545_), .Y(new_n4765_));
  AND2X1   g04572(.A(new_n4559_), .B(new_n4553_), .Y(new_n4766_));
  OR2X1    g04573(.A(new_n4766_), .B(new_n4765_), .Y(new_n4767_));
  OR2X1    g04574(.A(new_n4496_), .B(new_n4489_), .Y(new_n4768_));
  INVX1    g04575(.A(new_n4497_), .Y(new_n4769_));
  OAI21X1  g04576(.A0(new_n4503_), .A1(new_n4769_), .B0(new_n4768_), .Y(new_n4770_));
  XOR2X1   g04577(.A(new_n4770_), .B(new_n4767_), .Y(new_n4771_));
  XOR2X1   g04578(.A(new_n4771_), .B(new_n4764_), .Y(new_n4772_));
  XOR2X1   g04579(.A(new_n4772_), .B(new_n4760_), .Y(new_n4773_));
  XOR2X1   g04580(.A(new_n4773_), .B(new_n4758_), .Y(new_n4774_));
  XOR2X1   g04581(.A(new_n4774_), .B(new_n4692_), .Y(new_n4775_));
  XOR2X1   g04582(.A(new_n4775_), .B(new_n4665_), .Y(new_n4776_));
  XOR2X1   g04583(.A(new_n4776_), .B(new_n4623_), .Y(new_n4777_));
  INVX1    g04584(.A(new_n4617_), .Y(new_n4778_));
  OAI21X1  g04585(.A0(new_n4618_), .A1(new_n4470_), .B0(new_n4778_), .Y(new_n4779_));
  XOR2X1   g04586(.A(new_n4779_), .B(new_n4777_), .Y(\asquared[55] ));
  NOR2X1   g04587(.A(new_n4664_), .B(new_n4662_), .Y(new_n4781_));
  AOI21X1  g04588(.A0(new_n4775_), .A1(new_n4665_), .B0(new_n4781_), .Y(new_n4782_));
  AND2X1   g04589(.A(new_n4691_), .B(new_n4668_), .Y(new_n4783_));
  AOI21X1  g04590(.A0(new_n4774_), .A1(new_n4692_), .B0(new_n4783_), .Y(new_n4784_));
  NOR2X1   g04591(.A(new_n4772_), .B(new_n4760_), .Y(new_n4785_));
  AOI21X1  g04592(.A0(new_n4773_), .A1(new_n4758_), .B0(new_n4785_), .Y(new_n4786_));
  NOR2X1   g04593(.A(new_n4681_), .B(new_n4678_), .Y(new_n4787_));
  AOI21X1  g04594(.A0(new_n4690_), .A1(new_n4682_), .B0(new_n4787_), .Y(new_n4788_));
  NOR2X1   g04595(.A(new_n4688_), .B(new_n4686_), .Y(new_n4789_));
  AOI21X1  g04596(.A0(new_n4689_), .A1(new_n4684_), .B0(new_n4789_), .Y(new_n4790_));
  AOI22X1  g04597(.A0(\a[49] ), .A1(\a[6] ), .B0(\a[38] ), .B1(\a[17] ), .Y(new_n4791_));
  AND2X1   g04598(.A(\a[52] ), .B(\a[3] ), .Y(new_n4792_));
  INVX1    g04599(.A(new_n4792_), .Y(new_n4793_));
  NOR4X1   g04600(.A(new_n3915_), .B(new_n2519_), .C(new_n616_), .D(new_n230_), .Y(new_n4794_));
  NOR3X1   g04601(.A(new_n4793_), .B(new_n4794_), .C(new_n4791_), .Y(new_n4795_));
  NOR2X1   g04602(.A(new_n4795_), .B(new_n4794_), .Y(new_n4796_));
  INVX1    g04603(.A(new_n4796_), .Y(new_n4797_));
  OAI22X1  g04604(.A0(new_n4797_), .A1(new_n4791_), .B0(new_n4795_), .B1(new_n4793_), .Y(new_n4798_));
  NOR4X1   g04605(.A(new_n3460_), .B(new_n3036_), .C(new_n549_), .D(new_n341_), .Y(new_n4799_));
  AOI21X1  g04606(.A0(new_n4404_), .A1(new_n691_), .B0(new_n4799_), .Y(new_n4800_));
  NOR4X1   g04607(.A(new_n3460_), .B(new_n3081_), .C(new_n490_), .D(new_n341_), .Y(new_n4801_));
  OR2X1    g04608(.A(new_n4801_), .B(new_n4800_), .Y(new_n4802_));
  AND2X1   g04609(.A(\a[40] ), .B(\a[15] ), .Y(new_n4803_));
  OAI22X1  g04610(.A0(new_n3460_), .A1(new_n341_), .B0(new_n3081_), .B1(new_n490_), .Y(new_n4804_));
  AND2X1   g04611(.A(new_n4404_), .B(new_n691_), .Y(new_n4805_));
  NOR3X1   g04612(.A(new_n4801_), .B(new_n4805_), .C(new_n4799_), .Y(new_n4806_));
  AOI22X1  g04613(.A0(new_n4806_), .A1(new_n4804_), .B0(new_n4803_), .B1(new_n4802_), .Y(new_n4807_));
  XOR2X1   g04614(.A(new_n4807_), .B(new_n4798_), .Y(new_n4808_));
  NOR2X1   g04615(.A(new_n4501_), .B(new_n4495_), .Y(new_n4809_));
  AOI21X1  g04616(.A0(new_n4685_), .A1(new_n4551_), .B0(new_n4809_), .Y(new_n4810_));
  XOR2X1   g04617(.A(new_n4810_), .B(new_n4808_), .Y(new_n4811_));
  AND2X1   g04618(.A(new_n4770_), .B(new_n4767_), .Y(new_n4812_));
  AOI21X1  g04619(.A0(new_n4771_), .A1(new_n4763_), .B0(new_n4812_), .Y(new_n4813_));
  XOR2X1   g04620(.A(new_n4813_), .B(new_n4811_), .Y(new_n4814_));
  XOR2X1   g04621(.A(new_n4814_), .B(new_n4790_), .Y(new_n4815_));
  XOR2X1   g04622(.A(new_n4815_), .B(new_n4788_), .Y(new_n4816_));
  XOR2X1   g04623(.A(new_n4816_), .B(new_n4786_), .Y(new_n4817_));
  XOR2X1   g04624(.A(new_n4817_), .B(new_n4784_), .Y(new_n4818_));
  INVX1    g04625(.A(new_n4818_), .Y(new_n4819_));
  AND2X1   g04626(.A(new_n4533_), .B(new_n4514_), .Y(new_n4820_));
  AOI21X1  g04627(.A0(new_n4683_), .A1(new_n4558_), .B0(new_n4820_), .Y(new_n4821_));
  AND2X1   g04628(.A(new_n4523_), .B(new_n4761_), .Y(new_n4822_));
  AOI21X1  g04629(.A0(new_n4762_), .A1(new_n4543_), .B0(new_n4822_), .Y(new_n4823_));
  XOR2X1   g04630(.A(new_n4823_), .B(new_n4821_), .Y(new_n4824_));
  NAND4X1  g04631(.A(\a[53] ), .B(\a[28] ), .C(\a[26] ), .D(\a[1] ), .Y(new_n4825_));
  AND2X1   g04632(.A(\a[54] ), .B(\a[28] ), .Y(new_n4826_));
  AOI21X1  g04633(.A0(\a[54] ), .A1(\a[1] ), .B0(\a[28] ), .Y(new_n4827_));
  AOI21X1  g04634(.A0(new_n4826_), .A1(\a[1] ), .B0(new_n4827_), .Y(new_n4828_));
  XOR2X1   g04635(.A(new_n4828_), .B(new_n4825_), .Y(new_n4829_));
  XOR2X1   g04636(.A(new_n4829_), .B(new_n4708_), .Y(new_n4830_));
  XOR2X1   g04637(.A(new_n4830_), .B(new_n4824_), .Y(new_n4831_));
  NAND2X1  g04638(.A(new_n4726_), .B(new_n4723_), .Y(new_n4832_));
  OAI21X1  g04639(.A0(new_n4757_), .A1(new_n4727_), .B0(new_n4832_), .Y(new_n4833_));
  XOR2X1   g04640(.A(new_n4833_), .B(new_n4831_), .Y(new_n4834_));
  INVX1    g04641(.A(\a[54] ), .Y(new_n4835_));
  NOR3X1   g04642(.A(new_n4636_), .B(new_n4835_), .C(new_n194_), .Y(new_n4836_));
  NOR2X1   g04643(.A(new_n4640_), .B(new_n4638_), .Y(new_n4837_));
  NOR2X1   g04644(.A(new_n4837_), .B(new_n4836_), .Y(new_n4838_));
  XOR2X1   g04645(.A(new_n4838_), .B(new_n4742_), .Y(new_n4839_));
  AND2X1   g04646(.A(\a[50] ), .B(\a[5] ), .Y(new_n4840_));
  INVX1    g04647(.A(new_n4840_), .Y(new_n4841_));
  AND2X1   g04648(.A(new_n3330_), .B(new_n855_), .Y(new_n4842_));
  AOI22X1  g04649(.A0(\a[37] ), .A1(\a[18] ), .B0(\a[36] ), .B1(\a[19] ), .Y(new_n4843_));
  NOR3X1   g04650(.A(new_n4843_), .B(new_n4842_), .C(new_n4841_), .Y(new_n4844_));
  INVX1    g04651(.A(new_n4843_), .Y(new_n4845_));
  AOI21X1  g04652(.A0(new_n4845_), .A1(new_n4840_), .B0(new_n4842_), .Y(new_n4846_));
  NAND2X1  g04653(.A(new_n4846_), .B(new_n4845_), .Y(new_n4847_));
  OAI21X1  g04654(.A0(new_n4844_), .A1(new_n4841_), .B0(new_n4847_), .Y(new_n4848_));
  XOR2X1   g04655(.A(new_n4848_), .B(new_n4839_), .Y(new_n4849_));
  XOR2X1   g04656(.A(new_n4753_), .B(new_n4732_), .Y(new_n4850_));
  XOR2X1   g04657(.A(new_n4850_), .B(new_n4700_), .Y(new_n4851_));
  AND2X1   g04658(.A(new_n4657_), .B(new_n4649_), .Y(new_n4852_));
  AOI21X1  g04659(.A0(new_n4658_), .A1(new_n4641_), .B0(new_n4852_), .Y(new_n4853_));
  XOR2X1   g04660(.A(new_n4853_), .B(new_n4851_), .Y(new_n4854_));
  XOR2X1   g04661(.A(new_n4854_), .B(new_n4849_), .Y(new_n4855_));
  XOR2X1   g04662(.A(new_n4855_), .B(new_n4834_), .Y(new_n4856_));
  NOR2X1   g04663(.A(new_n4628_), .B(new_n4626_), .Y(new_n4857_));
  INVX1    g04664(.A(new_n4661_), .Y(new_n4858_));
  AOI21X1  g04665(.A0(new_n4858_), .A1(new_n4629_), .B0(new_n4857_), .Y(new_n4859_));
  XOR2X1   g04666(.A(new_n4859_), .B(new_n4856_), .Y(new_n4860_));
  INVX1    g04667(.A(new_n4659_), .Y(new_n4861_));
  OR2X1    g04668(.A(new_n4861_), .B(new_n4635_), .Y(new_n4862_));
  INVX1    g04669(.A(new_n4660_), .Y(new_n4863_));
  NAND2X1  g04670(.A(new_n4863_), .B(new_n4633_), .Y(new_n4864_));
  AND2X1   g04671(.A(new_n4864_), .B(new_n4862_), .Y(new_n4865_));
  XOR2X1   g04672(.A(new_n4655_), .B(new_n4646_), .Y(new_n4866_));
  XOR2X1   g04673(.A(new_n4866_), .B(new_n4721_), .Y(new_n4867_));
  INVX1    g04674(.A(new_n4867_), .Y(new_n4868_));
  AND2X1   g04675(.A(new_n4711_), .B(new_n4703_), .Y(new_n4869_));
  AOI21X1  g04676(.A0(new_n4722_), .A1(new_n4712_), .B0(new_n4869_), .Y(new_n4870_));
  AND2X1   g04677(.A(new_n4745_), .B(new_n4735_), .Y(new_n4871_));
  AOI21X1  g04678(.A0(new_n4755_), .A1(new_n4746_), .B0(new_n4871_), .Y(new_n4872_));
  XOR2X1   g04679(.A(new_n4872_), .B(new_n4870_), .Y(new_n4873_));
  XOR2X1   g04680(.A(new_n4873_), .B(new_n4868_), .Y(new_n4874_));
  XOR2X1   g04681(.A(new_n4874_), .B(new_n4865_), .Y(new_n4875_));
  INVX1    g04682(.A(new_n4875_), .Y(new_n4876_));
  NAND4X1  g04683(.A(\a[45] ), .B(\a[44] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n4877_));
  NAND4X1  g04684(.A(\a[45] ), .B(\a[42] ), .C(\a[13] ), .D(\a[10] ), .Y(new_n4878_));
  AOI22X1  g04685(.A0(new_n4878_), .A1(new_n4877_), .B0(new_n3208_), .B1(new_n634_), .Y(new_n4879_));
  AOI21X1  g04686(.A0(new_n3208_), .A1(new_n634_), .B0(new_n4879_), .Y(new_n4880_));
  AOI22X1  g04687(.A0(\a[44] ), .A1(\a[11] ), .B0(\a[42] ), .B1(\a[13] ), .Y(new_n4881_));
  INVX1    g04688(.A(new_n4881_), .Y(new_n4882_));
  NOR3X1   g04689(.A(new_n4879_), .B(new_n3811_), .C(new_n570_), .Y(new_n4883_));
  AOI21X1  g04690(.A0(new_n4882_), .A1(new_n4880_), .B0(new_n4883_), .Y(new_n4884_));
  NAND2X1  g04691(.A(\a[43] ), .B(\a[12] ), .Y(new_n4885_));
  AOI22X1  g04692(.A0(\a[29] ), .A1(\a[26] ), .B0(\a[28] ), .B1(\a[27] ), .Y(new_n4886_));
  NOR4X1   g04693(.A(new_n1803_), .B(new_n1431_), .C(new_n1679_), .D(new_n1263_), .Y(new_n4887_));
  NOR3X1   g04694(.A(new_n4886_), .B(new_n4887_), .C(new_n4885_), .Y(new_n4888_));
  OR2X1    g04695(.A(new_n4888_), .B(new_n4887_), .Y(new_n4889_));
  OAI22X1  g04696(.A0(new_n4889_), .A1(new_n4886_), .B0(new_n4888_), .B1(new_n4885_), .Y(new_n4890_));
  XOR2X1   g04697(.A(new_n4890_), .B(new_n4884_), .Y(new_n4891_));
  AND2X1   g04698(.A(\a[39] ), .B(\a[16] ), .Y(new_n4892_));
  AOI22X1  g04699(.A0(\a[48] ), .A1(\a[7] ), .B0(\a[47] ), .B1(\a[8] ), .Y(new_n4893_));
  INVX1    g04700(.A(new_n4893_), .Y(new_n4894_));
  NAND4X1  g04701(.A(\a[48] ), .B(\a[47] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n4895_));
  NAND3X1  g04702(.A(new_n4894_), .B(new_n4895_), .C(new_n4892_), .Y(new_n4896_));
  AOI22X1  g04703(.A0(new_n4894_), .A1(new_n4892_), .B0(new_n4272_), .B1(new_n325_), .Y(new_n4897_));
  AOI22X1  g04704(.A0(new_n4897_), .A1(new_n4894_), .B0(new_n4896_), .B1(new_n4892_), .Y(new_n4898_));
  XOR2X1   g04705(.A(new_n4898_), .B(new_n4891_), .Y(new_n4899_));
  INVX1    g04706(.A(new_n4899_), .Y(new_n4900_));
  NAND2X1  g04707(.A(new_n4676_), .B(new_n4673_), .Y(new_n4901_));
  OAI21X1  g04708(.A0(new_n4672_), .A1(new_n4670_), .B0(new_n4901_), .Y(new_n4902_));
  XOR2X1   g04709(.A(new_n4902_), .B(new_n4900_), .Y(new_n4903_));
  AND2X1   g04710(.A(\a[53] ), .B(\a[51] ), .Y(new_n4904_));
  AND2X1   g04711(.A(new_n4904_), .B(new_n235_), .Y(new_n4905_));
  INVX1    g04712(.A(\a[55] ), .Y(new_n4906_));
  AOI22X1  g04713(.A0(new_n210_), .A1(\a[51] ), .B0(new_n197_), .B1(\a[53] ), .Y(new_n4907_));
  NOR3X1   g04714(.A(new_n4907_), .B(new_n4905_), .C(new_n4906_), .Y(new_n4908_));
  NOR2X1   g04715(.A(new_n4908_), .B(new_n4905_), .Y(new_n4909_));
  AOI22X1  g04716(.A0(\a[53] ), .A1(\a[2] ), .B0(\a[51] ), .B1(\a[4] ), .Y(new_n4910_));
  INVX1    g04717(.A(new_n4910_), .Y(new_n4911_));
  NOR3X1   g04718(.A(new_n4908_), .B(new_n4906_), .C(new_n194_), .Y(new_n4912_));
  AOI21X1  g04719(.A0(new_n4911_), .A1(new_n4909_), .B0(new_n4912_), .Y(new_n4913_));
  INVX1    g04720(.A(new_n2120_), .Y(new_n4914_));
  INVX1    g04721(.A(new_n2361_), .Y(new_n4915_));
  OAI22X1  g04722(.A0(new_n4915_), .A1(new_n1794_), .B0(new_n4914_), .B1(new_n2135_), .Y(new_n4916_));
  OAI21X1  g04723(.A0(new_n2919_), .A1(new_n1397_), .B0(new_n4916_), .Y(new_n4917_));
  AND2X1   g04724(.A(\a[35] ), .B(\a[20] ), .Y(new_n4918_));
  AOI21X1  g04725(.A0(new_n2918_), .A1(new_n1154_), .B0(new_n4916_), .Y(new_n4919_));
  OAI22X1  g04726(.A0(new_n2028_), .A1(new_n1098_), .B0(new_n1851_), .B1(new_n1086_), .Y(new_n4920_));
  AOI22X1  g04727(.A0(new_n4920_), .A1(new_n4919_), .B0(new_n4918_), .B1(new_n4917_), .Y(new_n4921_));
  XOR2X1   g04728(.A(new_n4921_), .B(new_n4913_), .Y(new_n4922_));
  INVX1    g04729(.A(new_n1787_), .Y(new_n4923_));
  OAI22X1  g04730(.A0(new_n2672_), .A1(new_n1652_), .B0(new_n4923_), .B1(new_n2706_), .Y(new_n4924_));
  OAI21X1  g04731(.A0(new_n2076_), .A1(new_n1772_), .B0(new_n4924_), .Y(new_n4925_));
  AND2X1   g04732(.A(\a[32] ), .B(\a[23] ), .Y(new_n4926_));
  AOI21X1  g04733(.A0(new_n2075_), .A1(new_n1532_), .B0(new_n4924_), .Y(new_n4927_));
  OAI22X1  g04734(.A0(new_n1704_), .A1(new_n1185_), .B0(new_n1684_), .B1(new_n1326_), .Y(new_n4928_));
  AOI22X1  g04735(.A0(new_n4928_), .A1(new_n4927_), .B0(new_n4926_), .B1(new_n4925_), .Y(new_n4929_));
  XOR2X1   g04736(.A(new_n4929_), .B(new_n4922_), .Y(new_n4930_));
  XOR2X1   g04737(.A(new_n4930_), .B(new_n4903_), .Y(new_n4931_));
  XOR2X1   g04738(.A(new_n4931_), .B(new_n4876_), .Y(new_n4932_));
  XOR2X1   g04739(.A(new_n4932_), .B(new_n4860_), .Y(new_n4933_));
  XOR2X1   g04740(.A(new_n4933_), .B(new_n4819_), .Y(new_n4934_));
  XOR2X1   g04741(.A(new_n4934_), .B(new_n4782_), .Y(new_n4935_));
  AND2X1   g04742(.A(new_n4776_), .B(new_n4623_), .Y(new_n4936_));
  NOR3X1   g04743(.A(new_n4776_), .B(new_n4622_), .C(new_n4621_), .Y(new_n4937_));
  INVX1    g04744(.A(new_n4937_), .Y(new_n4938_));
  AOI21X1  g04745(.A0(new_n4779_), .A1(new_n4938_), .B0(new_n4936_), .Y(new_n4939_));
  XOR2X1   g04746(.A(new_n4939_), .B(new_n4935_), .Y(\asquared[56] ));
  INVX1    g04747(.A(new_n4817_), .Y(new_n4941_));
  NOR2X1   g04748(.A(new_n4941_), .B(new_n4784_), .Y(new_n4942_));
  AOI21X1  g04749(.A0(new_n4933_), .A1(new_n4819_), .B0(new_n4942_), .Y(new_n4943_));
  INVX1    g04750(.A(new_n4943_), .Y(new_n4944_));
  NOR2X1   g04751(.A(new_n4853_), .B(new_n4851_), .Y(new_n4945_));
  AOI21X1  g04752(.A0(new_n4854_), .A1(new_n4849_), .B0(new_n4945_), .Y(new_n4946_));
  NAND4X1  g04753(.A(new_n4828_), .B(new_n1996_), .C(\a[53] ), .D(\a[1] ), .Y(new_n4947_));
  OAI21X1  g04754(.A0(new_n4829_), .A1(new_n4708_), .B0(new_n4947_), .Y(new_n4948_));
  AOI22X1  g04755(.A0(\a[51] ), .A1(\a[5] ), .B0(\a[38] ), .B1(\a[18] ), .Y(new_n4949_));
  AND2X1   g04756(.A(\a[35] ), .B(\a[21] ), .Y(new_n4950_));
  NOR4X1   g04757(.A(new_n4349_), .B(new_n2519_), .C(new_n675_), .D(new_n255_), .Y(new_n4951_));
  OAI21X1  g04758(.A0(new_n4949_), .A1(new_n4951_), .B0(new_n4950_), .Y(new_n4952_));
  INVX1    g04759(.A(new_n4949_), .Y(new_n4953_));
  AOI21X1  g04760(.A0(new_n4953_), .A1(new_n4950_), .B0(new_n4951_), .Y(new_n4954_));
  INVX1    g04761(.A(new_n4954_), .Y(new_n4955_));
  OAI21X1  g04762(.A0(new_n4955_), .A1(new_n4949_), .B0(new_n4952_), .Y(new_n4956_));
  XOR2X1   g04763(.A(new_n4956_), .B(new_n4948_), .Y(new_n4957_));
  INVX1    g04764(.A(new_n4957_), .Y(new_n4958_));
  AND2X1   g04765(.A(new_n4753_), .B(new_n4732_), .Y(new_n4959_));
  AOI21X1  g04766(.A0(new_n4850_), .A1(new_n4701_), .B0(new_n4959_), .Y(new_n4960_));
  XOR2X1   g04767(.A(new_n4960_), .B(new_n4958_), .Y(new_n4961_));
  INVX1    g04768(.A(new_n4961_), .Y(new_n4962_));
  NOR2X1   g04769(.A(new_n4872_), .B(new_n4870_), .Y(new_n4963_));
  AOI21X1  g04770(.A0(new_n4873_), .A1(new_n4867_), .B0(new_n4963_), .Y(new_n4964_));
  XOR2X1   g04771(.A(new_n4964_), .B(new_n4962_), .Y(new_n4965_));
  INVX1    g04772(.A(new_n4965_), .Y(new_n4966_));
  XOR2X1   g04773(.A(new_n4966_), .B(new_n4946_), .Y(new_n4967_));
  INVX1    g04774(.A(new_n4967_), .Y(new_n4968_));
  AND2X1   g04775(.A(new_n4833_), .B(new_n4831_), .Y(new_n4969_));
  AOI21X1  g04776(.A0(new_n4855_), .A1(new_n4834_), .B0(new_n4969_), .Y(new_n4970_));
  XOR2X1   g04777(.A(new_n4970_), .B(new_n4968_), .Y(new_n4971_));
  INVX1    g04778(.A(new_n4971_), .Y(new_n4972_));
  AOI21X1  g04779(.A0(new_n4864_), .A1(new_n4862_), .B0(new_n4874_), .Y(new_n4973_));
  AOI21X1  g04780(.A0(new_n4931_), .A1(new_n4875_), .B0(new_n4973_), .Y(new_n4974_));
  XOR2X1   g04781(.A(new_n4974_), .B(new_n4972_), .Y(new_n4975_));
  INVX1    g04782(.A(new_n4856_), .Y(new_n4976_));
  OR2X1    g04783(.A(new_n4859_), .B(new_n4976_), .Y(new_n4977_));
  OR2X1    g04784(.A(new_n4932_), .B(new_n4860_), .Y(new_n4978_));
  AND2X1   g04785(.A(new_n4978_), .B(new_n4977_), .Y(new_n4979_));
  OR2X1    g04786(.A(new_n4979_), .B(new_n4975_), .Y(new_n4980_));
  AOI22X1  g04787(.A0(\a[49] ), .A1(\a[7] ), .B0(\a[39] ), .B1(\a[17] ), .Y(new_n4981_));
  NOR4X1   g04788(.A(new_n3915_), .B(new_n2652_), .C(new_n616_), .D(new_n532_), .Y(new_n4982_));
  INVX1    g04789(.A(\a[50] ), .Y(new_n4983_));
  NOR4X1   g04790(.A(new_n4983_), .B(new_n2652_), .C(new_n616_), .D(new_n230_), .Y(new_n4984_));
  AOI21X1  g04791(.A0(new_n4321_), .A1(new_n375_), .B0(new_n4984_), .Y(new_n4985_));
  NOR2X1   g04792(.A(new_n4985_), .B(new_n4982_), .Y(new_n4986_));
  INVX1    g04793(.A(new_n4982_), .Y(new_n4987_));
  AND2X1   g04794(.A(new_n4985_), .B(new_n4987_), .Y(new_n4988_));
  INVX1    g04795(.A(new_n4988_), .Y(new_n4989_));
  NAND2X1  g04796(.A(\a[50] ), .B(\a[6] ), .Y(new_n4990_));
  OAI22X1  g04797(.A0(new_n4990_), .A1(new_n4986_), .B0(new_n4989_), .B1(new_n4981_), .Y(new_n4991_));
  AND2X1   g04798(.A(\a[44] ), .B(\a[43] ), .Y(new_n4992_));
  NAND4X1  g04799(.A(\a[45] ), .B(\a[43] ), .C(\a[13] ), .D(\a[11] ), .Y(new_n4993_));
  NAND4X1  g04800(.A(\a[45] ), .B(\a[44] ), .C(\a[12] ), .D(\a[11] ), .Y(new_n4994_));
  AOI22X1  g04801(.A0(new_n4994_), .A1(new_n4993_), .B0(new_n4992_), .B1(new_n586_), .Y(new_n4995_));
  NAND2X1  g04802(.A(\a[45] ), .B(\a[11] ), .Y(new_n4996_));
  AOI22X1  g04803(.A0(\a[44] ), .A1(\a[12] ), .B0(\a[43] ), .B1(\a[13] ), .Y(new_n4997_));
  AOI21X1  g04804(.A0(new_n4992_), .A1(new_n586_), .B0(new_n4995_), .Y(new_n4998_));
  INVX1    g04805(.A(new_n4998_), .Y(new_n4999_));
  OAI22X1  g04806(.A0(new_n4999_), .A1(new_n4997_), .B0(new_n4996_), .B1(new_n4995_), .Y(new_n5000_));
  XOR2X1   g04807(.A(new_n5000_), .B(new_n4991_), .Y(new_n5001_));
  AND2X1   g04808(.A(\a[40] ), .B(\a[16] ), .Y(new_n5002_));
  NOR4X1   g04809(.A(new_n3926_), .B(new_n3081_), .C(new_n549_), .D(new_n413_), .Y(new_n5003_));
  AND2X1   g04810(.A(\a[48] ), .B(\a[40] ), .Y(new_n5004_));
  AOI22X1  g04811(.A0(new_n5004_), .A1(new_n1110_), .B0(new_n4404_), .B1(new_n689_), .Y(new_n5005_));
  OAI21X1  g04812(.A0(new_n5005_), .A1(new_n5003_), .B0(new_n5002_), .Y(new_n5006_));
  INVX1    g04813(.A(new_n5003_), .Y(new_n5007_));
  AND2X1   g04814(.A(new_n5005_), .B(new_n5007_), .Y(new_n5008_));
  INVX1    g04815(.A(new_n5008_), .Y(new_n5009_));
  AOI22X1  g04816(.A0(\a[48] ), .A1(\a[8] ), .B0(\a[41] ), .B1(\a[15] ), .Y(new_n5010_));
  OAI21X1  g04817(.A0(new_n5010_), .A1(new_n5009_), .B0(new_n5006_), .Y(new_n5011_));
  INVX1    g04818(.A(new_n5011_), .Y(new_n5012_));
  XOR2X1   g04819(.A(new_n5012_), .B(new_n5001_), .Y(new_n5013_));
  AND2X1   g04820(.A(new_n4695_), .B(new_n2134_), .Y(new_n5014_));
  NOR4X1   g04821(.A(new_n2583_), .B(new_n1851_), .C(new_n1216_), .D(new_n934_), .Y(new_n5015_));
  OAI22X1  g04822(.A0(new_n5015_), .A1(new_n5014_), .B0(new_n2919_), .B1(new_n1395_), .Y(new_n5016_));
  OAI21X1  g04823(.A0(new_n2919_), .A1(new_n1395_), .B0(new_n5016_), .Y(new_n5017_));
  AOI22X1  g04824(.A0(\a[34] ), .A1(\a[22] ), .B0(\a[33] ), .B1(\a[23] ), .Y(new_n5018_));
  NAND3X1  g04825(.A(new_n5016_), .B(\a[36] ), .C(\a[20] ), .Y(new_n5019_));
  OAI21X1  g04826(.A0(new_n5018_), .A1(new_n5017_), .B0(new_n5019_), .Y(new_n5020_));
  AOI22X1  g04827(.A0(new_n2671_), .A1(new_n1532_), .B0(new_n1787_), .B1(new_n1650_), .Y(new_n5021_));
  AOI21X1  g04828(.A0(new_n2075_), .A1(new_n1770_), .B0(new_n5021_), .Y(new_n5022_));
  NAND2X1  g04829(.A(\a[32] ), .B(\a[24] ), .Y(new_n5023_));
  OAI21X1  g04830(.A0(new_n2076_), .A1(new_n1771_), .B0(new_n5021_), .Y(new_n5024_));
  AOI22X1  g04831(.A0(\a[31] ), .A1(\a[25] ), .B0(\a[30] ), .B1(\a[26] ), .Y(new_n5025_));
  OAI22X1  g04832(.A0(new_n5025_), .A1(new_n5024_), .B0(new_n5023_), .B1(new_n5022_), .Y(new_n5026_));
  XOR2X1   g04833(.A(new_n5026_), .B(new_n5020_), .Y(new_n5027_));
  NOR3X1   g04834(.A(new_n4403_), .B(new_n3460_), .C(new_n490_), .Y(new_n5028_));
  NOR4X1   g04835(.A(new_n4041_), .B(new_n3096_), .C(new_n490_), .D(new_n341_), .Y(new_n5029_));
  AOI21X1  g04836(.A0(new_n3893_), .A1(new_n881_), .B0(new_n5029_), .Y(new_n5030_));
  AND2X1   g04837(.A(\a[47] ), .B(\a[9] ), .Y(new_n5031_));
  OAI21X1  g04838(.A0(new_n5030_), .A1(new_n5028_), .B0(new_n5031_), .Y(new_n5032_));
  NOR2X1   g04839(.A(new_n5030_), .B(new_n5028_), .Y(new_n5033_));
  NOR2X1   g04840(.A(new_n5033_), .B(new_n5028_), .Y(new_n5034_));
  INVX1    g04841(.A(new_n5034_), .Y(new_n5035_));
  AOI22X1  g04842(.A0(\a[46] ), .A1(\a[10] ), .B0(\a[42] ), .B1(\a[14] ), .Y(new_n5036_));
  OAI21X1  g04843(.A0(new_n5036_), .A1(new_n5035_), .B0(new_n5032_), .Y(new_n5037_));
  INVX1    g04844(.A(new_n5037_), .Y(new_n5038_));
  XOR2X1   g04845(.A(new_n5038_), .B(new_n5027_), .Y(new_n5039_));
  XOR2X1   g04846(.A(new_n5039_), .B(new_n5013_), .Y(new_n5040_));
  AND2X1   g04847(.A(new_n4826_), .B(\a[1] ), .Y(new_n5041_));
  AND2X1   g04848(.A(\a[56] ), .B(\a[54] ), .Y(new_n5042_));
  AOI22X1  g04849(.A0(\a[56] ), .A1(\a[0] ), .B0(\a[54] ), .B1(\a[2] ), .Y(new_n5043_));
  AOI21X1  g04850(.A0(new_n5042_), .A1(new_n197_), .B0(new_n5043_), .Y(new_n5044_));
  XOR2X1   g04851(.A(new_n5044_), .B(new_n5041_), .Y(new_n5045_));
  INVX1    g04852(.A(new_n5045_), .Y(new_n5046_));
  XOR2X1   g04853(.A(new_n5046_), .B(new_n4897_), .Y(new_n5047_));
  AND2X1   g04854(.A(\a[53] ), .B(\a[52] ), .Y(new_n5048_));
  AND2X1   g04855(.A(\a[53] ), .B(\a[37] ), .Y(new_n5049_));
  AOI22X1  g04856(.A0(new_n5049_), .A1(new_n942_), .B0(new_n5048_), .B1(new_n294_), .Y(new_n5050_));
  NOR4X1   g04857(.A(new_n4354_), .B(new_n2345_), .C(new_n752_), .D(new_n340_), .Y(new_n5051_));
  OR2X1    g04858(.A(new_n5051_), .B(new_n5050_), .Y(new_n5052_));
  AND2X1   g04859(.A(\a[53] ), .B(\a[3] ), .Y(new_n5053_));
  INVX1    g04860(.A(new_n5051_), .Y(new_n5054_));
  AND2X1   g04861(.A(new_n5054_), .B(new_n5050_), .Y(new_n5055_));
  OAI22X1  g04862(.A0(new_n4354_), .A1(new_n340_), .B0(new_n2345_), .B1(new_n752_), .Y(new_n5056_));
  AOI22X1  g04863(.A0(new_n5056_), .A1(new_n5055_), .B0(new_n5053_), .B1(new_n5052_), .Y(new_n5057_));
  XOR2X1   g04864(.A(new_n5057_), .B(new_n5047_), .Y(new_n5058_));
  INVX1    g04865(.A(new_n5058_), .Y(new_n5059_));
  XOR2X1   g04866(.A(new_n5059_), .B(new_n5040_), .Y(new_n5060_));
  INVX1    g04867(.A(new_n4811_), .Y(new_n5061_));
  OR2X1    g04868(.A(new_n4813_), .B(new_n5061_), .Y(new_n5062_));
  OAI21X1  g04869(.A0(new_n4814_), .A1(new_n4790_), .B0(new_n5062_), .Y(new_n5063_));
  XOR2X1   g04870(.A(new_n4927_), .B(new_n4919_), .Y(new_n5064_));
  XOR2X1   g04871(.A(new_n5064_), .B(new_n4797_), .Y(new_n5065_));
  INVX1    g04872(.A(new_n5065_), .Y(new_n5066_));
  INVX1    g04873(.A(new_n4884_), .Y(new_n5067_));
  AND2X1   g04874(.A(new_n4890_), .B(new_n5067_), .Y(new_n5068_));
  NOR2X1   g04875(.A(new_n4898_), .B(new_n4891_), .Y(new_n5069_));
  NOR2X1   g04876(.A(new_n5069_), .B(new_n5068_), .Y(new_n5070_));
  INVX1    g04877(.A(new_n5070_), .Y(new_n5071_));
  AND2X1   g04878(.A(\a[55] ), .B(\a[1] ), .Y(new_n5072_));
  XOR2X1   g04879(.A(new_n5072_), .B(new_n1484_), .Y(new_n5073_));
  INVX1    g04880(.A(new_n5073_), .Y(new_n5074_));
  NOR3X1   g04881(.A(new_n5074_), .B(new_n4888_), .C(new_n4887_), .Y(new_n5075_));
  XOR2X1   g04882(.A(new_n5074_), .B(new_n4889_), .Y(new_n5076_));
  OAI21X1  g04883(.A0(new_n4888_), .A1(new_n4887_), .B0(new_n5074_), .Y(new_n5077_));
  NAND2X1  g04884(.A(new_n5077_), .B(new_n4880_), .Y(new_n5078_));
  OAI22X1  g04885(.A0(new_n5078_), .A1(new_n5075_), .B0(new_n5076_), .B1(new_n4880_), .Y(new_n5079_));
  XOR2X1   g04886(.A(new_n5079_), .B(new_n5071_), .Y(new_n5080_));
  XOR2X1   g04887(.A(new_n5080_), .B(new_n5066_), .Y(new_n5081_));
  INVX1    g04888(.A(new_n5081_), .Y(new_n5082_));
  XOR2X1   g04889(.A(new_n5082_), .B(new_n5063_), .Y(new_n5083_));
  XOR2X1   g04890(.A(new_n5083_), .B(new_n5060_), .Y(new_n5084_));
  AND2X1   g04891(.A(new_n4690_), .B(new_n4682_), .Y(new_n5085_));
  OAI21X1  g04892(.A0(new_n5085_), .A1(new_n4787_), .B0(new_n4815_), .Y(new_n5086_));
  OAI21X1  g04893(.A0(new_n4816_), .A1(new_n4786_), .B0(new_n5086_), .Y(new_n5087_));
  XOR2X1   g04894(.A(new_n4909_), .B(new_n4846_), .Y(new_n5088_));
  INVX1    g04895(.A(new_n5088_), .Y(new_n5089_));
  XOR2X1   g04896(.A(new_n5089_), .B(new_n4806_), .Y(new_n5090_));
  INVX1    g04897(.A(new_n5090_), .Y(new_n5091_));
  INVX1    g04898(.A(new_n4798_), .Y(new_n5092_));
  OR2X1    g04899(.A(new_n4807_), .B(new_n5092_), .Y(new_n5093_));
  OAI21X1  g04900(.A0(new_n4810_), .A1(new_n4808_), .B0(new_n5093_), .Y(new_n5094_));
  XOR2X1   g04901(.A(new_n5094_), .B(new_n5091_), .Y(new_n5095_));
  NOR2X1   g04902(.A(new_n4823_), .B(new_n4821_), .Y(new_n5096_));
  AOI21X1  g04903(.A0(new_n4830_), .A1(new_n4824_), .B0(new_n5096_), .Y(new_n5097_));
  XOR2X1   g04904(.A(new_n5097_), .B(new_n5095_), .Y(new_n5098_));
  AND2X1   g04905(.A(new_n4655_), .B(new_n4646_), .Y(new_n5099_));
  AOI21X1  g04906(.A0(new_n4866_), .A1(new_n4721_), .B0(new_n5099_), .Y(new_n5100_));
  NOR2X1   g04907(.A(new_n4838_), .B(new_n4742_), .Y(new_n5101_));
  AOI21X1  g04908(.A0(new_n4848_), .A1(new_n4839_), .B0(new_n5101_), .Y(new_n5102_));
  XOR2X1   g04909(.A(new_n5102_), .B(new_n5100_), .Y(new_n5103_));
  OR2X1    g04910(.A(new_n4921_), .B(new_n4913_), .Y(new_n5104_));
  INVX1    g04911(.A(new_n4922_), .Y(new_n5105_));
  OAI21X1  g04912(.A0(new_n4929_), .A1(new_n5105_), .B0(new_n5104_), .Y(new_n5106_));
  XOR2X1   g04913(.A(new_n5106_), .B(new_n5103_), .Y(new_n5107_));
  AND2X1   g04914(.A(new_n4902_), .B(new_n4899_), .Y(new_n5108_));
  NOR2X1   g04915(.A(new_n4930_), .B(new_n4903_), .Y(new_n5109_));
  NOR2X1   g04916(.A(new_n5109_), .B(new_n5108_), .Y(new_n5110_));
  OR2X1    g04917(.A(new_n5110_), .B(new_n5107_), .Y(new_n5111_));
  INVX1    g04918(.A(new_n5110_), .Y(new_n5112_));
  XOR2X1   g04919(.A(new_n5112_), .B(new_n5107_), .Y(new_n5113_));
  AOI21X1  g04920(.A0(new_n5110_), .A1(new_n5107_), .B0(new_n5098_), .Y(new_n5114_));
  AOI22X1  g04921(.A0(new_n5114_), .A1(new_n5111_), .B0(new_n5113_), .B1(new_n5098_), .Y(new_n5115_));
  XOR2X1   g04922(.A(new_n5115_), .B(new_n5087_), .Y(new_n5116_));
  XOR2X1   g04923(.A(new_n5116_), .B(new_n5084_), .Y(new_n5117_));
  NAND3X1  g04924(.A(new_n4975_), .B(new_n4978_), .C(new_n4977_), .Y(new_n5118_));
  AOI21X1  g04925(.A0(new_n4980_), .A1(new_n5118_), .B0(new_n5117_), .Y(new_n5119_));
  AND2X1   g04926(.A(new_n5118_), .B(new_n5117_), .Y(new_n5120_));
  AOI21X1  g04927(.A0(new_n5120_), .A1(new_n4980_), .B0(new_n5119_), .Y(new_n5121_));
  XOR2X1   g04928(.A(new_n5121_), .B(new_n4944_), .Y(new_n5122_));
  INVX1    g04929(.A(new_n4934_), .Y(new_n5123_));
  NOR2X1   g04930(.A(new_n5123_), .B(new_n4782_), .Y(new_n5124_));
  INVX1    g04931(.A(new_n5124_), .Y(new_n5125_));
  AND2X1   g04932(.A(new_n5123_), .B(new_n4782_), .Y(new_n5126_));
  OAI21X1  g04933(.A0(new_n4939_), .A1(new_n5126_), .B0(new_n5125_), .Y(new_n5127_));
  XOR2X1   g04934(.A(new_n5127_), .B(new_n5122_), .Y(\asquared[57] ));
  INVX1    g04935(.A(new_n4975_), .Y(new_n5129_));
  AOI21X1  g04936(.A0(new_n4978_), .A1(new_n4977_), .B0(new_n5129_), .Y(new_n5130_));
  NOR2X1   g04937(.A(new_n5119_), .B(new_n5130_), .Y(new_n5131_));
  INVX1    g04938(.A(new_n5084_), .Y(new_n5132_));
  AND2X1   g04939(.A(new_n5115_), .B(new_n5087_), .Y(new_n5133_));
  AOI21X1  g04940(.A0(new_n5116_), .A1(new_n5132_), .B0(new_n5133_), .Y(new_n5134_));
  INVX1    g04941(.A(new_n5060_), .Y(new_n5135_));
  NAND2X1  g04942(.A(new_n5081_), .B(new_n5063_), .Y(new_n5136_));
  OAI21X1  g04943(.A0(new_n5083_), .A1(new_n5135_), .B0(new_n5136_), .Y(new_n5137_));
  AND2X1   g04944(.A(new_n5112_), .B(new_n5107_), .Y(new_n5138_));
  AND2X1   g04945(.A(new_n5113_), .B(new_n5098_), .Y(new_n5139_));
  OR2X1    g04946(.A(new_n5139_), .B(new_n5138_), .Y(new_n5140_));
  NAND2X1  g04947(.A(new_n5094_), .B(new_n5090_), .Y(new_n5141_));
  OAI21X1  g04948(.A0(new_n5097_), .A1(new_n5095_), .B0(new_n5141_), .Y(new_n5142_));
  OR2X1    g04949(.A(new_n5079_), .B(new_n5070_), .Y(new_n5143_));
  OAI21X1  g04950(.A0(new_n5080_), .A1(new_n5066_), .B0(new_n5143_), .Y(new_n5144_));
  XOR2X1   g04951(.A(new_n5144_), .B(new_n5142_), .Y(new_n5145_));
  NAND4X1  g04952(.A(\a[55] ), .B(\a[29] ), .C(\a[27] ), .D(\a[1] ), .Y(new_n5146_));
  AND2X1   g04953(.A(\a[57] ), .B(\a[0] ), .Y(new_n5147_));
  XOR2X1   g04954(.A(new_n5147_), .B(new_n5146_), .Y(new_n5148_));
  AND2X1   g04955(.A(\a[56] ), .B(\a[1] ), .Y(new_n5149_));
  XOR2X1   g04956(.A(new_n5149_), .B(new_n1803_), .Y(new_n5150_));
  INVX1    g04957(.A(new_n5150_), .Y(new_n5151_));
  XOR2X1   g04958(.A(new_n5151_), .B(new_n5148_), .Y(new_n5152_));
  NOR2X1   g04959(.A(new_n4927_), .B(new_n4919_), .Y(new_n5153_));
  AOI21X1  g04960(.A0(new_n5064_), .A1(new_n4797_), .B0(new_n5153_), .Y(new_n5154_));
  XOR2X1   g04961(.A(new_n5154_), .B(new_n5152_), .Y(new_n5155_));
  OAI22X1  g04962(.A0(new_n4908_), .A1(new_n4905_), .B0(new_n4844_), .B1(new_n4842_), .Y(new_n5156_));
  OAI21X1  g04963(.A0(new_n5089_), .A1(new_n4806_), .B0(new_n5156_), .Y(new_n5157_));
  XOR2X1   g04964(.A(new_n5157_), .B(new_n5155_), .Y(new_n5158_));
  XOR2X1   g04965(.A(new_n5158_), .B(new_n5145_), .Y(new_n5159_));
  XOR2X1   g04966(.A(new_n5159_), .B(new_n5140_), .Y(new_n5160_));
  XOR2X1   g04967(.A(new_n5160_), .B(new_n5137_), .Y(new_n5161_));
  NAND2X1  g04968(.A(new_n5161_), .B(new_n5134_), .Y(new_n5162_));
  OR2X1    g04969(.A(new_n4970_), .B(new_n4968_), .Y(new_n5163_));
  OAI21X1  g04970(.A0(new_n4974_), .A1(new_n4972_), .B0(new_n5163_), .Y(new_n5164_));
  OAI21X1  g04971(.A0(new_n4888_), .A1(new_n4887_), .B0(new_n5073_), .Y(new_n5165_));
  OAI21X1  g04972(.A0(new_n5076_), .A1(new_n4880_), .B0(new_n5165_), .Y(new_n5166_));
  OR2X1    g04973(.A(new_n5046_), .B(new_n4897_), .Y(new_n5167_));
  AND2X1   g04974(.A(new_n5046_), .B(new_n4897_), .Y(new_n5168_));
  OAI21X1  g04975(.A0(new_n5057_), .A1(new_n5168_), .B0(new_n5167_), .Y(new_n5169_));
  XOR2X1   g04976(.A(new_n5169_), .B(new_n5166_), .Y(new_n5170_));
  AND2X1   g04977(.A(new_n5026_), .B(new_n5020_), .Y(new_n5171_));
  AND2X1   g04978(.A(new_n5037_), .B(new_n5027_), .Y(new_n5172_));
  OR2X1    g04979(.A(new_n5172_), .B(new_n5171_), .Y(new_n5173_));
  XOR2X1   g04980(.A(new_n5173_), .B(new_n5170_), .Y(new_n5174_));
  NAND2X1  g04981(.A(new_n5059_), .B(new_n5040_), .Y(new_n5175_));
  OR2X1    g04982(.A(new_n5039_), .B(new_n5013_), .Y(new_n5176_));
  AND2X1   g04983(.A(new_n5176_), .B(new_n5175_), .Y(new_n5177_));
  XOR2X1   g04984(.A(new_n5177_), .B(new_n5174_), .Y(new_n5178_));
  AND2X1   g04985(.A(new_n5000_), .B(new_n4991_), .Y(new_n5179_));
  AOI21X1  g04986(.A0(new_n5011_), .A1(new_n5001_), .B0(new_n5179_), .Y(new_n5180_));
  XOR2X1   g04987(.A(new_n5024_), .B(new_n5009_), .Y(new_n5181_));
  XOR2X1   g04988(.A(new_n5181_), .B(new_n4988_), .Y(new_n5182_));
  INVX1    g04989(.A(new_n5055_), .Y(new_n5183_));
  XOR2X1   g04990(.A(new_n5183_), .B(new_n5017_), .Y(new_n5184_));
  AOI22X1  g04991(.A0(new_n5044_), .A1(new_n5041_), .B0(new_n5042_), .B1(new_n197_), .Y(new_n5185_));
  INVX1    g04992(.A(new_n5185_), .Y(new_n5186_));
  XOR2X1   g04993(.A(new_n5186_), .B(new_n5184_), .Y(new_n5187_));
  INVX1    g04994(.A(new_n5187_), .Y(new_n5188_));
  XOR2X1   g04995(.A(new_n5188_), .B(new_n5182_), .Y(new_n5189_));
  INVX1    g04996(.A(new_n5189_), .Y(new_n5190_));
  XOR2X1   g04997(.A(new_n5190_), .B(new_n5180_), .Y(new_n5191_));
  INVX1    g04998(.A(new_n5191_), .Y(new_n5192_));
  XOR2X1   g04999(.A(new_n5192_), .B(new_n5178_), .Y(new_n5193_));
  XOR2X1   g05000(.A(new_n5193_), .B(new_n5164_), .Y(new_n5194_));
  OR2X1    g05001(.A(new_n4964_), .B(new_n4962_), .Y(new_n5195_));
  OAI21X1  g05002(.A0(new_n4966_), .A1(new_n4946_), .B0(new_n5195_), .Y(new_n5196_));
  XOR2X1   g05003(.A(new_n4954_), .B(new_n5034_), .Y(new_n5197_));
  XOR2X1   g05004(.A(new_n5197_), .B(new_n4999_), .Y(new_n5198_));
  INVX1    g05005(.A(new_n5198_), .Y(new_n5199_));
  NAND2X1  g05006(.A(new_n4956_), .B(new_n4948_), .Y(new_n5200_));
  OAI21X1  g05007(.A0(new_n4960_), .A1(new_n4958_), .B0(new_n5200_), .Y(new_n5201_));
  XOR2X1   g05008(.A(new_n5201_), .B(new_n5199_), .Y(new_n5202_));
  NAND2X1  g05009(.A(\a[49] ), .B(\a[16] ), .Y(new_n5203_));
  NOR3X1   g05010(.A(new_n5203_), .B(new_n3081_), .C(new_n413_), .Y(new_n5204_));
  NAND4X1  g05011(.A(\a[50] ), .B(\a[49] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n5205_));
  NAND4X1  g05012(.A(\a[50] ), .B(\a[41] ), .C(\a[16] ), .D(\a[7] ), .Y(new_n5206_));
  AOI21X1  g05013(.A0(new_n5206_), .A1(new_n5205_), .B0(new_n5204_), .Y(new_n5207_));
  OR2X1    g05014(.A(new_n5207_), .B(new_n5204_), .Y(new_n5208_));
  AOI22X1  g05015(.A0(\a[49] ), .A1(\a[8] ), .B0(\a[41] ), .B1(\a[16] ), .Y(new_n5209_));
  NAND2X1  g05016(.A(\a[50] ), .B(\a[7] ), .Y(new_n5210_));
  OAI22X1  g05017(.A0(new_n5210_), .A1(new_n5207_), .B0(new_n5209_), .B1(new_n5208_), .Y(new_n5211_));
  NAND4X1  g05018(.A(\a[36] ), .B(\a[34] ), .C(\a[23] ), .D(\a[21] ), .Y(new_n5212_));
  NAND4X1  g05019(.A(\a[36] ), .B(\a[35] ), .C(\a[22] ), .D(\a[21] ), .Y(new_n5213_));
  AOI22X1  g05020(.A0(new_n5213_), .A1(new_n5212_), .B0(new_n2361_), .B1(new_n1394_), .Y(new_n5214_));
  NAND2X1  g05021(.A(\a[36] ), .B(\a[21] ), .Y(new_n5215_));
  AOI22X1  g05022(.A0(\a[35] ), .A1(\a[22] ), .B0(\a[34] ), .B1(\a[23] ), .Y(new_n5216_));
  AOI21X1  g05023(.A0(new_n2361_), .A1(new_n1394_), .B0(new_n5214_), .Y(new_n5217_));
  INVX1    g05024(.A(new_n5217_), .Y(new_n5218_));
  OAI22X1  g05025(.A0(new_n5218_), .A1(new_n5216_), .B0(new_n5215_), .B1(new_n5214_), .Y(new_n5219_));
  XOR2X1   g05026(.A(new_n5219_), .B(new_n5211_), .Y(new_n5220_));
  NAND4X1  g05027(.A(\a[32] ), .B(\a[31] ), .C(\a[26] ), .D(\a[25] ), .Y(new_n5221_));
  OAI22X1  g05028(.A0(new_n2675_), .A1(new_n1772_), .B0(new_n2673_), .B1(new_n1651_), .Y(new_n5222_));
  AND2X1   g05029(.A(new_n5222_), .B(new_n5221_), .Y(new_n5223_));
  AND2X1   g05030(.A(\a[33] ), .B(\a[24] ), .Y(new_n5224_));
  INVX1    g05031(.A(new_n5224_), .Y(new_n5225_));
  AOI21X1  g05032(.A0(new_n2671_), .A1(new_n1770_), .B0(new_n5222_), .Y(new_n5226_));
  INVX1    g05033(.A(new_n5226_), .Y(new_n5227_));
  AOI22X1  g05034(.A0(\a[32] ), .A1(\a[25] ), .B0(\a[31] ), .B1(\a[26] ), .Y(new_n5228_));
  OAI22X1  g05035(.A0(new_n5228_), .A1(new_n5227_), .B0(new_n5225_), .B1(new_n5223_), .Y(new_n5229_));
  INVX1    g05036(.A(new_n5229_), .Y(new_n5230_));
  XOR2X1   g05037(.A(new_n5230_), .B(new_n5220_), .Y(new_n5231_));
  XOR2X1   g05038(.A(new_n5231_), .B(new_n5202_), .Y(new_n5232_));
  XOR2X1   g05039(.A(new_n5232_), .B(new_n5196_), .Y(new_n5233_));
  NOR2X1   g05040(.A(new_n5102_), .B(new_n5100_), .Y(new_n5234_));
  AOI21X1  g05041(.A0(new_n5106_), .A1(new_n5103_), .B0(new_n5234_), .Y(new_n5235_));
  AND2X1   g05042(.A(\a[55] ), .B(\a[53] ), .Y(new_n5236_));
  INVX1    g05043(.A(new_n5236_), .Y(new_n5237_));
  AND2X1   g05044(.A(\a[54] ), .B(\a[53] ), .Y(new_n5238_));
  INVX1    g05045(.A(new_n5238_), .Y(new_n5239_));
  AND2X1   g05046(.A(\a[55] ), .B(\a[54] ), .Y(new_n5240_));
  INVX1    g05047(.A(new_n5240_), .Y(new_n5241_));
  OAI22X1  g05048(.A0(new_n5241_), .A1(new_n249_), .B0(new_n5239_), .B1(new_n217_), .Y(new_n5242_));
  OAI21X1  g05049(.A0(new_n5237_), .A1(new_n584_), .B0(new_n5242_), .Y(new_n5243_));
  AOI21X1  g05050(.A0(new_n5236_), .A1(new_n235_), .B0(new_n5242_), .Y(new_n5244_));
  INVX1    g05051(.A(\a[53] ), .Y(new_n5245_));
  OAI22X1  g05052(.A0(new_n4906_), .A1(new_n200_), .B0(new_n5245_), .B1(new_n340_), .Y(new_n5246_));
  AND2X1   g05053(.A(\a[54] ), .B(\a[3] ), .Y(new_n5247_));
  AOI22X1  g05054(.A0(new_n5247_), .A1(new_n5243_), .B0(new_n5246_), .B1(new_n5244_), .Y(new_n5248_));
  AND2X1   g05055(.A(\a[52] ), .B(\a[5] ), .Y(new_n5249_));
  INVX1    g05056(.A(new_n5249_), .Y(new_n5250_));
  AOI22X1  g05057(.A0(\a[38] ), .A1(\a[19] ), .B0(\a[37] ), .B1(\a[20] ), .Y(new_n5251_));
  AND2X1   g05058(.A(new_n3164_), .B(new_n1099_), .Y(new_n5252_));
  NOR3X1   g05059(.A(new_n5251_), .B(new_n5252_), .C(new_n5250_), .Y(new_n5253_));
  INVX1    g05060(.A(new_n5251_), .Y(new_n5254_));
  AOI21X1  g05061(.A0(new_n5254_), .A1(new_n5249_), .B0(new_n5252_), .Y(new_n5255_));
  INVX1    g05062(.A(new_n5255_), .Y(new_n5256_));
  OAI22X1  g05063(.A0(new_n5256_), .A1(new_n5251_), .B0(new_n5253_), .B1(new_n5250_), .Y(new_n5257_));
  XOR2X1   g05064(.A(new_n5257_), .B(new_n5248_), .Y(new_n5258_));
  AND2X1   g05065(.A(\a[42] ), .B(\a[15] ), .Y(new_n5259_));
  AOI22X1  g05066(.A0(\a[48] ), .A1(\a[9] ), .B0(\a[47] ), .B1(\a[10] ), .Y(new_n5260_));
  INVX1    g05067(.A(new_n5260_), .Y(new_n5261_));
  NAND4X1  g05068(.A(\a[48] ), .B(\a[47] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n5262_));
  NAND3X1  g05069(.A(new_n5261_), .B(new_n5262_), .C(new_n5259_), .Y(new_n5263_));
  AOI22X1  g05070(.A0(new_n5261_), .A1(new_n5259_), .B0(new_n4272_), .B1(new_n881_), .Y(new_n5264_));
  AOI22X1  g05071(.A0(new_n5264_), .A1(new_n5261_), .B0(new_n5263_), .B1(new_n5259_), .Y(new_n5265_));
  XOR2X1   g05072(.A(new_n5265_), .B(new_n5258_), .Y(new_n5266_));
  INVX1    g05073(.A(new_n5266_), .Y(new_n5267_));
  INVX1    g05074(.A(\a[44] ), .Y(new_n5268_));
  OAI22X1  g05075(.A0(new_n3460_), .A1(new_n488_), .B0(new_n5268_), .B1(new_n591_), .Y(new_n5269_));
  AND2X1   g05076(.A(\a[46] ), .B(\a[44] ), .Y(new_n5270_));
  NAND4X1  g05077(.A(\a[44] ), .B(\a[43] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n5271_));
  NAND4X1  g05078(.A(\a[46] ), .B(\a[43] ), .C(\a[14] ), .D(\a[11] ), .Y(new_n5272_));
  AOI22X1  g05079(.A0(new_n5272_), .A1(new_n5271_), .B0(new_n5270_), .B1(new_n634_), .Y(new_n5273_));
  AOI21X1  g05080(.A0(new_n5270_), .A1(new_n634_), .B0(new_n5273_), .Y(new_n5274_));
  NOR3X1   g05081(.A(new_n5273_), .B(new_n3037_), .C(new_n490_), .Y(new_n5275_));
  AOI21X1  g05082(.A0(new_n5274_), .A1(new_n5269_), .B0(new_n5275_), .Y(new_n5276_));
  AND2X1   g05083(.A(\a[45] ), .B(\a[12] ), .Y(new_n5277_));
  INVX1    g05084(.A(new_n5277_), .Y(new_n5278_));
  AOI22X1  g05085(.A0(\a[30] ), .A1(\a[27] ), .B0(\a[29] ), .B1(\a[28] ), .Y(new_n5279_));
  AND2X1   g05086(.A(new_n2196_), .B(new_n1671_), .Y(new_n5280_));
  NOR3X1   g05087(.A(new_n5279_), .B(new_n5280_), .C(new_n5278_), .Y(new_n5281_));
  INVX1    g05088(.A(new_n5279_), .Y(new_n5282_));
  AOI21X1  g05089(.A0(new_n5282_), .A1(new_n5277_), .B0(new_n5280_), .Y(new_n5283_));
  INVX1    g05090(.A(new_n5283_), .Y(new_n5284_));
  OAI22X1  g05091(.A0(new_n5284_), .A1(new_n5279_), .B0(new_n5281_), .B1(new_n5278_), .Y(new_n5285_));
  XOR2X1   g05092(.A(new_n5285_), .B(new_n5276_), .Y(new_n5286_));
  INVX1    g05093(.A(new_n5286_), .Y(new_n5287_));
  NOR4X1   g05094(.A(new_n4349_), .B(new_n3036_), .C(new_n616_), .D(new_n230_), .Y(new_n5288_));
  AND2X1   g05095(.A(\a[18] ), .B(\a[6] ), .Y(new_n5289_));
  AND2X1   g05096(.A(\a[51] ), .B(\a[39] ), .Y(new_n5290_));
  AOI22X1  g05097(.A0(new_n5290_), .A1(new_n5289_), .B0(new_n4077_), .B1(new_n796_), .Y(new_n5291_));
  OR2X1    g05098(.A(new_n5291_), .B(new_n5288_), .Y(new_n5292_));
  AND2X1   g05099(.A(\a[39] ), .B(\a[18] ), .Y(new_n5293_));
  INVX1    g05100(.A(new_n5288_), .Y(new_n5294_));
  AND2X1   g05101(.A(new_n5291_), .B(new_n5294_), .Y(new_n5295_));
  OAI22X1  g05102(.A0(new_n4349_), .A1(new_n230_), .B0(new_n3036_), .B1(new_n616_), .Y(new_n5296_));
  AOI22X1  g05103(.A0(new_n5296_), .A1(new_n5295_), .B0(new_n5293_), .B1(new_n5292_), .Y(new_n5297_));
  XOR2X1   g05104(.A(new_n5297_), .B(new_n5287_), .Y(new_n5298_));
  XOR2X1   g05105(.A(new_n5298_), .B(new_n5267_), .Y(new_n5299_));
  INVX1    g05106(.A(new_n5299_), .Y(new_n5300_));
  XOR2X1   g05107(.A(new_n5300_), .B(new_n5235_), .Y(new_n5301_));
  INVX1    g05108(.A(new_n5301_), .Y(new_n5302_));
  XOR2X1   g05109(.A(new_n5302_), .B(new_n5233_), .Y(new_n5303_));
  XOR2X1   g05110(.A(new_n5303_), .B(new_n5194_), .Y(new_n5304_));
  OR2X1    g05111(.A(new_n5161_), .B(new_n5134_), .Y(new_n5305_));
  AOI21X1  g05112(.A0(new_n5162_), .A1(new_n5305_), .B0(new_n5304_), .Y(new_n5306_));
  AND2X1   g05113(.A(new_n5305_), .B(new_n5304_), .Y(new_n5307_));
  AOI21X1  g05114(.A0(new_n5307_), .A1(new_n5162_), .B0(new_n5306_), .Y(new_n5308_));
  XOR2X1   g05115(.A(new_n5308_), .B(new_n5131_), .Y(new_n5309_));
  AND2X1   g05116(.A(new_n5121_), .B(new_n4944_), .Y(new_n5310_));
  NOR2X1   g05117(.A(new_n5121_), .B(new_n4944_), .Y(new_n5311_));
  INVX1    g05118(.A(new_n5311_), .Y(new_n5312_));
  AOI21X1  g05119(.A0(new_n5127_), .A1(new_n5312_), .B0(new_n5310_), .Y(new_n5313_));
  XOR2X1   g05120(.A(new_n5313_), .B(new_n5309_), .Y(\asquared[58] ));
  INVX1    g05121(.A(new_n5134_), .Y(new_n5315_));
  AOI21X1  g05122(.A0(new_n5161_), .A1(new_n5315_), .B0(new_n5306_), .Y(new_n5316_));
  AND2X1   g05123(.A(new_n5193_), .B(new_n5164_), .Y(new_n5317_));
  INVX1    g05124(.A(new_n5317_), .Y(new_n5318_));
  INVX1    g05125(.A(new_n5194_), .Y(new_n5319_));
  OAI21X1  g05126(.A0(new_n5303_), .A1(new_n5319_), .B0(new_n5318_), .Y(new_n5320_));
  INVX1    g05127(.A(new_n5177_), .Y(new_n5321_));
  NOR2X1   g05128(.A(new_n5192_), .B(new_n5178_), .Y(new_n5322_));
  AOI21X1  g05129(.A0(new_n5321_), .A1(new_n5174_), .B0(new_n5322_), .Y(new_n5323_));
  NAND2X1  g05130(.A(new_n5201_), .B(new_n5198_), .Y(new_n5324_));
  OAI21X1  g05131(.A0(new_n5231_), .A1(new_n5202_), .B0(new_n5324_), .Y(new_n5325_));
  NOR2X1   g05132(.A(new_n4954_), .B(new_n5034_), .Y(new_n5326_));
  AOI21X1  g05133(.A0(new_n5197_), .A1(new_n4999_), .B0(new_n5326_), .Y(new_n5327_));
  AND2X1   g05134(.A(new_n5183_), .B(new_n5017_), .Y(new_n5328_));
  AOI21X1  g05135(.A0(new_n5186_), .A1(new_n5184_), .B0(new_n5328_), .Y(new_n5329_));
  XOR2X1   g05136(.A(new_n5329_), .B(new_n5327_), .Y(new_n5330_));
  INVX1    g05137(.A(new_n5330_), .Y(new_n5331_));
  AND2X1   g05138(.A(new_n5024_), .B(new_n5009_), .Y(new_n5332_));
  AOI21X1  g05139(.A0(new_n5181_), .A1(new_n4989_), .B0(new_n5332_), .Y(new_n5333_));
  XOR2X1   g05140(.A(new_n5333_), .B(new_n5331_), .Y(new_n5334_));
  OR2X1    g05141(.A(new_n5188_), .B(new_n5182_), .Y(new_n5335_));
  OAI21X1  g05142(.A0(new_n5190_), .A1(new_n5180_), .B0(new_n5335_), .Y(new_n5336_));
  XOR2X1   g05143(.A(new_n5336_), .B(new_n5334_), .Y(new_n5337_));
  XOR2X1   g05144(.A(new_n5337_), .B(new_n5325_), .Y(new_n5338_));
  XOR2X1   g05145(.A(new_n5338_), .B(new_n5323_), .Y(new_n5339_));
  AND2X1   g05146(.A(new_n5232_), .B(new_n5196_), .Y(new_n5340_));
  AOI21X1  g05147(.A0(new_n5301_), .A1(new_n5233_), .B0(new_n5340_), .Y(new_n5341_));
  XOR2X1   g05148(.A(new_n5341_), .B(new_n5339_), .Y(new_n5342_));
  XOR2X1   g05149(.A(new_n5342_), .B(new_n5320_), .Y(new_n5343_));
  AND2X1   g05150(.A(new_n5159_), .B(new_n5140_), .Y(new_n5344_));
  AOI21X1  g05151(.A0(new_n5160_), .A1(new_n5137_), .B0(new_n5344_), .Y(new_n5345_));
  OR2X1    g05152(.A(new_n5298_), .B(new_n5267_), .Y(new_n5346_));
  OAI21X1  g05153(.A0(new_n5300_), .A1(new_n5235_), .B0(new_n5346_), .Y(new_n5347_));
  AND2X1   g05154(.A(new_n5274_), .B(new_n5269_), .Y(new_n5348_));
  OAI21X1  g05155(.A0(new_n5275_), .A1(new_n5348_), .B0(new_n5285_), .Y(new_n5349_));
  OAI21X1  g05156(.A0(new_n5297_), .A1(new_n5286_), .B0(new_n5349_), .Y(new_n5350_));
  INVX1    g05157(.A(new_n5257_), .Y(new_n5351_));
  OR2X1    g05158(.A(new_n5351_), .B(new_n5248_), .Y(new_n5352_));
  OAI21X1  g05159(.A0(new_n5265_), .A1(new_n5258_), .B0(new_n5352_), .Y(new_n5353_));
  AND2X1   g05160(.A(new_n5149_), .B(\a[29] ), .Y(new_n5354_));
  AND2X1   g05161(.A(\a[57] ), .B(\a[1] ), .Y(new_n5355_));
  XOR2X1   g05162(.A(new_n5355_), .B(new_n2198_), .Y(new_n5356_));
  XOR2X1   g05163(.A(new_n5356_), .B(new_n5354_), .Y(new_n5357_));
  XOR2X1   g05164(.A(new_n5357_), .B(new_n5284_), .Y(new_n5358_));
  INVX1    g05165(.A(new_n5358_), .Y(new_n5359_));
  OR2X1    g05166(.A(new_n5359_), .B(new_n5353_), .Y(new_n5360_));
  XOR2X1   g05167(.A(new_n5358_), .B(new_n5353_), .Y(new_n5361_));
  AOI21X1  g05168(.A0(new_n5359_), .A1(new_n5353_), .B0(new_n5350_), .Y(new_n5362_));
  AOI22X1  g05169(.A0(new_n5362_), .A1(new_n5360_), .B0(new_n5361_), .B1(new_n5350_), .Y(new_n5363_));
  XOR2X1   g05170(.A(new_n5363_), .B(new_n5347_), .Y(new_n5364_));
  AND2X1   g05171(.A(new_n5219_), .B(new_n5211_), .Y(new_n5365_));
  AOI21X1  g05172(.A0(new_n5229_), .A1(new_n5220_), .B0(new_n5365_), .Y(new_n5366_));
  XOR2X1   g05173(.A(new_n5264_), .B(new_n5226_), .Y(new_n5367_));
  XOR2X1   g05174(.A(new_n5367_), .B(new_n5217_), .Y(new_n5368_));
  INVX1    g05175(.A(new_n5274_), .Y(new_n5369_));
  XOR2X1   g05176(.A(new_n5255_), .B(new_n5244_), .Y(new_n5370_));
  XOR2X1   g05177(.A(new_n5370_), .B(new_n5369_), .Y(new_n5371_));
  INVX1    g05178(.A(new_n5371_), .Y(new_n5372_));
  XOR2X1   g05179(.A(new_n5372_), .B(new_n5368_), .Y(new_n5373_));
  INVX1    g05180(.A(new_n5373_), .Y(new_n5374_));
  XOR2X1   g05181(.A(new_n5374_), .B(new_n5366_), .Y(new_n5375_));
  INVX1    g05182(.A(new_n5375_), .Y(new_n5376_));
  XOR2X1   g05183(.A(new_n5376_), .B(new_n5364_), .Y(new_n5377_));
  XOR2X1   g05184(.A(new_n5377_), .B(new_n5345_), .Y(new_n5378_));
  INVX1    g05185(.A(\a[58] ), .Y(new_n5379_));
  NOR4X1   g05186(.A(new_n5379_), .B(new_n4835_), .C(new_n340_), .D(new_n194_), .Y(new_n5380_));
  AND2X1   g05187(.A(\a[58] ), .B(\a[56] ), .Y(new_n5381_));
  AOI22X1  g05188(.A0(new_n5381_), .A1(new_n197_), .B0(new_n5042_), .B1(new_n235_), .Y(new_n5382_));
  OR2X1    g05189(.A(new_n5382_), .B(new_n5380_), .Y(new_n5383_));
  INVX1    g05190(.A(new_n5380_), .Y(new_n5384_));
  AND2X1   g05191(.A(new_n5382_), .B(new_n5384_), .Y(new_n5385_));
  OAI22X1  g05192(.A0(new_n5379_), .A1(new_n194_), .B0(new_n4835_), .B1(new_n340_), .Y(new_n5386_));
  AND2X1   g05193(.A(\a[56] ), .B(\a[2] ), .Y(new_n5387_));
  AOI22X1  g05194(.A0(new_n5387_), .A1(new_n5383_), .B0(new_n5386_), .B1(new_n5385_), .Y(new_n5388_));
  AND2X1   g05195(.A(\a[53] ), .B(\a[5] ), .Y(new_n5389_));
  INVX1    g05196(.A(new_n5389_), .Y(new_n5390_));
  AOI22X1  g05197(.A0(\a[38] ), .A1(\a[20] ), .B0(\a[37] ), .B1(\a[21] ), .Y(new_n5391_));
  AND2X1   g05198(.A(new_n3164_), .B(new_n1236_), .Y(new_n5392_));
  NOR3X1   g05199(.A(new_n5391_), .B(new_n5392_), .C(new_n5390_), .Y(new_n5393_));
  INVX1    g05200(.A(new_n5391_), .Y(new_n5394_));
  AOI21X1  g05201(.A0(new_n5394_), .A1(new_n5389_), .B0(new_n5392_), .Y(new_n5395_));
  INVX1    g05202(.A(new_n5395_), .Y(new_n5396_));
  OAI22X1  g05203(.A0(new_n5396_), .A1(new_n5391_), .B0(new_n5393_), .B1(new_n5390_), .Y(new_n5397_));
  XOR2X1   g05204(.A(new_n5397_), .B(new_n5388_), .Y(new_n5398_));
  AND2X1   g05205(.A(\a[49] ), .B(\a[42] ), .Y(new_n5399_));
  NAND4X1  g05206(.A(\a[42] ), .B(\a[41] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n5400_));
  NAND4X1  g05207(.A(\a[49] ), .B(\a[41] ), .C(\a[17] ), .D(\a[9] ), .Y(new_n5401_));
  AOI22X1  g05208(.A0(new_n5401_), .A1(new_n5400_), .B0(new_n5399_), .B1(new_n657_), .Y(new_n5402_));
  NOR3X1   g05209(.A(new_n5402_), .B(new_n3081_), .C(new_n616_), .Y(new_n5403_));
  OAI22X1  g05210(.A0(new_n3915_), .A1(new_n341_), .B0(new_n3096_), .B1(new_n571_), .Y(new_n5404_));
  AND2X1   g05211(.A(new_n5399_), .B(new_n657_), .Y(new_n5405_));
  NOR2X1   g05212(.A(new_n5402_), .B(new_n5405_), .Y(new_n5406_));
  AOI21X1  g05213(.A0(new_n5406_), .A1(new_n5404_), .B0(new_n5403_), .Y(new_n5407_));
  XOR2X1   g05214(.A(new_n5407_), .B(new_n5398_), .Y(new_n5408_));
  AOI22X1  g05215(.A0(\a[51] ), .A1(\a[7] ), .B0(\a[50] ), .B1(\a[8] ), .Y(new_n5409_));
  AND2X1   g05216(.A(\a[40] ), .B(\a[18] ), .Y(new_n5410_));
  INVX1    g05217(.A(new_n5410_), .Y(new_n5411_));
  AND2X1   g05218(.A(new_n4484_), .B(new_n325_), .Y(new_n5412_));
  NOR3X1   g05219(.A(new_n5411_), .B(new_n5412_), .C(new_n5409_), .Y(new_n5413_));
  NOR2X1   g05220(.A(new_n5413_), .B(new_n5412_), .Y(new_n5414_));
  INVX1    g05221(.A(new_n5414_), .Y(new_n5415_));
  OAI22X1  g05222(.A0(new_n5415_), .A1(new_n5409_), .B0(new_n5413_), .B1(new_n5411_), .Y(new_n5416_));
  INVX1    g05223(.A(new_n2682_), .Y(new_n5417_));
  INVX1    g05224(.A(new_n4695_), .Y(new_n5418_));
  OAI22X1  g05225(.A0(new_n5418_), .A1(new_n1531_), .B0(new_n5417_), .B1(new_n1395_), .Y(new_n5419_));
  OAI21X1  g05226(.A0(new_n4915_), .A1(new_n1652_), .B0(new_n5419_), .Y(new_n5420_));
  AND2X1   g05227(.A(\a[36] ), .B(\a[22] ), .Y(new_n5421_));
  AOI21X1  g05228(.A0(new_n2361_), .A1(new_n1219_), .B0(new_n5419_), .Y(new_n5422_));
  OAI22X1  g05229(.A0(new_n2557_), .A1(new_n1216_), .B0(new_n2028_), .B1(new_n1185_), .Y(new_n5423_));
  AOI22X1  g05230(.A0(new_n5423_), .A1(new_n5422_), .B0(new_n5421_), .B1(new_n5420_), .Y(new_n5424_));
  XOR2X1   g05231(.A(new_n5424_), .B(new_n5416_), .Y(new_n5425_));
  INVX1    g05232(.A(new_n5425_), .Y(new_n5426_));
  OAI22X1  g05233(.A0(new_n2675_), .A1(new_n1771_), .B0(new_n3484_), .B1(new_n2673_), .Y(new_n5427_));
  OAI21X1  g05234(.A0(new_n2672_), .A1(new_n3483_), .B0(new_n5427_), .Y(new_n5428_));
  AOI21X1  g05235(.A0(new_n2671_), .A1(new_n1995_), .B0(new_n5427_), .Y(new_n5429_));
  OAI22X1  g05236(.A0(new_n2219_), .A1(new_n1263_), .B0(new_n1704_), .B1(new_n1679_), .Y(new_n5430_));
  AOI22X1  g05237(.A0(new_n5430_), .A1(new_n5429_), .B0(new_n5428_), .B1(new_n2346_), .Y(new_n5431_));
  XOR2X1   g05238(.A(new_n5431_), .B(new_n5426_), .Y(new_n5432_));
  XOR2X1   g05239(.A(new_n5432_), .B(new_n5408_), .Y(new_n5433_));
  AND2X1   g05240(.A(new_n5169_), .B(new_n5166_), .Y(new_n5434_));
  AOI21X1  g05241(.A0(new_n5173_), .A1(new_n5170_), .B0(new_n5434_), .Y(new_n5435_));
  XOR2X1   g05242(.A(new_n5435_), .B(new_n5433_), .Y(new_n5436_));
  AND2X1   g05243(.A(new_n5144_), .B(new_n5142_), .Y(new_n5437_));
  AOI21X1  g05244(.A0(new_n5158_), .A1(new_n5145_), .B0(new_n5437_), .Y(new_n5438_));
  INVX1    g05245(.A(new_n5295_), .Y(new_n5439_));
  XOR2X1   g05246(.A(new_n5439_), .B(new_n5208_), .Y(new_n5440_));
  INVX1    g05247(.A(\a[57] ), .Y(new_n5441_));
  NOR3X1   g05248(.A(new_n5146_), .B(new_n5441_), .C(new_n194_), .Y(new_n5442_));
  NOR2X1   g05249(.A(new_n5150_), .B(new_n5148_), .Y(new_n5443_));
  NOR2X1   g05250(.A(new_n5443_), .B(new_n5442_), .Y(new_n5444_));
  XOR2X1   g05251(.A(new_n5444_), .B(new_n5440_), .Y(new_n5445_));
  NOR2X1   g05252(.A(new_n5154_), .B(new_n5152_), .Y(new_n5446_));
  AOI21X1  g05253(.A0(new_n5157_), .A1(new_n5155_), .B0(new_n5446_), .Y(new_n5447_));
  XOR2X1   g05254(.A(new_n5447_), .B(new_n5445_), .Y(new_n5448_));
  NOR3X1   g05255(.A(new_n633_), .B(new_n4041_), .C(new_n3037_), .Y(new_n5449_));
  NAND4X1  g05256(.A(\a[48] ), .B(\a[47] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n5450_));
  NAND4X1  g05257(.A(\a[48] ), .B(\a[43] ), .C(\a[15] ), .D(\a[10] ), .Y(new_n5451_));
  AOI21X1  g05258(.A0(new_n5451_), .A1(new_n5450_), .B0(new_n5449_), .Y(new_n5452_));
  OR2X1    g05259(.A(new_n5452_), .B(new_n5449_), .Y(new_n5453_));
  AOI22X1  g05260(.A0(\a[47] ), .A1(\a[11] ), .B0(\a[43] ), .B1(\a[15] ), .Y(new_n5454_));
  NAND2X1  g05261(.A(\a[48] ), .B(\a[10] ), .Y(new_n5455_));
  OAI22X1  g05262(.A0(new_n5455_), .A1(new_n5452_), .B0(new_n5454_), .B1(new_n5453_), .Y(new_n5456_));
  NAND4X1  g05263(.A(\a[46] ), .B(\a[44] ), .C(\a[14] ), .D(\a[12] ), .Y(new_n5457_));
  NAND4X1  g05264(.A(\a[45] ), .B(\a[44] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n5458_));
  AOI22X1  g05265(.A0(new_n5458_), .A1(new_n5457_), .B0(new_n3809_), .B1(new_n586_), .Y(new_n5459_));
  NAND4X1  g05266(.A(\a[46] ), .B(\a[45] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n5460_));
  NAND3X1  g05267(.A(new_n5458_), .B(new_n5457_), .C(new_n5460_), .Y(new_n5461_));
  AOI22X1  g05268(.A0(\a[46] ), .A1(\a[12] ), .B0(\a[45] ), .B1(\a[13] ), .Y(new_n5462_));
  OAI22X1  g05269(.A0(new_n5462_), .A1(new_n5461_), .B0(new_n5459_), .B1(new_n4518_), .Y(new_n5463_));
  XOR2X1   g05270(.A(new_n5463_), .B(new_n5456_), .Y(new_n5464_));
  AOI22X1  g05271(.A0(\a[52] ), .A1(\a[6] ), .B0(\a[39] ), .B1(\a[19] ), .Y(new_n5465_));
  AND2X1   g05272(.A(\a[55] ), .B(\a[3] ), .Y(new_n5466_));
  NOR4X1   g05273(.A(new_n4354_), .B(new_n2652_), .C(new_n752_), .D(new_n230_), .Y(new_n5467_));
  OAI21X1  g05274(.A0(new_n5465_), .A1(new_n5467_), .B0(new_n5466_), .Y(new_n5468_));
  INVX1    g05275(.A(new_n5465_), .Y(new_n5469_));
  AOI21X1  g05276(.A0(new_n5469_), .A1(new_n5466_), .B0(new_n5467_), .Y(new_n5470_));
  INVX1    g05277(.A(new_n5470_), .Y(new_n5471_));
  OAI21X1  g05278(.A0(new_n5471_), .A1(new_n5465_), .B0(new_n5468_), .Y(new_n5472_));
  XOR2X1   g05279(.A(new_n5472_), .B(new_n5464_), .Y(new_n5473_));
  XOR2X1   g05280(.A(new_n5473_), .B(new_n5448_), .Y(new_n5474_));
  XOR2X1   g05281(.A(new_n5474_), .B(new_n5438_), .Y(new_n5475_));
  XOR2X1   g05282(.A(new_n5475_), .B(new_n5436_), .Y(new_n5476_));
  XOR2X1   g05283(.A(new_n5476_), .B(new_n5378_), .Y(new_n5477_));
  XOR2X1   g05284(.A(new_n5477_), .B(new_n5343_), .Y(new_n5478_));
  NOR2X1   g05285(.A(new_n5478_), .B(new_n5316_), .Y(new_n5479_));
  INVX1    g05286(.A(new_n5479_), .Y(new_n5480_));
  OAI21X1  g05287(.A0(new_n5119_), .A1(new_n5130_), .B0(new_n5308_), .Y(new_n5481_));
  NOR3X1   g05288(.A(new_n5308_), .B(new_n5119_), .C(new_n5130_), .Y(new_n5482_));
  OAI21X1  g05289(.A0(new_n5313_), .A1(new_n5482_), .B0(new_n5481_), .Y(new_n5483_));
  AND2X1   g05290(.A(new_n5478_), .B(new_n5316_), .Y(new_n5484_));
  INVX1    g05291(.A(new_n5484_), .Y(new_n5485_));
  AOI21X1  g05292(.A0(new_n5485_), .A1(new_n5480_), .B0(new_n5483_), .Y(new_n5486_));
  AND2X1   g05293(.A(new_n5485_), .B(new_n5483_), .Y(new_n5487_));
  AOI21X1  g05294(.A0(new_n5487_), .A1(new_n5480_), .B0(new_n5486_), .Y(\asquared[59] ));
  NOR2X1   g05295(.A(new_n5377_), .B(new_n5345_), .Y(new_n5489_));
  INVX1    g05296(.A(new_n5489_), .Y(new_n5490_));
  INVX1    g05297(.A(new_n5378_), .Y(new_n5491_));
  OAI21X1  g05298(.A0(new_n5476_), .A1(new_n5491_), .B0(new_n5490_), .Y(new_n5492_));
  INVX1    g05299(.A(new_n5436_), .Y(new_n5493_));
  INVX1    g05300(.A(new_n5474_), .Y(new_n5494_));
  OR2X1    g05301(.A(new_n5494_), .B(new_n5438_), .Y(new_n5495_));
  OAI21X1  g05302(.A0(new_n5475_), .A1(new_n5493_), .B0(new_n5495_), .Y(new_n5496_));
  NAND2X1  g05303(.A(new_n5363_), .B(new_n5347_), .Y(new_n5497_));
  NOR2X1   g05304(.A(new_n5363_), .B(new_n5347_), .Y(new_n5498_));
  OAI21X1  g05305(.A0(new_n5376_), .A1(new_n5498_), .B0(new_n5497_), .Y(new_n5499_));
  NOR2X1   g05306(.A(new_n5447_), .B(new_n5445_), .Y(new_n5500_));
  AOI21X1  g05307(.A0(new_n5473_), .A1(new_n5448_), .B0(new_n5500_), .Y(new_n5501_));
  AND2X1   g05308(.A(new_n5439_), .B(new_n5208_), .Y(new_n5502_));
  INVX1    g05309(.A(new_n5444_), .Y(new_n5503_));
  AOI21X1  g05310(.A0(new_n5503_), .A1(new_n5440_), .B0(new_n5502_), .Y(new_n5504_));
  NOR2X1   g05311(.A(new_n5255_), .B(new_n5244_), .Y(new_n5505_));
  AOI21X1  g05312(.A0(new_n5370_), .A1(new_n5369_), .B0(new_n5505_), .Y(new_n5506_));
  XOR2X1   g05313(.A(new_n5506_), .B(new_n5504_), .Y(new_n5507_));
  INVX1    g05314(.A(new_n5507_), .Y(new_n5508_));
  NOR2X1   g05315(.A(new_n5264_), .B(new_n5226_), .Y(new_n5509_));
  AOI21X1  g05316(.A0(new_n5367_), .A1(new_n5218_), .B0(new_n5509_), .Y(new_n5510_));
  XOR2X1   g05317(.A(new_n5510_), .B(new_n5508_), .Y(new_n5511_));
  INVX1    g05318(.A(new_n5511_), .Y(new_n5512_));
  OR2X1    g05319(.A(new_n5372_), .B(new_n5368_), .Y(new_n5513_));
  OAI21X1  g05320(.A0(new_n5374_), .A1(new_n5366_), .B0(new_n5513_), .Y(new_n5514_));
  XOR2X1   g05321(.A(new_n5514_), .B(new_n5512_), .Y(new_n5515_));
  XOR2X1   g05322(.A(new_n5515_), .B(new_n5501_), .Y(new_n5516_));
  XOR2X1   g05323(.A(new_n5516_), .B(new_n5499_), .Y(new_n5517_));
  XOR2X1   g05324(.A(new_n5517_), .B(new_n5496_), .Y(new_n5518_));
  XOR2X1   g05325(.A(new_n5518_), .B(new_n5492_), .Y(new_n5519_));
  AND2X1   g05326(.A(new_n5336_), .B(new_n5334_), .Y(new_n5520_));
  AOI21X1  g05327(.A0(new_n5337_), .A1(new_n5325_), .B0(new_n5520_), .Y(new_n5521_));
  AND2X1   g05328(.A(new_n5358_), .B(new_n5353_), .Y(new_n5522_));
  AOI21X1  g05329(.A0(new_n5361_), .A1(new_n5350_), .B0(new_n5522_), .Y(new_n5523_));
  NAND4X1  g05330(.A(\a[48] ), .B(\a[47] ), .C(\a[12] ), .D(\a[11] ), .Y(new_n5524_));
  NAND4X1  g05331(.A(\a[48] ), .B(\a[45] ), .C(\a[14] ), .D(\a[11] ), .Y(new_n5525_));
  AOI22X1  g05332(.A0(new_n5525_), .A1(new_n5524_), .B0(new_n3557_), .B1(new_n1282_), .Y(new_n5526_));
  AOI21X1  g05333(.A0(new_n3557_), .A1(new_n1282_), .B0(new_n5526_), .Y(new_n5527_));
  OAI22X1  g05334(.A0(new_n4041_), .A1(new_n453_), .B0(new_n3811_), .B1(new_n490_), .Y(new_n5528_));
  NOR3X1   g05335(.A(new_n5526_), .B(new_n3926_), .C(new_n488_), .Y(new_n5529_));
  AOI21X1  g05336(.A0(new_n5528_), .A1(new_n5527_), .B0(new_n5529_), .Y(new_n5530_));
  AND2X1   g05337(.A(\a[46] ), .B(\a[13] ), .Y(new_n5531_));
  INVX1    g05338(.A(new_n5531_), .Y(new_n5532_));
  AOI22X1  g05339(.A0(\a[31] ), .A1(\a[28] ), .B0(\a[30] ), .B1(\a[29] ), .Y(new_n5533_));
  NOR4X1   g05340(.A(new_n1704_), .B(new_n1684_), .C(new_n1803_), .D(new_n1431_), .Y(new_n5534_));
  NOR3X1   g05341(.A(new_n5533_), .B(new_n5534_), .C(new_n5532_), .Y(new_n5535_));
  INVX1    g05342(.A(new_n5533_), .Y(new_n5536_));
  AOI21X1  g05343(.A0(new_n5536_), .A1(new_n5531_), .B0(new_n5534_), .Y(new_n5537_));
  INVX1    g05344(.A(new_n5537_), .Y(new_n5538_));
  OAI22X1  g05345(.A0(new_n5538_), .A1(new_n5533_), .B0(new_n5535_), .B1(new_n5532_), .Y(new_n5539_));
  XOR2X1   g05346(.A(new_n5539_), .B(new_n5530_), .Y(new_n5540_));
  AND2X1   g05347(.A(\a[51] ), .B(\a[8] ), .Y(new_n5541_));
  AOI22X1  g05348(.A0(\a[43] ), .A1(\a[16] ), .B0(\a[42] ), .B1(\a[17] ), .Y(new_n5542_));
  INVX1    g05349(.A(new_n5542_), .Y(new_n5543_));
  NAND4X1  g05350(.A(\a[43] ), .B(\a[42] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n5544_));
  NAND3X1  g05351(.A(new_n5543_), .B(new_n5544_), .C(new_n5541_), .Y(new_n5545_));
  AOI22X1  g05352(.A0(new_n5543_), .A1(new_n5541_), .B0(new_n3462_), .B1(new_n792_), .Y(new_n5546_));
  AOI22X1  g05353(.A0(new_n5546_), .A1(new_n5543_), .B0(new_n5545_), .B1(new_n5541_), .Y(new_n5547_));
  XOR2X1   g05354(.A(new_n5547_), .B(new_n5540_), .Y(new_n5548_));
  INVX1    g05355(.A(new_n5429_), .Y(new_n5549_));
  AND2X1   g05356(.A(new_n5355_), .B(new_n2198_), .Y(new_n5550_));
  AOI22X1  g05357(.A0(\a[57] ), .A1(\a[2] ), .B0(\a[56] ), .B1(\a[3] ), .Y(new_n5551_));
  INVX1    g05358(.A(new_n5551_), .Y(new_n5552_));
  NAND2X1  g05359(.A(\a[57] ), .B(\a[1] ), .Y(new_n5553_));
  AND2X1   g05360(.A(\a[57] ), .B(\a[56] ), .Y(new_n5554_));
  AND2X1   g05361(.A(new_n5554_), .B(new_n231_), .Y(new_n5555_));
  OR4X1    g05362(.A(new_n5555_), .B(new_n5551_), .C(new_n5553_), .D(new_n2199_), .Y(new_n5556_));
  AOI21X1  g05363(.A0(new_n5552_), .A1(new_n5550_), .B0(new_n5555_), .Y(new_n5557_));
  AOI22X1  g05364(.A0(new_n5557_), .A1(new_n5552_), .B0(new_n5556_), .B1(new_n5550_), .Y(new_n5558_));
  XOR2X1   g05365(.A(new_n5558_), .B(new_n5549_), .Y(new_n5559_));
  AND2X1   g05366(.A(\a[40] ), .B(\a[4] ), .Y(new_n5560_));
  AND2X1   g05367(.A(\a[55] ), .B(\a[19] ), .Y(new_n5561_));
  AOI22X1  g05368(.A0(new_n5561_), .A1(new_n5560_), .B0(new_n5240_), .B1(new_n218_), .Y(new_n5562_));
  NOR4X1   g05369(.A(new_n4835_), .B(new_n3036_), .C(new_n752_), .D(new_n255_), .Y(new_n5563_));
  OR2X1    g05370(.A(new_n5563_), .B(new_n5562_), .Y(new_n5564_));
  AND2X1   g05371(.A(\a[55] ), .B(\a[4] ), .Y(new_n5565_));
  INVX1    g05372(.A(new_n5563_), .Y(new_n5566_));
  AND2X1   g05373(.A(new_n5566_), .B(new_n5562_), .Y(new_n5567_));
  OAI22X1  g05374(.A0(new_n4835_), .A1(new_n255_), .B0(new_n3036_), .B1(new_n752_), .Y(new_n5568_));
  AOI22X1  g05375(.A0(new_n5568_), .A1(new_n5567_), .B0(new_n5565_), .B1(new_n5564_), .Y(new_n5569_));
  XOR2X1   g05376(.A(new_n5569_), .B(new_n5559_), .Y(new_n5570_));
  XOR2X1   g05377(.A(new_n5570_), .B(new_n5548_), .Y(new_n5571_));
  XOR2X1   g05378(.A(new_n5571_), .B(new_n5523_), .Y(new_n5572_));
  XOR2X1   g05379(.A(new_n5572_), .B(new_n5521_), .Y(new_n5573_));
  AND2X1   g05380(.A(\a[52] ), .B(\a[18] ), .Y(new_n5574_));
  NAND4X1  g05381(.A(\a[53] ), .B(\a[41] ), .C(\a[18] ), .D(\a[6] ), .Y(new_n5575_));
  NAND4X1  g05382(.A(\a[53] ), .B(\a[52] ), .C(\a[7] ), .D(\a[6] ), .Y(new_n5576_));
  AOI22X1  g05383(.A0(new_n5576_), .A1(new_n5575_), .B0(new_n5574_), .B1(new_n3718_), .Y(new_n5577_));
  NAND4X1  g05384(.A(\a[52] ), .B(\a[41] ), .C(\a[18] ), .D(\a[7] ), .Y(new_n5578_));
  NAND3X1  g05385(.A(new_n5576_), .B(new_n5575_), .C(new_n5578_), .Y(new_n5579_));
  AOI22X1  g05386(.A0(\a[52] ), .A1(\a[7] ), .B0(\a[41] ), .B1(\a[18] ), .Y(new_n5580_));
  NAND2X1  g05387(.A(\a[53] ), .B(\a[6] ), .Y(new_n5581_));
  OAI22X1  g05388(.A0(new_n5581_), .A1(new_n5577_), .B0(new_n5580_), .B1(new_n5579_), .Y(new_n5582_));
  NOR3X1   g05389(.A(new_n544_), .B(new_n3915_), .C(new_n5268_), .Y(new_n5583_));
  NAND4X1  g05390(.A(\a[50] ), .B(\a[44] ), .C(\a[15] ), .D(\a[9] ), .Y(new_n5584_));
  NAND4X1  g05391(.A(\a[50] ), .B(\a[49] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n5585_));
  AOI21X1  g05392(.A0(new_n5585_), .A1(new_n5584_), .B0(new_n5583_), .Y(new_n5586_));
  NAND2X1  g05393(.A(\a[50] ), .B(\a[9] ), .Y(new_n5587_));
  AOI22X1  g05394(.A0(\a[49] ), .A1(\a[10] ), .B0(\a[44] ), .B1(\a[15] ), .Y(new_n5588_));
  NOR2X1   g05395(.A(new_n5586_), .B(new_n5583_), .Y(new_n5589_));
  INVX1    g05396(.A(new_n5589_), .Y(new_n5590_));
  OAI22X1  g05397(.A0(new_n5590_), .A1(new_n5588_), .B0(new_n5587_), .B1(new_n5586_), .Y(new_n5591_));
  XOR2X1   g05398(.A(new_n5591_), .B(new_n5582_), .Y(new_n5592_));
  NOR2X1   g05399(.A(new_n5356_), .B(new_n5354_), .Y(new_n5593_));
  NAND2X1  g05400(.A(new_n5356_), .B(new_n5354_), .Y(new_n5594_));
  OAI21X1  g05401(.A0(new_n5593_), .A1(new_n5283_), .B0(new_n5594_), .Y(new_n5595_));
  XOR2X1   g05402(.A(new_n5595_), .B(new_n5592_), .Y(new_n5596_));
  OR2X1    g05403(.A(new_n5329_), .B(new_n5327_), .Y(new_n5597_));
  OAI21X1  g05404(.A0(new_n5333_), .A1(new_n5331_), .B0(new_n5597_), .Y(new_n5598_));
  XOR2X1   g05405(.A(new_n5598_), .B(new_n5596_), .Y(new_n5599_));
  NAND4X1  g05406(.A(\a[39] ), .B(\a[37] ), .C(\a[22] ), .D(\a[20] ), .Y(new_n5600_));
  NAND4X1  g05407(.A(\a[39] ), .B(\a[38] ), .C(\a[21] ), .D(\a[20] ), .Y(new_n5601_));
  AOI22X1  g05408(.A0(new_n5601_), .A1(new_n5600_), .B0(new_n3164_), .B1(new_n1154_), .Y(new_n5602_));
  NAND4X1  g05409(.A(\a[38] ), .B(\a[37] ), .C(\a[22] ), .D(\a[21] ), .Y(new_n5603_));
  NAND3X1  g05410(.A(new_n5601_), .B(new_n5600_), .C(new_n5603_), .Y(new_n5604_));
  AOI22X1  g05411(.A0(\a[38] ), .A1(\a[21] ), .B0(\a[37] ), .B1(\a[22] ), .Y(new_n5605_));
  NAND2X1  g05412(.A(\a[39] ), .B(\a[20] ), .Y(new_n5606_));
  OAI22X1  g05413(.A0(new_n5606_), .A1(new_n5602_), .B0(new_n5605_), .B1(new_n5604_), .Y(new_n5607_));
  NAND4X1  g05414(.A(\a[36] ), .B(\a[34] ), .C(\a[25] ), .D(\a[23] ), .Y(new_n5608_));
  NAND4X1  g05415(.A(\a[36] ), .B(\a[35] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n5609_));
  AOI22X1  g05416(.A0(new_n5609_), .A1(new_n5608_), .B0(new_n2361_), .B1(new_n1532_), .Y(new_n5610_));
  NAND2X1  g05417(.A(\a[36] ), .B(\a[23] ), .Y(new_n5611_));
  AOI22X1  g05418(.A0(\a[35] ), .A1(\a[24] ), .B0(\a[34] ), .B1(\a[25] ), .Y(new_n5612_));
  AOI21X1  g05419(.A0(new_n2361_), .A1(new_n1532_), .B0(new_n5610_), .Y(new_n5613_));
  INVX1    g05420(.A(new_n5613_), .Y(new_n5614_));
  OAI22X1  g05421(.A0(new_n5614_), .A1(new_n5612_), .B0(new_n5611_), .B1(new_n5610_), .Y(new_n5615_));
  XOR2X1   g05422(.A(new_n5615_), .B(new_n5607_), .Y(new_n5616_));
  INVX1    g05423(.A(\a[59] ), .Y(new_n5617_));
  NOR4X1   g05424(.A(new_n5617_), .B(new_n2219_), .C(new_n1679_), .D(new_n194_), .Y(new_n5618_));
  NAND4X1  g05425(.A(\a[33] ), .B(\a[32] ), .C(\a[27] ), .D(\a[26] ), .Y(new_n5619_));
  NAND4X1  g05426(.A(\a[59] ), .B(\a[33] ), .C(\a[26] ), .D(\a[0] ), .Y(new_n5620_));
  AOI21X1  g05427(.A0(new_n5620_), .A1(new_n5619_), .B0(new_n5618_), .Y(new_n5621_));
  NAND2X1  g05428(.A(\a[33] ), .B(\a[26] ), .Y(new_n5622_));
  OR2X1    g05429(.A(new_n5621_), .B(new_n5618_), .Y(new_n5623_));
  AOI22X1  g05430(.A0(\a[59] ), .A1(\a[0] ), .B0(\a[32] ), .B1(\a[27] ), .Y(new_n5624_));
  OAI22X1  g05431(.A0(new_n5624_), .A1(new_n5623_), .B0(new_n5622_), .B1(new_n5621_), .Y(new_n5625_));
  XOR2X1   g05432(.A(new_n5625_), .B(new_n5616_), .Y(new_n5626_));
  XOR2X1   g05433(.A(new_n5626_), .B(new_n5599_), .Y(new_n5627_));
  XOR2X1   g05434(.A(new_n5627_), .B(new_n5573_), .Y(new_n5628_));
  AND2X1   g05435(.A(new_n5321_), .B(new_n5174_), .Y(new_n5629_));
  OAI21X1  g05436(.A0(new_n5322_), .A1(new_n5629_), .B0(new_n5338_), .Y(new_n5630_));
  OAI21X1  g05437(.A0(new_n5341_), .A1(new_n5339_), .B0(new_n5630_), .Y(new_n5631_));
  AND2X1   g05438(.A(new_n5463_), .B(new_n5456_), .Y(new_n5632_));
  AND2X1   g05439(.A(new_n5472_), .B(new_n5464_), .Y(new_n5633_));
  OR2X1    g05440(.A(new_n5633_), .B(new_n5632_), .Y(new_n5634_));
  INVX1    g05441(.A(new_n5416_), .Y(new_n5635_));
  OR2X1    g05442(.A(new_n5424_), .B(new_n5635_), .Y(new_n5636_));
  OAI21X1  g05443(.A0(new_n5431_), .A1(new_n5425_), .B0(new_n5636_), .Y(new_n5637_));
  XOR2X1   g05444(.A(new_n5637_), .B(new_n5634_), .Y(new_n5638_));
  INVX1    g05445(.A(new_n5397_), .Y(new_n5639_));
  OR2X1    g05446(.A(new_n5639_), .B(new_n5388_), .Y(new_n5640_));
  OAI21X1  g05447(.A0(new_n5407_), .A1(new_n5398_), .B0(new_n5640_), .Y(new_n5641_));
  XOR2X1   g05448(.A(new_n5641_), .B(new_n5638_), .Y(new_n5642_));
  XOR2X1   g05449(.A(new_n5431_), .B(new_n5425_), .Y(new_n5643_));
  NAND2X1  g05450(.A(new_n5643_), .B(new_n5408_), .Y(new_n5644_));
  OAI21X1  g05451(.A0(new_n5435_), .A1(new_n5433_), .B0(new_n5644_), .Y(new_n5645_));
  INVX1    g05452(.A(new_n5406_), .Y(new_n5646_));
  XOR2X1   g05453(.A(new_n5470_), .B(new_n5385_), .Y(new_n5647_));
  XOR2X1   g05454(.A(new_n5647_), .B(new_n5646_), .Y(new_n5648_));
  XOR2X1   g05455(.A(new_n5422_), .B(new_n5395_), .Y(new_n5649_));
  XOR2X1   g05456(.A(new_n5649_), .B(new_n5415_), .Y(new_n5650_));
  AOI21X1  g05457(.A0(\a[58] ), .A1(\a[1] ), .B0(\a[30] ), .Y(new_n5651_));
  AOI21X1  g05458(.A0(new_n1724_), .A1(\a[58] ), .B0(new_n5651_), .Y(new_n5652_));
  XOR2X1   g05459(.A(new_n5652_), .B(new_n5461_), .Y(new_n5653_));
  XOR2X1   g05460(.A(new_n5653_), .B(new_n5453_), .Y(new_n5654_));
  XOR2X1   g05461(.A(new_n5654_), .B(new_n5650_), .Y(new_n5655_));
  AND2X1   g05462(.A(new_n5655_), .B(new_n5648_), .Y(new_n5656_));
  INVX1    g05463(.A(new_n5650_), .Y(new_n5657_));
  NOR2X1   g05464(.A(new_n5654_), .B(new_n5657_), .Y(new_n5658_));
  AND2X1   g05465(.A(new_n5654_), .B(new_n5657_), .Y(new_n5659_));
  NOR3X1   g05466(.A(new_n5659_), .B(new_n5658_), .C(new_n5648_), .Y(new_n5660_));
  NOR2X1   g05467(.A(new_n5660_), .B(new_n5656_), .Y(new_n5661_));
  INVX1    g05468(.A(new_n5661_), .Y(new_n5662_));
  OR2X1    g05469(.A(new_n5662_), .B(new_n5645_), .Y(new_n5663_));
  XOR2X1   g05470(.A(new_n5661_), .B(new_n5645_), .Y(new_n5664_));
  AOI21X1  g05471(.A0(new_n5662_), .A1(new_n5645_), .B0(new_n5642_), .Y(new_n5665_));
  AOI22X1  g05472(.A0(new_n5665_), .A1(new_n5663_), .B0(new_n5664_), .B1(new_n5642_), .Y(new_n5666_));
  XOR2X1   g05473(.A(new_n5666_), .B(new_n5631_), .Y(new_n5667_));
  XOR2X1   g05474(.A(new_n5667_), .B(new_n5628_), .Y(new_n5668_));
  XOR2X1   g05475(.A(new_n5668_), .B(new_n5519_), .Y(new_n5669_));
  AND2X1   g05476(.A(new_n5342_), .B(new_n5320_), .Y(new_n5670_));
  INVX1    g05477(.A(new_n5477_), .Y(new_n5671_));
  AOI21X1  g05478(.A0(new_n5671_), .A1(new_n5343_), .B0(new_n5670_), .Y(new_n5672_));
  XOR2X1   g05479(.A(new_n5672_), .B(new_n5669_), .Y(new_n5673_));
  AOI21X1  g05480(.A0(new_n5485_), .A1(new_n5483_), .B0(new_n5479_), .Y(new_n5674_));
  XOR2X1   g05481(.A(new_n5674_), .B(new_n5673_), .Y(\asquared[60] ));
  AND2X1   g05482(.A(new_n5518_), .B(new_n5492_), .Y(new_n5676_));
  AOI21X1  g05483(.A0(new_n5668_), .A1(new_n5519_), .B0(new_n5676_), .Y(new_n5677_));
  INVX1    g05484(.A(new_n5677_), .Y(new_n5678_));
  AND2X1   g05485(.A(new_n5666_), .B(new_n5631_), .Y(new_n5679_));
  AOI21X1  g05486(.A0(new_n5667_), .A1(new_n5628_), .B0(new_n5679_), .Y(new_n5680_));
  NOR2X1   g05487(.A(new_n5572_), .B(new_n5521_), .Y(new_n5681_));
  AOI21X1  g05488(.A0(new_n5627_), .A1(new_n5573_), .B0(new_n5681_), .Y(new_n5682_));
  INVX1    g05489(.A(new_n5682_), .Y(new_n5683_));
  AND2X1   g05490(.A(new_n5661_), .B(new_n5645_), .Y(new_n5684_));
  AOI21X1  g05491(.A0(new_n5664_), .A1(new_n5642_), .B0(new_n5684_), .Y(new_n5685_));
  NOR2X1   g05492(.A(new_n5422_), .B(new_n5395_), .Y(new_n5686_));
  AOI21X1  g05493(.A0(new_n5649_), .A1(new_n5415_), .B0(new_n5686_), .Y(new_n5687_));
  AOI21X1  g05494(.A0(new_n5383_), .A1(new_n5384_), .B0(new_n5470_), .Y(new_n5688_));
  AOI21X1  g05495(.A0(new_n5647_), .A1(new_n5646_), .B0(new_n5688_), .Y(new_n5689_));
  XOR2X1   g05496(.A(new_n5689_), .B(new_n5687_), .Y(new_n5690_));
  OR2X1    g05497(.A(new_n5558_), .B(new_n5429_), .Y(new_n5691_));
  OAI21X1  g05498(.A0(new_n5569_), .A1(new_n5559_), .B0(new_n5691_), .Y(new_n5692_));
  XOR2X1   g05499(.A(new_n5692_), .B(new_n5690_), .Y(new_n5693_));
  INVX1    g05500(.A(new_n5693_), .Y(new_n5694_));
  AND2X1   g05501(.A(new_n5637_), .B(new_n5634_), .Y(new_n5695_));
  AOI21X1  g05502(.A0(new_n5641_), .A1(new_n5638_), .B0(new_n5695_), .Y(new_n5696_));
  XOR2X1   g05503(.A(new_n5696_), .B(new_n5694_), .Y(new_n5697_));
  AND2X1   g05504(.A(new_n5598_), .B(new_n5596_), .Y(new_n5698_));
  AOI21X1  g05505(.A0(new_n5626_), .A1(new_n5599_), .B0(new_n5698_), .Y(new_n5699_));
  XOR2X1   g05506(.A(new_n5699_), .B(new_n5697_), .Y(new_n5700_));
  XOR2X1   g05507(.A(new_n5700_), .B(new_n5685_), .Y(new_n5701_));
  XOR2X1   g05508(.A(new_n5701_), .B(new_n5683_), .Y(new_n5702_));
  XOR2X1   g05509(.A(new_n5702_), .B(new_n5680_), .Y(new_n5703_));
  AND2X1   g05510(.A(new_n5654_), .B(new_n5650_), .Y(new_n5704_));
  OR2X1    g05511(.A(new_n5656_), .B(new_n5704_), .Y(new_n5705_));
  NAND3X1  g05512(.A(\a[58] ), .B(\a[30] ), .C(\a[1] ), .Y(new_n5706_));
  AND2X1   g05513(.A(\a[60] ), .B(\a[0] ), .Y(new_n5707_));
  XOR2X1   g05514(.A(new_n5707_), .B(new_n5706_), .Y(new_n5708_));
  AND2X1   g05515(.A(\a[59] ), .B(\a[1] ), .Y(new_n5709_));
  XOR2X1   g05516(.A(new_n5709_), .B(new_n2430_), .Y(new_n5710_));
  XOR2X1   g05517(.A(new_n5710_), .B(new_n5708_), .Y(new_n5711_));
  NAND4X1  g05518(.A(\a[33] ), .B(\a[32] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n5712_));
  NAND4X1  g05519(.A(\a[37] ), .B(\a[33] ), .C(\a[27] ), .D(\a[23] ), .Y(new_n5713_));
  NOR4X1   g05520(.A(new_n2345_), .B(new_n2219_), .C(new_n1431_), .D(new_n1216_), .Y(new_n5714_));
  AOI21X1  g05521(.A0(new_n5713_), .A1(new_n5712_), .B0(new_n5714_), .Y(new_n5715_));
  NAND2X1  g05522(.A(\a[33] ), .B(\a[27] ), .Y(new_n5716_));
  OR2X1    g05523(.A(new_n5715_), .B(new_n5714_), .Y(new_n5717_));
  AOI22X1  g05524(.A0(\a[37] ), .A1(\a[23] ), .B0(\a[32] ), .B1(\a[28] ), .Y(new_n5718_));
  OAI22X1  g05525(.A0(new_n5718_), .A1(new_n5717_), .B0(new_n5716_), .B1(new_n5715_), .Y(new_n5719_));
  XOR2X1   g05526(.A(new_n5719_), .B(new_n5711_), .Y(new_n5720_));
  NAND2X1  g05527(.A(new_n5652_), .B(new_n5461_), .Y(new_n5721_));
  OAI21X1  g05528(.A0(new_n5452_), .A1(new_n5449_), .B0(new_n5653_), .Y(new_n5722_));
  NAND2X1  g05529(.A(new_n5722_), .B(new_n5721_), .Y(new_n5723_));
  XOR2X1   g05530(.A(new_n5723_), .B(new_n5720_), .Y(new_n5724_));
  INVX1    g05531(.A(new_n5724_), .Y(new_n5725_));
  NOR4X1   g05532(.A(new_n4354_), .B(new_n3096_), .C(new_n675_), .D(new_n413_), .Y(new_n5726_));
  NAND4X1  g05533(.A(\a[53] ), .B(\a[52] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n5727_));
  NAND4X1  g05534(.A(\a[53] ), .B(\a[42] ), .C(\a[18] ), .D(\a[7] ), .Y(new_n5728_));
  AOI21X1  g05535(.A0(new_n5728_), .A1(new_n5727_), .B0(new_n5726_), .Y(new_n5729_));
  OR2X1    g05536(.A(new_n5729_), .B(new_n5726_), .Y(new_n5730_));
  AOI22X1  g05537(.A0(\a[52] ), .A1(\a[8] ), .B0(\a[42] ), .B1(\a[18] ), .Y(new_n5731_));
  NAND2X1  g05538(.A(\a[53] ), .B(\a[7] ), .Y(new_n5732_));
  OAI22X1  g05539(.A0(new_n5732_), .A1(new_n5729_), .B0(new_n5731_), .B1(new_n5730_), .Y(new_n5733_));
  AND2X1   g05540(.A(\a[46] ), .B(\a[14] ), .Y(new_n5734_));
  INVX1    g05541(.A(new_n5734_), .Y(new_n5735_));
  NAND4X1  g05542(.A(\a[48] ), .B(\a[46] ), .C(\a[14] ), .D(\a[12] ), .Y(new_n5736_));
  NAND4X1  g05543(.A(\a[47] ), .B(\a[46] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n5737_));
  AOI22X1  g05544(.A0(new_n5737_), .A1(new_n5736_), .B0(new_n4272_), .B1(new_n586_), .Y(new_n5738_));
  AOI21X1  g05545(.A0(new_n4272_), .A1(new_n586_), .B0(new_n5738_), .Y(new_n5739_));
  INVX1    g05546(.A(new_n5739_), .Y(new_n5740_));
  AOI22X1  g05547(.A0(\a[48] ), .A1(\a[12] ), .B0(\a[47] ), .B1(\a[13] ), .Y(new_n5741_));
  OAI22X1  g05548(.A0(new_n5741_), .A1(new_n5740_), .B0(new_n5738_), .B1(new_n5735_), .Y(new_n5742_));
  XOR2X1   g05549(.A(new_n5742_), .B(new_n5733_), .Y(new_n5743_));
  AND2X1   g05550(.A(\a[19] ), .B(\a[5] ), .Y(new_n5744_));
  AND2X1   g05551(.A(\a[55] ), .B(\a[41] ), .Y(new_n5745_));
  AOI22X1  g05552(.A0(new_n5745_), .A1(new_n5744_), .B0(new_n5240_), .B1(new_n295_), .Y(new_n5746_));
  NOR4X1   g05553(.A(new_n4835_), .B(new_n3081_), .C(new_n752_), .D(new_n230_), .Y(new_n5747_));
  AND2X1   g05554(.A(\a[55] ), .B(\a[5] ), .Y(new_n5748_));
  OAI21X1  g05555(.A0(new_n5747_), .A1(new_n5746_), .B0(new_n5748_), .Y(new_n5749_));
  INVX1    g05556(.A(new_n5747_), .Y(new_n5750_));
  AND2X1   g05557(.A(new_n5750_), .B(new_n5746_), .Y(new_n5751_));
  INVX1    g05558(.A(new_n5751_), .Y(new_n5752_));
  AOI22X1  g05559(.A0(\a[54] ), .A1(\a[6] ), .B0(\a[41] ), .B1(\a[19] ), .Y(new_n5753_));
  OAI21X1  g05560(.A0(new_n5753_), .A1(new_n5752_), .B0(new_n5749_), .Y(new_n5754_));
  INVX1    g05561(.A(new_n5754_), .Y(new_n5755_));
  XOR2X1   g05562(.A(new_n5755_), .B(new_n5743_), .Y(new_n5756_));
  XOR2X1   g05563(.A(new_n5756_), .B(new_n5725_), .Y(new_n5757_));
  XOR2X1   g05564(.A(new_n5757_), .B(new_n5705_), .Y(new_n5758_));
  INVX1    g05565(.A(new_n5758_), .Y(new_n5759_));
  NAND2X1  g05566(.A(new_n5514_), .B(new_n5511_), .Y(new_n5760_));
  OAI21X1  g05567(.A0(new_n5515_), .A1(new_n5501_), .B0(new_n5760_), .Y(new_n5761_));
  NAND4X1  g05568(.A(\a[58] ), .B(\a[56] ), .C(\a[4] ), .D(\a[2] ), .Y(new_n5762_));
  NAND4X1  g05569(.A(\a[58] ), .B(\a[57] ), .C(\a[3] ), .D(\a[2] ), .Y(new_n5763_));
  AOI22X1  g05570(.A0(new_n5763_), .A1(new_n5762_), .B0(new_n5554_), .B1(new_n294_), .Y(new_n5764_));
  NAND4X1  g05571(.A(\a[57] ), .B(\a[56] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n5765_));
  NAND3X1  g05572(.A(new_n5763_), .B(new_n5762_), .C(new_n5765_), .Y(new_n5766_));
  AOI22X1  g05573(.A0(\a[57] ), .A1(\a[3] ), .B0(\a[56] ), .B1(\a[4] ), .Y(new_n5767_));
  NAND2X1  g05574(.A(\a[58] ), .B(\a[2] ), .Y(new_n5768_));
  OAI22X1  g05575(.A0(new_n5768_), .A1(new_n5764_), .B0(new_n5767_), .B1(new_n5766_), .Y(new_n5769_));
  NAND4X1  g05576(.A(\a[40] ), .B(\a[38] ), .C(\a[22] ), .D(\a[20] ), .Y(new_n5770_));
  NAND4X1  g05577(.A(\a[40] ), .B(\a[39] ), .C(\a[21] ), .D(\a[20] ), .Y(new_n5771_));
  AOI22X1  g05578(.A0(new_n5771_), .A1(new_n5770_), .B0(new_n3503_), .B1(new_n1154_), .Y(new_n5772_));
  NAND2X1  g05579(.A(\a[40] ), .B(\a[20] ), .Y(new_n5773_));
  AOI22X1  g05580(.A0(\a[39] ), .A1(\a[21] ), .B0(\a[38] ), .B1(\a[22] ), .Y(new_n5774_));
  AOI21X1  g05581(.A0(new_n3503_), .A1(new_n1154_), .B0(new_n5772_), .Y(new_n5775_));
  INVX1    g05582(.A(new_n5775_), .Y(new_n5776_));
  OAI22X1  g05583(.A0(new_n5776_), .A1(new_n5774_), .B0(new_n5773_), .B1(new_n5772_), .Y(new_n5777_));
  XOR2X1   g05584(.A(new_n5777_), .B(new_n5769_), .Y(new_n5778_));
  AOI22X1  g05585(.A0(new_n4695_), .A1(new_n1650_), .B0(new_n2682_), .B1(new_n1532_), .Y(new_n5779_));
  AOI21X1  g05586(.A0(new_n2361_), .A1(new_n1770_), .B0(new_n5779_), .Y(new_n5780_));
  AND2X1   g05587(.A(\a[36] ), .B(\a[24] ), .Y(new_n5781_));
  INVX1    g05588(.A(new_n5781_), .Y(new_n5782_));
  AOI21X1  g05589(.A0(new_n2361_), .A1(new_n1770_), .B0(new_n5780_), .Y(new_n5783_));
  INVX1    g05590(.A(new_n5783_), .Y(new_n5784_));
  AOI22X1  g05591(.A0(\a[35] ), .A1(\a[25] ), .B0(\a[34] ), .B1(\a[26] ), .Y(new_n5785_));
  OAI22X1  g05592(.A0(new_n5785_), .A1(new_n5784_), .B0(new_n5782_), .B1(new_n5780_), .Y(new_n5786_));
  XOR2X1   g05593(.A(new_n5786_), .B(new_n5778_), .Y(new_n5787_));
  NOR2X1   g05594(.A(new_n5506_), .B(new_n5504_), .Y(new_n5788_));
  INVX1    g05595(.A(new_n5788_), .Y(new_n5789_));
  OAI21X1  g05596(.A0(new_n5510_), .A1(new_n5508_), .B0(new_n5789_), .Y(new_n5790_));
  INVX1    g05597(.A(new_n5790_), .Y(new_n5791_));
  XOR2X1   g05598(.A(new_n5791_), .B(new_n5787_), .Y(new_n5792_));
  NOR4X1   g05599(.A(new_n4349_), .B(new_n5268_), .C(new_n571_), .D(new_n341_), .Y(new_n5793_));
  AND2X1   g05600(.A(\a[51] ), .B(\a[17] ), .Y(new_n5794_));
  AOI22X1  g05601(.A0(new_n5794_), .A1(new_n4442_), .B0(new_n4992_), .B1(new_n792_), .Y(new_n5795_));
  AND2X1   g05602(.A(\a[43] ), .B(\a[17] ), .Y(new_n5796_));
  OAI21X1  g05603(.A0(new_n5795_), .A1(new_n5793_), .B0(new_n5796_), .Y(new_n5797_));
  INVX1    g05604(.A(new_n5793_), .Y(new_n5798_));
  AND2X1   g05605(.A(new_n5795_), .B(new_n5798_), .Y(new_n5799_));
  INVX1    g05606(.A(new_n5799_), .Y(new_n5800_));
  AOI22X1  g05607(.A0(\a[51] ), .A1(\a[9] ), .B0(\a[44] ), .B1(\a[16] ), .Y(new_n5801_));
  OAI21X1  g05608(.A0(new_n5801_), .A1(new_n5800_), .B0(new_n5797_), .Y(new_n5802_));
  XOR2X1   g05609(.A(new_n5802_), .B(new_n5527_), .Y(new_n5803_));
  NOR3X1   g05610(.A(new_n633_), .B(new_n3915_), .C(new_n3811_), .Y(new_n5804_));
  NOR3X1   g05611(.A(new_n544_), .B(new_n4983_), .C(new_n3811_), .Y(new_n5805_));
  AOI21X1  g05612(.A0(new_n4321_), .A1(new_n1002_), .B0(new_n5805_), .Y(new_n5806_));
  OR2X1    g05613(.A(new_n5806_), .B(new_n5804_), .Y(new_n5807_));
  AND2X1   g05614(.A(\a[50] ), .B(\a[10] ), .Y(new_n5808_));
  OAI22X1  g05615(.A0(new_n3915_), .A1(new_n488_), .B0(new_n3811_), .B1(new_n549_), .Y(new_n5809_));
  INVX1    g05616(.A(new_n5804_), .Y(new_n5810_));
  AND2X1   g05617(.A(new_n5806_), .B(new_n5810_), .Y(new_n5811_));
  AOI22X1  g05618(.A0(new_n5811_), .A1(new_n5809_), .B0(new_n5808_), .B1(new_n5807_), .Y(new_n5812_));
  XOR2X1   g05619(.A(new_n5812_), .B(new_n5803_), .Y(new_n5813_));
  INVX1    g05620(.A(new_n5813_), .Y(new_n5814_));
  XOR2X1   g05621(.A(new_n5814_), .B(new_n5792_), .Y(new_n5815_));
  XOR2X1   g05622(.A(new_n5815_), .B(new_n5761_), .Y(new_n5816_));
  XOR2X1   g05623(.A(new_n5816_), .B(new_n5759_), .Y(new_n5817_));
  AND2X1   g05624(.A(new_n5516_), .B(new_n5499_), .Y(new_n5818_));
  AOI21X1  g05625(.A0(new_n5517_), .A1(new_n5496_), .B0(new_n5818_), .Y(new_n5819_));
  AND2X1   g05626(.A(new_n5591_), .B(new_n5582_), .Y(new_n5820_));
  AOI21X1  g05627(.A0(new_n5595_), .A1(new_n5592_), .B0(new_n5820_), .Y(new_n5821_));
  INVX1    g05628(.A(new_n5567_), .Y(new_n5822_));
  XOR2X1   g05629(.A(new_n5604_), .B(new_n5822_), .Y(new_n5823_));
  XOR2X1   g05630(.A(new_n5823_), .B(new_n5613_), .Y(new_n5824_));
  INVX1    g05631(.A(new_n5557_), .Y(new_n5825_));
  XOR2X1   g05632(.A(new_n5623_), .B(new_n5825_), .Y(new_n5826_));
  XOR2X1   g05633(.A(new_n5826_), .B(new_n5590_), .Y(new_n5827_));
  INVX1    g05634(.A(new_n5827_), .Y(new_n5828_));
  XOR2X1   g05635(.A(new_n5828_), .B(new_n5824_), .Y(new_n5829_));
  INVX1    g05636(.A(new_n5829_), .Y(new_n5830_));
  XOR2X1   g05637(.A(new_n5830_), .B(new_n5821_), .Y(new_n5831_));
  NOR2X1   g05638(.A(new_n5570_), .B(new_n5548_), .Y(new_n5832_));
  NAND2X1  g05639(.A(new_n5570_), .B(new_n5548_), .Y(new_n5833_));
  OAI21X1  g05640(.A0(new_n5832_), .A1(new_n5523_), .B0(new_n5833_), .Y(new_n5834_));
  AND2X1   g05641(.A(new_n5831_), .B(new_n5834_), .Y(new_n5835_));
  INVX1    g05642(.A(new_n5835_), .Y(new_n5836_));
  NAND2X1  g05643(.A(new_n5836_), .B(new_n5831_), .Y(new_n5837_));
  INVX1    g05644(.A(new_n5546_), .Y(new_n5838_));
  XOR2X1   g05645(.A(new_n5579_), .B(new_n5838_), .Y(new_n5839_));
  XOR2X1   g05646(.A(new_n5839_), .B(new_n5537_), .Y(new_n5840_));
  AND2X1   g05647(.A(new_n5615_), .B(new_n5607_), .Y(new_n5841_));
  AOI21X1  g05648(.A0(new_n5625_), .A1(new_n5616_), .B0(new_n5841_), .Y(new_n5842_));
  XOR2X1   g05649(.A(new_n5842_), .B(new_n5840_), .Y(new_n5843_));
  AND2X1   g05650(.A(new_n5528_), .B(new_n5527_), .Y(new_n5844_));
  OAI21X1  g05651(.A0(new_n5529_), .A1(new_n5844_), .B0(new_n5539_), .Y(new_n5845_));
  OAI21X1  g05652(.A0(new_n5547_), .A1(new_n5540_), .B0(new_n5845_), .Y(new_n5846_));
  XOR2X1   g05653(.A(new_n5846_), .B(new_n5843_), .Y(new_n5847_));
  XOR2X1   g05654(.A(new_n5831_), .B(new_n5834_), .Y(new_n5848_));
  AND2X1   g05655(.A(new_n5848_), .B(new_n5847_), .Y(new_n5849_));
  AOI21X1  g05656(.A0(new_n5836_), .A1(new_n5834_), .B0(new_n5847_), .Y(new_n5850_));
  AOI21X1  g05657(.A0(new_n5850_), .A1(new_n5837_), .B0(new_n5849_), .Y(new_n5851_));
  AND2X1   g05658(.A(new_n5851_), .B(new_n5819_), .Y(new_n5852_));
  XOR2X1   g05659(.A(new_n5851_), .B(new_n5819_), .Y(new_n5853_));
  OAI21X1  g05660(.A0(new_n5851_), .A1(new_n5819_), .B0(new_n5817_), .Y(new_n5854_));
  OAI22X1  g05661(.A0(new_n5854_), .A1(new_n5852_), .B0(new_n5853_), .B1(new_n5817_), .Y(new_n5855_));
  XOR2X1   g05662(.A(new_n5855_), .B(new_n5703_), .Y(new_n5856_));
  XOR2X1   g05663(.A(new_n5856_), .B(new_n5678_), .Y(new_n5857_));
  INVX1    g05664(.A(new_n5519_), .Y(new_n5858_));
  XOR2X1   g05665(.A(new_n5668_), .B(new_n5858_), .Y(new_n5859_));
  AND2X1   g05666(.A(new_n5672_), .B(new_n5859_), .Y(new_n5860_));
  OR2X1    g05667(.A(new_n5672_), .B(new_n5859_), .Y(new_n5861_));
  OAI21X1  g05668(.A0(new_n5674_), .A1(new_n5860_), .B0(new_n5861_), .Y(new_n5862_));
  XOR2X1   g05669(.A(new_n5862_), .B(new_n5857_), .Y(\asquared[61] ));
  INVX1    g05670(.A(new_n5702_), .Y(new_n5864_));
  OR2X1    g05671(.A(new_n5864_), .B(new_n5680_), .Y(new_n5865_));
  OAI21X1  g05672(.A0(new_n5855_), .A1(new_n5703_), .B0(new_n5865_), .Y(new_n5866_));
  AND2X1   g05673(.A(new_n5815_), .B(new_n5761_), .Y(new_n5867_));
  AND2X1   g05674(.A(new_n5816_), .B(new_n5758_), .Y(new_n5868_));
  OR2X1    g05675(.A(new_n5868_), .B(new_n5867_), .Y(new_n5869_));
  NOR2X1   g05676(.A(new_n5842_), .B(new_n5840_), .Y(new_n5870_));
  AOI21X1  g05677(.A0(new_n5846_), .A1(new_n5843_), .B0(new_n5870_), .Y(new_n5871_));
  AOI22X1  g05678(.A0(\a[54] ), .A1(\a[7] ), .B0(\a[53] ), .B1(\a[8] ), .Y(new_n5872_));
  AND2X1   g05679(.A(\a[42] ), .B(\a[19] ), .Y(new_n5873_));
  INVX1    g05680(.A(new_n5873_), .Y(new_n5874_));
  AND2X1   g05681(.A(new_n5238_), .B(new_n325_), .Y(new_n5875_));
  NOR3X1   g05682(.A(new_n5874_), .B(new_n5875_), .C(new_n5872_), .Y(new_n5876_));
  NOR2X1   g05683(.A(new_n5876_), .B(new_n5875_), .Y(new_n5877_));
  INVX1    g05684(.A(new_n5877_), .Y(new_n5878_));
  OAI22X1  g05685(.A0(new_n5878_), .A1(new_n5872_), .B0(new_n5876_), .B1(new_n5874_), .Y(new_n5879_));
  AND2X1   g05686(.A(\a[52] ), .B(\a[44] ), .Y(new_n5880_));
  AND2X1   g05687(.A(new_n5880_), .B(new_n1226_), .Y(new_n5881_));
  AOI22X1  g05688(.A0(new_n5574_), .A1(new_n4442_), .B0(new_n4992_), .B1(new_n796_), .Y(new_n5882_));
  OR2X1    g05689(.A(new_n5882_), .B(new_n5881_), .Y(new_n5883_));
  AND2X1   g05690(.A(\a[43] ), .B(\a[18] ), .Y(new_n5884_));
  INVX1    g05691(.A(new_n5880_), .Y(new_n5885_));
  OAI21X1  g05692(.A0(new_n5885_), .A1(new_n1227_), .B0(new_n5882_), .Y(new_n5886_));
  INVX1    g05693(.A(new_n5886_), .Y(new_n5887_));
  OAI22X1  g05694(.A0(new_n4354_), .A1(new_n341_), .B0(new_n5268_), .B1(new_n616_), .Y(new_n5888_));
  AOI22X1  g05695(.A0(new_n5888_), .A1(new_n5887_), .B0(new_n5884_), .B1(new_n5883_), .Y(new_n5889_));
  XOR2X1   g05696(.A(new_n5889_), .B(new_n5879_), .Y(new_n5890_));
  OAI22X1  g05697(.A0(new_n4915_), .A1(new_n3483_), .B0(new_n4914_), .B1(new_n3570_), .Y(new_n5891_));
  OAI21X1  g05698(.A0(new_n2919_), .A1(new_n1672_), .B0(new_n5891_), .Y(new_n5892_));
  AND2X1   g05699(.A(\a[35] ), .B(\a[26] ), .Y(new_n5893_));
  AOI21X1  g05700(.A0(new_n2918_), .A1(new_n1671_), .B0(new_n5891_), .Y(new_n5894_));
  OAI22X1  g05701(.A0(new_n2028_), .A1(new_n1679_), .B0(new_n1851_), .B1(new_n1431_), .Y(new_n5895_));
  AOI22X1  g05702(.A0(new_n5895_), .A1(new_n5894_), .B0(new_n5893_), .B1(new_n5892_), .Y(new_n5896_));
  XOR2X1   g05703(.A(new_n5896_), .B(new_n5890_), .Y(new_n5897_));
  INVX1    g05704(.A(new_n5897_), .Y(new_n5898_));
  OR2X1    g05705(.A(new_n5828_), .B(new_n5824_), .Y(new_n5899_));
  OAI21X1  g05706(.A0(new_n5830_), .A1(new_n5821_), .B0(new_n5899_), .Y(new_n5900_));
  XOR2X1   g05707(.A(new_n5900_), .B(new_n5898_), .Y(new_n5901_));
  XOR2X1   g05708(.A(new_n5901_), .B(new_n5871_), .Y(new_n5902_));
  AND2X1   g05709(.A(new_n5790_), .B(new_n5787_), .Y(new_n5903_));
  NOR2X1   g05710(.A(new_n5814_), .B(new_n5792_), .Y(new_n5904_));
  OR2X1    g05711(.A(new_n5904_), .B(new_n5903_), .Y(new_n5905_));
  AND2X1   g05712(.A(new_n5623_), .B(new_n5825_), .Y(new_n5906_));
  AOI21X1  g05713(.A0(new_n5826_), .A1(new_n5590_), .B0(new_n5906_), .Y(new_n5907_));
  AND2X1   g05714(.A(new_n5579_), .B(new_n5838_), .Y(new_n5908_));
  AOI21X1  g05715(.A0(new_n5839_), .A1(new_n5538_), .B0(new_n5908_), .Y(new_n5909_));
  AND2X1   g05716(.A(\a[38] ), .B(\a[23] ), .Y(new_n5910_));
  INVX1    g05717(.A(new_n5910_), .Y(new_n5911_));
  AOI22X1  g05718(.A0(\a[58] ), .A1(\a[3] ), .B0(\a[57] ), .B1(\a[4] ), .Y(new_n5912_));
  NOR3X1   g05719(.A(new_n217_), .B(new_n5379_), .C(new_n5441_), .Y(new_n5913_));
  NOR3X1   g05720(.A(new_n5912_), .B(new_n5913_), .C(new_n5911_), .Y(new_n5914_));
  INVX1    g05721(.A(new_n5912_), .Y(new_n5915_));
  AOI21X1  g05722(.A0(new_n5915_), .A1(new_n5910_), .B0(new_n5913_), .Y(new_n5916_));
  INVX1    g05723(.A(new_n5916_), .Y(new_n5917_));
  OAI22X1  g05724(.A0(new_n5917_), .A1(new_n5912_), .B0(new_n5914_), .B1(new_n5911_), .Y(new_n5918_));
  XOR2X1   g05725(.A(new_n5918_), .B(new_n5909_), .Y(new_n5919_));
  XOR2X1   g05726(.A(new_n5919_), .B(new_n5907_), .Y(new_n5920_));
  INVX1    g05727(.A(new_n5802_), .Y(new_n5921_));
  OR2X1    g05728(.A(new_n5812_), .B(new_n5803_), .Y(new_n5922_));
  OAI21X1  g05729(.A0(new_n5921_), .A1(new_n5527_), .B0(new_n5922_), .Y(new_n5923_));
  AND2X1   g05730(.A(new_n5604_), .B(new_n5822_), .Y(new_n5924_));
  AOI21X1  g05731(.A0(new_n5823_), .A1(new_n5614_), .B0(new_n5924_), .Y(new_n5925_));
  AND2X1   g05732(.A(new_n5709_), .B(new_n2429_), .Y(new_n5926_));
  AND2X1   g05733(.A(\a[60] ), .B(\a[1] ), .Y(new_n5927_));
  XOR2X1   g05734(.A(new_n5927_), .B(\a[31] ), .Y(new_n5928_));
  XOR2X1   g05735(.A(new_n5928_), .B(new_n5926_), .Y(new_n5929_));
  XOR2X1   g05736(.A(new_n5929_), .B(new_n5739_), .Y(new_n5930_));
  XOR2X1   g05737(.A(new_n5930_), .B(new_n5925_), .Y(new_n5931_));
  XOR2X1   g05738(.A(new_n5931_), .B(new_n5923_), .Y(new_n5932_));
  XOR2X1   g05739(.A(new_n5932_), .B(new_n5920_), .Y(new_n5933_));
  AND2X1   g05740(.A(new_n5932_), .B(new_n5920_), .Y(new_n5934_));
  INVX1    g05741(.A(new_n5934_), .Y(new_n5935_));
  AND2X1   g05742(.A(new_n5935_), .B(new_n5920_), .Y(new_n5936_));
  AND2X1   g05743(.A(new_n5935_), .B(new_n5932_), .Y(new_n5937_));
  NOR4X1   g05744(.A(new_n5937_), .B(new_n5936_), .C(new_n5904_), .D(new_n5903_), .Y(new_n5938_));
  AOI21X1  g05745(.A0(new_n5933_), .A1(new_n5905_), .B0(new_n5938_), .Y(new_n5939_));
  XOR2X1   g05746(.A(new_n5939_), .B(new_n5902_), .Y(new_n5940_));
  XOR2X1   g05747(.A(new_n5940_), .B(new_n5869_), .Y(new_n5941_));
  AND2X1   g05748(.A(new_n5850_), .B(new_n5837_), .Y(new_n5942_));
  NOR3X1   g05749(.A(new_n5942_), .B(new_n5849_), .C(new_n5819_), .Y(new_n5943_));
  NOR2X1   g05750(.A(new_n5853_), .B(new_n5817_), .Y(new_n5944_));
  OAI21X1  g05751(.A0(new_n5944_), .A1(new_n5943_), .B0(new_n5941_), .Y(new_n5945_));
  NAND2X1  g05752(.A(new_n5945_), .B(new_n5941_), .Y(new_n5946_));
  NOR2X1   g05753(.A(new_n5944_), .B(new_n5943_), .Y(new_n5947_));
  XOR2X1   g05754(.A(new_n5941_), .B(new_n5947_), .Y(new_n5948_));
  NOR2X1   g05755(.A(new_n5756_), .B(new_n5725_), .Y(new_n5949_));
  AOI21X1  g05756(.A0(new_n5757_), .A1(new_n5705_), .B0(new_n5949_), .Y(new_n5950_));
  XOR2X1   g05757(.A(new_n5800_), .B(new_n5730_), .Y(new_n5951_));
  INVX1    g05758(.A(\a[60] ), .Y(new_n5952_));
  NOR3X1   g05759(.A(new_n5706_), .B(new_n5952_), .C(new_n194_), .Y(new_n5953_));
  NOR2X1   g05760(.A(new_n5710_), .B(new_n5708_), .Y(new_n5954_));
  NOR2X1   g05761(.A(new_n5954_), .B(new_n5953_), .Y(new_n5955_));
  INVX1    g05762(.A(new_n5955_), .Y(new_n5956_));
  XOR2X1   g05763(.A(new_n5956_), .B(new_n5951_), .Y(new_n5957_));
  INVX1    g05764(.A(new_n5957_), .Y(new_n5958_));
  AND2X1   g05765(.A(new_n5742_), .B(new_n5733_), .Y(new_n5959_));
  AOI21X1  g05766(.A0(new_n5754_), .A1(new_n5743_), .B0(new_n5959_), .Y(new_n5960_));
  XOR2X1   g05767(.A(new_n5960_), .B(new_n5958_), .Y(new_n5961_));
  AND2X1   g05768(.A(new_n5719_), .B(new_n5711_), .Y(new_n5962_));
  AOI21X1  g05769(.A0(new_n5723_), .A1(new_n5720_), .B0(new_n5962_), .Y(new_n5963_));
  XOR2X1   g05770(.A(new_n5963_), .B(new_n5961_), .Y(new_n5964_));
  AND2X1   g05771(.A(new_n5777_), .B(new_n5769_), .Y(new_n5965_));
  AOI21X1  g05772(.A0(new_n5786_), .A1(new_n5778_), .B0(new_n5965_), .Y(new_n5966_));
  XOR2X1   g05773(.A(new_n5784_), .B(new_n5717_), .Y(new_n5967_));
  XOR2X1   g05774(.A(new_n5967_), .B(new_n5775_), .Y(new_n5968_));
  INVX1    g05775(.A(new_n5811_), .Y(new_n5969_));
  XOR2X1   g05776(.A(new_n5766_), .B(new_n5752_), .Y(new_n5970_));
  XOR2X1   g05777(.A(new_n5970_), .B(new_n5969_), .Y(new_n5971_));
  INVX1    g05778(.A(new_n5971_), .Y(new_n5972_));
  XOR2X1   g05779(.A(new_n5972_), .B(new_n5968_), .Y(new_n5973_));
  XOR2X1   g05780(.A(new_n5973_), .B(new_n5966_), .Y(new_n5974_));
  AND2X1   g05781(.A(new_n5974_), .B(new_n5964_), .Y(new_n5975_));
  NOR2X1   g05782(.A(new_n5974_), .B(new_n5964_), .Y(new_n5976_));
  NOR3X1   g05783(.A(new_n5976_), .B(new_n5975_), .C(new_n5950_), .Y(new_n5977_));
  OR2X1    g05784(.A(new_n5977_), .B(new_n5976_), .Y(new_n5978_));
  OAI22X1  g05785(.A0(new_n5978_), .A1(new_n5975_), .B0(new_n5977_), .B1(new_n5950_), .Y(new_n5979_));
  NOR2X1   g05786(.A(new_n5700_), .B(new_n5685_), .Y(new_n5980_));
  AOI21X1  g05787(.A0(new_n5701_), .A1(new_n5683_), .B0(new_n5980_), .Y(new_n5981_));
  XOR2X1   g05788(.A(new_n5981_), .B(new_n5979_), .Y(new_n5982_));
  OR2X1    g05789(.A(new_n5849_), .B(new_n5835_), .Y(new_n5983_));
  NOR2X1   g05790(.A(new_n5696_), .B(new_n5694_), .Y(new_n5984_));
  INVX1    g05791(.A(new_n5984_), .Y(new_n5985_));
  INVX1    g05792(.A(new_n5697_), .Y(new_n5986_));
  OAI21X1  g05793(.A0(new_n5699_), .A1(new_n5986_), .B0(new_n5985_), .Y(new_n5987_));
  NAND2X1  g05794(.A(\a[45] ), .B(\a[16] ), .Y(new_n5988_));
  NAND4X1  g05795(.A(\a[51] ), .B(\a[46] ), .C(\a[15] ), .D(\a[10] ), .Y(new_n5989_));
  NAND4X1  g05796(.A(\a[46] ), .B(\a[45] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n5990_));
  NAND4X1  g05797(.A(\a[51] ), .B(\a[45] ), .C(\a[16] ), .D(\a[10] ), .Y(new_n5991_));
  NAND2X1  g05798(.A(new_n5991_), .B(new_n5990_), .Y(new_n5992_));
  AND2X1   g05799(.A(new_n5992_), .B(new_n5989_), .Y(new_n5993_));
  NAND3X1  g05800(.A(new_n5991_), .B(new_n5990_), .C(new_n5989_), .Y(new_n5994_));
  AOI22X1  g05801(.A0(\a[51] ), .A1(\a[10] ), .B0(\a[46] ), .B1(\a[15] ), .Y(new_n5995_));
  OAI22X1  g05802(.A0(new_n5995_), .A1(new_n5994_), .B0(new_n5993_), .B1(new_n5988_), .Y(new_n5996_));
  NOR3X1   g05803(.A(new_n585_), .B(new_n3915_), .C(new_n4041_), .Y(new_n5997_));
  NAND4X1  g05804(.A(\a[50] ), .B(\a[47] ), .C(\a[14] ), .D(\a[11] ), .Y(new_n5998_));
  NAND4X1  g05805(.A(\a[50] ), .B(\a[49] ), .C(\a[12] ), .D(\a[11] ), .Y(new_n5999_));
  AOI21X1  g05806(.A0(new_n5999_), .A1(new_n5998_), .B0(new_n5997_), .Y(new_n6000_));
  NAND2X1  g05807(.A(\a[50] ), .B(\a[11] ), .Y(new_n6001_));
  NOR2X1   g05808(.A(new_n6000_), .B(new_n5997_), .Y(new_n6002_));
  INVX1    g05809(.A(new_n6002_), .Y(new_n6003_));
  AOI22X1  g05810(.A0(\a[49] ), .A1(\a[12] ), .B0(\a[47] ), .B1(\a[14] ), .Y(new_n6004_));
  OAI22X1  g05811(.A0(new_n6004_), .A1(new_n6003_), .B0(new_n6001_), .B1(new_n6000_), .Y(new_n6005_));
  XOR2X1   g05812(.A(new_n6005_), .B(new_n5996_), .Y(new_n6006_));
  AOI22X1  g05813(.A0(\a[32] ), .A1(\a[29] ), .B0(\a[31] ), .B1(\a[30] ), .Y(new_n6007_));
  AND2X1   g05814(.A(\a[48] ), .B(\a[13] ), .Y(new_n6008_));
  AND2X1   g05815(.A(new_n2671_), .B(new_n2196_), .Y(new_n6009_));
  OAI21X1  g05816(.A0(new_n6007_), .A1(new_n6009_), .B0(new_n6008_), .Y(new_n6010_));
  INVX1    g05817(.A(new_n6007_), .Y(new_n6011_));
  AOI21X1  g05818(.A0(new_n6011_), .A1(new_n6008_), .B0(new_n6009_), .Y(new_n6012_));
  INVX1    g05819(.A(new_n6012_), .Y(new_n6013_));
  OAI21X1  g05820(.A0(new_n6013_), .A1(new_n6007_), .B0(new_n6010_), .Y(new_n6014_));
  XOR2X1   g05821(.A(new_n6014_), .B(new_n6006_), .Y(new_n6015_));
  NOR2X1   g05822(.A(new_n5689_), .B(new_n5687_), .Y(new_n6016_));
  AOI21X1  g05823(.A0(new_n5692_), .A1(new_n5690_), .B0(new_n6016_), .Y(new_n6017_));
  XOR2X1   g05824(.A(new_n6017_), .B(new_n6015_), .Y(new_n6018_));
  AND2X1   g05825(.A(\a[59] ), .B(\a[5] ), .Y(new_n6019_));
  AND2X1   g05826(.A(\a[61] ), .B(\a[59] ), .Y(new_n6020_));
  AND2X1   g05827(.A(new_n6020_), .B(new_n197_), .Y(new_n6021_));
  INVX1    g05828(.A(\a[56] ), .Y(new_n6022_));
  INVX1    g05829(.A(\a[61] ), .Y(new_n6023_));
  NOR4X1   g05830(.A(new_n6023_), .B(new_n6022_), .C(new_n255_), .D(new_n194_), .Y(new_n6024_));
  NOR2X1   g05831(.A(new_n6024_), .B(new_n6021_), .Y(new_n6025_));
  AOI21X1  g05832(.A0(new_n6019_), .A1(new_n5387_), .B0(new_n6025_), .Y(new_n6026_));
  AOI21X1  g05833(.A0(new_n6019_), .A1(new_n5387_), .B0(new_n6026_), .Y(new_n6027_));
  OAI22X1  g05834(.A0(new_n5617_), .A1(new_n200_), .B0(new_n6022_), .B1(new_n255_), .Y(new_n6028_));
  NOR3X1   g05835(.A(new_n6026_), .B(new_n6023_), .C(new_n194_), .Y(new_n6029_));
  AOI21X1  g05836(.A0(new_n6028_), .A1(new_n6027_), .B0(new_n6029_), .Y(new_n6030_));
  AND2X1   g05837(.A(\a[55] ), .B(\a[6] ), .Y(new_n6031_));
  INVX1    g05838(.A(new_n6031_), .Y(new_n6032_));
  AOI22X1  g05839(.A0(\a[41] ), .A1(\a[20] ), .B0(\a[40] ), .B1(\a[21] ), .Y(new_n6033_));
  AND2X1   g05840(.A(new_n4404_), .B(new_n1236_), .Y(new_n6034_));
  NOR3X1   g05841(.A(new_n6033_), .B(new_n6034_), .C(new_n6032_), .Y(new_n6035_));
  INVX1    g05842(.A(new_n6033_), .Y(new_n6036_));
  AOI21X1  g05843(.A0(new_n6036_), .A1(new_n6031_), .B0(new_n6034_), .Y(new_n6037_));
  INVX1    g05844(.A(new_n6037_), .Y(new_n6038_));
  OAI22X1  g05845(.A0(new_n6038_), .A1(new_n6033_), .B0(new_n6035_), .B1(new_n6032_), .Y(new_n6039_));
  XOR2X1   g05846(.A(new_n6039_), .B(new_n6030_), .Y(new_n6040_));
  INVX1    g05847(.A(new_n6040_), .Y(new_n6041_));
  NAND4X1  g05848(.A(\a[39] ), .B(\a[36] ), .C(\a[25] ), .D(\a[22] ), .Y(new_n6042_));
  NAND4X1  g05849(.A(\a[39] ), .B(\a[37] ), .C(\a[24] ), .D(\a[22] ), .Y(new_n6043_));
  AOI22X1  g05850(.A0(new_n6043_), .A1(new_n6042_), .B0(new_n3330_), .B1(new_n1532_), .Y(new_n6044_));
  NOR3X1   g05851(.A(new_n6044_), .B(new_n2652_), .C(new_n1086_), .Y(new_n6045_));
  OAI22X1  g05852(.A0(new_n2345_), .A1(new_n1185_), .B0(new_n2583_), .B1(new_n1326_), .Y(new_n6046_));
  AOI21X1  g05853(.A0(new_n3330_), .A1(new_n1532_), .B0(new_n6044_), .Y(new_n6047_));
  AOI21X1  g05854(.A0(new_n6047_), .A1(new_n6046_), .B0(new_n6045_), .Y(new_n6048_));
  XOR2X1   g05855(.A(new_n6048_), .B(new_n6041_), .Y(new_n6049_));
  XOR2X1   g05856(.A(new_n6049_), .B(new_n6018_), .Y(new_n6050_));
  XOR2X1   g05857(.A(new_n6050_), .B(new_n5987_), .Y(new_n6051_));
  XOR2X1   g05858(.A(new_n6051_), .B(new_n5983_), .Y(new_n6052_));
  XOR2X1   g05859(.A(new_n6052_), .B(new_n5982_), .Y(new_n6053_));
  NOR2X1   g05860(.A(new_n6053_), .B(new_n5948_), .Y(new_n6054_));
  OR2X1    g05861(.A(new_n5941_), .B(new_n5947_), .Y(new_n6055_));
  AND2X1   g05862(.A(new_n6053_), .B(new_n6055_), .Y(new_n6056_));
  AOI21X1  g05863(.A0(new_n6056_), .A1(new_n5946_), .B0(new_n6054_), .Y(new_n6057_));
  AND2X1   g05864(.A(new_n6057_), .B(new_n5866_), .Y(new_n6058_));
  NOR2X1   g05865(.A(new_n6057_), .B(new_n5866_), .Y(new_n6059_));
  OR2X1    g05866(.A(new_n6059_), .B(new_n6058_), .Y(new_n6060_));
  NOR2X1   g05867(.A(new_n5856_), .B(new_n5678_), .Y(new_n6061_));
  INVX1    g05868(.A(new_n6061_), .Y(new_n6062_));
  AND2X1   g05869(.A(new_n5856_), .B(new_n5678_), .Y(new_n6063_));
  AOI21X1  g05870(.A0(new_n5862_), .A1(new_n6062_), .B0(new_n6063_), .Y(new_n6064_));
  XOR2X1   g05871(.A(new_n6064_), .B(new_n6060_), .Y(\asquared[62] ));
  OAI21X1  g05872(.A0(new_n6053_), .A1(new_n5948_), .B0(new_n5945_), .Y(new_n6066_));
  AND2X1   g05873(.A(new_n5766_), .B(new_n5752_), .Y(new_n6067_));
  AOI21X1  g05874(.A0(new_n5970_), .A1(new_n5969_), .B0(new_n6067_), .Y(new_n6068_));
  INVX1    g05875(.A(new_n6068_), .Y(new_n6069_));
  INVX1    g05876(.A(new_n6039_), .Y(new_n6070_));
  OR2X1    g05877(.A(new_n6070_), .B(new_n6030_), .Y(new_n6071_));
  OAI21X1  g05878(.A0(new_n6048_), .A1(new_n6040_), .B0(new_n6071_), .Y(new_n6072_));
  XOR2X1   g05879(.A(new_n6072_), .B(new_n6069_), .Y(new_n6073_));
  AND2X1   g05880(.A(new_n6005_), .B(new_n5996_), .Y(new_n6074_));
  AOI21X1  g05881(.A0(new_n6014_), .A1(new_n6006_), .B0(new_n6074_), .Y(new_n6075_));
  XOR2X1   g05882(.A(new_n6075_), .B(new_n6073_), .Y(new_n6076_));
  XOR2X1   g05883(.A(new_n6037_), .B(new_n6027_), .Y(new_n6077_));
  XOR2X1   g05884(.A(new_n6077_), .B(new_n5878_), .Y(new_n6078_));
  INVX1    g05885(.A(new_n6078_), .Y(new_n6079_));
  INVX1    g05886(.A(new_n6047_), .Y(new_n6080_));
  XOR2X1   g05887(.A(new_n5916_), .B(new_n5894_), .Y(new_n6081_));
  XOR2X1   g05888(.A(new_n6081_), .B(new_n6080_), .Y(new_n6082_));
  AND2X1   g05889(.A(\a[61] ), .B(\a[1] ), .Y(new_n6083_));
  XOR2X1   g05890(.A(new_n6083_), .B(new_n1787_), .Y(new_n6084_));
  INVX1    g05891(.A(new_n6084_), .Y(new_n6085_));
  XOR2X1   g05892(.A(new_n6085_), .B(new_n6012_), .Y(new_n6086_));
  INVX1    g05893(.A(new_n6086_), .Y(new_n6087_));
  XOR2X1   g05894(.A(new_n6087_), .B(new_n6002_), .Y(new_n6088_));
  XOR2X1   g05895(.A(new_n6088_), .B(new_n6082_), .Y(new_n6089_));
  XOR2X1   g05896(.A(new_n6089_), .B(new_n6079_), .Y(new_n6090_));
  XOR2X1   g05897(.A(new_n6090_), .B(new_n6076_), .Y(new_n6091_));
  NAND2X1  g05898(.A(new_n5900_), .B(new_n5897_), .Y(new_n6092_));
  OAI21X1  g05899(.A0(new_n5901_), .A1(new_n5871_), .B0(new_n6092_), .Y(new_n6093_));
  XOR2X1   g05900(.A(new_n6093_), .B(new_n6091_), .Y(new_n6094_));
  AND2X1   g05901(.A(new_n5972_), .B(new_n5968_), .Y(new_n6095_));
  OR2X1    g05902(.A(new_n5972_), .B(new_n5968_), .Y(new_n6096_));
  OAI21X1  g05903(.A0(new_n6095_), .A1(new_n5966_), .B0(new_n6096_), .Y(new_n6097_));
  NOR2X1   g05904(.A(new_n5930_), .B(new_n5925_), .Y(new_n6098_));
  AOI21X1  g05905(.A0(new_n5931_), .A1(new_n5923_), .B0(new_n6098_), .Y(new_n6099_));
  XOR2X1   g05906(.A(new_n6099_), .B(new_n6097_), .Y(new_n6100_));
  NOR2X1   g05907(.A(new_n5960_), .B(new_n5958_), .Y(new_n6101_));
  INVX1    g05908(.A(new_n6101_), .Y(new_n6102_));
  INVX1    g05909(.A(new_n5961_), .Y(new_n6103_));
  OAI21X1  g05910(.A0(new_n5963_), .A1(new_n6103_), .B0(new_n6102_), .Y(new_n6104_));
  XOR2X1   g05911(.A(new_n6104_), .B(new_n6100_), .Y(new_n6105_));
  AND2X1   g05912(.A(new_n6050_), .B(new_n5987_), .Y(new_n6106_));
  AOI21X1  g05913(.A0(new_n6051_), .A1(new_n5983_), .B0(new_n6106_), .Y(new_n6107_));
  XOR2X1   g05914(.A(new_n6107_), .B(new_n6105_), .Y(new_n6108_));
  XOR2X1   g05915(.A(new_n6108_), .B(new_n6094_), .Y(new_n6109_));
  INVX1    g05916(.A(new_n5981_), .Y(new_n6110_));
  AND2X1   g05917(.A(new_n6110_), .B(new_n5979_), .Y(new_n6111_));
  INVX1    g05918(.A(new_n6052_), .Y(new_n6112_));
  NOR2X1   g05919(.A(new_n6112_), .B(new_n5982_), .Y(new_n6113_));
  OAI21X1  g05920(.A0(new_n6113_), .A1(new_n6111_), .B0(new_n6109_), .Y(new_n6114_));
  NAND2X1  g05921(.A(new_n6114_), .B(new_n6109_), .Y(new_n6115_));
  AND2X1   g05922(.A(new_n5939_), .B(new_n5902_), .Y(new_n6116_));
  AOI21X1  g05923(.A0(new_n5940_), .A1(new_n5869_), .B0(new_n6116_), .Y(new_n6117_));
  XOR2X1   g05924(.A(new_n5994_), .B(new_n5886_), .Y(new_n6118_));
  AND2X1   g05925(.A(\a[58] ), .B(\a[57] ), .Y(new_n6119_));
  AND2X1   g05926(.A(\a[59] ), .B(\a[57] ), .Y(new_n6120_));
  AND2X1   g05927(.A(\a[59] ), .B(\a[58] ), .Y(new_n6121_));
  AOI22X1  g05928(.A0(new_n6121_), .A1(new_n294_), .B0(new_n6120_), .B1(new_n272_), .Y(new_n6122_));
  AOI21X1  g05929(.A0(new_n6119_), .A1(new_n218_), .B0(new_n6122_), .Y(new_n6123_));
  NAND2X1  g05930(.A(\a[59] ), .B(\a[3] ), .Y(new_n6124_));
  NAND4X1  g05931(.A(\a[58] ), .B(\a[57] ), .C(\a[5] ), .D(\a[4] ), .Y(new_n6125_));
  AND2X1   g05932(.A(new_n6122_), .B(new_n6125_), .Y(new_n6126_));
  INVX1    g05933(.A(new_n6126_), .Y(new_n6127_));
  AOI22X1  g05934(.A0(\a[58] ), .A1(\a[4] ), .B0(\a[57] ), .B1(\a[5] ), .Y(new_n6128_));
  OAI22X1  g05935(.A0(new_n6128_), .A1(new_n6127_), .B0(new_n6124_), .B1(new_n6123_), .Y(new_n6129_));
  XOR2X1   g05936(.A(new_n6129_), .B(new_n6118_), .Y(new_n6130_));
  INVX1    g05937(.A(new_n5879_), .Y(new_n6131_));
  OR2X1    g05938(.A(new_n5889_), .B(new_n6131_), .Y(new_n6132_));
  OAI21X1  g05939(.A0(new_n5896_), .A1(new_n5890_), .B0(new_n6132_), .Y(new_n6133_));
  XOR2X1   g05940(.A(new_n6133_), .B(new_n6130_), .Y(new_n6134_));
  INVX1    g05941(.A(new_n5918_), .Y(new_n6135_));
  OR2X1    g05942(.A(new_n6135_), .B(new_n5909_), .Y(new_n6136_));
  OAI21X1  g05943(.A0(new_n5919_), .A1(new_n5907_), .B0(new_n6136_), .Y(new_n6137_));
  XOR2X1   g05944(.A(new_n6137_), .B(new_n6134_), .Y(new_n6138_));
  AND2X1   g05945(.A(new_n5800_), .B(new_n5730_), .Y(new_n6139_));
  AOI21X1  g05946(.A0(new_n5956_), .A1(new_n5951_), .B0(new_n6139_), .Y(new_n6140_));
  AND2X1   g05947(.A(new_n5928_), .B(new_n5926_), .Y(new_n6141_));
  AOI21X1  g05948(.A0(new_n5929_), .A1(new_n5740_), .B0(new_n6141_), .Y(new_n6142_));
  XOR2X1   g05949(.A(new_n6142_), .B(new_n6140_), .Y(new_n6143_));
  INVX1    g05950(.A(new_n6143_), .Y(new_n6144_));
  AND2X1   g05951(.A(new_n5784_), .B(new_n5717_), .Y(new_n6145_));
  AOI21X1  g05952(.A0(new_n5967_), .A1(new_n5776_), .B0(new_n6145_), .Y(new_n6146_));
  XOR2X1   g05953(.A(new_n6146_), .B(new_n6144_), .Y(new_n6147_));
  INVX1    g05954(.A(new_n6015_), .Y(new_n6148_));
  NOR2X1   g05955(.A(new_n6017_), .B(new_n6148_), .Y(new_n6149_));
  NOR2X1   g05956(.A(new_n6049_), .B(new_n6018_), .Y(new_n6150_));
  NOR2X1   g05957(.A(new_n6150_), .B(new_n6149_), .Y(new_n6151_));
  OR2X1    g05958(.A(new_n6151_), .B(new_n6147_), .Y(new_n6152_));
  INVX1    g05959(.A(new_n6147_), .Y(new_n6153_));
  XOR2X1   g05960(.A(new_n6151_), .B(new_n6153_), .Y(new_n6154_));
  AOI21X1  g05961(.A0(new_n6151_), .A1(new_n6147_), .B0(new_n6138_), .Y(new_n6155_));
  AOI22X1  g05962(.A0(new_n6155_), .A1(new_n6152_), .B0(new_n6154_), .B1(new_n6138_), .Y(new_n6156_));
  XOR2X1   g05963(.A(new_n6156_), .B(new_n6117_), .Y(new_n6157_));
  AOI21X1  g05964(.A0(new_n5933_), .A1(new_n5905_), .B0(new_n5934_), .Y(new_n6158_));
  AOI22X1  g05965(.A0(\a[54] ), .A1(\a[8] ), .B0(\a[44] ), .B1(\a[18] ), .Y(new_n6159_));
  NOR4X1   g05966(.A(new_n4835_), .B(new_n5268_), .C(new_n675_), .D(new_n413_), .Y(new_n6160_));
  NAND4X1  g05967(.A(\a[44] ), .B(\a[43] ), .C(\a[19] ), .D(\a[18] ), .Y(new_n6161_));
  NAND4X1  g05968(.A(\a[54] ), .B(\a[43] ), .C(\a[19] ), .D(\a[8] ), .Y(new_n6162_));
  AOI21X1  g05969(.A0(new_n6162_), .A1(new_n6161_), .B0(new_n6160_), .Y(new_n6163_));
  NOR2X1   g05970(.A(new_n6163_), .B(new_n6160_), .Y(new_n6164_));
  INVX1    g05971(.A(new_n6164_), .Y(new_n6165_));
  NAND2X1  g05972(.A(\a[43] ), .B(\a[19] ), .Y(new_n6166_));
  OAI22X1  g05973(.A0(new_n6166_), .A1(new_n6163_), .B0(new_n6165_), .B1(new_n6159_), .Y(new_n6167_));
  AOI22X1  g05974(.A0(new_n2361_), .A1(new_n1671_), .B0(new_n2120_), .B1(new_n1484_), .Y(new_n6168_));
  AOI21X1  g05975(.A0(new_n2918_), .A1(new_n1674_), .B0(new_n6168_), .Y(new_n6169_));
  NAND2X1  g05976(.A(\a[35] ), .B(\a[27] ), .Y(new_n6170_));
  OAI21X1  g05977(.A0(new_n2919_), .A1(new_n1675_), .B0(new_n6168_), .Y(new_n6171_));
  AOI22X1  g05978(.A0(\a[34] ), .A1(\a[28] ), .B0(\a[33] ), .B1(\a[29] ), .Y(new_n6172_));
  OAI22X1  g05979(.A0(new_n6172_), .A1(new_n6171_), .B0(new_n6170_), .B1(new_n6169_), .Y(new_n6173_));
  XOR2X1   g05980(.A(new_n6173_), .B(new_n6167_), .Y(new_n6174_));
  AOI22X1  g05981(.A0(new_n4077_), .A1(new_n1394_), .B0(new_n2663_), .B1(new_n1530_), .Y(new_n6175_));
  AOI21X1  g05982(.A0(new_n3503_), .A1(new_n1219_), .B0(new_n6175_), .Y(new_n6176_));
  AND2X1   g05983(.A(\a[40] ), .B(\a[22] ), .Y(new_n6177_));
  INVX1    g05984(.A(new_n6177_), .Y(new_n6178_));
  INVX1    g05985(.A(new_n2663_), .Y(new_n6179_));
  INVX1    g05986(.A(new_n4077_), .Y(new_n6180_));
  OAI22X1  g05987(.A0(new_n6180_), .A1(new_n1395_), .B0(new_n6179_), .B1(new_n1531_), .Y(new_n6181_));
  AOI21X1  g05988(.A0(new_n3503_), .A1(new_n1219_), .B0(new_n6181_), .Y(new_n6182_));
  INVX1    g05989(.A(new_n6182_), .Y(new_n6183_));
  AOI22X1  g05990(.A0(\a[39] ), .A1(\a[23] ), .B0(\a[38] ), .B1(\a[24] ), .Y(new_n6184_));
  OAI22X1  g05991(.A0(new_n6184_), .A1(new_n6183_), .B0(new_n6178_), .B1(new_n6176_), .Y(new_n6185_));
  INVX1    g05992(.A(new_n6185_), .Y(new_n6186_));
  XOR2X1   g05993(.A(new_n6186_), .B(new_n6174_), .Y(new_n6187_));
  AOI22X1  g05994(.A0(\a[62] ), .A1(\a[0] ), .B0(\a[60] ), .B1(\a[2] ), .Y(new_n6188_));
  INVX1    g05995(.A(new_n6188_), .Y(new_n6189_));
  AND2X1   g05996(.A(new_n5927_), .B(\a[31] ), .Y(new_n6190_));
  AND2X1   g05997(.A(\a[62] ), .B(\a[60] ), .Y(new_n6191_));
  AND2X1   g05998(.A(new_n6191_), .B(new_n197_), .Y(new_n6192_));
  AOI21X1  g05999(.A0(new_n6189_), .A1(new_n6190_), .B0(new_n6192_), .Y(new_n6193_));
  NAND2X1  g06000(.A(new_n6193_), .B(new_n6189_), .Y(new_n6194_));
  OAI21X1  g06001(.A0(new_n6192_), .A1(new_n6188_), .B0(new_n6190_), .Y(new_n6195_));
  AND2X1   g06002(.A(new_n6195_), .B(new_n6194_), .Y(new_n6196_));
  AND2X1   g06003(.A(\a[41] ), .B(\a[21] ), .Y(new_n6197_));
  AOI22X1  g06004(.A0(\a[37] ), .A1(\a[25] ), .B0(\a[36] ), .B1(\a[26] ), .Y(new_n6198_));
  INVX1    g06005(.A(new_n6198_), .Y(new_n6199_));
  NAND4X1  g06006(.A(\a[37] ), .B(\a[36] ), .C(\a[26] ), .D(\a[25] ), .Y(new_n6200_));
  NAND3X1  g06007(.A(new_n6199_), .B(new_n6200_), .C(new_n6197_), .Y(new_n6201_));
  AOI22X1  g06008(.A0(new_n6199_), .A1(new_n6197_), .B0(new_n3330_), .B1(new_n1770_), .Y(new_n6202_));
  AOI22X1  g06009(.A0(new_n6202_), .A1(new_n6199_), .B0(new_n6201_), .B1(new_n6197_), .Y(new_n6203_));
  XOR2X1   g06010(.A(new_n6203_), .B(new_n6196_), .Y(new_n6204_));
  NOR4X1   g06011(.A(new_n4354_), .B(new_n3811_), .C(new_n616_), .D(new_n570_), .Y(new_n6205_));
  AND2X1   g06012(.A(\a[53] ), .B(\a[17] ), .Y(new_n6206_));
  AOI22X1  g06013(.A0(new_n6206_), .A1(new_n4747_), .B0(new_n5048_), .B1(new_n881_), .Y(new_n6207_));
  OR2X1    g06014(.A(new_n6207_), .B(new_n6205_), .Y(new_n6208_));
  AND2X1   g06015(.A(\a[53] ), .B(\a[9] ), .Y(new_n6209_));
  INVX1    g06016(.A(new_n6205_), .Y(new_n6210_));
  AND2X1   g06017(.A(new_n6207_), .B(new_n6210_), .Y(new_n6211_));
  OAI22X1  g06018(.A0(new_n4354_), .A1(new_n570_), .B0(new_n3811_), .B1(new_n616_), .Y(new_n6212_));
  AOI22X1  g06019(.A0(new_n6212_), .A1(new_n6211_), .B0(new_n6209_), .B1(new_n6208_), .Y(new_n6213_));
  XOR2X1   g06020(.A(new_n6213_), .B(new_n6204_), .Y(new_n6214_));
  NOR3X1   g06021(.A(new_n633_), .B(new_n4349_), .C(new_n4041_), .Y(new_n6215_));
  AND2X1   g06022(.A(\a[51] ), .B(\a[46] ), .Y(new_n6216_));
  AOI22X1  g06023(.A0(new_n6216_), .A1(new_n1345_), .B0(new_n3893_), .B1(new_n689_), .Y(new_n6217_));
  NOR2X1   g06024(.A(new_n6217_), .B(new_n6215_), .Y(new_n6218_));
  INVX1    g06025(.A(new_n6215_), .Y(new_n6219_));
  AND2X1   g06026(.A(new_n6217_), .B(new_n6219_), .Y(new_n6220_));
  INVX1    g06027(.A(new_n6220_), .Y(new_n6221_));
  AOI22X1  g06028(.A0(\a[51] ), .A1(\a[11] ), .B0(\a[47] ), .B1(\a[15] ), .Y(new_n6222_));
  NAND2X1  g06029(.A(\a[46] ), .B(\a[16] ), .Y(new_n6223_));
  OAI22X1  g06030(.A0(new_n6223_), .A1(new_n6218_), .B0(new_n6222_), .B1(new_n6221_), .Y(new_n6224_));
  NAND4X1  g06031(.A(\a[50] ), .B(\a[48] ), .C(\a[14] ), .D(\a[12] ), .Y(new_n6225_));
  NAND4X1  g06032(.A(\a[50] ), .B(\a[49] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n6226_));
  AOI22X1  g06033(.A0(new_n6226_), .A1(new_n6225_), .B0(new_n4274_), .B1(new_n582_), .Y(new_n6227_));
  NAND2X1  g06034(.A(\a[50] ), .B(\a[12] ), .Y(new_n6228_));
  AOI22X1  g06035(.A0(\a[49] ), .A1(\a[13] ), .B0(\a[48] ), .B1(\a[14] ), .Y(new_n6229_));
  AOI21X1  g06036(.A0(new_n4274_), .A1(new_n582_), .B0(new_n6227_), .Y(new_n6230_));
  INVX1    g06037(.A(new_n6230_), .Y(new_n6231_));
  OAI22X1  g06038(.A0(new_n6231_), .A1(new_n6229_), .B0(new_n6228_), .B1(new_n6227_), .Y(new_n6232_));
  XOR2X1   g06039(.A(new_n6232_), .B(new_n6224_), .Y(new_n6233_));
  AND2X1   g06040(.A(\a[42] ), .B(\a[20] ), .Y(new_n6234_));
  INVX1    g06041(.A(new_n6234_), .Y(new_n6235_));
  AOI22X1  g06042(.A0(\a[56] ), .A1(\a[6] ), .B0(\a[55] ), .B1(\a[7] ), .Y(new_n6236_));
  AND2X1   g06043(.A(\a[56] ), .B(\a[55] ), .Y(new_n6237_));
  AND2X1   g06044(.A(new_n6237_), .B(new_n375_), .Y(new_n6238_));
  NOR3X1   g06045(.A(new_n6236_), .B(new_n6238_), .C(new_n6235_), .Y(new_n6239_));
  INVX1    g06046(.A(new_n6236_), .Y(new_n6240_));
  AOI21X1  g06047(.A0(new_n6240_), .A1(new_n6234_), .B0(new_n6238_), .Y(new_n6241_));
  INVX1    g06048(.A(new_n6241_), .Y(new_n6242_));
  OAI22X1  g06049(.A0(new_n6242_), .A1(new_n6236_), .B0(new_n6239_), .B1(new_n6235_), .Y(new_n6243_));
  INVX1    g06050(.A(new_n6243_), .Y(new_n6244_));
  XOR2X1   g06051(.A(new_n6244_), .B(new_n6233_), .Y(new_n6245_));
  XOR2X1   g06052(.A(new_n6245_), .B(new_n6214_), .Y(new_n6246_));
  INVX1    g06053(.A(new_n6246_), .Y(new_n6247_));
  XOR2X1   g06054(.A(new_n6247_), .B(new_n6187_), .Y(new_n6248_));
  XOR2X1   g06055(.A(new_n6248_), .B(new_n6158_), .Y(new_n6249_));
  XOR2X1   g06056(.A(new_n6249_), .B(new_n5978_), .Y(new_n6250_));
  INVX1    g06057(.A(new_n6250_), .Y(new_n6251_));
  XOR2X1   g06058(.A(new_n6251_), .B(new_n6157_), .Y(new_n6252_));
  NOR2X1   g06059(.A(new_n6113_), .B(new_n6111_), .Y(new_n6253_));
  XOR2X1   g06060(.A(new_n6109_), .B(new_n6253_), .Y(new_n6254_));
  NOR2X1   g06061(.A(new_n6254_), .B(new_n6252_), .Y(new_n6255_));
  OR2X1    g06062(.A(new_n6109_), .B(new_n6253_), .Y(new_n6256_));
  AND2X1   g06063(.A(new_n6256_), .B(new_n6252_), .Y(new_n6257_));
  AOI21X1  g06064(.A0(new_n6257_), .A1(new_n6115_), .B0(new_n6255_), .Y(new_n6258_));
  AND2X1   g06065(.A(new_n6258_), .B(new_n6066_), .Y(new_n6259_));
  INVX1    g06066(.A(new_n6259_), .Y(new_n6260_));
  INVX1    g06067(.A(new_n6058_), .Y(new_n6261_));
  OAI21X1  g06068(.A0(new_n6064_), .A1(new_n6059_), .B0(new_n6261_), .Y(new_n6262_));
  NOR2X1   g06069(.A(new_n6258_), .B(new_n6066_), .Y(new_n6263_));
  INVX1    g06070(.A(new_n6263_), .Y(new_n6264_));
  AOI21X1  g06071(.A0(new_n6264_), .A1(new_n6260_), .B0(new_n6262_), .Y(new_n6265_));
  AND2X1   g06072(.A(new_n6264_), .B(new_n6262_), .Y(new_n6266_));
  AOI21X1  g06073(.A0(new_n6266_), .A1(new_n6260_), .B0(new_n6265_), .Y(\asquared[63] ));
  AOI21X1  g06074(.A0(new_n6264_), .A1(new_n6262_), .B0(new_n6259_), .Y(new_n6268_));
  OAI21X1  g06075(.A0(new_n6254_), .A1(new_n6252_), .B0(new_n6114_), .Y(new_n6269_));
  INVX1    g06076(.A(new_n6248_), .Y(new_n6270_));
  NOR2X1   g06077(.A(new_n6270_), .B(new_n6158_), .Y(new_n6271_));
  INVX1    g06078(.A(new_n6249_), .Y(new_n6272_));
  AOI21X1  g06079(.A0(new_n6272_), .A1(new_n5978_), .B0(new_n6271_), .Y(new_n6273_));
  AND2X1   g06080(.A(new_n6088_), .B(new_n6082_), .Y(new_n6274_));
  AOI21X1  g06081(.A0(new_n6089_), .A1(new_n6078_), .B0(new_n6274_), .Y(new_n6275_));
  AND2X1   g06082(.A(new_n6072_), .B(new_n6069_), .Y(new_n6276_));
  INVX1    g06083(.A(new_n6075_), .Y(new_n6277_));
  AOI21X1  g06084(.A0(new_n6277_), .A1(new_n6073_), .B0(new_n6276_), .Y(new_n6278_));
  XOR2X1   g06085(.A(new_n6278_), .B(new_n6275_), .Y(new_n6279_));
  INVX1    g06086(.A(new_n6279_), .Y(new_n6280_));
  AND2X1   g06087(.A(new_n6133_), .B(new_n6130_), .Y(new_n6281_));
  AOI21X1  g06088(.A0(new_n6137_), .A1(new_n6134_), .B0(new_n6281_), .Y(new_n6282_));
  XOR2X1   g06089(.A(new_n6282_), .B(new_n6280_), .Y(new_n6283_));
  AND2X1   g06090(.A(new_n5994_), .B(new_n5886_), .Y(new_n6284_));
  AOI21X1  g06091(.A0(new_n6129_), .A1(new_n6118_), .B0(new_n6284_), .Y(new_n6285_));
  NOR2X1   g06092(.A(new_n5916_), .B(new_n5894_), .Y(new_n6286_));
  AOI21X1  g06093(.A0(new_n6081_), .A1(new_n6080_), .B0(new_n6286_), .Y(new_n6287_));
  XOR2X1   g06094(.A(new_n6287_), .B(new_n6285_), .Y(new_n6288_));
  OR2X1    g06095(.A(new_n6085_), .B(new_n6012_), .Y(new_n6289_));
  OAI21X1  g06096(.A0(new_n6087_), .A1(new_n6002_), .B0(new_n6289_), .Y(new_n6290_));
  XOR2X1   g06097(.A(new_n6290_), .B(new_n6288_), .Y(new_n6291_));
  OR2X1    g06098(.A(new_n6245_), .B(new_n6214_), .Y(new_n6292_));
  OAI21X1  g06099(.A0(new_n6247_), .A1(new_n6187_), .B0(new_n6292_), .Y(new_n6293_));
  XOR2X1   g06100(.A(new_n6293_), .B(new_n6291_), .Y(new_n6294_));
  XOR2X1   g06101(.A(new_n6241_), .B(new_n6182_), .Y(new_n6295_));
  XOR2X1   g06102(.A(new_n6295_), .B(new_n6230_), .Y(new_n6296_));
  INVX1    g06103(.A(new_n6193_), .Y(new_n6297_));
  XOR2X1   g06104(.A(new_n6202_), .B(new_n6126_), .Y(new_n6298_));
  XOR2X1   g06105(.A(new_n6298_), .B(new_n6297_), .Y(new_n6299_));
  NOR2X1   g06106(.A(new_n6037_), .B(new_n6027_), .Y(new_n6300_));
  AOI21X1  g06107(.A0(new_n6077_), .A1(new_n5878_), .B0(new_n6300_), .Y(new_n6301_));
  XOR2X1   g06108(.A(new_n6301_), .B(new_n6299_), .Y(new_n6302_));
  XOR2X1   g06109(.A(new_n6302_), .B(new_n6296_), .Y(new_n6303_));
  XOR2X1   g06110(.A(new_n6303_), .B(new_n6294_), .Y(new_n6304_));
  NOR2X1   g06111(.A(new_n6304_), .B(new_n6283_), .Y(new_n6305_));
  AND2X1   g06112(.A(new_n6304_), .B(new_n6283_), .Y(new_n6306_));
  NOR3X1   g06113(.A(new_n6305_), .B(new_n6306_), .C(new_n6273_), .Y(new_n6307_));
  OR2X1    g06114(.A(new_n6307_), .B(new_n6306_), .Y(new_n6308_));
  OAI22X1  g06115(.A0(new_n6308_), .A1(new_n6305_), .B0(new_n6307_), .B1(new_n6273_), .Y(new_n6309_));
  AND2X1   g06116(.A(new_n6154_), .B(new_n6138_), .Y(new_n6310_));
  AND2X1   g06117(.A(new_n6155_), .B(new_n6152_), .Y(new_n6311_));
  NOR3X1   g06118(.A(new_n6311_), .B(new_n6310_), .C(new_n6117_), .Y(new_n6312_));
  NOR2X1   g06119(.A(new_n6250_), .B(new_n6157_), .Y(new_n6313_));
  NOR2X1   g06120(.A(new_n6313_), .B(new_n6312_), .Y(new_n6314_));
  XOR2X1   g06121(.A(new_n6314_), .B(new_n6309_), .Y(new_n6315_));
  NOR2X1   g06122(.A(new_n6107_), .B(new_n6105_), .Y(new_n6316_));
  AOI21X1  g06123(.A0(new_n6108_), .A1(new_n6094_), .B0(new_n6316_), .Y(new_n6317_));
  INVX1    g06124(.A(new_n6317_), .Y(new_n6318_));
  AND2X1   g06125(.A(new_n5931_), .B(new_n5923_), .Y(new_n6319_));
  OAI21X1  g06126(.A0(new_n6319_), .A1(new_n6098_), .B0(new_n6097_), .Y(new_n6320_));
  INVX1    g06127(.A(new_n6104_), .Y(new_n6321_));
  OAI21X1  g06128(.A0(new_n6321_), .A1(new_n6100_), .B0(new_n6320_), .Y(new_n6322_));
  INVX1    g06129(.A(new_n6211_), .Y(new_n6323_));
  XOR2X1   g06130(.A(new_n6323_), .B(new_n6171_), .Y(new_n6324_));
  XOR2X1   g06131(.A(new_n6324_), .B(new_n6164_), .Y(new_n6325_));
  AND2X1   g06132(.A(new_n6173_), .B(new_n6167_), .Y(new_n6326_));
  AOI21X1  g06133(.A0(new_n6185_), .A1(new_n6174_), .B0(new_n6326_), .Y(new_n6327_));
  XOR2X1   g06134(.A(new_n6327_), .B(new_n6325_), .Y(new_n6328_));
  AND2X1   g06135(.A(new_n6232_), .B(new_n6224_), .Y(new_n6329_));
  AND2X1   g06136(.A(new_n6243_), .B(new_n6233_), .Y(new_n6330_));
  OR2X1    g06137(.A(new_n6330_), .B(new_n6329_), .Y(new_n6331_));
  XOR2X1   g06138(.A(new_n6331_), .B(new_n6328_), .Y(new_n6332_));
  OR2X1    g06139(.A(new_n6142_), .B(new_n6140_), .Y(new_n6333_));
  OAI21X1  g06140(.A0(new_n6146_), .A1(new_n6144_), .B0(new_n6333_), .Y(new_n6334_));
  OR2X1    g06141(.A(new_n6203_), .B(new_n6196_), .Y(new_n6335_));
  INVX1    g06142(.A(new_n6204_), .Y(new_n6336_));
  OAI21X1  g06143(.A0(new_n6213_), .A1(new_n6336_), .B0(new_n6335_), .Y(new_n6337_));
  XOR2X1   g06144(.A(new_n6337_), .B(new_n6334_), .Y(new_n6338_));
  NAND4X1  g06145(.A(\a[61] ), .B(\a[32] ), .C(\a[30] ), .D(\a[1] ), .Y(new_n6339_));
  AND2X1   g06146(.A(\a[63] ), .B(\a[0] ), .Y(new_n6340_));
  XOR2X1   g06147(.A(new_n6340_), .B(new_n6339_), .Y(new_n6341_));
  AOI21X1  g06148(.A0(\a[62] ), .A1(\a[1] ), .B0(new_n2219_), .Y(new_n6342_));
  AOI21X1  g06149(.A0(\a[62] ), .A1(\a[32] ), .B0(new_n202_), .Y(new_n6343_));
  AOI21X1  g06150(.A0(new_n6343_), .A1(\a[62] ), .B0(new_n6342_), .Y(new_n6344_));
  XOR2X1   g06151(.A(new_n6344_), .B(new_n6341_), .Y(new_n6345_));
  NAND4X1  g06152(.A(\a[39] ), .B(\a[37] ), .C(\a[26] ), .D(\a[24] ), .Y(new_n6346_));
  NAND4X1  g06153(.A(\a[39] ), .B(\a[38] ), .C(\a[25] ), .D(\a[24] ), .Y(new_n6347_));
  AOI22X1  g06154(.A0(new_n6347_), .A1(new_n6346_), .B0(new_n3164_), .B1(new_n1770_), .Y(new_n6348_));
  NAND4X1  g06155(.A(\a[38] ), .B(\a[37] ), .C(\a[26] ), .D(\a[25] ), .Y(new_n6349_));
  NAND3X1  g06156(.A(new_n6347_), .B(new_n6346_), .C(new_n6349_), .Y(new_n6350_));
  AOI22X1  g06157(.A0(\a[38] ), .A1(\a[25] ), .B0(\a[37] ), .B1(\a[26] ), .Y(new_n6351_));
  NAND2X1  g06158(.A(\a[39] ), .B(\a[24] ), .Y(new_n6352_));
  OAI22X1  g06159(.A0(new_n6352_), .A1(new_n6348_), .B0(new_n6351_), .B1(new_n6350_), .Y(new_n6353_));
  AOI22X1  g06160(.A0(new_n4695_), .A1(new_n1484_), .B0(new_n2682_), .B1(new_n1671_), .Y(new_n6354_));
  AOI21X1  g06161(.A0(new_n2361_), .A1(new_n1674_), .B0(new_n6354_), .Y(new_n6355_));
  NAND2X1  g06162(.A(\a[36] ), .B(\a[27] ), .Y(new_n6356_));
  AOI22X1  g06163(.A0(\a[35] ), .A1(\a[28] ), .B0(\a[34] ), .B1(\a[29] ), .Y(new_n6357_));
  AOI21X1  g06164(.A0(new_n2361_), .A1(new_n1674_), .B0(new_n6355_), .Y(new_n6358_));
  INVX1    g06165(.A(new_n6358_), .Y(new_n6359_));
  OAI22X1  g06166(.A0(new_n6359_), .A1(new_n6357_), .B0(new_n6356_), .B1(new_n6355_), .Y(new_n6360_));
  XOR2X1   g06167(.A(new_n6360_), .B(new_n6353_), .Y(new_n6361_));
  XOR2X1   g06168(.A(new_n6361_), .B(new_n6345_), .Y(new_n6362_));
  XOR2X1   g06169(.A(new_n6362_), .B(new_n6338_), .Y(new_n6363_));
  XOR2X1   g06170(.A(new_n6363_), .B(new_n6332_), .Y(new_n6364_));
  XOR2X1   g06171(.A(new_n6364_), .B(new_n6322_), .Y(new_n6365_));
  XOR2X1   g06172(.A(new_n6365_), .B(new_n6318_), .Y(new_n6366_));
  NOR2X1   g06173(.A(new_n6090_), .B(new_n6076_), .Y(new_n6367_));
  AOI21X1  g06174(.A0(new_n6093_), .A1(new_n6091_), .B0(new_n6367_), .Y(new_n6368_));
  NOR2X1   g06175(.A(new_n6151_), .B(new_n6153_), .Y(new_n6369_));
  OR2X1    g06176(.A(new_n6310_), .B(new_n6369_), .Y(new_n6370_));
  AND2X1   g06177(.A(\a[54] ), .B(\a[46] ), .Y(new_n6371_));
  NAND4X1  g06178(.A(\a[54] ), .B(\a[45] ), .C(\a[18] ), .D(\a[9] ), .Y(new_n6372_));
  NAND4X1  g06179(.A(\a[46] ), .B(\a[45] ), .C(\a[18] ), .D(\a[17] ), .Y(new_n6373_));
  AOI22X1  g06180(.A0(new_n6373_), .A1(new_n6372_), .B0(new_n6371_), .B1(new_n1226_), .Y(new_n6374_));
  NAND4X1  g06181(.A(\a[54] ), .B(\a[46] ), .C(\a[17] ), .D(\a[9] ), .Y(new_n6375_));
  NAND3X1  g06182(.A(new_n6373_), .B(new_n6372_), .C(new_n6375_), .Y(new_n6376_));
  AOI22X1  g06183(.A0(\a[54] ), .A1(\a[9] ), .B0(\a[46] ), .B1(\a[17] ), .Y(new_n6377_));
  NAND2X1  g06184(.A(\a[45] ), .B(\a[18] ), .Y(new_n6378_));
  OAI22X1  g06185(.A0(new_n6378_), .A1(new_n6374_), .B0(new_n6377_), .B1(new_n6376_), .Y(new_n6379_));
  NOR4X1   g06186(.A(new_n4354_), .B(new_n4041_), .C(new_n571_), .D(new_n488_), .Y(new_n6380_));
  NOR4X1   g06187(.A(new_n5245_), .B(new_n4041_), .C(new_n571_), .D(new_n570_), .Y(new_n6381_));
  AOI21X1  g06188(.A0(new_n5048_), .A1(new_n1002_), .B0(new_n6381_), .Y(new_n6382_));
  NOR2X1   g06189(.A(new_n6382_), .B(new_n6380_), .Y(new_n6383_));
  NAND2X1  g06190(.A(\a[53] ), .B(\a[10] ), .Y(new_n6384_));
  AOI22X1  g06191(.A0(\a[52] ), .A1(\a[11] ), .B0(\a[47] ), .B1(\a[16] ), .Y(new_n6385_));
  NOR2X1   g06192(.A(new_n6383_), .B(new_n6380_), .Y(new_n6386_));
  INVX1    g06193(.A(new_n6386_), .Y(new_n6387_));
  OAI22X1  g06194(.A0(new_n6387_), .A1(new_n6385_), .B0(new_n6384_), .B1(new_n6383_), .Y(new_n6388_));
  XOR2X1   g06195(.A(new_n6388_), .B(new_n6379_), .Y(new_n6389_));
  AND2X1   g06196(.A(\a[48] ), .B(\a[15] ), .Y(new_n6390_));
  INVX1    g06197(.A(new_n6390_), .Y(new_n6391_));
  NAND4X1  g06198(.A(\a[50] ), .B(\a[48] ), .C(\a[15] ), .D(\a[13] ), .Y(new_n6392_));
  NAND4X1  g06199(.A(\a[51] ), .B(\a[48] ), .C(\a[15] ), .D(\a[12] ), .Y(new_n6393_));
  AOI22X1  g06200(.A0(new_n6393_), .A1(new_n6392_), .B0(new_n4484_), .B1(new_n586_), .Y(new_n6394_));
  AOI21X1  g06201(.A0(new_n4484_), .A1(new_n586_), .B0(new_n6394_), .Y(new_n6395_));
  INVX1    g06202(.A(new_n6395_), .Y(new_n6396_));
  AOI22X1  g06203(.A0(\a[51] ), .A1(\a[12] ), .B0(\a[50] ), .B1(\a[13] ), .Y(new_n6397_));
  OAI22X1  g06204(.A0(new_n6397_), .A1(new_n6396_), .B0(new_n6394_), .B1(new_n6391_), .Y(new_n6398_));
  INVX1    g06205(.A(new_n6398_), .Y(new_n6399_));
  XOR2X1   g06206(.A(new_n6399_), .B(new_n6389_), .Y(new_n6400_));
  AOI22X1  g06207(.A0(\a[57] ), .A1(\a[6] ), .B0(\a[43] ), .B1(\a[20] ), .Y(new_n6401_));
  AND2X1   g06208(.A(\a[40] ), .B(\a[23] ), .Y(new_n6402_));
  INVX1    g06209(.A(new_n6402_), .Y(new_n6403_));
  NOR4X1   g06210(.A(new_n5441_), .B(new_n3037_), .C(new_n934_), .D(new_n230_), .Y(new_n6404_));
  NOR3X1   g06211(.A(new_n6403_), .B(new_n6404_), .C(new_n6401_), .Y(new_n6405_));
  NOR2X1   g06212(.A(new_n6405_), .B(new_n6404_), .Y(new_n6406_));
  INVX1    g06213(.A(new_n6406_), .Y(new_n6407_));
  OAI22X1  g06214(.A0(new_n6407_), .A1(new_n6401_), .B0(new_n6405_), .B1(new_n6403_), .Y(new_n6408_));
  AND2X1   g06215(.A(\a[49] ), .B(\a[14] ), .Y(new_n6409_));
  AOI22X1  g06216(.A0(\a[33] ), .A1(\a[30] ), .B0(\a[32] ), .B1(\a[31] ), .Y(new_n6410_));
  INVX1    g06217(.A(new_n6410_), .Y(new_n6411_));
  NOR4X1   g06218(.A(new_n1851_), .B(new_n2219_), .C(new_n1704_), .D(new_n1684_), .Y(new_n6412_));
  OR4X1    g06219(.A(new_n6410_), .B(new_n6412_), .C(new_n3915_), .D(new_n490_), .Y(new_n6413_));
  AOI21X1  g06220(.A0(new_n6411_), .A1(new_n6409_), .B0(new_n6412_), .Y(new_n6414_));
  AOI22X1  g06221(.A0(new_n6414_), .A1(new_n6411_), .B0(new_n6413_), .B1(new_n6409_), .Y(new_n6415_));
  XOR2X1   g06222(.A(new_n6415_), .B(new_n6408_), .Y(new_n6416_));
  NOR4X1   g06223(.A(new_n4906_), .B(new_n5268_), .C(new_n752_), .D(new_n413_), .Y(new_n6417_));
  NAND4X1  g06224(.A(\a[56] ), .B(\a[55] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n6418_));
  NAND4X1  g06225(.A(\a[56] ), .B(\a[44] ), .C(\a[19] ), .D(\a[7] ), .Y(new_n6419_));
  AOI21X1  g06226(.A0(new_n6419_), .A1(new_n6418_), .B0(new_n6417_), .Y(new_n6420_));
  NOR3X1   g06227(.A(new_n6420_), .B(new_n6022_), .C(new_n532_), .Y(new_n6421_));
  OAI22X1  g06228(.A0(new_n4906_), .A1(new_n413_), .B0(new_n5268_), .B1(new_n752_), .Y(new_n6422_));
  NOR2X1   g06229(.A(new_n6420_), .B(new_n6417_), .Y(new_n6423_));
  AOI21X1  g06230(.A0(new_n6423_), .A1(new_n6422_), .B0(new_n6421_), .Y(new_n6424_));
  XOR2X1   g06231(.A(new_n6424_), .B(new_n6416_), .Y(new_n6425_));
  INVX1    g06232(.A(new_n6425_), .Y(new_n6426_));
  AND2X1   g06233(.A(\a[60] ), .B(\a[59] ), .Y(new_n6427_));
  AND2X1   g06234(.A(\a[61] ), .B(\a[60] ), .Y(new_n6428_));
  AOI22X1  g06235(.A0(new_n6428_), .A1(new_n231_), .B0(new_n6020_), .B1(new_n235_), .Y(new_n6429_));
  AOI21X1  g06236(.A0(new_n6427_), .A1(new_n294_), .B0(new_n6429_), .Y(new_n6430_));
  AND2X1   g06237(.A(\a[61] ), .B(\a[2] ), .Y(new_n6431_));
  INVX1    g06238(.A(new_n6431_), .Y(new_n6432_));
  AOI21X1  g06239(.A0(new_n6427_), .A1(new_n294_), .B0(new_n6430_), .Y(new_n6433_));
  INVX1    g06240(.A(new_n6433_), .Y(new_n6434_));
  AOI22X1  g06241(.A0(\a[60] ), .A1(\a[3] ), .B0(\a[59] ), .B1(\a[4] ), .Y(new_n6435_));
  OAI22X1  g06242(.A0(new_n6435_), .A1(new_n6434_), .B0(new_n6432_), .B1(new_n6430_), .Y(new_n6436_));
  XOR2X1   g06243(.A(new_n6436_), .B(new_n6220_), .Y(new_n6437_));
  AOI22X1  g06244(.A0(\a[42] ), .A1(\a[21] ), .B0(\a[41] ), .B1(\a[22] ), .Y(new_n6438_));
  AND2X1   g06245(.A(\a[58] ), .B(\a[5] ), .Y(new_n6439_));
  AND2X1   g06246(.A(new_n3607_), .B(new_n1154_), .Y(new_n6440_));
  OAI21X1  g06247(.A0(new_n6438_), .A1(new_n6440_), .B0(new_n6439_), .Y(new_n6441_));
  INVX1    g06248(.A(new_n6438_), .Y(new_n6442_));
  AOI21X1  g06249(.A0(new_n6442_), .A1(new_n6439_), .B0(new_n6440_), .Y(new_n6443_));
  INVX1    g06250(.A(new_n6443_), .Y(new_n6444_));
  OAI21X1  g06251(.A0(new_n6444_), .A1(new_n6438_), .B0(new_n6441_), .Y(new_n6445_));
  INVX1    g06252(.A(new_n6445_), .Y(new_n6446_));
  XOR2X1   g06253(.A(new_n6446_), .B(new_n6437_), .Y(new_n6447_));
  XOR2X1   g06254(.A(new_n6447_), .B(new_n6426_), .Y(new_n6448_));
  XOR2X1   g06255(.A(new_n6448_), .B(new_n6400_), .Y(new_n6449_));
  XOR2X1   g06256(.A(new_n6449_), .B(new_n6370_), .Y(new_n6450_));
  XOR2X1   g06257(.A(new_n6450_), .B(new_n6368_), .Y(new_n6451_));
  XOR2X1   g06258(.A(new_n6451_), .B(new_n6366_), .Y(new_n6452_));
  XOR2X1   g06259(.A(new_n6452_), .B(new_n6315_), .Y(new_n6453_));
  NOR2X1   g06260(.A(new_n6453_), .B(new_n6269_), .Y(new_n6454_));
  AND2X1   g06261(.A(new_n6453_), .B(new_n6269_), .Y(new_n6455_));
  OR2X1    g06262(.A(new_n6455_), .B(new_n6454_), .Y(new_n6456_));
  XOR2X1   g06263(.A(new_n6456_), .B(new_n6268_), .Y(\asquared[64] ));
  AND2X1   g06264(.A(new_n6365_), .B(new_n6318_), .Y(new_n6458_));
  INVX1    g06265(.A(new_n6458_), .Y(new_n6459_));
  INVX1    g06266(.A(new_n6366_), .Y(new_n6460_));
  OAI21X1  g06267(.A0(new_n6451_), .A1(new_n6460_), .B0(new_n6459_), .Y(new_n6461_));
  OAI21X1  g06268(.A0(new_n6310_), .A1(new_n6369_), .B0(new_n6449_), .Y(new_n6462_));
  INVX1    g06269(.A(new_n6450_), .Y(new_n6463_));
  OAI21X1  g06270(.A0(new_n6463_), .A1(new_n6368_), .B0(new_n6462_), .Y(new_n6464_));
  AND2X1   g06271(.A(new_n6363_), .B(new_n6332_), .Y(new_n6465_));
  AOI21X1  g06272(.A0(new_n6364_), .A1(new_n6322_), .B0(new_n6465_), .Y(new_n6466_));
  NAND2X1  g06273(.A(new_n6447_), .B(new_n6425_), .Y(new_n6467_));
  OAI21X1  g06274(.A0(new_n6448_), .A1(new_n6400_), .B0(new_n6467_), .Y(new_n6468_));
  AND2X1   g06275(.A(new_n6337_), .B(new_n6334_), .Y(new_n6469_));
  AOI21X1  g06276(.A0(new_n6362_), .A1(new_n6338_), .B0(new_n6469_), .Y(new_n6470_));
  XOR2X1   g06277(.A(new_n6470_), .B(new_n6468_), .Y(new_n6471_));
  AND2X1   g06278(.A(new_n6360_), .B(new_n6353_), .Y(new_n6472_));
  AOI21X1  g06279(.A0(new_n6361_), .A1(new_n6345_), .B0(new_n6472_), .Y(new_n6473_));
  XOR2X1   g06280(.A(new_n6407_), .B(new_n6376_), .Y(new_n6474_));
  XOR2X1   g06281(.A(new_n6474_), .B(new_n6358_), .Y(new_n6475_));
  INVX1    g06282(.A(new_n6423_), .Y(new_n6476_));
  XOR2X1   g06283(.A(new_n6443_), .B(new_n6433_), .Y(new_n6477_));
  XOR2X1   g06284(.A(new_n6477_), .B(new_n6476_), .Y(new_n6478_));
  INVX1    g06285(.A(new_n6478_), .Y(new_n6479_));
  XOR2X1   g06286(.A(new_n6479_), .B(new_n6475_), .Y(new_n6480_));
  INVX1    g06287(.A(new_n6480_), .Y(new_n6481_));
  XOR2X1   g06288(.A(new_n6481_), .B(new_n6473_), .Y(new_n6482_));
  INVX1    g06289(.A(new_n6482_), .Y(new_n6483_));
  XOR2X1   g06290(.A(new_n6483_), .B(new_n6471_), .Y(new_n6484_));
  XOR2X1   g06291(.A(new_n6484_), .B(new_n6466_), .Y(new_n6485_));
  XOR2X1   g06292(.A(new_n6485_), .B(new_n6464_), .Y(new_n6486_));
  XOR2X1   g06293(.A(new_n6486_), .B(new_n6461_), .Y(new_n6487_));
  AND2X1   g06294(.A(new_n6293_), .B(new_n6291_), .Y(new_n6488_));
  AOI21X1  g06295(.A0(new_n6303_), .A1(new_n6294_), .B0(new_n6488_), .Y(new_n6489_));
  AOI22X1  g06296(.A0(\a[57] ), .A1(\a[7] ), .B0(\a[47] ), .B1(\a[17] ), .Y(new_n6490_));
  NOR4X1   g06297(.A(new_n5441_), .B(new_n4041_), .C(new_n616_), .D(new_n532_), .Y(new_n6491_));
  NAND4X1  g06298(.A(\a[58] ), .B(\a[47] ), .C(\a[17] ), .D(\a[6] ), .Y(new_n6492_));
  NAND4X1  g06299(.A(\a[58] ), .B(\a[57] ), .C(\a[7] ), .D(\a[6] ), .Y(new_n6493_));
  AOI21X1  g06300(.A0(new_n6493_), .A1(new_n6492_), .B0(new_n6491_), .Y(new_n6494_));
  NOR2X1   g06301(.A(new_n6494_), .B(new_n6491_), .Y(new_n6495_));
  INVX1    g06302(.A(new_n6495_), .Y(new_n6496_));
  NAND2X1  g06303(.A(\a[58] ), .B(\a[6] ), .Y(new_n6497_));
  OAI22X1  g06304(.A0(new_n6497_), .A1(new_n6494_), .B0(new_n6496_), .B1(new_n6490_), .Y(new_n6498_));
  AOI22X1  g06305(.A0(new_n4992_), .A1(new_n1236_), .B0(new_n3208_), .B1(new_n2134_), .Y(new_n6499_));
  AOI21X1  g06306(.A0(new_n3462_), .A1(new_n1154_), .B0(new_n6499_), .Y(new_n6500_));
  NAND2X1  g06307(.A(\a[44] ), .B(\a[20] ), .Y(new_n6501_));
  INVX1    g06308(.A(new_n3462_), .Y(new_n6502_));
  OAI21X1  g06309(.A0(new_n6502_), .A1(new_n1397_), .B0(new_n6499_), .Y(new_n6503_));
  AOI22X1  g06310(.A0(\a[43] ), .A1(\a[21] ), .B0(\a[42] ), .B1(\a[22] ), .Y(new_n6504_));
  OAI22X1  g06311(.A0(new_n6504_), .A1(new_n6503_), .B0(new_n6501_), .B1(new_n6500_), .Y(new_n6505_));
  XOR2X1   g06312(.A(new_n6505_), .B(new_n6498_), .Y(new_n6506_));
  AOI22X1  g06313(.A0(new_n4404_), .A1(new_n1219_), .B0(new_n2847_), .B1(new_n1134_), .Y(new_n6507_));
  AOI21X1  g06314(.A0(new_n4077_), .A1(new_n1532_), .B0(new_n6507_), .Y(new_n6508_));
  AND2X1   g06315(.A(\a[41] ), .B(\a[23] ), .Y(new_n6509_));
  INVX1    g06316(.A(new_n6509_), .Y(new_n6510_));
  AOI21X1  g06317(.A0(new_n4077_), .A1(new_n1532_), .B0(new_n6508_), .Y(new_n6511_));
  INVX1    g06318(.A(new_n6511_), .Y(new_n6512_));
  AOI22X1  g06319(.A0(\a[40] ), .A1(\a[24] ), .B0(\a[39] ), .B1(\a[25] ), .Y(new_n6513_));
  OAI22X1  g06320(.A0(new_n6513_), .A1(new_n6512_), .B0(new_n6510_), .B1(new_n6508_), .Y(new_n6514_));
  XOR2X1   g06321(.A(new_n6514_), .B(new_n6506_), .Y(new_n6515_));
  AOI22X1  g06322(.A0(\a[56] ), .A1(\a[8] ), .B0(\a[48] ), .B1(\a[16] ), .Y(new_n6516_));
  AND2X1   g06323(.A(\a[38] ), .B(\a[26] ), .Y(new_n6517_));
  INVX1    g06324(.A(new_n6517_), .Y(new_n6518_));
  NOR4X1   g06325(.A(new_n6022_), .B(new_n3926_), .C(new_n571_), .D(new_n413_), .Y(new_n6519_));
  NOR3X1   g06326(.A(new_n6518_), .B(new_n6519_), .C(new_n6516_), .Y(new_n6520_));
  NOR2X1   g06327(.A(new_n6520_), .B(new_n6519_), .Y(new_n6521_));
  INVX1    g06328(.A(new_n6521_), .Y(new_n6522_));
  OAI22X1  g06329(.A0(new_n6522_), .A1(new_n6516_), .B0(new_n6520_), .B1(new_n6518_), .Y(new_n6523_));
  AND2X1   g06330(.A(\a[37] ), .B(\a[27] ), .Y(new_n6524_));
  INVX1    g06331(.A(new_n3330_), .Y(new_n6525_));
  AND2X1   g06332(.A(\a[37] ), .B(\a[35] ), .Y(new_n6526_));
  INVX1    g06333(.A(new_n6526_), .Y(new_n6527_));
  OAI22X1  g06334(.A0(new_n6527_), .A1(new_n1673_), .B0(new_n6525_), .B1(new_n1672_), .Y(new_n6528_));
  OAI21X1  g06335(.A0(new_n5417_), .A1(new_n1675_), .B0(new_n6528_), .Y(new_n6529_));
  AOI21X1  g06336(.A0(new_n2682_), .A1(new_n1674_), .B0(new_n6528_), .Y(new_n6530_));
  OAI22X1  g06337(.A0(new_n2583_), .A1(new_n1431_), .B0(new_n2557_), .B1(new_n1803_), .Y(new_n6531_));
  AOI22X1  g06338(.A0(new_n6531_), .A1(new_n6530_), .B0(new_n6529_), .B1(new_n6524_), .Y(new_n6532_));
  XOR2X1   g06339(.A(new_n6532_), .B(new_n6523_), .Y(new_n6533_));
  AND2X1   g06340(.A(\a[50] ), .B(\a[14] ), .Y(new_n6534_));
  AOI22X1  g06341(.A0(\a[34] ), .A1(\a[30] ), .B0(\a[33] ), .B1(\a[31] ), .Y(new_n6535_));
  INVX1    g06342(.A(new_n6535_), .Y(new_n6536_));
  NAND4X1  g06343(.A(\a[34] ), .B(\a[33] ), .C(\a[31] ), .D(\a[30] ), .Y(new_n6537_));
  NAND3X1  g06344(.A(new_n6536_), .B(new_n6537_), .C(new_n6534_), .Y(new_n6538_));
  AOI22X1  g06345(.A0(new_n6536_), .A1(new_n6534_), .B0(new_n2918_), .B1(new_n2075_), .Y(new_n6539_));
  AOI22X1  g06346(.A0(new_n6539_), .A1(new_n6536_), .B0(new_n6538_), .B1(new_n6534_), .Y(new_n6540_));
  XOR2X1   g06347(.A(new_n6540_), .B(new_n6533_), .Y(new_n6541_));
  AOI22X1  g06348(.A0(\a[46] ), .A1(\a[18] ), .B0(\a[45] ), .B1(\a[19] ), .Y(new_n6542_));
  AND2X1   g06349(.A(new_n3809_), .B(new_n855_), .Y(new_n6543_));
  OAI21X1  g06350(.A0(new_n6543_), .A1(new_n6542_), .B0(new_n6019_), .Y(new_n6544_));
  INVX1    g06351(.A(new_n6542_), .Y(new_n6545_));
  AOI21X1  g06352(.A0(new_n6545_), .A1(new_n6019_), .B0(new_n6543_), .Y(new_n6546_));
  INVX1    g06353(.A(new_n6546_), .Y(new_n6547_));
  OAI21X1  g06354(.A0(new_n6547_), .A1(new_n6542_), .B0(new_n6544_), .Y(new_n6548_));
  INVX1    g06355(.A(\a[63] ), .Y(new_n6549_));
  NOR3X1   g06356(.A(new_n6339_), .B(new_n6549_), .C(new_n194_), .Y(new_n6550_));
  NOR2X1   g06357(.A(new_n6344_), .B(new_n6341_), .Y(new_n6551_));
  NOR2X1   g06358(.A(new_n6551_), .B(new_n6550_), .Y(new_n6552_));
  XOR2X1   g06359(.A(new_n6552_), .B(new_n6548_), .Y(new_n6553_));
  INVX1    g06360(.A(new_n6428_), .Y(new_n6554_));
  INVX1    g06361(.A(new_n6191_), .Y(new_n6555_));
  AND2X1   g06362(.A(\a[62] ), .B(\a[61] ), .Y(new_n6556_));
  INVX1    g06363(.A(new_n6556_), .Y(new_n6557_));
  OAI22X1  g06364(.A0(new_n6557_), .A1(new_n249_), .B0(new_n6555_), .B1(new_n584_), .Y(new_n6558_));
  OAI21X1  g06365(.A0(new_n6554_), .A1(new_n217_), .B0(new_n6558_), .Y(new_n6559_));
  AND2X1   g06366(.A(\a[62] ), .B(\a[2] ), .Y(new_n6560_));
  AOI21X1  g06367(.A0(new_n6428_), .A1(new_n294_), .B0(new_n6558_), .Y(new_n6561_));
  OAI22X1  g06368(.A0(new_n6023_), .A1(new_n223_), .B0(new_n5952_), .B1(new_n340_), .Y(new_n6562_));
  AOI22X1  g06369(.A0(new_n6562_), .A1(new_n6561_), .B0(new_n6560_), .B1(new_n6559_), .Y(new_n6563_));
  XOR2X1   g06370(.A(new_n6563_), .B(new_n6553_), .Y(new_n6564_));
  INVX1    g06371(.A(new_n6564_), .Y(new_n6565_));
  XOR2X1   g06372(.A(new_n6565_), .B(new_n6541_), .Y(new_n6566_));
  XOR2X1   g06373(.A(new_n6566_), .B(new_n6515_), .Y(new_n6567_));
  XOR2X1   g06374(.A(new_n6567_), .B(new_n6489_), .Y(new_n6568_));
  NOR2X1   g06375(.A(new_n6241_), .B(new_n6182_), .Y(new_n6569_));
  AOI21X1  g06376(.A0(new_n6295_), .A1(new_n6231_), .B0(new_n6569_), .Y(new_n6570_));
  AND2X1   g06377(.A(new_n6323_), .B(new_n6171_), .Y(new_n6571_));
  AOI21X1  g06378(.A0(new_n6324_), .A1(new_n6165_), .B0(new_n6571_), .Y(new_n6572_));
  XOR2X1   g06379(.A(new_n6572_), .B(new_n6570_), .Y(new_n6573_));
  AOI21X1  g06380(.A0(new_n6122_), .A1(new_n6125_), .B0(new_n6202_), .Y(new_n6574_));
  AOI21X1  g06381(.A0(new_n6298_), .A1(new_n6297_), .B0(new_n6574_), .Y(new_n6575_));
  XOR2X1   g06382(.A(new_n6575_), .B(new_n6573_), .Y(new_n6576_));
  NOR2X1   g06383(.A(new_n6327_), .B(new_n6325_), .Y(new_n6577_));
  AOI21X1  g06384(.A0(new_n6331_), .A1(new_n6328_), .B0(new_n6577_), .Y(new_n6578_));
  INVX1    g06385(.A(new_n6299_), .Y(new_n6579_));
  NOR2X1   g06386(.A(new_n6301_), .B(new_n6579_), .Y(new_n6580_));
  NOR2X1   g06387(.A(new_n6302_), .B(new_n6296_), .Y(new_n6581_));
  NOR2X1   g06388(.A(new_n6581_), .B(new_n6580_), .Y(new_n6582_));
  INVX1    g06389(.A(new_n6582_), .Y(new_n6583_));
  XOR2X1   g06390(.A(new_n6583_), .B(new_n6578_), .Y(new_n6584_));
  XOR2X1   g06391(.A(new_n6584_), .B(new_n6576_), .Y(new_n6585_));
  XOR2X1   g06392(.A(new_n6585_), .B(new_n6568_), .Y(new_n6586_));
  XOR2X1   g06393(.A(new_n6396_), .B(new_n6350_), .Y(new_n6587_));
  XOR2X1   g06394(.A(new_n6587_), .B(new_n6387_), .Y(new_n6588_));
  INVX1    g06395(.A(new_n6408_), .Y(new_n6589_));
  OR2X1    g06396(.A(new_n6424_), .B(new_n6416_), .Y(new_n6590_));
  OAI21X1  g06397(.A0(new_n6415_), .A1(new_n6589_), .B0(new_n6590_), .Y(new_n6591_));
  XOR2X1   g06398(.A(new_n6591_), .B(new_n6588_), .Y(new_n6592_));
  AND2X1   g06399(.A(new_n6388_), .B(new_n6379_), .Y(new_n6593_));
  AND2X1   g06400(.A(new_n6398_), .B(new_n6389_), .Y(new_n6594_));
  OR2X1    g06401(.A(new_n6594_), .B(new_n6593_), .Y(new_n6595_));
  XOR2X1   g06402(.A(new_n6595_), .B(new_n6592_), .Y(new_n6596_));
  INVX1    g06403(.A(new_n6596_), .Y(new_n6597_));
  OR2X1    g06404(.A(new_n6278_), .B(new_n6275_), .Y(new_n6598_));
  OAI21X1  g06405(.A0(new_n6282_), .A1(new_n6280_), .B0(new_n6598_), .Y(new_n6599_));
  XOR2X1   g06406(.A(new_n6599_), .B(new_n6597_), .Y(new_n6600_));
  NOR2X1   g06407(.A(new_n6287_), .B(new_n6285_), .Y(new_n6601_));
  AOI21X1  g06408(.A0(new_n6290_), .A1(new_n6288_), .B0(new_n6601_), .Y(new_n6602_));
  NOR2X1   g06409(.A(new_n6446_), .B(new_n6437_), .Y(new_n6603_));
  AOI21X1  g06410(.A0(new_n6436_), .A1(new_n6221_), .B0(new_n6603_), .Y(new_n6604_));
  XOR2X1   g06411(.A(new_n6604_), .B(new_n6602_), .Y(new_n6605_));
  INVX1    g06412(.A(\a[62] ), .Y(new_n6606_));
  NOR4X1   g06413(.A(\a[63] ), .B(new_n6606_), .C(new_n2219_), .D(new_n202_), .Y(new_n6607_));
  AOI21X1  g06414(.A0(new_n6343_), .A1(\a[63] ), .B0(new_n6607_), .Y(new_n6608_));
  XOR2X1   g06415(.A(new_n6608_), .B(new_n6414_), .Y(new_n6609_));
  NOR4X1   g06416(.A(new_n4835_), .B(new_n3915_), .C(new_n549_), .D(new_n570_), .Y(new_n6610_));
  NAND4X1  g06417(.A(\a[55] ), .B(\a[49] ), .C(\a[15] ), .D(\a[9] ), .Y(new_n6611_));
  NAND4X1  g06418(.A(\a[55] ), .B(\a[54] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n6612_));
  AOI21X1  g06419(.A0(new_n6612_), .A1(new_n6611_), .B0(new_n6610_), .Y(new_n6613_));
  OR2X1    g06420(.A(new_n6613_), .B(new_n6610_), .Y(new_n6614_));
  AOI22X1  g06421(.A0(\a[54] ), .A1(\a[10] ), .B0(\a[49] ), .B1(\a[15] ), .Y(new_n6615_));
  NAND2X1  g06422(.A(\a[55] ), .B(\a[9] ), .Y(new_n6616_));
  OAI22X1  g06423(.A0(new_n6616_), .A1(new_n6613_), .B0(new_n6615_), .B1(new_n6614_), .Y(new_n6617_));
  NAND4X1  g06424(.A(\a[53] ), .B(\a[51] ), .C(\a[13] ), .D(\a[11] ), .Y(new_n6618_));
  NAND4X1  g06425(.A(\a[52] ), .B(\a[51] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n6619_));
  AOI22X1  g06426(.A0(new_n6619_), .A1(new_n6618_), .B0(new_n5048_), .B1(new_n482_), .Y(new_n6620_));
  NAND2X1  g06427(.A(\a[51] ), .B(\a[13] ), .Y(new_n6621_));
  AOI22X1  g06428(.A0(\a[53] ), .A1(\a[11] ), .B0(\a[52] ), .B1(\a[12] ), .Y(new_n6622_));
  AOI21X1  g06429(.A0(new_n5048_), .A1(new_n482_), .B0(new_n6620_), .Y(new_n6623_));
  INVX1    g06430(.A(new_n6623_), .Y(new_n6624_));
  OAI22X1  g06431(.A0(new_n6624_), .A1(new_n6622_), .B0(new_n6621_), .B1(new_n6620_), .Y(new_n6625_));
  XOR2X1   g06432(.A(new_n6625_), .B(new_n6617_), .Y(new_n6626_));
  XOR2X1   g06433(.A(new_n6626_), .B(new_n6609_), .Y(new_n6627_));
  INVX1    g06434(.A(new_n6627_), .Y(new_n6628_));
  XOR2X1   g06435(.A(new_n6628_), .B(new_n6605_), .Y(new_n6629_));
  XOR2X1   g06436(.A(new_n6629_), .B(new_n6600_), .Y(new_n6630_));
  XOR2X1   g06437(.A(new_n6630_), .B(new_n6308_), .Y(new_n6631_));
  XOR2X1   g06438(.A(new_n6631_), .B(new_n6586_), .Y(new_n6632_));
  XOR2X1   g06439(.A(new_n6632_), .B(new_n6487_), .Y(new_n6633_));
  OAI21X1  g06440(.A0(new_n6313_), .A1(new_n6312_), .B0(new_n6309_), .Y(new_n6634_));
  OR2X1    g06441(.A(new_n6452_), .B(new_n6315_), .Y(new_n6635_));
  AND2X1   g06442(.A(new_n6635_), .B(new_n6634_), .Y(new_n6636_));
  NOR2X1   g06443(.A(new_n6636_), .B(new_n6633_), .Y(new_n6637_));
  INVX1    g06444(.A(new_n6637_), .Y(new_n6638_));
  NAND2X1  g06445(.A(new_n6453_), .B(new_n6269_), .Y(new_n6639_));
  OAI21X1  g06446(.A0(new_n6454_), .A1(new_n6268_), .B0(new_n6639_), .Y(new_n6640_));
  AND2X1   g06447(.A(new_n6636_), .B(new_n6633_), .Y(new_n6641_));
  INVX1    g06448(.A(new_n6641_), .Y(new_n6642_));
  AOI21X1  g06449(.A0(new_n6638_), .A1(new_n6642_), .B0(new_n6640_), .Y(new_n6643_));
  AND2X1   g06450(.A(new_n6642_), .B(new_n6640_), .Y(new_n6644_));
  AOI21X1  g06451(.A0(new_n6644_), .A1(new_n6638_), .B0(new_n6643_), .Y(\asquared[65] ));
  AOI21X1  g06452(.A0(new_n6642_), .A1(new_n6640_), .B0(new_n6637_), .Y(new_n6646_));
  INVX1    g06453(.A(new_n6461_), .Y(new_n6647_));
  INVX1    g06454(.A(new_n6487_), .Y(new_n6648_));
  NAND2X1  g06455(.A(new_n6632_), .B(new_n6648_), .Y(new_n6649_));
  OAI21X1  g06456(.A0(new_n6486_), .A1(new_n6647_), .B0(new_n6649_), .Y(new_n6650_));
  AND2X1   g06457(.A(new_n6630_), .B(new_n6308_), .Y(new_n6651_));
  AOI21X1  g06458(.A0(new_n6631_), .A1(new_n6586_), .B0(new_n6651_), .Y(new_n6652_));
  NOR2X1   g06459(.A(new_n6567_), .B(new_n6489_), .Y(new_n6653_));
  AOI21X1  g06460(.A0(new_n6585_), .A1(new_n6568_), .B0(new_n6653_), .Y(new_n6654_));
  NAND2X1  g06461(.A(new_n6599_), .B(new_n6596_), .Y(new_n6655_));
  OAI21X1  g06462(.A0(new_n6629_), .A1(new_n6600_), .B0(new_n6655_), .Y(new_n6656_));
  INVX1    g06463(.A(new_n6515_), .Y(new_n6657_));
  NAND2X1  g06464(.A(new_n6564_), .B(new_n6541_), .Y(new_n6658_));
  OAI21X1  g06465(.A0(new_n6566_), .A1(new_n6657_), .B0(new_n6658_), .Y(new_n6659_));
  NAND2X1  g06466(.A(new_n6627_), .B(new_n6605_), .Y(new_n6660_));
  OAI21X1  g06467(.A0(new_n6604_), .A1(new_n6602_), .B0(new_n6660_), .Y(new_n6661_));
  XOR2X1   g06468(.A(new_n6661_), .B(new_n6659_), .Y(new_n6662_));
  AND2X1   g06469(.A(new_n6625_), .B(new_n6617_), .Y(new_n6663_));
  AOI21X1  g06470(.A0(new_n6626_), .A1(new_n6609_), .B0(new_n6663_), .Y(new_n6664_));
  XOR2X1   g06471(.A(new_n6614_), .B(new_n6512_), .Y(new_n6665_));
  XOR2X1   g06472(.A(new_n6665_), .B(new_n6495_), .Y(new_n6666_));
  XOR2X1   g06473(.A(new_n6561_), .B(new_n6546_), .Y(new_n6667_));
  XOR2X1   g06474(.A(new_n6667_), .B(new_n6522_), .Y(new_n6668_));
  INVX1    g06475(.A(new_n6668_), .Y(new_n6669_));
  XOR2X1   g06476(.A(new_n6669_), .B(new_n6666_), .Y(new_n6670_));
  INVX1    g06477(.A(new_n6670_), .Y(new_n6671_));
  XOR2X1   g06478(.A(new_n6671_), .B(new_n6664_), .Y(new_n6672_));
  XOR2X1   g06479(.A(new_n6672_), .B(new_n6662_), .Y(new_n6673_));
  INVX1    g06480(.A(new_n6673_), .Y(new_n6674_));
  XOR2X1   g06481(.A(new_n6674_), .B(new_n6656_), .Y(new_n6675_));
  XOR2X1   g06482(.A(new_n6675_), .B(new_n6654_), .Y(new_n6676_));
  XOR2X1   g06483(.A(new_n6676_), .B(new_n6652_), .Y(new_n6677_));
  INVX1    g06484(.A(new_n6484_), .Y(new_n6678_));
  NOR2X1   g06485(.A(new_n6678_), .B(new_n6466_), .Y(new_n6679_));
  INVX1    g06486(.A(new_n6485_), .Y(new_n6680_));
  AOI21X1  g06487(.A0(new_n6680_), .A1(new_n6464_), .B0(new_n6679_), .Y(new_n6681_));
  AND2X1   g06488(.A(new_n6572_), .B(new_n6570_), .Y(new_n6682_));
  OR2X1    g06489(.A(new_n6572_), .B(new_n6570_), .Y(new_n6683_));
  OAI21X1  g06490(.A0(new_n6575_), .A1(new_n6682_), .B0(new_n6683_), .Y(new_n6684_));
  OAI21X1  g06491(.A0(new_n6551_), .A1(new_n6550_), .B0(new_n6548_), .Y(new_n6685_));
  OAI21X1  g06492(.A0(new_n6563_), .A1(new_n6553_), .B0(new_n6685_), .Y(new_n6686_));
  XOR2X1   g06493(.A(new_n6686_), .B(new_n6684_), .Y(new_n6687_));
  AND2X1   g06494(.A(\a[63] ), .B(\a[61] ), .Y(new_n6688_));
  NAND2X1  g06495(.A(\a[61] ), .B(\a[4] ), .Y(new_n6689_));
  NAND2X1  g06496(.A(\a[63] ), .B(\a[2] ), .Y(new_n6690_));
  AOI22X1  g06497(.A0(new_n6690_), .A1(new_n6689_), .B0(new_n6688_), .B1(new_n235_), .Y(new_n6691_));
  XOR2X1   g06498(.A(new_n6691_), .B(new_n6539_), .Y(new_n6692_));
  NOR4X1   g06499(.A(new_n4354_), .B(new_n4041_), .C(new_n675_), .D(new_n591_), .Y(new_n6693_));
  NAND4X1  g06500(.A(\a[53] ), .B(\a[52] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n6694_));
  NAND4X1  g06501(.A(\a[53] ), .B(\a[47] ), .C(\a[18] ), .D(\a[12] ), .Y(new_n6695_));
  AOI21X1  g06502(.A0(new_n6695_), .A1(new_n6694_), .B0(new_n6693_), .Y(new_n6696_));
  OR2X1    g06503(.A(new_n6696_), .B(new_n6693_), .Y(new_n6697_));
  AOI22X1  g06504(.A0(\a[52] ), .A1(\a[13] ), .B0(\a[47] ), .B1(\a[18] ), .Y(new_n6698_));
  NAND2X1  g06505(.A(\a[53] ), .B(\a[12] ), .Y(new_n6699_));
  OAI22X1  g06506(.A0(new_n6699_), .A1(new_n6696_), .B0(new_n6698_), .B1(new_n6697_), .Y(new_n6700_));
  NAND4X1  g06507(.A(\a[51] ), .B(\a[49] ), .C(\a[16] ), .D(\a[14] ), .Y(new_n6701_));
  NAND4X1  g06508(.A(\a[50] ), .B(\a[49] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n6702_));
  AOI22X1  g06509(.A0(new_n6702_), .A1(new_n6701_), .B0(new_n4484_), .B1(new_n691_), .Y(new_n6703_));
  AOI22X1  g06510(.A0(\a[51] ), .A1(\a[14] ), .B0(\a[50] ), .B1(\a[15] ), .Y(new_n6704_));
  AOI21X1  g06511(.A0(new_n4484_), .A1(new_n691_), .B0(new_n6703_), .Y(new_n6705_));
  INVX1    g06512(.A(new_n6705_), .Y(new_n6706_));
  OAI22X1  g06513(.A0(new_n6706_), .A1(new_n6704_), .B0(new_n6703_), .B1(new_n5203_), .Y(new_n6707_));
  XOR2X1   g06514(.A(new_n6707_), .B(new_n6700_), .Y(new_n6708_));
  XOR2X1   g06515(.A(new_n6708_), .B(new_n6692_), .Y(new_n6709_));
  XOR2X1   g06516(.A(new_n6709_), .B(new_n6687_), .Y(new_n6710_));
  INVX1    g06517(.A(new_n6530_), .Y(new_n6711_));
  XOR2X1   g06518(.A(new_n6711_), .B(new_n6503_), .Y(new_n6712_));
  XOR2X1   g06519(.A(new_n6712_), .B(new_n6624_), .Y(new_n6713_));
  INVX1    g06520(.A(new_n6523_), .Y(new_n6714_));
  OR2X1    g06521(.A(new_n6532_), .B(new_n6714_), .Y(new_n6715_));
  OAI21X1  g06522(.A0(new_n6540_), .A1(new_n6533_), .B0(new_n6715_), .Y(new_n6716_));
  XOR2X1   g06523(.A(new_n6716_), .B(new_n6713_), .Y(new_n6717_));
  AND2X1   g06524(.A(new_n6505_), .B(new_n6498_), .Y(new_n6718_));
  AND2X1   g06525(.A(new_n6514_), .B(new_n6506_), .Y(new_n6719_));
  OR2X1    g06526(.A(new_n6719_), .B(new_n6718_), .Y(new_n6720_));
  XOR2X1   g06527(.A(new_n6720_), .B(new_n6717_), .Y(new_n6721_));
  INVX1    g06528(.A(new_n6721_), .Y(new_n6722_));
  OR2X1    g06529(.A(new_n6582_), .B(new_n6578_), .Y(new_n6723_));
  OAI21X1  g06530(.A0(new_n6584_), .A1(new_n6576_), .B0(new_n6723_), .Y(new_n6724_));
  XOR2X1   g06531(.A(new_n6724_), .B(new_n6722_), .Y(new_n6725_));
  XOR2X1   g06532(.A(new_n6725_), .B(new_n6710_), .Y(new_n6726_));
  XOR2X1   g06533(.A(new_n6726_), .B(new_n6681_), .Y(new_n6727_));
  AND2X1   g06534(.A(new_n6362_), .B(new_n6338_), .Y(new_n6728_));
  OAI21X1  g06535(.A0(new_n6728_), .A1(new_n6469_), .B0(new_n6468_), .Y(new_n6729_));
  OAI21X1  g06536(.A0(new_n6483_), .A1(new_n6471_), .B0(new_n6729_), .Y(new_n6730_));
  NOR4X1   g06537(.A(new_n4906_), .B(new_n3811_), .C(new_n934_), .D(new_n570_), .Y(new_n6731_));
  NAND4X1  g06538(.A(\a[56] ), .B(\a[45] ), .C(\a[20] ), .D(\a[9] ), .Y(new_n6732_));
  NAND4X1  g06539(.A(\a[56] ), .B(\a[55] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n6733_));
  AOI21X1  g06540(.A0(new_n6733_), .A1(new_n6732_), .B0(new_n6731_), .Y(new_n6734_));
  OR2X1    g06541(.A(new_n6734_), .B(new_n6731_), .Y(new_n6735_));
  AOI22X1  g06542(.A0(\a[55] ), .A1(\a[10] ), .B0(\a[45] ), .B1(\a[20] ), .Y(new_n6736_));
  NAND2X1  g06543(.A(\a[56] ), .B(\a[9] ), .Y(new_n6737_));
  OAI22X1  g06544(.A0(new_n6737_), .A1(new_n6734_), .B0(new_n6736_), .B1(new_n6735_), .Y(new_n6738_));
  NAND4X1  g06545(.A(\a[42] ), .B(\a[40] ), .C(\a[25] ), .D(\a[23] ), .Y(new_n6739_));
  NAND4X1  g06546(.A(\a[42] ), .B(\a[41] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n6740_));
  AOI22X1  g06547(.A0(new_n6740_), .A1(new_n6739_), .B0(new_n4404_), .B1(new_n1532_), .Y(new_n6741_));
  NAND2X1  g06548(.A(\a[42] ), .B(\a[23] ), .Y(new_n6742_));
  AOI22X1  g06549(.A0(\a[41] ), .A1(\a[24] ), .B0(\a[40] ), .B1(\a[25] ), .Y(new_n6743_));
  AOI21X1  g06550(.A0(new_n4404_), .A1(new_n1532_), .B0(new_n6741_), .Y(new_n6744_));
  INVX1    g06551(.A(new_n6744_), .Y(new_n6745_));
  OAI22X1  g06552(.A0(new_n6745_), .A1(new_n6743_), .B0(new_n6742_), .B1(new_n6741_), .Y(new_n6746_));
  XOR2X1   g06553(.A(new_n6746_), .B(new_n6738_), .Y(new_n6747_));
  AOI22X1  g06554(.A0(new_n3730_), .A1(new_n1996_), .B0(new_n3503_), .B1(new_n1995_), .Y(new_n6748_));
  AOI21X1  g06555(.A0(new_n3164_), .A1(new_n1671_), .B0(new_n6748_), .Y(new_n6749_));
  AND2X1   g06556(.A(\a[39] ), .B(\a[26] ), .Y(new_n6750_));
  INVX1    g06557(.A(new_n6750_), .Y(new_n6751_));
  OAI22X1  g06558(.A0(new_n3731_), .A1(new_n3570_), .B0(new_n3729_), .B1(new_n3483_), .Y(new_n6752_));
  AOI21X1  g06559(.A0(new_n3164_), .A1(new_n1671_), .B0(new_n6752_), .Y(new_n6753_));
  INVX1    g06560(.A(new_n6753_), .Y(new_n6754_));
  AOI22X1  g06561(.A0(\a[38] ), .A1(\a[27] ), .B0(\a[37] ), .B1(\a[28] ), .Y(new_n6755_));
  OAI22X1  g06562(.A0(new_n6755_), .A1(new_n6754_), .B0(new_n6751_), .B1(new_n6749_), .Y(new_n6756_));
  INVX1    g06563(.A(new_n6756_), .Y(new_n6757_));
  XOR2X1   g06564(.A(new_n6757_), .B(new_n6747_), .Y(new_n6758_));
  AOI22X1  g06565(.A0(\a[54] ), .A1(\a[11] ), .B0(\a[46] ), .B1(\a[19] ), .Y(new_n6759_));
  AND2X1   g06566(.A(\a[36] ), .B(\a[29] ), .Y(new_n6760_));
  INVX1    g06567(.A(new_n6760_), .Y(new_n6761_));
  NOR4X1   g06568(.A(new_n4835_), .B(new_n3460_), .C(new_n752_), .D(new_n488_), .Y(new_n6762_));
  NOR3X1   g06569(.A(new_n6761_), .B(new_n6762_), .C(new_n6759_), .Y(new_n6763_));
  NOR2X1   g06570(.A(new_n6763_), .B(new_n6762_), .Y(new_n6764_));
  INVX1    g06571(.A(new_n6764_), .Y(new_n6765_));
  OAI22X1  g06572(.A0(new_n6765_), .A1(new_n6759_), .B0(new_n6763_), .B1(new_n6761_), .Y(new_n6766_));
  NAND4X1  g06573(.A(\a[35] ), .B(\a[33] ), .C(\a[32] ), .D(\a[30] ), .Y(new_n6767_));
  OAI21X1  g06574(.A0(new_n4915_), .A1(new_n2076_), .B0(new_n6767_), .Y(new_n6768_));
  OAI21X1  g06575(.A0(new_n2919_), .A1(new_n2672_), .B0(new_n6768_), .Y(new_n6769_));
  AOI21X1  g06576(.A0(new_n2918_), .A1(new_n2671_), .B0(new_n6768_), .Y(new_n6770_));
  OAI22X1  g06577(.A0(new_n2028_), .A1(new_n1704_), .B0(new_n1851_), .B1(new_n2219_), .Y(new_n6771_));
  AOI22X1  g06578(.A0(new_n6771_), .A1(new_n6770_), .B0(new_n6769_), .B1(new_n2779_), .Y(new_n6772_));
  XOR2X1   g06579(.A(new_n6772_), .B(new_n6766_), .Y(new_n6773_));
  AND2X1   g06580(.A(\a[48] ), .B(\a[17] ), .Y(new_n6774_));
  NOR3X1   g06581(.A(new_n6606_), .B(new_n1851_), .C(new_n223_), .Y(new_n6775_));
  AOI21X1  g06582(.A0(\a[62] ), .A1(\a[3] ), .B0(\a[33] ), .Y(new_n6776_));
  OR4X1    g06583(.A(new_n6776_), .B(new_n6775_), .C(new_n3926_), .D(new_n616_), .Y(new_n6777_));
  NOR3X1   g06584(.A(new_n6776_), .B(new_n6775_), .C(new_n6774_), .Y(new_n6778_));
  AOI21X1  g06585(.A0(new_n6777_), .A1(new_n6774_), .B0(new_n6778_), .Y(new_n6779_));
  XOR2X1   g06586(.A(new_n6779_), .B(new_n6773_), .Y(new_n6780_));
  AOI22X1  g06587(.A0(\a[44] ), .A1(\a[21] ), .B0(\a[43] ), .B1(\a[22] ), .Y(new_n6781_));
  AND2X1   g06588(.A(\a[57] ), .B(\a[8] ), .Y(new_n6782_));
  AND2X1   g06589(.A(new_n4992_), .B(new_n1154_), .Y(new_n6783_));
  OAI21X1  g06590(.A0(new_n6781_), .A1(new_n6783_), .B0(new_n6782_), .Y(new_n6784_));
  INVX1    g06591(.A(new_n6781_), .Y(new_n6785_));
  AOI21X1  g06592(.A0(new_n6785_), .A1(new_n6782_), .B0(new_n6783_), .Y(new_n6786_));
  INVX1    g06593(.A(new_n6786_), .Y(new_n6787_));
  OAI21X1  g06594(.A0(new_n6787_), .A1(new_n6781_), .B0(new_n6784_), .Y(new_n6788_));
  AND2X1   g06595(.A(\a[63] ), .B(\a[62] ), .Y(new_n6789_));
  NOR2X1   g06596(.A(new_n6608_), .B(new_n6414_), .Y(new_n6790_));
  AOI21X1  g06597(.A0(new_n6789_), .A1(new_n1913_), .B0(new_n6790_), .Y(new_n6791_));
  XOR2X1   g06598(.A(new_n6791_), .B(new_n6788_), .Y(new_n6792_));
  INVX1    g06599(.A(new_n6121_), .Y(new_n6793_));
  INVX1    g06600(.A(new_n6427_), .Y(new_n6794_));
  AND2X1   g06601(.A(\a[60] ), .B(\a[58] ), .Y(new_n6795_));
  INVX1    g06602(.A(new_n6795_), .Y(new_n6796_));
  OAI22X1  g06603(.A0(new_n6796_), .A1(new_n678_), .B0(new_n6794_), .B1(new_n444_), .Y(new_n6797_));
  OAI21X1  g06604(.A0(new_n6793_), .A1(new_n376_), .B0(new_n6797_), .Y(new_n6798_));
  AND2X1   g06605(.A(\a[60] ), .B(\a[5] ), .Y(new_n6799_));
  AOI21X1  g06606(.A0(new_n6121_), .A1(new_n375_), .B0(new_n6797_), .Y(new_n6800_));
  OAI22X1  g06607(.A0(new_n5617_), .A1(new_n230_), .B0(new_n5379_), .B1(new_n532_), .Y(new_n6801_));
  AOI22X1  g06608(.A0(new_n6801_), .A1(new_n6800_), .B0(new_n6799_), .B1(new_n6798_), .Y(new_n6802_));
  XOR2X1   g06609(.A(new_n6802_), .B(new_n6792_), .Y(new_n6803_));
  INVX1    g06610(.A(new_n6803_), .Y(new_n6804_));
  XOR2X1   g06611(.A(new_n6804_), .B(new_n6780_), .Y(new_n6805_));
  XOR2X1   g06612(.A(new_n6805_), .B(new_n6758_), .Y(new_n6806_));
  XOR2X1   g06613(.A(new_n6806_), .B(new_n6730_), .Y(new_n6807_));
  AND2X1   g06614(.A(new_n6396_), .B(new_n6350_), .Y(new_n6808_));
  AOI21X1  g06615(.A0(new_n6587_), .A1(new_n6387_), .B0(new_n6808_), .Y(new_n6809_));
  AND2X1   g06616(.A(new_n6407_), .B(new_n6376_), .Y(new_n6810_));
  AOI21X1  g06617(.A0(new_n6474_), .A1(new_n6359_), .B0(new_n6810_), .Y(new_n6811_));
  XOR2X1   g06618(.A(new_n6811_), .B(new_n6809_), .Y(new_n6812_));
  INVX1    g06619(.A(new_n6812_), .Y(new_n6813_));
  NOR2X1   g06620(.A(new_n6443_), .B(new_n6433_), .Y(new_n6814_));
  AOI21X1  g06621(.A0(new_n6477_), .A1(new_n6476_), .B0(new_n6814_), .Y(new_n6815_));
  XOR2X1   g06622(.A(new_n6815_), .B(new_n6813_), .Y(new_n6816_));
  OR2X1    g06623(.A(new_n6479_), .B(new_n6475_), .Y(new_n6817_));
  OAI21X1  g06624(.A0(new_n6481_), .A1(new_n6473_), .B0(new_n6817_), .Y(new_n6818_));
  AND2X1   g06625(.A(new_n6591_), .B(new_n6588_), .Y(new_n6819_));
  AOI21X1  g06626(.A0(new_n6595_), .A1(new_n6592_), .B0(new_n6819_), .Y(new_n6820_));
  XOR2X1   g06627(.A(new_n6820_), .B(new_n6818_), .Y(new_n6821_));
  XOR2X1   g06628(.A(new_n6821_), .B(new_n6816_), .Y(new_n6822_));
  XOR2X1   g06629(.A(new_n6822_), .B(new_n6807_), .Y(new_n6823_));
  INVX1    g06630(.A(new_n6823_), .Y(new_n6824_));
  XOR2X1   g06631(.A(new_n6824_), .B(new_n6727_), .Y(new_n6825_));
  XOR2X1   g06632(.A(new_n6825_), .B(new_n6677_), .Y(new_n6826_));
  AND2X1   g06633(.A(new_n6826_), .B(new_n6650_), .Y(new_n6827_));
  NOR2X1   g06634(.A(new_n6826_), .B(new_n6650_), .Y(new_n6828_));
  OR2X1    g06635(.A(new_n6828_), .B(new_n6827_), .Y(new_n6829_));
  XOR2X1   g06636(.A(new_n6829_), .B(new_n6646_), .Y(\asquared[66] ));
  INVX1    g06637(.A(new_n6827_), .Y(new_n6831_));
  OAI21X1  g06638(.A0(new_n6828_), .A1(new_n6646_), .B0(new_n6831_), .Y(new_n6832_));
  INVX1    g06639(.A(new_n6652_), .Y(new_n6833_));
  NOR2X1   g06640(.A(new_n6825_), .B(new_n6677_), .Y(new_n6834_));
  AOI21X1  g06641(.A0(new_n6676_), .A1(new_n6833_), .B0(new_n6834_), .Y(new_n6835_));
  INVX1    g06642(.A(new_n6726_), .Y(new_n6836_));
  NOR2X1   g06643(.A(new_n6836_), .B(new_n6681_), .Y(new_n6837_));
  NOR2X1   g06644(.A(new_n6823_), .B(new_n6727_), .Y(new_n6838_));
  NOR2X1   g06645(.A(new_n6838_), .B(new_n6837_), .Y(new_n6839_));
  INVX1    g06646(.A(new_n6821_), .Y(new_n6840_));
  INVX1    g06647(.A(new_n6818_), .Y(new_n6841_));
  NOR2X1   g06648(.A(new_n6820_), .B(new_n6841_), .Y(new_n6842_));
  AOI21X1  g06649(.A0(new_n6840_), .A1(new_n6816_), .B0(new_n6842_), .Y(new_n6843_));
  INVX1    g06650(.A(new_n6539_), .Y(new_n6844_));
  AOI22X1  g06651(.A0(new_n6691_), .A1(new_n6844_), .B0(new_n6688_), .B1(new_n235_), .Y(new_n6845_));
  XOR2X1   g06652(.A(new_n6845_), .B(new_n6753_), .Y(new_n6846_));
  OAI22X1  g06653(.A0(new_n6796_), .A1(new_n280_), .B0(new_n6794_), .B1(new_n376_), .Y(new_n6847_));
  OAI21X1  g06654(.A0(new_n6793_), .A1(new_n445_), .B0(new_n6847_), .Y(new_n6848_));
  AND2X1   g06655(.A(\a[60] ), .B(\a[6] ), .Y(new_n6849_));
  AOI21X1  g06656(.A0(new_n6121_), .A1(new_n325_), .B0(new_n6847_), .Y(new_n6850_));
  OAI22X1  g06657(.A0(new_n5617_), .A1(new_n532_), .B0(new_n5379_), .B1(new_n413_), .Y(new_n6851_));
  AOI22X1  g06658(.A0(new_n6851_), .A1(new_n6850_), .B0(new_n6849_), .B1(new_n6848_), .Y(new_n6852_));
  XOR2X1   g06659(.A(new_n6852_), .B(new_n6846_), .Y(new_n6853_));
  INVX1    g06660(.A(new_n6692_), .Y(new_n6854_));
  AND2X1   g06661(.A(new_n6707_), .B(new_n6700_), .Y(new_n6855_));
  AOI21X1  g06662(.A0(new_n6708_), .A1(new_n6854_), .B0(new_n6855_), .Y(new_n6856_));
  XOR2X1   g06663(.A(new_n6856_), .B(new_n6853_), .Y(new_n6857_));
  OR2X1    g06664(.A(new_n6811_), .B(new_n6809_), .Y(new_n6858_));
  OAI21X1  g06665(.A0(new_n6815_), .A1(new_n6813_), .B0(new_n6858_), .Y(new_n6859_));
  XOR2X1   g06666(.A(new_n6859_), .B(new_n6857_), .Y(new_n6860_));
  NOR3X1   g06667(.A(new_n6776_), .B(new_n3926_), .C(new_n616_), .Y(new_n6861_));
  NOR2X1   g06668(.A(new_n6861_), .B(new_n6775_), .Y(new_n6862_));
  XOR2X1   g06669(.A(new_n6862_), .B(new_n6770_), .Y(new_n6863_));
  XOR2X1   g06670(.A(new_n6863_), .B(new_n6705_), .Y(new_n6864_));
  XOR2X1   g06671(.A(new_n6800_), .B(new_n6786_), .Y(new_n6865_));
  XOR2X1   g06672(.A(new_n6865_), .B(new_n6765_), .Y(new_n6866_));
  INVX1    g06673(.A(new_n6766_), .Y(new_n6867_));
  OR2X1    g06674(.A(new_n6772_), .B(new_n6867_), .Y(new_n6868_));
  OAI21X1  g06675(.A0(new_n6779_), .A1(new_n6773_), .B0(new_n6868_), .Y(new_n6869_));
  XOR2X1   g06676(.A(new_n6869_), .B(new_n6866_), .Y(new_n6870_));
  INVX1    g06677(.A(new_n6870_), .Y(new_n6871_));
  XOR2X1   g06678(.A(new_n6871_), .B(new_n6864_), .Y(new_n6872_));
  XOR2X1   g06679(.A(new_n6872_), .B(new_n6860_), .Y(new_n6873_));
  INVX1    g06680(.A(new_n6873_), .Y(new_n6874_));
  XOR2X1   g06681(.A(new_n6874_), .B(new_n6843_), .Y(new_n6875_));
  NOR2X1   g06682(.A(new_n6725_), .B(new_n6710_), .Y(new_n6876_));
  AOI21X1  g06683(.A0(new_n6724_), .A1(new_n6721_), .B0(new_n6876_), .Y(new_n6877_));
  XOR2X1   g06684(.A(new_n6735_), .B(new_n6697_), .Y(new_n6878_));
  XOR2X1   g06685(.A(new_n6878_), .B(new_n6744_), .Y(new_n6879_));
  INVX1    g06686(.A(new_n6791_), .Y(new_n6880_));
  NOR2X1   g06687(.A(new_n6802_), .B(new_n6792_), .Y(new_n6881_));
  AOI21X1  g06688(.A0(new_n6880_), .A1(new_n6788_), .B0(new_n6881_), .Y(new_n6882_));
  XOR2X1   g06689(.A(new_n6882_), .B(new_n6879_), .Y(new_n6883_));
  AND2X1   g06690(.A(new_n6746_), .B(new_n6738_), .Y(new_n6884_));
  AND2X1   g06691(.A(new_n6756_), .B(new_n6747_), .Y(new_n6885_));
  OR2X1    g06692(.A(new_n6885_), .B(new_n6884_), .Y(new_n6886_));
  XOR2X1   g06693(.A(new_n6886_), .B(new_n6883_), .Y(new_n6887_));
  NAND2X1  g06694(.A(new_n6803_), .B(new_n6780_), .Y(new_n6888_));
  OAI21X1  g06695(.A0(new_n6805_), .A1(new_n6758_), .B0(new_n6888_), .Y(new_n6889_));
  AND2X1   g06696(.A(new_n6686_), .B(new_n6684_), .Y(new_n6890_));
  INVX1    g06697(.A(new_n6709_), .Y(new_n6891_));
  AOI21X1  g06698(.A0(new_n6891_), .A1(new_n6687_), .B0(new_n6890_), .Y(new_n6892_));
  INVX1    g06699(.A(new_n6892_), .Y(new_n6893_));
  XOR2X1   g06700(.A(new_n6893_), .B(new_n6889_), .Y(new_n6894_));
  XOR2X1   g06701(.A(new_n6894_), .B(new_n6887_), .Y(new_n6895_));
  XOR2X1   g06702(.A(new_n6895_), .B(new_n6877_), .Y(new_n6896_));
  XOR2X1   g06703(.A(new_n6896_), .B(new_n6875_), .Y(new_n6897_));
  XOR2X1   g06704(.A(new_n6897_), .B(new_n6839_), .Y(new_n6898_));
  INVX1    g06705(.A(new_n6898_), .Y(new_n6899_));
  NAND2X1  g06706(.A(new_n6673_), .B(new_n6656_), .Y(new_n6900_));
  OAI21X1  g06707(.A0(new_n6675_), .A1(new_n6654_), .B0(new_n6900_), .Y(new_n6901_));
  NAND2X1  g06708(.A(new_n6806_), .B(new_n6730_), .Y(new_n6902_));
  INVX1    g06709(.A(new_n6807_), .Y(new_n6903_));
  OAI21X1  g06710(.A0(new_n6822_), .A1(new_n6903_), .B0(new_n6902_), .Y(new_n6904_));
  XOR2X1   g06711(.A(new_n6904_), .B(new_n6901_), .Y(new_n6905_));
  AND2X1   g06712(.A(new_n6661_), .B(new_n6659_), .Y(new_n6906_));
  AOI21X1  g06713(.A0(new_n6672_), .A1(new_n6662_), .B0(new_n6906_), .Y(new_n6907_));
  NAND4X1  g06714(.A(\a[63] ), .B(\a[61] ), .C(\a[5] ), .D(\a[3] ), .Y(new_n6908_));
  NAND4X1  g06715(.A(\a[63] ), .B(\a[62] ), .C(\a[4] ), .D(\a[3] ), .Y(new_n6909_));
  AOI22X1  g06716(.A0(new_n6909_), .A1(new_n6908_), .B0(new_n6556_), .B1(new_n218_), .Y(new_n6910_));
  NAND4X1  g06717(.A(\a[62] ), .B(\a[61] ), .C(\a[5] ), .D(\a[4] ), .Y(new_n6911_));
  NAND3X1  g06718(.A(new_n6909_), .B(new_n6908_), .C(new_n6911_), .Y(new_n6912_));
  AOI22X1  g06719(.A0(\a[62] ), .A1(\a[4] ), .B0(\a[61] ), .B1(\a[5] ), .Y(new_n6913_));
  NAND2X1  g06720(.A(\a[63] ), .B(\a[3] ), .Y(new_n6914_));
  OAI22X1  g06721(.A0(new_n6914_), .A1(new_n6910_), .B0(new_n6913_), .B1(new_n6912_), .Y(new_n6915_));
  NAND4X1  g06722(.A(\a[39] ), .B(\a[37] ), .C(\a[29] ), .D(\a[27] ), .Y(new_n6916_));
  NAND4X1  g06723(.A(\a[39] ), .B(\a[38] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n6917_));
  AOI22X1  g06724(.A0(new_n6917_), .A1(new_n6916_), .B0(new_n3164_), .B1(new_n1674_), .Y(new_n6918_));
  NAND2X1  g06725(.A(\a[39] ), .B(\a[27] ), .Y(new_n6919_));
  AOI22X1  g06726(.A0(\a[38] ), .A1(\a[28] ), .B0(\a[37] ), .B1(\a[29] ), .Y(new_n6920_));
  AOI21X1  g06727(.A0(new_n3164_), .A1(new_n1674_), .B0(new_n6918_), .Y(new_n6921_));
  INVX1    g06728(.A(new_n6921_), .Y(new_n6922_));
  OAI22X1  g06729(.A0(new_n6922_), .A1(new_n6920_), .B0(new_n6919_), .B1(new_n6918_), .Y(new_n6923_));
  XOR2X1   g06730(.A(new_n6923_), .B(new_n6915_), .Y(new_n6924_));
  NOR4X1   g06731(.A(new_n4835_), .B(new_n4041_), .C(new_n752_), .D(new_n453_), .Y(new_n6925_));
  AND2X1   g06732(.A(\a[47] ), .B(\a[11] ), .Y(new_n6926_));
  AOI22X1  g06733(.A0(new_n5561_), .A1(new_n6926_), .B0(new_n5240_), .B1(new_n482_), .Y(new_n6927_));
  AND2X1   g06734(.A(\a[55] ), .B(\a[11] ), .Y(new_n6928_));
  OAI21X1  g06735(.A0(new_n6927_), .A1(new_n6925_), .B0(new_n6928_), .Y(new_n6929_));
  INVX1    g06736(.A(new_n6925_), .Y(new_n6930_));
  AND2X1   g06737(.A(new_n6927_), .B(new_n6930_), .Y(new_n6931_));
  INVX1    g06738(.A(new_n6931_), .Y(new_n6932_));
  AOI22X1  g06739(.A0(\a[54] ), .A1(\a[12] ), .B0(\a[47] ), .B1(\a[19] ), .Y(new_n6933_));
  OAI21X1  g06740(.A0(new_n6933_), .A1(new_n6932_), .B0(new_n6929_), .Y(new_n6934_));
  INVX1    g06741(.A(new_n6934_), .Y(new_n6935_));
  XOR2X1   g06742(.A(new_n6935_), .B(new_n6924_), .Y(new_n6936_));
  AND2X1   g06743(.A(\a[57] ), .B(\a[24] ), .Y(new_n6937_));
  NAND4X1  g06744(.A(\a[57] ), .B(\a[43] ), .C(\a[23] ), .D(\a[9] ), .Y(new_n6938_));
  NAND4X1  g06745(.A(\a[43] ), .B(\a[42] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n6939_));
  AOI22X1  g06746(.A0(new_n6939_), .A1(new_n6938_), .B0(new_n6937_), .B1(new_n4227_), .Y(new_n6940_));
  NAND4X1  g06747(.A(\a[57] ), .B(\a[42] ), .C(\a[24] ), .D(\a[9] ), .Y(new_n6941_));
  NAND3X1  g06748(.A(new_n6939_), .B(new_n6938_), .C(new_n6941_), .Y(new_n6942_));
  AOI22X1  g06749(.A0(\a[57] ), .A1(\a[9] ), .B0(\a[42] ), .B1(\a[24] ), .Y(new_n6943_));
  NAND2X1  g06750(.A(\a[43] ), .B(\a[23] ), .Y(new_n6944_));
  OAI22X1  g06751(.A0(new_n6944_), .A1(new_n6940_), .B0(new_n6943_), .B1(new_n6942_), .Y(new_n6945_));
  NAND4X1  g06752(.A(\a[46] ), .B(\a[44] ), .C(\a[22] ), .D(\a[20] ), .Y(new_n6946_));
  NAND4X1  g06753(.A(\a[46] ), .B(\a[45] ), .C(\a[21] ), .D(\a[20] ), .Y(new_n6947_));
  AOI22X1  g06754(.A0(new_n6947_), .A1(new_n6946_), .B0(new_n3918_), .B1(new_n1154_), .Y(new_n6948_));
  NAND2X1  g06755(.A(\a[46] ), .B(\a[20] ), .Y(new_n6949_));
  AOI22X1  g06756(.A0(\a[45] ), .A1(\a[21] ), .B0(\a[44] ), .B1(\a[22] ), .Y(new_n6950_));
  AOI21X1  g06757(.A0(new_n3918_), .A1(new_n1154_), .B0(new_n6948_), .Y(new_n6951_));
  INVX1    g06758(.A(new_n6951_), .Y(new_n6952_));
  OAI22X1  g06759(.A0(new_n6952_), .A1(new_n6950_), .B0(new_n6949_), .B1(new_n6948_), .Y(new_n6953_));
  XOR2X1   g06760(.A(new_n6953_), .B(new_n6945_), .Y(new_n6954_));
  AND2X1   g06761(.A(\a[56] ), .B(\a[10] ), .Y(new_n6955_));
  INVX1    g06762(.A(new_n6955_), .Y(new_n6956_));
  AOI22X1  g06763(.A0(\a[41] ), .A1(\a[25] ), .B0(\a[40] ), .B1(\a[26] ), .Y(new_n6957_));
  AND2X1   g06764(.A(new_n4404_), .B(new_n1770_), .Y(new_n6958_));
  NOR3X1   g06765(.A(new_n6957_), .B(new_n6958_), .C(new_n6956_), .Y(new_n6959_));
  NOR2X1   g06766(.A(new_n6959_), .B(new_n6958_), .Y(new_n6960_));
  INVX1    g06767(.A(new_n6960_), .Y(new_n6961_));
  OAI22X1  g06768(.A0(new_n6961_), .A1(new_n6957_), .B0(new_n6959_), .B1(new_n6956_), .Y(new_n6962_));
  XOR2X1   g06769(.A(new_n6962_), .B(new_n6954_), .Y(new_n6963_));
  AOI22X1  g06770(.A0(\a[53] ), .A1(\a[13] ), .B0(\a[51] ), .B1(\a[15] ), .Y(new_n6964_));
  AND2X1   g06771(.A(\a[48] ), .B(\a[18] ), .Y(new_n6965_));
  INVX1    g06772(.A(new_n6965_), .Y(new_n6966_));
  AND2X1   g06773(.A(new_n4904_), .B(new_n639_), .Y(new_n6967_));
  NOR3X1   g06774(.A(new_n6966_), .B(new_n6967_), .C(new_n6964_), .Y(new_n6968_));
  INVX1    g06775(.A(new_n6964_), .Y(new_n6969_));
  AOI21X1  g06776(.A0(new_n6965_), .A1(new_n6969_), .B0(new_n6967_), .Y(new_n6970_));
  INVX1    g06777(.A(new_n6970_), .Y(new_n6971_));
  OAI22X1  g06778(.A0(new_n6971_), .A1(new_n6964_), .B0(new_n6968_), .B1(new_n6966_), .Y(new_n6972_));
  AND2X1   g06779(.A(\a[52] ), .B(\a[14] ), .Y(new_n6973_));
  AOI22X1  g06780(.A0(\a[36] ), .A1(\a[30] ), .B0(\a[35] ), .B1(\a[31] ), .Y(new_n6974_));
  INVX1    g06781(.A(new_n6974_), .Y(new_n6975_));
  NAND4X1  g06782(.A(\a[36] ), .B(\a[35] ), .C(\a[31] ), .D(\a[30] ), .Y(new_n6976_));
  NAND3X1  g06783(.A(new_n6975_), .B(new_n6976_), .C(new_n6973_), .Y(new_n6977_));
  AOI22X1  g06784(.A0(new_n6975_), .A1(new_n6973_), .B0(new_n2682_), .B1(new_n2075_), .Y(new_n6978_));
  AOI22X1  g06785(.A0(new_n6978_), .A1(new_n6975_), .B0(new_n6977_), .B1(new_n6973_), .Y(new_n6979_));
  XOR2X1   g06786(.A(new_n6979_), .B(new_n6972_), .Y(new_n6980_));
  AOI22X1  g06787(.A0(\a[50] ), .A1(\a[16] ), .B0(\a[49] ), .B1(\a[17] ), .Y(new_n6981_));
  INVX1    g06788(.A(new_n6981_), .Y(new_n6982_));
  NAND4X1  g06789(.A(\a[50] ), .B(\a[49] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n6983_));
  AOI21X1  g06790(.A0(new_n6982_), .A1(new_n6983_), .B0(new_n2920_), .Y(new_n6984_));
  AOI22X1  g06791(.A0(new_n6982_), .A1(new_n2820_), .B0(new_n4321_), .B1(new_n792_), .Y(new_n6985_));
  AOI21X1  g06792(.A0(new_n6985_), .A1(new_n6982_), .B0(new_n6984_), .Y(new_n6986_));
  XOR2X1   g06793(.A(new_n6986_), .B(new_n6980_), .Y(new_n6987_));
  INVX1    g06794(.A(new_n6987_), .Y(new_n6988_));
  XOR2X1   g06795(.A(new_n6988_), .B(new_n6963_), .Y(new_n6989_));
  XOR2X1   g06796(.A(new_n6989_), .B(new_n6936_), .Y(new_n6990_));
  XOR2X1   g06797(.A(new_n6990_), .B(new_n6907_), .Y(new_n6991_));
  AND2X1   g06798(.A(new_n6614_), .B(new_n6512_), .Y(new_n6992_));
  AOI21X1  g06799(.A0(new_n6665_), .A1(new_n6496_), .B0(new_n6992_), .Y(new_n6993_));
  NOR2X1   g06800(.A(new_n6561_), .B(new_n6546_), .Y(new_n6994_));
  AOI21X1  g06801(.A0(new_n6667_), .A1(new_n6522_), .B0(new_n6994_), .Y(new_n6995_));
  XOR2X1   g06802(.A(new_n6995_), .B(new_n6993_), .Y(new_n6996_));
  INVX1    g06803(.A(new_n6996_), .Y(new_n6997_));
  AND2X1   g06804(.A(new_n6711_), .B(new_n6503_), .Y(new_n6998_));
  AOI21X1  g06805(.A0(new_n6712_), .A1(new_n6624_), .B0(new_n6998_), .Y(new_n6999_));
  XOR2X1   g06806(.A(new_n6999_), .B(new_n6997_), .Y(new_n7000_));
  OR2X1    g06807(.A(new_n6669_), .B(new_n6666_), .Y(new_n7001_));
  OAI21X1  g06808(.A0(new_n6671_), .A1(new_n6664_), .B0(new_n7001_), .Y(new_n7002_));
  AND2X1   g06809(.A(new_n6716_), .B(new_n6713_), .Y(new_n7003_));
  AOI21X1  g06810(.A0(new_n6720_), .A1(new_n6717_), .B0(new_n7003_), .Y(new_n7004_));
  XOR2X1   g06811(.A(new_n7004_), .B(new_n7002_), .Y(new_n7005_));
  XOR2X1   g06812(.A(new_n7005_), .B(new_n7000_), .Y(new_n7006_));
  XOR2X1   g06813(.A(new_n7006_), .B(new_n6991_), .Y(new_n7007_));
  XOR2X1   g06814(.A(new_n7007_), .B(new_n6905_), .Y(new_n7008_));
  XOR2X1   g06815(.A(new_n7008_), .B(new_n6899_), .Y(new_n7009_));
  XOR2X1   g06816(.A(new_n7009_), .B(new_n6835_), .Y(new_n7010_));
  XOR2X1   g06817(.A(new_n7010_), .B(new_n6832_), .Y(\asquared[67] ));
  NAND2X1  g06818(.A(new_n7008_), .B(new_n6898_), .Y(new_n7012_));
  OAI21X1  g06819(.A0(new_n6897_), .A1(new_n6839_), .B0(new_n7012_), .Y(new_n7013_));
  AND2X1   g06820(.A(new_n6904_), .B(new_n6901_), .Y(new_n7014_));
  AOI21X1  g06821(.A0(new_n7007_), .A1(new_n6905_), .B0(new_n7014_), .Y(new_n7015_));
  NAND2X1  g06822(.A(new_n6872_), .B(new_n6860_), .Y(new_n7016_));
  OAI21X1  g06823(.A0(new_n6874_), .A1(new_n6843_), .B0(new_n7016_), .Y(new_n7017_));
  INVX1    g06824(.A(new_n7005_), .Y(new_n7018_));
  INVX1    g06825(.A(new_n7002_), .Y(new_n7019_));
  NOR2X1   g06826(.A(new_n7004_), .B(new_n7019_), .Y(new_n7020_));
  AOI21X1  g06827(.A0(new_n7018_), .A1(new_n7000_), .B0(new_n7020_), .Y(new_n7021_));
  AND2X1   g06828(.A(new_n6953_), .B(new_n6945_), .Y(new_n7022_));
  AOI21X1  g06829(.A0(new_n6962_), .A1(new_n6954_), .B0(new_n7022_), .Y(new_n7023_));
  AND2X1   g06830(.A(new_n6845_), .B(new_n6753_), .Y(new_n7024_));
  OR2X1    g06831(.A(new_n6845_), .B(new_n6753_), .Y(new_n7025_));
  OAI21X1  g06832(.A0(new_n6852_), .A1(new_n7024_), .B0(new_n7025_), .Y(new_n7026_));
  INVX1    g06833(.A(new_n7026_), .Y(new_n7027_));
  XOR2X1   g06834(.A(new_n7027_), .B(new_n7023_), .Y(new_n7028_));
  AND2X1   g06835(.A(new_n6923_), .B(new_n6915_), .Y(new_n7029_));
  AOI21X1  g06836(.A0(new_n6934_), .A1(new_n6924_), .B0(new_n7029_), .Y(new_n7030_));
  XOR2X1   g06837(.A(new_n7030_), .B(new_n7028_), .Y(new_n7031_));
  INVX1    g06838(.A(new_n6850_), .Y(new_n7032_));
  XOR2X1   g06839(.A(new_n6912_), .B(new_n7032_), .Y(new_n7033_));
  XOR2X1   g06840(.A(new_n7033_), .B(new_n6921_), .Y(new_n7034_));
  XOR2X1   g06841(.A(new_n6961_), .B(new_n6942_), .Y(new_n7035_));
  XOR2X1   g06842(.A(new_n7035_), .B(new_n6951_), .Y(new_n7036_));
  AND2X1   g06843(.A(\a[61] ), .B(\a[6] ), .Y(new_n7037_));
  INVX1    g06844(.A(new_n7037_), .Y(new_n7038_));
  XOR2X1   g06845(.A(new_n7038_), .B(new_n6985_), .Y(new_n7039_));
  INVX1    g06846(.A(new_n7039_), .Y(new_n7040_));
  XOR2X1   g06847(.A(new_n7040_), .B(new_n6978_), .Y(new_n7041_));
  INVX1    g06848(.A(new_n7041_), .Y(new_n7042_));
  XOR2X1   g06849(.A(new_n7042_), .B(new_n7036_), .Y(new_n7043_));
  INVX1    g06850(.A(new_n7043_), .Y(new_n7044_));
  XOR2X1   g06851(.A(new_n7044_), .B(new_n7034_), .Y(new_n7045_));
  INVX1    g06852(.A(new_n7045_), .Y(new_n7046_));
  XOR2X1   g06853(.A(new_n7046_), .B(new_n7031_), .Y(new_n7047_));
  INVX1    g06854(.A(new_n7047_), .Y(new_n7048_));
  XOR2X1   g06855(.A(new_n7048_), .B(new_n7021_), .Y(new_n7049_));
  XOR2X1   g06856(.A(new_n7049_), .B(new_n7017_), .Y(new_n7050_));
  XOR2X1   g06857(.A(new_n6971_), .B(new_n6931_), .Y(new_n7051_));
  AND2X1   g06858(.A(\a[56] ), .B(\a[20] ), .Y(new_n7052_));
  NAND4X1  g06859(.A(\a[57] ), .B(\a[56] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n7053_));
  NAND4X1  g06860(.A(\a[57] ), .B(\a[47] ), .C(\a[20] ), .D(\a[10] ), .Y(new_n7054_));
  AOI22X1  g06861(.A0(new_n7054_), .A1(new_n7053_), .B0(new_n7052_), .B1(new_n6926_), .Y(new_n7055_));
  AND2X1   g06862(.A(\a[57] ), .B(\a[10] ), .Y(new_n7056_));
  INVX1    g06863(.A(new_n7056_), .Y(new_n7057_));
  AOI21X1  g06864(.A0(new_n7052_), .A1(new_n6926_), .B0(new_n7055_), .Y(new_n7058_));
  INVX1    g06865(.A(new_n7058_), .Y(new_n7059_));
  AOI22X1  g06866(.A0(\a[56] ), .A1(\a[11] ), .B0(\a[47] ), .B1(\a[20] ), .Y(new_n7060_));
  OAI22X1  g06867(.A0(new_n7060_), .A1(new_n7059_), .B0(new_n7057_), .B1(new_n7055_), .Y(new_n7061_));
  XOR2X1   g06868(.A(new_n7061_), .B(new_n7051_), .Y(new_n7062_));
  INVX1    g06869(.A(new_n6972_), .Y(new_n7063_));
  OR2X1    g06870(.A(new_n6979_), .B(new_n7063_), .Y(new_n7064_));
  OR2X1    g06871(.A(new_n6986_), .B(new_n6980_), .Y(new_n7065_));
  AND2X1   g06872(.A(new_n7065_), .B(new_n7064_), .Y(new_n7066_));
  XOR2X1   g06873(.A(new_n7066_), .B(new_n7062_), .Y(new_n7067_));
  INVX1    g06874(.A(new_n7067_), .Y(new_n7068_));
  OR2X1    g06875(.A(new_n6995_), .B(new_n6993_), .Y(new_n7069_));
  OAI21X1  g06876(.A0(new_n6999_), .A1(new_n6997_), .B0(new_n7069_), .Y(new_n7070_));
  XOR2X1   g06877(.A(new_n7070_), .B(new_n7068_), .Y(new_n7071_));
  NOR2X1   g06878(.A(new_n6989_), .B(new_n6936_), .Y(new_n7072_));
  AOI21X1  g06879(.A0(new_n6987_), .A1(new_n6963_), .B0(new_n7072_), .Y(new_n7073_));
  INVX1    g06880(.A(new_n7073_), .Y(new_n7074_));
  NOR2X1   g06881(.A(new_n6856_), .B(new_n6853_), .Y(new_n7075_));
  AOI21X1  g06882(.A0(new_n6859_), .A1(new_n6857_), .B0(new_n7075_), .Y(new_n7076_));
  XOR2X1   g06883(.A(new_n7076_), .B(new_n7074_), .Y(new_n7077_));
  XOR2X1   g06884(.A(new_n7077_), .B(new_n7071_), .Y(new_n7078_));
  XOR2X1   g06885(.A(new_n7078_), .B(new_n7050_), .Y(new_n7079_));
  INVX1    g06886(.A(new_n7079_), .Y(new_n7080_));
  XOR2X1   g06887(.A(new_n7080_), .B(new_n7015_), .Y(new_n7081_));
  NOR2X1   g06888(.A(new_n7080_), .B(new_n7015_), .Y(new_n7082_));
  AND2X1   g06889(.A(new_n7080_), .B(new_n7015_), .Y(new_n7083_));
  INVX1    g06890(.A(new_n6875_), .Y(new_n7084_));
  AND2X1   g06891(.A(new_n6724_), .B(new_n6721_), .Y(new_n7085_));
  OAI21X1  g06892(.A0(new_n6876_), .A1(new_n7085_), .B0(new_n6895_), .Y(new_n7086_));
  OAI21X1  g06893(.A0(new_n6896_), .A1(new_n7084_), .B0(new_n7086_), .Y(new_n7087_));
  INVX1    g06894(.A(new_n6990_), .Y(new_n7088_));
  OR2X1    g06895(.A(new_n7088_), .B(new_n6907_), .Y(new_n7089_));
  OAI21X1  g06896(.A0(new_n7006_), .A1(new_n6991_), .B0(new_n7089_), .Y(new_n7090_));
  XOR2X1   g06897(.A(new_n7090_), .B(new_n7087_), .Y(new_n7091_));
  AND2X1   g06898(.A(new_n6893_), .B(new_n6889_), .Y(new_n7092_));
  AOI21X1  g06899(.A0(new_n6894_), .A1(new_n6887_), .B0(new_n7092_), .Y(new_n7093_));
  NOR4X1   g06900(.A(new_n5245_), .B(new_n4983_), .C(new_n616_), .D(new_n490_), .Y(new_n7094_));
  AND2X1   g06901(.A(\a[53] ), .B(\a[48] ), .Y(new_n7095_));
  AOI22X1  g06902(.A0(new_n7095_), .A1(\a[14] ), .B0(new_n4035_), .B1(\a[17] ), .Y(new_n7096_));
  NOR3X1   g06903(.A(new_n7096_), .B(new_n7094_), .C(new_n752_), .Y(new_n7097_));
  NOR2X1   g06904(.A(new_n7097_), .B(new_n7094_), .Y(new_n7098_));
  AOI22X1  g06905(.A0(\a[53] ), .A1(\a[14] ), .B0(\a[50] ), .B1(\a[17] ), .Y(new_n7099_));
  INVX1    g06906(.A(new_n7099_), .Y(new_n7100_));
  NOR3X1   g06907(.A(new_n7097_), .B(new_n3926_), .C(new_n752_), .Y(new_n7101_));
  AOI21X1  g06908(.A0(new_n7100_), .A1(new_n7098_), .B0(new_n7101_), .Y(new_n7102_));
  AND2X1   g06909(.A(new_n3607_), .B(new_n1770_), .Y(new_n7103_));
  NOR4X1   g06910(.A(new_n3460_), .B(new_n3096_), .C(new_n1326_), .D(new_n1098_), .Y(new_n7104_));
  NOR2X1   g06911(.A(new_n7104_), .B(new_n7103_), .Y(new_n7105_));
  NOR4X1   g06912(.A(new_n3460_), .B(new_n3081_), .C(new_n1263_), .D(new_n1098_), .Y(new_n7106_));
  NOR2X1   g06913(.A(new_n7106_), .B(new_n7105_), .Y(new_n7107_));
  NOR3X1   g06914(.A(new_n7107_), .B(new_n3096_), .C(new_n1326_), .Y(new_n7108_));
  NOR3X1   g06915(.A(new_n7106_), .B(new_n7104_), .C(new_n7103_), .Y(new_n7109_));
  OAI22X1  g06916(.A0(new_n3460_), .A1(new_n1098_), .B0(new_n3081_), .B1(new_n1263_), .Y(new_n7110_));
  AOI21X1  g06917(.A0(new_n7110_), .A1(new_n7109_), .B0(new_n7108_), .Y(new_n7111_));
  XOR2X1   g06918(.A(new_n7111_), .B(new_n7102_), .Y(new_n7112_));
  AND2X1   g06919(.A(\a[63] ), .B(\a[4] ), .Y(new_n7113_));
  AOI22X1  g06920(.A0(\a[40] ), .A1(\a[27] ), .B0(\a[39] ), .B1(\a[28] ), .Y(new_n7114_));
  INVX1    g06921(.A(new_n7114_), .Y(new_n7115_));
  NAND4X1  g06922(.A(\a[40] ), .B(\a[39] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n7116_));
  NAND3X1  g06923(.A(new_n7115_), .B(new_n7116_), .C(new_n7113_), .Y(new_n7117_));
  AOI22X1  g06924(.A0(new_n7115_), .A1(new_n7113_), .B0(new_n4077_), .B1(new_n1671_), .Y(new_n7118_));
  AOI22X1  g06925(.A0(new_n7118_), .A1(new_n7115_), .B0(new_n7117_), .B1(new_n7113_), .Y(new_n7119_));
  XOR2X1   g06926(.A(new_n7119_), .B(new_n7112_), .Y(new_n7120_));
  INVX1    g06927(.A(new_n7120_), .Y(new_n7121_));
  AOI21X1  g06928(.A0(\a[62] ), .A1(\a[5] ), .B0(\a[34] ), .Y(new_n7122_));
  AND2X1   g06929(.A(\a[49] ), .B(\a[18] ), .Y(new_n7123_));
  INVX1    g06930(.A(new_n7123_), .Y(new_n7124_));
  AND2X1   g06931(.A(new_n2573_), .B(\a[62] ), .Y(new_n7125_));
  NOR3X1   g06932(.A(new_n7124_), .B(new_n7125_), .C(new_n7122_), .Y(new_n7126_));
  INVX1    g06933(.A(new_n7122_), .Y(new_n7127_));
  AOI21X1  g06934(.A0(new_n7123_), .A1(new_n7127_), .B0(new_n7125_), .Y(new_n7128_));
  INVX1    g06935(.A(new_n7128_), .Y(new_n7129_));
  OAI22X1  g06936(.A0(new_n7129_), .A1(new_n7122_), .B0(new_n7126_), .B1(new_n7124_), .Y(new_n7130_));
  NAND4X1  g06937(.A(\a[36] ), .B(\a[34] ), .C(\a[33] ), .D(\a[31] ), .Y(new_n7131_));
  OAI21X1  g06938(.A0(new_n5417_), .A1(new_n2672_), .B0(new_n7131_), .Y(new_n7132_));
  OAI21X1  g06939(.A0(new_n4915_), .A1(new_n2675_), .B0(new_n7132_), .Y(new_n7133_));
  AOI21X1  g06940(.A0(new_n2361_), .A1(new_n2674_), .B0(new_n7132_), .Y(new_n7134_));
  OAI22X1  g06941(.A0(new_n2557_), .A1(new_n2219_), .B0(new_n2028_), .B1(new_n1851_), .Y(new_n7135_));
  AOI22X1  g06942(.A0(new_n7135_), .A1(new_n7134_), .B0(new_n7133_), .B1(new_n2907_), .Y(new_n7136_));
  XOR2X1   g06943(.A(new_n7136_), .B(new_n7130_), .Y(new_n7137_));
  AND2X1   g06944(.A(\a[38] ), .B(\a[29] ), .Y(new_n7138_));
  AOI22X1  g06945(.A0(\a[55] ), .A1(\a[12] ), .B0(\a[54] ), .B1(\a[13] ), .Y(new_n7139_));
  INVX1    g06946(.A(new_n7139_), .Y(new_n7140_));
  NAND4X1  g06947(.A(\a[55] ), .B(\a[54] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n7141_));
  NAND3X1  g06948(.A(new_n7140_), .B(new_n7141_), .C(new_n7138_), .Y(new_n7142_));
  AOI22X1  g06949(.A0(new_n7140_), .A1(new_n7138_), .B0(new_n5240_), .B1(new_n586_), .Y(new_n7143_));
  AOI22X1  g06950(.A0(new_n7143_), .A1(new_n7140_), .B0(new_n7142_), .B1(new_n7138_), .Y(new_n7144_));
  XOR2X1   g06951(.A(new_n7144_), .B(new_n7137_), .Y(new_n7145_));
  AOI22X1  g06952(.A0(\a[59] ), .A1(\a[8] ), .B0(\a[58] ), .B1(\a[9] ), .Y(new_n7146_));
  NAND4X1  g06953(.A(\a[60] ), .B(\a[58] ), .C(\a[9] ), .D(\a[7] ), .Y(new_n7147_));
  NAND4X1  g06954(.A(\a[60] ), .B(\a[59] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n7148_));
  AOI22X1  g06955(.A0(new_n7148_), .A1(new_n7147_), .B0(new_n6121_), .B1(new_n1030_), .Y(new_n7149_));
  AOI21X1  g06956(.A0(new_n6121_), .A1(new_n1030_), .B0(new_n7149_), .Y(new_n7150_));
  INVX1    g06957(.A(new_n7150_), .Y(new_n7151_));
  NAND2X1  g06958(.A(\a[60] ), .B(\a[7] ), .Y(new_n7152_));
  OAI22X1  g06959(.A0(new_n7152_), .A1(new_n7149_), .B0(new_n7151_), .B1(new_n7146_), .Y(new_n7153_));
  NAND4X1  g06960(.A(\a[45] ), .B(\a[43] ), .C(\a[24] ), .D(\a[22] ), .Y(new_n7154_));
  NAND4X1  g06961(.A(\a[45] ), .B(\a[44] ), .C(\a[23] ), .D(\a[22] ), .Y(new_n7155_));
  AOI22X1  g06962(.A0(new_n7155_), .A1(new_n7154_), .B0(new_n4992_), .B1(new_n1219_), .Y(new_n7156_));
  NAND2X1  g06963(.A(\a[45] ), .B(\a[22] ), .Y(new_n7157_));
  NAND4X1  g06964(.A(\a[44] ), .B(\a[43] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n7158_));
  NAND3X1  g06965(.A(new_n7155_), .B(new_n7154_), .C(new_n7158_), .Y(new_n7159_));
  AOI22X1  g06966(.A0(\a[44] ), .A1(\a[23] ), .B0(\a[43] ), .B1(\a[24] ), .Y(new_n7160_));
  OAI22X1  g06967(.A0(new_n7160_), .A1(new_n7159_), .B0(new_n7157_), .B1(new_n7156_), .Y(new_n7161_));
  XOR2X1   g06968(.A(new_n7161_), .B(new_n7153_), .Y(new_n7162_));
  NOR3X1   g06969(.A(new_n3296_), .B(new_n4354_), .C(new_n2345_), .Y(new_n7163_));
  AND2X1   g06970(.A(\a[52] ), .B(\a[51] ), .Y(new_n7164_));
  AND2X1   g06971(.A(new_n7164_), .B(new_n689_), .Y(new_n7165_));
  OR2X1    g06972(.A(new_n7165_), .B(new_n7163_), .Y(new_n7166_));
  NOR4X1   g06973(.A(new_n4349_), .B(new_n2345_), .C(new_n1684_), .D(new_n571_), .Y(new_n7167_));
  INVX1    g06974(.A(new_n7167_), .Y(new_n7168_));
  AND2X1   g06975(.A(new_n7168_), .B(new_n7166_), .Y(new_n7169_));
  AND2X1   g06976(.A(\a[52] ), .B(\a[15] ), .Y(new_n7170_));
  INVX1    g06977(.A(new_n7170_), .Y(new_n7171_));
  AOI22X1  g06978(.A0(\a[51] ), .A1(\a[16] ), .B0(\a[37] ), .B1(\a[30] ), .Y(new_n7172_));
  NOR3X1   g06979(.A(new_n7167_), .B(new_n7165_), .C(new_n7163_), .Y(new_n7173_));
  INVX1    g06980(.A(new_n7173_), .Y(new_n7174_));
  OAI22X1  g06981(.A0(new_n7174_), .A1(new_n7172_), .B0(new_n7171_), .B1(new_n7169_), .Y(new_n7175_));
  INVX1    g06982(.A(new_n7175_), .Y(new_n7176_));
  XOR2X1   g06983(.A(new_n7176_), .B(new_n7162_), .Y(new_n7177_));
  XOR2X1   g06984(.A(new_n7177_), .B(new_n7145_), .Y(new_n7178_));
  XOR2X1   g06985(.A(new_n7178_), .B(new_n7121_), .Y(new_n7179_));
  XOR2X1   g06986(.A(new_n7179_), .B(new_n7093_), .Y(new_n7180_));
  NOR2X1   g06987(.A(new_n6800_), .B(new_n6786_), .Y(new_n7181_));
  AOI21X1  g06988(.A0(new_n6865_), .A1(new_n6765_), .B0(new_n7181_), .Y(new_n7182_));
  AND2X1   g06989(.A(new_n6735_), .B(new_n6697_), .Y(new_n7183_));
  AOI21X1  g06990(.A0(new_n6878_), .A1(new_n6745_), .B0(new_n7183_), .Y(new_n7184_));
  XOR2X1   g06991(.A(new_n7184_), .B(new_n7182_), .Y(new_n7185_));
  NOR2X1   g06992(.A(new_n6862_), .B(new_n6770_), .Y(new_n7186_));
  AOI21X1  g06993(.A0(new_n6863_), .A1(new_n6706_), .B0(new_n7186_), .Y(new_n7187_));
  XOR2X1   g06994(.A(new_n7187_), .B(new_n7185_), .Y(new_n7188_));
  AND2X1   g06995(.A(new_n6869_), .B(new_n6866_), .Y(new_n7189_));
  INVX1    g06996(.A(new_n7189_), .Y(new_n7190_));
  OAI21X1  g06997(.A0(new_n6871_), .A1(new_n6864_), .B0(new_n7190_), .Y(new_n7191_));
  NOR2X1   g06998(.A(new_n6882_), .B(new_n6879_), .Y(new_n7192_));
  AOI21X1  g06999(.A0(new_n6886_), .A1(new_n6883_), .B0(new_n7192_), .Y(new_n7193_));
  XOR2X1   g07000(.A(new_n7193_), .B(new_n7191_), .Y(new_n7194_));
  XOR2X1   g07001(.A(new_n7194_), .B(new_n7188_), .Y(new_n7195_));
  XOR2X1   g07002(.A(new_n7195_), .B(new_n7180_), .Y(new_n7196_));
  NOR2X1   g07003(.A(new_n7196_), .B(new_n7091_), .Y(new_n7197_));
  AND2X1   g07004(.A(new_n7196_), .B(new_n7091_), .Y(new_n7198_));
  NOR4X1   g07005(.A(new_n7198_), .B(new_n7197_), .C(new_n7083_), .D(new_n7082_), .Y(new_n7199_));
  INVX1    g07006(.A(new_n7199_), .Y(new_n7200_));
  NOR3X1   g07007(.A(new_n7198_), .B(new_n7197_), .C(new_n7081_), .Y(new_n7201_));
  AOI21X1  g07008(.A0(new_n7200_), .A1(new_n7081_), .B0(new_n7201_), .Y(new_n7202_));
  XOR2X1   g07009(.A(new_n7202_), .B(new_n7013_), .Y(new_n7203_));
  NOR2X1   g07010(.A(new_n7009_), .B(new_n6835_), .Y(new_n7204_));
  NAND2X1  g07011(.A(new_n7009_), .B(new_n6835_), .Y(new_n7205_));
  AOI21X1  g07012(.A0(new_n7205_), .A1(new_n6832_), .B0(new_n7204_), .Y(new_n7206_));
  XOR2X1   g07013(.A(new_n7206_), .B(new_n7203_), .Y(\asquared[68] ));
  AND2X1   g07014(.A(new_n7090_), .B(new_n7087_), .Y(new_n7208_));
  OR2X1    g07015(.A(new_n7198_), .B(new_n7208_), .Y(new_n7209_));
  AND2X1   g07016(.A(new_n6886_), .B(new_n6883_), .Y(new_n7210_));
  OAI21X1  g07017(.A0(new_n7210_), .A1(new_n7192_), .B0(new_n7191_), .Y(new_n7211_));
  OAI21X1  g07018(.A0(new_n7194_), .A1(new_n7188_), .B0(new_n7211_), .Y(new_n7212_));
  INVX1    g07019(.A(new_n7143_), .Y(new_n7213_));
  XOR2X1   g07020(.A(new_n7109_), .B(new_n7098_), .Y(new_n7214_));
  XOR2X1   g07021(.A(new_n7214_), .B(new_n7213_), .Y(new_n7215_));
  OR2X1    g07022(.A(new_n7111_), .B(new_n7102_), .Y(new_n7216_));
  INVX1    g07023(.A(new_n7112_), .Y(new_n7217_));
  OAI21X1  g07024(.A0(new_n7119_), .A1(new_n7217_), .B0(new_n7216_), .Y(new_n7218_));
  INVX1    g07025(.A(new_n7130_), .Y(new_n7219_));
  OR2X1    g07026(.A(new_n7136_), .B(new_n7219_), .Y(new_n7220_));
  OAI21X1  g07027(.A0(new_n7144_), .A1(new_n7137_), .B0(new_n7220_), .Y(new_n7221_));
  XOR2X1   g07028(.A(new_n7221_), .B(new_n7218_), .Y(new_n7222_));
  XOR2X1   g07029(.A(new_n7222_), .B(new_n7215_), .Y(new_n7223_));
  AND2X1   g07030(.A(new_n7184_), .B(new_n7182_), .Y(new_n7224_));
  OR2X1    g07031(.A(new_n7184_), .B(new_n7182_), .Y(new_n7225_));
  OAI21X1  g07032(.A0(new_n7187_), .A1(new_n7224_), .B0(new_n7225_), .Y(new_n7226_));
  XOR2X1   g07033(.A(new_n7159_), .B(new_n7059_), .Y(new_n7227_));
  XOR2X1   g07034(.A(new_n7227_), .B(new_n7150_), .Y(new_n7228_));
  XOR2X1   g07035(.A(new_n7134_), .B(new_n7118_), .Y(new_n7229_));
  XOR2X1   g07036(.A(new_n7229_), .B(new_n7173_), .Y(new_n7230_));
  XOR2X1   g07037(.A(new_n7230_), .B(new_n7228_), .Y(new_n7231_));
  XOR2X1   g07038(.A(new_n7231_), .B(new_n7226_), .Y(new_n7232_));
  XOR2X1   g07039(.A(new_n7232_), .B(new_n7223_), .Y(new_n7233_));
  XOR2X1   g07040(.A(new_n7233_), .B(new_n7212_), .Y(new_n7234_));
  OR2X1    g07041(.A(new_n7046_), .B(new_n7031_), .Y(new_n7235_));
  OAI21X1  g07042(.A0(new_n7048_), .A1(new_n7021_), .B0(new_n7235_), .Y(new_n7236_));
  INVX1    g07043(.A(new_n7145_), .Y(new_n7237_));
  OR2X1    g07044(.A(new_n7177_), .B(new_n7237_), .Y(new_n7238_));
  OAI21X1  g07045(.A0(new_n7178_), .A1(new_n7120_), .B0(new_n7238_), .Y(new_n7239_));
  NAND3X1  g07046(.A(new_n6970_), .B(new_n6927_), .C(new_n6930_), .Y(new_n7240_));
  AOI21X1  g07047(.A0(new_n6927_), .A1(new_n6930_), .B0(new_n6970_), .Y(new_n7241_));
  AOI21X1  g07048(.A0(new_n7061_), .A1(new_n7240_), .B0(new_n7241_), .Y(new_n7242_));
  AND2X1   g07049(.A(new_n6961_), .B(new_n6942_), .Y(new_n7243_));
  AOI21X1  g07050(.A0(new_n7035_), .A1(new_n6952_), .B0(new_n7243_), .Y(new_n7244_));
  XOR2X1   g07051(.A(new_n7244_), .B(new_n7242_), .Y(new_n7245_));
  AND2X1   g07052(.A(new_n7161_), .B(new_n7153_), .Y(new_n7246_));
  AOI21X1  g07053(.A0(new_n7175_), .A1(new_n7162_), .B0(new_n7246_), .Y(new_n7247_));
  XOR2X1   g07054(.A(new_n7247_), .B(new_n7245_), .Y(new_n7248_));
  NAND2X1  g07055(.A(\a[60] ), .B(\a[8] ), .Y(new_n7249_));
  NAND2X1  g07056(.A(\a[61] ), .B(\a[7] ), .Y(new_n7250_));
  AOI22X1  g07057(.A0(new_n7250_), .A1(new_n7249_), .B0(new_n6428_), .B1(new_n325_), .Y(new_n7251_));
  XOR2X1   g07058(.A(new_n7251_), .B(new_n7128_), .Y(new_n7252_));
  INVX1    g07059(.A(new_n7252_), .Y(new_n7253_));
  OR2X1    g07060(.A(new_n7038_), .B(new_n6985_), .Y(new_n7254_));
  OAI21X1  g07061(.A0(new_n7040_), .A1(new_n6978_), .B0(new_n7254_), .Y(new_n7255_));
  XOR2X1   g07062(.A(new_n7255_), .B(new_n7253_), .Y(new_n7256_));
  AND2X1   g07063(.A(new_n6912_), .B(new_n7032_), .Y(new_n7257_));
  AOI21X1  g07064(.A0(new_n7033_), .A1(new_n6922_), .B0(new_n7257_), .Y(new_n7258_));
  XOR2X1   g07065(.A(new_n7258_), .B(new_n7256_), .Y(new_n7259_));
  XOR2X1   g07066(.A(new_n7259_), .B(new_n7248_), .Y(new_n7260_));
  XOR2X1   g07067(.A(new_n7260_), .B(new_n7239_), .Y(new_n7261_));
  XOR2X1   g07068(.A(new_n7261_), .B(new_n7236_), .Y(new_n7262_));
  INVX1    g07069(.A(new_n7262_), .Y(new_n7263_));
  XOR2X1   g07070(.A(new_n7263_), .B(new_n7234_), .Y(new_n7264_));
  XOR2X1   g07071(.A(new_n7264_), .B(new_n7209_), .Y(new_n7265_));
  AND2X1   g07072(.A(new_n7049_), .B(new_n7017_), .Y(new_n7266_));
  AND2X1   g07073(.A(new_n7078_), .B(new_n7050_), .Y(new_n7267_));
  OR2X1    g07074(.A(new_n7267_), .B(new_n7266_), .Y(new_n7268_));
  NOR2X1   g07075(.A(new_n7179_), .B(new_n7093_), .Y(new_n7269_));
  AOI21X1  g07076(.A0(new_n7195_), .A1(new_n7180_), .B0(new_n7269_), .Y(new_n7270_));
  OR2X1    g07077(.A(new_n7076_), .B(new_n7073_), .Y(new_n7271_));
  OAI21X1  g07078(.A0(new_n7077_), .A1(new_n7071_), .B0(new_n7271_), .Y(new_n7272_));
  NOR2X1   g07079(.A(new_n7042_), .B(new_n7036_), .Y(new_n7273_));
  INVX1    g07080(.A(new_n7273_), .Y(new_n7274_));
  OAI21X1  g07081(.A0(new_n7044_), .A1(new_n7034_), .B0(new_n7274_), .Y(new_n7275_));
  NOR2X1   g07082(.A(new_n7027_), .B(new_n7023_), .Y(new_n7276_));
  INVX1    g07083(.A(new_n7030_), .Y(new_n7277_));
  AOI21X1  g07084(.A0(new_n7277_), .A1(new_n7028_), .B0(new_n7276_), .Y(new_n7278_));
  XOR2X1   g07085(.A(new_n7278_), .B(new_n7275_), .Y(new_n7279_));
  AOI21X1  g07086(.A0(new_n7065_), .A1(new_n7064_), .B0(new_n7062_), .Y(new_n7280_));
  AOI21X1  g07087(.A0(new_n7070_), .A1(new_n7067_), .B0(new_n7280_), .Y(new_n7281_));
  XOR2X1   g07088(.A(new_n7281_), .B(new_n7279_), .Y(new_n7282_));
  NAND4X1  g07089(.A(\a[59] ), .B(\a[57] ), .C(\a[11] ), .D(\a[9] ), .Y(new_n7283_));
  NAND4X1  g07090(.A(\a[59] ), .B(\a[58] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n7284_));
  AOI22X1  g07091(.A0(new_n7284_), .A1(new_n7283_), .B0(new_n6119_), .B1(new_n1002_), .Y(new_n7285_));
  NAND4X1  g07092(.A(\a[58] ), .B(\a[57] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n7286_));
  NAND3X1  g07093(.A(new_n7284_), .B(new_n7283_), .C(new_n7286_), .Y(new_n7287_));
  AOI22X1  g07094(.A0(\a[58] ), .A1(\a[10] ), .B0(\a[57] ), .B1(\a[11] ), .Y(new_n7288_));
  NAND2X1  g07095(.A(\a[59] ), .B(\a[9] ), .Y(new_n7289_));
  OAI22X1  g07096(.A0(new_n7289_), .A1(new_n7285_), .B0(new_n7288_), .B1(new_n7287_), .Y(new_n7290_));
  AOI22X1  g07097(.A0(new_n4404_), .A1(new_n1671_), .B0(new_n2847_), .B1(new_n1484_), .Y(new_n7291_));
  AOI21X1  g07098(.A0(new_n4077_), .A1(new_n1674_), .B0(new_n7291_), .Y(new_n7292_));
  NAND2X1  g07099(.A(\a[41] ), .B(\a[27] ), .Y(new_n7293_));
  AOI22X1  g07100(.A0(\a[40] ), .A1(\a[28] ), .B0(\a[39] ), .B1(\a[29] ), .Y(new_n7294_));
  AOI21X1  g07101(.A0(new_n4077_), .A1(new_n1674_), .B0(new_n7292_), .Y(new_n7295_));
  INVX1    g07102(.A(new_n7295_), .Y(new_n7296_));
  OAI22X1  g07103(.A0(new_n7296_), .A1(new_n7294_), .B0(new_n7293_), .B1(new_n7292_), .Y(new_n7297_));
  XOR2X1   g07104(.A(new_n7297_), .B(new_n7290_), .Y(new_n7298_));
  AND2X1   g07105(.A(\a[47] ), .B(\a[21] ), .Y(new_n7299_));
  INVX1    g07106(.A(new_n7299_), .Y(new_n7300_));
  AOI22X1  g07107(.A0(\a[63] ), .A1(\a[5] ), .B0(\a[62] ), .B1(\a[6] ), .Y(new_n7301_));
  AND2X1   g07108(.A(new_n6789_), .B(new_n295_), .Y(new_n7302_));
  NOR3X1   g07109(.A(new_n7301_), .B(new_n7302_), .C(new_n7300_), .Y(new_n7303_));
  NOR2X1   g07110(.A(new_n7303_), .B(new_n7302_), .Y(new_n7304_));
  INVX1    g07111(.A(new_n7304_), .Y(new_n7305_));
  OAI22X1  g07112(.A0(new_n7305_), .A1(new_n7301_), .B0(new_n7303_), .B1(new_n7300_), .Y(new_n7306_));
  XOR2X1   g07113(.A(new_n7306_), .B(new_n7298_), .Y(new_n7307_));
  INVX1    g07114(.A(new_n7307_), .Y(new_n7308_));
  AOI22X1  g07115(.A0(\a[50] ), .A1(\a[18] ), .B0(\a[49] ), .B1(\a[19] ), .Y(new_n7309_));
  AND2X1   g07116(.A(new_n4321_), .B(new_n855_), .Y(new_n7310_));
  NOR3X1   g07117(.A(new_n7310_), .B(new_n7309_), .C(new_n4914_), .Y(new_n7311_));
  INVX1    g07118(.A(new_n7309_), .Y(new_n7312_));
  AOI21X1  g07119(.A0(new_n7312_), .A1(new_n2120_), .B0(new_n7310_), .Y(new_n7313_));
  INVX1    g07120(.A(new_n7313_), .Y(new_n7314_));
  OAI22X1  g07121(.A0(new_n7314_), .A1(new_n7309_), .B0(new_n7311_), .B1(new_n4914_), .Y(new_n7315_));
  INVX1    g07122(.A(new_n2484_), .Y(new_n7316_));
  INVX1    g07123(.A(new_n3164_), .Y(new_n7317_));
  OAI22X1  g07124(.A0(new_n7317_), .A1(new_n2076_), .B0(new_n7316_), .B1(new_n4923_), .Y(new_n7318_));
  OAI21X1  g07125(.A0(new_n2672_), .A1(new_n6525_), .B0(new_n7318_), .Y(new_n7319_));
  AND2X1   g07126(.A(\a[38] ), .B(\a[30] ), .Y(new_n7320_));
  AOI21X1  g07127(.A0(new_n2671_), .A1(new_n3330_), .B0(new_n7318_), .Y(new_n7321_));
  OAI22X1  g07128(.A0(new_n2345_), .A1(new_n1704_), .B0(new_n2583_), .B1(new_n2219_), .Y(new_n7322_));
  AOI22X1  g07129(.A0(new_n7322_), .A1(new_n7321_), .B0(new_n7320_), .B1(new_n7319_), .Y(new_n7323_));
  XOR2X1   g07130(.A(new_n7323_), .B(new_n7315_), .Y(new_n7324_));
  AND2X1   g07131(.A(\a[56] ), .B(\a[12] ), .Y(new_n7325_));
  AOI22X1  g07132(.A0(new_n7325_), .A1(new_n5794_), .B0(new_n6237_), .B1(new_n586_), .Y(new_n7326_));
  NOR4X1   g07133(.A(new_n4906_), .B(new_n4349_), .C(new_n616_), .D(new_n591_), .Y(new_n7327_));
  OR2X1    g07134(.A(new_n7327_), .B(new_n7326_), .Y(new_n7328_));
  INVX1    g07135(.A(new_n7327_), .Y(new_n7329_));
  AND2X1   g07136(.A(new_n7329_), .B(new_n7326_), .Y(new_n7330_));
  OAI22X1  g07137(.A0(new_n4906_), .A1(new_n591_), .B0(new_n4349_), .B1(new_n616_), .Y(new_n7331_));
  AOI22X1  g07138(.A0(new_n7331_), .A1(new_n7330_), .B0(new_n7328_), .B1(new_n7325_), .Y(new_n7332_));
  XOR2X1   g07139(.A(new_n7332_), .B(new_n7324_), .Y(new_n7333_));
  INVX1    g07140(.A(new_n7333_), .Y(new_n7334_));
  OAI22X1  g07141(.A0(new_n5245_), .A1(new_n549_), .B0(new_n4354_), .B1(new_n571_), .Y(new_n7335_));
  INVX1    g07142(.A(new_n5048_), .Y(new_n7336_));
  AND2X1   g07143(.A(\a[54] ), .B(\a[52] ), .Y(new_n7337_));
  INVX1    g07144(.A(new_n7337_), .Y(new_n7338_));
  OAI22X1  g07145(.A0(new_n7338_), .A1(new_n1025_), .B0(new_n5239_), .B1(new_n867_), .Y(new_n7339_));
  OAI21X1  g07146(.A0(new_n7336_), .A1(new_n1024_), .B0(new_n7339_), .Y(new_n7340_));
  AOI21X1  g07147(.A0(new_n5048_), .A1(new_n689_), .B0(new_n7339_), .Y(new_n7341_));
  AND2X1   g07148(.A(\a[54] ), .B(\a[14] ), .Y(new_n7342_));
  AOI22X1  g07149(.A0(new_n7342_), .A1(new_n7340_), .B0(new_n7341_), .B1(new_n7335_), .Y(new_n7343_));
  AND2X1   g07150(.A(\a[48] ), .B(\a[20] ), .Y(new_n7344_));
  INVX1    g07151(.A(new_n7344_), .Y(new_n7345_));
  AOI22X1  g07152(.A0(\a[46] ), .A1(\a[22] ), .B0(\a[45] ), .B1(\a[23] ), .Y(new_n7346_));
  AND2X1   g07153(.A(new_n3809_), .B(new_n1394_), .Y(new_n7347_));
  NOR3X1   g07154(.A(new_n7347_), .B(new_n7346_), .C(new_n7345_), .Y(new_n7348_));
  NOR2X1   g07155(.A(new_n7348_), .B(new_n7347_), .Y(new_n7349_));
  INVX1    g07156(.A(new_n7349_), .Y(new_n7350_));
  OAI22X1  g07157(.A0(new_n7350_), .A1(new_n7346_), .B0(new_n7348_), .B1(new_n7345_), .Y(new_n7351_));
  XOR2X1   g07158(.A(new_n7351_), .B(new_n7343_), .Y(new_n7352_));
  INVX1    g07159(.A(new_n4992_), .Y(new_n7353_));
  OAI22X1  g07160(.A0(new_n7353_), .A1(new_n1772_), .B0(new_n3212_), .B1(new_n1651_), .Y(new_n7354_));
  OAI21X1  g07161(.A0(new_n6502_), .A1(new_n1771_), .B0(new_n7354_), .Y(new_n7355_));
  AND2X1   g07162(.A(\a[44] ), .B(\a[24] ), .Y(new_n7356_));
  AOI21X1  g07163(.A0(new_n3462_), .A1(new_n1770_), .B0(new_n7354_), .Y(new_n7357_));
  OAI22X1  g07164(.A0(new_n3037_), .A1(new_n1326_), .B0(new_n3096_), .B1(new_n1263_), .Y(new_n7358_));
  AOI22X1  g07165(.A0(new_n7358_), .A1(new_n7357_), .B0(new_n7356_), .B1(new_n7355_), .Y(new_n7359_));
  XOR2X1   g07166(.A(new_n7359_), .B(new_n7352_), .Y(new_n7360_));
  XOR2X1   g07167(.A(new_n7360_), .B(new_n7334_), .Y(new_n7361_));
  XOR2X1   g07168(.A(new_n7361_), .B(new_n7308_), .Y(new_n7362_));
  XOR2X1   g07169(.A(new_n7362_), .B(new_n7282_), .Y(new_n7363_));
  INVX1    g07170(.A(new_n7363_), .Y(new_n7364_));
  XOR2X1   g07171(.A(new_n7364_), .B(new_n7272_), .Y(new_n7365_));
  XOR2X1   g07172(.A(new_n7365_), .B(new_n7270_), .Y(new_n7366_));
  XOR2X1   g07173(.A(new_n7366_), .B(new_n7268_), .Y(new_n7367_));
  XOR2X1   g07174(.A(new_n7367_), .B(new_n7265_), .Y(new_n7368_));
  NOR2X1   g07175(.A(new_n7199_), .B(new_n7082_), .Y(new_n7369_));
  XOR2X1   g07176(.A(new_n7369_), .B(new_n7368_), .Y(new_n7370_));
  INVX1    g07177(.A(new_n7202_), .Y(new_n7371_));
  NAND2X1  g07178(.A(new_n7371_), .B(new_n7013_), .Y(new_n7372_));
  NOR2X1   g07179(.A(new_n7371_), .B(new_n7013_), .Y(new_n7373_));
  OAI21X1  g07180(.A0(new_n7206_), .A1(new_n7373_), .B0(new_n7372_), .Y(new_n7374_));
  XOR2X1   g07181(.A(new_n7374_), .B(new_n7370_), .Y(\asquared[69] ));
  NOR2X1   g07182(.A(new_n7365_), .B(new_n7270_), .Y(new_n7376_));
  AOI21X1  g07183(.A0(new_n7366_), .A1(new_n7268_), .B0(new_n7376_), .Y(new_n7377_));
  INVX1    g07184(.A(new_n7377_), .Y(new_n7378_));
  AND2X1   g07185(.A(new_n7232_), .B(new_n7223_), .Y(new_n7379_));
  AOI21X1  g07186(.A0(new_n7233_), .A1(new_n7212_), .B0(new_n7379_), .Y(new_n7380_));
  NOR2X1   g07187(.A(new_n7361_), .B(new_n7308_), .Y(new_n7381_));
  AOI21X1  g07188(.A0(new_n7360_), .A1(new_n7333_), .B0(new_n7381_), .Y(new_n7382_));
  NOR2X1   g07189(.A(new_n7230_), .B(new_n7228_), .Y(new_n7383_));
  AOI21X1  g07190(.A0(new_n7231_), .A1(new_n7226_), .B0(new_n7383_), .Y(new_n7384_));
  XOR2X1   g07191(.A(new_n7357_), .B(new_n7330_), .Y(new_n7385_));
  XOR2X1   g07192(.A(new_n7385_), .B(new_n7295_), .Y(new_n7386_));
  NOR2X1   g07193(.A(new_n7134_), .B(new_n7118_), .Y(new_n7387_));
  AOI21X1  g07194(.A0(new_n7229_), .A1(new_n7174_), .B0(new_n7387_), .Y(new_n7388_));
  NOR2X1   g07195(.A(new_n7109_), .B(new_n7098_), .Y(new_n7389_));
  AOI21X1  g07196(.A0(new_n7214_), .A1(new_n7213_), .B0(new_n7389_), .Y(new_n7390_));
  XOR2X1   g07197(.A(new_n7390_), .B(new_n7388_), .Y(new_n7391_));
  XOR2X1   g07198(.A(new_n7391_), .B(new_n7386_), .Y(new_n7392_));
  XOR2X1   g07199(.A(new_n7392_), .B(new_n7384_), .Y(new_n7393_));
  XOR2X1   g07200(.A(new_n7393_), .B(new_n7382_), .Y(new_n7394_));
  XOR2X1   g07201(.A(new_n7394_), .B(new_n7380_), .Y(new_n7395_));
  AND2X1   g07202(.A(new_n7277_), .B(new_n7028_), .Y(new_n7396_));
  OAI21X1  g07203(.A0(new_n7396_), .A1(new_n7276_), .B0(new_n7275_), .Y(new_n7397_));
  OAI21X1  g07204(.A0(new_n7281_), .A1(new_n7279_), .B0(new_n7397_), .Y(new_n7398_));
  INVX1    g07205(.A(new_n7315_), .Y(new_n7399_));
  OR2X1    g07206(.A(new_n7323_), .B(new_n7399_), .Y(new_n7400_));
  OAI21X1  g07207(.A0(new_n7332_), .A1(new_n7324_), .B0(new_n7400_), .Y(new_n7401_));
  INVX1    g07208(.A(new_n7351_), .Y(new_n7402_));
  OR2X1    g07209(.A(new_n7402_), .B(new_n7343_), .Y(new_n7403_));
  OAI21X1  g07210(.A0(new_n7359_), .A1(new_n7352_), .B0(new_n7403_), .Y(new_n7404_));
  XOR2X1   g07211(.A(new_n7404_), .B(new_n7401_), .Y(new_n7405_));
  NOR2X1   g07212(.A(new_n7255_), .B(new_n7253_), .Y(new_n7406_));
  NAND2X1  g07213(.A(new_n7255_), .B(new_n7253_), .Y(new_n7407_));
  OAI21X1  g07214(.A0(new_n7258_), .A1(new_n7406_), .B0(new_n7407_), .Y(new_n7408_));
  XOR2X1   g07215(.A(new_n7408_), .B(new_n7405_), .Y(new_n7409_));
  XOR2X1   g07216(.A(new_n7305_), .B(new_n7287_), .Y(new_n7410_));
  XOR2X1   g07217(.A(new_n7410_), .B(new_n7350_), .Y(new_n7411_));
  XOR2X1   g07218(.A(new_n7321_), .B(new_n7313_), .Y(new_n7412_));
  XOR2X1   g07219(.A(new_n7412_), .B(new_n7341_), .Y(new_n7413_));
  AND2X1   g07220(.A(new_n7297_), .B(new_n7290_), .Y(new_n7414_));
  AOI21X1  g07221(.A0(new_n7306_), .A1(new_n7298_), .B0(new_n7414_), .Y(new_n7415_));
  XOR2X1   g07222(.A(new_n7415_), .B(new_n7413_), .Y(new_n7416_));
  XOR2X1   g07223(.A(new_n7416_), .B(new_n7411_), .Y(new_n7417_));
  XOR2X1   g07224(.A(new_n7417_), .B(new_n7409_), .Y(new_n7418_));
  XOR2X1   g07225(.A(new_n7418_), .B(new_n7398_), .Y(new_n7419_));
  XOR2X1   g07226(.A(new_n7419_), .B(new_n7395_), .Y(new_n7420_));
  XOR2X1   g07227(.A(new_n7420_), .B(new_n7378_), .Y(new_n7421_));
  AND2X1   g07228(.A(new_n7261_), .B(new_n7236_), .Y(new_n7422_));
  AOI21X1  g07229(.A0(new_n7262_), .A1(new_n7234_), .B0(new_n7422_), .Y(new_n7423_));
  AND2X1   g07230(.A(new_n7362_), .B(new_n7282_), .Y(new_n7424_));
  AOI21X1  g07231(.A0(new_n7363_), .A1(new_n7272_), .B0(new_n7424_), .Y(new_n7425_));
  XOR2X1   g07232(.A(new_n7425_), .B(new_n7423_), .Y(new_n7426_));
  NAND4X1  g07233(.A(\a[52] ), .B(\a[50] ), .C(\a[19] ), .D(\a[17] ), .Y(new_n7427_));
  NAND4X1  g07234(.A(\a[51] ), .B(\a[50] ), .C(\a[19] ), .D(\a[18] ), .Y(new_n7428_));
  AOI22X1  g07235(.A0(new_n7428_), .A1(new_n7427_), .B0(new_n7164_), .B1(new_n796_), .Y(new_n7429_));
  NAND4X1  g07236(.A(\a[52] ), .B(\a[51] ), .C(\a[18] ), .D(\a[17] ), .Y(new_n7430_));
  NAND3X1  g07237(.A(new_n7428_), .B(new_n7427_), .C(new_n7430_), .Y(new_n7431_));
  AOI22X1  g07238(.A0(\a[52] ), .A1(\a[17] ), .B0(\a[51] ), .B1(\a[18] ), .Y(new_n7432_));
  NAND2X1  g07239(.A(\a[50] ), .B(\a[19] ), .Y(new_n7433_));
  OAI22X1  g07240(.A0(new_n7433_), .A1(new_n7429_), .B0(new_n7432_), .B1(new_n7431_), .Y(new_n7434_));
  NAND4X1  g07241(.A(\a[41] ), .B(\a[39] ), .C(\a[30] ), .D(\a[28] ), .Y(new_n7435_));
  NAND4X1  g07242(.A(\a[41] ), .B(\a[40] ), .C(\a[29] ), .D(\a[28] ), .Y(new_n7436_));
  AOI22X1  g07243(.A0(new_n7436_), .A1(new_n7435_), .B0(new_n4077_), .B1(new_n2196_), .Y(new_n7437_));
  NAND2X1  g07244(.A(\a[41] ), .B(\a[28] ), .Y(new_n7438_));
  NAND4X1  g07245(.A(\a[40] ), .B(\a[39] ), .C(\a[30] ), .D(\a[29] ), .Y(new_n7439_));
  NAND3X1  g07246(.A(new_n7436_), .B(new_n7435_), .C(new_n7439_), .Y(new_n7440_));
  AOI22X1  g07247(.A0(\a[40] ), .A1(\a[29] ), .B0(\a[39] ), .B1(\a[30] ), .Y(new_n7441_));
  OAI22X1  g07248(.A0(new_n7441_), .A1(new_n7440_), .B0(new_n7438_), .B1(new_n7437_), .Y(new_n7442_));
  XOR2X1   g07249(.A(new_n7442_), .B(new_n7434_), .Y(new_n7443_));
  AND2X1   g07250(.A(new_n7159_), .B(new_n7059_), .Y(new_n7444_));
  AOI21X1  g07251(.A0(new_n7227_), .A1(new_n7151_), .B0(new_n7444_), .Y(new_n7445_));
  XOR2X1   g07252(.A(new_n7445_), .B(new_n7443_), .Y(new_n7446_));
  AND2X1   g07253(.A(\a[35] ), .B(\a[7] ), .Y(new_n7447_));
  AOI21X1  g07254(.A0(new_n7447_), .A1(\a[62] ), .B0(new_n2361_), .Y(new_n7448_));
  INVX1    g07255(.A(new_n7448_), .Y(new_n7449_));
  AOI21X1  g07256(.A0(\a[62] ), .A1(\a[7] ), .B0(\a[35] ), .Y(new_n7450_));
  NAND4X1  g07257(.A(\a[62] ), .B(\a[35] ), .C(\a[34] ), .D(\a[7] ), .Y(new_n7451_));
  OAI21X1  g07258(.A0(new_n7450_), .A1(new_n7449_), .B0(new_n7451_), .Y(new_n7452_));
  NAND4X1  g07259(.A(\a[38] ), .B(\a[36] ), .C(\a[33] ), .D(\a[31] ), .Y(new_n7453_));
  NAND4X1  g07260(.A(\a[38] ), .B(\a[37] ), .C(\a[32] ), .D(\a[31] ), .Y(new_n7454_));
  AOI22X1  g07261(.A0(new_n7454_), .A1(new_n7453_), .B0(new_n3330_), .B1(new_n2674_), .Y(new_n7455_));
  NAND2X1  g07262(.A(\a[38] ), .B(\a[31] ), .Y(new_n7456_));
  AOI21X1  g07263(.A0(new_n3330_), .A1(new_n2674_), .B0(new_n7455_), .Y(new_n7457_));
  INVX1    g07264(.A(new_n7457_), .Y(new_n7458_));
  AOI22X1  g07265(.A0(\a[37] ), .A1(\a[32] ), .B0(\a[36] ), .B1(\a[33] ), .Y(new_n7459_));
  OAI22X1  g07266(.A0(new_n7459_), .A1(new_n7458_), .B0(new_n7456_), .B1(new_n7455_), .Y(new_n7460_));
  XOR2X1   g07267(.A(new_n7460_), .B(new_n7452_), .Y(new_n7461_));
  AND2X1   g07268(.A(\a[49] ), .B(\a[15] ), .Y(new_n7462_));
  AND2X1   g07269(.A(\a[54] ), .B(\a[20] ), .Y(new_n7463_));
  AOI22X1  g07270(.A0(new_n7463_), .A1(new_n7462_), .B0(new_n5238_), .B1(new_n689_), .Y(new_n7464_));
  NOR4X1   g07271(.A(new_n5245_), .B(new_n3915_), .C(new_n934_), .D(new_n571_), .Y(new_n7465_));
  OR2X1    g07272(.A(new_n7465_), .B(new_n7464_), .Y(new_n7466_));
  AND2X1   g07273(.A(\a[54] ), .B(\a[15] ), .Y(new_n7467_));
  INVX1    g07274(.A(new_n7465_), .Y(new_n7468_));
  AND2X1   g07275(.A(new_n7468_), .B(new_n7464_), .Y(new_n7469_));
  OAI22X1  g07276(.A0(new_n5245_), .A1(new_n571_), .B0(new_n3915_), .B1(new_n934_), .Y(new_n7470_));
  AOI22X1  g07277(.A0(new_n7470_), .A1(new_n7469_), .B0(new_n7467_), .B1(new_n7466_), .Y(new_n7471_));
  XOR2X1   g07278(.A(new_n7471_), .B(new_n7461_), .Y(new_n7472_));
  NAND2X1  g07279(.A(new_n7472_), .B(new_n7446_), .Y(new_n7473_));
  AND2X1   g07280(.A(new_n7221_), .B(new_n7218_), .Y(new_n7474_));
  AOI21X1  g07281(.A0(new_n7222_), .A1(new_n7215_), .B0(new_n7474_), .Y(new_n7475_));
  XOR2X1   g07282(.A(new_n7472_), .B(new_n7446_), .Y(new_n7476_));
  NOR2X1   g07283(.A(new_n7476_), .B(new_n7475_), .Y(new_n7477_));
  INVX1    g07284(.A(new_n7475_), .Y(new_n7478_));
  NOR2X1   g07285(.A(new_n7472_), .B(new_n7446_), .Y(new_n7479_));
  AOI21X1  g07286(.A0(new_n7473_), .A1(new_n7478_), .B0(new_n7479_), .Y(new_n7480_));
  AOI21X1  g07287(.A0(new_n7480_), .A1(new_n7473_), .B0(new_n7477_), .Y(new_n7481_));
  NOR2X1   g07288(.A(new_n7259_), .B(new_n7248_), .Y(new_n7482_));
  AOI21X1  g07289(.A0(new_n7260_), .A1(new_n7239_), .B0(new_n7482_), .Y(new_n7483_));
  XOR2X1   g07290(.A(new_n7483_), .B(new_n7481_), .Y(new_n7484_));
  NAND4X1  g07291(.A(\a[61] ), .B(\a[59] ), .C(\a[10] ), .D(\a[8] ), .Y(new_n7485_));
  NAND4X1  g07292(.A(\a[61] ), .B(\a[60] ), .C(\a[9] ), .D(\a[8] ), .Y(new_n7486_));
  AOI22X1  g07293(.A0(new_n7486_), .A1(new_n7485_), .B0(new_n6427_), .B1(new_n881_), .Y(new_n7487_));
  NAND4X1  g07294(.A(\a[60] ), .B(\a[59] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n7488_));
  NAND3X1  g07295(.A(new_n7486_), .B(new_n7485_), .C(new_n7488_), .Y(new_n7489_));
  AOI22X1  g07296(.A0(\a[60] ), .A1(\a[9] ), .B0(\a[59] ), .B1(\a[10] ), .Y(new_n7490_));
  NAND2X1  g07297(.A(\a[61] ), .B(\a[8] ), .Y(new_n7491_));
  OAI22X1  g07298(.A0(new_n7491_), .A1(new_n7487_), .B0(new_n7490_), .B1(new_n7489_), .Y(new_n7492_));
  NAND4X1  g07299(.A(\a[46] ), .B(\a[44] ), .C(\a[25] ), .D(\a[23] ), .Y(new_n7493_));
  NAND4X1  g07300(.A(\a[46] ), .B(\a[45] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n7494_));
  AOI22X1  g07301(.A0(new_n7494_), .A1(new_n7493_), .B0(new_n3918_), .B1(new_n1532_), .Y(new_n7495_));
  NAND2X1  g07302(.A(\a[46] ), .B(\a[23] ), .Y(new_n7496_));
  AOI22X1  g07303(.A0(\a[45] ), .A1(\a[24] ), .B0(\a[44] ), .B1(\a[25] ), .Y(new_n7497_));
  AOI21X1  g07304(.A0(new_n3918_), .A1(new_n1532_), .B0(new_n7495_), .Y(new_n7498_));
  INVX1    g07305(.A(new_n7498_), .Y(new_n7499_));
  OAI22X1  g07306(.A0(new_n7499_), .A1(new_n7497_), .B0(new_n7496_), .B1(new_n7495_), .Y(new_n7500_));
  XOR2X1   g07307(.A(new_n7500_), .B(new_n7492_), .Y(new_n7501_));
  NAND2X1  g07308(.A(\a[63] ), .B(\a[6] ), .Y(new_n7502_));
  AOI22X1  g07309(.A0(\a[43] ), .A1(\a[26] ), .B0(\a[42] ), .B1(\a[27] ), .Y(new_n7503_));
  AND2X1   g07310(.A(new_n3462_), .B(new_n1995_), .Y(new_n7504_));
  NOR3X1   g07311(.A(new_n7503_), .B(new_n7504_), .C(new_n7502_), .Y(new_n7505_));
  OAI22X1  g07312(.A0(new_n7503_), .A1(new_n7502_), .B0(new_n6502_), .B1(new_n3483_), .Y(new_n7506_));
  OAI22X1  g07313(.A0(new_n7506_), .A1(new_n7503_), .B0(new_n7505_), .B1(new_n7502_), .Y(new_n7507_));
  XOR2X1   g07314(.A(new_n7507_), .B(new_n7501_), .Y(new_n7508_));
  AND2X1   g07315(.A(new_n7244_), .B(new_n7242_), .Y(new_n7509_));
  OR2X1    g07316(.A(new_n7244_), .B(new_n7242_), .Y(new_n7510_));
  OAI21X1  g07317(.A0(new_n7247_), .A1(new_n7509_), .B0(new_n7510_), .Y(new_n7511_));
  XOR2X1   g07318(.A(new_n7511_), .B(new_n7508_), .Y(new_n7512_));
  NAND4X1  g07319(.A(\a[58] ), .B(\a[56] ), .C(\a[13] ), .D(\a[11] ), .Y(new_n7513_));
  NAND4X1  g07320(.A(\a[58] ), .B(\a[57] ), .C(\a[12] ), .D(\a[11] ), .Y(new_n7514_));
  AOI22X1  g07321(.A0(new_n7514_), .A1(new_n7513_), .B0(new_n5554_), .B1(new_n586_), .Y(new_n7515_));
  AND2X1   g07322(.A(\a[58] ), .B(\a[11] ), .Y(new_n7516_));
  INVX1    g07323(.A(new_n7516_), .Y(new_n7517_));
  AOI21X1  g07324(.A0(new_n5554_), .A1(new_n586_), .B0(new_n7515_), .Y(new_n7518_));
  INVX1    g07325(.A(new_n7518_), .Y(new_n7519_));
  AOI22X1  g07326(.A0(\a[57] ), .A1(\a[12] ), .B0(\a[56] ), .B1(\a[13] ), .Y(new_n7520_));
  OAI22X1  g07327(.A0(new_n7520_), .A1(new_n7519_), .B0(new_n7517_), .B1(new_n7515_), .Y(new_n7521_));
  AOI22X1  g07328(.A0(new_n7251_), .A1(new_n7129_), .B0(new_n6428_), .B1(new_n325_), .Y(new_n7522_));
  XOR2X1   g07329(.A(new_n7522_), .B(new_n7521_), .Y(new_n7523_));
  AND2X1   g07330(.A(\a[55] ), .B(\a[14] ), .Y(new_n7524_));
  AOI22X1  g07331(.A0(\a[48] ), .A1(\a[21] ), .B0(\a[47] ), .B1(\a[22] ), .Y(new_n7525_));
  INVX1    g07332(.A(new_n7525_), .Y(new_n7526_));
  NAND4X1  g07333(.A(\a[48] ), .B(\a[47] ), .C(\a[22] ), .D(\a[21] ), .Y(new_n7527_));
  NAND3X1  g07334(.A(new_n7526_), .B(new_n7527_), .C(new_n7524_), .Y(new_n7528_));
  AOI22X1  g07335(.A0(new_n7526_), .A1(new_n7524_), .B0(new_n4272_), .B1(new_n1154_), .Y(new_n7529_));
  AOI22X1  g07336(.A0(new_n7529_), .A1(new_n7526_), .B0(new_n7528_), .B1(new_n7524_), .Y(new_n7530_));
  XOR2X1   g07337(.A(new_n7530_), .B(new_n7523_), .Y(new_n7531_));
  XOR2X1   g07338(.A(new_n7531_), .B(new_n7512_), .Y(new_n7532_));
  XOR2X1   g07339(.A(new_n7532_), .B(new_n7484_), .Y(new_n7533_));
  XOR2X1   g07340(.A(new_n7533_), .B(new_n7426_), .Y(new_n7534_));
  XOR2X1   g07341(.A(new_n7534_), .B(new_n7421_), .Y(new_n7535_));
  AOI21X1  g07342(.A0(new_n7196_), .A1(new_n7091_), .B0(new_n7208_), .Y(new_n7536_));
  NOR2X1   g07343(.A(new_n7264_), .B(new_n7536_), .Y(new_n7537_));
  INVX1    g07344(.A(new_n7265_), .Y(new_n7538_));
  AOI21X1  g07345(.A0(new_n7367_), .A1(new_n7538_), .B0(new_n7537_), .Y(new_n7539_));
  XOR2X1   g07346(.A(new_n7539_), .B(new_n7535_), .Y(new_n7540_));
  AND2X1   g07347(.A(new_n7369_), .B(new_n7368_), .Y(new_n7541_));
  INVX1    g07348(.A(new_n7541_), .Y(new_n7542_));
  NOR2X1   g07349(.A(new_n7369_), .B(new_n7368_), .Y(new_n7543_));
  AOI21X1  g07350(.A0(new_n7374_), .A1(new_n7542_), .B0(new_n7543_), .Y(new_n7544_));
  XOR2X1   g07351(.A(new_n7544_), .B(new_n7540_), .Y(\asquared[70] ));
  AND2X1   g07352(.A(new_n7420_), .B(new_n7378_), .Y(new_n7546_));
  AND2X1   g07353(.A(new_n7534_), .B(new_n7421_), .Y(new_n7547_));
  OR2X1    g07354(.A(new_n7547_), .B(new_n7546_), .Y(new_n7548_));
  NOR2X1   g07355(.A(new_n7425_), .B(new_n7423_), .Y(new_n7549_));
  AOI21X1  g07356(.A0(new_n7533_), .A1(new_n7426_), .B0(new_n7549_), .Y(new_n7550_));
  AND2X1   g07357(.A(new_n7417_), .B(new_n7409_), .Y(new_n7551_));
  AOI21X1  g07358(.A0(new_n7418_), .A1(new_n7398_), .B0(new_n7551_), .Y(new_n7552_));
  AND2X1   g07359(.A(new_n7511_), .B(new_n7508_), .Y(new_n7553_));
  AOI21X1  g07360(.A0(new_n7531_), .A1(new_n7512_), .B0(new_n7553_), .Y(new_n7554_));
  AND2X1   g07361(.A(new_n7404_), .B(new_n7401_), .Y(new_n7555_));
  AOI21X1  g07362(.A0(new_n7408_), .A1(new_n7405_), .B0(new_n7555_), .Y(new_n7556_));
  INVX1    g07363(.A(new_n7529_), .Y(new_n7557_));
  XOR2X1   g07364(.A(new_n7519_), .B(new_n7489_), .Y(new_n7558_));
  XOR2X1   g07365(.A(new_n7558_), .B(new_n7557_), .Y(new_n7559_));
  AND2X1   g07366(.A(new_n7305_), .B(new_n7287_), .Y(new_n7560_));
  AOI21X1  g07367(.A0(new_n7410_), .A1(new_n7350_), .B0(new_n7560_), .Y(new_n7561_));
  NOR2X1   g07368(.A(new_n7357_), .B(new_n7330_), .Y(new_n7562_));
  AOI21X1  g07369(.A0(new_n7385_), .A1(new_n7296_), .B0(new_n7562_), .Y(new_n7563_));
  XOR2X1   g07370(.A(new_n7563_), .B(new_n7561_), .Y(new_n7564_));
  XOR2X1   g07371(.A(new_n7564_), .B(new_n7559_), .Y(new_n7565_));
  XOR2X1   g07372(.A(new_n7565_), .B(new_n7556_), .Y(new_n7566_));
  XOR2X1   g07373(.A(new_n7566_), .B(new_n7554_), .Y(new_n7567_));
  XOR2X1   g07374(.A(new_n7567_), .B(new_n7552_), .Y(new_n7568_));
  INVX1    g07375(.A(new_n7568_), .Y(new_n7569_));
  NOR2X1   g07376(.A(new_n7483_), .B(new_n7481_), .Y(new_n7570_));
  AOI21X1  g07377(.A0(new_n7532_), .A1(new_n7484_), .B0(new_n7570_), .Y(new_n7571_));
  XOR2X1   g07378(.A(new_n7571_), .B(new_n7569_), .Y(new_n7572_));
  NOR2X1   g07379(.A(new_n7550_), .B(new_n7572_), .Y(new_n7573_));
  OR2X1    g07380(.A(new_n7573_), .B(new_n7550_), .Y(new_n7574_));
  NAND2X1  g07381(.A(new_n7419_), .B(new_n7395_), .Y(new_n7575_));
  OAI21X1  g07382(.A0(new_n7394_), .A1(new_n7380_), .B0(new_n7575_), .Y(new_n7576_));
  XOR2X1   g07383(.A(new_n7506_), .B(new_n7440_), .Y(new_n7577_));
  XOR2X1   g07384(.A(new_n7577_), .B(new_n7499_), .Y(new_n7578_));
  AOI21X1  g07385(.A0(\a[62] ), .A1(\a[8] ), .B0(new_n7449_), .Y(new_n7579_));
  NOR3X1   g07386(.A(new_n7448_), .B(new_n6606_), .C(new_n413_), .Y(new_n7580_));
  NOR3X1   g07387(.A(new_n7579_), .B(new_n7580_), .C(new_n7457_), .Y(new_n7581_));
  NOR2X1   g07388(.A(new_n7581_), .B(new_n7580_), .Y(new_n7582_));
  INVX1    g07389(.A(new_n7582_), .Y(new_n7583_));
  OAI22X1  g07390(.A0(new_n7583_), .A1(new_n7579_), .B0(new_n7581_), .B1(new_n7457_), .Y(new_n7584_));
  XOR2X1   g07391(.A(new_n7584_), .B(new_n7578_), .Y(new_n7585_));
  INVX1    g07392(.A(new_n7585_), .Y(new_n7586_));
  NAND2X1  g07393(.A(new_n7442_), .B(new_n7434_), .Y(new_n7587_));
  INVX1    g07394(.A(new_n7443_), .Y(new_n7588_));
  OAI21X1  g07395(.A0(new_n7445_), .A1(new_n7588_), .B0(new_n7587_), .Y(new_n7589_));
  XOR2X1   g07396(.A(new_n7589_), .B(new_n7586_), .Y(new_n7590_));
  AND2X1   g07397(.A(new_n7500_), .B(new_n7492_), .Y(new_n7591_));
  AOI21X1  g07398(.A0(new_n7507_), .A1(new_n7501_), .B0(new_n7591_), .Y(new_n7592_));
  INVX1    g07399(.A(new_n7521_), .Y(new_n7593_));
  OR2X1    g07400(.A(new_n7530_), .B(new_n7523_), .Y(new_n7594_));
  OAI21X1  g07401(.A0(new_n7522_), .A1(new_n7593_), .B0(new_n7594_), .Y(new_n7595_));
  XOR2X1   g07402(.A(new_n7595_), .B(new_n7592_), .Y(new_n7596_));
  AND2X1   g07403(.A(new_n7460_), .B(new_n7452_), .Y(new_n7597_));
  INVX1    g07404(.A(new_n7597_), .Y(new_n7598_));
  INVX1    g07405(.A(new_n7461_), .Y(new_n7599_));
  OAI21X1  g07406(.A0(new_n7471_), .A1(new_n7599_), .B0(new_n7598_), .Y(new_n7600_));
  INVX1    g07407(.A(new_n7600_), .Y(new_n7601_));
  XOR2X1   g07408(.A(new_n7601_), .B(new_n7596_), .Y(new_n7602_));
  XOR2X1   g07409(.A(new_n7602_), .B(new_n7480_), .Y(new_n7603_));
  XOR2X1   g07410(.A(new_n7603_), .B(new_n7590_), .Y(new_n7604_));
  XOR2X1   g07411(.A(new_n7604_), .B(new_n7576_), .Y(new_n7605_));
  NOR2X1   g07412(.A(new_n7415_), .B(new_n7413_), .Y(new_n7606_));
  AOI21X1  g07413(.A0(new_n7416_), .A1(new_n7411_), .B0(new_n7606_), .Y(new_n7607_));
  AOI22X1  g07414(.A0(\a[63] ), .A1(\a[7] ), .B0(\a[47] ), .B1(\a[23] ), .Y(new_n7608_));
  AND2X1   g07415(.A(\a[42] ), .B(\a[28] ), .Y(new_n7609_));
  INVX1    g07416(.A(new_n7609_), .Y(new_n7610_));
  NOR4X1   g07417(.A(new_n6549_), .B(new_n4041_), .C(new_n1216_), .D(new_n532_), .Y(new_n7611_));
  NOR3X1   g07418(.A(new_n7610_), .B(new_n7611_), .C(new_n7608_), .Y(new_n7612_));
  INVX1    g07419(.A(new_n7608_), .Y(new_n7613_));
  AOI21X1  g07420(.A0(new_n7609_), .A1(new_n7613_), .B0(new_n7611_), .Y(new_n7614_));
  INVX1    g07421(.A(new_n7614_), .Y(new_n7615_));
  OAI22X1  g07422(.A0(new_n7615_), .A1(new_n7608_), .B0(new_n7612_), .B1(new_n7610_), .Y(new_n7616_));
  INVX1    g07423(.A(new_n2847_), .Y(new_n7617_));
  INVX1    g07424(.A(new_n4404_), .Y(new_n7618_));
  OAI22X1  g07425(.A0(new_n7618_), .A1(new_n2197_), .B0(new_n7617_), .B1(new_n2430_), .Y(new_n7619_));
  OAI21X1  g07426(.A0(new_n6180_), .A1(new_n2076_), .B0(new_n7619_), .Y(new_n7620_));
  AND2X1   g07427(.A(\a[41] ), .B(\a[29] ), .Y(new_n7621_));
  AOI21X1  g07428(.A0(new_n4077_), .A1(new_n2075_), .B0(new_n7619_), .Y(new_n7622_));
  OAI22X1  g07429(.A0(new_n3036_), .A1(new_n1684_), .B0(new_n2652_), .B1(new_n1704_), .Y(new_n7623_));
  AOI22X1  g07430(.A0(new_n7623_), .A1(new_n7622_), .B0(new_n7621_), .B1(new_n7620_), .Y(new_n7624_));
  XOR2X1   g07431(.A(new_n7624_), .B(new_n7616_), .Y(new_n7625_));
  INVX1    g07432(.A(new_n7341_), .Y(new_n7626_));
  NOR2X1   g07433(.A(new_n7321_), .B(new_n7313_), .Y(new_n7627_));
  AOI21X1  g07434(.A0(new_n7412_), .A1(new_n7626_), .B0(new_n7627_), .Y(new_n7628_));
  XOR2X1   g07435(.A(new_n7628_), .B(new_n7625_), .Y(new_n7629_));
  INVX1    g07436(.A(new_n7629_), .Y(new_n7630_));
  AOI22X1  g07437(.A0(\a[56] ), .A1(\a[14] ), .B0(\a[55] ), .B1(\a[15] ), .Y(new_n7631_));
  AND2X1   g07438(.A(\a[48] ), .B(\a[22] ), .Y(new_n7632_));
  INVX1    g07439(.A(new_n7632_), .Y(new_n7633_));
  AND2X1   g07440(.A(new_n6237_), .B(new_n691_), .Y(new_n7634_));
  NOR3X1   g07441(.A(new_n7633_), .B(new_n7634_), .C(new_n7631_), .Y(new_n7635_));
  INVX1    g07442(.A(new_n7631_), .Y(new_n7636_));
  AOI21X1  g07443(.A0(new_n7632_), .A1(new_n7636_), .B0(new_n7634_), .Y(new_n7637_));
  INVX1    g07444(.A(new_n7637_), .Y(new_n7638_));
  OAI22X1  g07445(.A0(new_n7638_), .A1(new_n7631_), .B0(new_n7635_), .B1(new_n7633_), .Y(new_n7639_));
  AND2X1   g07446(.A(\a[45] ), .B(\a[43] ), .Y(new_n7640_));
  INVX1    g07447(.A(new_n7640_), .Y(new_n7641_));
  INVX1    g07448(.A(new_n3918_), .Y(new_n7642_));
  OAI22X1  g07449(.A0(new_n7642_), .A1(new_n1771_), .B0(new_n7641_), .B1(new_n3484_), .Y(new_n7643_));
  OAI21X1  g07450(.A0(new_n7353_), .A1(new_n3483_), .B0(new_n7643_), .Y(new_n7644_));
  AND2X1   g07451(.A(\a[45] ), .B(\a[25] ), .Y(new_n7645_));
  OAI22X1  g07452(.A0(new_n5268_), .A1(new_n1263_), .B0(new_n3037_), .B1(new_n1679_), .Y(new_n7646_));
  AOI21X1  g07453(.A0(new_n4992_), .A1(new_n1995_), .B0(new_n7643_), .Y(new_n7647_));
  AOI22X1  g07454(.A0(new_n7647_), .A1(new_n7646_), .B0(new_n7645_), .B1(new_n7644_), .Y(new_n7648_));
  XOR2X1   g07455(.A(new_n7648_), .B(new_n7639_), .Y(new_n7649_));
  INVX1    g07456(.A(new_n7649_), .Y(new_n7650_));
  INVX1    g07457(.A(new_n4484_), .Y(new_n7651_));
  INVX1    g07458(.A(new_n4321_), .Y(new_n7652_));
  NAND2X1  g07459(.A(\a[51] ), .B(\a[49] ), .Y(new_n7653_));
  OAI22X1  g07460(.A0(new_n7653_), .A1(new_n1149_), .B0(new_n7652_), .B1(new_n1794_), .Y(new_n7654_));
  OAI21X1  g07461(.A0(new_n7651_), .A1(new_n1521_), .B0(new_n7654_), .Y(new_n7655_));
  AND2X1   g07462(.A(\a[49] ), .B(\a[21] ), .Y(new_n7656_));
  AOI21X1  g07463(.A0(new_n4484_), .A1(new_n1099_), .B0(new_n7654_), .Y(new_n7657_));
  OAI22X1  g07464(.A0(new_n4349_), .A1(new_n752_), .B0(new_n4983_), .B1(new_n934_), .Y(new_n7658_));
  AOI22X1  g07465(.A0(new_n7658_), .A1(new_n7657_), .B0(new_n7656_), .B1(new_n7655_), .Y(new_n7659_));
  XOR2X1   g07466(.A(new_n7659_), .B(new_n7650_), .Y(new_n7660_));
  AND2X1   g07467(.A(new_n7660_), .B(new_n7630_), .Y(new_n7661_));
  XOR2X1   g07468(.A(new_n7660_), .B(new_n7630_), .Y(new_n7662_));
  OR2X1    g07469(.A(new_n7660_), .B(new_n7630_), .Y(new_n7663_));
  OAI21X1  g07470(.A0(new_n7661_), .A1(new_n7607_), .B0(new_n7663_), .Y(new_n7664_));
  OAI22X1  g07471(.A0(new_n7664_), .A1(new_n7661_), .B0(new_n7662_), .B1(new_n7607_), .Y(new_n7665_));
  OR2X1    g07472(.A(new_n7392_), .B(new_n7384_), .Y(new_n7666_));
  AND2X1   g07473(.A(new_n7392_), .B(new_n7384_), .Y(new_n7667_));
  OAI21X1  g07474(.A0(new_n7667_), .A1(new_n7382_), .B0(new_n7666_), .Y(new_n7668_));
  NAND4X1  g07475(.A(\a[61] ), .B(\a[59] ), .C(\a[11] ), .D(\a[9] ), .Y(new_n7669_));
  NAND4X1  g07476(.A(\a[61] ), .B(\a[60] ), .C(\a[10] ), .D(\a[9] ), .Y(new_n7670_));
  AOI22X1  g07477(.A0(new_n7670_), .A1(new_n7669_), .B0(new_n6427_), .B1(new_n1002_), .Y(new_n7671_));
  NAND4X1  g07478(.A(\a[60] ), .B(\a[59] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n7672_));
  NAND3X1  g07479(.A(new_n7670_), .B(new_n7669_), .C(new_n7672_), .Y(new_n7673_));
  AOI22X1  g07480(.A0(\a[60] ), .A1(\a[10] ), .B0(\a[59] ), .B1(\a[11] ), .Y(new_n7674_));
  NAND2X1  g07481(.A(\a[61] ), .B(\a[9] ), .Y(new_n7675_));
  OAI22X1  g07482(.A0(new_n7675_), .A1(new_n7671_), .B0(new_n7674_), .B1(new_n7673_), .Y(new_n7676_));
  INVX1    g07483(.A(new_n5574_), .Y(new_n7677_));
  NAND4X1  g07484(.A(\a[54] ), .B(\a[52] ), .C(\a[18] ), .D(\a[16] ), .Y(new_n7678_));
  NAND4X1  g07485(.A(\a[53] ), .B(\a[52] ), .C(\a[18] ), .D(\a[17] ), .Y(new_n7679_));
  AOI22X1  g07486(.A0(new_n7679_), .A1(new_n7678_), .B0(new_n5238_), .B1(new_n792_), .Y(new_n7680_));
  NAND4X1  g07487(.A(\a[54] ), .B(\a[53] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n7681_));
  NAND3X1  g07488(.A(new_n7679_), .B(new_n7678_), .C(new_n7681_), .Y(new_n7682_));
  AOI22X1  g07489(.A0(\a[54] ), .A1(\a[16] ), .B0(\a[53] ), .B1(\a[17] ), .Y(new_n7683_));
  OAI22X1  g07490(.A0(new_n7683_), .A1(new_n7682_), .B0(new_n7680_), .B1(new_n7677_), .Y(new_n7684_));
  XOR2X1   g07491(.A(new_n7684_), .B(new_n7676_), .Y(new_n7685_));
  NAND4X1  g07492(.A(\a[58] ), .B(\a[57] ), .C(\a[13] ), .D(\a[12] ), .Y(new_n7686_));
  NAND4X1  g07493(.A(\a[58] ), .B(\a[46] ), .C(\a[24] ), .D(\a[12] ), .Y(new_n7687_));
  AOI22X1  g07494(.A0(new_n7687_), .A1(new_n7686_), .B0(new_n6937_), .B1(new_n5531_), .Y(new_n7688_));
  NAND2X1  g07495(.A(\a[58] ), .B(\a[12] ), .Y(new_n7689_));
  AND2X1   g07496(.A(new_n6937_), .B(new_n5531_), .Y(new_n7690_));
  OR2X1    g07497(.A(new_n7688_), .B(new_n7690_), .Y(new_n7691_));
  AOI22X1  g07498(.A0(\a[57] ), .A1(\a[13] ), .B0(\a[46] ), .B1(\a[24] ), .Y(new_n7692_));
  OAI22X1  g07499(.A0(new_n7692_), .A1(new_n7691_), .B0(new_n7689_), .B1(new_n7688_), .Y(new_n7693_));
  XOR2X1   g07500(.A(new_n7693_), .B(new_n7685_), .Y(new_n7694_));
  INVX1    g07501(.A(new_n7469_), .Y(new_n7695_));
  XOR2X1   g07502(.A(new_n7695_), .B(new_n7431_), .Y(new_n7696_));
  AND2X1   g07503(.A(new_n3164_), .B(new_n2674_), .Y(new_n7697_));
  NOR4X1   g07504(.A(new_n2519_), .B(new_n2583_), .C(new_n2028_), .D(new_n2219_), .Y(new_n7698_));
  OAI22X1  g07505(.A0(new_n7698_), .A1(new_n7697_), .B0(new_n2919_), .B1(new_n6525_), .Y(new_n7699_));
  NAND3X1  g07506(.A(new_n7699_), .B(\a[38] ), .C(\a[32] ), .Y(new_n7700_));
  OAI21X1  g07507(.A0(new_n2919_), .A1(new_n6525_), .B0(new_n7699_), .Y(new_n7701_));
  AOI22X1  g07508(.A0(\a[37] ), .A1(\a[33] ), .B0(\a[36] ), .B1(\a[34] ), .Y(new_n7702_));
  OAI21X1  g07509(.A0(new_n7702_), .A1(new_n7701_), .B0(new_n7700_), .Y(new_n7703_));
  XOR2X1   g07510(.A(new_n7703_), .B(new_n7696_), .Y(new_n7704_));
  AND2X1   g07511(.A(new_n7390_), .B(new_n7388_), .Y(new_n7705_));
  OR2X1    g07512(.A(new_n7390_), .B(new_n7388_), .Y(new_n7706_));
  OAI21X1  g07513(.A0(new_n7705_), .A1(new_n7386_), .B0(new_n7706_), .Y(new_n7707_));
  XOR2X1   g07514(.A(new_n7707_), .B(new_n7704_), .Y(new_n7708_));
  XOR2X1   g07515(.A(new_n7708_), .B(new_n7694_), .Y(new_n7709_));
  XOR2X1   g07516(.A(new_n7709_), .B(new_n7668_), .Y(new_n7710_));
  XOR2X1   g07517(.A(new_n7710_), .B(new_n7665_), .Y(new_n7711_));
  XOR2X1   g07518(.A(new_n7711_), .B(new_n7605_), .Y(new_n7712_));
  XOR2X1   g07519(.A(new_n7550_), .B(new_n7572_), .Y(new_n7713_));
  AND2X1   g07520(.A(new_n7713_), .B(new_n7712_), .Y(new_n7714_));
  XOR2X1   g07521(.A(new_n7571_), .B(new_n7568_), .Y(new_n7715_));
  AOI21X1  g07522(.A0(new_n7550_), .A1(new_n7715_), .B0(new_n7712_), .Y(new_n7716_));
  AOI21X1  g07523(.A0(new_n7716_), .A1(new_n7574_), .B0(new_n7714_), .Y(new_n7717_));
  AND2X1   g07524(.A(new_n7717_), .B(new_n7548_), .Y(new_n7718_));
  INVX1    g07525(.A(new_n7718_), .Y(new_n7719_));
  INVX1    g07526(.A(new_n7535_), .Y(new_n7720_));
  NOR2X1   g07527(.A(new_n7539_), .B(new_n7720_), .Y(new_n7721_));
  INVX1    g07528(.A(new_n7721_), .Y(new_n7722_));
  AND2X1   g07529(.A(new_n7539_), .B(new_n7720_), .Y(new_n7723_));
  OAI21X1  g07530(.A0(new_n7544_), .A1(new_n7723_), .B0(new_n7722_), .Y(new_n7724_));
  NOR3X1   g07531(.A(new_n7717_), .B(new_n7547_), .C(new_n7546_), .Y(new_n7725_));
  INVX1    g07532(.A(new_n7725_), .Y(new_n7726_));
  AOI21X1  g07533(.A0(new_n7719_), .A1(new_n7726_), .B0(new_n7724_), .Y(new_n7727_));
  AND2X1   g07534(.A(new_n7726_), .B(new_n7724_), .Y(new_n7728_));
  AOI21X1  g07535(.A0(new_n7728_), .A1(new_n7719_), .B0(new_n7727_), .Y(\asquared[71] ));
  AOI21X1  g07536(.A0(new_n7726_), .A1(new_n7724_), .B0(new_n7718_), .Y(new_n7730_));
  OR2X1    g07537(.A(new_n7714_), .B(new_n7573_), .Y(new_n7731_));
  AND2X1   g07538(.A(new_n7709_), .B(new_n7668_), .Y(new_n7732_));
  AOI21X1  g07539(.A0(new_n7710_), .A1(new_n7665_), .B0(new_n7732_), .Y(new_n7733_));
  AND2X1   g07540(.A(new_n7695_), .B(new_n7431_), .Y(new_n7734_));
  AOI21X1  g07541(.A0(new_n7703_), .A1(new_n7696_), .B0(new_n7734_), .Y(new_n7735_));
  XOR2X1   g07542(.A(new_n7735_), .B(new_n7583_), .Y(new_n7736_));
  AND2X1   g07543(.A(new_n7506_), .B(new_n7440_), .Y(new_n7737_));
  AOI21X1  g07544(.A0(new_n7577_), .A1(new_n7499_), .B0(new_n7737_), .Y(new_n7738_));
  XOR2X1   g07545(.A(new_n7738_), .B(new_n7736_), .Y(new_n7739_));
  AND2X1   g07546(.A(new_n7584_), .B(new_n7578_), .Y(new_n7740_));
  AOI21X1  g07547(.A0(new_n7589_), .A1(new_n7585_), .B0(new_n7740_), .Y(new_n7741_));
  XOR2X1   g07548(.A(new_n7741_), .B(new_n7739_), .Y(new_n7742_));
  AND2X1   g07549(.A(new_n7707_), .B(new_n7704_), .Y(new_n7743_));
  AOI21X1  g07550(.A0(new_n7708_), .A1(new_n7694_), .B0(new_n7743_), .Y(new_n7744_));
  XOR2X1   g07551(.A(new_n7744_), .B(new_n7742_), .Y(new_n7745_));
  INVX1    g07552(.A(new_n7745_), .Y(new_n7746_));
  INVX1    g07553(.A(new_n7602_), .Y(new_n7747_));
  OR2X1    g07554(.A(new_n7747_), .B(new_n7480_), .Y(new_n7748_));
  OAI21X1  g07555(.A0(new_n7603_), .A1(new_n7590_), .B0(new_n7748_), .Y(new_n7749_));
  XOR2X1   g07556(.A(new_n7749_), .B(new_n7746_), .Y(new_n7750_));
  XOR2X1   g07557(.A(new_n7750_), .B(new_n7733_), .Y(new_n7751_));
  AND2X1   g07558(.A(new_n7604_), .B(new_n7576_), .Y(new_n7752_));
  AOI21X1  g07559(.A0(new_n7711_), .A1(new_n7605_), .B0(new_n7752_), .Y(new_n7753_));
  XOR2X1   g07560(.A(new_n7753_), .B(new_n7751_), .Y(new_n7754_));
  INVX1    g07561(.A(new_n7567_), .Y(new_n7755_));
  NOR2X1   g07562(.A(new_n7755_), .B(new_n7552_), .Y(new_n7756_));
  INVX1    g07563(.A(new_n7756_), .Y(new_n7757_));
  OAI21X1  g07564(.A0(new_n7571_), .A1(new_n7568_), .B0(new_n7757_), .Y(new_n7758_));
  AND2X1   g07565(.A(new_n7684_), .B(new_n7676_), .Y(new_n7759_));
  AOI21X1  g07566(.A0(new_n7693_), .A1(new_n7685_), .B0(new_n7759_), .Y(new_n7760_));
  AND2X1   g07567(.A(new_n7519_), .B(new_n7489_), .Y(new_n7761_));
  AOI21X1  g07568(.A0(new_n7558_), .A1(new_n7557_), .B0(new_n7761_), .Y(new_n7762_));
  XOR2X1   g07569(.A(new_n7762_), .B(new_n7760_), .Y(new_n7763_));
  INVX1    g07570(.A(new_n7639_), .Y(new_n7764_));
  OR2X1    g07571(.A(new_n7648_), .B(new_n7764_), .Y(new_n7765_));
  OAI21X1  g07572(.A0(new_n7659_), .A1(new_n7649_), .B0(new_n7765_), .Y(new_n7766_));
  XOR2X1   g07573(.A(new_n7766_), .B(new_n7763_), .Y(new_n7767_));
  XOR2X1   g07574(.A(new_n7767_), .B(new_n7664_), .Y(new_n7768_));
  INVX1    g07575(.A(new_n7616_), .Y(new_n7769_));
  OR2X1    g07576(.A(new_n7624_), .B(new_n7769_), .Y(new_n7770_));
  OAI21X1  g07577(.A0(new_n7628_), .A1(new_n7625_), .B0(new_n7770_), .Y(new_n7771_));
  XOR2X1   g07578(.A(new_n7691_), .B(new_n7673_), .Y(new_n7772_));
  XOR2X1   g07579(.A(new_n7772_), .B(new_n7647_), .Y(new_n7773_));
  XOR2X1   g07580(.A(new_n7637_), .B(new_n7622_), .Y(new_n7774_));
  XOR2X1   g07581(.A(new_n7774_), .B(new_n7614_), .Y(new_n7775_));
  XOR2X1   g07582(.A(new_n7775_), .B(new_n7773_), .Y(new_n7776_));
  XOR2X1   g07583(.A(new_n7776_), .B(new_n7771_), .Y(new_n7777_));
  XOR2X1   g07584(.A(new_n7777_), .B(new_n7768_), .Y(new_n7778_));
  XOR2X1   g07585(.A(new_n7778_), .B(new_n7758_), .Y(new_n7779_));
  INVX1    g07586(.A(new_n7779_), .Y(new_n7780_));
  INVX1    g07587(.A(new_n7565_), .Y(new_n7781_));
  OR2X1    g07588(.A(new_n7781_), .B(new_n7556_), .Y(new_n7782_));
  OAI21X1  g07589(.A0(new_n7566_), .A1(new_n7554_), .B0(new_n7782_), .Y(new_n7783_));
  AOI21X1  g07590(.A0(\a[62] ), .A1(\a[9] ), .B0(\a[36] ), .Y(new_n7784_));
  AND2X1   g07591(.A(\a[49] ), .B(\a[22] ), .Y(new_n7785_));
  INVX1    g07592(.A(new_n7785_), .Y(new_n7786_));
  NOR3X1   g07593(.A(new_n6606_), .B(new_n2583_), .C(new_n341_), .Y(new_n7787_));
  NOR3X1   g07594(.A(new_n7786_), .B(new_n7787_), .C(new_n7784_), .Y(new_n7788_));
  INVX1    g07595(.A(new_n7784_), .Y(new_n7789_));
  AOI21X1  g07596(.A0(new_n7785_), .A1(new_n7789_), .B0(new_n7787_), .Y(new_n7790_));
  INVX1    g07597(.A(new_n7790_), .Y(new_n7791_));
  OAI22X1  g07598(.A0(new_n7791_), .A1(new_n7784_), .B0(new_n7788_), .B1(new_n7786_), .Y(new_n7792_));
  INVX1    g07599(.A(new_n7164_), .Y(new_n7793_));
  NAND2X1  g07600(.A(\a[52] ), .B(\a[50] ), .Y(new_n7794_));
  OAI22X1  g07601(.A0(new_n7794_), .A1(new_n1149_), .B0(new_n7651_), .B1(new_n1794_), .Y(new_n7795_));
  OAI21X1  g07602(.A0(new_n7793_), .A1(new_n1521_), .B0(new_n7795_), .Y(new_n7796_));
  AND2X1   g07603(.A(\a[50] ), .B(\a[21] ), .Y(new_n7797_));
  OAI22X1  g07604(.A0(new_n4354_), .A1(new_n752_), .B0(new_n4349_), .B1(new_n934_), .Y(new_n7798_));
  AOI21X1  g07605(.A0(new_n7164_), .A1(new_n1099_), .B0(new_n7795_), .Y(new_n7799_));
  AOI22X1  g07606(.A0(new_n7799_), .A1(new_n7798_), .B0(new_n7797_), .B1(new_n7796_), .Y(new_n7800_));
  XOR2X1   g07607(.A(new_n7800_), .B(new_n7792_), .Y(new_n7801_));
  AND2X1   g07608(.A(\a[37] ), .B(\a[34] ), .Y(new_n7802_));
  AND2X1   g07609(.A(new_n7802_), .B(new_n2682_), .Y(new_n7803_));
  AOI22X1  g07610(.A0(new_n3164_), .A1(new_n2918_), .B0(new_n3163_), .B1(new_n2682_), .Y(new_n7804_));
  OR2X1    g07611(.A(new_n7804_), .B(new_n7803_), .Y(new_n7805_));
  NAND4X1  g07612(.A(\a[37] ), .B(\a[36] ), .C(\a[35] ), .D(\a[34] ), .Y(new_n7806_));
  AND2X1   g07613(.A(new_n7804_), .B(new_n7806_), .Y(new_n7807_));
  OR2X1    g07614(.A(new_n7802_), .B(new_n2682_), .Y(new_n7808_));
  AOI22X1  g07615(.A0(new_n7808_), .A1(new_n7807_), .B0(new_n7805_), .B1(new_n3163_), .Y(new_n7809_));
  XOR2X1   g07616(.A(new_n7809_), .B(new_n7801_), .Y(new_n7810_));
  XOR2X1   g07617(.A(new_n7701_), .B(new_n7682_), .Y(new_n7811_));
  NAND4X1  g07618(.A(\a[63] ), .B(\a[60] ), .C(\a[11] ), .D(\a[8] ), .Y(new_n7812_));
  NAND4X1  g07619(.A(\a[61] ), .B(\a[60] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n7813_));
  AOI22X1  g07620(.A0(new_n7813_), .A1(new_n7812_), .B0(new_n6688_), .B1(new_n324_), .Y(new_n7814_));
  AND2X1   g07621(.A(\a[60] ), .B(\a[11] ), .Y(new_n7815_));
  INVX1    g07622(.A(new_n7815_), .Y(new_n7816_));
  AOI22X1  g07623(.A0(\a[63] ), .A1(\a[8] ), .B0(\a[61] ), .B1(\a[10] ), .Y(new_n7817_));
  AOI21X1  g07624(.A0(new_n6688_), .A1(new_n324_), .B0(new_n7814_), .Y(new_n7818_));
  INVX1    g07625(.A(new_n7818_), .Y(new_n7819_));
  OAI22X1  g07626(.A0(new_n7819_), .A1(new_n7817_), .B0(new_n7816_), .B1(new_n7814_), .Y(new_n7820_));
  INVX1    g07627(.A(new_n7820_), .Y(new_n7821_));
  XOR2X1   g07628(.A(new_n7821_), .B(new_n7811_), .Y(new_n7822_));
  NOR2X1   g07629(.A(new_n7563_), .B(new_n7561_), .Y(new_n7823_));
  AOI21X1  g07630(.A0(new_n7564_), .A1(new_n7559_), .B0(new_n7823_), .Y(new_n7824_));
  XOR2X1   g07631(.A(new_n7824_), .B(new_n7822_), .Y(new_n7825_));
  XOR2X1   g07632(.A(new_n7825_), .B(new_n7810_), .Y(new_n7826_));
  XOR2X1   g07633(.A(new_n7826_), .B(new_n7783_), .Y(new_n7827_));
  INVX1    g07634(.A(new_n7592_), .Y(new_n7828_));
  NAND2X1  g07635(.A(new_n7595_), .B(new_n7828_), .Y(new_n7829_));
  OAI21X1  g07636(.A0(new_n7601_), .A1(new_n7596_), .B0(new_n7829_), .Y(new_n7830_));
  AOI22X1  g07637(.A0(new_n4992_), .A1(new_n1671_), .B0(new_n3208_), .B1(new_n1484_), .Y(new_n7831_));
  AOI21X1  g07638(.A0(new_n3462_), .A1(new_n1674_), .B0(new_n7831_), .Y(new_n7832_));
  OAI21X1  g07639(.A0(new_n6502_), .A1(new_n1675_), .B0(new_n7831_), .Y(new_n7833_));
  AOI22X1  g07640(.A0(\a[43] ), .A1(\a[28] ), .B0(\a[42] ), .B1(\a[29] ), .Y(new_n7834_));
  NAND2X1  g07641(.A(\a[44] ), .B(\a[27] ), .Y(new_n7835_));
  OAI22X1  g07642(.A0(new_n7835_), .A1(new_n7832_), .B0(new_n7834_), .B1(new_n7833_), .Y(new_n7836_));
  NAND4X1  g07643(.A(\a[41] ), .B(\a[39] ), .C(\a[32] ), .D(\a[30] ), .Y(new_n7837_));
  NAND4X1  g07644(.A(\a[41] ), .B(\a[40] ), .C(\a[31] ), .D(\a[30] ), .Y(new_n7838_));
  AOI22X1  g07645(.A0(new_n7838_), .A1(new_n7837_), .B0(new_n4077_), .B1(new_n2671_), .Y(new_n7839_));
  NAND2X1  g07646(.A(\a[41] ), .B(\a[30] ), .Y(new_n7840_));
  AOI22X1  g07647(.A0(\a[40] ), .A1(\a[31] ), .B0(\a[39] ), .B1(\a[32] ), .Y(new_n7841_));
  AOI21X1  g07648(.A0(new_n4077_), .A1(new_n2671_), .B0(new_n7839_), .Y(new_n7842_));
  INVX1    g07649(.A(new_n7842_), .Y(new_n7843_));
  OAI22X1  g07650(.A0(new_n7843_), .A1(new_n7841_), .B0(new_n7840_), .B1(new_n7839_), .Y(new_n7844_));
  XOR2X1   g07651(.A(new_n7844_), .B(new_n7836_), .Y(new_n7845_));
  NAND2X1  g07652(.A(\a[48] ), .B(\a[23] ), .Y(new_n7846_));
  AOI22X1  g07653(.A0(\a[54] ), .A1(\a[17] ), .B0(\a[53] ), .B1(\a[18] ), .Y(new_n7847_));
  AND2X1   g07654(.A(new_n5238_), .B(new_n796_), .Y(new_n7848_));
  NOR3X1   g07655(.A(new_n7847_), .B(new_n7848_), .C(new_n7846_), .Y(new_n7849_));
  OAI22X1  g07656(.A0(new_n7847_), .A1(new_n7846_), .B0(new_n5239_), .B1(new_n797_), .Y(new_n7850_));
  OAI22X1  g07657(.A0(new_n7850_), .A1(new_n7847_), .B0(new_n7849_), .B1(new_n7846_), .Y(new_n7851_));
  XOR2X1   g07658(.A(new_n7851_), .B(new_n7845_), .Y(new_n7852_));
  INVX1    g07659(.A(new_n7657_), .Y(new_n7853_));
  NAND2X1  g07660(.A(\a[58] ), .B(\a[13] ), .Y(new_n7854_));
  NAND2X1  g07661(.A(\a[59] ), .B(\a[12] ), .Y(new_n7855_));
  AOI22X1  g07662(.A0(new_n7855_), .A1(new_n7854_), .B0(new_n6121_), .B1(new_n586_), .Y(new_n7856_));
  XOR2X1   g07663(.A(new_n7856_), .B(new_n7853_), .Y(new_n7857_));
  NAND4X1  g07664(.A(\a[57] ), .B(\a[55] ), .C(\a[16] ), .D(\a[14] ), .Y(new_n7858_));
  NAND4X1  g07665(.A(\a[57] ), .B(\a[56] ), .C(\a[15] ), .D(\a[14] ), .Y(new_n7859_));
  AOI22X1  g07666(.A0(new_n7859_), .A1(new_n7858_), .B0(new_n6237_), .B1(new_n689_), .Y(new_n7860_));
  NAND4X1  g07667(.A(\a[56] ), .B(\a[55] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n7861_));
  NAND3X1  g07668(.A(new_n7859_), .B(new_n7858_), .C(new_n7861_), .Y(new_n7862_));
  AOI22X1  g07669(.A0(\a[56] ), .A1(\a[15] ), .B0(\a[55] ), .B1(\a[16] ), .Y(new_n7863_));
  NAND2X1  g07670(.A(\a[57] ), .B(\a[14] ), .Y(new_n7864_));
  OAI22X1  g07671(.A0(new_n7864_), .A1(new_n7860_), .B0(new_n7863_), .B1(new_n7862_), .Y(new_n7865_));
  NAND4X1  g07672(.A(\a[47] ), .B(\a[45] ), .C(\a[26] ), .D(\a[24] ), .Y(new_n7866_));
  NAND4X1  g07673(.A(\a[47] ), .B(\a[46] ), .C(\a[25] ), .D(\a[24] ), .Y(new_n7867_));
  AOI22X1  g07674(.A0(new_n7867_), .A1(new_n7866_), .B0(new_n3809_), .B1(new_n1770_), .Y(new_n7868_));
  NAND2X1  g07675(.A(\a[47] ), .B(\a[24] ), .Y(new_n7869_));
  NAND4X1  g07676(.A(\a[46] ), .B(\a[45] ), .C(\a[26] ), .D(\a[25] ), .Y(new_n7870_));
  NAND3X1  g07677(.A(new_n7867_), .B(new_n7866_), .C(new_n7870_), .Y(new_n7871_));
  AOI22X1  g07678(.A0(\a[46] ), .A1(\a[25] ), .B0(\a[45] ), .B1(\a[26] ), .Y(new_n7872_));
  OAI22X1  g07679(.A0(new_n7872_), .A1(new_n7871_), .B0(new_n7869_), .B1(new_n7868_), .Y(new_n7873_));
  XOR2X1   g07680(.A(new_n7873_), .B(new_n7865_), .Y(new_n7874_));
  XOR2X1   g07681(.A(new_n7874_), .B(new_n7857_), .Y(new_n7875_));
  XOR2X1   g07682(.A(new_n7875_), .B(new_n7852_), .Y(new_n7876_));
  XOR2X1   g07683(.A(new_n7876_), .B(new_n7830_), .Y(new_n7877_));
  XOR2X1   g07684(.A(new_n7877_), .B(new_n7827_), .Y(new_n7878_));
  XOR2X1   g07685(.A(new_n7878_), .B(new_n7780_), .Y(new_n7879_));
  XOR2X1   g07686(.A(new_n7879_), .B(new_n7754_), .Y(new_n7880_));
  NOR2X1   g07687(.A(new_n7880_), .B(new_n7731_), .Y(new_n7881_));
  AND2X1   g07688(.A(new_n7880_), .B(new_n7731_), .Y(new_n7882_));
  OR2X1    g07689(.A(new_n7882_), .B(new_n7881_), .Y(new_n7883_));
  XOR2X1   g07690(.A(new_n7883_), .B(new_n7730_), .Y(\asquared[72] ));
  AND2X1   g07691(.A(new_n7826_), .B(new_n7783_), .Y(new_n7885_));
  AOI21X1  g07692(.A0(new_n7877_), .A1(new_n7827_), .B0(new_n7885_), .Y(new_n7886_));
  INVX1    g07693(.A(new_n7886_), .Y(new_n7887_));
  NOR2X1   g07694(.A(new_n7775_), .B(new_n7773_), .Y(new_n7888_));
  AOI21X1  g07695(.A0(new_n7776_), .A1(new_n7771_), .B0(new_n7888_), .Y(new_n7889_));
  AND2X1   g07696(.A(new_n7701_), .B(new_n7682_), .Y(new_n7890_));
  AOI21X1  g07697(.A0(new_n7820_), .A1(new_n7811_), .B0(new_n7890_), .Y(new_n7891_));
  NAND4X1  g07698(.A(\a[43] ), .B(\a[41] ), .C(\a[31] ), .D(\a[29] ), .Y(new_n7892_));
  NAND4X1  g07699(.A(\a[43] ), .B(\a[42] ), .C(\a[30] ), .D(\a[29] ), .Y(new_n7893_));
  AOI22X1  g07700(.A0(new_n7893_), .A1(new_n7892_), .B0(new_n3607_), .B1(new_n2075_), .Y(new_n7894_));
  AND2X1   g07701(.A(\a[43] ), .B(\a[29] ), .Y(new_n7895_));
  INVX1    g07702(.A(new_n7895_), .Y(new_n7896_));
  AOI22X1  g07703(.A0(\a[42] ), .A1(\a[30] ), .B0(\a[41] ), .B1(\a[31] ), .Y(new_n7897_));
  AOI21X1  g07704(.A0(new_n3607_), .A1(new_n2075_), .B0(new_n7894_), .Y(new_n7898_));
  INVX1    g07705(.A(new_n7898_), .Y(new_n7899_));
  OAI22X1  g07706(.A0(new_n7899_), .A1(new_n7897_), .B0(new_n7896_), .B1(new_n7894_), .Y(new_n7900_));
  XOR2X1   g07707(.A(new_n7900_), .B(new_n7891_), .Y(new_n7901_));
  INVX1    g07708(.A(new_n7901_), .Y(new_n7902_));
  NOR2X1   g07709(.A(new_n7637_), .B(new_n7622_), .Y(new_n7903_));
  AOI21X1  g07710(.A0(new_n7774_), .A1(new_n7615_), .B0(new_n7903_), .Y(new_n7904_));
  XOR2X1   g07711(.A(new_n7904_), .B(new_n7902_), .Y(new_n7905_));
  XOR2X1   g07712(.A(new_n7905_), .B(new_n7889_), .Y(new_n7906_));
  NOR2X1   g07713(.A(new_n7824_), .B(new_n7822_), .Y(new_n7907_));
  AOI21X1  g07714(.A0(new_n7825_), .A1(new_n7810_), .B0(new_n7907_), .Y(new_n7908_));
  XOR2X1   g07715(.A(new_n7908_), .B(new_n7906_), .Y(new_n7909_));
  AND2X1   g07716(.A(new_n7767_), .B(new_n7664_), .Y(new_n7910_));
  AOI21X1  g07717(.A0(new_n7777_), .A1(new_n7768_), .B0(new_n7910_), .Y(new_n7911_));
  XOR2X1   g07718(.A(new_n7911_), .B(new_n7909_), .Y(new_n7912_));
  XOR2X1   g07719(.A(new_n7912_), .B(new_n7887_), .Y(new_n7913_));
  AND2X1   g07720(.A(new_n7778_), .B(new_n7758_), .Y(new_n7914_));
  AOI21X1  g07721(.A0(new_n7878_), .A1(new_n7779_), .B0(new_n7914_), .Y(new_n7915_));
  XOR2X1   g07722(.A(new_n7915_), .B(new_n7913_), .Y(new_n7916_));
  NAND2X1  g07723(.A(new_n7749_), .B(new_n7745_), .Y(new_n7917_));
  OAI21X1  g07724(.A0(new_n7750_), .A1(new_n7733_), .B0(new_n7917_), .Y(new_n7918_));
  AND2X1   g07725(.A(new_n7844_), .B(new_n7836_), .Y(new_n7919_));
  AOI21X1  g07726(.A0(new_n7851_), .A1(new_n7845_), .B0(new_n7919_), .Y(new_n7920_));
  INVX1    g07727(.A(new_n7647_), .Y(new_n7921_));
  AND2X1   g07728(.A(new_n7691_), .B(new_n7673_), .Y(new_n7922_));
  AOI21X1  g07729(.A0(new_n7772_), .A1(new_n7921_), .B0(new_n7922_), .Y(new_n7923_));
  XOR2X1   g07730(.A(new_n7923_), .B(new_n7920_), .Y(new_n7924_));
  INVX1    g07731(.A(new_n7792_), .Y(new_n7925_));
  OR2X1    g07732(.A(new_n7800_), .B(new_n7925_), .Y(new_n7926_));
  OAI21X1  g07733(.A0(new_n7809_), .A1(new_n7801_), .B0(new_n7926_), .Y(new_n7927_));
  XOR2X1   g07734(.A(new_n7927_), .B(new_n7924_), .Y(new_n7928_));
  AND2X1   g07735(.A(new_n7875_), .B(new_n7852_), .Y(new_n7929_));
  AOI21X1  g07736(.A0(new_n7876_), .A1(new_n7830_), .B0(new_n7929_), .Y(new_n7930_));
  XOR2X1   g07737(.A(new_n7930_), .B(new_n7928_), .Y(new_n7931_));
  AND2X1   g07738(.A(new_n7873_), .B(new_n7865_), .Y(new_n7932_));
  AOI21X1  g07739(.A0(new_n7874_), .A1(new_n7857_), .B0(new_n7932_), .Y(new_n7933_));
  XOR2X1   g07740(.A(new_n7850_), .B(new_n7833_), .Y(new_n7934_));
  XOR2X1   g07741(.A(new_n7934_), .B(new_n7842_), .Y(new_n7935_));
  INVX1    g07742(.A(new_n7799_), .Y(new_n7936_));
  XOR2X1   g07743(.A(new_n7807_), .B(new_n7790_), .Y(new_n7937_));
  XOR2X1   g07744(.A(new_n7937_), .B(new_n7936_), .Y(new_n7938_));
  INVX1    g07745(.A(new_n7938_), .Y(new_n7939_));
  XOR2X1   g07746(.A(new_n7939_), .B(new_n7935_), .Y(new_n7940_));
  XOR2X1   g07747(.A(new_n7940_), .B(new_n7933_), .Y(new_n7941_));
  XOR2X1   g07748(.A(new_n7941_), .B(new_n7931_), .Y(new_n7942_));
  XOR2X1   g07749(.A(new_n7942_), .B(new_n7918_), .Y(new_n7943_));
  NOR2X1   g07750(.A(new_n7762_), .B(new_n7760_), .Y(new_n7944_));
  AOI21X1  g07751(.A0(new_n7766_), .A1(new_n7763_), .B0(new_n7944_), .Y(new_n7945_));
  AOI22X1  g07752(.A0(\a[56] ), .A1(\a[16] ), .B0(\a[49] ), .B1(\a[23] ), .Y(new_n7946_));
  AND2X1   g07753(.A(\a[40] ), .B(\a[32] ), .Y(new_n7947_));
  INVX1    g07754(.A(new_n7947_), .Y(new_n7948_));
  NOR4X1   g07755(.A(new_n6022_), .B(new_n3915_), .C(new_n1216_), .D(new_n571_), .Y(new_n7949_));
  NOR3X1   g07756(.A(new_n7948_), .B(new_n7949_), .C(new_n7946_), .Y(new_n7950_));
  INVX1    g07757(.A(new_n7946_), .Y(new_n7951_));
  AOI21X1  g07758(.A0(new_n7947_), .A1(new_n7951_), .B0(new_n7949_), .Y(new_n7952_));
  INVX1    g07759(.A(new_n7952_), .Y(new_n7953_));
  OAI22X1  g07760(.A0(new_n7953_), .A1(new_n7946_), .B0(new_n7950_), .B1(new_n7948_), .Y(new_n7954_));
  AOI22X1  g07761(.A0(\a[51] ), .A1(\a[21] ), .B0(\a[50] ), .B1(\a[22] ), .Y(new_n7955_));
  INVX1    g07762(.A(new_n7955_), .Y(new_n7956_));
  NAND4X1  g07763(.A(\a[51] ), .B(\a[50] ), .C(\a[22] ), .D(\a[21] ), .Y(new_n7957_));
  AOI21X1  g07764(.A0(new_n7956_), .A1(new_n7957_), .B0(new_n6527_), .Y(new_n7958_));
  AOI22X1  g07765(.A0(new_n7956_), .A1(new_n6526_), .B0(new_n4484_), .B1(new_n1154_), .Y(new_n7959_));
  AOI21X1  g07766(.A0(new_n7959_), .A1(new_n7956_), .B0(new_n7958_), .Y(new_n7960_));
  XOR2X1   g07767(.A(new_n7960_), .B(new_n7954_), .Y(new_n7961_));
  AND2X1   g07768(.A(\a[55] ), .B(\a[17] ), .Y(new_n7962_));
  AND2X1   g07769(.A(new_n5240_), .B(new_n796_), .Y(new_n7963_));
  NOR4X1   g07770(.A(new_n4906_), .B(new_n4354_), .C(new_n934_), .D(new_n616_), .Y(new_n7964_));
  OAI22X1  g07771(.A0(new_n7964_), .A1(new_n7963_), .B0(new_n7338_), .B1(new_n1520_), .Y(new_n7965_));
  OAI22X1  g07772(.A0(new_n4835_), .A1(new_n675_), .B0(new_n4354_), .B1(new_n934_), .Y(new_n7966_));
  OAI21X1  g07773(.A0(new_n7338_), .A1(new_n1520_), .B0(new_n7965_), .Y(new_n7967_));
  INVX1    g07774(.A(new_n7967_), .Y(new_n7968_));
  AOI22X1  g07775(.A0(new_n7968_), .A1(new_n7966_), .B0(new_n7965_), .B1(new_n7962_), .Y(new_n7969_));
  XOR2X1   g07776(.A(new_n7969_), .B(new_n7961_), .Y(new_n7970_));
  INVX1    g07777(.A(new_n7970_), .Y(new_n7971_));
  INVX1    g07778(.A(new_n6789_), .Y(new_n7972_));
  INVX1    g07779(.A(new_n6688_), .Y(new_n7973_));
  OAI22X1  g07780(.A0(new_n7973_), .A1(new_n1519_), .B0(new_n7972_), .B1(new_n735_), .Y(new_n7974_));
  OAI21X1  g07781(.A0(new_n6557_), .A1(new_n1517_), .B0(new_n7974_), .Y(new_n7975_));
  AOI21X1  g07782(.A0(new_n6556_), .A1(new_n1002_), .B0(new_n7974_), .Y(new_n7976_));
  OAI22X1  g07783(.A0(new_n6606_), .A1(new_n570_), .B0(new_n6023_), .B1(new_n488_), .Y(new_n7977_));
  AND2X1   g07784(.A(\a[63] ), .B(\a[9] ), .Y(new_n7978_));
  AOI22X1  g07785(.A0(new_n7978_), .A1(new_n7975_), .B0(new_n7977_), .B1(new_n7976_), .Y(new_n7979_));
  AOI22X1  g07786(.A0(new_n7856_), .A1(new_n7853_), .B0(new_n6121_), .B1(new_n586_), .Y(new_n7980_));
  AND2X1   g07787(.A(\a[60] ), .B(\a[12] ), .Y(new_n7981_));
  INVX1    g07788(.A(new_n7981_), .Y(new_n7982_));
  AOI22X1  g07789(.A0(\a[48] ), .A1(\a[24] ), .B0(\a[47] ), .B1(\a[25] ), .Y(new_n7983_));
  AND2X1   g07790(.A(new_n4272_), .B(new_n1532_), .Y(new_n7984_));
  NOR3X1   g07791(.A(new_n7983_), .B(new_n7984_), .C(new_n7982_), .Y(new_n7985_));
  INVX1    g07792(.A(new_n7983_), .Y(new_n7986_));
  AOI21X1  g07793(.A0(new_n7986_), .A1(new_n7981_), .B0(new_n7984_), .Y(new_n7987_));
  INVX1    g07794(.A(new_n7987_), .Y(new_n7988_));
  OAI22X1  g07795(.A0(new_n7988_), .A1(new_n7983_), .B0(new_n7985_), .B1(new_n7982_), .Y(new_n7989_));
  AND2X1   g07796(.A(new_n7989_), .B(new_n7980_), .Y(new_n7990_));
  XOR2X1   g07797(.A(new_n7989_), .B(new_n7980_), .Y(new_n7991_));
  OAI21X1  g07798(.A0(new_n7989_), .A1(new_n7980_), .B0(new_n7979_), .Y(new_n7992_));
  OAI22X1  g07799(.A0(new_n7992_), .A1(new_n7990_), .B0(new_n7991_), .B1(new_n7979_), .Y(new_n7993_));
  XOR2X1   g07800(.A(new_n7993_), .B(new_n7971_), .Y(new_n7994_));
  INVX1    g07801(.A(new_n7994_), .Y(new_n7995_));
  XOR2X1   g07802(.A(new_n7995_), .B(new_n7945_), .Y(new_n7996_));
  AND2X1   g07803(.A(new_n7589_), .B(new_n7585_), .Y(new_n7997_));
  OAI21X1  g07804(.A0(new_n7997_), .A1(new_n7740_), .B0(new_n7739_), .Y(new_n7998_));
  OAI21X1  g07805(.A0(new_n7744_), .A1(new_n7742_), .B0(new_n7998_), .Y(new_n7999_));
  XOR2X1   g07806(.A(new_n7871_), .B(new_n7862_), .Y(new_n8000_));
  XOR2X1   g07807(.A(new_n8000_), .B(new_n7819_), .Y(new_n8001_));
  INVX1    g07808(.A(new_n8001_), .Y(new_n8002_));
  OR2X1    g07809(.A(new_n7735_), .B(new_n7582_), .Y(new_n8003_));
  OAI21X1  g07810(.A0(new_n7738_), .A1(new_n7736_), .B0(new_n8003_), .Y(new_n8004_));
  XOR2X1   g07811(.A(new_n8004_), .B(new_n8002_), .Y(new_n8005_));
  NAND4X1  g07812(.A(\a[59] ), .B(\a[57] ), .C(\a[15] ), .D(\a[13] ), .Y(new_n8006_));
  NAND4X1  g07813(.A(\a[59] ), .B(\a[58] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n8007_));
  AOI22X1  g07814(.A0(new_n8007_), .A1(new_n8006_), .B0(new_n6119_), .B1(new_n691_), .Y(new_n8008_));
  NAND4X1  g07815(.A(\a[58] ), .B(\a[57] ), .C(\a[15] ), .D(\a[14] ), .Y(new_n8009_));
  NAND3X1  g07816(.A(new_n8007_), .B(new_n8006_), .C(new_n8009_), .Y(new_n8010_));
  AOI22X1  g07817(.A0(\a[58] ), .A1(\a[14] ), .B0(\a[57] ), .B1(\a[15] ), .Y(new_n8011_));
  NAND2X1  g07818(.A(\a[59] ), .B(\a[13] ), .Y(new_n8012_));
  OAI22X1  g07819(.A0(new_n8012_), .A1(new_n8008_), .B0(new_n8011_), .B1(new_n8010_), .Y(new_n8013_));
  NAND4X1  g07820(.A(\a[46] ), .B(\a[44] ), .C(\a[28] ), .D(\a[26] ), .Y(new_n8014_));
  NAND4X1  g07821(.A(\a[46] ), .B(\a[45] ), .C(\a[27] ), .D(\a[26] ), .Y(new_n8015_));
  AOI22X1  g07822(.A0(new_n8015_), .A1(new_n8014_), .B0(new_n3918_), .B1(new_n1671_), .Y(new_n8016_));
  NAND2X1  g07823(.A(\a[46] ), .B(\a[26] ), .Y(new_n8017_));
  NAND4X1  g07824(.A(\a[45] ), .B(\a[44] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n8018_));
  NAND3X1  g07825(.A(new_n8015_), .B(new_n8014_), .C(new_n8018_), .Y(new_n8019_));
  AOI22X1  g07826(.A0(\a[45] ), .A1(\a[27] ), .B0(\a[44] ), .B1(\a[28] ), .Y(new_n8020_));
  OAI22X1  g07827(.A0(new_n8020_), .A1(new_n8019_), .B0(new_n8017_), .B1(new_n8016_), .Y(new_n8021_));
  XOR2X1   g07828(.A(new_n8021_), .B(new_n8013_), .Y(new_n8022_));
  AND2X1   g07829(.A(\a[53] ), .B(\a[19] ), .Y(new_n8023_));
  INVX1    g07830(.A(new_n8023_), .Y(new_n8024_));
  AOI22X1  g07831(.A0(\a[39] ), .A1(\a[33] ), .B0(\a[38] ), .B1(\a[34] ), .Y(new_n8025_));
  AND2X1   g07832(.A(new_n3503_), .B(new_n2918_), .Y(new_n8026_));
  NOR3X1   g07833(.A(new_n8025_), .B(new_n8026_), .C(new_n8024_), .Y(new_n8027_));
  NOR2X1   g07834(.A(new_n8027_), .B(new_n8026_), .Y(new_n8028_));
  INVX1    g07835(.A(new_n8028_), .Y(new_n8029_));
  OAI22X1  g07836(.A0(new_n8029_), .A1(new_n8025_), .B0(new_n8027_), .B1(new_n8024_), .Y(new_n8030_));
  XOR2X1   g07837(.A(new_n8030_), .B(new_n8022_), .Y(new_n8031_));
  INVX1    g07838(.A(new_n8031_), .Y(new_n8032_));
  XOR2X1   g07839(.A(new_n8032_), .B(new_n8005_), .Y(new_n8033_));
  INVX1    g07840(.A(new_n8033_), .Y(new_n8034_));
  XOR2X1   g07841(.A(new_n8034_), .B(new_n7999_), .Y(new_n8035_));
  XOR2X1   g07842(.A(new_n8035_), .B(new_n7996_), .Y(new_n8036_));
  XOR2X1   g07843(.A(new_n8036_), .B(new_n7943_), .Y(new_n8037_));
  XOR2X1   g07844(.A(new_n8037_), .B(new_n7916_), .Y(new_n8038_));
  AND2X1   g07845(.A(new_n7711_), .B(new_n7605_), .Y(new_n8039_));
  OAI21X1  g07846(.A0(new_n8039_), .A1(new_n7752_), .B0(new_n7751_), .Y(new_n8040_));
  OAI21X1  g07847(.A0(new_n7879_), .A1(new_n7754_), .B0(new_n8040_), .Y(new_n8041_));
  AND2X1   g07848(.A(new_n8041_), .B(new_n8038_), .Y(new_n8042_));
  INVX1    g07849(.A(new_n8042_), .Y(new_n8043_));
  INVX1    g07850(.A(new_n7882_), .Y(new_n8044_));
  OAI21X1  g07851(.A0(new_n7881_), .A1(new_n7730_), .B0(new_n8044_), .Y(new_n8045_));
  NOR2X1   g07852(.A(new_n8041_), .B(new_n8038_), .Y(new_n8046_));
  INVX1    g07853(.A(new_n8046_), .Y(new_n8047_));
  AOI21X1  g07854(.A0(new_n8043_), .A1(new_n8047_), .B0(new_n8045_), .Y(new_n8048_));
  AND2X1   g07855(.A(new_n8047_), .B(new_n8045_), .Y(new_n8049_));
  AOI21X1  g07856(.A0(new_n8049_), .A1(new_n8043_), .B0(new_n8048_), .Y(\asquared[73] ));
  AOI21X1  g07857(.A0(new_n8047_), .A1(new_n8045_), .B0(new_n8042_), .Y(new_n8051_));
  INVX1    g07858(.A(new_n7913_), .Y(new_n8052_));
  OR2X1    g07859(.A(new_n7915_), .B(new_n8052_), .Y(new_n8053_));
  OAI21X1  g07860(.A0(new_n8037_), .A1(new_n7916_), .B0(new_n8053_), .Y(new_n8054_));
  AND2X1   g07861(.A(new_n7942_), .B(new_n7918_), .Y(new_n8055_));
  INVX1    g07862(.A(new_n8036_), .Y(new_n8056_));
  AOI21X1  g07863(.A0(new_n8056_), .A1(new_n7943_), .B0(new_n8055_), .Y(new_n8057_));
  AND2X1   g07864(.A(new_n8033_), .B(new_n7999_), .Y(new_n8058_));
  XOR2X1   g07865(.A(new_n8033_), .B(new_n7999_), .Y(new_n8059_));
  AOI21X1  g07866(.A0(new_n8059_), .A1(new_n7996_), .B0(new_n8058_), .Y(new_n8060_));
  INVX1    g07867(.A(new_n7928_), .Y(new_n8061_));
  OR2X1    g07868(.A(new_n7930_), .B(new_n8061_), .Y(new_n8062_));
  OAI21X1  g07869(.A0(new_n7941_), .A1(new_n7931_), .B0(new_n8062_), .Y(new_n8063_));
  NOR2X1   g07870(.A(new_n8032_), .B(new_n8005_), .Y(new_n8064_));
  AOI21X1  g07871(.A0(new_n8004_), .A1(new_n8001_), .B0(new_n8064_), .Y(new_n8065_));
  AND2X1   g07872(.A(new_n7871_), .B(new_n7862_), .Y(new_n8066_));
  AOI21X1  g07873(.A0(new_n8000_), .A1(new_n7819_), .B0(new_n8066_), .Y(new_n8067_));
  NAND4X1  g07874(.A(\a[41] ), .B(\a[40] ), .C(\a[33] ), .D(\a[32] ), .Y(new_n8068_));
  INVX1    g07875(.A(new_n3607_), .Y(new_n8069_));
  AND2X1   g07876(.A(\a[42] ), .B(\a[40] ), .Y(new_n8070_));
  INVX1    g07877(.A(new_n8070_), .Y(new_n8071_));
  OAI22X1  g07878(.A0(new_n8071_), .A1(new_n2673_), .B0(new_n8069_), .B1(new_n2672_), .Y(new_n8072_));
  AND2X1   g07879(.A(new_n8072_), .B(new_n8068_), .Y(new_n8073_));
  AND2X1   g07880(.A(\a[42] ), .B(\a[31] ), .Y(new_n8074_));
  INVX1    g07881(.A(new_n8074_), .Y(new_n8075_));
  AOI21X1  g07882(.A0(new_n4404_), .A1(new_n2674_), .B0(new_n8072_), .Y(new_n8076_));
  INVX1    g07883(.A(new_n8076_), .Y(new_n8077_));
  AOI22X1  g07884(.A0(\a[41] ), .A1(\a[32] ), .B0(\a[40] ), .B1(\a[33] ), .Y(new_n8078_));
  OAI22X1  g07885(.A0(new_n8078_), .A1(new_n8077_), .B0(new_n8075_), .B1(new_n8073_), .Y(new_n8079_));
  XOR2X1   g07886(.A(new_n8079_), .B(new_n8067_), .Y(new_n8080_));
  AND2X1   g07887(.A(new_n7850_), .B(new_n7833_), .Y(new_n8081_));
  AOI21X1  g07888(.A0(new_n7934_), .A1(new_n7843_), .B0(new_n8081_), .Y(new_n8082_));
  XOR2X1   g07889(.A(new_n8082_), .B(new_n8080_), .Y(new_n8083_));
  INVX1    g07890(.A(new_n8083_), .Y(new_n8084_));
  OR2X1    g07891(.A(new_n7939_), .B(new_n7935_), .Y(new_n8085_));
  AND2X1   g07892(.A(new_n7939_), .B(new_n7935_), .Y(new_n8086_));
  OAI21X1  g07893(.A0(new_n8086_), .A1(new_n7933_), .B0(new_n8085_), .Y(new_n8087_));
  XOR2X1   g07894(.A(new_n8087_), .B(new_n8084_), .Y(new_n8088_));
  XOR2X1   g07895(.A(new_n8088_), .B(new_n8065_), .Y(new_n8089_));
  INVX1    g07896(.A(new_n8089_), .Y(new_n8090_));
  XOR2X1   g07897(.A(new_n8090_), .B(new_n8063_), .Y(new_n8091_));
  XOR2X1   g07898(.A(new_n8091_), .B(new_n8060_), .Y(new_n8092_));
  XOR2X1   g07899(.A(new_n8092_), .B(new_n8057_), .Y(new_n8093_));
  NOR2X1   g07900(.A(new_n7911_), .B(new_n7909_), .Y(new_n8094_));
  AOI21X1  g07901(.A0(new_n7912_), .A1(new_n7887_), .B0(new_n8094_), .Y(new_n8095_));
  INVX1    g07902(.A(new_n7980_), .Y(new_n8096_));
  NOR2X1   g07903(.A(new_n7991_), .B(new_n7979_), .Y(new_n8097_));
  AOI21X1  g07904(.A0(new_n7989_), .A1(new_n8096_), .B0(new_n8097_), .Y(new_n8098_));
  NOR2X1   g07905(.A(new_n7807_), .B(new_n7790_), .Y(new_n8099_));
  AOI21X1  g07906(.A0(new_n7937_), .A1(new_n7936_), .B0(new_n8099_), .Y(new_n8100_));
  XOR2X1   g07907(.A(new_n8100_), .B(new_n8098_), .Y(new_n8101_));
  AND2X1   g07908(.A(new_n8021_), .B(new_n8013_), .Y(new_n8102_));
  AND2X1   g07909(.A(new_n8030_), .B(new_n8022_), .Y(new_n8103_));
  OR2X1    g07910(.A(new_n8103_), .B(new_n8102_), .Y(new_n8104_));
  XOR2X1   g07911(.A(new_n8104_), .B(new_n8101_), .Y(new_n8105_));
  INVX1    g07912(.A(new_n8105_), .Y(new_n8106_));
  OR2X1    g07913(.A(new_n7993_), .B(new_n7971_), .Y(new_n8107_));
  OAI21X1  g07914(.A0(new_n7995_), .A1(new_n7945_), .B0(new_n8107_), .Y(new_n8108_));
  XOR2X1   g07915(.A(new_n8108_), .B(new_n8106_), .Y(new_n8109_));
  INVX1    g07916(.A(new_n7954_), .Y(new_n8110_));
  OR2X1    g07917(.A(new_n7969_), .B(new_n7961_), .Y(new_n8111_));
  OAI21X1  g07918(.A0(new_n7960_), .A1(new_n8110_), .B0(new_n8111_), .Y(new_n8112_));
  NAND2X1  g07919(.A(\a[60] ), .B(\a[13] ), .Y(new_n8113_));
  XOR2X1   g07920(.A(new_n8113_), .B(new_n7959_), .Y(new_n8114_));
  XOR2X1   g07921(.A(new_n8114_), .B(new_n8029_), .Y(new_n8115_));
  INVX1    g07922(.A(new_n8115_), .Y(new_n8116_));
  XOR2X1   g07923(.A(new_n7987_), .B(new_n7976_), .Y(new_n8117_));
  XOR2X1   g07924(.A(new_n8117_), .B(new_n7968_), .Y(new_n8118_));
  XOR2X1   g07925(.A(new_n8118_), .B(new_n8116_), .Y(new_n8119_));
  XOR2X1   g07926(.A(new_n8119_), .B(new_n8112_), .Y(new_n8120_));
  INVX1    g07927(.A(new_n8120_), .Y(new_n8121_));
  XOR2X1   g07928(.A(new_n8121_), .B(new_n8109_), .Y(new_n8122_));
  INVX1    g07929(.A(new_n8122_), .Y(new_n8123_));
  XOR2X1   g07930(.A(new_n8123_), .B(new_n8095_), .Y(new_n8124_));
  AOI21X1  g07931(.A0(\a[62] ), .A1(\a[11] ), .B0(\a[37] ), .Y(new_n8125_));
  AND2X1   g07932(.A(\a[50] ), .B(\a[23] ), .Y(new_n8126_));
  INVX1    g07933(.A(new_n8126_), .Y(new_n8127_));
  AND2X1   g07934(.A(new_n3161_), .B(\a[62] ), .Y(new_n8128_));
  NOR3X1   g07935(.A(new_n8127_), .B(new_n8128_), .C(new_n8125_), .Y(new_n8129_));
  INVX1    g07936(.A(new_n8125_), .Y(new_n8130_));
  AOI21X1  g07937(.A0(new_n8126_), .A1(new_n8130_), .B0(new_n8128_), .Y(new_n8131_));
  INVX1    g07938(.A(new_n8131_), .Y(new_n8132_));
  OAI22X1  g07939(.A0(new_n8132_), .A1(new_n8125_), .B0(new_n8129_), .B1(new_n8127_), .Y(new_n8133_));
  NOR4X1   g07940(.A(new_n4835_), .B(new_n3915_), .C(new_n1185_), .D(new_n752_), .Y(new_n8134_));
  AND2X1   g07941(.A(\a[24] ), .B(\a[18] ), .Y(new_n8135_));
  AND2X1   g07942(.A(\a[55] ), .B(\a[49] ), .Y(new_n8136_));
  AOI22X1  g07943(.A0(new_n8136_), .A1(new_n8135_), .B0(new_n5240_), .B1(new_n855_), .Y(new_n8137_));
  OR2X1    g07944(.A(new_n8137_), .B(new_n8134_), .Y(new_n8138_));
  AND2X1   g07945(.A(\a[55] ), .B(\a[18] ), .Y(new_n8139_));
  INVX1    g07946(.A(new_n8134_), .Y(new_n8140_));
  AND2X1   g07947(.A(new_n8137_), .B(new_n8140_), .Y(new_n8141_));
  OAI22X1  g07948(.A0(new_n4835_), .A1(new_n752_), .B0(new_n3915_), .B1(new_n1185_), .Y(new_n8142_));
  AOI22X1  g07949(.A0(new_n8142_), .A1(new_n8141_), .B0(new_n8139_), .B1(new_n8138_), .Y(new_n8143_));
  XOR2X1   g07950(.A(new_n8143_), .B(new_n8133_), .Y(new_n8144_));
  INVX1    g07951(.A(new_n4904_), .Y(new_n8145_));
  OAI22X1  g07952(.A0(new_n8145_), .A1(new_n2135_), .B0(new_n7793_), .B1(new_n1397_), .Y(new_n8146_));
  OAI21X1  g07953(.A0(new_n7336_), .A1(new_n1794_), .B0(new_n8146_), .Y(new_n8147_));
  AND2X1   g07954(.A(\a[51] ), .B(\a[22] ), .Y(new_n8148_));
  AOI21X1  g07955(.A0(new_n5048_), .A1(new_n1236_), .B0(new_n8146_), .Y(new_n8149_));
  OAI22X1  g07956(.A0(new_n5245_), .A1(new_n934_), .B0(new_n4354_), .B1(new_n1098_), .Y(new_n8150_));
  AOI22X1  g07957(.A0(new_n8150_), .A1(new_n8149_), .B0(new_n8148_), .B1(new_n8147_), .Y(new_n8151_));
  XOR2X1   g07958(.A(new_n8151_), .B(new_n8144_), .Y(new_n8152_));
  OAI22X1  g07959(.A0(new_n5379_), .A1(new_n549_), .B0(new_n5441_), .B1(new_n571_), .Y(new_n8153_));
  INVX1    g07960(.A(new_n6119_), .Y(new_n8154_));
  INVX1    g07961(.A(new_n6120_), .Y(new_n8155_));
  OAI22X1  g07962(.A0(new_n6793_), .A1(new_n867_), .B0(new_n8155_), .B1(new_n1025_), .Y(new_n8156_));
  OAI21X1  g07963(.A0(new_n8154_), .A1(new_n1024_), .B0(new_n8156_), .Y(new_n8157_));
  AOI21X1  g07964(.A0(new_n6119_), .A1(new_n689_), .B0(new_n8156_), .Y(new_n8158_));
  AND2X1   g07965(.A(\a[59] ), .B(\a[14] ), .Y(new_n8159_));
  AOI22X1  g07966(.A0(new_n8159_), .A1(new_n8157_), .B0(new_n8158_), .B1(new_n8153_), .Y(new_n8160_));
  AND2X1   g07967(.A(\a[56] ), .B(\a[17] ), .Y(new_n8161_));
  AOI22X1  g07968(.A0(\a[47] ), .A1(\a[26] ), .B0(\a[46] ), .B1(\a[27] ), .Y(new_n8162_));
  INVX1    g07969(.A(new_n8162_), .Y(new_n8163_));
  NAND4X1  g07970(.A(\a[47] ), .B(\a[46] ), .C(\a[27] ), .D(\a[26] ), .Y(new_n8164_));
  NAND3X1  g07971(.A(new_n8163_), .B(new_n8164_), .C(new_n8161_), .Y(new_n8165_));
  AOI22X1  g07972(.A0(new_n8163_), .A1(new_n8161_), .B0(new_n3893_), .B1(new_n1995_), .Y(new_n8166_));
  AOI22X1  g07973(.A0(new_n8166_), .A1(new_n8163_), .B0(new_n8165_), .B1(new_n8161_), .Y(new_n8167_));
  XOR2X1   g07974(.A(new_n8167_), .B(new_n7952_), .Y(new_n8168_));
  XOR2X1   g07975(.A(new_n8168_), .B(new_n8160_), .Y(new_n8169_));
  XOR2X1   g07976(.A(new_n8169_), .B(new_n8152_), .Y(new_n8170_));
  NOR2X1   g07977(.A(new_n7923_), .B(new_n7920_), .Y(new_n8171_));
  AOI21X1  g07978(.A0(new_n7927_), .A1(new_n7924_), .B0(new_n8171_), .Y(new_n8172_));
  XOR2X1   g07979(.A(new_n8172_), .B(new_n8170_), .Y(new_n8173_));
  NOR2X1   g07980(.A(new_n7905_), .B(new_n7889_), .Y(new_n8174_));
  INVX1    g07981(.A(new_n7908_), .Y(new_n8175_));
  AOI21X1  g07982(.A0(new_n8175_), .A1(new_n7906_), .B0(new_n8174_), .Y(new_n8176_));
  XOR2X1   g07983(.A(new_n8019_), .B(new_n8010_), .Y(new_n8177_));
  XOR2X1   g07984(.A(new_n8177_), .B(new_n7899_), .Y(new_n8178_));
  INVX1    g07985(.A(new_n8178_), .Y(new_n8179_));
  INVX1    g07986(.A(new_n7900_), .Y(new_n8180_));
  OR2X1    g07987(.A(new_n8180_), .B(new_n7891_), .Y(new_n8181_));
  OAI21X1  g07988(.A0(new_n7904_), .A1(new_n7901_), .B0(new_n8181_), .Y(new_n8182_));
  XOR2X1   g07989(.A(new_n8182_), .B(new_n8179_), .Y(new_n8183_));
  AOI22X1  g07990(.A0(\a[63] ), .A1(\a[10] ), .B0(\a[61] ), .B1(\a[12] ), .Y(new_n8184_));
  AND2X1   g07991(.A(\a[48] ), .B(\a[25] ), .Y(new_n8185_));
  INVX1    g07992(.A(new_n8185_), .Y(new_n8186_));
  AND2X1   g07993(.A(new_n6688_), .B(new_n396_), .Y(new_n8187_));
  NOR3X1   g07994(.A(new_n8186_), .B(new_n8187_), .C(new_n8184_), .Y(new_n8188_));
  NOR2X1   g07995(.A(new_n8188_), .B(new_n8187_), .Y(new_n8189_));
  INVX1    g07996(.A(new_n8189_), .Y(new_n8190_));
  OAI22X1  g07997(.A0(new_n8190_), .A1(new_n8184_), .B0(new_n8188_), .B1(new_n8186_), .Y(new_n8191_));
  OAI22X1  g07998(.A0(new_n7642_), .A1(new_n1675_), .B0(new_n7641_), .B1(new_n2199_), .Y(new_n8192_));
  OAI21X1  g07999(.A0(new_n7353_), .A1(new_n2197_), .B0(new_n8192_), .Y(new_n8193_));
  AND2X1   g08000(.A(\a[45] ), .B(\a[28] ), .Y(new_n8194_));
  AOI21X1  g08001(.A0(new_n4992_), .A1(new_n2196_), .B0(new_n8192_), .Y(new_n8195_));
  OAI22X1  g08002(.A0(new_n5268_), .A1(new_n1803_), .B0(new_n3037_), .B1(new_n1684_), .Y(new_n8196_));
  AOI22X1  g08003(.A0(new_n8196_), .A1(new_n8195_), .B0(new_n8194_), .B1(new_n8193_), .Y(new_n8197_));
  XOR2X1   g08004(.A(new_n8197_), .B(new_n8191_), .Y(new_n8198_));
  NAND4X1  g08005(.A(\a[39] ), .B(\a[37] ), .C(\a[36] ), .D(\a[34] ), .Y(new_n8199_));
  OAI21X1  g08006(.A0(new_n3729_), .A1(new_n4915_), .B0(new_n8199_), .Y(new_n8200_));
  OAI21X1  g08007(.A0(new_n7317_), .A1(new_n5417_), .B0(new_n8200_), .Y(new_n8201_));
  AOI21X1  g08008(.A0(new_n3164_), .A1(new_n2682_), .B0(new_n8200_), .Y(new_n8202_));
  OAI22X1  g08009(.A0(new_n2519_), .A1(new_n2557_), .B0(new_n2345_), .B1(new_n2583_), .Y(new_n8203_));
  AOI22X1  g08010(.A0(new_n8203_), .A1(new_n8202_), .B0(new_n8201_), .B1(new_n3285_), .Y(new_n8204_));
  XOR2X1   g08011(.A(new_n8204_), .B(new_n8198_), .Y(new_n8205_));
  INVX1    g08012(.A(new_n8205_), .Y(new_n8206_));
  XOR2X1   g08013(.A(new_n8206_), .B(new_n8183_), .Y(new_n8207_));
  XOR2X1   g08014(.A(new_n8207_), .B(new_n8176_), .Y(new_n8208_));
  XOR2X1   g08015(.A(new_n8208_), .B(new_n8173_), .Y(new_n8209_));
  XOR2X1   g08016(.A(new_n8209_), .B(new_n8124_), .Y(new_n8210_));
  XOR2X1   g08017(.A(new_n8210_), .B(new_n8093_), .Y(new_n8211_));
  NOR2X1   g08018(.A(new_n8211_), .B(new_n8054_), .Y(new_n8212_));
  AND2X1   g08019(.A(new_n8211_), .B(new_n8054_), .Y(new_n8213_));
  OR2X1    g08020(.A(new_n8213_), .B(new_n8212_), .Y(new_n8214_));
  XOR2X1   g08021(.A(new_n8214_), .B(new_n8051_), .Y(\asquared[74] ));
  INVX1    g08022(.A(new_n8092_), .Y(new_n8216_));
  OR2X1    g08023(.A(new_n8216_), .B(new_n8057_), .Y(new_n8217_));
  OAI21X1  g08024(.A0(new_n8210_), .A1(new_n8093_), .B0(new_n8217_), .Y(new_n8218_));
  AND2X1   g08025(.A(new_n8089_), .B(new_n8063_), .Y(new_n8219_));
  INVX1    g08026(.A(new_n8219_), .Y(new_n8220_));
  OAI21X1  g08027(.A0(new_n8091_), .A1(new_n8060_), .B0(new_n8220_), .Y(new_n8221_));
  XOR2X1   g08028(.A(new_n8202_), .B(new_n8076_), .Y(new_n8222_));
  AOI22X1  g08029(.A0(new_n6795_), .A1(new_n690_), .B0(new_n6427_), .B1(new_n691_), .Y(new_n8223_));
  AOI21X1  g08030(.A0(new_n6121_), .A1(new_n689_), .B0(new_n8223_), .Y(new_n8224_));
  AND2X1   g08031(.A(\a[60] ), .B(\a[14] ), .Y(new_n8225_));
  INVX1    g08032(.A(new_n8225_), .Y(new_n8226_));
  AOI22X1  g08033(.A0(\a[59] ), .A1(\a[15] ), .B0(\a[58] ), .B1(\a[16] ), .Y(new_n8227_));
  AOI21X1  g08034(.A0(new_n6121_), .A1(new_n689_), .B0(new_n8224_), .Y(new_n8228_));
  INVX1    g08035(.A(new_n8228_), .Y(new_n8229_));
  OAI22X1  g08036(.A0(new_n8229_), .A1(new_n8227_), .B0(new_n8226_), .B1(new_n8224_), .Y(new_n8230_));
  XOR2X1   g08037(.A(new_n8230_), .B(new_n8222_), .Y(new_n8231_));
  INVX1    g08038(.A(new_n8133_), .Y(new_n8232_));
  OR2X1    g08039(.A(new_n8143_), .B(new_n8232_), .Y(new_n8233_));
  OAI21X1  g08040(.A0(new_n8151_), .A1(new_n8144_), .B0(new_n8233_), .Y(new_n8234_));
  XOR2X1   g08041(.A(new_n8234_), .B(new_n8231_), .Y(new_n8235_));
  AND2X1   g08042(.A(new_n8000_), .B(new_n7819_), .Y(new_n8236_));
  OAI21X1  g08043(.A0(new_n8236_), .A1(new_n8066_), .B0(new_n8079_), .Y(new_n8237_));
  OAI21X1  g08044(.A0(new_n8082_), .A1(new_n8080_), .B0(new_n8237_), .Y(new_n8238_));
  XOR2X1   g08045(.A(new_n8238_), .B(new_n8235_), .Y(new_n8239_));
  INVX1    g08046(.A(new_n8239_), .Y(new_n8240_));
  INVX1    g08047(.A(new_n8152_), .Y(new_n8241_));
  OR2X1    g08048(.A(new_n8169_), .B(new_n8241_), .Y(new_n8242_));
  OAI21X1  g08049(.A0(new_n8172_), .A1(new_n8170_), .B0(new_n8242_), .Y(new_n8243_));
  AND2X1   g08050(.A(new_n8182_), .B(new_n8178_), .Y(new_n8244_));
  NOR2X1   g08051(.A(new_n8206_), .B(new_n8183_), .Y(new_n8245_));
  NOR2X1   g08052(.A(new_n8245_), .B(new_n8244_), .Y(new_n8246_));
  XOR2X1   g08053(.A(new_n8246_), .B(new_n8243_), .Y(new_n8247_));
  XOR2X1   g08054(.A(new_n8247_), .B(new_n8240_), .Y(new_n8248_));
  INVX1    g08055(.A(new_n8248_), .Y(new_n8249_));
  XOR2X1   g08056(.A(new_n8249_), .B(new_n8221_), .Y(new_n8250_));
  NAND2X1  g08057(.A(new_n8087_), .B(new_n8083_), .Y(new_n8251_));
  OAI21X1  g08058(.A0(new_n8088_), .A1(new_n8065_), .B0(new_n8251_), .Y(new_n8252_));
  XOR2X1   g08059(.A(new_n8195_), .B(new_n8166_), .Y(new_n8253_));
  XOR2X1   g08060(.A(new_n8253_), .B(new_n8158_), .Y(new_n8254_));
  XOR2X1   g08061(.A(new_n8149_), .B(new_n8141_), .Y(new_n8255_));
  XOR2X1   g08062(.A(new_n8255_), .B(new_n8190_), .Y(new_n8256_));
  INVX1    g08063(.A(new_n8191_), .Y(new_n8257_));
  OR2X1    g08064(.A(new_n8197_), .B(new_n8257_), .Y(new_n8258_));
  OAI21X1  g08065(.A0(new_n8204_), .A1(new_n8198_), .B0(new_n8258_), .Y(new_n8259_));
  XOR2X1   g08066(.A(new_n8259_), .B(new_n8256_), .Y(new_n8260_));
  INVX1    g08067(.A(new_n8260_), .Y(new_n8261_));
  XOR2X1   g08068(.A(new_n8261_), .B(new_n8254_), .Y(new_n8262_));
  XOR2X1   g08069(.A(new_n8262_), .B(new_n8252_), .Y(new_n8263_));
  AND2X1   g08070(.A(\a[61] ), .B(\a[13] ), .Y(new_n8264_));
  AND2X1   g08071(.A(\a[62] ), .B(\a[12] ), .Y(new_n8265_));
  OAI22X1  g08072(.A0(new_n8265_), .A1(new_n8264_), .B0(new_n6557_), .B1(new_n587_), .Y(new_n8266_));
  XOR2X1   g08073(.A(new_n8266_), .B(new_n8132_), .Y(new_n8267_));
  NOR4X1   g08074(.A(new_n5441_), .B(new_n5268_), .C(new_n1684_), .D(new_n616_), .Y(new_n8268_));
  NAND4X1  g08075(.A(\a[45] ), .B(\a[44] ), .C(\a[30] ), .D(\a[29] ), .Y(new_n8269_));
  NAND4X1  g08076(.A(\a[57] ), .B(\a[45] ), .C(\a[29] ), .D(\a[17] ), .Y(new_n8270_));
  AOI21X1  g08077(.A0(new_n8270_), .A1(new_n8269_), .B0(new_n8268_), .Y(new_n8271_));
  NAND2X1  g08078(.A(\a[45] ), .B(\a[29] ), .Y(new_n8272_));
  OR2X1    g08079(.A(new_n8271_), .B(new_n8268_), .Y(new_n8273_));
  AOI22X1  g08080(.A0(\a[57] ), .A1(\a[17] ), .B0(\a[44] ), .B1(\a[30] ), .Y(new_n8274_));
  OAI22X1  g08081(.A0(new_n8274_), .A1(new_n8273_), .B0(new_n8272_), .B1(new_n8271_), .Y(new_n8275_));
  XOR2X1   g08082(.A(new_n8275_), .B(new_n8267_), .Y(new_n8276_));
  AND2X1   g08083(.A(new_n8019_), .B(new_n8010_), .Y(new_n8277_));
  AOI21X1  g08084(.A0(new_n8177_), .A1(new_n7899_), .B0(new_n8277_), .Y(new_n8278_));
  XOR2X1   g08085(.A(new_n8278_), .B(new_n8276_), .Y(new_n8279_));
  AOI22X1  g08086(.A0(\a[43] ), .A1(\a[31] ), .B0(\a[42] ), .B1(\a[32] ), .Y(new_n8280_));
  AND2X1   g08087(.A(\a[63] ), .B(\a[11] ), .Y(new_n8281_));
  INVX1    g08088(.A(new_n8281_), .Y(new_n8282_));
  AND2X1   g08089(.A(new_n3462_), .B(new_n2671_), .Y(new_n8283_));
  NOR3X1   g08090(.A(new_n8282_), .B(new_n8283_), .C(new_n8280_), .Y(new_n8284_));
  INVX1    g08091(.A(new_n8280_), .Y(new_n8285_));
  AOI21X1  g08092(.A0(new_n8281_), .A1(new_n8285_), .B0(new_n8283_), .Y(new_n8286_));
  INVX1    g08093(.A(new_n8286_), .Y(new_n8287_));
  OAI22X1  g08094(.A0(new_n8287_), .A1(new_n8280_), .B0(new_n8284_), .B1(new_n8282_), .Y(new_n8288_));
  AND2X1   g08095(.A(\a[41] ), .B(\a[33] ), .Y(new_n8289_));
  NOR4X1   g08096(.A(new_n6022_), .B(new_n3915_), .C(new_n1326_), .D(new_n675_), .Y(new_n8290_));
  AOI22X1  g08097(.A0(\a[56] ), .A1(\a[18] ), .B0(\a[49] ), .B1(\a[25] ), .Y(new_n8291_));
  OR4X1    g08098(.A(new_n8291_), .B(new_n8290_), .C(new_n3081_), .D(new_n1851_), .Y(new_n8292_));
  NOR3X1   g08099(.A(new_n8291_), .B(new_n8290_), .C(new_n8289_), .Y(new_n8293_));
  AOI21X1  g08100(.A0(new_n8292_), .A1(new_n8289_), .B0(new_n8293_), .Y(new_n8294_));
  XOR2X1   g08101(.A(new_n8294_), .B(new_n8288_), .Y(new_n8295_));
  INVX1    g08102(.A(new_n3893_), .Y(new_n8296_));
  INVX1    g08103(.A(new_n4272_), .Y(new_n8297_));
  AND2X1   g08104(.A(\a[48] ), .B(\a[46] ), .Y(new_n8298_));
  INVX1    g08105(.A(new_n8298_), .Y(new_n8299_));
  OAI22X1  g08106(.A0(new_n8299_), .A1(new_n3570_), .B0(new_n8297_), .B1(new_n3483_), .Y(new_n8300_));
  OAI21X1  g08107(.A0(new_n8296_), .A1(new_n1672_), .B0(new_n8300_), .Y(new_n8301_));
  AND2X1   g08108(.A(\a[48] ), .B(\a[26] ), .Y(new_n8302_));
  AOI21X1  g08109(.A0(new_n3893_), .A1(new_n1671_), .B0(new_n8300_), .Y(new_n8303_));
  OAI22X1  g08110(.A0(new_n4041_), .A1(new_n1679_), .B0(new_n3460_), .B1(new_n1431_), .Y(new_n8304_));
  AOI22X1  g08111(.A0(new_n8304_), .A1(new_n8303_), .B0(new_n8302_), .B1(new_n8301_), .Y(new_n8305_));
  XOR2X1   g08112(.A(new_n8305_), .B(new_n8295_), .Y(new_n8306_));
  OAI22X1  g08113(.A0(new_n4906_), .A1(new_n752_), .B0(new_n5245_), .B1(new_n1098_), .Y(new_n8307_));
  NAND4X1  g08114(.A(\a[55] ), .B(\a[52] ), .C(\a[22] ), .D(\a[19] ), .Y(new_n8308_));
  NAND4X1  g08115(.A(\a[53] ), .B(\a[52] ), .C(\a[22] ), .D(\a[21] ), .Y(new_n8309_));
  AOI22X1  g08116(.A0(new_n8309_), .A1(new_n8308_), .B0(new_n5236_), .B1(new_n1148_), .Y(new_n8310_));
  AOI21X1  g08117(.A0(new_n5236_), .A1(new_n1148_), .B0(new_n8310_), .Y(new_n8311_));
  NOR3X1   g08118(.A(new_n8310_), .B(new_n4354_), .C(new_n1086_), .Y(new_n8312_));
  AOI21X1  g08119(.A0(new_n8311_), .A1(new_n8307_), .B0(new_n8312_), .Y(new_n8313_));
  INVX1    g08120(.A(new_n7463_), .Y(new_n8314_));
  AOI22X1  g08121(.A0(\a[40] ), .A1(\a[34] ), .B0(\a[39] ), .B1(\a[35] ), .Y(new_n8315_));
  AND2X1   g08122(.A(new_n4077_), .B(new_n2361_), .Y(new_n8316_));
  NOR3X1   g08123(.A(new_n8315_), .B(new_n8316_), .C(new_n8314_), .Y(new_n8317_));
  INVX1    g08124(.A(new_n8315_), .Y(new_n8318_));
  AOI21X1  g08125(.A0(new_n8318_), .A1(new_n7463_), .B0(new_n8316_), .Y(new_n8319_));
  INVX1    g08126(.A(new_n8319_), .Y(new_n8320_));
  OAI22X1  g08127(.A0(new_n8320_), .A1(new_n8315_), .B0(new_n8317_), .B1(new_n8314_), .Y(new_n8321_));
  XOR2X1   g08128(.A(new_n8321_), .B(new_n8313_), .Y(new_n8322_));
  AOI22X1  g08129(.A0(\a[51] ), .A1(\a[23] ), .B0(\a[50] ), .B1(\a[24] ), .Y(new_n8323_));
  INVX1    g08130(.A(new_n8323_), .Y(new_n8324_));
  NAND4X1  g08131(.A(\a[51] ), .B(\a[50] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n8325_));
  AOI21X1  g08132(.A0(new_n8324_), .A1(new_n8325_), .B0(new_n7316_), .Y(new_n8326_));
  AOI22X1  g08133(.A0(new_n8324_), .A1(new_n2484_), .B0(new_n4484_), .B1(new_n1219_), .Y(new_n8327_));
  AOI21X1  g08134(.A0(new_n8327_), .A1(new_n8324_), .B0(new_n8326_), .Y(new_n8328_));
  XOR2X1   g08135(.A(new_n8328_), .B(new_n8322_), .Y(new_n8329_));
  INVX1    g08136(.A(new_n8329_), .Y(new_n8330_));
  XOR2X1   g08137(.A(new_n8330_), .B(new_n8306_), .Y(new_n8331_));
  XOR2X1   g08138(.A(new_n8331_), .B(new_n8279_), .Y(new_n8332_));
  XOR2X1   g08139(.A(new_n8332_), .B(new_n8263_), .Y(new_n8333_));
  INVX1    g08140(.A(new_n8333_), .Y(new_n8334_));
  XOR2X1   g08141(.A(new_n8334_), .B(new_n8250_), .Y(new_n8335_));
  INVX1    g08142(.A(new_n8335_), .Y(new_n8336_));
  AND2X1   g08143(.A(new_n8123_), .B(new_n8095_), .Y(new_n8337_));
  OR2X1    g08144(.A(new_n8123_), .B(new_n8095_), .Y(new_n8338_));
  OAI21X1  g08145(.A0(new_n8209_), .A1(new_n8337_), .B0(new_n8338_), .Y(new_n8339_));
  INVX1    g08146(.A(new_n8207_), .Y(new_n8340_));
  NOR2X1   g08147(.A(new_n8340_), .B(new_n8176_), .Y(new_n8341_));
  INVX1    g08148(.A(new_n8208_), .Y(new_n8342_));
  AOI21X1  g08149(.A0(new_n8342_), .A1(new_n8173_), .B0(new_n8341_), .Y(new_n8343_));
  NAND2X1  g08150(.A(new_n8108_), .B(new_n8105_), .Y(new_n8344_));
  OAI21X1  g08151(.A0(new_n8121_), .A1(new_n8109_), .B0(new_n8344_), .Y(new_n8345_));
  NOR2X1   g08152(.A(new_n7987_), .B(new_n7976_), .Y(new_n8346_));
  AOI21X1  g08153(.A0(new_n8117_), .A1(new_n7967_), .B0(new_n8346_), .Y(new_n8347_));
  NOR2X1   g08154(.A(new_n8113_), .B(new_n7959_), .Y(new_n8348_));
  AOI21X1  g08155(.A0(new_n8114_), .A1(new_n8029_), .B0(new_n8348_), .Y(new_n8349_));
  XOR2X1   g08156(.A(new_n8349_), .B(new_n8347_), .Y(new_n8350_));
  INVX1    g08157(.A(new_n8350_), .Y(new_n8351_));
  OR2X1    g08158(.A(new_n8167_), .B(new_n7952_), .Y(new_n8352_));
  AND2X1   g08159(.A(new_n8167_), .B(new_n7952_), .Y(new_n8353_));
  OAI21X1  g08160(.A0(new_n8353_), .A1(new_n8160_), .B0(new_n8352_), .Y(new_n8354_));
  XOR2X1   g08161(.A(new_n8354_), .B(new_n8351_), .Y(new_n8355_));
  NOR2X1   g08162(.A(new_n8118_), .B(new_n8116_), .Y(new_n8356_));
  AOI21X1  g08163(.A0(new_n8119_), .A1(new_n8112_), .B0(new_n8356_), .Y(new_n8357_));
  NOR2X1   g08164(.A(new_n8100_), .B(new_n8098_), .Y(new_n8358_));
  AOI21X1  g08165(.A0(new_n8104_), .A1(new_n8101_), .B0(new_n8358_), .Y(new_n8359_));
  XOR2X1   g08166(.A(new_n8359_), .B(new_n8357_), .Y(new_n8360_));
  INVX1    g08167(.A(new_n8360_), .Y(new_n8361_));
  XOR2X1   g08168(.A(new_n8361_), .B(new_n8355_), .Y(new_n8362_));
  INVX1    g08169(.A(new_n8362_), .Y(new_n8363_));
  XOR2X1   g08170(.A(new_n8363_), .B(new_n8345_), .Y(new_n8364_));
  XOR2X1   g08171(.A(new_n8364_), .B(new_n8343_), .Y(new_n8365_));
  XOR2X1   g08172(.A(new_n8365_), .B(new_n8339_), .Y(new_n8366_));
  XOR2X1   g08173(.A(new_n8366_), .B(new_n8336_), .Y(new_n8367_));
  XOR2X1   g08174(.A(new_n8367_), .B(new_n8218_), .Y(new_n8368_));
  INVX1    g08175(.A(new_n8213_), .Y(new_n8369_));
  OAI21X1  g08176(.A0(new_n8212_), .A1(new_n8051_), .B0(new_n8369_), .Y(new_n8370_));
  XOR2X1   g08177(.A(new_n8370_), .B(new_n8368_), .Y(\asquared[75] ));
  AND2X1   g08178(.A(new_n8365_), .B(new_n8339_), .Y(new_n8372_));
  AOI21X1  g08179(.A0(new_n8366_), .A1(new_n8336_), .B0(new_n8372_), .Y(new_n8373_));
  NAND2X1  g08180(.A(new_n8362_), .B(new_n8345_), .Y(new_n8374_));
  OAI21X1  g08181(.A0(new_n8364_), .A1(new_n8343_), .B0(new_n8374_), .Y(new_n8375_));
  NOR2X1   g08182(.A(new_n8202_), .B(new_n8076_), .Y(new_n8376_));
  AOI21X1  g08183(.A0(new_n8230_), .A1(new_n8222_), .B0(new_n8376_), .Y(new_n8377_));
  NOR2X1   g08184(.A(new_n8149_), .B(new_n8141_), .Y(new_n8378_));
  AOI21X1  g08185(.A0(new_n8255_), .A1(new_n8190_), .B0(new_n8378_), .Y(new_n8379_));
  XOR2X1   g08186(.A(new_n8379_), .B(new_n8377_), .Y(new_n8380_));
  INVX1    g08187(.A(new_n8158_), .Y(new_n8381_));
  NOR2X1   g08188(.A(new_n8195_), .B(new_n8166_), .Y(new_n8382_));
  AOI21X1  g08189(.A0(new_n8253_), .A1(new_n8381_), .B0(new_n8382_), .Y(new_n8383_));
  XOR2X1   g08190(.A(new_n8383_), .B(new_n8380_), .Y(new_n8384_));
  XOR2X1   g08191(.A(new_n8329_), .B(new_n8306_), .Y(new_n8385_));
  AND2X1   g08192(.A(new_n8329_), .B(new_n8306_), .Y(new_n8386_));
  AOI21X1  g08193(.A0(new_n8385_), .A1(new_n8279_), .B0(new_n8386_), .Y(new_n8387_));
  XOR2X1   g08194(.A(new_n8387_), .B(new_n8384_), .Y(new_n8388_));
  INVX1    g08195(.A(new_n8267_), .Y(new_n8389_));
  NAND2X1  g08196(.A(new_n8275_), .B(new_n8389_), .Y(new_n8390_));
  OAI21X1  g08197(.A0(new_n8278_), .A1(new_n8276_), .B0(new_n8390_), .Y(new_n8391_));
  XOR2X1   g08198(.A(new_n8327_), .B(new_n8319_), .Y(new_n8392_));
  XOR2X1   g08199(.A(new_n8392_), .B(new_n8311_), .Y(new_n8393_));
  NOR3X1   g08200(.A(new_n8291_), .B(new_n3081_), .C(new_n1851_), .Y(new_n8394_));
  NOR2X1   g08201(.A(new_n8394_), .B(new_n8290_), .Y(new_n8395_));
  XOR2X1   g08202(.A(new_n8395_), .B(new_n8286_), .Y(new_n8396_));
  OAI22X1  g08203(.A0(new_n8266_), .A1(new_n8131_), .B0(new_n6557_), .B1(new_n587_), .Y(new_n8397_));
  INVX1    g08204(.A(new_n8397_), .Y(new_n8398_));
  XOR2X1   g08205(.A(new_n8398_), .B(new_n8396_), .Y(new_n8399_));
  XOR2X1   g08206(.A(new_n8399_), .B(new_n8393_), .Y(new_n8400_));
  XOR2X1   g08207(.A(new_n8400_), .B(new_n8391_), .Y(new_n8401_));
  XOR2X1   g08208(.A(new_n8401_), .B(new_n8388_), .Y(new_n8402_));
  XOR2X1   g08209(.A(new_n8402_), .B(new_n8375_), .Y(new_n8403_));
  INVX1    g08210(.A(new_n8403_), .Y(new_n8404_));
  NOR2X1   g08211(.A(new_n8359_), .B(new_n8357_), .Y(new_n8405_));
  INVX1    g08212(.A(new_n8405_), .Y(new_n8406_));
  OAI21X1  g08213(.A0(new_n8361_), .A1(new_n8355_), .B0(new_n8406_), .Y(new_n8407_));
  INVX1    g08214(.A(new_n8303_), .Y(new_n8408_));
  XOR2X1   g08215(.A(new_n8408_), .B(new_n8273_), .Y(new_n8409_));
  XOR2X1   g08216(.A(new_n8409_), .B(new_n8229_), .Y(new_n8410_));
  AND2X1   g08217(.A(new_n8311_), .B(new_n8307_), .Y(new_n8411_));
  OAI21X1  g08218(.A0(new_n8312_), .A1(new_n8411_), .B0(new_n8321_), .Y(new_n8412_));
  OAI21X1  g08219(.A0(new_n8328_), .A1(new_n8322_), .B0(new_n8412_), .Y(new_n8413_));
  AND2X1   g08220(.A(new_n8292_), .B(new_n8289_), .Y(new_n8414_));
  OAI21X1  g08221(.A0(new_n8293_), .A1(new_n8414_), .B0(new_n8288_), .Y(new_n8415_));
  OR2X1    g08222(.A(new_n8305_), .B(new_n8295_), .Y(new_n8416_));
  AND2X1   g08223(.A(new_n8416_), .B(new_n8415_), .Y(new_n8417_));
  INVX1    g08224(.A(new_n8417_), .Y(new_n8418_));
  XOR2X1   g08225(.A(new_n8418_), .B(new_n8413_), .Y(new_n8419_));
  XOR2X1   g08226(.A(new_n8419_), .B(new_n8410_), .Y(new_n8420_));
  XOR2X1   g08227(.A(new_n8420_), .B(new_n8407_), .Y(new_n8421_));
  AOI22X1  g08228(.A0(\a[63] ), .A1(\a[12] ), .B0(\a[56] ), .B1(\a[19] ), .Y(new_n8422_));
  AND2X1   g08229(.A(\a[45] ), .B(\a[30] ), .Y(new_n8423_));
  INVX1    g08230(.A(new_n8423_), .Y(new_n8424_));
  AND2X1   g08231(.A(\a[63] ), .B(\a[19] ), .Y(new_n8425_));
  AND2X1   g08232(.A(new_n8425_), .B(new_n7325_), .Y(new_n8426_));
  NOR3X1   g08233(.A(new_n8424_), .B(new_n8426_), .C(new_n8422_), .Y(new_n8427_));
  NOR2X1   g08234(.A(new_n8427_), .B(new_n8426_), .Y(new_n8428_));
  INVX1    g08235(.A(new_n8428_), .Y(new_n8429_));
  OAI22X1  g08236(.A0(new_n8429_), .A1(new_n8422_), .B0(new_n8427_), .B1(new_n8424_), .Y(new_n8430_));
  AND2X1   g08237(.A(\a[52] ), .B(\a[23] ), .Y(new_n8431_));
  AOI22X1  g08238(.A0(\a[40] ), .A1(\a[35] ), .B0(\a[39] ), .B1(\a[36] ), .Y(new_n8432_));
  INVX1    g08239(.A(new_n8432_), .Y(new_n8433_));
  NAND4X1  g08240(.A(\a[40] ), .B(\a[39] ), .C(\a[36] ), .D(\a[35] ), .Y(new_n8434_));
  NAND3X1  g08241(.A(new_n8433_), .B(new_n8434_), .C(new_n8431_), .Y(new_n8435_));
  AOI22X1  g08242(.A0(new_n8433_), .A1(new_n8431_), .B0(new_n4077_), .B1(new_n2682_), .Y(new_n8436_));
  AOI22X1  g08243(.A0(new_n8436_), .A1(new_n8433_), .B0(new_n8435_), .B1(new_n8431_), .Y(new_n8437_));
  XOR2X1   g08244(.A(new_n8437_), .B(new_n8430_), .Y(new_n8438_));
  NAND3X1  g08245(.A(\a[62] ), .B(\a[38] ), .C(\a[13] ), .Y(new_n8439_));
  NOR3X1   g08246(.A(new_n8439_), .B(new_n2519_), .C(new_n2345_), .Y(new_n8440_));
  AND2X1   g08247(.A(new_n8439_), .B(new_n7317_), .Y(new_n8441_));
  OAI21X1  g08248(.A0(new_n6606_), .A1(new_n591_), .B0(new_n2519_), .Y(new_n8442_));
  AOI21X1  g08249(.A0(new_n8442_), .A1(new_n8441_), .B0(new_n8440_), .Y(new_n8443_));
  XOR2X1   g08250(.A(new_n8443_), .B(new_n8438_), .Y(new_n8444_));
  INVX1    g08251(.A(new_n8444_), .Y(new_n8445_));
  NOR2X1   g08252(.A(new_n8349_), .B(new_n8347_), .Y(new_n8446_));
  AOI21X1  g08253(.A0(new_n8354_), .A1(new_n8350_), .B0(new_n8446_), .Y(new_n8447_));
  XOR2X1   g08254(.A(new_n8447_), .B(new_n8445_), .Y(new_n8448_));
  INVX1    g08255(.A(new_n8448_), .Y(new_n8449_));
  NAND4X1  g08256(.A(\a[61] ), .B(\a[59] ), .C(\a[16] ), .D(\a[14] ), .Y(new_n8450_));
  NAND4X1  g08257(.A(\a[61] ), .B(\a[60] ), .C(\a[15] ), .D(\a[14] ), .Y(new_n8451_));
  AOI22X1  g08258(.A0(new_n8451_), .A1(new_n8450_), .B0(new_n6427_), .B1(new_n689_), .Y(new_n8452_));
  NAND4X1  g08259(.A(\a[60] ), .B(\a[59] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n8453_));
  NAND3X1  g08260(.A(new_n8451_), .B(new_n8450_), .C(new_n8453_), .Y(new_n8454_));
  AOI22X1  g08261(.A0(\a[60] ), .A1(\a[15] ), .B0(\a[59] ), .B1(\a[16] ), .Y(new_n8455_));
  NAND2X1  g08262(.A(\a[61] ), .B(\a[14] ), .Y(new_n8456_));
  OAI22X1  g08263(.A0(new_n8456_), .A1(new_n8452_), .B0(new_n8455_), .B1(new_n8454_), .Y(new_n8457_));
  NAND2X1  g08264(.A(\a[58] ), .B(\a[17] ), .Y(new_n8458_));
  NOR4X1   g08265(.A(new_n5441_), .B(new_n3915_), .C(new_n1263_), .D(new_n675_), .Y(new_n8459_));
  NAND4X1  g08266(.A(\a[58] ), .B(\a[49] ), .C(\a[26] ), .D(\a[17] ), .Y(new_n8460_));
  NAND4X1  g08267(.A(\a[58] ), .B(\a[57] ), .C(\a[18] ), .D(\a[17] ), .Y(new_n8461_));
  AOI21X1  g08268(.A0(new_n8461_), .A1(new_n8460_), .B0(new_n8459_), .Y(new_n8462_));
  OR2X1    g08269(.A(new_n8462_), .B(new_n8459_), .Y(new_n8463_));
  AOI22X1  g08270(.A0(\a[57] ), .A1(\a[18] ), .B0(\a[49] ), .B1(\a[26] ), .Y(new_n8464_));
  OAI22X1  g08271(.A0(new_n8464_), .A1(new_n8463_), .B0(new_n8462_), .B1(new_n8458_), .Y(new_n8465_));
  XOR2X1   g08272(.A(new_n8465_), .B(new_n8457_), .Y(new_n8466_));
  AOI22X1  g08273(.A0(new_n8298_), .A1(new_n1484_), .B0(new_n4272_), .B1(new_n1671_), .Y(new_n8467_));
  AOI21X1  g08274(.A0(new_n3893_), .A1(new_n1674_), .B0(new_n8467_), .Y(new_n8468_));
  AND2X1   g08275(.A(\a[48] ), .B(\a[27] ), .Y(new_n8469_));
  INVX1    g08276(.A(new_n8469_), .Y(new_n8470_));
  OAI22X1  g08277(.A0(new_n8299_), .A1(new_n1673_), .B0(new_n8297_), .B1(new_n1672_), .Y(new_n8471_));
  AOI21X1  g08278(.A0(new_n3893_), .A1(new_n1674_), .B0(new_n8471_), .Y(new_n8472_));
  INVX1    g08279(.A(new_n8472_), .Y(new_n8473_));
  AOI22X1  g08280(.A0(\a[47] ), .A1(\a[28] ), .B0(\a[46] ), .B1(\a[29] ), .Y(new_n8474_));
  OAI22X1  g08281(.A0(new_n8474_), .A1(new_n8473_), .B0(new_n8470_), .B1(new_n8468_), .Y(new_n8475_));
  INVX1    g08282(.A(new_n8475_), .Y(new_n8476_));
  XOR2X1   g08283(.A(new_n8476_), .B(new_n8466_), .Y(new_n8477_));
  XOR2X1   g08284(.A(new_n8477_), .B(new_n8449_), .Y(new_n8478_));
  INVX1    g08285(.A(new_n8478_), .Y(new_n8479_));
  XOR2X1   g08286(.A(new_n8479_), .B(new_n8421_), .Y(new_n8480_));
  XOR2X1   g08287(.A(new_n8480_), .B(new_n8404_), .Y(new_n8481_));
  AND2X1   g08288(.A(new_n8234_), .B(new_n8231_), .Y(new_n8482_));
  AOI21X1  g08289(.A0(new_n8238_), .A1(new_n8235_), .B0(new_n8482_), .Y(new_n8483_));
  AOI22X1  g08290(.A0(\a[55] ), .A1(\a[20] ), .B0(\a[50] ), .B1(\a[25] ), .Y(new_n8484_));
  AND2X1   g08291(.A(\a[41] ), .B(\a[34] ), .Y(new_n8485_));
  INVX1    g08292(.A(new_n8485_), .Y(new_n8486_));
  NOR4X1   g08293(.A(new_n4906_), .B(new_n4983_), .C(new_n1326_), .D(new_n934_), .Y(new_n8487_));
  NOR3X1   g08294(.A(new_n8486_), .B(new_n8487_), .C(new_n8484_), .Y(new_n8488_));
  INVX1    g08295(.A(new_n8484_), .Y(new_n8489_));
  AOI21X1  g08296(.A0(new_n8485_), .A1(new_n8489_), .B0(new_n8487_), .Y(new_n8490_));
  INVX1    g08297(.A(new_n8490_), .Y(new_n8491_));
  OAI22X1  g08298(.A0(new_n8491_), .A1(new_n8484_), .B0(new_n8488_), .B1(new_n8486_), .Y(new_n8492_));
  OAI22X1  g08299(.A0(new_n7353_), .A1(new_n2672_), .B0(new_n3212_), .B1(new_n2673_), .Y(new_n8493_));
  OAI21X1  g08300(.A0(new_n6502_), .A1(new_n2675_), .B0(new_n8493_), .Y(new_n8494_));
  AND2X1   g08301(.A(\a[44] ), .B(\a[31] ), .Y(new_n8495_));
  OAI22X1  g08302(.A0(new_n3037_), .A1(new_n2219_), .B0(new_n3096_), .B1(new_n1851_), .Y(new_n8496_));
  AOI21X1  g08303(.A0(new_n3462_), .A1(new_n2674_), .B0(new_n8493_), .Y(new_n8497_));
  AOI22X1  g08304(.A0(new_n8497_), .A1(new_n8496_), .B0(new_n8495_), .B1(new_n8494_), .Y(new_n8498_));
  XOR2X1   g08305(.A(new_n8498_), .B(new_n8492_), .Y(new_n8499_));
  NAND4X1  g08306(.A(\a[54] ), .B(\a[53] ), .C(\a[22] ), .D(\a[21] ), .Y(new_n8500_));
  NAND4X1  g08307(.A(\a[54] ), .B(\a[51] ), .C(\a[24] ), .D(\a[21] ), .Y(new_n8501_));
  AOI22X1  g08308(.A0(new_n8501_), .A1(new_n8500_), .B0(new_n4904_), .B1(new_n1530_), .Y(new_n8502_));
  NOR3X1   g08309(.A(new_n8502_), .B(new_n4835_), .C(new_n1098_), .Y(new_n8503_));
  AOI21X1  g08310(.A0(new_n4904_), .A1(new_n1530_), .B0(new_n8502_), .Y(new_n8504_));
  OAI22X1  g08311(.A0(new_n5245_), .A1(new_n1086_), .B0(new_n4349_), .B1(new_n1185_), .Y(new_n8505_));
  AOI21X1  g08312(.A0(new_n8505_), .A1(new_n8504_), .B0(new_n8503_), .Y(new_n8506_));
  XOR2X1   g08313(.A(new_n8506_), .B(new_n8499_), .Y(new_n8507_));
  NAND2X1  g08314(.A(new_n8259_), .B(new_n8256_), .Y(new_n8508_));
  OAI21X1  g08315(.A0(new_n8261_), .A1(new_n8254_), .B0(new_n8508_), .Y(new_n8509_));
  XOR2X1   g08316(.A(new_n8509_), .B(new_n8507_), .Y(new_n8510_));
  XOR2X1   g08317(.A(new_n8510_), .B(new_n8483_), .Y(new_n8511_));
  OAI21X1  g08318(.A0(new_n8245_), .A1(new_n8244_), .B0(new_n8243_), .Y(new_n8512_));
  OAI21X1  g08319(.A0(new_n8247_), .A1(new_n8240_), .B0(new_n8512_), .Y(new_n8513_));
  XOR2X1   g08320(.A(new_n8513_), .B(new_n8511_), .Y(new_n8514_));
  INVX1    g08321(.A(new_n8514_), .Y(new_n8515_));
  AND2X1   g08322(.A(new_n8262_), .B(new_n8252_), .Y(new_n8516_));
  INVX1    g08323(.A(new_n8332_), .Y(new_n8517_));
  AOI21X1  g08324(.A0(new_n8517_), .A1(new_n8263_), .B0(new_n8516_), .Y(new_n8518_));
  XOR2X1   g08325(.A(new_n8518_), .B(new_n8515_), .Y(new_n8519_));
  NOR2X1   g08326(.A(new_n8333_), .B(new_n8250_), .Y(new_n8520_));
  AOI21X1  g08327(.A0(new_n8248_), .A1(new_n8221_), .B0(new_n8520_), .Y(new_n8521_));
  XOR2X1   g08328(.A(new_n8521_), .B(new_n8519_), .Y(new_n8522_));
  XOR2X1   g08329(.A(new_n8522_), .B(new_n8481_), .Y(new_n8523_));
  XOR2X1   g08330(.A(new_n8523_), .B(new_n8373_), .Y(new_n8524_));
  OR2X1    g08331(.A(new_n8367_), .B(new_n8218_), .Y(new_n8525_));
  AND2X1   g08332(.A(new_n8367_), .B(new_n8218_), .Y(new_n8526_));
  AOI21X1  g08333(.A0(new_n8370_), .A1(new_n8525_), .B0(new_n8526_), .Y(new_n8527_));
  XOR2X1   g08334(.A(new_n8527_), .B(new_n8524_), .Y(\asquared[76] ));
  INVX1    g08335(.A(new_n8523_), .Y(new_n8529_));
  OR2X1    g08336(.A(new_n8529_), .B(new_n8373_), .Y(new_n8530_));
  AND2X1   g08337(.A(new_n8529_), .B(new_n8373_), .Y(new_n8531_));
  OAI21X1  g08338(.A0(new_n8527_), .A1(new_n8531_), .B0(new_n8530_), .Y(new_n8532_));
  NOR2X1   g08339(.A(new_n8521_), .B(new_n8519_), .Y(new_n8533_));
  AOI21X1  g08340(.A0(new_n8522_), .A1(new_n8481_), .B0(new_n8533_), .Y(new_n8534_));
  AND2X1   g08341(.A(new_n8402_), .B(new_n8375_), .Y(new_n8535_));
  INVX1    g08342(.A(new_n8535_), .Y(new_n8536_));
  OAI21X1  g08343(.A0(new_n8480_), .A1(new_n8404_), .B0(new_n8536_), .Y(new_n8537_));
  NAND2X1  g08344(.A(new_n8420_), .B(new_n8407_), .Y(new_n8538_));
  NOR2X1   g08345(.A(new_n8420_), .B(new_n8407_), .Y(new_n8539_));
  OAI21X1  g08346(.A0(new_n8479_), .A1(new_n8539_), .B0(new_n8538_), .Y(new_n8540_));
  NOR2X1   g08347(.A(new_n8387_), .B(new_n8384_), .Y(new_n8541_));
  AOI21X1  g08348(.A0(new_n8401_), .A1(new_n8388_), .B0(new_n8541_), .Y(new_n8542_));
  NOR2X1   g08349(.A(new_n8399_), .B(new_n8393_), .Y(new_n8543_));
  AOI21X1  g08350(.A0(new_n8400_), .A1(new_n8391_), .B0(new_n8543_), .Y(new_n8544_));
  AOI22X1  g08351(.A0(\a[45] ), .A1(\a[31] ), .B0(\a[44] ), .B1(\a[32] ), .Y(new_n8545_));
  AND2X1   g08352(.A(\a[63] ), .B(\a[13] ), .Y(new_n8546_));
  INVX1    g08353(.A(new_n8546_), .Y(new_n8547_));
  AND2X1   g08354(.A(new_n3918_), .B(new_n2671_), .Y(new_n8548_));
  NOR3X1   g08355(.A(new_n8547_), .B(new_n8548_), .C(new_n8545_), .Y(new_n8549_));
  NOR2X1   g08356(.A(new_n8549_), .B(new_n8548_), .Y(new_n8550_));
  INVX1    g08357(.A(new_n8550_), .Y(new_n8551_));
  OAI22X1  g08358(.A0(new_n8551_), .A1(new_n8545_), .B0(new_n8549_), .B1(new_n8547_), .Y(new_n8552_));
  NOR4X1   g08359(.A(new_n5441_), .B(new_n5245_), .C(new_n1216_), .D(new_n752_), .Y(new_n8553_));
  AOI22X1  g08360(.A0(\a[57] ), .A1(\a[19] ), .B0(\a[53] ), .B1(\a[23] ), .Y(new_n8554_));
  OR4X1    g08361(.A(new_n8554_), .B(new_n8553_), .C(new_n3037_), .D(new_n1851_), .Y(new_n8555_));
  NOR3X1   g08362(.A(new_n8554_), .B(new_n8553_), .C(new_n3744_), .Y(new_n8556_));
  AOI21X1  g08363(.A0(new_n8555_), .A1(new_n3744_), .B0(new_n8556_), .Y(new_n8557_));
  XOR2X1   g08364(.A(new_n8557_), .B(new_n8552_), .Y(new_n8558_));
  INVX1    g08365(.A(new_n5042_), .Y(new_n8559_));
  INVX1    g08366(.A(new_n6237_), .Y(new_n8560_));
  OAI22X1  g08367(.A0(new_n8560_), .A1(new_n1794_), .B0(new_n8559_), .B1(new_n2135_), .Y(new_n8561_));
  OAI21X1  g08368(.A0(new_n5241_), .A1(new_n1397_), .B0(new_n8561_), .Y(new_n8562_));
  AOI21X1  g08369(.A0(new_n5240_), .A1(new_n1154_), .B0(new_n8561_), .Y(new_n8563_));
  OAI22X1  g08370(.A0(new_n4906_), .A1(new_n1098_), .B0(new_n4835_), .B1(new_n1086_), .Y(new_n8564_));
  AOI22X1  g08371(.A0(new_n8564_), .A1(new_n8563_), .B0(new_n8562_), .B1(new_n7052_), .Y(new_n8565_));
  XOR2X1   g08372(.A(new_n8565_), .B(new_n8558_), .Y(new_n8566_));
  NAND2X1  g08373(.A(new_n8418_), .B(new_n8413_), .Y(new_n8567_));
  NAND2X1  g08374(.A(new_n8419_), .B(new_n8410_), .Y(new_n8568_));
  NAND2X1  g08375(.A(new_n8568_), .B(new_n8567_), .Y(new_n8569_));
  XOR2X1   g08376(.A(new_n8569_), .B(new_n8566_), .Y(new_n8570_));
  XOR2X1   g08377(.A(new_n8570_), .B(new_n8544_), .Y(new_n8571_));
  XOR2X1   g08378(.A(new_n8571_), .B(new_n8542_), .Y(new_n8572_));
  XOR2X1   g08379(.A(new_n8572_), .B(new_n8540_), .Y(new_n8573_));
  XOR2X1   g08380(.A(new_n8573_), .B(new_n8537_), .Y(new_n8574_));
  INVX1    g08381(.A(new_n8574_), .Y(new_n8575_));
  NAND2X1  g08382(.A(new_n8397_), .B(new_n8396_), .Y(new_n8576_));
  OAI21X1  g08383(.A0(new_n8395_), .A1(new_n8286_), .B0(new_n8576_), .Y(new_n8577_));
  AND2X1   g08384(.A(new_n8408_), .B(new_n8273_), .Y(new_n8578_));
  AOI21X1  g08385(.A0(new_n8409_), .A1(new_n8229_), .B0(new_n8578_), .Y(new_n8579_));
  XOR2X1   g08386(.A(new_n8579_), .B(new_n8577_), .Y(new_n8580_));
  INVX1    g08387(.A(new_n8311_), .Y(new_n8581_));
  NOR2X1   g08388(.A(new_n8327_), .B(new_n8319_), .Y(new_n8582_));
  AOI21X1  g08389(.A0(new_n8392_), .A1(new_n8581_), .B0(new_n8582_), .Y(new_n8583_));
  XOR2X1   g08390(.A(new_n8583_), .B(new_n8580_), .Y(new_n8584_));
  OR2X1    g08391(.A(new_n8447_), .B(new_n8445_), .Y(new_n8585_));
  OAI21X1  g08392(.A0(new_n8477_), .A1(new_n8449_), .B0(new_n8585_), .Y(new_n8586_));
  XOR2X1   g08393(.A(new_n8586_), .B(new_n8584_), .Y(new_n8587_));
  XOR2X1   g08394(.A(new_n8490_), .B(new_n8472_), .Y(new_n8588_));
  XOR2X1   g08395(.A(new_n8588_), .B(new_n8429_), .Y(new_n8589_));
  INVX1    g08396(.A(new_n8492_), .Y(new_n8590_));
  OR2X1    g08397(.A(new_n8498_), .B(new_n8590_), .Y(new_n8591_));
  OAI21X1  g08398(.A0(new_n8506_), .A1(new_n8499_), .B0(new_n8591_), .Y(new_n8592_));
  NAND2X1  g08399(.A(\a[62] ), .B(\a[14] ), .Y(new_n8593_));
  AND2X1   g08400(.A(new_n8593_), .B(new_n8441_), .Y(new_n8594_));
  AOI21X1  g08401(.A0(new_n8439_), .A1(new_n7317_), .B0(new_n8593_), .Y(new_n8595_));
  NOR3X1   g08402(.A(new_n8595_), .B(new_n8594_), .C(new_n8436_), .Y(new_n8596_));
  OR2X1    g08403(.A(new_n8596_), .B(new_n8595_), .Y(new_n8597_));
  OAI22X1  g08404(.A0(new_n8597_), .A1(new_n8594_), .B0(new_n8596_), .B1(new_n8436_), .Y(new_n8598_));
  XOR2X1   g08405(.A(new_n8598_), .B(new_n8592_), .Y(new_n8599_));
  XOR2X1   g08406(.A(new_n8599_), .B(new_n8589_), .Y(new_n8600_));
  XOR2X1   g08407(.A(new_n8600_), .B(new_n8587_), .Y(new_n8601_));
  INVX1    g08408(.A(new_n8511_), .Y(new_n8602_));
  NOR2X1   g08409(.A(new_n8518_), .B(new_n8514_), .Y(new_n8603_));
  AOI21X1  g08410(.A0(new_n8513_), .A1(new_n8602_), .B0(new_n8603_), .Y(new_n8604_));
  XOR2X1   g08411(.A(new_n8604_), .B(new_n8601_), .Y(new_n8605_));
  NAND2X1  g08412(.A(new_n8509_), .B(new_n8507_), .Y(new_n8606_));
  INVX1    g08413(.A(new_n8510_), .Y(new_n8607_));
  OAI21X1  g08414(.A0(new_n8607_), .A1(new_n8483_), .B0(new_n8606_), .Y(new_n8608_));
  XOR2X1   g08415(.A(new_n8463_), .B(new_n8454_), .Y(new_n8609_));
  XOR2X1   g08416(.A(new_n8609_), .B(new_n8497_), .Y(new_n8610_));
  AND2X1   g08417(.A(new_n8465_), .B(new_n8457_), .Y(new_n8611_));
  AND2X1   g08418(.A(new_n8475_), .B(new_n8466_), .Y(new_n8612_));
  OR2X1    g08419(.A(new_n8612_), .B(new_n8611_), .Y(new_n8613_));
  INVX1    g08420(.A(new_n8430_), .Y(new_n8614_));
  OR2X1    g08421(.A(new_n8437_), .B(new_n8614_), .Y(new_n8615_));
  OR2X1    g08422(.A(new_n8443_), .B(new_n8438_), .Y(new_n8616_));
  AND2X1   g08423(.A(new_n8616_), .B(new_n8615_), .Y(new_n8617_));
  INVX1    g08424(.A(new_n8617_), .Y(new_n8618_));
  XOR2X1   g08425(.A(new_n8618_), .B(new_n8613_), .Y(new_n8619_));
  INVX1    g08426(.A(new_n8619_), .Y(new_n8620_));
  XOR2X1   g08427(.A(new_n8620_), .B(new_n8610_), .Y(new_n8621_));
  XOR2X1   g08428(.A(new_n8621_), .B(new_n8608_), .Y(new_n8622_));
  INVX1    g08429(.A(new_n8622_), .Y(new_n8623_));
  NAND4X1  g08430(.A(\a[48] ), .B(\a[46] ), .C(\a[30] ), .D(\a[28] ), .Y(new_n8624_));
  NAND4X1  g08431(.A(\a[48] ), .B(\a[47] ), .C(\a[29] ), .D(\a[28] ), .Y(new_n8625_));
  AOI22X1  g08432(.A0(new_n8625_), .A1(new_n8624_), .B0(new_n3893_), .B1(new_n2196_), .Y(new_n8626_));
  NAND4X1  g08433(.A(\a[47] ), .B(\a[46] ), .C(\a[30] ), .D(\a[29] ), .Y(new_n8627_));
  NAND3X1  g08434(.A(new_n8625_), .B(new_n8624_), .C(new_n8627_), .Y(new_n8628_));
  AOI22X1  g08435(.A0(\a[47] ), .A1(\a[29] ), .B0(\a[46] ), .B1(\a[30] ), .Y(new_n8629_));
  NAND2X1  g08436(.A(\a[48] ), .B(\a[28] ), .Y(new_n8630_));
  OAI22X1  g08437(.A0(new_n8630_), .A1(new_n8626_), .B0(new_n8629_), .B1(new_n8628_), .Y(new_n8631_));
  NAND4X1  g08438(.A(\a[42] ), .B(\a[40] ), .C(\a[36] ), .D(\a[34] ), .Y(new_n8632_));
  NAND4X1  g08439(.A(\a[42] ), .B(\a[41] ), .C(\a[35] ), .D(\a[34] ), .Y(new_n8633_));
  AOI22X1  g08440(.A0(new_n8633_), .A1(new_n8632_), .B0(new_n4404_), .B1(new_n2682_), .Y(new_n8634_));
  NAND2X1  g08441(.A(\a[42] ), .B(\a[34] ), .Y(new_n8635_));
  AOI21X1  g08442(.A0(new_n4404_), .A1(new_n2682_), .B0(new_n8634_), .Y(new_n8636_));
  INVX1    g08443(.A(new_n8636_), .Y(new_n8637_));
  AOI22X1  g08444(.A0(\a[41] ), .A1(\a[35] ), .B0(\a[40] ), .B1(\a[36] ), .Y(new_n8638_));
  OAI22X1  g08445(.A0(new_n8638_), .A1(new_n8637_), .B0(new_n8635_), .B1(new_n8634_), .Y(new_n8639_));
  XOR2X1   g08446(.A(new_n8639_), .B(new_n8631_), .Y(new_n8640_));
  AOI22X1  g08447(.A0(\a[52] ), .A1(\a[24] ), .B0(\a[51] ), .B1(\a[25] ), .Y(new_n8641_));
  AND2X1   g08448(.A(new_n7164_), .B(new_n1532_), .Y(new_n8642_));
  NOR3X1   g08449(.A(new_n8641_), .B(new_n8642_), .C(new_n3731_), .Y(new_n8643_));
  NOR2X1   g08450(.A(new_n8643_), .B(new_n8642_), .Y(new_n8644_));
  INVX1    g08451(.A(new_n8644_), .Y(new_n8645_));
  OAI22X1  g08452(.A0(new_n8645_), .A1(new_n8641_), .B0(new_n8643_), .B1(new_n3731_), .Y(new_n8646_));
  XOR2X1   g08453(.A(new_n8646_), .B(new_n8640_), .Y(new_n8647_));
  AND2X1   g08454(.A(new_n8379_), .B(new_n8377_), .Y(new_n8648_));
  OR2X1    g08455(.A(new_n8379_), .B(new_n8377_), .Y(new_n8649_));
  OAI21X1  g08456(.A0(new_n8383_), .A1(new_n8648_), .B0(new_n8649_), .Y(new_n8650_));
  XOR2X1   g08457(.A(new_n8650_), .B(new_n8647_), .Y(new_n8651_));
  NAND4X1  g08458(.A(\a[61] ), .B(\a[59] ), .C(\a[17] ), .D(\a[15] ), .Y(new_n8652_));
  NAND4X1  g08459(.A(\a[61] ), .B(\a[60] ), .C(\a[16] ), .D(\a[15] ), .Y(new_n8653_));
  AOI22X1  g08460(.A0(new_n8653_), .A1(new_n8652_), .B0(new_n6427_), .B1(new_n792_), .Y(new_n8654_));
  AND2X1   g08461(.A(\a[61] ), .B(\a[15] ), .Y(new_n8655_));
  INVX1    g08462(.A(new_n8655_), .Y(new_n8656_));
  AOI21X1  g08463(.A0(new_n6427_), .A1(new_n792_), .B0(new_n8654_), .Y(new_n8657_));
  INVX1    g08464(.A(new_n8657_), .Y(new_n8658_));
  AOI22X1  g08465(.A0(\a[60] ), .A1(\a[16] ), .B0(\a[59] ), .B1(\a[17] ), .Y(new_n8659_));
  OAI22X1  g08466(.A0(new_n8659_), .A1(new_n8658_), .B0(new_n8656_), .B1(new_n8654_), .Y(new_n8660_));
  XOR2X1   g08467(.A(new_n8660_), .B(new_n8504_), .Y(new_n8661_));
  AND2X1   g08468(.A(\a[58] ), .B(\a[18] ), .Y(new_n8662_));
  AOI22X1  g08469(.A0(\a[50] ), .A1(\a[26] ), .B0(\a[49] ), .B1(\a[27] ), .Y(new_n8663_));
  INVX1    g08470(.A(new_n8663_), .Y(new_n8664_));
  NAND4X1  g08471(.A(\a[50] ), .B(\a[49] ), .C(\a[27] ), .D(\a[26] ), .Y(new_n8665_));
  NAND3X1  g08472(.A(new_n8664_), .B(new_n8665_), .C(new_n8662_), .Y(new_n8666_));
  AOI22X1  g08473(.A0(new_n8664_), .A1(new_n8662_), .B0(new_n4321_), .B1(new_n1995_), .Y(new_n8667_));
  AOI22X1  g08474(.A0(new_n8667_), .A1(new_n8664_), .B0(new_n8666_), .B1(new_n8662_), .Y(new_n8668_));
  XOR2X1   g08475(.A(new_n8668_), .B(new_n8661_), .Y(new_n8669_));
  XOR2X1   g08476(.A(new_n8669_), .B(new_n8651_), .Y(new_n8670_));
  XOR2X1   g08477(.A(new_n8670_), .B(new_n8623_), .Y(new_n8671_));
  XOR2X1   g08478(.A(new_n8671_), .B(new_n8605_), .Y(new_n8672_));
  XOR2X1   g08479(.A(new_n8672_), .B(new_n8575_), .Y(new_n8673_));
  XOR2X1   g08480(.A(new_n8673_), .B(new_n8534_), .Y(new_n8674_));
  XOR2X1   g08481(.A(new_n8674_), .B(new_n8532_), .Y(\asquared[77] ));
  AND2X1   g08482(.A(new_n8573_), .B(new_n8537_), .Y(new_n8676_));
  AOI21X1  g08483(.A0(new_n8672_), .A1(new_n8574_), .B0(new_n8676_), .Y(new_n8677_));
  INVX1    g08484(.A(new_n8601_), .Y(new_n8678_));
  NOR2X1   g08485(.A(new_n8604_), .B(new_n8678_), .Y(new_n8679_));
  NOR2X1   g08486(.A(new_n8671_), .B(new_n8605_), .Y(new_n8680_));
  NOR2X1   g08487(.A(new_n8680_), .B(new_n8679_), .Y(new_n8681_));
  AND2X1   g08488(.A(new_n8621_), .B(new_n8608_), .Y(new_n8682_));
  AND2X1   g08489(.A(new_n8670_), .B(new_n8622_), .Y(new_n8683_));
  OR2X1    g08490(.A(new_n8683_), .B(new_n8682_), .Y(new_n8684_));
  AND2X1   g08491(.A(new_n8586_), .B(new_n8584_), .Y(new_n8685_));
  AOI21X1  g08492(.A0(new_n8600_), .A1(new_n8587_), .B0(new_n8685_), .Y(new_n8686_));
  AND2X1   g08493(.A(new_n8598_), .B(new_n8592_), .Y(new_n8687_));
  AOI21X1  g08494(.A0(new_n8599_), .A1(new_n8589_), .B0(new_n8687_), .Y(new_n8688_));
  AOI22X1  g08495(.A0(\a[55] ), .A1(\a[22] ), .B0(\a[51] ), .B1(\a[26] ), .Y(new_n8689_));
  AND2X1   g08496(.A(\a[43] ), .B(\a[34] ), .Y(new_n8690_));
  INVX1    g08497(.A(new_n8690_), .Y(new_n8691_));
  NOR4X1   g08498(.A(new_n4906_), .B(new_n4349_), .C(new_n1263_), .D(new_n1086_), .Y(new_n8692_));
  NOR3X1   g08499(.A(new_n8691_), .B(new_n8692_), .C(new_n8689_), .Y(new_n8693_));
  NOR2X1   g08500(.A(new_n8693_), .B(new_n8692_), .Y(new_n8694_));
  INVX1    g08501(.A(new_n8694_), .Y(new_n8695_));
  OAI22X1  g08502(.A0(new_n8695_), .A1(new_n8689_), .B0(new_n8693_), .B1(new_n8691_), .Y(new_n8696_));
  OAI22X1  g08503(.A0(new_n7338_), .A1(new_n2706_), .B0(new_n7336_), .B1(new_n1772_), .Y(new_n8697_));
  OAI21X1  g08504(.A0(new_n5239_), .A1(new_n1652_), .B0(new_n8697_), .Y(new_n8698_));
  AND2X1   g08505(.A(\a[52] ), .B(\a[25] ), .Y(new_n8699_));
  OAI22X1  g08506(.A0(new_n4835_), .A1(new_n1216_), .B0(new_n5245_), .B1(new_n1185_), .Y(new_n8700_));
  AOI21X1  g08507(.A0(new_n5238_), .A1(new_n1219_), .B0(new_n8697_), .Y(new_n8701_));
  AOI22X1  g08508(.A0(new_n8701_), .A1(new_n8700_), .B0(new_n8699_), .B1(new_n8698_), .Y(new_n8702_));
  XOR2X1   g08509(.A(new_n8702_), .B(new_n8696_), .Y(new_n8703_));
  AND2X1   g08510(.A(\a[61] ), .B(\a[16] ), .Y(new_n8704_));
  AOI22X1  g08511(.A0(\a[45] ), .A1(\a[32] ), .B0(\a[44] ), .B1(\a[33] ), .Y(new_n8705_));
  INVX1    g08512(.A(new_n8705_), .Y(new_n8706_));
  NAND4X1  g08513(.A(\a[45] ), .B(\a[44] ), .C(\a[33] ), .D(\a[32] ), .Y(new_n8707_));
  NAND3X1  g08514(.A(new_n8706_), .B(new_n8707_), .C(new_n8704_), .Y(new_n8708_));
  AOI22X1  g08515(.A0(new_n8706_), .A1(new_n8704_), .B0(new_n3918_), .B1(new_n2674_), .Y(new_n8709_));
  AOI22X1  g08516(.A0(new_n8709_), .A1(new_n8706_), .B0(new_n8708_), .B1(new_n8704_), .Y(new_n8710_));
  XOR2X1   g08517(.A(new_n8710_), .B(new_n8703_), .Y(new_n8711_));
  INVX1    g08518(.A(new_n8711_), .Y(new_n8712_));
  NAND2X1  g08519(.A(new_n8618_), .B(new_n8613_), .Y(new_n8713_));
  OAI21X1  g08520(.A0(new_n8620_), .A1(new_n8610_), .B0(new_n8713_), .Y(new_n8714_));
  AND2X1   g08521(.A(new_n8714_), .B(new_n8712_), .Y(new_n8715_));
  XOR2X1   g08522(.A(new_n8714_), .B(new_n8712_), .Y(new_n8716_));
  OAI21X1  g08523(.A0(new_n8714_), .A1(new_n8712_), .B0(new_n8688_), .Y(new_n8717_));
  OAI22X1  g08524(.A0(new_n8717_), .A1(new_n8715_), .B0(new_n8716_), .B1(new_n8688_), .Y(new_n8718_));
  XOR2X1   g08525(.A(new_n8718_), .B(new_n8686_), .Y(new_n8719_));
  XOR2X1   g08526(.A(new_n8719_), .B(new_n8684_), .Y(new_n8720_));
  XOR2X1   g08527(.A(new_n8720_), .B(new_n8681_), .Y(new_n8721_));
  NOR2X1   g08528(.A(new_n8571_), .B(new_n8542_), .Y(new_n8722_));
  AOI21X1  g08529(.A0(new_n8572_), .A1(new_n8540_), .B0(new_n8722_), .Y(new_n8723_));
  NAND2X1  g08530(.A(\a[59] ), .B(\a[18] ), .Y(new_n8724_));
  NAND2X1  g08531(.A(\a[60] ), .B(\a[17] ), .Y(new_n8725_));
  AOI22X1  g08532(.A0(new_n8725_), .A1(new_n8724_), .B0(new_n6427_), .B1(new_n796_), .Y(new_n8726_));
  XOR2X1   g08533(.A(new_n8726_), .B(new_n8644_), .Y(new_n8727_));
  INVX1    g08534(.A(new_n8497_), .Y(new_n8728_));
  AND2X1   g08535(.A(new_n8463_), .B(new_n8454_), .Y(new_n8729_));
  AOI21X1  g08536(.A0(new_n8609_), .A1(new_n8728_), .B0(new_n8729_), .Y(new_n8730_));
  XOR2X1   g08537(.A(new_n8730_), .B(new_n8727_), .Y(new_n8731_));
  NOR2X1   g08538(.A(new_n8490_), .B(new_n8472_), .Y(new_n8732_));
  AOI21X1  g08539(.A0(new_n8588_), .A1(new_n8429_), .B0(new_n8732_), .Y(new_n8733_));
  XOR2X1   g08540(.A(new_n8733_), .B(new_n8731_), .Y(new_n8734_));
  AND2X1   g08541(.A(new_n8650_), .B(new_n8647_), .Y(new_n8735_));
  AOI21X1  g08542(.A0(new_n8669_), .A1(new_n8651_), .B0(new_n8735_), .Y(new_n8736_));
  XOR2X1   g08543(.A(new_n8736_), .B(new_n8734_), .Y(new_n8737_));
  INVX1    g08544(.A(new_n8563_), .Y(new_n8738_));
  XOR2X1   g08545(.A(new_n8628_), .B(new_n8738_), .Y(new_n8739_));
  XOR2X1   g08546(.A(new_n8739_), .B(new_n8551_), .Y(new_n8740_));
  NOR3X1   g08547(.A(new_n8554_), .B(new_n3037_), .C(new_n1851_), .Y(new_n8741_));
  NOR2X1   g08548(.A(new_n8741_), .B(new_n8553_), .Y(new_n8742_));
  INVX1    g08549(.A(new_n8742_), .Y(new_n8743_));
  XOR2X1   g08550(.A(new_n8667_), .B(new_n8657_), .Y(new_n8744_));
  XOR2X1   g08551(.A(new_n8744_), .B(new_n8743_), .Y(new_n8745_));
  INVX1    g08552(.A(new_n8552_), .Y(new_n8746_));
  OR2X1    g08553(.A(new_n8565_), .B(new_n8558_), .Y(new_n8747_));
  OAI21X1  g08554(.A0(new_n8557_), .A1(new_n8746_), .B0(new_n8747_), .Y(new_n8748_));
  XOR2X1   g08555(.A(new_n8748_), .B(new_n8745_), .Y(new_n8749_));
  XOR2X1   g08556(.A(new_n8749_), .B(new_n8740_), .Y(new_n8750_));
  XOR2X1   g08557(.A(new_n8750_), .B(new_n8737_), .Y(new_n8751_));
  XOR2X1   g08558(.A(new_n8751_), .B(new_n8723_), .Y(new_n8752_));
  INVX1    g08559(.A(new_n8660_), .Y(new_n8753_));
  OR2X1    g08560(.A(new_n8668_), .B(new_n8661_), .Y(new_n8754_));
  OAI21X1  g08561(.A0(new_n8753_), .A1(new_n8504_), .B0(new_n8754_), .Y(new_n8755_));
  XOR2X1   g08562(.A(new_n8755_), .B(new_n8597_), .Y(new_n8756_));
  AND2X1   g08563(.A(new_n8639_), .B(new_n8631_), .Y(new_n8757_));
  AND2X1   g08564(.A(new_n8646_), .B(new_n8640_), .Y(new_n8758_));
  OR2X1    g08565(.A(new_n8758_), .B(new_n8757_), .Y(new_n8759_));
  XOR2X1   g08566(.A(new_n8759_), .B(new_n8756_), .Y(new_n8760_));
  NAND2X1  g08567(.A(new_n8569_), .B(new_n8566_), .Y(new_n8761_));
  NOR2X1   g08568(.A(new_n8569_), .B(new_n8566_), .Y(new_n8762_));
  OAI21X1  g08569(.A0(new_n8762_), .A1(new_n8544_), .B0(new_n8761_), .Y(new_n8763_));
  XOR2X1   g08570(.A(new_n8763_), .B(new_n8760_), .Y(new_n8764_));
  NAND2X1  g08571(.A(\a[47] ), .B(\a[30] ), .Y(new_n8765_));
  AND2X1   g08572(.A(\a[63] ), .B(\a[31] ), .Y(new_n8766_));
  NAND4X1  g08573(.A(\a[47] ), .B(\a[46] ), .C(\a[31] ), .D(\a[30] ), .Y(new_n8767_));
  NAND4X1  g08574(.A(\a[63] ), .B(\a[47] ), .C(\a[30] ), .D(\a[14] ), .Y(new_n8768_));
  AOI22X1  g08575(.A0(new_n8768_), .A1(new_n8767_), .B0(new_n8766_), .B1(new_n5734_), .Y(new_n8769_));
  NAND4X1  g08576(.A(\a[63] ), .B(\a[46] ), .C(\a[31] ), .D(\a[14] ), .Y(new_n8770_));
  NAND3X1  g08577(.A(new_n8768_), .B(new_n8767_), .C(new_n8770_), .Y(new_n8771_));
  AOI22X1  g08578(.A0(\a[63] ), .A1(\a[14] ), .B0(\a[46] ), .B1(\a[31] ), .Y(new_n8772_));
  OAI22X1  g08579(.A0(new_n8772_), .A1(new_n8771_), .B0(new_n8769_), .B1(new_n8765_), .Y(new_n8773_));
  NAND4X1  g08580(.A(\a[42] ), .B(\a[40] ), .C(\a[37] ), .D(\a[35] ), .Y(new_n8774_));
  NAND4X1  g08581(.A(\a[42] ), .B(\a[41] ), .C(\a[36] ), .D(\a[35] ), .Y(new_n8775_));
  AOI22X1  g08582(.A0(new_n8775_), .A1(new_n8774_), .B0(new_n4404_), .B1(new_n3330_), .Y(new_n8776_));
  NAND2X1  g08583(.A(\a[42] ), .B(\a[35] ), .Y(new_n8777_));
  NAND4X1  g08584(.A(\a[41] ), .B(\a[40] ), .C(\a[37] ), .D(\a[36] ), .Y(new_n8778_));
  NAND3X1  g08585(.A(new_n8775_), .B(new_n8774_), .C(new_n8778_), .Y(new_n8779_));
  AOI22X1  g08586(.A0(\a[41] ), .A1(\a[36] ), .B0(\a[40] ), .B1(\a[37] ), .Y(new_n8780_));
  OAI22X1  g08587(.A0(new_n8780_), .A1(new_n8779_), .B0(new_n8777_), .B1(new_n8776_), .Y(new_n8781_));
  XOR2X1   g08588(.A(new_n8781_), .B(new_n8773_), .Y(new_n8782_));
  NAND4X1  g08589(.A(\a[62] ), .B(\a[39] ), .C(\a[38] ), .D(\a[15] ), .Y(new_n8783_));
  AOI21X1  g08590(.A0(new_n4737_), .A1(\a[62] ), .B0(new_n3503_), .Y(new_n8784_));
  INVX1    g08591(.A(new_n8784_), .Y(new_n8785_));
  AOI21X1  g08592(.A0(\a[62] ), .A1(\a[15] ), .B0(\a[39] ), .Y(new_n8786_));
  OAI21X1  g08593(.A0(new_n8786_), .A1(new_n8785_), .B0(new_n8783_), .Y(new_n8787_));
  XOR2X1   g08594(.A(new_n8787_), .B(new_n8782_), .Y(new_n8788_));
  AND2X1   g08595(.A(new_n8409_), .B(new_n8229_), .Y(new_n8789_));
  OAI21X1  g08596(.A0(new_n8789_), .A1(new_n8578_), .B0(new_n8577_), .Y(new_n8790_));
  OAI21X1  g08597(.A0(new_n8583_), .A1(new_n8580_), .B0(new_n8790_), .Y(new_n8791_));
  XOR2X1   g08598(.A(new_n8791_), .B(new_n8788_), .Y(new_n8792_));
  NAND4X1  g08599(.A(\a[58] ), .B(\a[56] ), .C(\a[21] ), .D(\a[19] ), .Y(new_n8793_));
  NAND4X1  g08600(.A(\a[58] ), .B(\a[57] ), .C(\a[20] ), .D(\a[19] ), .Y(new_n8794_));
  AOI22X1  g08601(.A0(new_n8794_), .A1(new_n8793_), .B0(new_n5554_), .B1(new_n1236_), .Y(new_n8795_));
  NAND2X1  g08602(.A(\a[58] ), .B(\a[19] ), .Y(new_n8796_));
  NAND4X1  g08603(.A(\a[57] ), .B(\a[56] ), .C(\a[21] ), .D(\a[20] ), .Y(new_n8797_));
  NAND3X1  g08604(.A(new_n8794_), .B(new_n8793_), .C(new_n8797_), .Y(new_n8798_));
  AOI22X1  g08605(.A0(\a[57] ), .A1(\a[20] ), .B0(\a[56] ), .B1(\a[21] ), .Y(new_n8799_));
  OAI22X1  g08606(.A0(new_n8799_), .A1(new_n8798_), .B0(new_n8796_), .B1(new_n8795_), .Y(new_n8800_));
  XOR2X1   g08607(.A(new_n8800_), .B(new_n8636_), .Y(new_n8801_));
  INVX1    g08608(.A(new_n4035_), .Y(new_n8802_));
  OAI22X1  g08609(.A0(new_n7652_), .A1(new_n1672_), .B0(new_n8802_), .B1(new_n1673_), .Y(new_n8803_));
  OAI21X1  g08610(.A0(new_n4280_), .A1(new_n1675_), .B0(new_n8803_), .Y(new_n8804_));
  AND2X1   g08611(.A(\a[50] ), .B(\a[27] ), .Y(new_n8805_));
  AOI21X1  g08612(.A0(new_n4274_), .A1(new_n1674_), .B0(new_n8803_), .Y(new_n8806_));
  OAI22X1  g08613(.A0(new_n3915_), .A1(new_n1431_), .B0(new_n3926_), .B1(new_n1803_), .Y(new_n8807_));
  AOI22X1  g08614(.A0(new_n8807_), .A1(new_n8806_), .B0(new_n8805_), .B1(new_n8804_), .Y(new_n8808_));
  XOR2X1   g08615(.A(new_n8808_), .B(new_n8801_), .Y(new_n8809_));
  XOR2X1   g08616(.A(new_n8809_), .B(new_n8792_), .Y(new_n8810_));
  INVX1    g08617(.A(new_n8810_), .Y(new_n8811_));
  XOR2X1   g08618(.A(new_n8811_), .B(new_n8764_), .Y(new_n8812_));
  XOR2X1   g08619(.A(new_n8812_), .B(new_n8752_), .Y(new_n8813_));
  XOR2X1   g08620(.A(new_n8813_), .B(new_n8721_), .Y(new_n8814_));
  INVX1    g08621(.A(new_n8814_), .Y(new_n8815_));
  XOR2X1   g08622(.A(new_n8815_), .B(new_n8677_), .Y(new_n8816_));
  NOR2X1   g08623(.A(new_n8673_), .B(new_n8534_), .Y(new_n8817_));
  NAND2X1  g08624(.A(new_n8673_), .B(new_n8534_), .Y(new_n8818_));
  AOI21X1  g08625(.A0(new_n8818_), .A1(new_n8532_), .B0(new_n8817_), .Y(new_n8819_));
  XOR2X1   g08626(.A(new_n8819_), .B(new_n8816_), .Y(\asquared[78] ));
  OR2X1    g08627(.A(new_n8814_), .B(new_n8677_), .Y(new_n8821_));
  AND2X1   g08628(.A(new_n8814_), .B(new_n8677_), .Y(new_n8822_));
  OAI21X1  g08629(.A0(new_n8819_), .A1(new_n8822_), .B0(new_n8821_), .Y(new_n8823_));
  INVX1    g08630(.A(new_n8681_), .Y(new_n8824_));
  AND2X1   g08631(.A(new_n8720_), .B(new_n8824_), .Y(new_n8825_));
  OR2X1    g08632(.A(new_n8720_), .B(new_n8824_), .Y(new_n8826_));
  AOI21X1  g08633(.A0(new_n8813_), .A1(new_n8826_), .B0(new_n8825_), .Y(new_n8827_));
  AND2X1   g08634(.A(new_n8763_), .B(new_n8760_), .Y(new_n8828_));
  AOI21X1  g08635(.A0(new_n8810_), .A1(new_n8764_), .B0(new_n8828_), .Y(new_n8829_));
  NOR2X1   g08636(.A(new_n8736_), .B(new_n8734_), .Y(new_n8830_));
  AOI21X1  g08637(.A0(new_n8750_), .A1(new_n8737_), .B0(new_n8830_), .Y(new_n8831_));
  INVX1    g08638(.A(new_n8831_), .Y(new_n8832_));
  AND2X1   g08639(.A(new_n8755_), .B(new_n8597_), .Y(new_n8833_));
  AOI21X1  g08640(.A0(new_n8759_), .A1(new_n8756_), .B0(new_n8833_), .Y(new_n8834_));
  NAND4X1  g08641(.A(\a[60] ), .B(\a[57] ), .C(\a[21] ), .D(\a[18] ), .Y(new_n8835_));
  NAND4X1  g08642(.A(\a[60] ), .B(\a[59] ), .C(\a[19] ), .D(\a[18] ), .Y(new_n8836_));
  AOI22X1  g08643(.A0(new_n8836_), .A1(new_n8835_), .B0(new_n6120_), .B1(new_n1148_), .Y(new_n8837_));
  NAND4X1  g08644(.A(\a[59] ), .B(\a[57] ), .C(\a[21] ), .D(\a[19] ), .Y(new_n8838_));
  NAND3X1  g08645(.A(new_n8836_), .B(new_n8835_), .C(new_n8838_), .Y(new_n8839_));
  AOI22X1  g08646(.A0(\a[59] ), .A1(\a[19] ), .B0(\a[57] ), .B1(\a[21] ), .Y(new_n8840_));
  NAND2X1  g08647(.A(\a[60] ), .B(\a[18] ), .Y(new_n8841_));
  OAI22X1  g08648(.A0(new_n8841_), .A1(new_n8837_), .B0(new_n8840_), .B1(new_n8839_), .Y(new_n8842_));
  NAND4X1  g08649(.A(\a[51] ), .B(\a[49] ), .C(\a[29] ), .D(\a[27] ), .Y(new_n8843_));
  NAND4X1  g08650(.A(\a[51] ), .B(\a[50] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n8844_));
  AOI22X1  g08651(.A0(new_n8844_), .A1(new_n8843_), .B0(new_n4321_), .B1(new_n1674_), .Y(new_n8845_));
  NAND2X1  g08652(.A(\a[51] ), .B(\a[27] ), .Y(new_n8846_));
  NAND4X1  g08653(.A(\a[50] ), .B(\a[49] ), .C(\a[29] ), .D(\a[28] ), .Y(new_n8847_));
  NAND3X1  g08654(.A(new_n8844_), .B(new_n8843_), .C(new_n8847_), .Y(new_n8848_));
  AOI22X1  g08655(.A0(\a[50] ), .A1(\a[28] ), .B0(\a[49] ), .B1(\a[29] ), .Y(new_n8849_));
  OAI22X1  g08656(.A0(new_n8849_), .A1(new_n8848_), .B0(new_n8846_), .B1(new_n8845_), .Y(new_n8850_));
  XOR2X1   g08657(.A(new_n8850_), .B(new_n8842_), .Y(new_n8851_));
  AOI22X1  g08658(.A0(new_n6688_), .A1(new_n753_), .B0(new_n6789_), .B1(new_n689_), .Y(new_n8852_));
  AOI21X1  g08659(.A0(new_n6556_), .A1(new_n792_), .B0(new_n8852_), .Y(new_n8853_));
  AND2X1   g08660(.A(\a[63] ), .B(\a[15] ), .Y(new_n8854_));
  INVX1    g08661(.A(new_n8854_), .Y(new_n8855_));
  OAI22X1  g08662(.A0(new_n7973_), .A1(new_n2705_), .B0(new_n7972_), .B1(new_n1024_), .Y(new_n8856_));
  AOI21X1  g08663(.A0(new_n6556_), .A1(new_n792_), .B0(new_n8856_), .Y(new_n8857_));
  INVX1    g08664(.A(new_n8857_), .Y(new_n8858_));
  AOI22X1  g08665(.A0(\a[62] ), .A1(\a[16] ), .B0(\a[61] ), .B1(\a[17] ), .Y(new_n8859_));
  OAI22X1  g08666(.A0(new_n8859_), .A1(new_n8858_), .B0(new_n8855_), .B1(new_n8853_), .Y(new_n8860_));
  INVX1    g08667(.A(new_n8860_), .Y(new_n8861_));
  XOR2X1   g08668(.A(new_n8861_), .B(new_n8851_), .Y(new_n8862_));
  AOI22X1  g08669(.A0(\a[48] ), .A1(\a[30] ), .B0(\a[47] ), .B1(\a[31] ), .Y(new_n8863_));
  AND2X1   g08670(.A(\a[58] ), .B(\a[20] ), .Y(new_n8864_));
  INVX1    g08671(.A(new_n8864_), .Y(new_n8865_));
  AND2X1   g08672(.A(new_n4272_), .B(new_n2075_), .Y(new_n8866_));
  NOR3X1   g08673(.A(new_n8865_), .B(new_n8866_), .C(new_n8863_), .Y(new_n8867_));
  INVX1    g08674(.A(new_n8863_), .Y(new_n8868_));
  AOI21X1  g08675(.A0(new_n8864_), .A1(new_n8868_), .B0(new_n8866_), .Y(new_n8869_));
  INVX1    g08676(.A(new_n8869_), .Y(new_n8870_));
  OAI22X1  g08677(.A0(new_n8870_), .A1(new_n8863_), .B0(new_n8867_), .B1(new_n8865_), .Y(new_n8871_));
  OAI22X1  g08678(.A0(new_n3811_), .A1(new_n1851_), .B0(new_n5268_), .B1(new_n2028_), .Y(new_n8872_));
  INVX1    g08679(.A(new_n3809_), .Y(new_n8873_));
  INVX1    g08680(.A(new_n5270_), .Y(new_n8874_));
  OAI22X1  g08681(.A0(new_n8874_), .A1(new_n2920_), .B0(new_n8873_), .B1(new_n2675_), .Y(new_n8875_));
  OAI21X1  g08682(.A0(new_n7642_), .A1(new_n2919_), .B0(new_n8875_), .Y(new_n8876_));
  AOI21X1  g08683(.A0(new_n3918_), .A1(new_n2918_), .B0(new_n8875_), .Y(new_n8877_));
  AOI22X1  g08684(.A0(new_n8877_), .A1(new_n8872_), .B0(new_n8876_), .B1(new_n3808_), .Y(new_n8878_));
  XOR2X1   g08685(.A(new_n8878_), .B(new_n8871_), .Y(new_n8879_));
  NAND4X1  g08686(.A(\a[56] ), .B(\a[53] ), .C(\a[25] ), .D(\a[22] ), .Y(new_n8880_));
  NAND4X1  g08687(.A(\a[54] ), .B(\a[53] ), .C(\a[25] ), .D(\a[24] ), .Y(new_n8881_));
  AOI22X1  g08688(.A0(new_n8881_), .A1(new_n8880_), .B0(new_n5042_), .B1(new_n1530_), .Y(new_n8882_));
  NOR3X1   g08689(.A(new_n8882_), .B(new_n5245_), .C(new_n1326_), .Y(new_n8883_));
  OAI22X1  g08690(.A0(new_n6022_), .A1(new_n1086_), .B0(new_n4835_), .B1(new_n1185_), .Y(new_n8884_));
  AOI21X1  g08691(.A0(new_n5042_), .A1(new_n1530_), .B0(new_n8882_), .Y(new_n8885_));
  AOI21X1  g08692(.A0(new_n8885_), .A1(new_n8884_), .B0(new_n8883_), .Y(new_n8886_));
  XOR2X1   g08693(.A(new_n8886_), .B(new_n8879_), .Y(new_n8887_));
  XOR2X1   g08694(.A(new_n8887_), .B(new_n8862_), .Y(new_n8888_));
  XOR2X1   g08695(.A(new_n8888_), .B(new_n8834_), .Y(new_n8889_));
  XOR2X1   g08696(.A(new_n8889_), .B(new_n8832_), .Y(new_n8890_));
  INVX1    g08697(.A(new_n8890_), .Y(new_n8891_));
  XOR2X1   g08698(.A(new_n8891_), .B(new_n8829_), .Y(new_n8892_));
  INVX1    g08699(.A(new_n8892_), .Y(new_n8893_));
  INVX1    g08700(.A(new_n8723_), .Y(new_n8894_));
  NOR2X1   g08701(.A(new_n8812_), .B(new_n8752_), .Y(new_n8895_));
  AOI21X1  g08702(.A0(new_n8751_), .A1(new_n8894_), .B0(new_n8895_), .Y(new_n8896_));
  XOR2X1   g08703(.A(new_n8896_), .B(new_n8893_), .Y(new_n8897_));
  INVX1    g08704(.A(new_n8897_), .Y(new_n8898_));
  NOR2X1   g08705(.A(new_n8718_), .B(new_n8686_), .Y(new_n8899_));
  AOI21X1  g08706(.A0(new_n8719_), .A1(new_n8684_), .B0(new_n8899_), .Y(new_n8900_));
  NOR2X1   g08707(.A(new_n8808_), .B(new_n8801_), .Y(new_n8901_));
  AOI21X1  g08708(.A0(new_n8800_), .A1(new_n8637_), .B0(new_n8901_), .Y(new_n8902_));
  AND2X1   g08709(.A(new_n8781_), .B(new_n8773_), .Y(new_n8903_));
  AOI21X1  g08710(.A0(new_n8787_), .A1(new_n8782_), .B0(new_n8903_), .Y(new_n8904_));
  XOR2X1   g08711(.A(new_n8904_), .B(new_n8902_), .Y(new_n8905_));
  INVX1    g08712(.A(new_n8905_), .Y(new_n8906_));
  INVX1    g08713(.A(new_n8696_), .Y(new_n8907_));
  OR2X1    g08714(.A(new_n8702_), .B(new_n8907_), .Y(new_n8908_));
  OAI21X1  g08715(.A0(new_n8710_), .A1(new_n8703_), .B0(new_n8908_), .Y(new_n8909_));
  XOR2X1   g08716(.A(new_n8909_), .B(new_n8906_), .Y(new_n8910_));
  AND2X1   g08717(.A(new_n8748_), .B(new_n8745_), .Y(new_n8911_));
  AOI21X1  g08718(.A0(new_n8749_), .A1(new_n8740_), .B0(new_n8911_), .Y(new_n8912_));
  XOR2X1   g08719(.A(new_n8912_), .B(new_n8910_), .Y(new_n8913_));
  XOR2X1   g08720(.A(new_n8784_), .B(new_n8779_), .Y(new_n8914_));
  XOR2X1   g08721(.A(new_n8914_), .B(new_n8701_), .Y(new_n8915_));
  INVX1    g08722(.A(new_n8806_), .Y(new_n8916_));
  XOR2X1   g08723(.A(new_n8916_), .B(new_n8771_), .Y(new_n8917_));
  XOR2X1   g08724(.A(new_n8917_), .B(new_n8709_), .Y(new_n8918_));
  NOR2X1   g08725(.A(new_n8667_), .B(new_n8657_), .Y(new_n8919_));
  AOI21X1  g08726(.A0(new_n8744_), .A1(new_n8743_), .B0(new_n8919_), .Y(new_n8920_));
  XOR2X1   g08727(.A(new_n8920_), .B(new_n8918_), .Y(new_n8921_));
  XOR2X1   g08728(.A(new_n8921_), .B(new_n8915_), .Y(new_n8922_));
  XOR2X1   g08729(.A(new_n8922_), .B(new_n8913_), .Y(new_n8923_));
  XOR2X1   g08730(.A(new_n8923_), .B(new_n8900_), .Y(new_n8924_));
  NOR2X1   g08731(.A(new_n8716_), .B(new_n8688_), .Y(new_n8925_));
  AOI21X1  g08732(.A0(new_n8714_), .A1(new_n8711_), .B0(new_n8925_), .Y(new_n8926_));
  AND2X1   g08733(.A(new_n8791_), .B(new_n8788_), .Y(new_n8927_));
  AOI21X1  g08734(.A0(new_n8809_), .A1(new_n8792_), .B0(new_n8927_), .Y(new_n8928_));
  XOR2X1   g08735(.A(new_n8928_), .B(new_n8926_), .Y(new_n8929_));
  AOI22X1  g08736(.A0(\a[43] ), .A1(\a[35] ), .B0(\a[42] ), .B1(\a[36] ), .Y(new_n8930_));
  AND2X1   g08737(.A(\a[55] ), .B(\a[23] ), .Y(new_n8931_));
  INVX1    g08738(.A(new_n8931_), .Y(new_n8932_));
  AND2X1   g08739(.A(new_n3462_), .B(new_n2682_), .Y(new_n8933_));
  NOR3X1   g08740(.A(new_n8932_), .B(new_n8933_), .C(new_n8930_), .Y(new_n8934_));
  INVX1    g08741(.A(new_n8930_), .Y(new_n8935_));
  AOI21X1  g08742(.A0(new_n8931_), .A1(new_n8935_), .B0(new_n8933_), .Y(new_n8936_));
  INVX1    g08743(.A(new_n8936_), .Y(new_n8937_));
  OAI22X1  g08744(.A0(new_n8937_), .A1(new_n8930_), .B0(new_n8934_), .B1(new_n8932_), .Y(new_n8938_));
  AND2X1   g08745(.A(\a[52] ), .B(\a[26] ), .Y(new_n8939_));
  INVX1    g08746(.A(new_n8939_), .Y(new_n8940_));
  NAND4X1  g08747(.A(\a[52] ), .B(\a[41] ), .C(\a[37] ), .D(\a[26] ), .Y(new_n8941_));
  OAI21X1  g08748(.A0(new_n7618_), .A1(new_n7317_), .B0(new_n8941_), .Y(new_n8942_));
  OAI21X1  g08749(.A0(new_n8940_), .A1(new_n6179_), .B0(new_n8942_), .Y(new_n8943_));
  AOI21X1  g08750(.A0(new_n8939_), .A1(new_n2663_), .B0(new_n8942_), .Y(new_n8944_));
  OR2X1    g08751(.A(new_n8939_), .B(new_n2663_), .Y(new_n8945_));
  AOI22X1  g08752(.A0(new_n8945_), .A1(new_n8944_), .B0(new_n8943_), .B1(new_n4067_), .Y(new_n8946_));
  XOR2X1   g08753(.A(new_n8946_), .B(new_n8938_), .Y(new_n8947_));
  AND2X1   g08754(.A(new_n8628_), .B(new_n8738_), .Y(new_n8948_));
  AOI21X1  g08755(.A0(new_n8739_), .A1(new_n8551_), .B0(new_n8948_), .Y(new_n8949_));
  XOR2X1   g08756(.A(new_n8949_), .B(new_n8947_), .Y(new_n8950_));
  XOR2X1   g08757(.A(new_n8798_), .B(new_n8695_), .Y(new_n8951_));
  OAI21X1  g08758(.A0(new_n8643_), .A1(new_n8642_), .B0(new_n8726_), .Y(new_n8952_));
  OAI21X1  g08759(.A0(new_n6794_), .A1(new_n797_), .B0(new_n8952_), .Y(new_n8953_));
  XOR2X1   g08760(.A(new_n8953_), .B(new_n8951_), .Y(new_n8954_));
  AND2X1   g08761(.A(new_n8730_), .B(new_n8727_), .Y(new_n8955_));
  OR2X1    g08762(.A(new_n8730_), .B(new_n8727_), .Y(new_n8956_));
  OAI21X1  g08763(.A0(new_n8733_), .A1(new_n8955_), .B0(new_n8956_), .Y(new_n8957_));
  XOR2X1   g08764(.A(new_n8957_), .B(new_n8954_), .Y(new_n8958_));
  XOR2X1   g08765(.A(new_n8958_), .B(new_n8950_), .Y(new_n8959_));
  INVX1    g08766(.A(new_n8959_), .Y(new_n8960_));
  XOR2X1   g08767(.A(new_n8960_), .B(new_n8929_), .Y(new_n8961_));
  XOR2X1   g08768(.A(new_n8961_), .B(new_n8924_), .Y(new_n8962_));
  XOR2X1   g08769(.A(new_n8962_), .B(new_n8898_), .Y(new_n8963_));
  XOR2X1   g08770(.A(new_n8963_), .B(new_n8827_), .Y(new_n8964_));
  XOR2X1   g08771(.A(new_n8964_), .B(new_n8823_), .Y(\asquared[79] ));
  NOR2X1   g08772(.A(new_n8896_), .B(new_n8893_), .Y(new_n8966_));
  AOI21X1  g08773(.A0(new_n8962_), .A1(new_n8897_), .B0(new_n8966_), .Y(new_n8967_));
  NOR2X1   g08774(.A(new_n8912_), .B(new_n8910_), .Y(new_n8968_));
  AOI21X1  g08775(.A0(new_n8922_), .A1(new_n8913_), .B0(new_n8968_), .Y(new_n8969_));
  INVX1    g08776(.A(new_n8969_), .Y(new_n8970_));
  NAND2X1  g08777(.A(new_n8921_), .B(new_n8915_), .Y(new_n8971_));
  OAI21X1  g08778(.A0(new_n8920_), .A1(new_n8918_), .B0(new_n8971_), .Y(new_n8972_));
  NAND4X1  g08779(.A(\a[55] ), .B(\a[53] ), .C(\a[26] ), .D(\a[24] ), .Y(new_n8973_));
  NAND4X1  g08780(.A(\a[55] ), .B(\a[54] ), .C(\a[25] ), .D(\a[24] ), .Y(new_n8974_));
  AOI22X1  g08781(.A0(new_n8974_), .A1(new_n8973_), .B0(new_n5238_), .B1(new_n1770_), .Y(new_n8975_));
  NAND4X1  g08782(.A(\a[54] ), .B(\a[53] ), .C(\a[26] ), .D(\a[25] ), .Y(new_n8976_));
  NAND3X1  g08783(.A(new_n8974_), .B(new_n8973_), .C(new_n8976_), .Y(new_n8977_));
  AOI22X1  g08784(.A0(\a[54] ), .A1(\a[25] ), .B0(\a[53] ), .B1(\a[26] ), .Y(new_n8978_));
  NAND2X1  g08785(.A(\a[55] ), .B(\a[24] ), .Y(new_n8979_));
  OAI22X1  g08786(.A0(new_n8979_), .A1(new_n8975_), .B0(new_n8978_), .B1(new_n8977_), .Y(new_n8980_));
  NAND2X1  g08787(.A(\a[42] ), .B(\a[37] ), .Y(new_n8981_));
  NAND4X1  g08788(.A(\a[42] ), .B(\a[40] ), .C(\a[39] ), .D(\a[37] ), .Y(new_n8982_));
  NAND4X1  g08789(.A(\a[42] ), .B(\a[41] ), .C(\a[38] ), .D(\a[37] ), .Y(new_n8983_));
  AOI22X1  g08790(.A0(new_n8983_), .A1(new_n8982_), .B0(new_n4404_), .B1(new_n3503_), .Y(new_n8984_));
  AOI21X1  g08791(.A0(new_n4404_), .A1(new_n3503_), .B0(new_n8984_), .Y(new_n8985_));
  INVX1    g08792(.A(new_n8985_), .Y(new_n8986_));
  AOI22X1  g08793(.A0(\a[41] ), .A1(\a[38] ), .B0(\a[40] ), .B1(\a[39] ), .Y(new_n8987_));
  OAI22X1  g08794(.A0(new_n8987_), .A1(new_n8986_), .B0(new_n8984_), .B1(new_n8981_), .Y(new_n8988_));
  XOR2X1   g08795(.A(new_n8988_), .B(new_n8980_), .Y(new_n8989_));
  AND2X1   g08796(.A(\a[51] ), .B(\a[28] ), .Y(new_n8990_));
  INVX1    g08797(.A(new_n8990_), .Y(new_n8991_));
  AOI21X1  g08798(.A0(\a[62] ), .A1(\a[17] ), .B0(\a[40] ), .Y(new_n8992_));
  AND2X1   g08799(.A(\a[62] ), .B(\a[40] ), .Y(new_n8993_));
  AND2X1   g08800(.A(new_n8993_), .B(\a[17] ), .Y(new_n8994_));
  NOR3X1   g08801(.A(new_n8992_), .B(new_n8994_), .C(new_n8991_), .Y(new_n8995_));
  INVX1    g08802(.A(new_n8992_), .Y(new_n8996_));
  AOI21X1  g08803(.A0(new_n8996_), .A1(new_n8990_), .B0(new_n8994_), .Y(new_n8997_));
  INVX1    g08804(.A(new_n8997_), .Y(new_n8998_));
  OAI22X1  g08805(.A0(new_n8998_), .A1(new_n8992_), .B0(new_n8995_), .B1(new_n8991_), .Y(new_n8999_));
  INVX1    g08806(.A(new_n8999_), .Y(new_n9000_));
  XOR2X1   g08807(.A(new_n9000_), .B(new_n8989_), .Y(new_n9001_));
  OAI22X1  g08808(.A0(new_n6796_), .A1(new_n1149_), .B0(new_n6794_), .B1(new_n1521_), .Y(new_n9002_));
  OAI21X1  g08809(.A0(new_n6793_), .A1(new_n1794_), .B0(new_n9002_), .Y(new_n9003_));
  AOI21X1  g08810(.A0(new_n6121_), .A1(new_n1236_), .B0(new_n9002_), .Y(new_n9004_));
  OAI22X1  g08811(.A0(new_n5617_), .A1(new_n934_), .B0(new_n5379_), .B1(new_n1098_), .Y(new_n9005_));
  AND2X1   g08812(.A(\a[60] ), .B(\a[19] ), .Y(new_n9006_));
  AOI22X1  g08813(.A0(new_n9006_), .A1(new_n9003_), .B0(new_n9005_), .B1(new_n9004_), .Y(new_n9007_));
  AND2X1   g08814(.A(\a[57] ), .B(\a[22] ), .Y(new_n9008_));
  INVX1    g08815(.A(new_n9008_), .Y(new_n9009_));
  AOI22X1  g08816(.A0(\a[50] ), .A1(\a[29] ), .B0(\a[49] ), .B1(\a[30] ), .Y(new_n9010_));
  AND2X1   g08817(.A(new_n4321_), .B(new_n2196_), .Y(new_n9011_));
  NOR3X1   g08818(.A(new_n9010_), .B(new_n9011_), .C(new_n9009_), .Y(new_n9012_));
  INVX1    g08819(.A(new_n9010_), .Y(new_n9013_));
  AOI21X1  g08820(.A0(new_n9013_), .A1(new_n9008_), .B0(new_n9011_), .Y(new_n9014_));
  INVX1    g08821(.A(new_n9014_), .Y(new_n9015_));
  OAI22X1  g08822(.A0(new_n9015_), .A1(new_n9010_), .B0(new_n9012_), .B1(new_n9009_), .Y(new_n9016_));
  XOR2X1   g08823(.A(new_n9016_), .B(new_n9007_), .Y(new_n9017_));
  INVX1    g08824(.A(new_n9017_), .Y(new_n9018_));
  OAI22X1  g08825(.A0(new_n8299_), .A1(new_n2673_), .B0(new_n8297_), .B1(new_n2672_), .Y(new_n9019_));
  OAI21X1  g08826(.A0(new_n8296_), .A1(new_n2675_), .B0(new_n9019_), .Y(new_n9020_));
  AND2X1   g08827(.A(\a[48] ), .B(\a[31] ), .Y(new_n9021_));
  OAI22X1  g08828(.A0(new_n4041_), .A1(new_n2219_), .B0(new_n3460_), .B1(new_n1851_), .Y(new_n9022_));
  AOI21X1  g08829(.A0(new_n3893_), .A1(new_n2674_), .B0(new_n9019_), .Y(new_n9023_));
  AOI22X1  g08830(.A0(new_n9023_), .A1(new_n9022_), .B0(new_n9021_), .B1(new_n9020_), .Y(new_n9024_));
  XOR2X1   g08831(.A(new_n9024_), .B(new_n9018_), .Y(new_n9025_));
  XOR2X1   g08832(.A(new_n9025_), .B(new_n9001_), .Y(new_n9026_));
  XOR2X1   g08833(.A(new_n9026_), .B(new_n8972_), .Y(new_n9027_));
  XOR2X1   g08834(.A(new_n9027_), .B(new_n8970_), .Y(new_n9028_));
  INVX1    g08835(.A(new_n8709_), .Y(new_n9029_));
  AND2X1   g08836(.A(new_n8916_), .B(new_n8771_), .Y(new_n9030_));
  AOI21X1  g08837(.A0(new_n8917_), .A1(new_n9029_), .B0(new_n9030_), .Y(new_n9031_));
  NOR2X1   g08838(.A(new_n8914_), .B(new_n8701_), .Y(new_n9032_));
  AOI21X1  g08839(.A0(new_n8785_), .A1(new_n8779_), .B0(new_n9032_), .Y(new_n9033_));
  XOR2X1   g08840(.A(new_n9033_), .B(new_n9031_), .Y(new_n9034_));
  INVX1    g08841(.A(new_n9034_), .Y(new_n9035_));
  AND2X1   g08842(.A(new_n8850_), .B(new_n8842_), .Y(new_n9036_));
  AOI21X1  g08843(.A0(new_n8860_), .A1(new_n8851_), .B0(new_n9036_), .Y(new_n9037_));
  XOR2X1   g08844(.A(new_n9037_), .B(new_n9035_), .Y(new_n9038_));
  NOR2X1   g08845(.A(new_n8904_), .B(new_n8902_), .Y(new_n9039_));
  AOI21X1  g08846(.A0(new_n8909_), .A1(new_n8905_), .B0(new_n9039_), .Y(new_n9040_));
  XOR2X1   g08847(.A(new_n9040_), .B(new_n9038_), .Y(new_n9041_));
  AND2X1   g08848(.A(new_n8957_), .B(new_n8954_), .Y(new_n9042_));
  AOI21X1  g08849(.A0(new_n8958_), .A1(new_n8950_), .B0(new_n9042_), .Y(new_n9043_));
  XOR2X1   g08850(.A(new_n9043_), .B(new_n9041_), .Y(new_n9044_));
  XOR2X1   g08851(.A(new_n9044_), .B(new_n9028_), .Y(new_n9045_));
  INVX1    g08852(.A(new_n8923_), .Y(new_n9046_));
  OR2X1    g08853(.A(new_n9046_), .B(new_n8900_), .Y(new_n9047_));
  OAI21X1  g08854(.A0(new_n8961_), .A1(new_n8924_), .B0(new_n9047_), .Y(new_n9048_));
  INVX1    g08855(.A(new_n9048_), .Y(new_n9049_));
  OR2X1    g08856(.A(new_n9049_), .B(new_n9045_), .Y(new_n9050_));
  NAND2X1  g08857(.A(new_n8959_), .B(new_n8929_), .Y(new_n9051_));
  OAI21X1  g08858(.A0(new_n8928_), .A1(new_n8926_), .B0(new_n9051_), .Y(new_n9052_));
  XOR2X1   g08859(.A(new_n8860_), .B(new_n8851_), .Y(new_n9053_));
  NAND2X1  g08860(.A(new_n8887_), .B(new_n9053_), .Y(new_n9054_));
  OAI21X1  g08861(.A0(new_n8888_), .A1(new_n8834_), .B0(new_n9054_), .Y(new_n9055_));
  INVX1    g08862(.A(new_n8885_), .Y(new_n9056_));
  XOR2X1   g08863(.A(new_n8848_), .B(new_n8839_), .Y(new_n9057_));
  XOR2X1   g08864(.A(new_n9057_), .B(new_n9056_), .Y(new_n9058_));
  INVX1    g08865(.A(new_n9058_), .Y(new_n9059_));
  INVX1    g08866(.A(new_n8938_), .Y(new_n9060_));
  OR2X1    g08867(.A(new_n8946_), .B(new_n9060_), .Y(new_n9061_));
  OAI21X1  g08868(.A0(new_n8949_), .A1(new_n8947_), .B0(new_n9061_), .Y(new_n9062_));
  XOR2X1   g08869(.A(new_n9062_), .B(new_n9059_), .Y(new_n9063_));
  AOI22X1  g08870(.A0(\a[45] ), .A1(\a[34] ), .B0(\a[44] ), .B1(\a[35] ), .Y(new_n9064_));
  AND2X1   g08871(.A(\a[63] ), .B(\a[16] ), .Y(new_n9065_));
  INVX1    g08872(.A(new_n9065_), .Y(new_n9066_));
  AND2X1   g08873(.A(new_n3918_), .B(new_n2361_), .Y(new_n9067_));
  NOR3X1   g08874(.A(new_n9066_), .B(new_n9067_), .C(new_n9064_), .Y(new_n9068_));
  NOR2X1   g08875(.A(new_n9068_), .B(new_n9067_), .Y(new_n9069_));
  INVX1    g08876(.A(new_n9069_), .Y(new_n9070_));
  OAI22X1  g08877(.A0(new_n9070_), .A1(new_n9064_), .B0(new_n9068_), .B1(new_n9066_), .Y(new_n9071_));
  AND2X1   g08878(.A(\a[43] ), .B(\a[36] ), .Y(new_n9072_));
  AND2X1   g08879(.A(\a[56] ), .B(\a[27] ), .Y(new_n9073_));
  AND2X1   g08880(.A(new_n9073_), .B(new_n8431_), .Y(new_n9074_));
  AOI22X1  g08881(.A0(\a[56] ), .A1(\a[23] ), .B0(\a[52] ), .B1(\a[27] ), .Y(new_n9075_));
  OR4X1    g08882(.A(new_n9075_), .B(new_n9074_), .C(new_n3037_), .D(new_n2583_), .Y(new_n9076_));
  NOR3X1   g08883(.A(new_n9075_), .B(new_n9074_), .C(new_n9072_), .Y(new_n9077_));
  AOI21X1  g08884(.A0(new_n9076_), .A1(new_n9072_), .B0(new_n9077_), .Y(new_n9078_));
  XOR2X1   g08885(.A(new_n9078_), .B(new_n9071_), .Y(new_n9079_));
  AND2X1   g08886(.A(new_n8798_), .B(new_n8695_), .Y(new_n9080_));
  AOI21X1  g08887(.A0(new_n8953_), .A1(new_n8951_), .B0(new_n9080_), .Y(new_n9081_));
  XOR2X1   g08888(.A(new_n9081_), .B(new_n9079_), .Y(new_n9082_));
  INVX1    g08889(.A(new_n9082_), .Y(new_n9083_));
  XOR2X1   g08890(.A(new_n9083_), .B(new_n9063_), .Y(new_n9084_));
  XOR2X1   g08891(.A(new_n9084_), .B(new_n9055_), .Y(new_n9085_));
  INVX1    g08892(.A(new_n8871_), .Y(new_n9086_));
  OR2X1    g08893(.A(new_n8878_), .B(new_n9086_), .Y(new_n9087_));
  OAI21X1  g08894(.A0(new_n8886_), .A1(new_n8879_), .B0(new_n9087_), .Y(new_n9088_));
  AND2X1   g08895(.A(\a[61] ), .B(\a[18] ), .Y(new_n9089_));
  XOR2X1   g08896(.A(new_n9089_), .B(new_n8944_), .Y(new_n9090_));
  XOR2X1   g08897(.A(new_n9090_), .B(new_n8937_), .Y(new_n9091_));
  XOR2X1   g08898(.A(new_n8869_), .B(new_n8857_), .Y(new_n9092_));
  XOR2X1   g08899(.A(new_n9092_), .B(new_n8877_), .Y(new_n9093_));
  XOR2X1   g08900(.A(new_n9093_), .B(new_n9091_), .Y(new_n9094_));
  XOR2X1   g08901(.A(new_n9094_), .B(new_n9088_), .Y(new_n9095_));
  XOR2X1   g08902(.A(new_n9095_), .B(new_n9085_), .Y(new_n9096_));
  XOR2X1   g08903(.A(new_n9096_), .B(new_n9052_), .Y(new_n9097_));
  NAND2X1  g08904(.A(new_n8889_), .B(new_n8832_), .Y(new_n9098_));
  OAI21X1  g08905(.A0(new_n8891_), .A1(new_n8829_), .B0(new_n9098_), .Y(new_n9099_));
  XOR2X1   g08906(.A(new_n9099_), .B(new_n9097_), .Y(new_n9100_));
  XOR2X1   g08907(.A(new_n9048_), .B(new_n9045_), .Y(new_n9101_));
  AND2X1   g08908(.A(new_n9101_), .B(new_n9100_), .Y(new_n9102_));
  AOI21X1  g08909(.A0(new_n9049_), .A1(new_n9045_), .B0(new_n9100_), .Y(new_n9103_));
  AOI21X1  g08910(.A0(new_n9103_), .A1(new_n9050_), .B0(new_n9102_), .Y(new_n9104_));
  XOR2X1   g08911(.A(new_n9104_), .B(new_n8967_), .Y(new_n9105_));
  NOR2X1   g08912(.A(new_n8963_), .B(new_n8827_), .Y(new_n9106_));
  NAND2X1  g08913(.A(new_n8963_), .B(new_n8827_), .Y(new_n9107_));
  AOI21X1  g08914(.A0(new_n9107_), .A1(new_n8823_), .B0(new_n9106_), .Y(new_n9108_));
  XOR2X1   g08915(.A(new_n9108_), .B(new_n9105_), .Y(\asquared[80] ));
  AOI21X1  g08916(.A0(new_n9048_), .A1(new_n9045_), .B0(new_n9102_), .Y(new_n9110_));
  AND2X1   g08917(.A(new_n9096_), .B(new_n9052_), .Y(new_n9111_));
  AOI21X1  g08918(.A0(new_n9099_), .A1(new_n9097_), .B0(new_n9111_), .Y(new_n9112_));
  INVX1    g08919(.A(new_n9112_), .Y(new_n9113_));
  AND2X1   g08920(.A(new_n9084_), .B(new_n9055_), .Y(new_n9114_));
  AND2X1   g08921(.A(new_n9095_), .B(new_n9085_), .Y(new_n9115_));
  OR2X1    g08922(.A(new_n9115_), .B(new_n9114_), .Y(new_n9116_));
  AND2X1   g08923(.A(new_n8909_), .B(new_n8905_), .Y(new_n9117_));
  OAI21X1  g08924(.A0(new_n9117_), .A1(new_n9039_), .B0(new_n9038_), .Y(new_n9118_));
  OAI21X1  g08925(.A0(new_n9043_), .A1(new_n9041_), .B0(new_n9118_), .Y(new_n9119_));
  AOI22X1  g08926(.A0(\a[63] ), .A1(\a[17] ), .B0(\a[51] ), .B1(\a[29] ), .Y(new_n9120_));
  AND2X1   g08927(.A(\a[47] ), .B(\a[33] ), .Y(new_n9121_));
  INVX1    g08928(.A(new_n9121_), .Y(new_n9122_));
  NOR4X1   g08929(.A(new_n6549_), .B(new_n4349_), .C(new_n1803_), .D(new_n616_), .Y(new_n9123_));
  NOR3X1   g08930(.A(new_n9122_), .B(new_n9123_), .C(new_n9120_), .Y(new_n9124_));
  INVX1    g08931(.A(new_n9120_), .Y(new_n9125_));
  AOI21X1  g08932(.A0(new_n9121_), .A1(new_n9125_), .B0(new_n9123_), .Y(new_n9126_));
  INVX1    g08933(.A(new_n9126_), .Y(new_n9127_));
  OAI22X1  g08934(.A0(new_n9127_), .A1(new_n9120_), .B0(new_n9124_), .B1(new_n9122_), .Y(new_n9128_));
  OAI22X1  g08935(.A0(new_n8874_), .A1(new_n5418_), .B0(new_n8873_), .B1(new_n4915_), .Y(new_n9129_));
  OAI21X1  g08936(.A0(new_n7642_), .A1(new_n5417_), .B0(new_n9129_), .Y(new_n9130_));
  AND2X1   g08937(.A(\a[46] ), .B(\a[34] ), .Y(new_n9131_));
  AOI21X1  g08938(.A0(new_n3918_), .A1(new_n2682_), .B0(new_n9129_), .Y(new_n9132_));
  OAI21X1  g08939(.A0(new_n5268_), .A1(new_n2583_), .B0(new_n4009_), .Y(new_n9133_));
  AOI22X1  g08940(.A0(new_n9133_), .A1(new_n9132_), .B0(new_n9131_), .B1(new_n9130_), .Y(new_n9134_));
  XOR2X1   g08941(.A(new_n9134_), .B(new_n9128_), .Y(new_n9135_));
  AND2X1   g08942(.A(\a[61] ), .B(\a[19] ), .Y(new_n9136_));
  AND2X1   g08943(.A(\a[62] ), .B(\a[18] ), .Y(new_n9137_));
  OAI22X1  g08944(.A0(new_n9137_), .A1(new_n9136_), .B0(new_n6557_), .B1(new_n1518_), .Y(new_n9138_));
  XOR2X1   g08945(.A(new_n9138_), .B(new_n8998_), .Y(new_n9139_));
  INVX1    g08946(.A(new_n9139_), .Y(new_n9140_));
  XOR2X1   g08947(.A(new_n9140_), .B(new_n9135_), .Y(new_n9141_));
  AND2X1   g08948(.A(new_n6121_), .B(new_n1154_), .Y(new_n9142_));
  AOI22X1  g08949(.A0(new_n6795_), .A1(new_n2134_), .B0(new_n6427_), .B1(new_n1236_), .Y(new_n9143_));
  AOI22X1  g08950(.A0(\a[59] ), .A1(\a[21] ), .B0(\a[58] ), .B1(\a[22] ), .Y(new_n9144_));
  AOI21X1  g08951(.A0(new_n6121_), .A1(new_n1154_), .B0(new_n9144_), .Y(new_n9145_));
  AND2X1   g08952(.A(\a[60] ), .B(\a[20] ), .Y(new_n9146_));
  OAI22X1  g08953(.A0(new_n9146_), .A1(new_n9145_), .B0(new_n9143_), .B1(new_n9142_), .Y(new_n9147_));
  XOR2X1   g08954(.A(new_n9147_), .B(new_n8985_), .Y(new_n9148_));
  OAI22X1  g08955(.A0(new_n7652_), .A1(new_n2076_), .B0(new_n8802_), .B1(new_n4923_), .Y(new_n9149_));
  OAI21X1  g08956(.A0(new_n4280_), .A1(new_n2672_), .B0(new_n9149_), .Y(new_n9150_));
  AND2X1   g08957(.A(\a[50] ), .B(\a[30] ), .Y(new_n9151_));
  AOI21X1  g08958(.A0(new_n4274_), .A1(new_n2671_), .B0(new_n9149_), .Y(new_n9152_));
  OAI22X1  g08959(.A0(new_n3915_), .A1(new_n1704_), .B0(new_n3926_), .B1(new_n2219_), .Y(new_n9153_));
  AOI22X1  g08960(.A0(new_n9153_), .A1(new_n9152_), .B0(new_n9151_), .B1(new_n9150_), .Y(new_n9154_));
  XOR2X1   g08961(.A(new_n9154_), .B(new_n9148_), .Y(new_n9155_));
  OAI22X1  g08962(.A0(new_n6022_), .A1(new_n1185_), .B0(new_n4835_), .B1(new_n1263_), .Y(new_n9156_));
  NAND4X1  g08963(.A(\a[57] ), .B(\a[54] ), .C(\a[26] ), .D(\a[23] ), .Y(new_n9157_));
  NAND4X1  g08964(.A(\a[57] ), .B(\a[56] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n9158_));
  AOI22X1  g08965(.A0(new_n9158_), .A1(new_n9157_), .B0(new_n5042_), .B1(new_n1650_), .Y(new_n9159_));
  AOI21X1  g08966(.A0(new_n5042_), .A1(new_n1650_), .B0(new_n9159_), .Y(new_n9160_));
  NOR3X1   g08967(.A(new_n9159_), .B(new_n5441_), .C(new_n1216_), .Y(new_n9161_));
  AOI21X1  g08968(.A0(new_n9160_), .A1(new_n9156_), .B0(new_n9161_), .Y(new_n9162_));
  AND2X1   g08969(.A(\a[55] ), .B(\a[25] ), .Y(new_n9163_));
  INVX1    g08970(.A(new_n9163_), .Y(new_n9164_));
  AOI22X1  g08971(.A0(\a[43] ), .A1(\a[37] ), .B0(\a[42] ), .B1(\a[38] ), .Y(new_n9165_));
  AND2X1   g08972(.A(new_n3462_), .B(new_n3164_), .Y(new_n9166_));
  NOR3X1   g08973(.A(new_n9165_), .B(new_n9166_), .C(new_n9164_), .Y(new_n9167_));
  INVX1    g08974(.A(new_n9165_), .Y(new_n9168_));
  AOI21X1  g08975(.A0(new_n9168_), .A1(new_n9163_), .B0(new_n9166_), .Y(new_n9169_));
  INVX1    g08976(.A(new_n9169_), .Y(new_n9170_));
  OAI22X1  g08977(.A0(new_n9170_), .A1(new_n9165_), .B0(new_n9167_), .B1(new_n9164_), .Y(new_n9171_));
  XOR2X1   g08978(.A(new_n9171_), .B(new_n9162_), .Y(new_n9172_));
  AOI22X1  g08979(.A0(\a[53] ), .A1(\a[27] ), .B0(\a[52] ), .B1(\a[28] ), .Y(new_n9173_));
  INVX1    g08980(.A(new_n9173_), .Y(new_n9174_));
  NAND4X1  g08981(.A(\a[53] ), .B(\a[52] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n9175_));
  AOI21X1  g08982(.A0(new_n9174_), .A1(new_n9175_), .B0(new_n7617_), .Y(new_n9176_));
  AOI22X1  g08983(.A0(new_n9174_), .A1(new_n2847_), .B0(new_n5048_), .B1(new_n1671_), .Y(new_n9177_));
  AOI21X1  g08984(.A0(new_n9177_), .A1(new_n9174_), .B0(new_n9176_), .Y(new_n9178_));
  XOR2X1   g08985(.A(new_n9178_), .B(new_n9172_), .Y(new_n9179_));
  XOR2X1   g08986(.A(new_n9179_), .B(new_n9155_), .Y(new_n9180_));
  XOR2X1   g08987(.A(new_n9180_), .B(new_n9141_), .Y(new_n9181_));
  XOR2X1   g08988(.A(new_n9181_), .B(new_n9119_), .Y(new_n9182_));
  XOR2X1   g08989(.A(new_n9182_), .B(new_n9116_), .Y(new_n9183_));
  XOR2X1   g08990(.A(new_n9183_), .B(new_n9113_), .Y(new_n9184_));
  INVX1    g08991(.A(new_n9184_), .Y(new_n9185_));
  AND2X1   g08992(.A(new_n9027_), .B(new_n8970_), .Y(new_n9186_));
  AOI21X1  g08993(.A0(new_n9044_), .A1(new_n9028_), .B0(new_n9186_), .Y(new_n9187_));
  NOR2X1   g08994(.A(new_n9025_), .B(new_n9001_), .Y(new_n9188_));
  AOI21X1  g08995(.A0(new_n9026_), .A1(new_n8972_), .B0(new_n9188_), .Y(new_n9189_));
  NOR3X1   g08996(.A(new_n9075_), .B(new_n3037_), .C(new_n2583_), .Y(new_n9190_));
  NOR2X1   g08997(.A(new_n9190_), .B(new_n9074_), .Y(new_n9191_));
  INVX1    g08998(.A(new_n9191_), .Y(new_n9192_));
  XOR2X1   g08999(.A(new_n8977_), .B(new_n9070_), .Y(new_n9193_));
  XOR2X1   g09000(.A(new_n9193_), .B(new_n9192_), .Y(new_n9194_));
  AND2X1   g09001(.A(new_n9076_), .B(new_n9072_), .Y(new_n9195_));
  OAI21X1  g09002(.A0(new_n9077_), .A1(new_n9195_), .B0(new_n9071_), .Y(new_n9196_));
  OAI21X1  g09003(.A0(new_n9081_), .A1(new_n9079_), .B0(new_n9196_), .Y(new_n9197_));
  XOR2X1   g09004(.A(new_n9197_), .B(new_n9194_), .Y(new_n9198_));
  NOR2X1   g09005(.A(new_n9033_), .B(new_n9031_), .Y(new_n9199_));
  NOR2X1   g09006(.A(new_n9037_), .B(new_n9035_), .Y(new_n9200_));
  NOR2X1   g09007(.A(new_n9200_), .B(new_n9199_), .Y(new_n9201_));
  XOR2X1   g09008(.A(new_n9201_), .B(new_n9198_), .Y(new_n9202_));
  XOR2X1   g09009(.A(new_n9202_), .B(new_n9189_), .Y(new_n9203_));
  INVX1    g09010(.A(new_n9203_), .Y(new_n9204_));
  INVX1    g09011(.A(new_n9023_), .Y(new_n9205_));
  XOR2X1   g09012(.A(new_n9014_), .B(new_n9004_), .Y(new_n9206_));
  XOR2X1   g09013(.A(new_n9206_), .B(new_n9205_), .Y(new_n9207_));
  INVX1    g09014(.A(new_n9207_), .Y(new_n9208_));
  AND2X1   g09015(.A(new_n8988_), .B(new_n8980_), .Y(new_n9209_));
  AND2X1   g09016(.A(new_n8999_), .B(new_n8989_), .Y(new_n9210_));
  OR2X1    g09017(.A(new_n9210_), .B(new_n9209_), .Y(new_n9211_));
  INVX1    g09018(.A(new_n9016_), .Y(new_n9212_));
  OR2X1    g09019(.A(new_n9212_), .B(new_n9007_), .Y(new_n9213_));
  OAI21X1  g09020(.A0(new_n9024_), .A1(new_n9017_), .B0(new_n9213_), .Y(new_n9214_));
  XOR2X1   g09021(.A(new_n9214_), .B(new_n9211_), .Y(new_n9215_));
  XOR2X1   g09022(.A(new_n9215_), .B(new_n9208_), .Y(new_n9216_));
  XOR2X1   g09023(.A(new_n9216_), .B(new_n9204_), .Y(new_n9217_));
  INVX1    g09024(.A(new_n9217_), .Y(new_n9218_));
  AND2X1   g09025(.A(new_n8848_), .B(new_n8839_), .Y(new_n9219_));
  AOI21X1  g09026(.A0(new_n9057_), .A1(new_n9056_), .B0(new_n9219_), .Y(new_n9220_));
  INVX1    g09027(.A(new_n8877_), .Y(new_n9221_));
  NOR2X1   g09028(.A(new_n8869_), .B(new_n8857_), .Y(new_n9222_));
  AOI21X1  g09029(.A0(new_n9092_), .A1(new_n9221_), .B0(new_n9222_), .Y(new_n9223_));
  XOR2X1   g09030(.A(new_n9223_), .B(new_n9220_), .Y(new_n9224_));
  INVX1    g09031(.A(new_n8944_), .Y(new_n9225_));
  NAND2X1  g09032(.A(new_n9089_), .B(new_n9225_), .Y(new_n9226_));
  OAI21X1  g09033(.A0(new_n9090_), .A1(new_n8936_), .B0(new_n9226_), .Y(new_n9227_));
  XOR2X1   g09034(.A(new_n9227_), .B(new_n9224_), .Y(new_n9228_));
  NOR2X1   g09035(.A(new_n9083_), .B(new_n9063_), .Y(new_n9229_));
  AOI21X1  g09036(.A0(new_n9062_), .A1(new_n9058_), .B0(new_n9229_), .Y(new_n9230_));
  NOR2X1   g09037(.A(new_n9093_), .B(new_n9091_), .Y(new_n9231_));
  AOI21X1  g09038(.A0(new_n9094_), .A1(new_n9088_), .B0(new_n9231_), .Y(new_n9232_));
  XOR2X1   g09039(.A(new_n9232_), .B(new_n9230_), .Y(new_n9233_));
  XOR2X1   g09040(.A(new_n9233_), .B(new_n9228_), .Y(new_n9234_));
  XOR2X1   g09041(.A(new_n9234_), .B(new_n9218_), .Y(new_n9235_));
  XOR2X1   g09042(.A(new_n9235_), .B(new_n9187_), .Y(new_n9236_));
  XOR2X1   g09043(.A(new_n9236_), .B(new_n9185_), .Y(new_n9237_));
  NOR2X1   g09044(.A(new_n9237_), .B(new_n9110_), .Y(new_n9238_));
  INVX1    g09045(.A(new_n9238_), .Y(new_n9239_));
  INVX1    g09046(.A(new_n8967_), .Y(new_n9240_));
  NAND2X1  g09047(.A(new_n9104_), .B(new_n9240_), .Y(new_n9241_));
  NOR2X1   g09048(.A(new_n9104_), .B(new_n9240_), .Y(new_n9242_));
  OAI21X1  g09049(.A0(new_n9108_), .A1(new_n9242_), .B0(new_n9241_), .Y(new_n9243_));
  AND2X1   g09050(.A(new_n9237_), .B(new_n9110_), .Y(new_n9244_));
  INVX1    g09051(.A(new_n9244_), .Y(new_n9245_));
  AOI21X1  g09052(.A0(new_n9239_), .A1(new_n9245_), .B0(new_n9243_), .Y(new_n9246_));
  AND2X1   g09053(.A(new_n9245_), .B(new_n9243_), .Y(new_n9247_));
  AOI21X1  g09054(.A0(new_n9247_), .A1(new_n9239_), .B0(new_n9246_), .Y(\asquared[81] ));
  AOI21X1  g09055(.A0(new_n9245_), .A1(new_n9243_), .B0(new_n9238_), .Y(new_n9249_));
  NAND2X1  g09056(.A(new_n9234_), .B(new_n9217_), .Y(new_n9250_));
  OAI21X1  g09057(.A0(new_n9235_), .A1(new_n9187_), .B0(new_n9250_), .Y(new_n9251_));
  OR2X1    g09058(.A(new_n9202_), .B(new_n9189_), .Y(new_n9252_));
  OAI21X1  g09059(.A0(new_n9216_), .A1(new_n9204_), .B0(new_n9252_), .Y(new_n9253_));
  NOR2X1   g09060(.A(new_n9232_), .B(new_n9230_), .Y(new_n9254_));
  AOI21X1  g09061(.A0(new_n9233_), .A1(new_n9228_), .B0(new_n9254_), .Y(new_n9255_));
  AND2X1   g09062(.A(\a[62] ), .B(\a[41] ), .Y(new_n9256_));
  AOI21X1  g09063(.A0(new_n9256_), .A1(\a[19] ), .B0(new_n4404_), .Y(new_n9257_));
  INVX1    g09064(.A(new_n9257_), .Y(new_n9258_));
  AOI21X1  g09065(.A0(\a[62] ), .A1(\a[19] ), .B0(\a[41] ), .Y(new_n9259_));
  NAND4X1  g09066(.A(\a[62] ), .B(\a[41] ), .C(\a[40] ), .D(\a[19] ), .Y(new_n9260_));
  OAI21X1  g09067(.A0(new_n9259_), .A1(new_n9258_), .B0(new_n9260_), .Y(new_n9261_));
  NAND4X1  g09068(.A(\a[59] ), .B(\a[56] ), .C(\a[25] ), .D(\a[22] ), .Y(new_n9262_));
  NAND4X1  g09069(.A(\a[59] ), .B(\a[58] ), .C(\a[23] ), .D(\a[22] ), .Y(new_n9263_));
  AOI22X1  g09070(.A0(new_n9263_), .A1(new_n9262_), .B0(new_n5381_), .B1(new_n1134_), .Y(new_n9264_));
  NAND2X1  g09071(.A(\a[59] ), .B(\a[22] ), .Y(new_n9265_));
  NAND4X1  g09072(.A(\a[58] ), .B(\a[56] ), .C(\a[25] ), .D(\a[23] ), .Y(new_n9266_));
  NAND3X1  g09073(.A(new_n9263_), .B(new_n9262_), .C(new_n9266_), .Y(new_n9267_));
  AOI22X1  g09074(.A0(\a[58] ), .A1(\a[23] ), .B0(\a[56] ), .B1(\a[25] ), .Y(new_n9268_));
  OAI22X1  g09075(.A0(new_n9268_), .A1(new_n9267_), .B0(new_n9265_), .B1(new_n9264_), .Y(new_n9269_));
  XOR2X1   g09076(.A(new_n9269_), .B(new_n9261_), .Y(new_n9270_));
  AOI22X1  g09077(.A0(\a[48] ), .A1(\a[33] ), .B0(\a[47] ), .B1(\a[34] ), .Y(new_n9271_));
  INVX1    g09078(.A(new_n9271_), .Y(new_n9272_));
  NAND4X1  g09079(.A(\a[48] ), .B(\a[47] ), .C(\a[34] ), .D(\a[33] ), .Y(new_n9273_));
  NAND3X1  g09080(.A(new_n9272_), .B(new_n9273_), .C(new_n6937_), .Y(new_n9274_));
  AOI22X1  g09081(.A0(new_n9272_), .A1(new_n6937_), .B0(new_n4272_), .B1(new_n2918_), .Y(new_n9275_));
  AOI22X1  g09082(.A0(new_n9275_), .A1(new_n9272_), .B0(new_n9274_), .B1(new_n6937_), .Y(new_n9276_));
  XOR2X1   g09083(.A(new_n9276_), .B(new_n9270_), .Y(new_n9277_));
  NOR2X1   g09084(.A(new_n9223_), .B(new_n9220_), .Y(new_n9278_));
  AOI21X1  g09085(.A0(new_n9227_), .A1(new_n9224_), .B0(new_n9278_), .Y(new_n9279_));
  XOR2X1   g09086(.A(new_n9279_), .B(new_n9277_), .Y(new_n9280_));
  NAND4X1  g09087(.A(\a[63] ), .B(\a[60] ), .C(\a[21] ), .D(\a[18] ), .Y(new_n9281_));
  NAND4X1  g09088(.A(\a[63] ), .B(\a[61] ), .C(\a[20] ), .D(\a[18] ), .Y(new_n9282_));
  AOI22X1  g09089(.A0(new_n9282_), .A1(new_n9281_), .B0(new_n6428_), .B1(new_n1236_), .Y(new_n9283_));
  NAND4X1  g09090(.A(\a[61] ), .B(\a[60] ), .C(\a[21] ), .D(\a[20] ), .Y(new_n9284_));
  NAND3X1  g09091(.A(new_n9282_), .B(new_n9281_), .C(new_n9284_), .Y(new_n9285_));
  AOI22X1  g09092(.A0(\a[61] ), .A1(\a[20] ), .B0(\a[60] ), .B1(\a[21] ), .Y(new_n9286_));
  NAND2X1  g09093(.A(\a[63] ), .B(\a[18] ), .Y(new_n9287_));
  OAI22X1  g09094(.A0(new_n9287_), .A1(new_n9283_), .B0(new_n9286_), .B1(new_n9285_), .Y(new_n9288_));
  NAND2X1  g09095(.A(\a[46] ), .B(\a[35] ), .Y(new_n9289_));
  NAND4X1  g09096(.A(\a[46] ), .B(\a[45] ), .C(\a[36] ), .D(\a[35] ), .Y(new_n9290_));
  NAND4X1  g09097(.A(\a[46] ), .B(\a[44] ), .C(\a[37] ), .D(\a[35] ), .Y(new_n9291_));
  AOI22X1  g09098(.A0(new_n9291_), .A1(new_n9290_), .B0(new_n3918_), .B1(new_n3330_), .Y(new_n9292_));
  AOI22X1  g09099(.A0(\a[45] ), .A1(\a[36] ), .B0(\a[44] ), .B1(\a[37] ), .Y(new_n9293_));
  AOI21X1  g09100(.A0(new_n3918_), .A1(new_n3330_), .B0(new_n9292_), .Y(new_n9294_));
  INVX1    g09101(.A(new_n9294_), .Y(new_n9295_));
  OAI22X1  g09102(.A0(new_n9295_), .A1(new_n9293_), .B0(new_n9292_), .B1(new_n9289_), .Y(new_n9296_));
  XOR2X1   g09103(.A(new_n9296_), .B(new_n9288_), .Y(new_n9297_));
  AOI22X1  g09104(.A0(new_n8939_), .A1(\a[29] ), .B0(new_n1996_), .B1(\a[53] ), .Y(new_n9298_));
  AND2X1   g09105(.A(new_n5048_), .B(new_n1674_), .Y(new_n9299_));
  NOR3X1   g09106(.A(new_n9299_), .B(new_n9298_), .C(new_n4906_), .Y(new_n9300_));
  AND2X1   g09107(.A(\a[55] ), .B(\a[26] ), .Y(new_n9301_));
  INVX1    g09108(.A(new_n9301_), .Y(new_n9302_));
  AOI22X1  g09109(.A0(\a[53] ), .A1(\a[28] ), .B0(\a[52] ), .B1(\a[29] ), .Y(new_n9303_));
  NOR2X1   g09110(.A(new_n9300_), .B(new_n9299_), .Y(new_n9304_));
  INVX1    g09111(.A(new_n9304_), .Y(new_n9305_));
  OAI22X1  g09112(.A0(new_n9305_), .A1(new_n9303_), .B0(new_n9302_), .B1(new_n9300_), .Y(new_n9306_));
  INVX1    g09113(.A(new_n9306_), .Y(new_n9307_));
  XOR2X1   g09114(.A(new_n9307_), .B(new_n9297_), .Y(new_n9308_));
  XOR2X1   g09115(.A(new_n9308_), .B(new_n9280_), .Y(new_n9309_));
  XOR2X1   g09116(.A(new_n9309_), .B(new_n9255_), .Y(new_n9310_));
  XOR2X1   g09117(.A(new_n9310_), .B(new_n9253_), .Y(new_n9311_));
  XOR2X1   g09118(.A(new_n9311_), .B(new_n9251_), .Y(new_n9312_));
  AND2X1   g09119(.A(new_n9181_), .B(new_n9119_), .Y(new_n9313_));
  AOI21X1  g09120(.A0(new_n9182_), .A1(new_n9116_), .B0(new_n9313_), .Y(new_n9314_));
  NOR2X1   g09121(.A(new_n9014_), .B(new_n9004_), .Y(new_n9315_));
  AOI21X1  g09122(.A0(new_n9206_), .A1(new_n9205_), .B0(new_n9315_), .Y(new_n9316_));
  AND2X1   g09123(.A(\a[54] ), .B(\a[27] ), .Y(new_n9317_));
  AND2X1   g09124(.A(new_n3503_), .B(new_n3462_), .Y(new_n9318_));
  AOI22X1  g09125(.A0(\a[43] ), .A1(\a[38] ), .B0(\a[42] ), .B1(\a[39] ), .Y(new_n9319_));
  OAI21X1  g09126(.A0(new_n9319_), .A1(new_n9318_), .B0(new_n9317_), .Y(new_n9320_));
  INVX1    g09127(.A(new_n9319_), .Y(new_n9321_));
  AOI21X1  g09128(.A0(new_n9321_), .A1(new_n9317_), .B0(new_n9318_), .Y(new_n9322_));
  NAND2X1  g09129(.A(new_n9322_), .B(new_n9321_), .Y(new_n9323_));
  AND2X1   g09130(.A(new_n9323_), .B(new_n9320_), .Y(new_n9324_));
  XOR2X1   g09131(.A(new_n9324_), .B(new_n9316_), .Y(new_n9325_));
  AND2X1   g09132(.A(new_n8977_), .B(new_n9070_), .Y(new_n9326_));
  AOI21X1  g09133(.A0(new_n9193_), .A1(new_n9192_), .B0(new_n9326_), .Y(new_n9327_));
  XOR2X1   g09134(.A(new_n9327_), .B(new_n9325_), .Y(new_n9328_));
  NAND2X1  g09135(.A(new_n9197_), .B(new_n9194_), .Y(new_n9329_));
  OAI21X1  g09136(.A0(new_n9200_), .A1(new_n9199_), .B0(new_n9198_), .Y(new_n9330_));
  NAND2X1  g09137(.A(new_n9330_), .B(new_n9329_), .Y(new_n9331_));
  AND2X1   g09138(.A(new_n9214_), .B(new_n9211_), .Y(new_n9332_));
  AOI21X1  g09139(.A0(new_n9215_), .A1(new_n9207_), .B0(new_n9332_), .Y(new_n9333_));
  XOR2X1   g09140(.A(new_n9333_), .B(new_n9331_), .Y(new_n9334_));
  XOR2X1   g09141(.A(new_n9334_), .B(new_n9328_), .Y(new_n9335_));
  XOR2X1   g09142(.A(new_n9335_), .B(new_n9314_), .Y(new_n9336_));
  NOR2X1   g09143(.A(new_n9138_), .B(new_n8997_), .Y(new_n9337_));
  AOI21X1  g09144(.A0(new_n6556_), .A1(new_n855_), .B0(new_n9337_), .Y(new_n9338_));
  XOR2X1   g09145(.A(new_n9338_), .B(new_n9132_), .Y(new_n9339_));
  OAI22X1  g09146(.A0(new_n7653_), .A1(new_n4923_), .B0(new_n7651_), .B1(new_n2076_), .Y(new_n9340_));
  OAI21X1  g09147(.A0(new_n7652_), .A1(new_n2672_), .B0(new_n9340_), .Y(new_n9341_));
  AND2X1   g09148(.A(\a[51] ), .B(\a[30] ), .Y(new_n9342_));
  AOI21X1  g09149(.A0(new_n4321_), .A1(new_n2671_), .B0(new_n9340_), .Y(new_n9343_));
  OAI22X1  g09150(.A0(new_n4983_), .A1(new_n1704_), .B0(new_n3915_), .B1(new_n2219_), .Y(new_n9344_));
  AOI22X1  g09151(.A0(new_n9344_), .A1(new_n9343_), .B0(new_n9342_), .B1(new_n9341_), .Y(new_n9345_));
  XOR2X1   g09152(.A(new_n9345_), .B(new_n9339_), .Y(new_n9346_));
  XOR2X1   g09153(.A(new_n9152_), .B(new_n9126_), .Y(new_n9347_));
  OAI21X1  g09154(.A0(new_n6793_), .A1(new_n1397_), .B0(new_n9143_), .Y(new_n9348_));
  XOR2X1   g09155(.A(new_n9348_), .B(new_n9347_), .Y(new_n9349_));
  INVX1    g09156(.A(new_n9349_), .Y(new_n9350_));
  INVX1    g09157(.A(new_n9128_), .Y(new_n9351_));
  OR2X1    g09158(.A(new_n9134_), .B(new_n9351_), .Y(new_n9352_));
  OAI21X1  g09159(.A0(new_n9139_), .A1(new_n9135_), .B0(new_n9352_), .Y(new_n9353_));
  XOR2X1   g09160(.A(new_n9353_), .B(new_n9350_), .Y(new_n9354_));
  XOR2X1   g09161(.A(new_n9354_), .B(new_n9346_), .Y(new_n9355_));
  INVX1    g09162(.A(new_n9355_), .Y(new_n9356_));
  INVX1    g09163(.A(new_n9179_), .Y(new_n9357_));
  OR2X1    g09164(.A(new_n9180_), .B(new_n9141_), .Y(new_n9358_));
  OAI21X1  g09165(.A0(new_n9357_), .A1(new_n9155_), .B0(new_n9358_), .Y(new_n9359_));
  XOR2X1   g09166(.A(new_n9359_), .B(new_n9356_), .Y(new_n9360_));
  INVX1    g09167(.A(new_n9160_), .Y(new_n9361_));
  XOR2X1   g09168(.A(new_n9177_), .B(new_n9169_), .Y(new_n9362_));
  XOR2X1   g09169(.A(new_n9362_), .B(new_n9361_), .Y(new_n9363_));
  INVX1    g09170(.A(new_n9363_), .Y(new_n9364_));
  AND2X1   g09171(.A(new_n9160_), .B(new_n9156_), .Y(new_n9365_));
  OAI21X1  g09172(.A0(new_n9161_), .A1(new_n9365_), .B0(new_n9171_), .Y(new_n9366_));
  OAI21X1  g09173(.A0(new_n9178_), .A1(new_n9172_), .B0(new_n9366_), .Y(new_n9367_));
  OR2X1    g09174(.A(new_n9147_), .B(new_n8985_), .Y(new_n9368_));
  AND2X1   g09175(.A(new_n9147_), .B(new_n8985_), .Y(new_n9369_));
  OAI21X1  g09176(.A0(new_n9154_), .A1(new_n9369_), .B0(new_n9368_), .Y(new_n9370_));
  XOR2X1   g09177(.A(new_n9370_), .B(new_n9367_), .Y(new_n9371_));
  XOR2X1   g09178(.A(new_n9371_), .B(new_n9364_), .Y(new_n9372_));
  XOR2X1   g09179(.A(new_n9372_), .B(new_n9360_), .Y(new_n9373_));
  XOR2X1   g09180(.A(new_n9373_), .B(new_n9336_), .Y(new_n9374_));
  XOR2X1   g09181(.A(new_n9374_), .B(new_n9312_), .Y(new_n9375_));
  AND2X1   g09182(.A(new_n9183_), .B(new_n9113_), .Y(new_n9376_));
  AOI21X1  g09183(.A0(new_n9236_), .A1(new_n9184_), .B0(new_n9376_), .Y(new_n9377_));
  NOR2X1   g09184(.A(new_n9377_), .B(new_n9375_), .Y(new_n9378_));
  AND2X1   g09185(.A(new_n9377_), .B(new_n9375_), .Y(new_n9379_));
  OR2X1    g09186(.A(new_n9379_), .B(new_n9378_), .Y(new_n9380_));
  XOR2X1   g09187(.A(new_n9380_), .B(new_n9249_), .Y(\asquared[82] ));
  INVX1    g09188(.A(new_n9378_), .Y(new_n9382_));
  OAI21X1  g09189(.A0(new_n9379_), .A1(new_n9249_), .B0(new_n9382_), .Y(new_n9383_));
  AND2X1   g09190(.A(new_n9311_), .B(new_n9251_), .Y(new_n9384_));
  INVX1    g09191(.A(new_n9374_), .Y(new_n9385_));
  AOI21X1  g09192(.A0(new_n9385_), .A1(new_n9312_), .B0(new_n9384_), .Y(new_n9386_));
  INVX1    g09193(.A(new_n9314_), .Y(new_n9387_));
  AND2X1   g09194(.A(new_n9335_), .B(new_n9387_), .Y(new_n9388_));
  INVX1    g09195(.A(new_n9336_), .Y(new_n9389_));
  AOI21X1  g09196(.A0(new_n9373_), .A1(new_n9389_), .B0(new_n9388_), .Y(new_n9390_));
  NAND2X1  g09197(.A(new_n9359_), .B(new_n9355_), .Y(new_n9391_));
  OAI21X1  g09198(.A0(new_n9372_), .A1(new_n9360_), .B0(new_n9391_), .Y(new_n9392_));
  INVX1    g09199(.A(new_n9333_), .Y(new_n9393_));
  NAND2X1  g09200(.A(new_n9393_), .B(new_n9331_), .Y(new_n9394_));
  OAI21X1  g09201(.A0(new_n9334_), .A1(new_n9328_), .B0(new_n9394_), .Y(new_n9395_));
  NOR4X1   g09202(.A(new_n6023_), .B(new_n4349_), .C(new_n1704_), .D(new_n1098_), .Y(new_n9396_));
  NAND4X1  g09203(.A(\a[62] ), .B(\a[51] ), .C(\a[31] ), .D(\a[20] ), .Y(new_n9397_));
  NAND4X1  g09204(.A(\a[62] ), .B(\a[61] ), .C(\a[21] ), .D(\a[20] ), .Y(new_n9398_));
  AOI21X1  g09205(.A0(new_n9398_), .A1(new_n9397_), .B0(new_n9396_), .Y(new_n9399_));
  OR2X1    g09206(.A(new_n9399_), .B(new_n9396_), .Y(new_n9400_));
  AOI22X1  g09207(.A0(\a[61] ), .A1(\a[21] ), .B0(\a[51] ), .B1(\a[31] ), .Y(new_n9401_));
  NAND2X1  g09208(.A(\a[62] ), .B(\a[20] ), .Y(new_n9402_));
  OAI22X1  g09209(.A0(new_n9402_), .A1(new_n9399_), .B0(new_n9401_), .B1(new_n9400_), .Y(new_n9403_));
  NAND4X1  g09210(.A(\a[50] ), .B(\a[48] ), .C(\a[34] ), .D(\a[32] ), .Y(new_n9404_));
  NAND4X1  g09211(.A(\a[50] ), .B(\a[49] ), .C(\a[33] ), .D(\a[32] ), .Y(new_n9405_));
  AOI22X1  g09212(.A0(new_n9405_), .A1(new_n9404_), .B0(new_n4274_), .B1(new_n2918_), .Y(new_n9406_));
  NAND2X1  g09213(.A(\a[50] ), .B(\a[32] ), .Y(new_n9407_));
  NAND4X1  g09214(.A(\a[49] ), .B(\a[48] ), .C(\a[34] ), .D(\a[33] ), .Y(new_n9408_));
  NAND3X1  g09215(.A(new_n9405_), .B(new_n9404_), .C(new_n9408_), .Y(new_n9409_));
  AOI22X1  g09216(.A0(\a[49] ), .A1(\a[33] ), .B0(\a[48] ), .B1(\a[34] ), .Y(new_n9410_));
  OAI22X1  g09217(.A0(new_n9410_), .A1(new_n9409_), .B0(new_n9407_), .B1(new_n9406_), .Y(new_n9411_));
  XOR2X1   g09218(.A(new_n9411_), .B(new_n9403_), .Y(new_n9412_));
  AOI22X1  g09219(.A0(new_n6795_), .A1(new_n1530_), .B0(new_n6427_), .B1(new_n1394_), .Y(new_n9413_));
  AOI21X1  g09220(.A0(new_n6121_), .A1(new_n1219_), .B0(new_n9413_), .Y(new_n9414_));
  AND2X1   g09221(.A(\a[60] ), .B(\a[22] ), .Y(new_n9415_));
  INVX1    g09222(.A(new_n9415_), .Y(new_n9416_));
  OAI22X1  g09223(.A0(new_n6796_), .A1(new_n1531_), .B0(new_n6794_), .B1(new_n1395_), .Y(new_n9417_));
  AOI21X1  g09224(.A0(new_n6121_), .A1(new_n1219_), .B0(new_n9417_), .Y(new_n9418_));
  INVX1    g09225(.A(new_n9418_), .Y(new_n9419_));
  AOI22X1  g09226(.A0(\a[59] ), .A1(\a[23] ), .B0(\a[58] ), .B1(\a[24] ), .Y(new_n9420_));
  OAI22X1  g09227(.A0(new_n9420_), .A1(new_n9419_), .B0(new_n9416_), .B1(new_n9414_), .Y(new_n9421_));
  XOR2X1   g09228(.A(new_n9421_), .B(new_n9412_), .Y(new_n9422_));
  INVX1    g09229(.A(new_n9422_), .Y(new_n9423_));
  OR2X1    g09230(.A(new_n9324_), .B(new_n9316_), .Y(new_n9424_));
  INVX1    g09231(.A(new_n9325_), .Y(new_n9425_));
  OAI21X1  g09232(.A0(new_n9327_), .A1(new_n9425_), .B0(new_n9424_), .Y(new_n9426_));
  XOR2X1   g09233(.A(new_n9426_), .B(new_n9423_), .Y(new_n9427_));
  AOI22X1  g09234(.A0(\a[44] ), .A1(\a[38] ), .B0(\a[43] ), .B1(\a[39] ), .Y(new_n9428_));
  AND2X1   g09235(.A(\a[56] ), .B(\a[26] ), .Y(new_n9429_));
  INVX1    g09236(.A(new_n9429_), .Y(new_n9430_));
  AND2X1   g09237(.A(new_n4992_), .B(new_n3503_), .Y(new_n9431_));
  NOR3X1   g09238(.A(new_n9430_), .B(new_n9431_), .C(new_n9428_), .Y(new_n9432_));
  NOR2X1   g09239(.A(new_n9432_), .B(new_n9431_), .Y(new_n9433_));
  INVX1    g09240(.A(new_n9433_), .Y(new_n9434_));
  OAI22X1  g09241(.A0(new_n9434_), .A1(new_n9428_), .B0(new_n9432_), .B1(new_n9430_), .Y(new_n9435_));
  AOI22X1  g09242(.A0(\a[53] ), .A1(\a[29] ), .B0(\a[52] ), .B1(\a[30] ), .Y(new_n9436_));
  INVX1    g09243(.A(new_n9436_), .Y(new_n9437_));
  NAND4X1  g09244(.A(\a[53] ), .B(\a[52] ), .C(\a[30] ), .D(\a[29] ), .Y(new_n9438_));
  AOI21X1  g09245(.A0(new_n9437_), .A1(new_n9438_), .B0(new_n8071_), .Y(new_n9439_));
  AOI22X1  g09246(.A0(new_n9437_), .A1(new_n8070_), .B0(new_n5048_), .B1(new_n2196_), .Y(new_n9440_));
  AOI21X1  g09247(.A0(new_n9440_), .A1(new_n9437_), .B0(new_n9439_), .Y(new_n9441_));
  XOR2X1   g09248(.A(new_n9441_), .B(new_n9435_), .Y(new_n9442_));
  NAND4X1  g09249(.A(\a[47] ), .B(\a[45] ), .C(\a[37] ), .D(\a[35] ), .Y(new_n9443_));
  NAND4X1  g09250(.A(\a[47] ), .B(\a[46] ), .C(\a[36] ), .D(\a[35] ), .Y(new_n9444_));
  AOI22X1  g09251(.A0(new_n9444_), .A1(new_n9443_), .B0(new_n3809_), .B1(new_n3330_), .Y(new_n9445_));
  NOR3X1   g09252(.A(new_n9445_), .B(new_n4041_), .C(new_n2557_), .Y(new_n9446_));
  AOI21X1  g09253(.A0(new_n3809_), .A1(new_n3330_), .B0(new_n9445_), .Y(new_n9447_));
  OAI22X1  g09254(.A0(new_n3460_), .A1(new_n2583_), .B0(new_n3811_), .B1(new_n2345_), .Y(new_n9448_));
  AOI21X1  g09255(.A0(new_n9448_), .A1(new_n9447_), .B0(new_n9446_), .Y(new_n9449_));
  XOR2X1   g09256(.A(new_n9449_), .B(new_n9442_), .Y(new_n9450_));
  INVX1    g09257(.A(new_n9450_), .Y(new_n9451_));
  XOR2X1   g09258(.A(new_n9451_), .B(new_n9427_), .Y(new_n9452_));
  XOR2X1   g09259(.A(new_n9452_), .B(new_n9395_), .Y(new_n9453_));
  XOR2X1   g09260(.A(new_n9453_), .B(new_n9392_), .Y(new_n9454_));
  XOR2X1   g09261(.A(new_n9454_), .B(new_n9390_), .Y(new_n9455_));
  NOR2X1   g09262(.A(new_n9309_), .B(new_n9255_), .Y(new_n9456_));
  AOI21X1  g09263(.A0(new_n9310_), .A1(new_n9253_), .B0(new_n9456_), .Y(new_n9457_));
  NOR2X1   g09264(.A(new_n9152_), .B(new_n9126_), .Y(new_n9458_));
  AOI21X1  g09265(.A0(new_n9348_), .A1(new_n9347_), .B0(new_n9458_), .Y(new_n9459_));
  INVX1    g09266(.A(new_n4826_), .Y(new_n9460_));
  AND2X1   g09267(.A(\a[57] ), .B(\a[55] ), .Y(new_n9461_));
  NAND4X1  g09268(.A(\a[55] ), .B(\a[54] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n9462_));
  NAND4X1  g09269(.A(\a[57] ), .B(\a[54] ), .C(\a[28] ), .D(\a[25] ), .Y(new_n9463_));
  AOI22X1  g09270(.A0(new_n9463_), .A1(new_n9462_), .B0(new_n9461_), .B1(new_n1871_), .Y(new_n9464_));
  AOI22X1  g09271(.A0(\a[57] ), .A1(\a[25] ), .B0(\a[55] ), .B1(\a[27] ), .Y(new_n9465_));
  AOI21X1  g09272(.A0(new_n9461_), .A1(new_n1871_), .B0(new_n9464_), .Y(new_n9466_));
  INVX1    g09273(.A(new_n9466_), .Y(new_n9467_));
  OAI22X1  g09274(.A0(new_n9467_), .A1(new_n9465_), .B0(new_n9464_), .B1(new_n9460_), .Y(new_n9468_));
  XOR2X1   g09275(.A(new_n9468_), .B(new_n9459_), .Y(new_n9469_));
  NOR2X1   g09276(.A(new_n9177_), .B(new_n9169_), .Y(new_n9470_));
  AOI21X1  g09277(.A0(new_n9362_), .A1(new_n9361_), .B0(new_n9470_), .Y(new_n9471_));
  XOR2X1   g09278(.A(new_n9471_), .B(new_n9469_), .Y(new_n9472_));
  NAND2X1  g09279(.A(new_n9353_), .B(new_n9349_), .Y(new_n9473_));
  OAI21X1  g09280(.A0(new_n9354_), .A1(new_n9346_), .B0(new_n9473_), .Y(new_n9474_));
  AND2X1   g09281(.A(new_n9370_), .B(new_n9367_), .Y(new_n9475_));
  AOI21X1  g09282(.A0(new_n9371_), .A1(new_n9363_), .B0(new_n9475_), .Y(new_n9476_));
  XOR2X1   g09283(.A(new_n9476_), .B(new_n9474_), .Y(new_n9477_));
  XOR2X1   g09284(.A(new_n9477_), .B(new_n9472_), .Y(new_n9478_));
  XOR2X1   g09285(.A(new_n9478_), .B(new_n9457_), .Y(new_n9479_));
  NOR2X1   g09286(.A(new_n9279_), .B(new_n9277_), .Y(new_n9480_));
  INVX1    g09287(.A(new_n9480_), .Y(new_n9481_));
  INVX1    g09288(.A(new_n9280_), .Y(new_n9482_));
  OAI21X1  g09289(.A0(new_n9308_), .A1(new_n9482_), .B0(new_n9481_), .Y(new_n9483_));
  XOR2X1   g09290(.A(new_n9343_), .B(new_n9275_), .Y(new_n9484_));
  XOR2X1   g09291(.A(new_n9484_), .B(new_n9305_), .Y(new_n9485_));
  XOR2X1   g09292(.A(new_n9285_), .B(new_n9267_), .Y(new_n9486_));
  XOR2X1   g09293(.A(new_n9486_), .B(new_n9294_), .Y(new_n9487_));
  AND2X1   g09294(.A(new_n9296_), .B(new_n9288_), .Y(new_n9488_));
  AOI21X1  g09295(.A0(new_n9306_), .A1(new_n9297_), .B0(new_n9488_), .Y(new_n9489_));
  XOR2X1   g09296(.A(new_n9489_), .B(new_n9487_), .Y(new_n9490_));
  XOR2X1   g09297(.A(new_n9490_), .B(new_n9485_), .Y(new_n9491_));
  XOR2X1   g09298(.A(new_n9491_), .B(new_n9483_), .Y(new_n9492_));
  AND2X1   g09299(.A(new_n9338_), .B(new_n9132_), .Y(new_n9493_));
  OR2X1    g09300(.A(new_n9338_), .B(new_n9132_), .Y(new_n9494_));
  OAI21X1  g09301(.A0(new_n9345_), .A1(new_n9493_), .B0(new_n9494_), .Y(new_n9495_));
  AND2X1   g09302(.A(new_n9269_), .B(new_n9261_), .Y(new_n9496_));
  INVX1    g09303(.A(new_n9496_), .Y(new_n9497_));
  INVX1    g09304(.A(new_n9270_), .Y(new_n9498_));
  OAI21X1  g09305(.A0(new_n9276_), .A1(new_n9498_), .B0(new_n9497_), .Y(new_n9499_));
  INVX1    g09306(.A(new_n9499_), .Y(new_n9500_));
  XOR2X1   g09307(.A(new_n9500_), .B(new_n9495_), .Y(new_n9501_));
  INVX1    g09308(.A(new_n8425_), .Y(new_n9502_));
  XOR2X1   g09309(.A(new_n9257_), .B(new_n9502_), .Y(new_n9503_));
  XOR2X1   g09310(.A(new_n9503_), .B(new_n9322_), .Y(new_n9504_));
  XOR2X1   g09311(.A(new_n9504_), .B(new_n9501_), .Y(new_n9505_));
  XOR2X1   g09312(.A(new_n9505_), .B(new_n9492_), .Y(new_n9506_));
  XOR2X1   g09313(.A(new_n9506_), .B(new_n9479_), .Y(new_n9507_));
  XOR2X1   g09314(.A(new_n9507_), .B(new_n9455_), .Y(new_n9508_));
  XOR2X1   g09315(.A(new_n9508_), .B(new_n9386_), .Y(new_n9509_));
  XOR2X1   g09316(.A(new_n9509_), .B(new_n9383_), .Y(\asquared[83] ));
  INVX1    g09317(.A(new_n9454_), .Y(new_n9511_));
  NOR2X1   g09318(.A(new_n9511_), .B(new_n9390_), .Y(new_n9512_));
  INVX1    g09319(.A(new_n9455_), .Y(new_n9513_));
  AOI21X1  g09320(.A0(new_n9507_), .A1(new_n9513_), .B0(new_n9512_), .Y(new_n9514_));
  NOR2X1   g09321(.A(new_n9478_), .B(new_n9457_), .Y(new_n9515_));
  AOI21X1  g09322(.A0(new_n9506_), .A1(new_n9479_), .B0(new_n9515_), .Y(new_n9516_));
  AND2X1   g09323(.A(new_n9491_), .B(new_n9483_), .Y(new_n9517_));
  AOI21X1  g09324(.A0(new_n9505_), .A1(new_n9492_), .B0(new_n9517_), .Y(new_n9518_));
  INVX1    g09325(.A(new_n9518_), .Y(new_n9519_));
  INVX1    g09326(.A(new_n9472_), .Y(new_n9520_));
  INVX1    g09327(.A(new_n9476_), .Y(new_n9521_));
  NAND2X1  g09328(.A(new_n9521_), .B(new_n9474_), .Y(new_n9522_));
  OAI21X1  g09329(.A0(new_n9477_), .A1(new_n9520_), .B0(new_n9522_), .Y(new_n9523_));
  NAND3X1  g09330(.A(\a[62] ), .B(\a[42] ), .C(\a[21] ), .Y(new_n9524_));
  AND2X1   g09331(.A(new_n9524_), .B(new_n8069_), .Y(new_n9525_));
  OAI21X1  g09332(.A0(new_n6606_), .A1(new_n1098_), .B0(new_n3096_), .Y(new_n9526_));
  NOR3X1   g09333(.A(new_n9524_), .B(new_n3096_), .C(new_n3081_), .Y(new_n9527_));
  AOI21X1  g09334(.A0(new_n9526_), .A1(new_n9525_), .B0(new_n9527_), .Y(new_n9528_));
  AOI22X1  g09335(.A0(\a[44] ), .A1(\a[39] ), .B0(\a[43] ), .B1(\a[40] ), .Y(new_n9529_));
  AND2X1   g09336(.A(\a[54] ), .B(\a[29] ), .Y(new_n9530_));
  AND2X1   g09337(.A(new_n4992_), .B(new_n4077_), .Y(new_n9531_));
  OAI21X1  g09338(.A0(new_n9529_), .A1(new_n9531_), .B0(new_n9530_), .Y(new_n9532_));
  NOR3X1   g09339(.A(new_n9529_), .B(new_n4835_), .C(new_n1803_), .Y(new_n9533_));
  OR2X1    g09340(.A(new_n9533_), .B(new_n9531_), .Y(new_n9534_));
  OAI21X1  g09341(.A0(new_n9534_), .A1(new_n9529_), .B0(new_n9532_), .Y(new_n9535_));
  XOR2X1   g09342(.A(new_n9535_), .B(new_n9528_), .Y(new_n9536_));
  OAI22X1  g09343(.A0(new_n7652_), .A1(new_n2919_), .B0(new_n8802_), .B1(new_n4914_), .Y(new_n9537_));
  OAI21X1  g09344(.A0(new_n4280_), .A1(new_n4915_), .B0(new_n9537_), .Y(new_n9538_));
  AND2X1   g09345(.A(\a[50] ), .B(\a[33] ), .Y(new_n9539_));
  AOI21X1  g09346(.A0(new_n4274_), .A1(new_n2361_), .B0(new_n9537_), .Y(new_n9540_));
  OAI22X1  g09347(.A0(new_n3915_), .A1(new_n2028_), .B0(new_n3926_), .B1(new_n2557_), .Y(new_n9541_));
  AOI22X1  g09348(.A0(new_n9541_), .A1(new_n9540_), .B0(new_n9539_), .B1(new_n9538_), .Y(new_n9542_));
  XOR2X1   g09349(.A(new_n9542_), .B(new_n9536_), .Y(new_n9543_));
  INVX1    g09350(.A(new_n9543_), .Y(new_n9544_));
  INVX1    g09351(.A(new_n9468_), .Y(new_n9545_));
  OR2X1    g09352(.A(new_n9545_), .B(new_n9459_), .Y(new_n9546_));
  OAI21X1  g09353(.A0(new_n9471_), .A1(new_n9469_), .B0(new_n9546_), .Y(new_n9547_));
  XOR2X1   g09354(.A(new_n9547_), .B(new_n9544_), .Y(new_n9548_));
  AOI22X1  g09355(.A0(\a[57] ), .A1(\a[26] ), .B0(\a[51] ), .B1(\a[32] ), .Y(new_n9549_));
  AND2X1   g09356(.A(\a[57] ), .B(\a[51] ), .Y(new_n9550_));
  NAND4X1  g09357(.A(\a[58] ), .B(\a[57] ), .C(\a[26] ), .D(\a[25] ), .Y(new_n9551_));
  NAND4X1  g09358(.A(\a[58] ), .B(\a[51] ), .C(\a[32] ), .D(\a[25] ), .Y(new_n9552_));
  AOI22X1  g09359(.A0(new_n9552_), .A1(new_n9551_), .B0(new_n9550_), .B1(new_n2318_), .Y(new_n9553_));
  AOI21X1  g09360(.A0(new_n9550_), .A1(new_n2318_), .B0(new_n9553_), .Y(new_n9554_));
  INVX1    g09361(.A(new_n9554_), .Y(new_n9555_));
  NAND2X1  g09362(.A(\a[58] ), .B(\a[25] ), .Y(new_n9556_));
  OAI22X1  g09363(.A0(new_n9556_), .A1(new_n9553_), .B0(new_n9555_), .B1(new_n9549_), .Y(new_n9557_));
  NAND4X1  g09364(.A(\a[47] ), .B(\a[45] ), .C(\a[38] ), .D(\a[36] ), .Y(new_n9558_));
  NAND4X1  g09365(.A(\a[47] ), .B(\a[46] ), .C(\a[37] ), .D(\a[36] ), .Y(new_n9559_));
  AOI22X1  g09366(.A0(new_n9559_), .A1(new_n9558_), .B0(new_n3809_), .B1(new_n3164_), .Y(new_n9560_));
  NAND2X1  g09367(.A(\a[47] ), .B(\a[36] ), .Y(new_n9561_));
  NAND4X1  g09368(.A(\a[46] ), .B(\a[45] ), .C(\a[38] ), .D(\a[37] ), .Y(new_n9562_));
  NAND3X1  g09369(.A(new_n9559_), .B(new_n9558_), .C(new_n9562_), .Y(new_n9563_));
  AOI22X1  g09370(.A0(\a[46] ), .A1(\a[37] ), .B0(\a[45] ), .B1(\a[38] ), .Y(new_n9564_));
  OAI22X1  g09371(.A0(new_n9564_), .A1(new_n9563_), .B0(new_n9561_), .B1(new_n9560_), .Y(new_n9565_));
  XOR2X1   g09372(.A(new_n9565_), .B(new_n9557_), .Y(new_n9566_));
  INVX1    g09373(.A(new_n9073_), .Y(new_n9567_));
  AOI22X1  g09374(.A0(\a[63] ), .A1(\a[20] ), .B0(\a[61] ), .B1(\a[22] ), .Y(new_n9568_));
  AND2X1   g09375(.A(new_n6688_), .B(new_n2134_), .Y(new_n9569_));
  NOR3X1   g09376(.A(new_n9568_), .B(new_n9569_), .C(new_n9567_), .Y(new_n9570_));
  INVX1    g09377(.A(new_n9568_), .Y(new_n9571_));
  AOI21X1  g09378(.A0(new_n9571_), .A1(new_n9073_), .B0(new_n9569_), .Y(new_n9572_));
  INVX1    g09379(.A(new_n9572_), .Y(new_n9573_));
  OAI22X1  g09380(.A0(new_n9573_), .A1(new_n9568_), .B0(new_n9570_), .B1(new_n9567_), .Y(new_n9574_));
  INVX1    g09381(.A(new_n9574_), .Y(new_n9575_));
  XOR2X1   g09382(.A(new_n9575_), .B(new_n9566_), .Y(new_n9576_));
  XOR2X1   g09383(.A(new_n9576_), .B(new_n9548_), .Y(new_n9577_));
  XOR2X1   g09384(.A(new_n9577_), .B(new_n9523_), .Y(new_n9578_));
  XOR2X1   g09385(.A(new_n9578_), .B(new_n9519_), .Y(new_n9579_));
  INVX1    g09386(.A(new_n9579_), .Y(new_n9580_));
  XOR2X1   g09387(.A(new_n9580_), .B(new_n9516_), .Y(new_n9581_));
  AND2X1   g09388(.A(new_n9426_), .B(new_n9422_), .Y(new_n9582_));
  NOR2X1   g09389(.A(new_n9451_), .B(new_n9427_), .Y(new_n9583_));
  NOR2X1   g09390(.A(new_n9583_), .B(new_n9582_), .Y(new_n9584_));
  INVX1    g09391(.A(new_n9584_), .Y(new_n9585_));
  NOR2X1   g09392(.A(new_n9489_), .B(new_n9487_), .Y(new_n9586_));
  AOI21X1  g09393(.A0(new_n9490_), .A1(new_n9485_), .B0(new_n9586_), .Y(new_n9587_));
  XOR2X1   g09394(.A(new_n9587_), .B(new_n9585_), .Y(new_n9588_));
  XOR2X1   g09395(.A(new_n9447_), .B(new_n9418_), .Y(new_n9589_));
  XOR2X1   g09396(.A(new_n9589_), .B(new_n9434_), .Y(new_n9590_));
  INVX1    g09397(.A(new_n9590_), .Y(new_n9591_));
  XOR2X1   g09398(.A(new_n9409_), .B(new_n9400_), .Y(new_n9592_));
  XOR2X1   g09399(.A(new_n9592_), .B(new_n9467_), .Y(new_n9593_));
  AND2X1   g09400(.A(new_n9440_), .B(new_n9437_), .Y(new_n9594_));
  OAI21X1  g09401(.A0(new_n9594_), .A1(new_n9439_), .B0(new_n9435_), .Y(new_n9595_));
  OR2X1    g09402(.A(new_n9449_), .B(new_n9442_), .Y(new_n9596_));
  AND2X1   g09403(.A(new_n9596_), .B(new_n9595_), .Y(new_n9597_));
  XOR2X1   g09404(.A(new_n9597_), .B(new_n9593_), .Y(new_n9598_));
  XOR2X1   g09405(.A(new_n9598_), .B(new_n9591_), .Y(new_n9599_));
  XOR2X1   g09406(.A(new_n9599_), .B(new_n9588_), .Y(new_n9600_));
  AND2X1   g09407(.A(new_n9452_), .B(new_n9395_), .Y(new_n9601_));
  AOI21X1  g09408(.A0(new_n9453_), .A1(new_n9392_), .B0(new_n9601_), .Y(new_n9602_));
  NOR2X1   g09409(.A(new_n9343_), .B(new_n9275_), .Y(new_n9603_));
  AOI21X1  g09410(.A0(new_n9484_), .A1(new_n9305_), .B0(new_n9603_), .Y(new_n9604_));
  AND2X1   g09411(.A(new_n9285_), .B(new_n9267_), .Y(new_n9605_));
  AOI21X1  g09412(.A0(new_n9486_), .A1(new_n9295_), .B0(new_n9605_), .Y(new_n9606_));
  XOR2X1   g09413(.A(new_n9606_), .B(new_n9604_), .Y(new_n9607_));
  AND2X1   g09414(.A(new_n9411_), .B(new_n9403_), .Y(new_n9608_));
  AOI21X1  g09415(.A0(new_n9421_), .A1(new_n9412_), .B0(new_n9608_), .Y(new_n9609_));
  XOR2X1   g09416(.A(new_n9609_), .B(new_n9607_), .Y(new_n9610_));
  NAND2X1  g09417(.A(\a[59] ), .B(\a[24] ), .Y(new_n9611_));
  NAND2X1  g09418(.A(\a[60] ), .B(\a[23] ), .Y(new_n9612_));
  AOI22X1  g09419(.A0(new_n9612_), .A1(new_n9611_), .B0(new_n6427_), .B1(new_n1219_), .Y(new_n9613_));
  XOR2X1   g09420(.A(new_n9613_), .B(new_n9440_), .Y(new_n9614_));
  NAND4X1  g09421(.A(\a[53] ), .B(\a[52] ), .C(\a[31] ), .D(\a[30] ), .Y(new_n9615_));
  NAND4X1  g09422(.A(\a[55] ), .B(\a[52] ), .C(\a[31] ), .D(\a[28] ), .Y(new_n9616_));
  AOI22X1  g09423(.A0(new_n9616_), .A1(new_n9615_), .B0(new_n5236_), .B1(new_n2198_), .Y(new_n9617_));
  NAND2X1  g09424(.A(\a[52] ), .B(\a[31] ), .Y(new_n9618_));
  AOI22X1  g09425(.A0(\a[55] ), .A1(\a[28] ), .B0(\a[53] ), .B1(\a[30] ), .Y(new_n9619_));
  AOI21X1  g09426(.A0(new_n5236_), .A1(new_n2198_), .B0(new_n9617_), .Y(new_n9620_));
  INVX1    g09427(.A(new_n9620_), .Y(new_n9621_));
  OAI22X1  g09428(.A0(new_n9621_), .A1(new_n9619_), .B0(new_n9618_), .B1(new_n9617_), .Y(new_n9622_));
  XOR2X1   g09429(.A(new_n9622_), .B(new_n9614_), .Y(new_n9623_));
  INVX1    g09430(.A(new_n9623_), .Y(new_n9624_));
  OR2X1    g09431(.A(new_n9257_), .B(new_n9502_), .Y(new_n9625_));
  AND2X1   g09432(.A(new_n9257_), .B(new_n9502_), .Y(new_n9626_));
  OAI21X1  g09433(.A0(new_n9626_), .A1(new_n9322_), .B0(new_n9625_), .Y(new_n9627_));
  XOR2X1   g09434(.A(new_n9627_), .B(new_n9624_), .Y(new_n9628_));
  NAND2X1  g09435(.A(new_n9499_), .B(new_n9495_), .Y(new_n9629_));
  OAI21X1  g09436(.A0(new_n9504_), .A1(new_n9501_), .B0(new_n9629_), .Y(new_n9630_));
  XOR2X1   g09437(.A(new_n9630_), .B(new_n9628_), .Y(new_n9631_));
  INVX1    g09438(.A(new_n9631_), .Y(new_n9632_));
  XOR2X1   g09439(.A(new_n9632_), .B(new_n9610_), .Y(new_n9633_));
  INVX1    g09440(.A(new_n9633_), .Y(new_n9634_));
  XOR2X1   g09441(.A(new_n9634_), .B(new_n9602_), .Y(new_n9635_));
  XOR2X1   g09442(.A(new_n9635_), .B(new_n9600_), .Y(new_n9636_));
  XOR2X1   g09443(.A(new_n9636_), .B(new_n9581_), .Y(new_n9637_));
  NOR2X1   g09444(.A(new_n9637_), .B(new_n9514_), .Y(new_n9638_));
  AND2X1   g09445(.A(new_n9637_), .B(new_n9514_), .Y(new_n9639_));
  OR2X1    g09446(.A(new_n9639_), .B(new_n9638_), .Y(new_n9640_));
  NOR2X1   g09447(.A(new_n9508_), .B(new_n9386_), .Y(new_n9641_));
  AND2X1   g09448(.A(new_n9508_), .B(new_n9386_), .Y(new_n9642_));
  INVX1    g09449(.A(new_n9642_), .Y(new_n9643_));
  AOI21X1  g09450(.A0(new_n9643_), .A1(new_n9383_), .B0(new_n9641_), .Y(new_n9644_));
  XOR2X1   g09451(.A(new_n9644_), .B(new_n9640_), .Y(\asquared[84] ));
  INVX1    g09452(.A(new_n9638_), .Y(new_n9646_));
  OAI21X1  g09453(.A0(new_n9644_), .A1(new_n9639_), .B0(new_n9646_), .Y(new_n9647_));
  NOR2X1   g09454(.A(new_n9580_), .B(new_n9516_), .Y(new_n9648_));
  INVX1    g09455(.A(new_n9636_), .Y(new_n9649_));
  AOI21X1  g09456(.A0(new_n9649_), .A1(new_n9581_), .B0(new_n9648_), .Y(new_n9650_));
  INVX1    g09457(.A(new_n9600_), .Y(new_n9651_));
  NOR2X1   g09458(.A(new_n9634_), .B(new_n9602_), .Y(new_n9652_));
  AOI21X1  g09459(.A0(new_n9635_), .A1(new_n9651_), .B0(new_n9652_), .Y(new_n9653_));
  INVX1    g09460(.A(new_n9440_), .Y(new_n9654_));
  AOI22X1  g09461(.A0(new_n9613_), .A1(new_n9654_), .B0(new_n6427_), .B1(new_n1219_), .Y(new_n9655_));
  XOR2X1   g09462(.A(new_n9655_), .B(new_n9572_), .Y(new_n9656_));
  AND2X1   g09463(.A(\a[58] ), .B(\a[26] ), .Y(new_n9657_));
  AOI22X1  g09464(.A0(\a[53] ), .A1(\a[31] ), .B0(\a[52] ), .B1(\a[32] ), .Y(new_n9658_));
  INVX1    g09465(.A(new_n9658_), .Y(new_n9659_));
  NAND4X1  g09466(.A(\a[53] ), .B(\a[52] ), .C(\a[32] ), .D(\a[31] ), .Y(new_n9660_));
  NAND3X1  g09467(.A(new_n9659_), .B(new_n9660_), .C(new_n9657_), .Y(new_n9661_));
  AOI22X1  g09468(.A0(new_n9659_), .A1(new_n9657_), .B0(new_n5048_), .B1(new_n2671_), .Y(new_n9662_));
  AOI22X1  g09469(.A0(new_n9662_), .A1(new_n9659_), .B0(new_n9661_), .B1(new_n9657_), .Y(new_n9663_));
  XOR2X1   g09470(.A(new_n9663_), .B(new_n9656_), .Y(new_n9664_));
  INVX1    g09471(.A(new_n9614_), .Y(new_n9665_));
  AND2X1   g09472(.A(new_n9622_), .B(new_n9665_), .Y(new_n9666_));
  AOI21X1  g09473(.A0(new_n9627_), .A1(new_n9624_), .B0(new_n9666_), .Y(new_n9667_));
  XOR2X1   g09474(.A(new_n9667_), .B(new_n9664_), .Y(new_n9668_));
  AND2X1   g09475(.A(new_n9606_), .B(new_n9604_), .Y(new_n9669_));
  OR2X1    g09476(.A(new_n9606_), .B(new_n9604_), .Y(new_n9670_));
  OAI21X1  g09477(.A0(new_n9609_), .A1(new_n9669_), .B0(new_n9670_), .Y(new_n9671_));
  XOR2X1   g09478(.A(new_n9671_), .B(new_n9668_), .Y(new_n9672_));
  NAND2X1  g09479(.A(new_n9630_), .B(new_n9628_), .Y(new_n9673_));
  OAI21X1  g09480(.A0(new_n9632_), .A1(new_n9610_), .B0(new_n9673_), .Y(new_n9674_));
  XOR2X1   g09481(.A(new_n9674_), .B(new_n9672_), .Y(new_n9675_));
  OAI22X1  g09482(.A0(new_n7973_), .A1(new_n1396_), .B0(new_n7972_), .B1(new_n1397_), .Y(new_n9676_));
  OAI21X1  g09483(.A0(new_n6557_), .A1(new_n1395_), .B0(new_n9676_), .Y(new_n9677_));
  AOI21X1  g09484(.A0(new_n6556_), .A1(new_n1394_), .B0(new_n9676_), .Y(new_n9678_));
  OAI22X1  g09485(.A0(new_n6606_), .A1(new_n1086_), .B0(new_n6023_), .B1(new_n1216_), .Y(new_n9679_));
  AND2X1   g09486(.A(\a[63] ), .B(\a[21] ), .Y(new_n9680_));
  AOI22X1  g09487(.A0(new_n9680_), .A1(new_n9677_), .B0(new_n9679_), .B1(new_n9678_), .Y(new_n9681_));
  AND2X1   g09488(.A(\a[51] ), .B(\a[33] ), .Y(new_n9682_));
  INVX1    g09489(.A(new_n9682_), .Y(new_n9683_));
  AOI22X1  g09490(.A0(\a[60] ), .A1(\a[24] ), .B0(\a[59] ), .B1(\a[25] ), .Y(new_n9684_));
  AND2X1   g09491(.A(new_n6427_), .B(new_n1532_), .Y(new_n9685_));
  NOR3X1   g09492(.A(new_n9684_), .B(new_n9685_), .C(new_n9683_), .Y(new_n9686_));
  NOR2X1   g09493(.A(new_n9686_), .B(new_n9685_), .Y(new_n9687_));
  INVX1    g09494(.A(new_n9687_), .Y(new_n9688_));
  OAI22X1  g09495(.A0(new_n9688_), .A1(new_n9684_), .B0(new_n9686_), .B1(new_n9683_), .Y(new_n9689_));
  XOR2X1   g09496(.A(new_n9689_), .B(new_n9681_), .Y(new_n9690_));
  OAI22X1  g09497(.A0(new_n7652_), .A1(new_n4915_), .B0(new_n8802_), .B1(new_n5418_), .Y(new_n9691_));
  OAI21X1  g09498(.A0(new_n4280_), .A1(new_n5417_), .B0(new_n9691_), .Y(new_n9692_));
  AND2X1   g09499(.A(\a[50] ), .B(\a[34] ), .Y(new_n9693_));
  AOI21X1  g09500(.A0(new_n4274_), .A1(new_n2682_), .B0(new_n9691_), .Y(new_n9694_));
  OAI22X1  g09501(.A0(new_n3915_), .A1(new_n2557_), .B0(new_n3926_), .B1(new_n2583_), .Y(new_n9695_));
  AOI22X1  g09502(.A0(new_n9695_), .A1(new_n9694_), .B0(new_n9693_), .B1(new_n9692_), .Y(new_n9696_));
  XOR2X1   g09503(.A(new_n9696_), .B(new_n9690_), .Y(new_n9697_));
  AOI22X1  g09504(.A0(\a[55] ), .A1(\a[29] ), .B0(\a[46] ), .B1(\a[38] ), .Y(new_n9698_));
  NOR4X1   g09505(.A(new_n4906_), .B(new_n3460_), .C(new_n2519_), .D(new_n1803_), .Y(new_n9699_));
  AND2X1   g09506(.A(\a[46] ), .B(\a[28] ), .Y(new_n9700_));
  AND2X1   g09507(.A(\a[56] ), .B(\a[38] ), .Y(new_n9701_));
  AOI22X1  g09508(.A0(new_n9701_), .A1(new_n9700_), .B0(new_n6237_), .B1(new_n1674_), .Y(new_n9702_));
  NOR2X1   g09509(.A(new_n9702_), .B(new_n9699_), .Y(new_n9703_));
  INVX1    g09510(.A(new_n9699_), .Y(new_n9704_));
  AND2X1   g09511(.A(new_n9702_), .B(new_n9704_), .Y(new_n9705_));
  INVX1    g09512(.A(new_n9705_), .Y(new_n9706_));
  NAND2X1  g09513(.A(\a[56] ), .B(\a[28] ), .Y(new_n9707_));
  OAI22X1  g09514(.A0(new_n9707_), .A1(new_n9703_), .B0(new_n9706_), .B1(new_n9698_), .Y(new_n9708_));
  NAND4X1  g09515(.A(\a[45] ), .B(\a[43] ), .C(\a[41] ), .D(\a[39] ), .Y(new_n9709_));
  NAND4X1  g09516(.A(\a[45] ), .B(\a[44] ), .C(\a[40] ), .D(\a[39] ), .Y(new_n9710_));
  AOI22X1  g09517(.A0(new_n9710_), .A1(new_n9709_), .B0(new_n4404_), .B1(new_n4992_), .Y(new_n9711_));
  NAND2X1  g09518(.A(\a[45] ), .B(\a[39] ), .Y(new_n9712_));
  NAND4X1  g09519(.A(\a[44] ), .B(\a[43] ), .C(\a[41] ), .D(\a[40] ), .Y(new_n9713_));
  NAND3X1  g09520(.A(new_n9710_), .B(new_n9709_), .C(new_n9713_), .Y(new_n9714_));
  AOI22X1  g09521(.A0(\a[44] ), .A1(\a[40] ), .B0(\a[43] ), .B1(\a[41] ), .Y(new_n9715_));
  OAI22X1  g09522(.A0(new_n9715_), .A1(new_n9714_), .B0(new_n9712_), .B1(new_n9711_), .Y(new_n9716_));
  XOR2X1   g09523(.A(new_n9716_), .B(new_n9708_), .Y(new_n9717_));
  AND2X1   g09524(.A(\a[47] ), .B(\a[37] ), .Y(new_n9718_));
  INVX1    g09525(.A(new_n9718_), .Y(new_n9719_));
  AOI22X1  g09526(.A0(\a[57] ), .A1(\a[27] ), .B0(\a[54] ), .B1(\a[30] ), .Y(new_n9720_));
  NOR4X1   g09527(.A(new_n5441_), .B(new_n4835_), .C(new_n1684_), .D(new_n1679_), .Y(new_n9721_));
  NOR3X1   g09528(.A(new_n9720_), .B(new_n9721_), .C(new_n9719_), .Y(new_n9722_));
  INVX1    g09529(.A(new_n9720_), .Y(new_n9723_));
  AOI21X1  g09530(.A0(new_n9723_), .A1(new_n9718_), .B0(new_n9721_), .Y(new_n9724_));
  INVX1    g09531(.A(new_n9724_), .Y(new_n9725_));
  OAI22X1  g09532(.A0(new_n9725_), .A1(new_n9720_), .B0(new_n9722_), .B1(new_n9719_), .Y(new_n9726_));
  INVX1    g09533(.A(new_n9726_), .Y(new_n9727_));
  XOR2X1   g09534(.A(new_n9727_), .B(new_n9717_), .Y(new_n9728_));
  XOR2X1   g09535(.A(new_n9728_), .B(new_n9697_), .Y(new_n9729_));
  INVX1    g09536(.A(new_n9540_), .Y(new_n9730_));
  XOR2X1   g09537(.A(new_n9563_), .B(new_n9730_), .Y(new_n9731_));
  XOR2X1   g09538(.A(new_n9731_), .B(new_n9555_), .Y(new_n9732_));
  INVX1    g09539(.A(new_n9732_), .Y(new_n9733_));
  NOR2X1   g09540(.A(new_n9447_), .B(new_n9418_), .Y(new_n9734_));
  AOI21X1  g09541(.A0(new_n9589_), .A1(new_n9434_), .B0(new_n9734_), .Y(new_n9735_));
  AND2X1   g09542(.A(new_n9409_), .B(new_n9400_), .Y(new_n9736_));
  AOI21X1  g09543(.A0(new_n9592_), .A1(new_n9467_), .B0(new_n9736_), .Y(new_n9737_));
  XOR2X1   g09544(.A(new_n9737_), .B(new_n9735_), .Y(new_n9738_));
  XOR2X1   g09545(.A(new_n9738_), .B(new_n9733_), .Y(new_n9739_));
  XOR2X1   g09546(.A(new_n9739_), .B(new_n9729_), .Y(new_n9740_));
  XOR2X1   g09547(.A(new_n9740_), .B(new_n9675_), .Y(new_n9741_));
  XOR2X1   g09548(.A(new_n9741_), .B(new_n9653_), .Y(new_n9742_));
  NAND2X1  g09549(.A(new_n9577_), .B(new_n9523_), .Y(new_n9743_));
  NOR2X1   g09550(.A(new_n9577_), .B(new_n9523_), .Y(new_n9744_));
  OAI21X1  g09551(.A0(new_n9744_), .A1(new_n9518_), .B0(new_n9743_), .Y(new_n9745_));
  OR2X1    g09552(.A(new_n9587_), .B(new_n9584_), .Y(new_n9746_));
  INVX1    g09553(.A(new_n9599_), .Y(new_n9747_));
  OAI21X1  g09554(.A0(new_n9747_), .A1(new_n9588_), .B0(new_n9746_), .Y(new_n9748_));
  XOR2X1   g09555(.A(new_n9748_), .B(new_n9745_), .Y(new_n9749_));
  NAND2X1  g09556(.A(new_n9547_), .B(new_n9543_), .Y(new_n9750_));
  OAI21X1  g09557(.A0(new_n9576_), .A1(new_n9548_), .B0(new_n9750_), .Y(new_n9751_));
  INVX1    g09558(.A(new_n9593_), .Y(new_n9752_));
  OR2X1    g09559(.A(new_n9597_), .B(new_n9752_), .Y(new_n9753_));
  OAI21X1  g09560(.A0(new_n9598_), .A1(new_n9591_), .B0(new_n9753_), .Y(new_n9754_));
  XOR2X1   g09561(.A(new_n9754_), .B(new_n9751_), .Y(new_n9755_));
  XOR2X1   g09562(.A(new_n9534_), .B(new_n9525_), .Y(new_n9756_));
  XOR2X1   g09563(.A(new_n9756_), .B(new_n9620_), .Y(new_n9757_));
  AND2X1   g09564(.A(new_n9565_), .B(new_n9557_), .Y(new_n9758_));
  AND2X1   g09565(.A(new_n9574_), .B(new_n9566_), .Y(new_n9759_));
  OR2X1    g09566(.A(new_n9759_), .B(new_n9758_), .Y(new_n9760_));
  INVX1    g09567(.A(new_n9535_), .Y(new_n9761_));
  OR2X1    g09568(.A(new_n9542_), .B(new_n9536_), .Y(new_n9762_));
  OAI21X1  g09569(.A0(new_n9761_), .A1(new_n9528_), .B0(new_n9762_), .Y(new_n9763_));
  XOR2X1   g09570(.A(new_n9763_), .B(new_n9760_), .Y(new_n9764_));
  XOR2X1   g09571(.A(new_n9764_), .B(new_n9757_), .Y(new_n9765_));
  XOR2X1   g09572(.A(new_n9765_), .B(new_n9755_), .Y(new_n9766_));
  XOR2X1   g09573(.A(new_n9766_), .B(new_n9749_), .Y(new_n9767_));
  XOR2X1   g09574(.A(new_n9767_), .B(new_n9742_), .Y(new_n9768_));
  XOR2X1   g09575(.A(new_n9768_), .B(new_n9650_), .Y(new_n9769_));
  XOR2X1   g09576(.A(new_n9769_), .B(new_n9647_), .Y(\asquared[85] ));
  NOR2X1   g09577(.A(new_n9768_), .B(new_n9650_), .Y(new_n9771_));
  AND2X1   g09578(.A(new_n9768_), .B(new_n9650_), .Y(new_n9772_));
  INVX1    g09579(.A(new_n9772_), .Y(new_n9773_));
  AOI21X1  g09580(.A0(new_n9773_), .A1(new_n9647_), .B0(new_n9771_), .Y(new_n9774_));
  INVX1    g09581(.A(new_n9653_), .Y(new_n9775_));
  AND2X1   g09582(.A(new_n9741_), .B(new_n9775_), .Y(new_n9776_));
  INVX1    g09583(.A(new_n9742_), .Y(new_n9777_));
  AOI21X1  g09584(.A0(new_n9767_), .A1(new_n9777_), .B0(new_n9776_), .Y(new_n9778_));
  AND2X1   g09585(.A(new_n9748_), .B(new_n9745_), .Y(new_n9779_));
  AOI21X1  g09586(.A0(new_n9766_), .A1(new_n9749_), .B0(new_n9779_), .Y(new_n9780_));
  AOI22X1  g09587(.A0(\a[63] ), .A1(\a[22] ), .B0(\a[57] ), .B1(\a[28] ), .Y(new_n9781_));
  AND2X1   g09588(.A(\a[50] ), .B(\a[35] ), .Y(new_n9782_));
  INVX1    g09589(.A(new_n9782_), .Y(new_n9783_));
  NOR4X1   g09590(.A(new_n6549_), .B(new_n5441_), .C(new_n1431_), .D(new_n1086_), .Y(new_n9784_));
  NOR3X1   g09591(.A(new_n9783_), .B(new_n9784_), .C(new_n9781_), .Y(new_n9785_));
  INVX1    g09592(.A(new_n9781_), .Y(new_n9786_));
  AOI21X1  g09593(.A0(new_n9782_), .A1(new_n9786_), .B0(new_n9784_), .Y(new_n9787_));
  INVX1    g09594(.A(new_n9787_), .Y(new_n9788_));
  OAI22X1  g09595(.A0(new_n9788_), .A1(new_n9781_), .B0(new_n9785_), .B1(new_n9783_), .Y(new_n9789_));
  OAI22X1  g09596(.A0(new_n7336_), .A1(new_n2675_), .B0(new_n8145_), .B1(new_n2920_), .Y(new_n9790_));
  OAI21X1  g09597(.A0(new_n7793_), .A1(new_n2919_), .B0(new_n9790_), .Y(new_n9791_));
  AND2X1   g09598(.A(\a[53] ), .B(\a[32] ), .Y(new_n9792_));
  AOI21X1  g09599(.A0(new_n7164_), .A1(new_n2918_), .B0(new_n9790_), .Y(new_n9793_));
  OAI22X1  g09600(.A0(new_n4354_), .A1(new_n1851_), .B0(new_n4349_), .B1(new_n2028_), .Y(new_n9794_));
  AOI22X1  g09601(.A0(new_n9794_), .A1(new_n9793_), .B0(new_n9792_), .B1(new_n9791_), .Y(new_n9795_));
  XOR2X1   g09602(.A(new_n9795_), .B(new_n9789_), .Y(new_n9796_));
  OAI22X1  g09603(.A0(new_n8874_), .A1(new_n7617_), .B0(new_n8873_), .B1(new_n6180_), .Y(new_n9797_));
  OAI21X1  g09604(.A0(new_n7642_), .A1(new_n7618_), .B0(new_n9797_), .Y(new_n9798_));
  AND2X1   g09605(.A(\a[46] ), .B(\a[39] ), .Y(new_n9799_));
  AOI21X1  g09606(.A0(new_n3918_), .A1(new_n4404_), .B0(new_n9797_), .Y(new_n9800_));
  OAI22X1  g09607(.A0(new_n3811_), .A1(new_n3036_), .B0(new_n5268_), .B1(new_n3081_), .Y(new_n9801_));
  AOI22X1  g09608(.A0(new_n9801_), .A1(new_n9800_), .B0(new_n9799_), .B1(new_n9798_), .Y(new_n9802_));
  XOR2X1   g09609(.A(new_n9802_), .B(new_n9796_), .Y(new_n9803_));
  NAND3X1  g09610(.A(\a[62] ), .B(\a[43] ), .C(\a[23] ), .Y(new_n9804_));
  AND2X1   g09611(.A(new_n9804_), .B(new_n3462_), .Y(new_n9805_));
  AND2X1   g09612(.A(new_n9804_), .B(new_n6502_), .Y(new_n9806_));
  INVX1    g09613(.A(new_n9806_), .Y(new_n9807_));
  AOI21X1  g09614(.A0(\a[62] ), .A1(\a[23] ), .B0(\a[43] ), .Y(new_n9808_));
  OAI22X1  g09615(.A0(new_n9808_), .A1(new_n9807_), .B0(new_n9805_), .B1(new_n6502_), .Y(new_n9809_));
  INVX1    g09616(.A(new_n9809_), .Y(new_n9810_));
  NAND4X1  g09617(.A(\a[49] ), .B(\a[47] ), .C(\a[38] ), .D(\a[36] ), .Y(new_n9811_));
  NAND4X1  g09618(.A(\a[49] ), .B(\a[48] ), .C(\a[37] ), .D(\a[36] ), .Y(new_n9812_));
  AOI22X1  g09619(.A0(new_n9812_), .A1(new_n9811_), .B0(new_n4272_), .B1(new_n3164_), .Y(new_n9813_));
  NAND2X1  g09620(.A(\a[49] ), .B(\a[36] ), .Y(new_n9814_));
  AOI22X1  g09621(.A0(\a[48] ), .A1(\a[37] ), .B0(\a[47] ), .B1(\a[38] ), .Y(new_n9815_));
  AOI21X1  g09622(.A0(new_n4272_), .A1(new_n3164_), .B0(new_n9813_), .Y(new_n9816_));
  INVX1    g09623(.A(new_n9816_), .Y(new_n9817_));
  OAI22X1  g09624(.A0(new_n9817_), .A1(new_n9815_), .B0(new_n9814_), .B1(new_n9813_), .Y(new_n9818_));
  XOR2X1   g09625(.A(new_n9818_), .B(new_n9810_), .Y(new_n9819_));
  OAI22X1  g09626(.A0(new_n8560_), .A1(new_n2197_), .B0(new_n8559_), .B1(new_n2430_), .Y(new_n9820_));
  OAI21X1  g09627(.A0(new_n5241_), .A1(new_n2076_), .B0(new_n9820_), .Y(new_n9821_));
  AND2X1   g09628(.A(\a[56] ), .B(\a[29] ), .Y(new_n9822_));
  AOI21X1  g09629(.A0(new_n5240_), .A1(new_n2075_), .B0(new_n9820_), .Y(new_n9823_));
  OAI22X1  g09630(.A0(new_n4906_), .A1(new_n1684_), .B0(new_n4835_), .B1(new_n1704_), .Y(new_n9824_));
  AOI22X1  g09631(.A0(new_n9824_), .A1(new_n9823_), .B0(new_n9822_), .B1(new_n9821_), .Y(new_n9825_));
  XOR2X1   g09632(.A(new_n9825_), .B(new_n9819_), .Y(new_n9826_));
  XOR2X1   g09633(.A(new_n9826_), .B(new_n9803_), .Y(new_n9827_));
  AND2X1   g09634(.A(new_n9763_), .B(new_n9760_), .Y(new_n9828_));
  AND2X1   g09635(.A(new_n9764_), .B(new_n9757_), .Y(new_n9829_));
  OR2X1    g09636(.A(new_n9829_), .B(new_n9828_), .Y(new_n9830_));
  XOR2X1   g09637(.A(new_n9830_), .B(new_n9827_), .Y(new_n9831_));
  NOR2X1   g09638(.A(new_n9737_), .B(new_n9735_), .Y(new_n9832_));
  AOI21X1  g09639(.A0(new_n9738_), .A1(new_n9732_), .B0(new_n9832_), .Y(new_n9833_));
  NAND2X1  g09640(.A(\a[61] ), .B(\a[24] ), .Y(new_n9834_));
  XOR2X1   g09641(.A(new_n9834_), .B(new_n9714_), .Y(new_n9835_));
  XOR2X1   g09642(.A(new_n9835_), .B(new_n9705_), .Y(new_n9836_));
  XOR2X1   g09643(.A(new_n9724_), .B(new_n9662_), .Y(new_n9837_));
  NAND4X1  g09644(.A(\a[60] ), .B(\a[58] ), .C(\a[27] ), .D(\a[25] ), .Y(new_n9838_));
  NAND4X1  g09645(.A(\a[60] ), .B(\a[59] ), .C(\a[26] ), .D(\a[25] ), .Y(new_n9839_));
  AOI22X1  g09646(.A0(new_n9839_), .A1(new_n9838_), .B0(new_n6121_), .B1(new_n1995_), .Y(new_n9840_));
  NAND2X1  g09647(.A(\a[60] ), .B(\a[25] ), .Y(new_n9841_));
  NAND4X1  g09648(.A(\a[59] ), .B(\a[58] ), .C(\a[27] ), .D(\a[26] ), .Y(new_n9842_));
  NAND3X1  g09649(.A(new_n9839_), .B(new_n9838_), .C(new_n9842_), .Y(new_n9843_));
  AOI22X1  g09650(.A0(\a[59] ), .A1(\a[26] ), .B0(\a[58] ), .B1(\a[27] ), .Y(new_n9844_));
  OAI22X1  g09651(.A0(new_n9844_), .A1(new_n9843_), .B0(new_n9841_), .B1(new_n9840_), .Y(new_n9845_));
  XOR2X1   g09652(.A(new_n9845_), .B(new_n9837_), .Y(new_n9846_));
  NOR2X1   g09653(.A(new_n9846_), .B(new_n9836_), .Y(new_n9847_));
  XOR2X1   g09654(.A(new_n9846_), .B(new_n9836_), .Y(new_n9848_));
  NAND2X1  g09655(.A(new_n9846_), .B(new_n9836_), .Y(new_n9849_));
  OAI21X1  g09656(.A0(new_n9847_), .A1(new_n9833_), .B0(new_n9849_), .Y(new_n9850_));
  OAI22X1  g09657(.A0(new_n9850_), .A1(new_n9847_), .B0(new_n9848_), .B1(new_n9833_), .Y(new_n9851_));
  XOR2X1   g09658(.A(new_n9694_), .B(new_n9678_), .Y(new_n9852_));
  XOR2X1   g09659(.A(new_n9852_), .B(new_n9688_), .Y(new_n9853_));
  AND2X1   g09660(.A(new_n9716_), .B(new_n9708_), .Y(new_n9854_));
  AND2X1   g09661(.A(new_n9726_), .B(new_n9717_), .Y(new_n9855_));
  OR2X1    g09662(.A(new_n9855_), .B(new_n9854_), .Y(new_n9856_));
  INVX1    g09663(.A(new_n9689_), .Y(new_n9857_));
  OR2X1    g09664(.A(new_n9857_), .B(new_n9681_), .Y(new_n9858_));
  OAI21X1  g09665(.A0(new_n9696_), .A1(new_n9690_), .B0(new_n9858_), .Y(new_n9859_));
  XOR2X1   g09666(.A(new_n9859_), .B(new_n9856_), .Y(new_n9860_));
  XOR2X1   g09667(.A(new_n9860_), .B(new_n9853_), .Y(new_n9861_));
  XOR2X1   g09668(.A(new_n9861_), .B(new_n9851_), .Y(new_n9862_));
  XOR2X1   g09669(.A(new_n9862_), .B(new_n9831_), .Y(new_n9863_));
  XOR2X1   g09670(.A(new_n9863_), .B(new_n9780_), .Y(new_n9864_));
  AND2X1   g09671(.A(new_n9754_), .B(new_n9751_), .Y(new_n9865_));
  AOI21X1  g09672(.A0(new_n9765_), .A1(new_n9755_), .B0(new_n9865_), .Y(new_n9866_));
  INVX1    g09673(.A(new_n9866_), .Y(new_n9867_));
  AND2X1   g09674(.A(new_n9563_), .B(new_n9730_), .Y(new_n9868_));
  AOI21X1  g09675(.A0(new_n9731_), .A1(new_n9555_), .B0(new_n9868_), .Y(new_n9869_));
  INVX1    g09676(.A(new_n9525_), .Y(new_n9870_));
  NOR2X1   g09677(.A(new_n9756_), .B(new_n9620_), .Y(new_n9871_));
  AOI21X1  g09678(.A0(new_n9534_), .A1(new_n9870_), .B0(new_n9871_), .Y(new_n9872_));
  XOR2X1   g09679(.A(new_n9872_), .B(new_n9869_), .Y(new_n9873_));
  NOR2X1   g09680(.A(new_n9655_), .B(new_n9572_), .Y(new_n9874_));
  INVX1    g09681(.A(new_n9874_), .Y(new_n9875_));
  INVX1    g09682(.A(new_n9656_), .Y(new_n9876_));
  OAI21X1  g09683(.A0(new_n9663_), .A1(new_n9876_), .B0(new_n9875_), .Y(new_n9877_));
  INVX1    g09684(.A(new_n9877_), .Y(new_n9878_));
  XOR2X1   g09685(.A(new_n9878_), .B(new_n9873_), .Y(new_n9879_));
  NOR2X1   g09686(.A(new_n9667_), .B(new_n9664_), .Y(new_n9880_));
  AOI21X1  g09687(.A0(new_n9671_), .A1(new_n9668_), .B0(new_n9880_), .Y(new_n9881_));
  XOR2X1   g09688(.A(new_n9881_), .B(new_n9879_), .Y(new_n9882_));
  XOR2X1   g09689(.A(new_n9726_), .B(new_n9717_), .Y(new_n9883_));
  NAND2X1  g09690(.A(new_n9883_), .B(new_n9697_), .Y(new_n9884_));
  OAI21X1  g09691(.A0(new_n9739_), .A1(new_n9729_), .B0(new_n9884_), .Y(new_n9885_));
  XOR2X1   g09692(.A(new_n9885_), .B(new_n9882_), .Y(new_n9886_));
  XOR2X1   g09693(.A(new_n9886_), .B(new_n9867_), .Y(new_n9887_));
  INVX1    g09694(.A(new_n9887_), .Y(new_n9888_));
  AND2X1   g09695(.A(new_n9674_), .B(new_n9672_), .Y(new_n9889_));
  AOI21X1  g09696(.A0(new_n9740_), .A1(new_n9675_), .B0(new_n9889_), .Y(new_n9890_));
  XOR2X1   g09697(.A(new_n9890_), .B(new_n9888_), .Y(new_n9891_));
  XOR2X1   g09698(.A(new_n9891_), .B(new_n9864_), .Y(new_n9892_));
  NOR2X1   g09699(.A(new_n9892_), .B(new_n9778_), .Y(new_n9893_));
  AND2X1   g09700(.A(new_n9892_), .B(new_n9778_), .Y(new_n9894_));
  OR2X1    g09701(.A(new_n9894_), .B(new_n9893_), .Y(new_n9895_));
  XOR2X1   g09702(.A(new_n9895_), .B(new_n9774_), .Y(\asquared[86] ));
  INVX1    g09703(.A(new_n9863_), .Y(new_n9897_));
  OR2X1    g09704(.A(new_n9897_), .B(new_n9780_), .Y(new_n9898_));
  INVX1    g09705(.A(new_n9891_), .Y(new_n9899_));
  OAI21X1  g09706(.A0(new_n9899_), .A1(new_n9864_), .B0(new_n9898_), .Y(new_n9900_));
  NAND2X1  g09707(.A(new_n9845_), .B(new_n9837_), .Y(new_n9901_));
  OAI21X1  g09708(.A0(new_n9724_), .A1(new_n9662_), .B0(new_n9901_), .Y(new_n9902_));
  INVX1    g09709(.A(new_n9789_), .Y(new_n9903_));
  OR2X1    g09710(.A(new_n9795_), .B(new_n9903_), .Y(new_n9904_));
  OAI21X1  g09711(.A0(new_n9802_), .A1(new_n9796_), .B0(new_n9904_), .Y(new_n9905_));
  XOR2X1   g09712(.A(new_n9905_), .B(new_n9902_), .Y(new_n9906_));
  NAND2X1  g09713(.A(new_n9818_), .B(new_n9809_), .Y(new_n9907_));
  OAI21X1  g09714(.A0(new_n9825_), .A1(new_n9819_), .B0(new_n9907_), .Y(new_n9908_));
  XOR2X1   g09715(.A(new_n9908_), .B(new_n9906_), .Y(new_n9909_));
  NAND2X1  g09716(.A(new_n9877_), .B(new_n9873_), .Y(new_n9910_));
  OAI21X1  g09717(.A0(new_n9872_), .A1(new_n9869_), .B0(new_n9910_), .Y(new_n9911_));
  XOR2X1   g09718(.A(new_n9823_), .B(new_n9800_), .Y(new_n9912_));
  XOR2X1   g09719(.A(new_n9912_), .B(new_n9816_), .Y(new_n9913_));
  INVX1    g09720(.A(new_n9793_), .Y(new_n9914_));
  XOR2X1   g09721(.A(new_n9843_), .B(new_n9914_), .Y(new_n9915_));
  XOR2X1   g09722(.A(new_n9915_), .B(new_n9787_), .Y(new_n9916_));
  XOR2X1   g09723(.A(new_n9916_), .B(new_n9913_), .Y(new_n9917_));
  XOR2X1   g09724(.A(new_n9917_), .B(new_n9911_), .Y(new_n9918_));
  XOR2X1   g09725(.A(new_n9918_), .B(new_n9909_), .Y(new_n9919_));
  AND2X1   g09726(.A(new_n9859_), .B(new_n9856_), .Y(new_n9920_));
  AOI21X1  g09727(.A0(new_n9860_), .A1(new_n9853_), .B0(new_n9920_), .Y(new_n9921_));
  AOI22X1  g09728(.A0(\a[50] ), .A1(\a[36] ), .B0(\a[49] ), .B1(\a[37] ), .Y(new_n9922_));
  AND2X1   g09729(.A(\a[63] ), .B(\a[23] ), .Y(new_n9923_));
  INVX1    g09730(.A(new_n9923_), .Y(new_n9924_));
  AND2X1   g09731(.A(new_n4321_), .B(new_n3330_), .Y(new_n9925_));
  NOR3X1   g09732(.A(new_n9924_), .B(new_n9925_), .C(new_n9922_), .Y(new_n9926_));
  NOR2X1   g09733(.A(new_n9926_), .B(new_n9925_), .Y(new_n9927_));
  INVX1    g09734(.A(new_n9927_), .Y(new_n9928_));
  OAI22X1  g09735(.A0(new_n9928_), .A1(new_n9922_), .B0(new_n9926_), .B1(new_n9924_), .Y(new_n9929_));
  OAI22X1  g09736(.A0(new_n7336_), .A1(new_n2919_), .B0(new_n8145_), .B1(new_n4914_), .Y(new_n9930_));
  OAI21X1  g09737(.A0(new_n7793_), .A1(new_n4915_), .B0(new_n9930_), .Y(new_n9931_));
  AND2X1   g09738(.A(\a[53] ), .B(\a[33] ), .Y(new_n9932_));
  AOI21X1  g09739(.A0(new_n7164_), .A1(new_n2361_), .B0(new_n9930_), .Y(new_n9933_));
  OAI22X1  g09740(.A0(new_n4354_), .A1(new_n2028_), .B0(new_n4349_), .B1(new_n2557_), .Y(new_n9934_));
  AOI22X1  g09741(.A0(new_n9934_), .A1(new_n9933_), .B0(new_n9932_), .B1(new_n9931_), .Y(new_n9935_));
  XOR2X1   g09742(.A(new_n9935_), .B(new_n9929_), .Y(new_n9936_));
  AOI22X1  g09743(.A0(\a[57] ), .A1(\a[29] ), .B0(\a[55] ), .B1(\a[31] ), .Y(new_n9937_));
  INVX1    g09744(.A(new_n9937_), .Y(new_n9938_));
  NAND4X1  g09745(.A(\a[57] ), .B(\a[55] ), .C(\a[31] ), .D(\a[29] ), .Y(new_n9939_));
  NAND3X1  g09746(.A(new_n9938_), .B(new_n9939_), .C(new_n4713_), .Y(new_n9940_));
  AOI22X1  g09747(.A0(new_n9938_), .A1(new_n4713_), .B0(new_n9461_), .B1(new_n2429_), .Y(new_n9941_));
  AOI22X1  g09748(.A0(new_n9941_), .A1(new_n9938_), .B0(new_n9940_), .B1(new_n4713_), .Y(new_n9942_));
  XOR2X1   g09749(.A(new_n9942_), .B(new_n9936_), .Y(new_n9943_));
  INVX1    g09750(.A(new_n9943_), .Y(new_n9944_));
  NAND4X1  g09751(.A(\a[60] ), .B(\a[58] ), .C(\a[28] ), .D(\a[26] ), .Y(new_n9945_));
  NAND4X1  g09752(.A(\a[60] ), .B(\a[59] ), .C(\a[27] ), .D(\a[26] ), .Y(new_n9946_));
  AOI22X1  g09753(.A0(new_n9946_), .A1(new_n9945_), .B0(new_n6121_), .B1(new_n1671_), .Y(new_n9947_));
  NAND4X1  g09754(.A(\a[59] ), .B(\a[58] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n9948_));
  NAND3X1  g09755(.A(new_n9946_), .B(new_n9945_), .C(new_n9948_), .Y(new_n9949_));
  AOI22X1  g09756(.A0(\a[59] ), .A1(\a[27] ), .B0(\a[58] ), .B1(\a[28] ), .Y(new_n9950_));
  NAND2X1  g09757(.A(\a[60] ), .B(\a[26] ), .Y(new_n9951_));
  OAI22X1  g09758(.A0(new_n9951_), .A1(new_n9947_), .B0(new_n9950_), .B1(new_n9949_), .Y(new_n9952_));
  NAND2X1  g09759(.A(\a[45] ), .B(\a[41] ), .Y(new_n9953_));
  AND2X1   g09760(.A(\a[54] ), .B(\a[32] ), .Y(new_n9954_));
  NAND4X1  g09761(.A(\a[54] ), .B(\a[45] ), .C(\a[41] ), .D(\a[32] ), .Y(new_n9955_));
  NAND4X1  g09762(.A(\a[45] ), .B(\a[44] ), .C(\a[42] ), .D(\a[41] ), .Y(new_n9956_));
  AOI22X1  g09763(.A0(new_n9956_), .A1(new_n9955_), .B0(new_n9954_), .B1(new_n3208_), .Y(new_n9957_));
  NAND4X1  g09764(.A(\a[54] ), .B(\a[44] ), .C(\a[42] ), .D(\a[32] ), .Y(new_n9958_));
  NAND3X1  g09765(.A(new_n9956_), .B(new_n9955_), .C(new_n9958_), .Y(new_n9959_));
  AOI22X1  g09766(.A0(\a[54] ), .A1(\a[32] ), .B0(\a[44] ), .B1(\a[42] ), .Y(new_n9960_));
  OAI22X1  g09767(.A0(new_n9960_), .A1(new_n9959_), .B0(new_n9957_), .B1(new_n9953_), .Y(new_n9961_));
  XOR2X1   g09768(.A(new_n9961_), .B(new_n9952_), .Y(new_n9962_));
  AND2X1   g09769(.A(\a[56] ), .B(\a[30] ), .Y(new_n9963_));
  INVX1    g09770(.A(new_n9963_), .Y(new_n9964_));
  AOI22X1  g09771(.A0(\a[47] ), .A1(\a[39] ), .B0(\a[46] ), .B1(\a[40] ), .Y(new_n9965_));
  AND2X1   g09772(.A(new_n3893_), .B(new_n4077_), .Y(new_n9966_));
  NOR3X1   g09773(.A(new_n9965_), .B(new_n9966_), .C(new_n9964_), .Y(new_n9967_));
  NOR2X1   g09774(.A(new_n9967_), .B(new_n9966_), .Y(new_n9968_));
  INVX1    g09775(.A(new_n9968_), .Y(new_n9969_));
  OAI22X1  g09776(.A0(new_n9969_), .A1(new_n9965_), .B0(new_n9967_), .B1(new_n9964_), .Y(new_n9970_));
  XOR2X1   g09777(.A(new_n9970_), .B(new_n9962_), .Y(new_n9971_));
  XOR2X1   g09778(.A(new_n9971_), .B(new_n9944_), .Y(new_n9972_));
  XOR2X1   g09779(.A(new_n9972_), .B(new_n9921_), .Y(new_n9973_));
  XOR2X1   g09780(.A(new_n9973_), .B(new_n9919_), .Y(new_n9974_));
  AND2X1   g09781(.A(new_n9886_), .B(new_n9867_), .Y(new_n9975_));
  INVX1    g09782(.A(new_n9975_), .Y(new_n9976_));
  OAI21X1  g09783(.A0(new_n9890_), .A1(new_n9888_), .B0(new_n9976_), .Y(new_n9977_));
  AND2X1   g09784(.A(new_n9974_), .B(new_n9977_), .Y(new_n9978_));
  INVX1    g09785(.A(new_n9978_), .Y(new_n9979_));
  NAND2X1  g09786(.A(new_n9979_), .B(new_n9974_), .Y(new_n9980_));
  XOR2X1   g09787(.A(new_n9974_), .B(new_n9977_), .Y(new_n9981_));
  AND2X1   g09788(.A(new_n9861_), .B(new_n9851_), .Y(new_n9982_));
  AOI21X1  g09789(.A0(new_n9862_), .A1(new_n9831_), .B0(new_n9982_), .Y(new_n9983_));
  NOR2X1   g09790(.A(new_n9881_), .B(new_n9879_), .Y(new_n9984_));
  AOI21X1  g09791(.A0(new_n9885_), .A1(new_n9882_), .B0(new_n9984_), .Y(new_n9985_));
  XOR2X1   g09792(.A(new_n9985_), .B(new_n9983_), .Y(new_n9986_));
  AND2X1   g09793(.A(\a[61] ), .B(\a[25] ), .Y(new_n9987_));
  AND2X1   g09794(.A(\a[62] ), .B(\a[24] ), .Y(new_n9988_));
  OAI22X1  g09795(.A0(new_n9988_), .A1(new_n9987_), .B0(new_n6557_), .B1(new_n1772_), .Y(new_n9989_));
  XOR2X1   g09796(.A(new_n9989_), .B(new_n9807_), .Y(new_n9990_));
  INVX1    g09797(.A(new_n9990_), .Y(new_n9991_));
  NAND3X1  g09798(.A(new_n9714_), .B(\a[61] ), .C(\a[24] ), .Y(new_n9992_));
  OAI21X1  g09799(.A0(new_n9835_), .A1(new_n9705_), .B0(new_n9992_), .Y(new_n9993_));
  XOR2X1   g09800(.A(new_n9993_), .B(new_n9991_), .Y(new_n9994_));
  INVX1    g09801(.A(new_n9994_), .Y(new_n9995_));
  NOR2X1   g09802(.A(new_n9694_), .B(new_n9678_), .Y(new_n9996_));
  AOI21X1  g09803(.A0(new_n9852_), .A1(new_n9688_), .B0(new_n9996_), .Y(new_n9997_));
  XOR2X1   g09804(.A(new_n9997_), .B(new_n9995_), .Y(new_n9998_));
  INVX1    g09805(.A(new_n9998_), .Y(new_n9999_));
  XOR2X1   g09806(.A(new_n9999_), .B(new_n9850_), .Y(new_n10000_));
  AND2X1   g09807(.A(new_n9826_), .B(new_n9803_), .Y(new_n10001_));
  AOI21X1  g09808(.A0(new_n9830_), .A1(new_n9827_), .B0(new_n10001_), .Y(new_n10002_));
  XOR2X1   g09809(.A(new_n10002_), .B(new_n10000_), .Y(new_n10003_));
  XOR2X1   g09810(.A(new_n10003_), .B(new_n9986_), .Y(new_n10004_));
  AND2X1   g09811(.A(new_n10004_), .B(new_n9981_), .Y(new_n10005_));
  AOI21X1  g09812(.A0(new_n9979_), .A1(new_n9977_), .B0(new_n10004_), .Y(new_n10006_));
  AOI21X1  g09813(.A0(new_n10006_), .A1(new_n9980_), .B0(new_n10005_), .Y(new_n10007_));
  AND2X1   g09814(.A(new_n10007_), .B(new_n9900_), .Y(new_n10008_));
  INVX1    g09815(.A(new_n10008_), .Y(new_n10009_));
  INVX1    g09816(.A(new_n9893_), .Y(new_n10010_));
  OAI21X1  g09817(.A0(new_n9894_), .A1(new_n9774_), .B0(new_n10010_), .Y(new_n10011_));
  NOR2X1   g09818(.A(new_n10007_), .B(new_n9900_), .Y(new_n10012_));
  INVX1    g09819(.A(new_n10012_), .Y(new_n10013_));
  AOI21X1  g09820(.A0(new_n10009_), .A1(new_n10013_), .B0(new_n10011_), .Y(new_n10014_));
  AND2X1   g09821(.A(new_n10013_), .B(new_n10011_), .Y(new_n10015_));
  AOI21X1  g09822(.A0(new_n10015_), .A1(new_n10009_), .B0(new_n10014_), .Y(\asquared[87] ));
  AOI21X1  g09823(.A0(new_n10013_), .A1(new_n10011_), .B0(new_n10008_), .Y(new_n10017_));
  AND2X1   g09824(.A(new_n9971_), .B(new_n9943_), .Y(new_n10018_));
  INVX1    g09825(.A(new_n10018_), .Y(new_n10019_));
  OAI21X1  g09826(.A0(new_n9972_), .A1(new_n9921_), .B0(new_n10019_), .Y(new_n10020_));
  INVX1    g09827(.A(new_n10020_), .Y(new_n10021_));
  NOR2X1   g09828(.A(new_n9823_), .B(new_n9800_), .Y(new_n10022_));
  AOI21X1  g09829(.A0(new_n9912_), .A1(new_n9817_), .B0(new_n10022_), .Y(new_n10023_));
  INVX1    g09830(.A(new_n9929_), .Y(new_n10024_));
  OR2X1    g09831(.A(new_n9935_), .B(new_n10024_), .Y(new_n10025_));
  OR2X1    g09832(.A(new_n9942_), .B(new_n9936_), .Y(new_n10026_));
  AND2X1   g09833(.A(new_n10026_), .B(new_n10025_), .Y(new_n10027_));
  XOR2X1   g09834(.A(new_n10027_), .B(new_n10023_), .Y(new_n10028_));
  AND2X1   g09835(.A(new_n9961_), .B(new_n9952_), .Y(new_n10029_));
  AND2X1   g09836(.A(new_n9970_), .B(new_n9962_), .Y(new_n10030_));
  OR2X1    g09837(.A(new_n10030_), .B(new_n10029_), .Y(new_n10031_));
  XOR2X1   g09838(.A(new_n10031_), .B(new_n10028_), .Y(new_n10032_));
  XOR2X1   g09839(.A(new_n10032_), .B(new_n10021_), .Y(new_n10033_));
  AND2X1   g09840(.A(new_n9998_), .B(new_n9850_), .Y(new_n10034_));
  INVX1    g09841(.A(new_n10034_), .Y(new_n10035_));
  OAI21X1  g09842(.A0(new_n10002_), .A1(new_n10000_), .B0(new_n10035_), .Y(new_n10036_));
  INVX1    g09843(.A(new_n10036_), .Y(new_n10037_));
  XOR2X1   g09844(.A(new_n10037_), .B(new_n10033_), .Y(new_n10038_));
  NOR2X1   g09845(.A(new_n9985_), .B(new_n9983_), .Y(new_n10039_));
  AOI21X1  g09846(.A0(new_n10003_), .A1(new_n9986_), .B0(new_n10039_), .Y(new_n10040_));
  XOR2X1   g09847(.A(new_n10040_), .B(new_n10038_), .Y(new_n10041_));
  AND2X1   g09848(.A(new_n9918_), .B(new_n9909_), .Y(new_n10042_));
  AOI21X1  g09849(.A0(new_n9973_), .A1(new_n9919_), .B0(new_n10042_), .Y(new_n10043_));
  INVX1    g09850(.A(new_n10043_), .Y(new_n10044_));
  AND2X1   g09851(.A(\a[62] ), .B(\a[44] ), .Y(new_n10045_));
  AOI21X1  g09852(.A0(new_n10045_), .A1(\a[25] ), .B0(new_n7353_), .Y(new_n10046_));
  AOI21X1  g09853(.A0(new_n10045_), .A1(\a[25] ), .B0(new_n4992_), .Y(new_n10047_));
  INVX1    g09854(.A(new_n10047_), .Y(new_n10048_));
  AOI21X1  g09855(.A0(\a[62] ), .A1(\a[25] ), .B0(\a[44] ), .Y(new_n10049_));
  OAI22X1  g09856(.A0(new_n10049_), .A1(new_n10048_), .B0(new_n10046_), .B1(new_n7353_), .Y(new_n10050_));
  INVX1    g09857(.A(new_n10050_), .Y(new_n10051_));
  AOI22X1  g09858(.A0(\a[56] ), .A1(\a[31] ), .B0(\a[54] ), .B1(\a[33] ), .Y(new_n10052_));
  AND2X1   g09859(.A(\a[47] ), .B(\a[40] ), .Y(new_n10053_));
  NOR3X1   g09860(.A(new_n2673_), .B(new_n6022_), .C(new_n4835_), .Y(new_n10054_));
  OAI21X1  g09861(.A0(new_n10052_), .A1(new_n10054_), .B0(new_n10053_), .Y(new_n10055_));
  NOR3X1   g09862(.A(new_n10052_), .B(new_n4041_), .C(new_n3036_), .Y(new_n10056_));
  OR2X1    g09863(.A(new_n10056_), .B(new_n10054_), .Y(new_n10057_));
  OAI21X1  g09864(.A0(new_n10057_), .A1(new_n10052_), .B0(new_n10055_), .Y(new_n10058_));
  XOR2X1   g09865(.A(new_n10058_), .B(new_n10051_), .Y(new_n10059_));
  AND2X1   g09866(.A(new_n9843_), .B(new_n9914_), .Y(new_n10060_));
  AOI21X1  g09867(.A0(new_n9915_), .A1(new_n9788_), .B0(new_n10060_), .Y(new_n10061_));
  XOR2X1   g09868(.A(new_n10061_), .B(new_n10059_), .Y(new_n10062_));
  NAND4X1  g09869(.A(\a[63] ), .B(\a[61] ), .C(\a[26] ), .D(\a[24] ), .Y(new_n10063_));
  NAND4X1  g09870(.A(\a[63] ), .B(\a[60] ), .C(\a[27] ), .D(\a[24] ), .Y(new_n10064_));
  AOI22X1  g09871(.A0(new_n10064_), .A1(new_n10063_), .B0(new_n6428_), .B1(new_n1995_), .Y(new_n10065_));
  NAND4X1  g09872(.A(\a[61] ), .B(\a[60] ), .C(\a[27] ), .D(\a[26] ), .Y(new_n10066_));
  NAND3X1  g09873(.A(new_n10064_), .B(new_n10063_), .C(new_n10066_), .Y(new_n10067_));
  AOI22X1  g09874(.A0(\a[61] ), .A1(\a[26] ), .B0(\a[60] ), .B1(\a[27] ), .Y(new_n10068_));
  NAND2X1  g09875(.A(\a[63] ), .B(\a[24] ), .Y(new_n10069_));
  OAI22X1  g09876(.A0(new_n10069_), .A1(new_n10065_), .B0(new_n10068_), .B1(new_n10067_), .Y(new_n10070_));
  NAND4X1  g09877(.A(\a[50] ), .B(\a[48] ), .C(\a[39] ), .D(\a[37] ), .Y(new_n10071_));
  NAND4X1  g09878(.A(\a[50] ), .B(\a[49] ), .C(\a[38] ), .D(\a[37] ), .Y(new_n10072_));
  AOI22X1  g09879(.A0(new_n10072_), .A1(new_n10071_), .B0(new_n4274_), .B1(new_n3503_), .Y(new_n10073_));
  NAND2X1  g09880(.A(\a[50] ), .B(\a[37] ), .Y(new_n10074_));
  AOI22X1  g09881(.A0(\a[49] ), .A1(\a[38] ), .B0(\a[48] ), .B1(\a[39] ), .Y(new_n10075_));
  AOI21X1  g09882(.A0(new_n4274_), .A1(new_n3503_), .B0(new_n10073_), .Y(new_n10076_));
  INVX1    g09883(.A(new_n10076_), .Y(new_n10077_));
  OAI22X1  g09884(.A0(new_n10077_), .A1(new_n10075_), .B0(new_n10074_), .B1(new_n10073_), .Y(new_n10078_));
  XOR2X1   g09885(.A(new_n10078_), .B(new_n10070_), .Y(new_n10079_));
  AND2X1   g09886(.A(\a[55] ), .B(\a[32] ), .Y(new_n10080_));
  INVX1    g09887(.A(new_n10080_), .Y(new_n10081_));
  AOI22X1  g09888(.A0(\a[46] ), .A1(\a[41] ), .B0(\a[45] ), .B1(\a[42] ), .Y(new_n10082_));
  AND2X1   g09889(.A(new_n3809_), .B(new_n3607_), .Y(new_n10083_));
  NOR3X1   g09890(.A(new_n10082_), .B(new_n10083_), .C(new_n10081_), .Y(new_n10084_));
  NOR2X1   g09891(.A(new_n10084_), .B(new_n10083_), .Y(new_n10085_));
  INVX1    g09892(.A(new_n10085_), .Y(new_n10086_));
  OAI22X1  g09893(.A0(new_n10086_), .A1(new_n10082_), .B0(new_n10084_), .B1(new_n10081_), .Y(new_n10087_));
  XOR2X1   g09894(.A(new_n10087_), .B(new_n10079_), .Y(new_n10088_));
  XOR2X1   g09895(.A(new_n10088_), .B(new_n10062_), .Y(new_n10089_));
  NOR4X1   g09896(.A(new_n5441_), .B(new_n5245_), .C(new_n2028_), .D(new_n1684_), .Y(new_n10090_));
  NAND4X1  g09897(.A(\a[59] ), .B(\a[57] ), .C(\a[30] ), .D(\a[28] ), .Y(new_n10091_));
  NAND4X1  g09898(.A(\a[59] ), .B(\a[53] ), .C(\a[34] ), .D(\a[28] ), .Y(new_n10092_));
  AOI21X1  g09899(.A0(new_n10092_), .A1(new_n10091_), .B0(new_n10090_), .Y(new_n10093_));
  NAND2X1  g09900(.A(\a[59] ), .B(\a[28] ), .Y(new_n10094_));
  OR2X1    g09901(.A(new_n10093_), .B(new_n10090_), .Y(new_n10095_));
  AOI22X1  g09902(.A0(\a[57] ), .A1(\a[30] ), .B0(\a[53] ), .B1(\a[34] ), .Y(new_n10096_));
  OAI22X1  g09903(.A0(new_n10096_), .A1(new_n10095_), .B0(new_n10094_), .B1(new_n10093_), .Y(new_n10097_));
  OAI22X1  g09904(.A0(new_n9989_), .A1(new_n9806_), .B0(new_n6557_), .B1(new_n1772_), .Y(new_n10098_));
  INVX1    g09905(.A(new_n10098_), .Y(new_n10099_));
  XOR2X1   g09906(.A(new_n10099_), .B(new_n10097_), .Y(new_n10100_));
  AND2X1   g09907(.A(\a[52] ), .B(\a[29] ), .Y(new_n10101_));
  AND2X1   g09908(.A(\a[58] ), .B(\a[35] ), .Y(new_n10102_));
  AOI22X1  g09909(.A0(new_n10102_), .A1(new_n10101_), .B0(new_n7164_), .B1(new_n2682_), .Y(new_n10103_));
  NOR4X1   g09910(.A(new_n5379_), .B(new_n4349_), .C(new_n2583_), .D(new_n1803_), .Y(new_n10104_));
  NOR2X1   g09911(.A(new_n10104_), .B(new_n10103_), .Y(new_n10105_));
  NOR3X1   g09912(.A(new_n10105_), .B(new_n4354_), .C(new_n2557_), .Y(new_n10106_));
  INVX1    g09913(.A(new_n10104_), .Y(new_n10107_));
  AND2X1   g09914(.A(new_n10107_), .B(new_n10103_), .Y(new_n10108_));
  OAI22X1  g09915(.A0(new_n5379_), .A1(new_n1803_), .B0(new_n4349_), .B1(new_n2583_), .Y(new_n10109_));
  AOI21X1  g09916(.A0(new_n10109_), .A1(new_n10108_), .B0(new_n10106_), .Y(new_n10110_));
  XOR2X1   g09917(.A(new_n10110_), .B(new_n10100_), .Y(new_n10111_));
  XOR2X1   g09918(.A(new_n10111_), .B(new_n10089_), .Y(new_n10112_));
  XOR2X1   g09919(.A(new_n10112_), .B(new_n10044_), .Y(new_n10113_));
  INVX1    g09920(.A(new_n10113_), .Y(new_n10114_));
  NOR2X1   g09921(.A(new_n9916_), .B(new_n9913_), .Y(new_n10115_));
  AOI21X1  g09922(.A0(new_n9917_), .A1(new_n9911_), .B0(new_n10115_), .Y(new_n10116_));
  AND2X1   g09923(.A(new_n9905_), .B(new_n9902_), .Y(new_n10117_));
  AOI21X1  g09924(.A0(new_n9908_), .A1(new_n9906_), .B0(new_n10117_), .Y(new_n10118_));
  XOR2X1   g09925(.A(new_n10118_), .B(new_n10116_), .Y(new_n10119_));
  NAND2X1  g09926(.A(new_n9993_), .B(new_n9991_), .Y(new_n10120_));
  OAI21X1  g09927(.A0(new_n9997_), .A1(new_n9995_), .B0(new_n10120_), .Y(new_n10121_));
  INVX1    g09928(.A(new_n9941_), .Y(new_n10122_));
  XOR2X1   g09929(.A(new_n9969_), .B(new_n9959_), .Y(new_n10123_));
  XOR2X1   g09930(.A(new_n10123_), .B(new_n10122_), .Y(new_n10124_));
  INVX1    g09931(.A(new_n9933_), .Y(new_n10125_));
  XOR2X1   g09932(.A(new_n9949_), .B(new_n10125_), .Y(new_n10126_));
  XOR2X1   g09933(.A(new_n10126_), .B(new_n9928_), .Y(new_n10127_));
  XOR2X1   g09934(.A(new_n10127_), .B(new_n10124_), .Y(new_n10128_));
  XOR2X1   g09935(.A(new_n10128_), .B(new_n10121_), .Y(new_n10129_));
  XOR2X1   g09936(.A(new_n10129_), .B(new_n10119_), .Y(new_n10130_));
  XOR2X1   g09937(.A(new_n10130_), .B(new_n10114_), .Y(new_n10131_));
  XOR2X1   g09938(.A(new_n10131_), .B(new_n10041_), .Y(new_n10132_));
  NOR3X1   g09939(.A(new_n10132_), .B(new_n10005_), .C(new_n9978_), .Y(new_n10133_));
  OR2X1    g09940(.A(new_n10005_), .B(new_n9978_), .Y(new_n10134_));
  AND2X1   g09941(.A(new_n10132_), .B(new_n10134_), .Y(new_n10135_));
  OR2X1    g09942(.A(new_n10135_), .B(new_n10133_), .Y(new_n10136_));
  XOR2X1   g09943(.A(new_n10136_), .B(new_n10017_), .Y(\asquared[88] ));
  INVX1    g09944(.A(new_n10038_), .Y(new_n10138_));
  NOR2X1   g09945(.A(new_n10040_), .B(new_n10138_), .Y(new_n10139_));
  NOR2X1   g09946(.A(new_n10131_), .B(new_n10041_), .Y(new_n10140_));
  NOR2X1   g09947(.A(new_n10140_), .B(new_n10139_), .Y(new_n10141_));
  AND2X1   g09948(.A(new_n10112_), .B(new_n10044_), .Y(new_n10142_));
  AOI21X1  g09949(.A0(new_n10130_), .A1(new_n10113_), .B0(new_n10142_), .Y(new_n10143_));
  INVX1    g09950(.A(new_n10143_), .Y(new_n10144_));
  NOR2X1   g09951(.A(new_n10118_), .B(new_n10116_), .Y(new_n10145_));
  AOI21X1  g09952(.A0(new_n10129_), .A1(new_n10119_), .B0(new_n10145_), .Y(new_n10146_));
  AND2X1   g09953(.A(new_n9949_), .B(new_n10125_), .Y(new_n10147_));
  AOI21X1  g09954(.A0(new_n10126_), .A1(new_n9928_), .B0(new_n10147_), .Y(new_n10148_));
  NOR2X1   g09955(.A(new_n10110_), .B(new_n10100_), .Y(new_n10149_));
  AOI21X1  g09956(.A0(new_n10098_), .A1(new_n10097_), .B0(new_n10149_), .Y(new_n10150_));
  XOR2X1   g09957(.A(new_n10150_), .B(new_n10148_), .Y(new_n10151_));
  AND2X1   g09958(.A(new_n10078_), .B(new_n10070_), .Y(new_n10152_));
  AND2X1   g09959(.A(new_n10087_), .B(new_n10079_), .Y(new_n10153_));
  OR2X1    g09960(.A(new_n10153_), .B(new_n10152_), .Y(new_n10154_));
  XOR2X1   g09961(.A(new_n10154_), .B(new_n10151_), .Y(new_n10155_));
  INVX1    g09962(.A(new_n10155_), .Y(new_n10156_));
  NAND2X1  g09963(.A(new_n10088_), .B(new_n10062_), .Y(new_n10157_));
  NAND2X1  g09964(.A(new_n10111_), .B(new_n10089_), .Y(new_n10158_));
  NAND2X1  g09965(.A(new_n10158_), .B(new_n10157_), .Y(new_n10159_));
  XOR2X1   g09966(.A(new_n10159_), .B(new_n10156_), .Y(new_n10160_));
  XOR2X1   g09967(.A(new_n10160_), .B(new_n10146_), .Y(new_n10161_));
  XOR2X1   g09968(.A(new_n10161_), .B(new_n10144_), .Y(new_n10162_));
  NAND2X1  g09969(.A(new_n10032_), .B(new_n10020_), .Y(new_n10163_));
  OAI21X1  g09970(.A0(new_n10037_), .A1(new_n10033_), .B0(new_n10163_), .Y(new_n10164_));
  OAI22X1  g09971(.A0(new_n6557_), .A1(new_n3483_), .B0(new_n6555_), .B1(new_n3570_), .Y(new_n10165_));
  OAI21X1  g09972(.A0(new_n6554_), .A1(new_n1672_), .B0(new_n10165_), .Y(new_n10166_));
  AOI21X1  g09973(.A0(new_n6428_), .A1(new_n1671_), .B0(new_n10165_), .Y(new_n10167_));
  OAI22X1  g09974(.A0(new_n6023_), .A1(new_n1679_), .B0(new_n5952_), .B1(new_n1431_), .Y(new_n10168_));
  AND2X1   g09975(.A(\a[62] ), .B(\a[26] ), .Y(new_n10169_));
  AOI22X1  g09976(.A0(new_n10169_), .A1(new_n10166_), .B0(new_n10168_), .B1(new_n10167_), .Y(new_n10170_));
  AND2X1   g09977(.A(\a[57] ), .B(\a[31] ), .Y(new_n10171_));
  INVX1    g09978(.A(new_n10171_), .Y(new_n10172_));
  AOI22X1  g09979(.A0(\a[47] ), .A1(\a[41] ), .B0(\a[46] ), .B1(\a[42] ), .Y(new_n10173_));
  AND2X1   g09980(.A(new_n3893_), .B(new_n3607_), .Y(new_n10174_));
  NOR3X1   g09981(.A(new_n10173_), .B(new_n10174_), .C(new_n10172_), .Y(new_n10175_));
  INVX1    g09982(.A(new_n10173_), .Y(new_n10176_));
  AOI21X1  g09983(.A0(new_n10176_), .A1(new_n10171_), .B0(new_n10174_), .Y(new_n10177_));
  INVX1    g09984(.A(new_n10177_), .Y(new_n10178_));
  OAI22X1  g09985(.A0(new_n10178_), .A1(new_n10173_), .B0(new_n10175_), .B1(new_n10172_), .Y(new_n10179_));
  XOR2X1   g09986(.A(new_n10179_), .B(new_n10170_), .Y(new_n10180_));
  OAI22X1  g09987(.A0(new_n7336_), .A1(new_n5417_), .B0(new_n8145_), .B1(new_n6527_), .Y(new_n10181_));
  OAI21X1  g09988(.A0(new_n7793_), .A1(new_n6525_), .B0(new_n10181_), .Y(new_n10182_));
  AND2X1   g09989(.A(\a[53] ), .B(\a[35] ), .Y(new_n10183_));
  AOI21X1  g09990(.A0(new_n7164_), .A1(new_n3330_), .B0(new_n10181_), .Y(new_n10184_));
  OAI22X1  g09991(.A0(new_n4354_), .A1(new_n2583_), .B0(new_n4349_), .B1(new_n2345_), .Y(new_n10185_));
  AOI22X1  g09992(.A0(new_n10185_), .A1(new_n10184_), .B0(new_n10183_), .B1(new_n10182_), .Y(new_n10186_));
  XOR2X1   g09993(.A(new_n10186_), .B(new_n10180_), .Y(new_n10187_));
  AOI22X1  g09994(.A0(\a[50] ), .A1(\a[38] ), .B0(\a[49] ), .B1(\a[39] ), .Y(new_n10188_));
  AND2X1   g09995(.A(\a[59] ), .B(\a[29] ), .Y(new_n10189_));
  INVX1    g09996(.A(new_n10189_), .Y(new_n10190_));
  AND2X1   g09997(.A(new_n4321_), .B(new_n3503_), .Y(new_n10191_));
  NOR3X1   g09998(.A(new_n10190_), .B(new_n10191_), .C(new_n10188_), .Y(new_n10192_));
  INVX1    g09999(.A(new_n10188_), .Y(new_n10193_));
  AOI21X1  g10000(.A0(new_n10189_), .A1(new_n10193_), .B0(new_n10191_), .Y(new_n10194_));
  INVX1    g10001(.A(new_n10194_), .Y(new_n10195_));
  OAI22X1  g10002(.A0(new_n10195_), .A1(new_n10188_), .B0(new_n10192_), .B1(new_n10190_), .Y(new_n10196_));
  AOI22X1  g10003(.A0(\a[58] ), .A1(\a[30] ), .B0(\a[56] ), .B1(\a[32] ), .Y(new_n10197_));
  INVX1    g10004(.A(new_n10197_), .Y(new_n10198_));
  NAND4X1  g10005(.A(\a[58] ), .B(\a[56] ), .C(\a[32] ), .D(\a[30] ), .Y(new_n10199_));
  NAND3X1  g10006(.A(new_n10198_), .B(new_n10199_), .C(new_n5004_), .Y(new_n10200_));
  AOI22X1  g10007(.A0(new_n10198_), .A1(new_n5004_), .B0(new_n5381_), .B1(new_n1787_), .Y(new_n10201_));
  AOI22X1  g10008(.A0(new_n10201_), .A1(new_n10198_), .B0(new_n10200_), .B1(new_n5004_), .Y(new_n10202_));
  XOR2X1   g10009(.A(new_n10202_), .B(new_n10196_), .Y(new_n10203_));
  AND2X1   g10010(.A(new_n9969_), .B(new_n9959_), .Y(new_n10204_));
  AOI21X1  g10011(.A0(new_n10123_), .A1(new_n10122_), .B0(new_n10204_), .Y(new_n10205_));
  XOR2X1   g10012(.A(new_n10205_), .B(new_n10203_), .Y(new_n10206_));
  AND2X1   g10013(.A(\a[63] ), .B(\a[25] ), .Y(new_n10207_));
  XOR2X1   g10014(.A(new_n10207_), .B(new_n10048_), .Y(new_n10208_));
  XOR2X1   g10015(.A(new_n10208_), .B(new_n10086_), .Y(new_n10209_));
  XOR2X1   g10016(.A(new_n10209_), .B(new_n10206_), .Y(new_n10210_));
  XOR2X1   g10017(.A(new_n10210_), .B(new_n10187_), .Y(new_n10211_));
  XOR2X1   g10018(.A(new_n10211_), .B(new_n10164_), .Y(new_n10212_));
  INVX1    g10019(.A(new_n10212_), .Y(new_n10213_));
  AND2X1   g10020(.A(new_n10127_), .B(new_n10124_), .Y(new_n10214_));
  AOI21X1  g10021(.A0(new_n10128_), .A1(new_n10121_), .B0(new_n10214_), .Y(new_n10215_));
  AOI21X1  g10022(.A0(new_n10026_), .A1(new_n10025_), .B0(new_n10023_), .Y(new_n10216_));
  AOI21X1  g10023(.A0(new_n10031_), .A1(new_n10028_), .B0(new_n10216_), .Y(new_n10217_));
  XOR2X1   g10024(.A(new_n10217_), .B(new_n10215_), .Y(new_n10218_));
  XOR2X1   g10025(.A(new_n10095_), .B(new_n10067_), .Y(new_n10219_));
  XOR2X1   g10026(.A(new_n10219_), .B(new_n10076_), .Y(new_n10220_));
  XOR2X1   g10027(.A(new_n10108_), .B(new_n10057_), .Y(new_n10221_));
  AOI22X1  g10028(.A0(\a[55] ), .A1(\a[33] ), .B0(\a[54] ), .B1(\a[34] ), .Y(new_n10222_));
  AND2X1   g10029(.A(new_n5240_), .B(new_n2918_), .Y(new_n10223_));
  NOR3X1   g10030(.A(new_n10222_), .B(new_n10223_), .C(new_n7641_), .Y(new_n10224_));
  INVX1    g10031(.A(new_n10222_), .Y(new_n10225_));
  AOI21X1  g10032(.A0(new_n10225_), .A1(new_n7640_), .B0(new_n10223_), .Y(new_n10226_));
  INVX1    g10033(.A(new_n10226_), .Y(new_n10227_));
  OAI22X1  g10034(.A0(new_n10227_), .A1(new_n10222_), .B0(new_n10224_), .B1(new_n7641_), .Y(new_n10228_));
  XOR2X1   g10035(.A(new_n10228_), .B(new_n10221_), .Y(new_n10229_));
  AND2X1   g10036(.A(new_n10058_), .B(new_n10050_), .Y(new_n10230_));
  NOR2X1   g10037(.A(new_n10061_), .B(new_n10059_), .Y(new_n10231_));
  OR2X1    g10038(.A(new_n10231_), .B(new_n10230_), .Y(new_n10232_));
  XOR2X1   g10039(.A(new_n10232_), .B(new_n10229_), .Y(new_n10233_));
  XOR2X1   g10040(.A(new_n10233_), .B(new_n10220_), .Y(new_n10234_));
  XOR2X1   g10041(.A(new_n10234_), .B(new_n10218_), .Y(new_n10235_));
  XOR2X1   g10042(.A(new_n10235_), .B(new_n10213_), .Y(new_n10236_));
  XOR2X1   g10043(.A(new_n10236_), .B(new_n10162_), .Y(new_n10237_));
  XOR2X1   g10044(.A(new_n10237_), .B(new_n10141_), .Y(new_n10238_));
  INVX1    g10045(.A(new_n10135_), .Y(new_n10239_));
  OAI21X1  g10046(.A0(new_n10133_), .A1(new_n10017_), .B0(new_n10239_), .Y(new_n10240_));
  XOR2X1   g10047(.A(new_n10240_), .B(new_n10238_), .Y(\asquared[89] ));
  AND2X1   g10048(.A(new_n10161_), .B(new_n10144_), .Y(new_n10242_));
  INVX1    g10049(.A(new_n10242_), .Y(new_n10243_));
  INVX1    g10050(.A(new_n10162_), .Y(new_n10244_));
  OAI21X1  g10051(.A0(new_n10236_), .A1(new_n10244_), .B0(new_n10243_), .Y(new_n10245_));
  INVX1    g10052(.A(new_n10245_), .Y(new_n10246_));
  NOR2X1   g10053(.A(new_n10217_), .B(new_n10215_), .Y(new_n10247_));
  AOI21X1  g10054(.A0(new_n10234_), .A1(new_n10218_), .B0(new_n10247_), .Y(new_n10248_));
  AND2X1   g10055(.A(new_n10209_), .B(new_n10206_), .Y(new_n10249_));
  AOI21X1  g10056(.A0(new_n10210_), .A1(new_n10187_), .B0(new_n10249_), .Y(new_n10250_));
  INVX1    g10057(.A(new_n10250_), .Y(new_n10251_));
  INVX1    g10058(.A(new_n10196_), .Y(new_n10252_));
  OR2X1    g10059(.A(new_n10202_), .B(new_n10252_), .Y(new_n10253_));
  OAI21X1  g10060(.A0(new_n10205_), .A1(new_n10203_), .B0(new_n10253_), .Y(new_n10254_));
  INVX1    g10061(.A(new_n10179_), .Y(new_n10255_));
  OR2X1    g10062(.A(new_n10255_), .B(new_n10170_), .Y(new_n10256_));
  OAI21X1  g10063(.A0(new_n10186_), .A1(new_n10180_), .B0(new_n10256_), .Y(new_n10257_));
  XOR2X1   g10064(.A(new_n10257_), .B(new_n10254_), .Y(new_n10258_));
  XOR2X1   g10065(.A(new_n10194_), .B(new_n10178_), .Y(new_n10259_));
  AND2X1   g10066(.A(\a[63] ), .B(\a[26] ), .Y(new_n10260_));
  AOI22X1  g10067(.A0(\a[50] ), .A1(\a[39] ), .B0(\a[49] ), .B1(\a[40] ), .Y(new_n10261_));
  INVX1    g10068(.A(new_n10261_), .Y(new_n10262_));
  NAND4X1  g10069(.A(\a[50] ), .B(\a[49] ), .C(\a[40] ), .D(\a[39] ), .Y(new_n10263_));
  NAND3X1  g10070(.A(new_n10262_), .B(new_n10263_), .C(new_n10260_), .Y(new_n10264_));
  AOI22X1  g10071(.A0(new_n10262_), .A1(new_n10260_), .B0(new_n4321_), .B1(new_n4077_), .Y(new_n10265_));
  AOI22X1  g10072(.A0(new_n10265_), .A1(new_n10262_), .B0(new_n10264_), .B1(new_n10260_), .Y(new_n10266_));
  XOR2X1   g10073(.A(new_n10266_), .B(new_n10259_), .Y(new_n10267_));
  XOR2X1   g10074(.A(new_n10267_), .B(new_n10258_), .Y(new_n10268_));
  XOR2X1   g10075(.A(new_n10268_), .B(new_n10251_), .Y(new_n10269_));
  INVX1    g10076(.A(new_n10269_), .Y(new_n10270_));
  XOR2X1   g10077(.A(new_n10270_), .B(new_n10248_), .Y(new_n10271_));
  AND2X1   g10078(.A(new_n10211_), .B(new_n10164_), .Y(new_n10272_));
  AOI21X1  g10079(.A0(new_n10235_), .A1(new_n10212_), .B0(new_n10272_), .Y(new_n10273_));
  OR2X1    g10080(.A(new_n10273_), .B(new_n10271_), .Y(new_n10274_));
  NAND2X1  g10081(.A(new_n10159_), .B(new_n10155_), .Y(new_n10275_));
  OAI21X1  g10082(.A0(new_n10160_), .A1(new_n10146_), .B0(new_n10275_), .Y(new_n10276_));
  AOI22X1  g10083(.A0(\a[56] ), .A1(\a[33] ), .B0(\a[54] ), .B1(\a[35] ), .Y(new_n10277_));
  AND2X1   g10084(.A(\a[48] ), .B(\a[41] ), .Y(new_n10278_));
  INVX1    g10085(.A(new_n10278_), .Y(new_n10279_));
  AND2X1   g10086(.A(new_n5042_), .B(new_n2120_), .Y(new_n10280_));
  NOR3X1   g10087(.A(new_n10279_), .B(new_n10280_), .C(new_n10277_), .Y(new_n10281_));
  NOR2X1   g10088(.A(new_n10281_), .B(new_n10280_), .Y(new_n10282_));
  INVX1    g10089(.A(new_n10282_), .Y(new_n10283_));
  OAI22X1  g10090(.A0(new_n10283_), .A1(new_n10277_), .B0(new_n10281_), .B1(new_n10279_), .Y(new_n10284_));
  OAI22X1  g10091(.A0(new_n7336_), .A1(new_n6525_), .B0(new_n8145_), .B1(new_n7316_), .Y(new_n10285_));
  OAI21X1  g10092(.A0(new_n7793_), .A1(new_n7317_), .B0(new_n10285_), .Y(new_n10286_));
  AND2X1   g10093(.A(\a[53] ), .B(\a[36] ), .Y(new_n10287_));
  AOI21X1  g10094(.A0(new_n7164_), .A1(new_n3164_), .B0(new_n10285_), .Y(new_n10288_));
  OAI22X1  g10095(.A0(new_n4354_), .A1(new_n2345_), .B0(new_n4349_), .B1(new_n2519_), .Y(new_n10289_));
  AOI22X1  g10096(.A0(new_n10289_), .A1(new_n10288_), .B0(new_n10287_), .B1(new_n10286_), .Y(new_n10290_));
  XOR2X1   g10097(.A(new_n10290_), .B(new_n10284_), .Y(new_n10291_));
  OAI22X1  g10098(.A0(new_n6793_), .A1(new_n2076_), .B0(new_n8155_), .B1(new_n4923_), .Y(new_n10292_));
  OAI21X1  g10099(.A0(new_n8154_), .A1(new_n2672_), .B0(new_n10292_), .Y(new_n10293_));
  AND2X1   g10100(.A(\a[59] ), .B(\a[30] ), .Y(new_n10294_));
  AOI21X1  g10101(.A0(new_n6119_), .A1(new_n2671_), .B0(new_n10292_), .Y(new_n10295_));
  OAI22X1  g10102(.A0(new_n5379_), .A1(new_n1704_), .B0(new_n5441_), .B1(new_n2219_), .Y(new_n10296_));
  AOI22X1  g10103(.A0(new_n10296_), .A1(new_n10295_), .B0(new_n10294_), .B1(new_n10293_), .Y(new_n10297_));
  XOR2X1   g10104(.A(new_n10297_), .B(new_n10291_), .Y(new_n10298_));
  INVX1    g10105(.A(new_n10201_), .Y(new_n10299_));
  XOR2X1   g10106(.A(new_n10184_), .B(new_n10167_), .Y(new_n10300_));
  XOR2X1   g10107(.A(new_n10300_), .B(new_n10299_), .Y(new_n10301_));
  AND2X1   g10108(.A(\a[62] ), .B(\a[45] ), .Y(new_n10302_));
  AOI21X1  g10109(.A0(new_n10302_), .A1(\a[27] ), .B0(new_n7642_), .Y(new_n10303_));
  AOI21X1  g10110(.A0(new_n10302_), .A1(\a[27] ), .B0(new_n3918_), .Y(new_n10304_));
  INVX1    g10111(.A(new_n10304_), .Y(new_n10305_));
  AOI21X1  g10112(.A0(\a[62] ), .A1(\a[27] ), .B0(\a[45] ), .Y(new_n10306_));
  OAI22X1  g10113(.A0(new_n10306_), .A1(new_n10305_), .B0(new_n10303_), .B1(new_n7642_), .Y(new_n10307_));
  AND2X1   g10114(.A(\a[55] ), .B(\a[34] ), .Y(new_n10308_));
  AND2X1   g10115(.A(new_n3893_), .B(new_n3462_), .Y(new_n10309_));
  AOI22X1  g10116(.A0(\a[47] ), .A1(\a[42] ), .B0(\a[46] ), .B1(\a[43] ), .Y(new_n10310_));
  OR4X1    g10117(.A(new_n10310_), .B(new_n10309_), .C(new_n4906_), .D(new_n2028_), .Y(new_n10311_));
  NOR3X1   g10118(.A(new_n10310_), .B(new_n10309_), .C(new_n10308_), .Y(new_n10312_));
  AOI21X1  g10119(.A0(new_n10311_), .A1(new_n10308_), .B0(new_n10312_), .Y(new_n10313_));
  XOR2X1   g10120(.A(new_n10313_), .B(new_n10307_), .Y(new_n10314_));
  NAND2X1  g10121(.A(\a[60] ), .B(\a[29] ), .Y(new_n10315_));
  NAND2X1  g10122(.A(\a[61] ), .B(\a[28] ), .Y(new_n10316_));
  AOI22X1  g10123(.A0(new_n10316_), .A1(new_n10315_), .B0(new_n6428_), .B1(new_n1674_), .Y(new_n10317_));
  XOR2X1   g10124(.A(new_n10317_), .B(new_n10226_), .Y(new_n10318_));
  INVX1    g10125(.A(new_n10318_), .Y(new_n10319_));
  XOR2X1   g10126(.A(new_n10319_), .B(new_n10314_), .Y(new_n10320_));
  XOR2X1   g10127(.A(new_n10320_), .B(new_n10301_), .Y(new_n10321_));
  XOR2X1   g10128(.A(new_n10321_), .B(new_n10298_), .Y(new_n10322_));
  XOR2X1   g10129(.A(new_n10322_), .B(new_n10276_), .Y(new_n10323_));
  AND2X1   g10130(.A(new_n10095_), .B(new_n10067_), .Y(new_n10324_));
  AOI21X1  g10131(.A0(new_n10219_), .A1(new_n10077_), .B0(new_n10324_), .Y(new_n10325_));
  NAND2X1  g10132(.A(new_n10207_), .B(new_n10048_), .Y(new_n10326_));
  NOR2X1   g10133(.A(new_n10207_), .B(new_n10048_), .Y(new_n10327_));
  OAI21X1  g10134(.A0(new_n10327_), .A1(new_n10085_), .B0(new_n10326_), .Y(new_n10328_));
  XOR2X1   g10135(.A(new_n10328_), .B(new_n10325_), .Y(new_n10329_));
  OAI21X1  g10136(.A0(new_n10105_), .A1(new_n10104_), .B0(new_n10057_), .Y(new_n10330_));
  INVX1    g10137(.A(new_n10228_), .Y(new_n10331_));
  OAI21X1  g10138(.A0(new_n10331_), .A1(new_n10221_), .B0(new_n10330_), .Y(new_n10332_));
  XOR2X1   g10139(.A(new_n10332_), .B(new_n10329_), .Y(new_n10333_));
  NOR2X1   g10140(.A(new_n10150_), .B(new_n10148_), .Y(new_n10334_));
  AOI21X1  g10141(.A0(new_n10154_), .A1(new_n10151_), .B0(new_n10334_), .Y(new_n10335_));
  XOR2X1   g10142(.A(new_n10335_), .B(new_n10333_), .Y(new_n10336_));
  INVX1    g10143(.A(new_n10229_), .Y(new_n10337_));
  OAI21X1  g10144(.A0(new_n10231_), .A1(new_n10230_), .B0(new_n10337_), .Y(new_n10338_));
  OAI21X1  g10145(.A0(new_n10233_), .A1(new_n10220_), .B0(new_n10338_), .Y(new_n10339_));
  XOR2X1   g10146(.A(new_n10339_), .B(new_n10336_), .Y(new_n10340_));
  XOR2X1   g10147(.A(new_n10340_), .B(new_n10323_), .Y(new_n10341_));
  XOR2X1   g10148(.A(new_n10273_), .B(new_n10271_), .Y(new_n10342_));
  NOR2X1   g10149(.A(new_n10342_), .B(new_n10341_), .Y(new_n10343_));
  INVX1    g10150(.A(new_n10341_), .Y(new_n10344_));
  AOI21X1  g10151(.A0(new_n10273_), .A1(new_n10271_), .B0(new_n10344_), .Y(new_n10345_));
  AOI21X1  g10152(.A0(new_n10345_), .A1(new_n10274_), .B0(new_n10343_), .Y(new_n10346_));
  XOR2X1   g10153(.A(new_n10346_), .B(new_n10246_), .Y(new_n10347_));
  AND2X1   g10154(.A(new_n10237_), .B(new_n10141_), .Y(new_n10348_));
  INVX1    g10155(.A(new_n10348_), .Y(new_n10349_));
  NOR2X1   g10156(.A(new_n10237_), .B(new_n10141_), .Y(new_n10350_));
  AOI21X1  g10157(.A0(new_n10240_), .A1(new_n10349_), .B0(new_n10350_), .Y(new_n10351_));
  XOR2X1   g10158(.A(new_n10351_), .B(new_n10347_), .Y(\asquared[90] ));
  INVX1    g10159(.A(new_n10271_), .Y(new_n10353_));
  NOR2X1   g10160(.A(new_n10273_), .B(new_n10353_), .Y(new_n10354_));
  NOR2X1   g10161(.A(new_n10335_), .B(new_n10333_), .Y(new_n10355_));
  AOI21X1  g10162(.A0(new_n10339_), .A1(new_n10336_), .B0(new_n10355_), .Y(new_n10356_));
  INVX1    g10163(.A(new_n10301_), .Y(new_n10357_));
  NOR2X1   g10164(.A(new_n10320_), .B(new_n10357_), .Y(new_n10358_));
  INVX1    g10165(.A(new_n10321_), .Y(new_n10359_));
  AOI21X1  g10166(.A0(new_n10359_), .A1(new_n10298_), .B0(new_n10358_), .Y(new_n10360_));
  NOR3X1   g10167(.A(new_n10310_), .B(new_n4906_), .C(new_n2028_), .Y(new_n10361_));
  OR2X1    g10168(.A(new_n10361_), .B(new_n10309_), .Y(new_n10362_));
  XOR2X1   g10169(.A(new_n10362_), .B(new_n10305_), .Y(new_n10363_));
  XOR2X1   g10170(.A(new_n10363_), .B(new_n10283_), .Y(new_n10364_));
  AND2X1   g10171(.A(new_n10311_), .B(new_n10308_), .Y(new_n10365_));
  OAI21X1  g10172(.A0(new_n10312_), .A1(new_n10365_), .B0(new_n10307_), .Y(new_n10366_));
  OAI21X1  g10173(.A0(new_n10318_), .A1(new_n10314_), .B0(new_n10366_), .Y(new_n10367_));
  INVX1    g10174(.A(new_n10284_), .Y(new_n10368_));
  OR2X1    g10175(.A(new_n10290_), .B(new_n10368_), .Y(new_n10369_));
  OAI21X1  g10176(.A0(new_n10297_), .A1(new_n10291_), .B0(new_n10369_), .Y(new_n10370_));
  XOR2X1   g10177(.A(new_n10370_), .B(new_n10367_), .Y(new_n10371_));
  XOR2X1   g10178(.A(new_n10371_), .B(new_n10364_), .Y(new_n10372_));
  INVX1    g10179(.A(new_n10372_), .Y(new_n10373_));
  XOR2X1   g10180(.A(new_n10373_), .B(new_n10360_), .Y(new_n10374_));
  INVX1    g10181(.A(new_n10374_), .Y(new_n10375_));
  XOR2X1   g10182(.A(new_n10375_), .B(new_n10356_), .Y(new_n10376_));
  INVX1    g10183(.A(new_n10376_), .Y(new_n10377_));
  INVX1    g10184(.A(new_n10322_), .Y(new_n10378_));
  AND2X1   g10185(.A(new_n10378_), .B(new_n10276_), .Y(new_n10379_));
  INVX1    g10186(.A(new_n10323_), .Y(new_n10380_));
  AOI21X1  g10187(.A0(new_n10340_), .A1(new_n10380_), .B0(new_n10379_), .Y(new_n10381_));
  XOR2X1   g10188(.A(new_n10381_), .B(new_n10377_), .Y(new_n10382_));
  NAND2X1  g10189(.A(new_n10268_), .B(new_n10251_), .Y(new_n10383_));
  OAI21X1  g10190(.A0(new_n10270_), .A1(new_n10248_), .B0(new_n10383_), .Y(new_n10384_));
  INVX1    g10191(.A(new_n10265_), .Y(new_n10385_));
  XOR2X1   g10192(.A(new_n10295_), .B(new_n10288_), .Y(new_n10386_));
  XOR2X1   g10193(.A(new_n10386_), .B(new_n10385_), .Y(new_n10387_));
  AND2X1   g10194(.A(new_n10219_), .B(new_n10077_), .Y(new_n10388_));
  OAI21X1  g10195(.A0(new_n10388_), .A1(new_n10324_), .B0(new_n10328_), .Y(new_n10389_));
  INVX1    g10196(.A(new_n10332_), .Y(new_n10390_));
  OAI21X1  g10197(.A0(new_n10390_), .A1(new_n10329_), .B0(new_n10389_), .Y(new_n10391_));
  XOR2X1   g10198(.A(new_n10391_), .B(new_n10387_), .Y(new_n10392_));
  INVX1    g10199(.A(new_n10392_), .Y(new_n10393_));
  AOI22X1  g10200(.A0(\a[57] ), .A1(\a[33] ), .B0(\a[56] ), .B1(\a[34] ), .Y(new_n10394_));
  NAND4X1  g10201(.A(\a[57] ), .B(\a[55] ), .C(\a[35] ), .D(\a[33] ), .Y(new_n10395_));
  NAND4X1  g10202(.A(\a[56] ), .B(\a[55] ), .C(\a[35] ), .D(\a[34] ), .Y(new_n10396_));
  AOI22X1  g10203(.A0(new_n10396_), .A1(new_n10395_), .B0(new_n5554_), .B1(new_n2918_), .Y(new_n10397_));
  AOI21X1  g10204(.A0(new_n5554_), .A1(new_n2918_), .B0(new_n10397_), .Y(new_n10398_));
  INVX1    g10205(.A(new_n10398_), .Y(new_n10399_));
  NAND2X1  g10206(.A(\a[55] ), .B(\a[35] ), .Y(new_n10400_));
  OAI22X1  g10207(.A0(new_n10400_), .A1(new_n10397_), .B0(new_n10399_), .B1(new_n10394_), .Y(new_n10401_));
  NAND4X1  g10208(.A(\a[54] ), .B(\a[52] ), .C(\a[38] ), .D(\a[36] ), .Y(new_n10402_));
  NAND4X1  g10209(.A(\a[54] ), .B(\a[53] ), .C(\a[37] ), .D(\a[36] ), .Y(new_n10403_));
  AOI22X1  g10210(.A0(new_n10403_), .A1(new_n10402_), .B0(new_n5048_), .B1(new_n3164_), .Y(new_n10404_));
  NAND2X1  g10211(.A(\a[54] ), .B(\a[36] ), .Y(new_n10405_));
  NAND4X1  g10212(.A(\a[53] ), .B(\a[52] ), .C(\a[38] ), .D(\a[37] ), .Y(new_n10406_));
  NAND3X1  g10213(.A(new_n10403_), .B(new_n10402_), .C(new_n10406_), .Y(new_n10407_));
  AOI22X1  g10214(.A0(\a[53] ), .A1(\a[37] ), .B0(\a[52] ), .B1(\a[38] ), .Y(new_n10408_));
  OAI22X1  g10215(.A0(new_n10408_), .A1(new_n10407_), .B0(new_n10405_), .B1(new_n10404_), .Y(new_n10409_));
  XOR2X1   g10216(.A(new_n10409_), .B(new_n10401_), .Y(new_n10410_));
  AOI22X1  g10217(.A0(new_n8298_), .A1(new_n3208_), .B0(new_n4272_), .B1(new_n3462_), .Y(new_n10411_));
  AOI21X1  g10218(.A0(new_n3893_), .A1(new_n4992_), .B0(new_n10411_), .Y(new_n10412_));
  AND2X1   g10219(.A(\a[48] ), .B(\a[42] ), .Y(new_n10413_));
  INVX1    g10220(.A(new_n10413_), .Y(new_n10414_));
  OAI22X1  g10221(.A0(new_n8299_), .A1(new_n3212_), .B0(new_n8297_), .B1(new_n6502_), .Y(new_n10415_));
  AOI21X1  g10222(.A0(new_n3893_), .A1(new_n4992_), .B0(new_n10415_), .Y(new_n10416_));
  INVX1    g10223(.A(new_n10416_), .Y(new_n10417_));
  AOI22X1  g10224(.A0(\a[47] ), .A1(\a[43] ), .B0(\a[46] ), .B1(\a[44] ), .Y(new_n10418_));
  OAI22X1  g10225(.A0(new_n10418_), .A1(new_n10417_), .B0(new_n10414_), .B1(new_n10412_), .Y(new_n10419_));
  INVX1    g10226(.A(new_n10419_), .Y(new_n10420_));
  XOR2X1   g10227(.A(new_n10420_), .B(new_n10410_), .Y(new_n10421_));
  XOR2X1   g10228(.A(new_n10421_), .B(new_n10393_), .Y(new_n10422_));
  XOR2X1   g10229(.A(new_n10422_), .B(new_n10384_), .Y(new_n10423_));
  AND2X1   g10230(.A(new_n10257_), .B(new_n10254_), .Y(new_n10424_));
  AOI21X1  g10231(.A0(new_n10267_), .A1(new_n10258_), .B0(new_n10424_), .Y(new_n10425_));
  NOR2X1   g10232(.A(new_n10184_), .B(new_n10167_), .Y(new_n10426_));
  AOI21X1  g10233(.A0(new_n10300_), .A1(new_n10299_), .B0(new_n10426_), .Y(new_n10427_));
  OAI22X1  g10234(.A0(new_n7653_), .A1(new_n7617_), .B0(new_n7651_), .B1(new_n6180_), .Y(new_n10428_));
  OAI21X1  g10235(.A0(new_n7652_), .A1(new_n7618_), .B0(new_n10428_), .Y(new_n10429_));
  AND2X1   g10236(.A(new_n4321_), .B(new_n4404_), .Y(new_n10430_));
  NOR2X1   g10237(.A(new_n10428_), .B(new_n10430_), .Y(new_n10431_));
  OAI22X1  g10238(.A0(new_n4983_), .A1(new_n3036_), .B0(new_n3915_), .B1(new_n3081_), .Y(new_n10432_));
  AOI22X1  g10239(.A0(new_n10432_), .A1(new_n10431_), .B0(new_n10429_), .B1(new_n5290_), .Y(new_n10433_));
  XOR2X1   g10240(.A(new_n10433_), .B(new_n10427_), .Y(new_n10434_));
  OR2X1    g10241(.A(new_n10194_), .B(new_n10177_), .Y(new_n10435_));
  OAI21X1  g10242(.A0(new_n10266_), .A1(new_n10259_), .B0(new_n10435_), .Y(new_n10436_));
  XOR2X1   g10243(.A(new_n10436_), .B(new_n10434_), .Y(new_n10437_));
  AOI22X1  g10244(.A0(new_n10317_), .A1(new_n10227_), .B0(new_n6428_), .B1(new_n1674_), .Y(new_n10438_));
  AND2X1   g10245(.A(new_n6121_), .B(new_n2671_), .Y(new_n10439_));
  AOI22X1  g10246(.A0(new_n6795_), .A1(new_n1787_), .B0(new_n6427_), .B1(new_n2075_), .Y(new_n10440_));
  AOI22X1  g10247(.A0(\a[59] ), .A1(\a[31] ), .B0(\a[58] ), .B1(\a[32] ), .Y(new_n10441_));
  AOI21X1  g10248(.A0(new_n6121_), .A1(new_n2671_), .B0(new_n10441_), .Y(new_n10442_));
  AND2X1   g10249(.A(\a[60] ), .B(\a[30] ), .Y(new_n10443_));
  OAI22X1  g10250(.A0(new_n10443_), .A1(new_n10442_), .B0(new_n10440_), .B1(new_n10439_), .Y(new_n10444_));
  INVX1    g10251(.A(new_n10444_), .Y(new_n10445_));
  NAND2X1  g10252(.A(new_n10445_), .B(new_n10438_), .Y(new_n10446_));
  OAI22X1  g10253(.A0(new_n7973_), .A1(new_n1673_), .B0(new_n7972_), .B1(new_n1672_), .Y(new_n10447_));
  OAI21X1  g10254(.A0(new_n6557_), .A1(new_n1675_), .B0(new_n10447_), .Y(new_n10448_));
  AOI21X1  g10255(.A0(new_n6556_), .A1(new_n1674_), .B0(new_n10447_), .Y(new_n10449_));
  OAI22X1  g10256(.A0(new_n6606_), .A1(new_n1431_), .B0(new_n6023_), .B1(new_n1803_), .Y(new_n10450_));
  AND2X1   g10257(.A(\a[63] ), .B(\a[27] ), .Y(new_n10451_));
  AOI22X1  g10258(.A0(new_n10451_), .A1(new_n10448_), .B0(new_n10450_), .B1(new_n10449_), .Y(new_n10452_));
  OR2X1    g10259(.A(new_n10445_), .B(new_n10438_), .Y(new_n10453_));
  AOI21X1  g10260(.A0(new_n10446_), .A1(new_n10453_), .B0(new_n10452_), .Y(new_n10454_));
  AND2X1   g10261(.A(new_n10453_), .B(new_n10452_), .Y(new_n10455_));
  AOI21X1  g10262(.A0(new_n10455_), .A1(new_n10446_), .B0(new_n10454_), .Y(new_n10456_));
  XOR2X1   g10263(.A(new_n10456_), .B(new_n10437_), .Y(new_n10457_));
  XOR2X1   g10264(.A(new_n10457_), .B(new_n10425_), .Y(new_n10458_));
  XOR2X1   g10265(.A(new_n10458_), .B(new_n10423_), .Y(new_n10459_));
  INVX1    g10266(.A(new_n10459_), .Y(new_n10460_));
  XOR2X1   g10267(.A(new_n10460_), .B(new_n10382_), .Y(new_n10461_));
  OAI21X1  g10268(.A0(new_n10343_), .A1(new_n10354_), .B0(new_n10461_), .Y(new_n10462_));
  NAND2X1  g10269(.A(new_n10346_), .B(new_n10245_), .Y(new_n10463_));
  NOR2X1   g10270(.A(new_n10346_), .B(new_n10245_), .Y(new_n10464_));
  OAI21X1  g10271(.A0(new_n10351_), .A1(new_n10464_), .B0(new_n10463_), .Y(new_n10465_));
  NOR3X1   g10272(.A(new_n10461_), .B(new_n10343_), .C(new_n10354_), .Y(new_n10466_));
  INVX1    g10273(.A(new_n10466_), .Y(new_n10467_));
  AOI21X1  g10274(.A0(new_n10462_), .A1(new_n10467_), .B0(new_n10465_), .Y(new_n10468_));
  AND2X1   g10275(.A(new_n10467_), .B(new_n10465_), .Y(new_n10469_));
  AOI21X1  g10276(.A0(new_n10469_), .A1(new_n10462_), .B0(new_n10468_), .Y(\asquared[91] ));
  INVX1    g10277(.A(new_n10462_), .Y(new_n10471_));
  AOI21X1  g10278(.A0(new_n10467_), .A1(new_n10465_), .B0(new_n10471_), .Y(new_n10472_));
  NOR2X1   g10279(.A(new_n10381_), .B(new_n10377_), .Y(new_n10473_));
  AOI21X1  g10280(.A0(new_n10460_), .A1(new_n10382_), .B0(new_n10473_), .Y(new_n10474_));
  XOR2X1   g10281(.A(new_n10449_), .B(new_n10407_), .Y(new_n10475_));
  OAI21X1  g10282(.A0(new_n6793_), .A1(new_n2672_), .B0(new_n10440_), .Y(new_n10476_));
  XOR2X1   g10283(.A(new_n10476_), .B(new_n10475_), .Y(new_n10477_));
  NOR2X1   g10284(.A(new_n10433_), .B(new_n10427_), .Y(new_n10478_));
  AOI21X1  g10285(.A0(new_n10436_), .A1(new_n10434_), .B0(new_n10478_), .Y(new_n10479_));
  XOR2X1   g10286(.A(new_n10479_), .B(new_n10477_), .Y(new_n10480_));
  AOI22X1  g10287(.A0(\a[51] ), .A1(\a[40] ), .B0(\a[50] ), .B1(\a[41] ), .Y(new_n10481_));
  AND2X1   g10288(.A(\a[63] ), .B(\a[28] ), .Y(new_n10482_));
  INVX1    g10289(.A(new_n10482_), .Y(new_n10483_));
  AND2X1   g10290(.A(new_n4484_), .B(new_n4404_), .Y(new_n10484_));
  NOR3X1   g10291(.A(new_n10483_), .B(new_n10484_), .C(new_n10481_), .Y(new_n10485_));
  NOR2X1   g10292(.A(new_n10485_), .B(new_n10484_), .Y(new_n10486_));
  INVX1    g10293(.A(new_n10486_), .Y(new_n10487_));
  OAI22X1  g10294(.A0(new_n10487_), .A1(new_n10481_), .B0(new_n10485_), .B1(new_n10483_), .Y(new_n10488_));
  AND2X1   g10295(.A(\a[56] ), .B(\a[35] ), .Y(new_n10489_));
  AOI22X1  g10296(.A0(\a[48] ), .A1(\a[43] ), .B0(\a[47] ), .B1(\a[44] ), .Y(new_n10490_));
  INVX1    g10297(.A(new_n10490_), .Y(new_n10491_));
  NAND4X1  g10298(.A(\a[48] ), .B(\a[47] ), .C(\a[44] ), .D(\a[43] ), .Y(new_n10492_));
  NAND3X1  g10299(.A(new_n10491_), .B(new_n10492_), .C(new_n10489_), .Y(new_n10493_));
  AOI22X1  g10300(.A0(new_n10491_), .A1(new_n10489_), .B0(new_n4272_), .B1(new_n4992_), .Y(new_n10494_));
  AOI22X1  g10301(.A0(new_n10494_), .A1(new_n10491_), .B0(new_n10493_), .B1(new_n10489_), .Y(new_n10495_));
  XOR2X1   g10302(.A(new_n10495_), .B(new_n10488_), .Y(new_n10496_));
  NAND3X1  g10303(.A(\a[62] ), .B(\a[46] ), .C(\a[29] ), .Y(new_n10497_));
  NOR3X1   g10304(.A(new_n10497_), .B(new_n3460_), .C(new_n3811_), .Y(new_n10498_));
  AND2X1   g10305(.A(new_n10497_), .B(new_n8873_), .Y(new_n10499_));
  OAI21X1  g10306(.A0(new_n6606_), .A1(new_n1803_), .B0(new_n3460_), .Y(new_n10500_));
  AOI21X1  g10307(.A0(new_n10500_), .A1(new_n10499_), .B0(new_n10498_), .Y(new_n10501_));
  XOR2X1   g10308(.A(new_n10501_), .B(new_n10496_), .Y(new_n10502_));
  XOR2X1   g10309(.A(new_n10502_), .B(new_n10480_), .Y(new_n10503_));
  OR2X1    g10310(.A(new_n10373_), .B(new_n10360_), .Y(new_n10504_));
  OAI21X1  g10311(.A0(new_n10375_), .A1(new_n10356_), .B0(new_n10504_), .Y(new_n10505_));
  XOR2X1   g10312(.A(new_n10505_), .B(new_n10503_), .Y(new_n10506_));
  AND2X1   g10313(.A(new_n10362_), .B(new_n10305_), .Y(new_n10507_));
  AOI21X1  g10314(.A0(new_n10363_), .A1(new_n10283_), .B0(new_n10507_), .Y(new_n10508_));
  AOI22X1  g10315(.A0(\a[57] ), .A1(\a[34] ), .B0(\a[55] ), .B1(\a[36] ), .Y(new_n10509_));
  INVX1    g10316(.A(new_n10509_), .Y(new_n10510_));
  NAND4X1  g10317(.A(\a[57] ), .B(\a[55] ), .C(\a[36] ), .D(\a[34] ), .Y(new_n10511_));
  NAND3X1  g10318(.A(new_n10510_), .B(new_n10511_), .C(new_n5399_), .Y(new_n10512_));
  AOI22X1  g10319(.A0(new_n10510_), .A1(new_n5399_), .B0(new_n9461_), .B1(new_n4695_), .Y(new_n10513_));
  AOI22X1  g10320(.A0(new_n10513_), .A1(new_n10510_), .B0(new_n10512_), .B1(new_n5399_), .Y(new_n10514_));
  XOR2X1   g10321(.A(new_n10514_), .B(new_n10508_), .Y(new_n10515_));
  NOR2X1   g10322(.A(new_n10295_), .B(new_n10288_), .Y(new_n10516_));
  AOI21X1  g10323(.A0(new_n10386_), .A1(new_n10385_), .B0(new_n10516_), .Y(new_n10517_));
  XOR2X1   g10324(.A(new_n10517_), .B(new_n10515_), .Y(new_n10518_));
  AND2X1   g10325(.A(new_n10370_), .B(new_n10367_), .Y(new_n10519_));
  AOI21X1  g10326(.A0(new_n10371_), .A1(new_n10364_), .B0(new_n10519_), .Y(new_n10520_));
  OAI22X1  g10327(.A0(new_n6796_), .A1(new_n2673_), .B0(new_n6794_), .B1(new_n2672_), .Y(new_n10521_));
  OAI21X1  g10328(.A0(new_n6793_), .A1(new_n2675_), .B0(new_n10521_), .Y(new_n10522_));
  AOI21X1  g10329(.A0(new_n6121_), .A1(new_n2674_), .B0(new_n10521_), .Y(new_n10523_));
  OAI22X1  g10330(.A0(new_n5617_), .A1(new_n2219_), .B0(new_n5379_), .B1(new_n1851_), .Y(new_n10524_));
  AND2X1   g10331(.A(\a[60] ), .B(\a[31] ), .Y(new_n10525_));
  AOI22X1  g10332(.A0(new_n10525_), .A1(new_n10522_), .B0(new_n10524_), .B1(new_n10523_), .Y(new_n10526_));
  NAND4X1  g10333(.A(\a[54] ), .B(\a[52] ), .C(\a[39] ), .D(\a[37] ), .Y(new_n10527_));
  NAND4X1  g10334(.A(\a[54] ), .B(\a[53] ), .C(\a[38] ), .D(\a[37] ), .Y(new_n10528_));
  AOI22X1  g10335(.A0(new_n10528_), .A1(new_n10527_), .B0(new_n5048_), .B1(new_n3503_), .Y(new_n10529_));
  NAND2X1  g10336(.A(\a[54] ), .B(\a[37] ), .Y(new_n10530_));
  NAND4X1  g10337(.A(\a[53] ), .B(\a[52] ), .C(\a[39] ), .D(\a[38] ), .Y(new_n10531_));
  NAND3X1  g10338(.A(new_n10528_), .B(new_n10527_), .C(new_n10531_), .Y(new_n10532_));
  AOI22X1  g10339(.A0(\a[53] ), .A1(\a[38] ), .B0(\a[52] ), .B1(\a[39] ), .Y(new_n10533_));
  OAI22X1  g10340(.A0(new_n10533_), .A1(new_n10532_), .B0(new_n10530_), .B1(new_n10529_), .Y(new_n10534_));
  XOR2X1   g10341(.A(new_n10534_), .B(new_n10431_), .Y(new_n10535_));
  XOR2X1   g10342(.A(new_n10535_), .B(new_n10526_), .Y(new_n10536_));
  XOR2X1   g10343(.A(new_n10536_), .B(new_n10520_), .Y(new_n10537_));
  XOR2X1   g10344(.A(new_n10537_), .B(new_n10518_), .Y(new_n10538_));
  XOR2X1   g10345(.A(new_n10538_), .B(new_n10506_), .Y(new_n10539_));
  AND2X1   g10346(.A(new_n10422_), .B(new_n10384_), .Y(new_n10540_));
  INVX1    g10347(.A(new_n10540_), .Y(new_n10541_));
  INVX1    g10348(.A(new_n10423_), .Y(new_n10542_));
  OAI21X1  g10349(.A0(new_n10458_), .A1(new_n10542_), .B0(new_n10541_), .Y(new_n10543_));
  INVX1    g10350(.A(new_n10543_), .Y(new_n10544_));
  NAND2X1  g10351(.A(new_n10456_), .B(new_n10437_), .Y(new_n10545_));
  INVX1    g10352(.A(new_n10457_), .Y(new_n10546_));
  OAI21X1  g10353(.A0(new_n10546_), .A1(new_n10425_), .B0(new_n10545_), .Y(new_n10547_));
  NAND2X1  g10354(.A(new_n10391_), .B(new_n10387_), .Y(new_n10548_));
  OAI21X1  g10355(.A0(new_n10421_), .A1(new_n10393_), .B0(new_n10548_), .Y(new_n10549_));
  AND2X1   g10356(.A(\a[61] ), .B(\a[30] ), .Y(new_n10550_));
  INVX1    g10357(.A(new_n10550_), .Y(new_n10551_));
  XOR2X1   g10358(.A(new_n10551_), .B(new_n10416_), .Y(new_n10552_));
  XOR2X1   g10359(.A(new_n10552_), .B(new_n10399_), .Y(new_n10553_));
  INVX1    g10360(.A(new_n10553_), .Y(new_n10554_));
  AND2X1   g10361(.A(new_n10409_), .B(new_n10401_), .Y(new_n10555_));
  AND2X1   g10362(.A(new_n10419_), .B(new_n10410_), .Y(new_n10556_));
  NOR2X1   g10363(.A(new_n10444_), .B(new_n10438_), .Y(new_n10557_));
  OR4X1    g10364(.A(new_n10454_), .B(new_n10557_), .C(new_n10556_), .D(new_n10555_), .Y(new_n10558_));
  OAI22X1  g10365(.A0(new_n10454_), .A1(new_n10557_), .B0(new_n10556_), .B1(new_n10555_), .Y(new_n10559_));
  NAND2X1  g10366(.A(new_n10559_), .B(new_n10558_), .Y(new_n10560_));
  XOR2X1   g10367(.A(new_n10560_), .B(new_n10554_), .Y(new_n10561_));
  XOR2X1   g10368(.A(new_n10561_), .B(new_n10549_), .Y(new_n10562_));
  XOR2X1   g10369(.A(new_n10562_), .B(new_n10547_), .Y(new_n10563_));
  XOR2X1   g10370(.A(new_n10563_), .B(new_n10544_), .Y(new_n10564_));
  XOR2X1   g10371(.A(new_n10564_), .B(new_n10539_), .Y(new_n10565_));
  NOR2X1   g10372(.A(new_n10565_), .B(new_n10474_), .Y(new_n10566_));
  AND2X1   g10373(.A(new_n10565_), .B(new_n10474_), .Y(new_n10567_));
  OR2X1    g10374(.A(new_n10567_), .B(new_n10566_), .Y(new_n10568_));
  XOR2X1   g10375(.A(new_n10568_), .B(new_n10472_), .Y(\asquared[92] ));
  AND2X1   g10376(.A(new_n10561_), .B(new_n10549_), .Y(new_n10570_));
  AOI21X1  g10377(.A0(new_n10562_), .A1(new_n10547_), .B0(new_n10570_), .Y(new_n10571_));
  INVX1    g10378(.A(new_n10520_), .Y(new_n10572_));
  AND2X1   g10379(.A(new_n10536_), .B(new_n10572_), .Y(new_n10573_));
  NOR2X1   g10380(.A(new_n10537_), .B(new_n10518_), .Y(new_n10574_));
  NOR2X1   g10381(.A(new_n10574_), .B(new_n10573_), .Y(new_n10575_));
  OAI21X1  g10382(.A0(new_n10560_), .A1(new_n10554_), .B0(new_n10559_), .Y(new_n10576_));
  AND2X1   g10383(.A(\a[61] ), .B(\a[31] ), .Y(new_n10577_));
  AND2X1   g10384(.A(\a[62] ), .B(\a[30] ), .Y(new_n10578_));
  OAI22X1  g10385(.A0(new_n10578_), .A1(new_n10577_), .B0(new_n6557_), .B1(new_n2076_), .Y(new_n10579_));
  XOR2X1   g10386(.A(new_n10579_), .B(new_n10499_), .Y(new_n10580_));
  AOI22X1  g10387(.A0(new_n5048_), .A1(new_n4077_), .B0(new_n4904_), .B1(new_n2847_), .Y(new_n10581_));
  AOI21X1  g10388(.A0(new_n7164_), .A1(new_n4404_), .B0(new_n10581_), .Y(new_n10582_));
  NAND2X1  g10389(.A(\a[53] ), .B(\a[39] ), .Y(new_n10583_));
  AOI22X1  g10390(.A0(\a[52] ), .A1(\a[40] ), .B0(\a[51] ), .B1(\a[41] ), .Y(new_n10584_));
  AOI21X1  g10391(.A0(new_n7164_), .A1(new_n4404_), .B0(new_n10582_), .Y(new_n10585_));
  INVX1    g10392(.A(new_n10585_), .Y(new_n10586_));
  OAI22X1  g10393(.A0(new_n10586_), .A1(new_n10584_), .B0(new_n10583_), .B1(new_n10582_), .Y(new_n10587_));
  XOR2X1   g10394(.A(new_n10587_), .B(new_n10580_), .Y(new_n10588_));
  NAND2X1  g10395(.A(new_n10552_), .B(new_n10399_), .Y(new_n10589_));
  OAI21X1  g10396(.A0(new_n10551_), .A1(new_n10416_), .B0(new_n10589_), .Y(new_n10590_));
  XOR2X1   g10397(.A(new_n10590_), .B(new_n10588_), .Y(new_n10591_));
  NAND2X1  g10398(.A(\a[58] ), .B(\a[34] ), .Y(new_n10592_));
  NOR4X1   g10399(.A(new_n5441_), .B(new_n4983_), .C(new_n3096_), .D(new_n2557_), .Y(new_n10593_));
  NAND4X1  g10400(.A(\a[58] ), .B(\a[50] ), .C(\a[42] ), .D(\a[34] ), .Y(new_n10594_));
  NAND4X1  g10401(.A(\a[58] ), .B(\a[57] ), .C(\a[35] ), .D(\a[34] ), .Y(new_n10595_));
  AOI21X1  g10402(.A0(new_n10595_), .A1(new_n10594_), .B0(new_n10593_), .Y(new_n10596_));
  OR2X1    g10403(.A(new_n10596_), .B(new_n10593_), .Y(new_n10597_));
  AOI22X1  g10404(.A0(\a[57] ), .A1(\a[35] ), .B0(\a[50] ), .B1(\a[42] ), .Y(new_n10598_));
  OAI22X1  g10405(.A0(new_n10598_), .A1(new_n10597_), .B0(new_n10596_), .B1(new_n10592_), .Y(new_n10599_));
  NAND4X1  g10406(.A(\a[49] ), .B(\a[47] ), .C(\a[45] ), .D(\a[43] ), .Y(new_n10600_));
  NAND4X1  g10407(.A(\a[49] ), .B(\a[48] ), .C(\a[44] ), .D(\a[43] ), .Y(new_n10601_));
  AOI22X1  g10408(.A0(new_n10601_), .A1(new_n10600_), .B0(new_n4272_), .B1(new_n3918_), .Y(new_n10602_));
  NAND2X1  g10409(.A(\a[49] ), .B(\a[43] ), .Y(new_n10603_));
  NAND4X1  g10410(.A(\a[48] ), .B(\a[47] ), .C(\a[45] ), .D(\a[44] ), .Y(new_n10604_));
  NAND3X1  g10411(.A(new_n10601_), .B(new_n10600_), .C(new_n10604_), .Y(new_n10605_));
  AOI22X1  g10412(.A0(\a[48] ), .A1(\a[44] ), .B0(\a[47] ), .B1(\a[45] ), .Y(new_n10606_));
  OAI22X1  g10413(.A0(new_n10606_), .A1(new_n10605_), .B0(new_n10603_), .B1(new_n10602_), .Y(new_n10607_));
  XOR2X1   g10414(.A(new_n10607_), .B(new_n10599_), .Y(new_n10608_));
  AND2X1   g10415(.A(\a[56] ), .B(\a[36] ), .Y(new_n10609_));
  INVX1    g10416(.A(new_n10609_), .Y(new_n10610_));
  AOI22X1  g10417(.A0(\a[63] ), .A1(\a[29] ), .B0(\a[59] ), .B1(\a[33] ), .Y(new_n10611_));
  NOR4X1   g10418(.A(new_n6549_), .B(new_n5617_), .C(new_n1851_), .D(new_n1803_), .Y(new_n10612_));
  NOR3X1   g10419(.A(new_n10611_), .B(new_n10612_), .C(new_n10610_), .Y(new_n10613_));
  OR2X1    g10420(.A(new_n10613_), .B(new_n10612_), .Y(new_n10614_));
  OAI22X1  g10421(.A0(new_n10614_), .A1(new_n10611_), .B0(new_n10613_), .B1(new_n10610_), .Y(new_n10615_));
  XOR2X1   g10422(.A(new_n10615_), .B(new_n10608_), .Y(new_n10616_));
  XOR2X1   g10423(.A(new_n10616_), .B(new_n10591_), .Y(new_n10617_));
  XOR2X1   g10424(.A(new_n10617_), .B(new_n10576_), .Y(new_n10618_));
  XOR2X1   g10425(.A(new_n10618_), .B(new_n10575_), .Y(new_n10619_));
  XOR2X1   g10426(.A(new_n10619_), .B(new_n10571_), .Y(new_n10620_));
  AND2X1   g10427(.A(new_n10505_), .B(new_n10503_), .Y(new_n10621_));
  AND2X1   g10428(.A(new_n10538_), .B(new_n10506_), .Y(new_n10622_));
  OR2X1    g10429(.A(new_n10622_), .B(new_n10621_), .Y(new_n10623_));
  OAI21X1  g10430(.A0(new_n10428_), .A1(new_n10430_), .B0(new_n10534_), .Y(new_n10624_));
  OAI21X1  g10431(.A0(new_n10535_), .A1(new_n10526_), .B0(new_n10624_), .Y(new_n10625_));
  INVX1    g10432(.A(new_n10625_), .Y(new_n10626_));
  NAND4X1  g10433(.A(new_n10449_), .B(new_n10403_), .C(new_n10402_), .D(new_n10406_), .Y(new_n10627_));
  AOI21X1  g10434(.A0(new_n5048_), .A1(new_n3164_), .B0(new_n10404_), .Y(new_n10628_));
  NOR2X1   g10435(.A(new_n10449_), .B(new_n10628_), .Y(new_n10629_));
  AOI21X1  g10436(.A0(new_n10476_), .A1(new_n10627_), .B0(new_n10629_), .Y(new_n10630_));
  XOR2X1   g10437(.A(new_n10630_), .B(new_n10626_), .Y(new_n10631_));
  INVX1    g10438(.A(new_n10488_), .Y(new_n10632_));
  OR2X1    g10439(.A(new_n10495_), .B(new_n10632_), .Y(new_n10633_));
  OR2X1    g10440(.A(new_n10501_), .B(new_n10496_), .Y(new_n10634_));
  AND2X1   g10441(.A(new_n10634_), .B(new_n10633_), .Y(new_n10635_));
  XOR2X1   g10442(.A(new_n10635_), .B(new_n10631_), .Y(new_n10636_));
  NOR2X1   g10443(.A(new_n10479_), .B(new_n10477_), .Y(new_n10637_));
  AOI21X1  g10444(.A0(new_n10502_), .A1(new_n10480_), .B0(new_n10637_), .Y(new_n10638_));
  OR2X1    g10445(.A(new_n10514_), .B(new_n10508_), .Y(new_n10639_));
  INVX1    g10446(.A(new_n10515_), .Y(new_n10640_));
  OAI21X1  g10447(.A0(new_n10517_), .A1(new_n10640_), .B0(new_n10639_), .Y(new_n10641_));
  INVX1    g10448(.A(new_n10523_), .Y(new_n10642_));
  XOR2X1   g10449(.A(new_n10532_), .B(new_n10642_), .Y(new_n10643_));
  XOR2X1   g10450(.A(new_n10643_), .B(new_n10487_), .Y(new_n10644_));
  INVX1    g10451(.A(new_n10644_), .Y(new_n10645_));
  XOR2X1   g10452(.A(new_n10513_), .B(new_n10494_), .Y(new_n10646_));
  AND2X1   g10453(.A(\a[60] ), .B(\a[32] ), .Y(new_n10647_));
  AOI22X1  g10454(.A0(\a[55] ), .A1(\a[37] ), .B0(\a[54] ), .B1(\a[38] ), .Y(new_n10648_));
  INVX1    g10455(.A(new_n10648_), .Y(new_n10649_));
  NAND4X1  g10456(.A(\a[55] ), .B(\a[54] ), .C(\a[38] ), .D(\a[37] ), .Y(new_n10650_));
  NAND3X1  g10457(.A(new_n10650_), .B(new_n10649_), .C(new_n10647_), .Y(new_n10651_));
  AOI22X1  g10458(.A0(new_n10649_), .A1(new_n10647_), .B0(new_n5240_), .B1(new_n3164_), .Y(new_n10652_));
  AOI22X1  g10459(.A0(new_n10652_), .A1(new_n10649_), .B0(new_n10651_), .B1(new_n10647_), .Y(new_n10653_));
  XOR2X1   g10460(.A(new_n10653_), .B(new_n10646_), .Y(new_n10654_));
  XOR2X1   g10461(.A(new_n10654_), .B(new_n10645_), .Y(new_n10655_));
  XOR2X1   g10462(.A(new_n10655_), .B(new_n10641_), .Y(new_n10656_));
  XOR2X1   g10463(.A(new_n10656_), .B(new_n10638_), .Y(new_n10657_));
  XOR2X1   g10464(.A(new_n10657_), .B(new_n10636_), .Y(new_n10658_));
  XOR2X1   g10465(.A(new_n10658_), .B(new_n10623_), .Y(new_n10659_));
  XOR2X1   g10466(.A(new_n10659_), .B(new_n10620_), .Y(new_n10660_));
  INVX1    g10467(.A(new_n10539_), .Y(new_n10661_));
  NAND2X1  g10468(.A(new_n10563_), .B(new_n10543_), .Y(new_n10662_));
  OAI21X1  g10469(.A0(new_n10564_), .A1(new_n10661_), .B0(new_n10662_), .Y(new_n10663_));
  AND2X1   g10470(.A(new_n10663_), .B(new_n10660_), .Y(new_n10664_));
  INVX1    g10471(.A(new_n10664_), .Y(new_n10665_));
  INVX1    g10472(.A(new_n10566_), .Y(new_n10666_));
  OAI21X1  g10473(.A0(new_n10567_), .A1(new_n10472_), .B0(new_n10666_), .Y(new_n10667_));
  NOR2X1   g10474(.A(new_n10663_), .B(new_n10660_), .Y(new_n10668_));
  INVX1    g10475(.A(new_n10668_), .Y(new_n10669_));
  AOI21X1  g10476(.A0(new_n10665_), .A1(new_n10669_), .B0(new_n10667_), .Y(new_n10670_));
  AND2X1   g10477(.A(new_n10669_), .B(new_n10667_), .Y(new_n10671_));
  AOI21X1  g10478(.A0(new_n10671_), .A1(new_n10665_), .B0(new_n10670_), .Y(\asquared[93] ));
  AOI21X1  g10479(.A0(new_n10669_), .A1(new_n10667_), .B0(new_n10664_), .Y(new_n10673_));
  AND2X1   g10480(.A(new_n10658_), .B(new_n10623_), .Y(new_n10674_));
  AND2X1   g10481(.A(new_n10659_), .B(new_n10620_), .Y(new_n10675_));
  OR2X1    g10482(.A(new_n10675_), .B(new_n10674_), .Y(new_n10676_));
  OAI21X1  g10483(.A0(new_n10574_), .A1(new_n10573_), .B0(new_n10618_), .Y(new_n10677_));
  OAI21X1  g10484(.A0(new_n10619_), .A1(new_n10571_), .B0(new_n10677_), .Y(new_n10678_));
  AND2X1   g10485(.A(new_n10513_), .B(new_n10494_), .Y(new_n10679_));
  OR2X1    g10486(.A(new_n10513_), .B(new_n10494_), .Y(new_n10680_));
  OAI21X1  g10487(.A0(new_n10653_), .A1(new_n10679_), .B0(new_n10680_), .Y(new_n10681_));
  INVX1    g10488(.A(new_n10681_), .Y(new_n10682_));
  AND2X1   g10489(.A(new_n10532_), .B(new_n10642_), .Y(new_n10683_));
  AOI21X1  g10490(.A0(new_n10643_), .A1(new_n10487_), .B0(new_n10683_), .Y(new_n10684_));
  XOR2X1   g10491(.A(new_n10684_), .B(new_n10682_), .Y(new_n10685_));
  AND2X1   g10492(.A(new_n10607_), .B(new_n10599_), .Y(new_n10686_));
  AOI21X1  g10493(.A0(new_n10615_), .A1(new_n10608_), .B0(new_n10686_), .Y(new_n10687_));
  XOR2X1   g10494(.A(new_n10687_), .B(new_n10685_), .Y(new_n10688_));
  NOR2X1   g10495(.A(new_n10654_), .B(new_n10645_), .Y(new_n10689_));
  AOI21X1  g10496(.A0(new_n10655_), .A1(new_n10641_), .B0(new_n10689_), .Y(new_n10690_));
  XOR2X1   g10497(.A(new_n10690_), .B(new_n10688_), .Y(new_n10691_));
  AND2X1   g10498(.A(new_n10587_), .B(new_n10580_), .Y(new_n10692_));
  AOI21X1  g10499(.A0(new_n10590_), .A1(new_n10588_), .B0(new_n10692_), .Y(new_n10693_));
  XOR2X1   g10500(.A(new_n10605_), .B(new_n10597_), .Y(new_n10694_));
  XOR2X1   g10501(.A(new_n10694_), .B(new_n10585_), .Y(new_n10695_));
  INVX1    g10502(.A(new_n10652_), .Y(new_n10696_));
  XOR2X1   g10503(.A(new_n10696_), .B(new_n10614_), .Y(new_n10697_));
  OAI22X1  g10504(.A0(new_n10579_), .A1(new_n10499_), .B0(new_n6557_), .B1(new_n2076_), .Y(new_n10698_));
  XOR2X1   g10505(.A(new_n10698_), .B(new_n10697_), .Y(new_n10699_));
  XOR2X1   g10506(.A(new_n10699_), .B(new_n10695_), .Y(new_n10700_));
  XOR2X1   g10507(.A(new_n10700_), .B(new_n10693_), .Y(new_n10701_));
  XOR2X1   g10508(.A(new_n10701_), .B(new_n10691_), .Y(new_n10702_));
  XOR2X1   g10509(.A(new_n10702_), .B(new_n10678_), .Y(new_n10703_));
  INVX1    g10510(.A(new_n10656_), .Y(new_n10704_));
  OR2X1    g10511(.A(new_n10657_), .B(new_n10636_), .Y(new_n10705_));
  OAI21X1  g10512(.A0(new_n10704_), .A1(new_n10638_), .B0(new_n10705_), .Y(new_n10706_));
  AND2X1   g10513(.A(new_n10616_), .B(new_n10591_), .Y(new_n10707_));
  AOI21X1  g10514(.A0(new_n10617_), .A1(new_n10576_), .B0(new_n10707_), .Y(new_n10708_));
  NOR2X1   g10515(.A(new_n10630_), .B(new_n10626_), .Y(new_n10709_));
  INVX1    g10516(.A(new_n10635_), .Y(new_n10710_));
  AOI21X1  g10517(.A0(new_n10710_), .A1(new_n10631_), .B0(new_n10709_), .Y(new_n10711_));
  NAND4X1  g10518(.A(\a[63] ), .B(\a[60] ), .C(\a[33] ), .D(\a[30] ), .Y(new_n10712_));
  NAND4X1  g10519(.A(\a[63] ), .B(\a[61] ), .C(\a[32] ), .D(\a[30] ), .Y(new_n10713_));
  AOI22X1  g10520(.A0(new_n10713_), .A1(new_n10712_), .B0(new_n6428_), .B1(new_n2674_), .Y(new_n10714_));
  NAND4X1  g10521(.A(\a[61] ), .B(\a[60] ), .C(\a[33] ), .D(\a[32] ), .Y(new_n10715_));
  NAND3X1  g10522(.A(new_n10713_), .B(new_n10712_), .C(new_n10715_), .Y(new_n10716_));
  AOI22X1  g10523(.A0(\a[61] ), .A1(\a[32] ), .B0(\a[60] ), .B1(\a[33] ), .Y(new_n10717_));
  NAND2X1  g10524(.A(\a[63] ), .B(\a[30] ), .Y(new_n10718_));
  OAI22X1  g10525(.A0(new_n10718_), .A1(new_n10714_), .B0(new_n10717_), .B1(new_n10716_), .Y(new_n10719_));
  INVX1    g10526(.A(new_n10102_), .Y(new_n10720_));
  NAND4X1  g10527(.A(\a[57] ), .B(\a[54] ), .C(\a[39] ), .D(\a[36] ), .Y(new_n10721_));
  NAND4X1  g10528(.A(\a[58] ), .B(\a[57] ), .C(\a[36] ), .D(\a[35] ), .Y(new_n10722_));
  NAND4X1  g10529(.A(\a[58] ), .B(\a[54] ), .C(\a[39] ), .D(\a[35] ), .Y(new_n10723_));
  NAND2X1  g10530(.A(new_n10723_), .B(new_n10722_), .Y(new_n10724_));
  AND2X1   g10531(.A(new_n10724_), .B(new_n10721_), .Y(new_n10725_));
  NAND3X1  g10532(.A(new_n10723_), .B(new_n10722_), .C(new_n10721_), .Y(new_n10726_));
  AOI22X1  g10533(.A0(\a[57] ), .A1(\a[36] ), .B0(\a[54] ), .B1(\a[39] ), .Y(new_n10727_));
  OAI22X1  g10534(.A0(new_n10727_), .A1(new_n10726_), .B0(new_n10725_), .B1(new_n10720_), .Y(new_n10728_));
  XOR2X1   g10535(.A(new_n10728_), .B(new_n10719_), .Y(new_n10729_));
  AND2X1   g10536(.A(\a[59] ), .B(\a[34] ), .Y(new_n10730_));
  INVX1    g10537(.A(new_n10730_), .Y(new_n10731_));
  AOI22X1  g10538(.A0(\a[53] ), .A1(\a[40] ), .B0(\a[52] ), .B1(\a[41] ), .Y(new_n10732_));
  AND2X1   g10539(.A(new_n5048_), .B(new_n4404_), .Y(new_n10733_));
  NOR3X1   g10540(.A(new_n10732_), .B(new_n10733_), .C(new_n10731_), .Y(new_n10734_));
  NOR2X1   g10541(.A(new_n10734_), .B(new_n10733_), .Y(new_n10735_));
  INVX1    g10542(.A(new_n10735_), .Y(new_n10736_));
  OAI22X1  g10543(.A0(new_n10736_), .A1(new_n10732_), .B0(new_n10734_), .B1(new_n10731_), .Y(new_n10737_));
  XOR2X1   g10544(.A(new_n10737_), .B(new_n10729_), .Y(new_n10738_));
  INVX1    g10545(.A(new_n10738_), .Y(new_n10739_));
  AOI22X1  g10546(.A0(\a[55] ), .A1(\a[38] ), .B0(\a[48] ), .B1(\a[45] ), .Y(new_n10740_));
  NOR4X1   g10547(.A(new_n4906_), .B(new_n3926_), .C(new_n3811_), .D(new_n2519_), .Y(new_n10741_));
  NOR4X1   g10548(.A(new_n6022_), .B(new_n3926_), .C(new_n3811_), .D(new_n2345_), .Y(new_n10742_));
  AOI21X1  g10549(.A0(new_n6237_), .A1(new_n3164_), .B0(new_n10742_), .Y(new_n10743_));
  NOR2X1   g10550(.A(new_n10743_), .B(new_n10741_), .Y(new_n10744_));
  INVX1    g10551(.A(new_n10741_), .Y(new_n10745_));
  AND2X1   g10552(.A(new_n10743_), .B(new_n10745_), .Y(new_n10746_));
  INVX1    g10553(.A(new_n10746_), .Y(new_n10747_));
  NAND2X1  g10554(.A(\a[56] ), .B(\a[37] ), .Y(new_n10748_));
  OAI22X1  g10555(.A0(new_n10748_), .A1(new_n10744_), .B0(new_n10747_), .B1(new_n10740_), .Y(new_n10749_));
  NAND4X1  g10556(.A(\a[51] ), .B(\a[49] ), .C(\a[44] ), .D(\a[42] ), .Y(new_n10750_));
  NAND4X1  g10557(.A(\a[51] ), .B(\a[50] ), .C(\a[43] ), .D(\a[42] ), .Y(new_n10751_));
  AOI22X1  g10558(.A0(new_n10751_), .A1(new_n10750_), .B0(new_n4321_), .B1(new_n4992_), .Y(new_n10752_));
  NAND2X1  g10559(.A(\a[51] ), .B(\a[42] ), .Y(new_n10753_));
  AOI21X1  g10560(.A0(new_n4321_), .A1(new_n4992_), .B0(new_n10752_), .Y(new_n10754_));
  INVX1    g10561(.A(new_n10754_), .Y(new_n10755_));
  AOI22X1  g10562(.A0(\a[50] ), .A1(\a[43] ), .B0(\a[49] ), .B1(\a[44] ), .Y(new_n10756_));
  OAI22X1  g10563(.A0(new_n10756_), .A1(new_n10755_), .B0(new_n10753_), .B1(new_n10752_), .Y(new_n10757_));
  XOR2X1   g10564(.A(new_n10757_), .B(new_n10749_), .Y(new_n10758_));
  AND2X1   g10565(.A(\a[62] ), .B(\a[47] ), .Y(new_n10759_));
  AOI21X1  g10566(.A0(new_n10759_), .A1(\a[31] ), .B0(new_n8296_), .Y(new_n10760_));
  AOI21X1  g10567(.A0(new_n10759_), .A1(\a[31] ), .B0(new_n3893_), .Y(new_n10761_));
  INVX1    g10568(.A(new_n10761_), .Y(new_n10762_));
  AOI21X1  g10569(.A0(\a[62] ), .A1(\a[31] ), .B0(\a[47] ), .Y(new_n10763_));
  OAI22X1  g10570(.A0(new_n10763_), .A1(new_n10762_), .B0(new_n10760_), .B1(new_n8296_), .Y(new_n10764_));
  INVX1    g10571(.A(new_n10764_), .Y(new_n10765_));
  XOR2X1   g10572(.A(new_n10765_), .B(new_n10758_), .Y(new_n10766_));
  XOR2X1   g10573(.A(new_n10766_), .B(new_n10739_), .Y(new_n10767_));
  XOR2X1   g10574(.A(new_n10767_), .B(new_n10711_), .Y(new_n10768_));
  XOR2X1   g10575(.A(new_n10768_), .B(new_n10708_), .Y(new_n10769_));
  XOR2X1   g10576(.A(new_n10769_), .B(new_n10706_), .Y(new_n10770_));
  XOR2X1   g10577(.A(new_n10770_), .B(new_n10703_), .Y(new_n10771_));
  AND2X1   g10578(.A(new_n10771_), .B(new_n10676_), .Y(new_n10772_));
  NOR3X1   g10579(.A(new_n10771_), .B(new_n10675_), .C(new_n10674_), .Y(new_n10773_));
  OR2X1    g10580(.A(new_n10773_), .B(new_n10772_), .Y(new_n10774_));
  XOR2X1   g10581(.A(new_n10774_), .B(new_n10673_), .Y(\asquared[94] ));
  NOR2X1   g10582(.A(new_n10768_), .B(new_n10708_), .Y(new_n10776_));
  AOI21X1  g10583(.A0(new_n10769_), .A1(new_n10706_), .B0(new_n10776_), .Y(new_n10777_));
  AND2X1   g10584(.A(new_n10766_), .B(new_n10739_), .Y(new_n10778_));
  OR2X1    g10585(.A(new_n10766_), .B(new_n10739_), .Y(new_n10779_));
  OAI21X1  g10586(.A0(new_n10778_), .A1(new_n10711_), .B0(new_n10779_), .Y(new_n10780_));
  AND2X1   g10587(.A(new_n10696_), .B(new_n10614_), .Y(new_n10781_));
  AOI21X1  g10588(.A0(new_n10698_), .A1(new_n10697_), .B0(new_n10781_), .Y(new_n10782_));
  AND2X1   g10589(.A(new_n10605_), .B(new_n10597_), .Y(new_n10783_));
  AOI21X1  g10590(.A0(new_n10694_), .A1(new_n10586_), .B0(new_n10783_), .Y(new_n10784_));
  XOR2X1   g10591(.A(new_n10784_), .B(new_n10782_), .Y(new_n10785_));
  AND2X1   g10592(.A(new_n10728_), .B(new_n10719_), .Y(new_n10786_));
  AOI21X1  g10593(.A0(new_n10737_), .A1(new_n10729_), .B0(new_n10786_), .Y(new_n10787_));
  XOR2X1   g10594(.A(new_n10787_), .B(new_n10785_), .Y(new_n10788_));
  XOR2X1   g10595(.A(new_n10694_), .B(new_n10586_), .Y(new_n10789_));
  NOR2X1   g10596(.A(new_n10700_), .B(new_n10693_), .Y(new_n10790_));
  AOI21X1  g10597(.A0(new_n10699_), .A1(new_n10789_), .B0(new_n10790_), .Y(new_n10791_));
  XOR2X1   g10598(.A(new_n10791_), .B(new_n10788_), .Y(new_n10792_));
  INVX1    g10599(.A(new_n10792_), .Y(new_n10793_));
  XOR2X1   g10600(.A(new_n10793_), .B(new_n10780_), .Y(new_n10794_));
  XOR2X1   g10601(.A(new_n10794_), .B(new_n10777_), .Y(new_n10795_));
  NOR2X1   g10602(.A(new_n10690_), .B(new_n10688_), .Y(new_n10796_));
  AOI21X1  g10603(.A0(new_n10701_), .A1(new_n10691_), .B0(new_n10796_), .Y(new_n10797_));
  INVX1    g10604(.A(new_n10797_), .Y(new_n10798_));
  XOR2X1   g10605(.A(new_n10762_), .B(new_n8766_), .Y(new_n10799_));
  XOR2X1   g10606(.A(new_n10799_), .B(new_n10746_), .Y(new_n10800_));
  AND2X1   g10607(.A(new_n10757_), .B(new_n10749_), .Y(new_n10801_));
  AOI21X1  g10608(.A0(new_n10764_), .A1(new_n10758_), .B0(new_n10801_), .Y(new_n10802_));
  XOR2X1   g10609(.A(new_n10802_), .B(new_n10800_), .Y(new_n10803_));
  XOR2X1   g10610(.A(new_n10726_), .B(new_n10716_), .Y(new_n10804_));
  XOR2X1   g10611(.A(new_n10804_), .B(new_n10736_), .Y(new_n10805_));
  XOR2X1   g10612(.A(new_n10805_), .B(new_n10803_), .Y(new_n10806_));
  XOR2X1   g10613(.A(new_n10806_), .B(new_n10798_), .Y(new_n10807_));
  AOI22X1  g10614(.A0(\a[51] ), .A1(\a[43] ), .B0(\a[50] ), .B1(\a[44] ), .Y(new_n10808_));
  AND2X1   g10615(.A(\a[58] ), .B(\a[36] ), .Y(new_n10809_));
  INVX1    g10616(.A(new_n10809_), .Y(new_n10810_));
  AND2X1   g10617(.A(new_n4484_), .B(new_n4992_), .Y(new_n10811_));
  NOR3X1   g10618(.A(new_n10810_), .B(new_n10811_), .C(new_n10808_), .Y(new_n10812_));
  INVX1    g10619(.A(new_n10808_), .Y(new_n10813_));
  AOI21X1  g10620(.A0(new_n10809_), .A1(new_n10813_), .B0(new_n10811_), .Y(new_n10814_));
  INVX1    g10621(.A(new_n10814_), .Y(new_n10815_));
  OAI22X1  g10622(.A0(new_n10815_), .A1(new_n10808_), .B0(new_n10812_), .B1(new_n10810_), .Y(new_n10816_));
  OAI22X1  g10623(.A0(new_n7338_), .A1(new_n8071_), .B0(new_n5239_), .B1(new_n7618_), .Y(new_n10817_));
  OAI21X1  g10624(.A0(new_n7336_), .A1(new_n8069_), .B0(new_n10817_), .Y(new_n10818_));
  AND2X1   g10625(.A(\a[54] ), .B(\a[40] ), .Y(new_n10819_));
  OAI22X1  g10626(.A0(new_n5245_), .A1(new_n3081_), .B0(new_n4354_), .B1(new_n3096_), .Y(new_n10820_));
  AOI21X1  g10627(.A0(new_n5048_), .A1(new_n3607_), .B0(new_n10817_), .Y(new_n10821_));
  AOI22X1  g10628(.A0(new_n10821_), .A1(new_n10820_), .B0(new_n10819_), .B1(new_n10818_), .Y(new_n10822_));
  XOR2X1   g10629(.A(new_n10822_), .B(new_n10816_), .Y(new_n10823_));
  INVX1    g10630(.A(new_n10823_), .Y(new_n10824_));
  AND2X1   g10631(.A(\a[49] ), .B(\a[45] ), .Y(new_n10825_));
  NAND4X1  g10632(.A(\a[56] ), .B(\a[49] ), .C(\a[45] ), .D(\a[38] ), .Y(new_n10826_));
  OAI21X1  g10633(.A0(new_n4280_), .A1(new_n8873_), .B0(new_n10826_), .Y(new_n10827_));
  NAND4X1  g10634(.A(\a[56] ), .B(\a[48] ), .C(\a[46] ), .D(\a[38] ), .Y(new_n10828_));
  NAND2X1  g10635(.A(new_n10828_), .B(new_n10827_), .Y(new_n10829_));
  AOI21X1  g10636(.A0(new_n9701_), .A1(new_n8298_), .B0(new_n10827_), .Y(new_n10830_));
  OR2X1    g10637(.A(new_n9701_), .B(new_n8298_), .Y(new_n10831_));
  AOI22X1  g10638(.A0(new_n10831_), .A1(new_n10830_), .B0(new_n10829_), .B1(new_n10825_), .Y(new_n10832_));
  XOR2X1   g10639(.A(new_n10832_), .B(new_n10824_), .Y(new_n10833_));
  NOR2X1   g10640(.A(new_n10684_), .B(new_n10682_), .Y(new_n10834_));
  INVX1    g10641(.A(new_n10687_), .Y(new_n10835_));
  AOI21X1  g10642(.A0(new_n10835_), .A1(new_n10685_), .B0(new_n10834_), .Y(new_n10836_));
  XOR2X1   g10643(.A(new_n10836_), .B(new_n10833_), .Y(new_n10837_));
  NAND4X1  g10644(.A(\a[62] ), .B(\a[59] ), .C(\a[35] ), .D(\a[32] ), .Y(new_n10838_));
  NAND4X1  g10645(.A(\a[62] ), .B(\a[61] ), .C(\a[33] ), .D(\a[32] ), .Y(new_n10839_));
  AOI22X1  g10646(.A0(new_n10839_), .A1(new_n10838_), .B0(new_n6020_), .B1(new_n2120_), .Y(new_n10840_));
  AND2X1   g10647(.A(\a[62] ), .B(\a[32] ), .Y(new_n10841_));
  INVX1    g10648(.A(new_n10841_), .Y(new_n10842_));
  AOI21X1  g10649(.A0(new_n6020_), .A1(new_n2120_), .B0(new_n10840_), .Y(new_n10843_));
  INVX1    g10650(.A(new_n10843_), .Y(new_n10844_));
  AOI22X1  g10651(.A0(\a[61] ), .A1(\a[33] ), .B0(\a[59] ), .B1(\a[35] ), .Y(new_n10845_));
  OAI22X1  g10652(.A0(new_n10845_), .A1(new_n10844_), .B0(new_n10842_), .B1(new_n10840_), .Y(new_n10846_));
  XOR2X1   g10653(.A(new_n10846_), .B(new_n10754_), .Y(new_n10847_));
  AND2X1   g10654(.A(\a[60] ), .B(\a[57] ), .Y(new_n10848_));
  AOI22X1  g10655(.A0(new_n10848_), .A1(new_n7802_), .B0(new_n9461_), .B1(new_n3730_), .Y(new_n10849_));
  NOR4X1   g10656(.A(new_n5952_), .B(new_n4906_), .C(new_n2652_), .D(new_n2028_), .Y(new_n10850_));
  OR2X1    g10657(.A(new_n10850_), .B(new_n10849_), .Y(new_n10851_));
  AND2X1   g10658(.A(\a[57] ), .B(\a[37] ), .Y(new_n10852_));
  INVX1    g10659(.A(new_n10850_), .Y(new_n10853_));
  AND2X1   g10660(.A(new_n10853_), .B(new_n10849_), .Y(new_n10854_));
  OAI22X1  g10661(.A0(new_n5952_), .A1(new_n2028_), .B0(new_n4906_), .B1(new_n2652_), .Y(new_n10855_));
  AOI22X1  g10662(.A0(new_n10855_), .A1(new_n10854_), .B0(new_n10852_), .B1(new_n10851_), .Y(new_n10856_));
  XOR2X1   g10663(.A(new_n10856_), .B(new_n10847_), .Y(new_n10857_));
  XOR2X1   g10664(.A(new_n10857_), .B(new_n10837_), .Y(new_n10858_));
  XOR2X1   g10665(.A(new_n10858_), .B(new_n10807_), .Y(new_n10859_));
  XOR2X1   g10666(.A(new_n10859_), .B(new_n10795_), .Y(new_n10860_));
  INVX1    g10667(.A(new_n10860_), .Y(new_n10861_));
  AND2X1   g10668(.A(new_n10702_), .B(new_n10678_), .Y(new_n10862_));
  AOI21X1  g10669(.A0(new_n10770_), .A1(new_n10703_), .B0(new_n10862_), .Y(new_n10863_));
  XOR2X1   g10670(.A(new_n10863_), .B(new_n10861_), .Y(new_n10864_));
  INVX1    g10671(.A(new_n10772_), .Y(new_n10865_));
  OAI21X1  g10672(.A0(new_n10773_), .A1(new_n10673_), .B0(new_n10865_), .Y(new_n10866_));
  XOR2X1   g10673(.A(new_n10866_), .B(new_n10864_), .Y(\asquared[95] ));
  AND2X1   g10674(.A(new_n10806_), .B(new_n10798_), .Y(new_n10868_));
  AOI21X1  g10675(.A0(new_n10858_), .A1(new_n10807_), .B0(new_n10868_), .Y(new_n10869_));
  INVX1    g10676(.A(new_n10869_), .Y(new_n10870_));
  NOR2X1   g10677(.A(new_n10836_), .B(new_n10833_), .Y(new_n10871_));
  AOI21X1  g10678(.A0(new_n10857_), .A1(new_n10837_), .B0(new_n10871_), .Y(new_n10872_));
  NAND2X1  g10679(.A(\a[59] ), .B(\a[36] ), .Y(new_n10873_));
  NAND2X1  g10680(.A(\a[60] ), .B(\a[35] ), .Y(new_n10874_));
  AOI22X1  g10681(.A0(new_n10874_), .A1(new_n10873_), .B0(new_n6427_), .B1(new_n2682_), .Y(new_n10875_));
  XOR2X1   g10682(.A(new_n10875_), .B(new_n10830_), .Y(new_n10876_));
  NOR3X1   g10683(.A(new_n10761_), .B(new_n6549_), .C(new_n1704_), .Y(new_n10877_));
  AOI21X1  g10684(.A0(new_n10799_), .A1(new_n10747_), .B0(new_n10877_), .Y(new_n10878_));
  XOR2X1   g10685(.A(new_n10878_), .B(new_n10876_), .Y(new_n10879_));
  INVX1    g10686(.A(new_n10879_), .Y(new_n10880_));
  AND2X1   g10687(.A(new_n10726_), .B(new_n10716_), .Y(new_n10881_));
  AOI21X1  g10688(.A0(new_n10804_), .A1(new_n10736_), .B0(new_n10881_), .Y(new_n10882_));
  XOR2X1   g10689(.A(new_n10882_), .B(new_n10880_), .Y(new_n10883_));
  NOR2X1   g10690(.A(new_n10802_), .B(new_n10800_), .Y(new_n10884_));
  AOI21X1  g10691(.A0(new_n10805_), .A1(new_n10803_), .B0(new_n10884_), .Y(new_n10885_));
  XOR2X1   g10692(.A(new_n10885_), .B(new_n10883_), .Y(new_n10886_));
  XOR2X1   g10693(.A(new_n10886_), .B(new_n10872_), .Y(new_n10887_));
  XOR2X1   g10694(.A(new_n10887_), .B(new_n10870_), .Y(new_n10888_));
  NAND3X1  g10695(.A(\a[62] ), .B(\a[48] ), .C(\a[33] ), .Y(new_n10889_));
  AND2X1   g10696(.A(new_n10889_), .B(new_n8297_), .Y(new_n10890_));
  OAI21X1  g10697(.A0(new_n6606_), .A1(new_n1851_), .B0(new_n3926_), .Y(new_n10891_));
  NOR3X1   g10698(.A(new_n10889_), .B(new_n3926_), .C(new_n4041_), .Y(new_n10892_));
  AOI21X1  g10699(.A0(new_n10891_), .A1(new_n10890_), .B0(new_n10892_), .Y(new_n10893_));
  AOI22X1  g10700(.A0(\a[50] ), .A1(\a[45] ), .B0(\a[49] ), .B1(\a[46] ), .Y(new_n10894_));
  AND2X1   g10701(.A(\a[56] ), .B(\a[39] ), .Y(new_n10895_));
  AND2X1   g10702(.A(new_n4321_), .B(new_n3809_), .Y(new_n10896_));
  OAI21X1  g10703(.A0(new_n10896_), .A1(new_n10894_), .B0(new_n10895_), .Y(new_n10897_));
  INVX1    g10704(.A(new_n10895_), .Y(new_n10898_));
  OAI22X1  g10705(.A0(new_n10894_), .A1(new_n10898_), .B0(new_n7652_), .B1(new_n8873_), .Y(new_n10899_));
  OAI21X1  g10706(.A0(new_n10899_), .A1(new_n10894_), .B0(new_n10897_), .Y(new_n10900_));
  XOR2X1   g10707(.A(new_n10900_), .B(new_n10893_), .Y(new_n10901_));
  OAI22X1  g10708(.A0(new_n7336_), .A1(new_n6502_), .B0(new_n8145_), .B1(new_n3212_), .Y(new_n10902_));
  OAI21X1  g10709(.A0(new_n7793_), .A1(new_n7353_), .B0(new_n10902_), .Y(new_n10903_));
  AND2X1   g10710(.A(\a[53] ), .B(\a[42] ), .Y(new_n10904_));
  OAI22X1  g10711(.A0(new_n4354_), .A1(new_n3037_), .B0(new_n4349_), .B1(new_n5268_), .Y(new_n10905_));
  AOI21X1  g10712(.A0(new_n7164_), .A1(new_n4992_), .B0(new_n10902_), .Y(new_n10906_));
  AOI22X1  g10713(.A0(new_n10906_), .A1(new_n10905_), .B0(new_n10904_), .B1(new_n10903_), .Y(new_n10907_));
  XOR2X1   g10714(.A(new_n10907_), .B(new_n10901_), .Y(new_n10908_));
  AND2X1   g10715(.A(new_n10784_), .B(new_n10782_), .Y(new_n10909_));
  OR2X1    g10716(.A(new_n10784_), .B(new_n10782_), .Y(new_n10910_));
  OAI21X1  g10717(.A0(new_n10787_), .A1(new_n10909_), .B0(new_n10910_), .Y(new_n10911_));
  XOR2X1   g10718(.A(new_n10911_), .B(new_n10908_), .Y(new_n10912_));
  AOI22X1  g10719(.A0(\a[63] ), .A1(\a[32] ), .B0(\a[61] ), .B1(\a[34] ), .Y(new_n10913_));
  AND2X1   g10720(.A(\a[54] ), .B(\a[41] ), .Y(new_n10914_));
  INVX1    g10721(.A(new_n10914_), .Y(new_n10915_));
  AND2X1   g10722(.A(new_n6688_), .B(new_n2820_), .Y(new_n10916_));
  NOR3X1   g10723(.A(new_n10915_), .B(new_n10916_), .C(new_n10913_), .Y(new_n10917_));
  NOR2X1   g10724(.A(new_n10917_), .B(new_n10916_), .Y(new_n10918_));
  INVX1    g10725(.A(new_n10918_), .Y(new_n10919_));
  OAI22X1  g10726(.A0(new_n10919_), .A1(new_n10913_), .B0(new_n10917_), .B1(new_n10915_), .Y(new_n10920_));
  NAND4X1  g10727(.A(\a[58] ), .B(\a[55] ), .C(\a[40] ), .D(\a[37] ), .Y(new_n10921_));
  NAND4X1  g10728(.A(\a[58] ), .B(\a[57] ), .C(\a[38] ), .D(\a[37] ), .Y(new_n10922_));
  AOI22X1  g10729(.A0(new_n10922_), .A1(new_n10921_), .B0(new_n9461_), .B1(new_n2663_), .Y(new_n10923_));
  NAND2X1  g10730(.A(\a[58] ), .B(\a[37] ), .Y(new_n10924_));
  NAND4X1  g10731(.A(\a[57] ), .B(\a[55] ), .C(\a[40] ), .D(\a[38] ), .Y(new_n10925_));
  NAND3X1  g10732(.A(new_n10922_), .B(new_n10921_), .C(new_n10925_), .Y(new_n10926_));
  AOI22X1  g10733(.A0(\a[57] ), .A1(\a[38] ), .B0(\a[55] ), .B1(\a[40] ), .Y(new_n10927_));
  OAI22X1  g10734(.A0(new_n10927_), .A1(new_n10926_), .B0(new_n10924_), .B1(new_n10923_), .Y(new_n10928_));
  XOR2X1   g10735(.A(new_n10928_), .B(new_n10814_), .Y(new_n10929_));
  XOR2X1   g10736(.A(new_n10929_), .B(new_n10920_), .Y(new_n10930_));
  XOR2X1   g10737(.A(new_n10930_), .B(new_n10912_), .Y(new_n10931_));
  INVX1    g10738(.A(new_n10931_), .Y(new_n10932_));
  NOR2X1   g10739(.A(new_n10791_), .B(new_n10788_), .Y(new_n10933_));
  AOI21X1  g10740(.A0(new_n10792_), .A1(new_n10780_), .B0(new_n10933_), .Y(new_n10934_));
  INVX1    g10741(.A(new_n10821_), .Y(new_n10935_));
  XOR2X1   g10742(.A(new_n10854_), .B(new_n10843_), .Y(new_n10936_));
  XOR2X1   g10743(.A(new_n10936_), .B(new_n10935_), .Y(new_n10937_));
  INVX1    g10744(.A(new_n10816_), .Y(new_n10938_));
  OR2X1    g10745(.A(new_n10822_), .B(new_n10938_), .Y(new_n10939_));
  OAI21X1  g10746(.A0(new_n10832_), .A1(new_n10823_), .B0(new_n10939_), .Y(new_n10940_));
  NOR2X1   g10747(.A(new_n10856_), .B(new_n10847_), .Y(new_n10941_));
  AOI21X1  g10748(.A0(new_n10846_), .A1(new_n10755_), .B0(new_n10941_), .Y(new_n10942_));
  INVX1    g10749(.A(new_n10942_), .Y(new_n10943_));
  XOR2X1   g10750(.A(new_n10943_), .B(new_n10940_), .Y(new_n10944_));
  XOR2X1   g10751(.A(new_n10944_), .B(new_n10937_), .Y(new_n10945_));
  XOR2X1   g10752(.A(new_n10945_), .B(new_n10934_), .Y(new_n10946_));
  XOR2X1   g10753(.A(new_n10946_), .B(new_n10932_), .Y(new_n10947_));
  XOR2X1   g10754(.A(new_n10947_), .B(new_n10888_), .Y(new_n10948_));
  NOR2X1   g10755(.A(new_n10794_), .B(new_n10777_), .Y(new_n10949_));
  AOI21X1  g10756(.A0(new_n10859_), .A1(new_n10795_), .B0(new_n10949_), .Y(new_n10950_));
  NOR2X1   g10757(.A(new_n10950_), .B(new_n10948_), .Y(new_n10951_));
  AND2X1   g10758(.A(new_n10950_), .B(new_n10948_), .Y(new_n10952_));
  OR2X1    g10759(.A(new_n10952_), .B(new_n10951_), .Y(new_n10953_));
  AND2X1   g10760(.A(new_n10863_), .B(new_n10861_), .Y(new_n10954_));
  INVX1    g10761(.A(new_n10954_), .Y(new_n10955_));
  NOR2X1   g10762(.A(new_n10863_), .B(new_n10861_), .Y(new_n10956_));
  AOI21X1  g10763(.A0(new_n10866_), .A1(new_n10955_), .B0(new_n10956_), .Y(new_n10957_));
  XOR2X1   g10764(.A(new_n10957_), .B(new_n10953_), .Y(\asquared[96] ));
  NOR2X1   g10765(.A(new_n10887_), .B(new_n10870_), .Y(new_n10959_));
  NAND2X1  g10766(.A(new_n10887_), .B(new_n10870_), .Y(new_n10960_));
  OAI21X1  g10767(.A0(new_n10947_), .A1(new_n10959_), .B0(new_n10960_), .Y(new_n10961_));
  AND2X1   g10768(.A(new_n10911_), .B(new_n10908_), .Y(new_n10962_));
  INVX1    g10769(.A(new_n10962_), .Y(new_n10963_));
  INVX1    g10770(.A(new_n10912_), .Y(new_n10964_));
  OAI21X1  g10771(.A0(new_n10930_), .A1(new_n10964_), .B0(new_n10963_), .Y(new_n10965_));
  NAND4X1  g10772(.A(\a[59] ), .B(\a[56] ), .C(\a[40] ), .D(\a[37] ), .Y(new_n10966_));
  AND2X1   g10773(.A(\a[60] ), .B(\a[40] ), .Y(new_n10967_));
  AOI22X1  g10774(.A0(new_n10967_), .A1(new_n10609_), .B0(new_n6427_), .B1(new_n3330_), .Y(new_n10968_));
  AND2X1   g10775(.A(new_n10968_), .B(new_n10966_), .Y(new_n10969_));
  INVX1    g10776(.A(new_n10969_), .Y(new_n10970_));
  AOI22X1  g10777(.A0(\a[59] ), .A1(\a[37] ), .B0(\a[56] ), .B1(\a[40] ), .Y(new_n10971_));
  NOR4X1   g10778(.A(new_n5617_), .B(new_n6022_), .C(new_n3036_), .D(new_n2345_), .Y(new_n10972_));
  AND2X1   g10779(.A(\a[60] ), .B(\a[36] ), .Y(new_n10973_));
  OAI21X1  g10780(.A0(new_n10968_), .A1(new_n10972_), .B0(new_n10973_), .Y(new_n10974_));
  OAI21X1  g10781(.A0(new_n10971_), .A1(new_n10970_), .B0(new_n10974_), .Y(new_n10975_));
  AOI22X1  g10782(.A0(\a[58] ), .A1(\a[38] ), .B0(\a[57] ), .B1(\a[39] ), .Y(new_n10976_));
  AND2X1   g10783(.A(new_n6119_), .B(new_n3503_), .Y(new_n10977_));
  NOR3X1   g10784(.A(new_n10976_), .B(new_n10977_), .C(new_n5885_), .Y(new_n10978_));
  NOR2X1   g10785(.A(new_n10978_), .B(new_n10977_), .Y(new_n10979_));
  INVX1    g10786(.A(new_n10979_), .Y(new_n10980_));
  OAI22X1  g10787(.A0(new_n10980_), .A1(new_n10976_), .B0(new_n10978_), .B1(new_n5885_), .Y(new_n10981_));
  XOR2X1   g10788(.A(new_n10981_), .B(new_n10975_), .Y(new_n10982_));
  NAND4X1  g10789(.A(\a[51] ), .B(\a[49] ), .C(\a[47] ), .D(\a[45] ), .Y(new_n10983_));
  NAND4X1  g10790(.A(\a[51] ), .B(\a[50] ), .C(\a[46] ), .D(\a[45] ), .Y(new_n10984_));
  AOI22X1  g10791(.A0(new_n10984_), .A1(new_n10983_), .B0(new_n4321_), .B1(new_n3893_), .Y(new_n10985_));
  NOR3X1   g10792(.A(new_n10985_), .B(new_n4349_), .C(new_n3811_), .Y(new_n10986_));
  AOI21X1  g10793(.A0(new_n4321_), .A1(new_n3893_), .B0(new_n10985_), .Y(new_n10987_));
  OAI22X1  g10794(.A0(new_n4983_), .A1(new_n3460_), .B0(new_n3915_), .B1(new_n4041_), .Y(new_n10988_));
  AOI21X1  g10795(.A0(new_n10988_), .A1(new_n10987_), .B0(new_n10986_), .Y(new_n10989_));
  XOR2X1   g10796(.A(new_n10989_), .B(new_n10982_), .Y(new_n10990_));
  NAND2X1  g10797(.A(new_n10943_), .B(new_n10940_), .Y(new_n10991_));
  NAND2X1  g10798(.A(new_n10944_), .B(new_n10937_), .Y(new_n10992_));
  NAND2X1  g10799(.A(new_n10992_), .B(new_n10991_), .Y(new_n10993_));
  XOR2X1   g10800(.A(new_n10993_), .B(new_n10990_), .Y(new_n10994_));
  XOR2X1   g10801(.A(new_n10994_), .B(new_n10965_), .Y(new_n10995_));
  INVX1    g10802(.A(new_n10945_), .Y(new_n10996_));
  OR2X1    g10803(.A(new_n10996_), .B(new_n10934_), .Y(new_n10997_));
  OAI21X1  g10804(.A0(new_n10946_), .A1(new_n10931_), .B0(new_n10997_), .Y(new_n10998_));
  XOR2X1   g10805(.A(new_n10998_), .B(new_n10995_), .Y(new_n10999_));
  INVX1    g10806(.A(new_n10883_), .Y(new_n11000_));
  OR2X1    g10807(.A(new_n10885_), .B(new_n11000_), .Y(new_n11001_));
  OAI21X1  g10808(.A0(new_n10886_), .A1(new_n10872_), .B0(new_n11001_), .Y(new_n11002_));
  INVX1    g10809(.A(new_n10890_), .Y(new_n11003_));
  XOR2X1   g10810(.A(new_n10899_), .B(new_n11003_), .Y(new_n11004_));
  INVX1    g10811(.A(new_n11004_), .Y(new_n11005_));
  XOR2X1   g10812(.A(new_n11005_), .B(new_n10906_), .Y(new_n11006_));
  INVX1    g10813(.A(new_n10920_), .Y(new_n11007_));
  OAI21X1  g10814(.A0(new_n10812_), .A1(new_n10811_), .B0(new_n10928_), .Y(new_n11008_));
  OAI21X1  g10815(.A0(new_n10929_), .A1(new_n11007_), .B0(new_n11008_), .Y(new_n11009_));
  INVX1    g10816(.A(new_n10900_), .Y(new_n11010_));
  OR2X1    g10817(.A(new_n10907_), .B(new_n10901_), .Y(new_n11011_));
  OAI21X1  g10818(.A0(new_n11010_), .A1(new_n10893_), .B0(new_n11011_), .Y(new_n11012_));
  XOR2X1   g10819(.A(new_n11012_), .B(new_n11009_), .Y(new_n11013_));
  XOR2X1   g10820(.A(new_n11013_), .B(new_n11006_), .Y(new_n11014_));
  XOR2X1   g10821(.A(new_n11014_), .B(new_n11002_), .Y(new_n11015_));
  NAND4X1  g10822(.A(\a[63] ), .B(\a[61] ), .C(\a[35] ), .D(\a[33] ), .Y(new_n11016_));
  NAND4X1  g10823(.A(\a[63] ), .B(\a[62] ), .C(\a[34] ), .D(\a[33] ), .Y(new_n11017_));
  AOI22X1  g10824(.A0(new_n11017_), .A1(new_n11016_), .B0(new_n6556_), .B1(new_n2361_), .Y(new_n11018_));
  NAND4X1  g10825(.A(\a[62] ), .B(\a[61] ), .C(\a[35] ), .D(\a[34] ), .Y(new_n11019_));
  NAND3X1  g10826(.A(new_n11017_), .B(new_n11016_), .C(new_n11019_), .Y(new_n11020_));
  AOI22X1  g10827(.A0(\a[62] ), .A1(\a[34] ), .B0(\a[61] ), .B1(\a[35] ), .Y(new_n11021_));
  NAND2X1  g10828(.A(\a[63] ), .B(\a[33] ), .Y(new_n11022_));
  OAI22X1  g10829(.A0(new_n11022_), .A1(new_n11018_), .B0(new_n11021_), .B1(new_n11020_), .Y(new_n11023_));
  INVX1    g10830(.A(new_n5745_), .Y(new_n11024_));
  NAND4X1  g10831(.A(\a[55] ), .B(\a[53] ), .C(\a[43] ), .D(\a[41] ), .Y(new_n11025_));
  NAND4X1  g10832(.A(\a[55] ), .B(\a[54] ), .C(\a[42] ), .D(\a[41] ), .Y(new_n11026_));
  AOI22X1  g10833(.A0(new_n11026_), .A1(new_n11025_), .B0(new_n5238_), .B1(new_n3462_), .Y(new_n11027_));
  AOI22X1  g10834(.A0(\a[54] ), .A1(\a[42] ), .B0(\a[53] ), .B1(\a[43] ), .Y(new_n11028_));
  AOI21X1  g10835(.A0(new_n5238_), .A1(new_n3462_), .B0(new_n11027_), .Y(new_n11029_));
  INVX1    g10836(.A(new_n11029_), .Y(new_n11030_));
  OAI22X1  g10837(.A0(new_n11030_), .A1(new_n11028_), .B0(new_n11027_), .B1(new_n11024_), .Y(new_n11031_));
  XOR2X1   g10838(.A(new_n11031_), .B(new_n11023_), .Y(new_n11032_));
  AOI21X1  g10839(.A0(new_n10851_), .A1(new_n10853_), .B0(new_n10843_), .Y(new_n11033_));
  AOI21X1  g10840(.A0(new_n10936_), .A1(new_n10935_), .B0(new_n11033_), .Y(new_n11034_));
  XOR2X1   g10841(.A(new_n11034_), .B(new_n11032_), .Y(new_n11035_));
  XOR2X1   g10842(.A(new_n10926_), .B(new_n10919_), .Y(new_n11036_));
  INVX1    g10843(.A(new_n10830_), .Y(new_n11037_));
  AOI22X1  g10844(.A0(new_n10875_), .A1(new_n11037_), .B0(new_n6427_), .B1(new_n2682_), .Y(new_n11038_));
  INVX1    g10845(.A(new_n11038_), .Y(new_n11039_));
  XOR2X1   g10846(.A(new_n11039_), .B(new_n11036_), .Y(new_n11040_));
  OR2X1    g10847(.A(new_n10878_), .B(new_n10876_), .Y(new_n11041_));
  OAI21X1  g10848(.A0(new_n10882_), .A1(new_n10880_), .B0(new_n11041_), .Y(new_n11042_));
  XOR2X1   g10849(.A(new_n11042_), .B(new_n11040_), .Y(new_n11043_));
  XOR2X1   g10850(.A(new_n11043_), .B(new_n11035_), .Y(new_n11044_));
  XOR2X1   g10851(.A(new_n11044_), .B(new_n11015_), .Y(new_n11045_));
  OR2X1    g10852(.A(new_n11045_), .B(new_n10999_), .Y(new_n11046_));
  AND2X1   g10853(.A(new_n10998_), .B(new_n10995_), .Y(new_n11047_));
  OAI21X1  g10854(.A0(new_n10998_), .A1(new_n10995_), .B0(new_n11045_), .Y(new_n11048_));
  OR2X1    g10855(.A(new_n11048_), .B(new_n11047_), .Y(new_n11049_));
  AND2X1   g10856(.A(new_n11049_), .B(new_n11046_), .Y(new_n11050_));
  AND2X1   g10857(.A(new_n11050_), .B(new_n10961_), .Y(new_n11051_));
  INVX1    g10858(.A(new_n11051_), .Y(new_n11052_));
  INVX1    g10859(.A(new_n10951_), .Y(new_n11053_));
  OAI21X1  g10860(.A0(new_n10957_), .A1(new_n10952_), .B0(new_n11053_), .Y(new_n11054_));
  NOR2X1   g10861(.A(new_n11050_), .B(new_n10961_), .Y(new_n11055_));
  INVX1    g10862(.A(new_n11055_), .Y(new_n11056_));
  AOI21X1  g10863(.A0(new_n11052_), .A1(new_n11056_), .B0(new_n11054_), .Y(new_n11057_));
  AND2X1   g10864(.A(new_n11056_), .B(new_n11054_), .Y(new_n11058_));
  AOI21X1  g10865(.A0(new_n11058_), .A1(new_n11052_), .B0(new_n11057_), .Y(\asquared[97] ));
  AOI21X1  g10866(.A0(new_n11056_), .A1(new_n11054_), .B0(new_n11051_), .Y(new_n11060_));
  INVX1    g10867(.A(new_n10998_), .Y(new_n11061_));
  OAI21X1  g10868(.A0(new_n11061_), .A1(new_n10995_), .B0(new_n11046_), .Y(new_n11062_));
  AOI21X1  g10869(.A0(new_n10992_), .A1(new_n10991_), .B0(new_n10990_), .Y(new_n11063_));
  INVX1    g10870(.A(new_n10965_), .Y(new_n11064_));
  NOR2X1   g10871(.A(new_n10994_), .B(new_n11064_), .Y(new_n11065_));
  NOR2X1   g10872(.A(new_n11065_), .B(new_n11063_), .Y(new_n11066_));
  NAND2X1  g10873(.A(\a[61] ), .B(\a[36] ), .Y(new_n11067_));
  XOR2X1   g10874(.A(new_n11067_), .B(new_n10987_), .Y(new_n11068_));
  XOR2X1   g10875(.A(new_n11068_), .B(new_n10979_), .Y(new_n11069_));
  NAND2X1  g10876(.A(new_n10981_), .B(new_n10975_), .Y(new_n11070_));
  INVX1    g10877(.A(new_n10982_), .Y(new_n11071_));
  OAI21X1  g10878(.A0(new_n10989_), .A1(new_n11071_), .B0(new_n11070_), .Y(new_n11072_));
  AND2X1   g10879(.A(new_n10926_), .B(new_n10919_), .Y(new_n11073_));
  AOI21X1  g10880(.A0(new_n11039_), .A1(new_n11036_), .B0(new_n11073_), .Y(new_n11074_));
  XOR2X1   g10881(.A(new_n11074_), .B(new_n11072_), .Y(new_n11075_));
  XOR2X1   g10882(.A(new_n11075_), .B(new_n11069_), .Y(new_n11076_));
  NAND3X1  g10883(.A(\a[62] ), .B(\a[49] ), .C(\a[35] ), .Y(new_n11077_));
  AND2X1   g10884(.A(new_n11077_), .B(new_n4280_), .Y(new_n11078_));
  OAI21X1  g10885(.A0(new_n6606_), .A1(new_n2557_), .B0(new_n3915_), .Y(new_n11079_));
  NOR3X1   g10886(.A(new_n11077_), .B(new_n3915_), .C(new_n3926_), .Y(new_n11080_));
  AOI21X1  g10887(.A0(new_n11079_), .A1(new_n11078_), .B0(new_n11080_), .Y(new_n11081_));
  AND2X1   g10888(.A(\a[57] ), .B(\a[40] ), .Y(new_n11082_));
  AOI22X1  g10889(.A0(\a[51] ), .A1(\a[46] ), .B0(\a[50] ), .B1(\a[47] ), .Y(new_n11083_));
  INVX1    g10890(.A(new_n11083_), .Y(new_n11084_));
  NAND4X1  g10891(.A(\a[51] ), .B(\a[50] ), .C(\a[47] ), .D(\a[46] ), .Y(new_n11085_));
  NAND3X1  g10892(.A(new_n11084_), .B(new_n11085_), .C(new_n11082_), .Y(new_n11086_));
  AOI22X1  g10893(.A0(new_n11084_), .A1(new_n11082_), .B0(new_n4484_), .B1(new_n3893_), .Y(new_n11087_));
  AOI22X1  g10894(.A0(new_n11087_), .A1(new_n11084_), .B0(new_n11086_), .B1(new_n11082_), .Y(new_n11088_));
  XOR2X1   g10895(.A(new_n11088_), .B(new_n11081_), .Y(new_n11089_));
  NAND2X1  g10896(.A(new_n10899_), .B(new_n11003_), .Y(new_n11090_));
  OAI21X1  g10897(.A0(new_n11005_), .A1(new_n10906_), .B0(new_n11090_), .Y(new_n11091_));
  XOR2X1   g10898(.A(new_n11091_), .B(new_n11089_), .Y(new_n11092_));
  XOR2X1   g10899(.A(new_n11020_), .B(new_n10970_), .Y(new_n11093_));
  XOR2X1   g10900(.A(new_n11093_), .B(new_n11029_), .Y(new_n11094_));
  AND2X1   g10901(.A(new_n11031_), .B(new_n11023_), .Y(new_n11095_));
  INVX1    g10902(.A(new_n11034_), .Y(new_n11096_));
  AOI21X1  g10903(.A0(new_n11096_), .A1(new_n11032_), .B0(new_n11095_), .Y(new_n11097_));
  XOR2X1   g10904(.A(new_n11097_), .B(new_n11094_), .Y(new_n11098_));
  XOR2X1   g10905(.A(new_n11098_), .B(new_n11092_), .Y(new_n11099_));
  XOR2X1   g10906(.A(new_n11099_), .B(new_n11076_), .Y(new_n11100_));
  XOR2X1   g10907(.A(new_n11100_), .B(new_n11066_), .Y(new_n11101_));
  NOR2X1   g10908(.A(new_n11042_), .B(new_n11040_), .Y(new_n11102_));
  NAND2X1  g10909(.A(new_n11042_), .B(new_n11040_), .Y(new_n11103_));
  OAI21X1  g10910(.A0(new_n11102_), .A1(new_n11035_), .B0(new_n11103_), .Y(new_n11104_));
  NAND2X1  g10911(.A(\a[56] ), .B(\a[41] ), .Y(new_n11105_));
  NOR4X1   g10912(.A(new_n6549_), .B(new_n4906_), .C(new_n3096_), .D(new_n2028_), .Y(new_n11106_));
  NAND4X1  g10913(.A(\a[56] ), .B(\a[55] ), .C(\a[42] ), .D(\a[41] ), .Y(new_n11107_));
  NAND4X1  g10914(.A(\a[63] ), .B(\a[56] ), .C(\a[41] ), .D(\a[34] ), .Y(new_n11108_));
  AOI21X1  g10915(.A0(new_n11108_), .A1(new_n11107_), .B0(new_n11106_), .Y(new_n11109_));
  OR2X1    g10916(.A(new_n11109_), .B(new_n11106_), .Y(new_n11110_));
  AOI22X1  g10917(.A0(\a[63] ), .A1(\a[34] ), .B0(\a[55] ), .B1(\a[42] ), .Y(new_n11111_));
  OAI22X1  g10918(.A0(new_n11111_), .A1(new_n11110_), .B0(new_n11109_), .B1(new_n11105_), .Y(new_n11112_));
  NAND4X1  g10919(.A(\a[60] ), .B(\a[58] ), .C(\a[39] ), .D(\a[37] ), .Y(new_n11113_));
  NAND4X1  g10920(.A(\a[60] ), .B(\a[59] ), .C(\a[38] ), .D(\a[37] ), .Y(new_n11114_));
  AOI22X1  g10921(.A0(new_n11114_), .A1(new_n11113_), .B0(new_n6121_), .B1(new_n3503_), .Y(new_n11115_));
  NAND2X1  g10922(.A(\a[60] ), .B(\a[37] ), .Y(new_n11116_));
  NAND4X1  g10923(.A(\a[59] ), .B(\a[58] ), .C(\a[39] ), .D(\a[38] ), .Y(new_n11117_));
  NAND3X1  g10924(.A(new_n11114_), .B(new_n11113_), .C(new_n11117_), .Y(new_n11118_));
  AOI22X1  g10925(.A0(\a[59] ), .A1(\a[38] ), .B0(\a[58] ), .B1(\a[39] ), .Y(new_n11119_));
  OAI22X1  g10926(.A0(new_n11119_), .A1(new_n11118_), .B0(new_n11116_), .B1(new_n11115_), .Y(new_n11120_));
  XOR2X1   g10927(.A(new_n11120_), .B(new_n11112_), .Y(new_n11121_));
  AOI22X1  g10928(.A0(new_n7337_), .A1(new_n7640_), .B0(new_n5238_), .B1(new_n4992_), .Y(new_n11122_));
  AOI21X1  g10929(.A0(new_n5048_), .A1(new_n3918_), .B0(new_n11122_), .Y(new_n11123_));
  AND2X1   g10930(.A(\a[54] ), .B(\a[43] ), .Y(new_n11124_));
  INVX1    g10931(.A(new_n11124_), .Y(new_n11125_));
  AOI22X1  g10932(.A0(\a[53] ), .A1(\a[44] ), .B0(\a[52] ), .B1(\a[45] ), .Y(new_n11126_));
  OAI22X1  g10933(.A0(new_n7338_), .A1(new_n7641_), .B0(new_n5239_), .B1(new_n7353_), .Y(new_n11127_));
  AOI21X1  g10934(.A0(new_n5048_), .A1(new_n3918_), .B0(new_n11127_), .Y(new_n11128_));
  INVX1    g10935(.A(new_n11128_), .Y(new_n11129_));
  OAI22X1  g10936(.A0(new_n11129_), .A1(new_n11126_), .B0(new_n11125_), .B1(new_n11123_), .Y(new_n11130_));
  INVX1    g10937(.A(new_n11130_), .Y(new_n11131_));
  XOR2X1   g10938(.A(new_n11131_), .B(new_n11121_), .Y(new_n11132_));
  AND2X1   g10939(.A(new_n11012_), .B(new_n11009_), .Y(new_n11133_));
  AOI21X1  g10940(.A0(new_n11013_), .A1(new_n11006_), .B0(new_n11133_), .Y(new_n11134_));
  XOR2X1   g10941(.A(new_n11134_), .B(new_n11132_), .Y(new_n11135_));
  XOR2X1   g10942(.A(new_n11135_), .B(new_n11104_), .Y(new_n11136_));
  INVX1    g10943(.A(new_n11136_), .Y(new_n11137_));
  NAND2X1  g10944(.A(new_n11014_), .B(new_n11002_), .Y(new_n11138_));
  NOR2X1   g10945(.A(new_n11014_), .B(new_n11002_), .Y(new_n11139_));
  OAI21X1  g10946(.A0(new_n11044_), .A1(new_n11139_), .B0(new_n11138_), .Y(new_n11140_));
  XOR2X1   g10947(.A(new_n11140_), .B(new_n11137_), .Y(new_n11141_));
  XOR2X1   g10948(.A(new_n11141_), .B(new_n11101_), .Y(new_n11142_));
  AND2X1   g10949(.A(new_n11142_), .B(new_n11062_), .Y(new_n11143_));
  NOR2X1   g10950(.A(new_n11142_), .B(new_n11062_), .Y(new_n11144_));
  OR2X1    g10951(.A(new_n11144_), .B(new_n11143_), .Y(new_n11145_));
  XOR2X1   g10952(.A(new_n11145_), .B(new_n11060_), .Y(\asquared[98] ));
  NAND2X1  g10953(.A(new_n11140_), .B(new_n11136_), .Y(new_n11147_));
  OAI21X1  g10954(.A0(new_n11141_), .A1(new_n11101_), .B0(new_n11147_), .Y(new_n11148_));
  NOR2X1   g10955(.A(new_n11134_), .B(new_n11132_), .Y(new_n11149_));
  AOI21X1  g10956(.A0(new_n11135_), .A1(new_n11104_), .B0(new_n11149_), .Y(new_n11150_));
  AND2X1   g10957(.A(new_n11020_), .B(new_n10970_), .Y(new_n11151_));
  AOI21X1  g10958(.A0(new_n11093_), .A1(new_n11030_), .B0(new_n11151_), .Y(new_n11152_));
  NOR2X1   g10959(.A(new_n11067_), .B(new_n10987_), .Y(new_n11153_));
  AOI21X1  g10960(.A0(new_n11068_), .A1(new_n10980_), .B0(new_n11153_), .Y(new_n11154_));
  INVX1    g10961(.A(new_n11154_), .Y(new_n11155_));
  XOR2X1   g10962(.A(new_n11155_), .B(new_n11152_), .Y(new_n11156_));
  AND2X1   g10963(.A(new_n11120_), .B(new_n11112_), .Y(new_n11157_));
  AOI21X1  g10964(.A0(new_n11130_), .A1(new_n11121_), .B0(new_n11157_), .Y(new_n11158_));
  XOR2X1   g10965(.A(new_n11158_), .B(new_n11156_), .Y(new_n11159_));
  XOR2X1   g10966(.A(new_n11118_), .B(new_n11110_), .Y(new_n11160_));
  XOR2X1   g10967(.A(new_n11160_), .B(new_n11128_), .Y(new_n11161_));
  NOR2X1   g10968(.A(new_n11088_), .B(new_n11081_), .Y(new_n11162_));
  AOI21X1  g10969(.A0(new_n11091_), .A1(new_n11089_), .B0(new_n11162_), .Y(new_n11163_));
  XOR2X1   g10970(.A(new_n11163_), .B(new_n11161_), .Y(new_n11164_));
  AOI22X1  g10971(.A0(\a[59] ), .A1(\a[39] ), .B0(\a[58] ), .B1(\a[40] ), .Y(new_n11165_));
  AND2X1   g10972(.A(\a[53] ), .B(\a[45] ), .Y(new_n11166_));
  INVX1    g10973(.A(new_n11166_), .Y(new_n11167_));
  AND2X1   g10974(.A(new_n6121_), .B(new_n4077_), .Y(new_n11168_));
  NOR3X1   g10975(.A(new_n11167_), .B(new_n11168_), .C(new_n11165_), .Y(new_n11169_));
  INVX1    g10976(.A(new_n11165_), .Y(new_n11170_));
  AOI21X1  g10977(.A0(new_n11166_), .A1(new_n11170_), .B0(new_n11168_), .Y(new_n11171_));
  INVX1    g10978(.A(new_n11171_), .Y(new_n11172_));
  OAI22X1  g10979(.A0(new_n11172_), .A1(new_n11165_), .B0(new_n11169_), .B1(new_n11167_), .Y(new_n11173_));
  NAND4X1  g10980(.A(\a[52] ), .B(\a[51] ), .C(\a[47] ), .D(\a[46] ), .Y(new_n11174_));
  NAND4X1  g10981(.A(\a[52] ), .B(\a[50] ), .C(\a[48] ), .D(\a[46] ), .Y(new_n11175_));
  AOI22X1  g10982(.A0(new_n11175_), .A1(new_n11174_), .B0(new_n4484_), .B1(new_n4272_), .Y(new_n11176_));
  NOR3X1   g10983(.A(new_n11176_), .B(new_n4354_), .C(new_n3460_), .Y(new_n11177_));
  AOI21X1  g10984(.A0(new_n4484_), .A1(new_n4272_), .B0(new_n11176_), .Y(new_n11178_));
  OAI22X1  g10985(.A0(new_n4349_), .A1(new_n4041_), .B0(new_n4983_), .B1(new_n3926_), .Y(new_n11179_));
  AOI21X1  g10986(.A0(new_n11179_), .A1(new_n11178_), .B0(new_n11177_), .Y(new_n11180_));
  XOR2X1   g10987(.A(new_n11180_), .B(new_n11173_), .Y(new_n11181_));
  INVX1    g10988(.A(new_n11078_), .Y(new_n11182_));
  AOI22X1  g10989(.A0(\a[62] ), .A1(\a[36] ), .B0(\a[61] ), .B1(\a[37] ), .Y(new_n11183_));
  AOI21X1  g10990(.A0(new_n6556_), .A1(new_n3330_), .B0(new_n11183_), .Y(new_n11184_));
  XOR2X1   g10991(.A(new_n11184_), .B(new_n11182_), .Y(new_n11185_));
  INVX1    g10992(.A(new_n11185_), .Y(new_n11186_));
  XOR2X1   g10993(.A(new_n11186_), .B(new_n11181_), .Y(new_n11187_));
  XOR2X1   g10994(.A(new_n11187_), .B(new_n11164_), .Y(new_n11188_));
  NOR2X1   g10995(.A(new_n11188_), .B(new_n11159_), .Y(new_n11189_));
  XOR2X1   g10996(.A(new_n11188_), .B(new_n11159_), .Y(new_n11190_));
  NAND2X1  g10997(.A(new_n11188_), .B(new_n11159_), .Y(new_n11191_));
  OAI21X1  g10998(.A0(new_n11189_), .A1(new_n11150_), .B0(new_n11191_), .Y(new_n11192_));
  OAI22X1  g10999(.A0(new_n11192_), .A1(new_n11189_), .B0(new_n11190_), .B1(new_n11150_), .Y(new_n11193_));
  NOR2X1   g11000(.A(new_n11097_), .B(new_n11094_), .Y(new_n11194_));
  AOI21X1  g11001(.A0(new_n11098_), .A1(new_n11092_), .B0(new_n11194_), .Y(new_n11195_));
  INVX1    g11002(.A(new_n11087_), .Y(new_n11196_));
  AOI22X1  g11003(.A0(\a[55] ), .A1(\a[43] ), .B0(\a[54] ), .B1(\a[44] ), .Y(new_n11197_));
  AOI21X1  g11004(.A0(new_n5240_), .A1(new_n4992_), .B0(new_n11197_), .Y(new_n11198_));
  AND2X1   g11005(.A(\a[63] ), .B(\a[35] ), .Y(new_n11199_));
  XOR2X1   g11006(.A(new_n11199_), .B(new_n11198_), .Y(new_n11200_));
  XOR2X1   g11007(.A(new_n11200_), .B(new_n11196_), .Y(new_n11201_));
  AND2X1   g11008(.A(\a[60] ), .B(\a[38] ), .Y(new_n11202_));
  AOI22X1  g11009(.A0(\a[57] ), .A1(\a[41] ), .B0(\a[56] ), .B1(\a[42] ), .Y(new_n11203_));
  INVX1    g11010(.A(new_n11203_), .Y(new_n11204_));
  NAND4X1  g11011(.A(\a[57] ), .B(\a[56] ), .C(\a[42] ), .D(\a[41] ), .Y(new_n11205_));
  NAND3X1  g11012(.A(new_n11204_), .B(new_n11205_), .C(new_n11202_), .Y(new_n11206_));
  AOI22X1  g11013(.A0(new_n11204_), .A1(new_n11202_), .B0(new_n5554_), .B1(new_n3607_), .Y(new_n11207_));
  AOI22X1  g11014(.A0(new_n11207_), .A1(new_n11204_), .B0(new_n11206_), .B1(new_n11202_), .Y(new_n11208_));
  XOR2X1   g11015(.A(new_n11208_), .B(new_n11201_), .Y(new_n11209_));
  AND2X1   g11016(.A(new_n11039_), .B(new_n11036_), .Y(new_n11210_));
  OAI21X1  g11017(.A0(new_n11210_), .A1(new_n11073_), .B0(new_n11072_), .Y(new_n11211_));
  OAI21X1  g11018(.A0(new_n11075_), .A1(new_n11069_), .B0(new_n11211_), .Y(new_n11212_));
  AND2X1   g11019(.A(new_n11212_), .B(new_n11209_), .Y(new_n11213_));
  XOR2X1   g11020(.A(new_n11212_), .B(new_n11209_), .Y(new_n11214_));
  OAI21X1  g11021(.A0(new_n11212_), .A1(new_n11209_), .B0(new_n11195_), .Y(new_n11215_));
  OAI22X1  g11022(.A0(new_n11215_), .A1(new_n11213_), .B0(new_n11214_), .B1(new_n11195_), .Y(new_n11216_));
  AND2X1   g11023(.A(new_n11099_), .B(new_n11076_), .Y(new_n11217_));
  INVX1    g11024(.A(new_n11217_), .Y(new_n11218_));
  OAI21X1  g11025(.A0(new_n11065_), .A1(new_n11063_), .B0(new_n11100_), .Y(new_n11219_));
  AOI21X1  g11026(.A0(new_n11219_), .A1(new_n11218_), .B0(new_n11216_), .Y(new_n11220_));
  OR2X1    g11027(.A(new_n11220_), .B(new_n11216_), .Y(new_n11221_));
  AND2X1   g11028(.A(new_n11219_), .B(new_n11218_), .Y(new_n11222_));
  XOR2X1   g11029(.A(new_n11216_), .B(new_n11222_), .Y(new_n11223_));
  NOR2X1   g11030(.A(new_n11220_), .B(new_n11222_), .Y(new_n11224_));
  NOR2X1   g11031(.A(new_n11224_), .B(new_n11193_), .Y(new_n11225_));
  AOI22X1  g11032(.A0(new_n11225_), .A1(new_n11221_), .B0(new_n11223_), .B1(new_n11193_), .Y(new_n11226_));
  XOR2X1   g11033(.A(new_n11226_), .B(new_n11148_), .Y(new_n11227_));
  INVX1    g11034(.A(new_n11143_), .Y(new_n11228_));
  OAI21X1  g11035(.A0(new_n11144_), .A1(new_n11060_), .B0(new_n11228_), .Y(new_n11229_));
  XOR2X1   g11036(.A(new_n11229_), .B(new_n11227_), .Y(\asquared[99] ));
  AOI21X1  g11037(.A0(new_n11223_), .A1(new_n11193_), .B0(new_n11220_), .Y(new_n11231_));
  AOI22X1  g11038(.A0(\a[58] ), .A1(\a[41] ), .B0(\a[55] ), .B1(\a[44] ), .Y(new_n11232_));
  NOR4X1   g11039(.A(new_n5379_), .B(new_n4906_), .C(new_n5268_), .D(new_n3081_), .Y(new_n11233_));
  NAND4X1  g11040(.A(\a[59] ), .B(\a[58] ), .C(\a[41] ), .D(\a[40] ), .Y(new_n11234_));
  NAND4X1  g11041(.A(\a[59] ), .B(\a[55] ), .C(\a[44] ), .D(\a[40] ), .Y(new_n11235_));
  AOI21X1  g11042(.A0(new_n11235_), .A1(new_n11234_), .B0(new_n11233_), .Y(new_n11236_));
  NOR2X1   g11043(.A(new_n11236_), .B(new_n11233_), .Y(new_n11237_));
  INVX1    g11044(.A(new_n11237_), .Y(new_n11238_));
  NAND2X1  g11045(.A(\a[59] ), .B(\a[40] ), .Y(new_n11239_));
  OAI22X1  g11046(.A0(new_n11239_), .A1(new_n11236_), .B0(new_n11238_), .B1(new_n11232_), .Y(new_n11240_));
  NAND4X1  g11047(.A(\a[54] ), .B(\a[52] ), .C(\a[47] ), .D(\a[45] ), .Y(new_n11241_));
  NAND4X1  g11048(.A(\a[54] ), .B(\a[53] ), .C(\a[46] ), .D(\a[45] ), .Y(new_n11242_));
  AOI22X1  g11049(.A0(new_n11242_), .A1(new_n11241_), .B0(new_n5048_), .B1(new_n3893_), .Y(new_n11243_));
  NAND2X1  g11050(.A(\a[54] ), .B(\a[45] ), .Y(new_n11244_));
  NAND4X1  g11051(.A(\a[53] ), .B(\a[52] ), .C(\a[47] ), .D(\a[46] ), .Y(new_n11245_));
  NAND3X1  g11052(.A(new_n11242_), .B(new_n11241_), .C(new_n11245_), .Y(new_n11246_));
  AOI22X1  g11053(.A0(\a[53] ), .A1(\a[46] ), .B0(\a[52] ), .B1(\a[47] ), .Y(new_n11247_));
  OAI22X1  g11054(.A0(new_n11247_), .A1(new_n11246_), .B0(new_n11244_), .B1(new_n11243_), .Y(new_n11248_));
  XOR2X1   g11055(.A(new_n11248_), .B(new_n11240_), .Y(new_n11249_));
  AOI22X1  g11056(.A0(\a[57] ), .A1(\a[42] ), .B0(\a[56] ), .B1(\a[43] ), .Y(new_n11250_));
  AND2X1   g11057(.A(\a[51] ), .B(\a[48] ), .Y(new_n11251_));
  AND2X1   g11058(.A(new_n5554_), .B(new_n3462_), .Y(new_n11252_));
  OAI21X1  g11059(.A0(new_n11250_), .A1(new_n11252_), .B0(new_n11251_), .Y(new_n11253_));
  INVX1    g11060(.A(new_n11250_), .Y(new_n11254_));
  AOI21X1  g11061(.A0(new_n11254_), .A1(new_n11251_), .B0(new_n11252_), .Y(new_n11255_));
  INVX1    g11062(.A(new_n11255_), .Y(new_n11256_));
  OAI21X1  g11063(.A0(new_n11256_), .A1(new_n11250_), .B0(new_n11253_), .Y(new_n11257_));
  XOR2X1   g11064(.A(new_n11257_), .B(new_n11249_), .Y(new_n11258_));
  OR2X1    g11065(.A(new_n11154_), .B(new_n11152_), .Y(new_n11259_));
  OAI21X1  g11066(.A0(new_n11158_), .A1(new_n11156_), .B0(new_n11259_), .Y(new_n11260_));
  XOR2X1   g11067(.A(new_n11260_), .B(new_n11258_), .Y(new_n11261_));
  INVX1    g11068(.A(new_n11261_), .Y(new_n11262_));
  NOR2X1   g11069(.A(new_n11163_), .B(new_n11161_), .Y(new_n11263_));
  AOI21X1  g11070(.A0(new_n11187_), .A1(new_n11164_), .B0(new_n11263_), .Y(new_n11264_));
  XOR2X1   g11071(.A(new_n11264_), .B(new_n11262_), .Y(new_n11265_));
  INVX1    g11072(.A(new_n11265_), .Y(new_n11266_));
  AND2X1   g11073(.A(new_n11266_), .B(new_n11192_), .Y(new_n11267_));
  INVX1    g11074(.A(new_n11209_), .Y(new_n11268_));
  AND2X1   g11075(.A(new_n11212_), .B(new_n11268_), .Y(new_n11269_));
  NOR2X1   g11076(.A(new_n11214_), .B(new_n11195_), .Y(new_n11270_));
  OR2X1    g11077(.A(new_n11270_), .B(new_n11269_), .Y(new_n11271_));
  AND2X1   g11078(.A(new_n11118_), .B(new_n11110_), .Y(new_n11272_));
  AOI21X1  g11079(.A0(new_n11160_), .A1(new_n11129_), .B0(new_n11272_), .Y(new_n11273_));
  AND2X1   g11080(.A(\a[62] ), .B(\a[50] ), .Y(new_n11274_));
  AOI21X1  g11081(.A0(new_n11274_), .A1(\a[37] ), .B0(new_n7652_), .Y(new_n11275_));
  AOI21X1  g11082(.A0(new_n11274_), .A1(\a[37] ), .B0(new_n4321_), .Y(new_n11276_));
  INVX1    g11083(.A(new_n11276_), .Y(new_n11277_));
  AOI21X1  g11084(.A0(\a[62] ), .A1(\a[37] ), .B0(\a[50] ), .Y(new_n11278_));
  OAI22X1  g11085(.A0(new_n11278_), .A1(new_n11277_), .B0(new_n11275_), .B1(new_n7652_), .Y(new_n11279_));
  XOR2X1   g11086(.A(new_n11279_), .B(new_n11273_), .Y(new_n11280_));
  INVX1    g11087(.A(new_n11201_), .Y(new_n11281_));
  NOR2X1   g11088(.A(new_n11208_), .B(new_n11281_), .Y(new_n11282_));
  AOI21X1  g11089(.A0(new_n11200_), .A1(new_n11196_), .B0(new_n11282_), .Y(new_n11283_));
  XOR2X1   g11090(.A(new_n11283_), .B(new_n11280_), .Y(new_n11284_));
  INVX1    g11091(.A(new_n11284_), .Y(new_n11285_));
  AOI22X1  g11092(.A0(new_n11184_), .A1(new_n11182_), .B0(new_n6556_), .B1(new_n3330_), .Y(new_n11286_));
  XOR2X1   g11093(.A(new_n11286_), .B(new_n11207_), .Y(new_n11287_));
  NAND4X1  g11094(.A(\a[63] ), .B(\a[60] ), .C(\a[39] ), .D(\a[36] ), .Y(new_n11288_));
  OAI21X1  g11095(.A0(new_n7973_), .A1(new_n7316_), .B0(new_n11288_), .Y(new_n11289_));
  OAI21X1  g11096(.A0(new_n6554_), .A1(new_n3729_), .B0(new_n11289_), .Y(new_n11290_));
  AND2X1   g11097(.A(\a[63] ), .B(\a[36] ), .Y(new_n11291_));
  AOI21X1  g11098(.A0(new_n6428_), .A1(new_n3503_), .B0(new_n11289_), .Y(new_n11292_));
  OAI22X1  g11099(.A0(new_n6023_), .A1(new_n2519_), .B0(new_n5952_), .B1(new_n2652_), .Y(new_n11293_));
  AOI22X1  g11100(.A0(new_n11293_), .A1(new_n11292_), .B0(new_n11291_), .B1(new_n11290_), .Y(new_n11294_));
  XOR2X1   g11101(.A(new_n11294_), .B(new_n11287_), .Y(new_n11295_));
  XOR2X1   g11102(.A(new_n11178_), .B(new_n11171_), .Y(new_n11296_));
  INVX1    g11103(.A(new_n11199_), .Y(new_n11297_));
  OAI22X1  g11104(.A0(new_n11297_), .A1(new_n11197_), .B0(new_n5241_), .B1(new_n7353_), .Y(new_n11298_));
  XOR2X1   g11105(.A(new_n11298_), .B(new_n11296_), .Y(new_n11299_));
  AND2X1   g11106(.A(new_n11179_), .B(new_n11178_), .Y(new_n11300_));
  OAI21X1  g11107(.A0(new_n11300_), .A1(new_n11177_), .B0(new_n11173_), .Y(new_n11301_));
  OAI21X1  g11108(.A0(new_n11186_), .A1(new_n11181_), .B0(new_n11301_), .Y(new_n11302_));
  XOR2X1   g11109(.A(new_n11302_), .B(new_n11299_), .Y(new_n11303_));
  XOR2X1   g11110(.A(new_n11303_), .B(new_n11295_), .Y(new_n11304_));
  XOR2X1   g11111(.A(new_n11304_), .B(new_n11285_), .Y(new_n11305_));
  XOR2X1   g11112(.A(new_n11305_), .B(new_n11271_), .Y(new_n11306_));
  NOR2X1   g11113(.A(new_n11266_), .B(new_n11192_), .Y(new_n11307_));
  OAI21X1  g11114(.A0(new_n11267_), .A1(new_n11307_), .B0(new_n11306_), .Y(new_n11308_));
  OR2X1    g11115(.A(new_n11307_), .B(new_n11306_), .Y(new_n11309_));
  OAI21X1  g11116(.A0(new_n11309_), .A1(new_n11267_), .B0(new_n11308_), .Y(new_n11310_));
  NOR2X1   g11117(.A(new_n11310_), .B(new_n11231_), .Y(new_n11311_));
  AND2X1   g11118(.A(new_n11310_), .B(new_n11231_), .Y(new_n11312_));
  OR2X1    g11119(.A(new_n11312_), .B(new_n11311_), .Y(new_n11313_));
  NOR2X1   g11120(.A(new_n11226_), .B(new_n11148_), .Y(new_n11314_));
  INVX1    g11121(.A(new_n11314_), .Y(new_n11315_));
  AND2X1   g11122(.A(new_n11226_), .B(new_n11148_), .Y(new_n11316_));
  AOI21X1  g11123(.A0(new_n11229_), .A1(new_n11315_), .B0(new_n11316_), .Y(new_n11317_));
  XOR2X1   g11124(.A(new_n11317_), .B(new_n11313_), .Y(\asquared[100] ));
  INVX1    g11125(.A(new_n11308_), .Y(new_n11319_));
  AOI21X1  g11126(.A0(new_n11265_), .A1(new_n11192_), .B0(new_n11319_), .Y(new_n11320_));
  INVX1    g11127(.A(new_n11320_), .Y(new_n11321_));
  NOR2X1   g11128(.A(new_n11178_), .B(new_n11171_), .Y(new_n11322_));
  AOI21X1  g11129(.A0(new_n11298_), .A1(new_n11296_), .B0(new_n11322_), .Y(new_n11323_));
  OAI22X1  g11130(.A0(new_n7336_), .A1(new_n8297_), .B0(new_n8145_), .B1(new_n4279_), .Y(new_n11324_));
  OAI21X1  g11131(.A0(new_n7793_), .A1(new_n4280_), .B0(new_n11324_), .Y(new_n11325_));
  AND2X1   g11132(.A(\a[53] ), .B(\a[47] ), .Y(new_n11326_));
  AOI21X1  g11133(.A0(new_n7164_), .A1(new_n4274_), .B0(new_n11324_), .Y(new_n11327_));
  OAI21X1  g11134(.A0(new_n4354_), .A1(new_n3926_), .B0(new_n7653_), .Y(new_n11328_));
  AOI22X1  g11135(.A0(new_n11328_), .A1(new_n11327_), .B0(new_n11326_), .B1(new_n11325_), .Y(new_n11329_));
  XOR2X1   g11136(.A(new_n11329_), .B(new_n11323_), .Y(new_n11330_));
  AND2X1   g11137(.A(new_n11286_), .B(new_n11207_), .Y(new_n11331_));
  OR2X1    g11138(.A(new_n11286_), .B(new_n11207_), .Y(new_n11332_));
  OAI21X1  g11139(.A0(new_n11294_), .A1(new_n11331_), .B0(new_n11332_), .Y(new_n11333_));
  XOR2X1   g11140(.A(new_n11333_), .B(new_n11330_), .Y(new_n11334_));
  NAND2X1  g11141(.A(new_n11260_), .B(new_n11258_), .Y(new_n11335_));
  OAI21X1  g11142(.A0(new_n11264_), .A1(new_n11262_), .B0(new_n11335_), .Y(new_n11336_));
  XOR2X1   g11143(.A(new_n11336_), .B(new_n11334_), .Y(new_n11337_));
  INVX1    g11144(.A(new_n11292_), .Y(new_n11338_));
  XOR2X1   g11145(.A(new_n11246_), .B(new_n11338_), .Y(new_n11339_));
  XOR2X1   g11146(.A(new_n11339_), .B(new_n11237_), .Y(new_n11340_));
  AND2X1   g11147(.A(new_n11248_), .B(new_n11240_), .Y(new_n11341_));
  AOI21X1  g11148(.A0(new_n11257_), .A1(new_n11249_), .B0(new_n11341_), .Y(new_n11342_));
  XOR2X1   g11149(.A(new_n11342_), .B(new_n11340_), .Y(new_n11343_));
  AND2X1   g11150(.A(\a[63] ), .B(\a[37] ), .Y(new_n11344_));
  XOR2X1   g11151(.A(new_n11344_), .B(new_n11277_), .Y(new_n11345_));
  XOR2X1   g11152(.A(new_n11345_), .B(new_n11256_), .Y(new_n11346_));
  XOR2X1   g11153(.A(new_n11346_), .B(new_n11343_), .Y(new_n11347_));
  XOR2X1   g11154(.A(new_n11347_), .B(new_n11337_), .Y(new_n11348_));
  NOR2X1   g11155(.A(new_n11304_), .B(new_n11285_), .Y(new_n11349_));
  AOI21X1  g11156(.A0(new_n11305_), .A1(new_n11271_), .B0(new_n11349_), .Y(new_n11350_));
  NAND2X1  g11157(.A(\a[62] ), .B(\a[38] ), .Y(new_n11351_));
  NAND4X1  g11158(.A(\a[62] ), .B(\a[60] ), .C(\a[40] ), .D(\a[38] ), .Y(new_n11352_));
  NAND4X1  g11159(.A(\a[62] ), .B(\a[61] ), .C(\a[39] ), .D(\a[38] ), .Y(new_n11353_));
  AOI22X1  g11160(.A0(new_n11353_), .A1(new_n11352_), .B0(new_n6428_), .B1(new_n4077_), .Y(new_n11354_));
  NAND4X1  g11161(.A(\a[61] ), .B(\a[60] ), .C(\a[40] ), .D(\a[39] ), .Y(new_n11355_));
  NAND3X1  g11162(.A(new_n11353_), .B(new_n11352_), .C(new_n11355_), .Y(new_n11356_));
  AOI22X1  g11163(.A0(\a[61] ), .A1(\a[39] ), .B0(\a[60] ), .B1(\a[40] ), .Y(new_n11357_));
  OAI22X1  g11164(.A0(new_n11357_), .A1(new_n11356_), .B0(new_n11354_), .B1(new_n11351_), .Y(new_n11358_));
  NAND2X1  g11165(.A(\a[57] ), .B(\a[43] ), .Y(new_n11359_));
  NAND4X1  g11166(.A(\a[57] ), .B(\a[55] ), .C(\a[45] ), .D(\a[43] ), .Y(new_n11360_));
  NAND4X1  g11167(.A(\a[57] ), .B(\a[56] ), .C(\a[44] ), .D(\a[43] ), .Y(new_n11361_));
  AOI22X1  g11168(.A0(new_n11361_), .A1(new_n11360_), .B0(new_n6237_), .B1(new_n3918_), .Y(new_n11362_));
  AOI22X1  g11169(.A0(\a[56] ), .A1(\a[44] ), .B0(\a[55] ), .B1(\a[45] ), .Y(new_n11363_));
  AOI21X1  g11170(.A0(new_n6237_), .A1(new_n3918_), .B0(new_n11362_), .Y(new_n11364_));
  INVX1    g11171(.A(new_n11364_), .Y(new_n11365_));
  OAI22X1  g11172(.A0(new_n11365_), .A1(new_n11363_), .B0(new_n11362_), .B1(new_n11359_), .Y(new_n11366_));
  XOR2X1   g11173(.A(new_n11366_), .B(new_n11358_), .Y(new_n11367_));
  INVX1    g11174(.A(new_n6371_), .Y(new_n11368_));
  AOI22X1  g11175(.A0(\a[59] ), .A1(\a[41] ), .B0(\a[58] ), .B1(\a[42] ), .Y(new_n11369_));
  AND2X1   g11176(.A(new_n6121_), .B(new_n3607_), .Y(new_n11370_));
  NOR3X1   g11177(.A(new_n11369_), .B(new_n11370_), .C(new_n11368_), .Y(new_n11371_));
  NOR2X1   g11178(.A(new_n11371_), .B(new_n11370_), .Y(new_n11372_));
  INVX1    g11179(.A(new_n11372_), .Y(new_n11373_));
  OAI22X1  g11180(.A0(new_n11373_), .A1(new_n11369_), .B0(new_n11371_), .B1(new_n11368_), .Y(new_n11374_));
  XOR2X1   g11181(.A(new_n11374_), .B(new_n11367_), .Y(new_n11375_));
  INVX1    g11182(.A(new_n11375_), .Y(new_n11376_));
  INVX1    g11183(.A(new_n11279_), .Y(new_n11377_));
  OR2X1    g11184(.A(new_n11377_), .B(new_n11273_), .Y(new_n11378_));
  OR2X1    g11185(.A(new_n11283_), .B(new_n11280_), .Y(new_n11379_));
  AND2X1   g11186(.A(new_n11379_), .B(new_n11378_), .Y(new_n11380_));
  XOR2X1   g11187(.A(new_n11380_), .B(new_n11376_), .Y(new_n11381_));
  INVX1    g11188(.A(new_n11295_), .Y(new_n11382_));
  AND2X1   g11189(.A(new_n11302_), .B(new_n11299_), .Y(new_n11383_));
  AOI21X1  g11190(.A0(new_n11303_), .A1(new_n11382_), .B0(new_n11383_), .Y(new_n11384_));
  XOR2X1   g11191(.A(new_n11384_), .B(new_n11381_), .Y(new_n11385_));
  XOR2X1   g11192(.A(new_n11385_), .B(new_n11350_), .Y(new_n11386_));
  XOR2X1   g11193(.A(new_n11386_), .B(new_n11348_), .Y(new_n11387_));
  AND2X1   g11194(.A(new_n11387_), .B(new_n11321_), .Y(new_n11388_));
  INVX1    g11195(.A(new_n11388_), .Y(new_n11389_));
  INVX1    g11196(.A(new_n11311_), .Y(new_n11390_));
  OAI21X1  g11197(.A0(new_n11317_), .A1(new_n11312_), .B0(new_n11390_), .Y(new_n11391_));
  OR2X1    g11198(.A(new_n11387_), .B(new_n11321_), .Y(new_n11392_));
  AOI21X1  g11199(.A0(new_n11392_), .A1(new_n11389_), .B0(new_n11391_), .Y(new_n11393_));
  AND2X1   g11200(.A(new_n11392_), .B(new_n11391_), .Y(new_n11394_));
  AOI21X1  g11201(.A0(new_n11394_), .A1(new_n11389_), .B0(new_n11393_), .Y(\asquared[101] ));
  AOI21X1  g11202(.A0(new_n11392_), .A1(new_n11391_), .B0(new_n11388_), .Y(new_n11396_));
  NOR2X1   g11203(.A(new_n11385_), .B(new_n11350_), .Y(new_n11397_));
  AOI21X1  g11204(.A0(new_n11386_), .A1(new_n11348_), .B0(new_n11397_), .Y(new_n11398_));
  AND2X1   g11205(.A(new_n11336_), .B(new_n11334_), .Y(new_n11399_));
  AOI21X1  g11206(.A0(new_n11347_), .A1(new_n11337_), .B0(new_n11399_), .Y(new_n11400_));
  AOI22X1  g11207(.A0(\a[55] ), .A1(\a[46] ), .B0(\a[54] ), .B1(\a[47] ), .Y(new_n11401_));
  AND2X1   g11208(.A(\a[63] ), .B(\a[38] ), .Y(new_n11402_));
  INVX1    g11209(.A(new_n11402_), .Y(new_n11403_));
  AND2X1   g11210(.A(new_n5240_), .B(new_n3893_), .Y(new_n11404_));
  NOR3X1   g11211(.A(new_n11403_), .B(new_n11404_), .C(new_n11401_), .Y(new_n11405_));
  NOR2X1   g11212(.A(new_n11405_), .B(new_n11404_), .Y(new_n11406_));
  INVX1    g11213(.A(new_n11406_), .Y(new_n11407_));
  OAI22X1  g11214(.A0(new_n11407_), .A1(new_n11401_), .B0(new_n11405_), .B1(new_n11403_), .Y(new_n11408_));
  NAND4X1  g11215(.A(\a[59] ), .B(\a[56] ), .C(\a[45] ), .D(\a[42] ), .Y(new_n11409_));
  NAND4X1  g11216(.A(\a[59] ), .B(\a[58] ), .C(\a[43] ), .D(\a[42] ), .Y(new_n11410_));
  AOI22X1  g11217(.A0(new_n11410_), .A1(new_n11409_), .B0(new_n5381_), .B1(new_n7640_), .Y(new_n11411_));
  NOR3X1   g11218(.A(new_n11411_), .B(new_n5617_), .C(new_n3096_), .Y(new_n11412_));
  AOI21X1  g11219(.A0(new_n5381_), .A1(new_n7640_), .B0(new_n11411_), .Y(new_n11413_));
  OAI22X1  g11220(.A0(new_n5379_), .A1(new_n3037_), .B0(new_n6022_), .B1(new_n3811_), .Y(new_n11414_));
  AOI21X1  g11221(.A0(new_n11414_), .A1(new_n11413_), .B0(new_n11412_), .Y(new_n11415_));
  XOR2X1   g11222(.A(new_n11415_), .B(new_n11408_), .Y(new_n11416_));
  INVX1    g11223(.A(new_n11416_), .Y(new_n11417_));
  NOR4X1   g11224(.A(new_n5441_), .B(new_n4354_), .C(new_n3915_), .D(new_n5268_), .Y(new_n11418_));
  AND2X1   g11225(.A(\a[57] ), .B(\a[44] ), .Y(new_n11419_));
  AOI22X1  g11226(.A0(new_n11419_), .A1(new_n7095_), .B0(new_n5048_), .B1(new_n4274_), .Y(new_n11420_));
  NOR2X1   g11227(.A(new_n11420_), .B(new_n11418_), .Y(new_n11421_));
  NOR3X1   g11228(.A(new_n11421_), .B(new_n5245_), .C(new_n3926_), .Y(new_n11422_));
  NOR2X1   g11229(.A(new_n11421_), .B(new_n11418_), .Y(new_n11423_));
  OAI22X1  g11230(.A0(new_n5441_), .A1(new_n5268_), .B0(new_n4354_), .B1(new_n3915_), .Y(new_n11424_));
  AOI21X1  g11231(.A0(new_n11424_), .A1(new_n11423_), .B0(new_n11422_), .Y(new_n11425_));
  XOR2X1   g11232(.A(new_n11425_), .B(new_n11417_), .Y(new_n11426_));
  NOR2X1   g11233(.A(new_n11329_), .B(new_n11323_), .Y(new_n11427_));
  AOI21X1  g11234(.A0(new_n11333_), .A1(new_n11330_), .B0(new_n11427_), .Y(new_n11428_));
  XOR2X1   g11235(.A(new_n11428_), .B(new_n11426_), .Y(new_n11429_));
  NAND2X1  g11236(.A(new_n11344_), .B(new_n11277_), .Y(new_n11430_));
  NOR2X1   g11237(.A(new_n11344_), .B(new_n11277_), .Y(new_n11431_));
  OAI21X1  g11238(.A0(new_n11431_), .A1(new_n11255_), .B0(new_n11430_), .Y(new_n11432_));
  NAND2X1  g11239(.A(\a[60] ), .B(\a[41] ), .Y(new_n11433_));
  NAND2X1  g11240(.A(\a[61] ), .B(\a[40] ), .Y(new_n11434_));
  AOI22X1  g11241(.A0(new_n11434_), .A1(new_n11433_), .B0(new_n6428_), .B1(new_n4404_), .Y(new_n11435_));
  XOR2X1   g11242(.A(new_n11435_), .B(new_n11327_), .Y(new_n11436_));
  AOI21X1  g11243(.A0(new_n5290_), .A1(\a[62] ), .B0(new_n4484_), .Y(new_n11437_));
  OAI21X1  g11244(.A0(new_n6606_), .A1(new_n2652_), .B0(new_n4349_), .Y(new_n11438_));
  NOR4X1   g11245(.A(new_n6606_), .B(new_n4349_), .C(new_n4983_), .D(new_n2652_), .Y(new_n11439_));
  AOI21X1  g11246(.A0(new_n11438_), .A1(new_n11437_), .B0(new_n11439_), .Y(new_n11440_));
  XOR2X1   g11247(.A(new_n11440_), .B(new_n11436_), .Y(new_n11441_));
  XOR2X1   g11248(.A(new_n11441_), .B(new_n11432_), .Y(new_n11442_));
  XOR2X1   g11249(.A(new_n11442_), .B(new_n11429_), .Y(new_n11443_));
  XOR2X1   g11250(.A(new_n11443_), .B(new_n11400_), .Y(new_n11444_));
  AOI21X1  g11251(.A0(new_n11379_), .A1(new_n11378_), .B0(new_n11376_), .Y(new_n11445_));
  INVX1    g11252(.A(new_n11445_), .Y(new_n11446_));
  INVX1    g11253(.A(new_n11381_), .Y(new_n11447_));
  OAI21X1  g11254(.A0(new_n11384_), .A1(new_n11447_), .B0(new_n11446_), .Y(new_n11448_));
  NOR2X1   g11255(.A(new_n11342_), .B(new_n11340_), .Y(new_n11449_));
  AOI21X1  g11256(.A0(new_n11346_), .A1(new_n11343_), .B0(new_n11449_), .Y(new_n11450_));
  XOR2X1   g11257(.A(new_n11450_), .B(new_n11448_), .Y(new_n11451_));
  XOR2X1   g11258(.A(new_n11373_), .B(new_n11356_), .Y(new_n11452_));
  XOR2X1   g11259(.A(new_n11452_), .B(new_n11365_), .Y(new_n11453_));
  AND2X1   g11260(.A(new_n11366_), .B(new_n11358_), .Y(new_n11454_));
  AOI21X1  g11261(.A0(new_n11374_), .A1(new_n11367_), .B0(new_n11454_), .Y(new_n11455_));
  AND2X1   g11262(.A(new_n11246_), .B(new_n11338_), .Y(new_n11456_));
  AOI21X1  g11263(.A0(new_n11339_), .A1(new_n11238_), .B0(new_n11456_), .Y(new_n11457_));
  XOR2X1   g11264(.A(new_n11457_), .B(new_n11455_), .Y(new_n11458_));
  XOR2X1   g11265(.A(new_n11458_), .B(new_n11453_), .Y(new_n11459_));
  XOR2X1   g11266(.A(new_n11459_), .B(new_n11451_), .Y(new_n11460_));
  INVX1    g11267(.A(new_n11460_), .Y(new_n11461_));
  XOR2X1   g11268(.A(new_n11461_), .B(new_n11444_), .Y(new_n11462_));
  NOR2X1   g11269(.A(new_n11462_), .B(new_n11398_), .Y(new_n11463_));
  AND2X1   g11270(.A(new_n11462_), .B(new_n11398_), .Y(new_n11464_));
  OR2X1    g11271(.A(new_n11464_), .B(new_n11463_), .Y(new_n11465_));
  XOR2X1   g11272(.A(new_n11465_), .B(new_n11396_), .Y(\asquared[102] ));
  INVX1    g11273(.A(new_n11443_), .Y(new_n11467_));
  OR2X1    g11274(.A(new_n11467_), .B(new_n11400_), .Y(new_n11468_));
  OAI21X1  g11275(.A0(new_n11460_), .A1(new_n11444_), .B0(new_n11468_), .Y(new_n11469_));
  AND2X1   g11276(.A(new_n11346_), .B(new_n11343_), .Y(new_n11470_));
  OAI21X1  g11277(.A0(new_n11470_), .A1(new_n11449_), .B0(new_n11448_), .Y(new_n11471_));
  INVX1    g11278(.A(new_n11459_), .Y(new_n11472_));
  OAI21X1  g11279(.A0(new_n11472_), .A1(new_n11451_), .B0(new_n11471_), .Y(new_n11473_));
  INVX1    g11280(.A(new_n11327_), .Y(new_n11474_));
  AOI22X1  g11281(.A0(new_n11435_), .A1(new_n11474_), .B0(new_n6428_), .B1(new_n4404_), .Y(new_n11475_));
  XOR2X1   g11282(.A(new_n11475_), .B(new_n11413_), .Y(new_n11476_));
  NAND4X1  g11283(.A(\a[63] ), .B(\a[60] ), .C(\a[42] ), .D(\a[39] ), .Y(new_n11477_));
  NAND4X1  g11284(.A(\a[63] ), .B(\a[61] ), .C(\a[41] ), .D(\a[39] ), .Y(new_n11478_));
  AOI22X1  g11285(.A0(new_n11478_), .A1(new_n11477_), .B0(new_n6428_), .B1(new_n3607_), .Y(new_n11479_));
  NOR3X1   g11286(.A(new_n11479_), .B(new_n6549_), .C(new_n2652_), .Y(new_n11480_));
  AOI21X1  g11287(.A0(new_n6428_), .A1(new_n3607_), .B0(new_n11479_), .Y(new_n11481_));
  OAI22X1  g11288(.A0(new_n6023_), .A1(new_n3081_), .B0(new_n5952_), .B1(new_n3096_), .Y(new_n11482_));
  AOI21X1  g11289(.A0(new_n11482_), .A1(new_n11481_), .B0(new_n11480_), .Y(new_n11483_));
  XOR2X1   g11290(.A(new_n11483_), .B(new_n11476_), .Y(new_n11484_));
  NOR2X1   g11291(.A(new_n11440_), .B(new_n11436_), .Y(new_n11485_));
  AOI21X1  g11292(.A0(new_n11441_), .A1(new_n11432_), .B0(new_n11485_), .Y(new_n11486_));
  XOR2X1   g11293(.A(new_n11486_), .B(new_n11484_), .Y(new_n11487_));
  INVX1    g11294(.A(new_n8993_), .Y(new_n11488_));
  AOI22X1  g11295(.A0(\a[59] ), .A1(\a[43] ), .B0(\a[58] ), .B1(\a[44] ), .Y(new_n11489_));
  AND2X1   g11296(.A(new_n6121_), .B(new_n4992_), .Y(new_n11490_));
  NOR3X1   g11297(.A(new_n11490_), .B(new_n11489_), .C(new_n11488_), .Y(new_n11491_));
  INVX1    g11298(.A(new_n11489_), .Y(new_n11492_));
  AOI21X1  g11299(.A0(new_n11492_), .A1(new_n8993_), .B0(new_n11490_), .Y(new_n11493_));
  INVX1    g11300(.A(new_n11493_), .Y(new_n11494_));
  OAI22X1  g11301(.A0(new_n11494_), .A1(new_n11489_), .B0(new_n11491_), .B1(new_n11488_), .Y(new_n11495_));
  INVX1    g11302(.A(new_n5554_), .Y(new_n11496_));
  NAND4X1  g11303(.A(\a[57] ), .B(\a[55] ), .C(\a[47] ), .D(\a[45] ), .Y(new_n11497_));
  OAI21X1  g11304(.A0(new_n11496_), .A1(new_n8873_), .B0(new_n11497_), .Y(new_n11498_));
  OAI21X1  g11305(.A0(new_n8560_), .A1(new_n8296_), .B0(new_n11498_), .Y(new_n11499_));
  AND2X1   g11306(.A(\a[57] ), .B(\a[45] ), .Y(new_n11500_));
  OAI22X1  g11307(.A0(new_n6022_), .A1(new_n3460_), .B0(new_n4906_), .B1(new_n4041_), .Y(new_n11501_));
  AOI21X1  g11308(.A0(new_n6237_), .A1(new_n3893_), .B0(new_n11498_), .Y(new_n11502_));
  AOI22X1  g11309(.A0(new_n11502_), .A1(new_n11501_), .B0(new_n11500_), .B1(new_n11499_), .Y(new_n11503_));
  XOR2X1   g11310(.A(new_n11503_), .B(new_n11495_), .Y(new_n11504_));
  OAI22X1  g11311(.A0(new_n7338_), .A1(new_n8802_), .B0(new_n5239_), .B1(new_n4280_), .Y(new_n11505_));
  OAI21X1  g11312(.A0(new_n7336_), .A1(new_n7652_), .B0(new_n11505_), .Y(new_n11506_));
  AND2X1   g11313(.A(\a[54] ), .B(\a[48] ), .Y(new_n11507_));
  AOI21X1  g11314(.A0(new_n5048_), .A1(new_n4321_), .B0(new_n11505_), .Y(new_n11508_));
  OAI21X1  g11315(.A0(new_n5245_), .A1(new_n3915_), .B0(new_n7794_), .Y(new_n11509_));
  AOI22X1  g11316(.A0(new_n11509_), .A1(new_n11508_), .B0(new_n11507_), .B1(new_n11506_), .Y(new_n11510_));
  XOR2X1   g11317(.A(new_n11510_), .B(new_n11504_), .Y(new_n11511_));
  XOR2X1   g11318(.A(new_n11511_), .B(new_n11487_), .Y(new_n11512_));
  XOR2X1   g11319(.A(new_n11512_), .B(new_n11473_), .Y(new_n11513_));
  XOR2X1   g11320(.A(new_n11437_), .B(new_n11423_), .Y(new_n11514_));
  XOR2X1   g11321(.A(new_n11514_), .B(new_n11407_), .Y(new_n11515_));
  INVX1    g11322(.A(new_n11515_), .Y(new_n11516_));
  AND2X1   g11323(.A(new_n11373_), .B(new_n11356_), .Y(new_n11517_));
  AOI21X1  g11324(.A0(new_n11452_), .A1(new_n11365_), .B0(new_n11517_), .Y(new_n11518_));
  XOR2X1   g11325(.A(new_n11518_), .B(new_n11516_), .Y(new_n11519_));
  INVX1    g11326(.A(new_n11519_), .Y(new_n11520_));
  AND2X1   g11327(.A(new_n11414_), .B(new_n11413_), .Y(new_n11521_));
  OAI21X1  g11328(.A0(new_n11521_), .A1(new_n11412_), .B0(new_n11408_), .Y(new_n11522_));
  OAI21X1  g11329(.A0(new_n11425_), .A1(new_n11416_), .B0(new_n11522_), .Y(new_n11523_));
  XOR2X1   g11330(.A(new_n11523_), .B(new_n11520_), .Y(new_n11524_));
  NOR2X1   g11331(.A(new_n11428_), .B(new_n11426_), .Y(new_n11525_));
  AOI21X1  g11332(.A0(new_n11442_), .A1(new_n11429_), .B0(new_n11525_), .Y(new_n11526_));
  INVX1    g11333(.A(new_n11526_), .Y(new_n11527_));
  NOR2X1   g11334(.A(new_n11457_), .B(new_n11455_), .Y(new_n11528_));
  AOI21X1  g11335(.A0(new_n11458_), .A1(new_n11453_), .B0(new_n11528_), .Y(new_n11529_));
  XOR2X1   g11336(.A(new_n11529_), .B(new_n11527_), .Y(new_n11530_));
  XOR2X1   g11337(.A(new_n11530_), .B(new_n11524_), .Y(new_n11531_));
  XOR2X1   g11338(.A(new_n11531_), .B(new_n11513_), .Y(new_n11532_));
  AND2X1   g11339(.A(new_n11532_), .B(new_n11469_), .Y(new_n11533_));
  INVX1    g11340(.A(new_n11533_), .Y(new_n11534_));
  INVX1    g11341(.A(new_n11463_), .Y(new_n11535_));
  OAI21X1  g11342(.A0(new_n11464_), .A1(new_n11396_), .B0(new_n11535_), .Y(new_n11536_));
  NOR2X1   g11343(.A(new_n11532_), .B(new_n11469_), .Y(new_n11537_));
  INVX1    g11344(.A(new_n11537_), .Y(new_n11538_));
  AOI21X1  g11345(.A0(new_n11534_), .A1(new_n11538_), .B0(new_n11536_), .Y(new_n11539_));
  AND2X1   g11346(.A(new_n11538_), .B(new_n11536_), .Y(new_n11540_));
  AOI21X1  g11347(.A0(new_n11540_), .A1(new_n11534_), .B0(new_n11539_), .Y(\asquared[103] ));
  AOI21X1  g11348(.A0(new_n11538_), .A1(new_n11536_), .B0(new_n11533_), .Y(new_n11542_));
  NOR2X1   g11349(.A(new_n11529_), .B(new_n11526_), .Y(new_n11543_));
  INVX1    g11350(.A(new_n11543_), .Y(new_n11544_));
  OAI21X1  g11351(.A0(new_n11530_), .A1(new_n11524_), .B0(new_n11544_), .Y(new_n11545_));
  AOI22X1  g11352(.A0(\a[57] ), .A1(\a[46] ), .B0(\a[56] ), .B1(\a[47] ), .Y(new_n11546_));
  AND2X1   g11353(.A(\a[60] ), .B(\a[43] ), .Y(new_n11547_));
  INVX1    g11354(.A(new_n11547_), .Y(new_n11548_));
  AND2X1   g11355(.A(new_n5554_), .B(new_n3893_), .Y(new_n11549_));
  NOR3X1   g11356(.A(new_n11548_), .B(new_n11549_), .C(new_n11546_), .Y(new_n11550_));
  INVX1    g11357(.A(new_n11546_), .Y(new_n11551_));
  AOI21X1  g11358(.A0(new_n11547_), .A1(new_n11551_), .B0(new_n11549_), .Y(new_n11552_));
  INVX1    g11359(.A(new_n11552_), .Y(new_n11553_));
  OAI22X1  g11360(.A0(new_n11553_), .A1(new_n11546_), .B0(new_n11550_), .B1(new_n11548_), .Y(new_n11554_));
  OAI22X1  g11361(.A0(new_n5241_), .A1(new_n4280_), .B0(new_n5237_), .B1(new_n8802_), .Y(new_n11555_));
  OAI21X1  g11362(.A0(new_n5239_), .A1(new_n7652_), .B0(new_n11555_), .Y(new_n11556_));
  AND2X1   g11363(.A(\a[55] ), .B(\a[48] ), .Y(new_n11557_));
  AOI21X1  g11364(.A0(new_n5238_), .A1(new_n4321_), .B0(new_n11555_), .Y(new_n11558_));
  OAI22X1  g11365(.A0(new_n4835_), .A1(new_n3915_), .B0(new_n5245_), .B1(new_n4983_), .Y(new_n11559_));
  AOI22X1  g11366(.A0(new_n11559_), .A1(new_n11558_), .B0(new_n11557_), .B1(new_n11556_), .Y(new_n11560_));
  XOR2X1   g11367(.A(new_n11560_), .B(new_n11554_), .Y(new_n11561_));
  NOR4X1   g11368(.A(new_n6606_), .B(new_n4354_), .C(new_n4349_), .D(new_n3081_), .Y(new_n11562_));
  OAI21X1  g11369(.A0(new_n9256_), .A1(\a[51] ), .B0(\a[52] ), .Y(new_n11563_));
  OR2X1    g11370(.A(new_n9256_), .B(\a[52] ), .Y(new_n11564_));
  AOI21X1  g11371(.A0(new_n11564_), .A1(new_n11563_), .B0(new_n11562_), .Y(new_n11565_));
  XOR2X1   g11372(.A(new_n11565_), .B(new_n11561_), .Y(new_n11566_));
  INVX1    g11373(.A(new_n11566_), .Y(new_n11567_));
  AND2X1   g11374(.A(\a[63] ), .B(\a[40] ), .Y(new_n11568_));
  XOR2X1   g11375(.A(new_n11568_), .B(new_n11508_), .Y(new_n11569_));
  XOR2X1   g11376(.A(new_n11569_), .B(new_n11502_), .Y(new_n11570_));
  XOR2X1   g11377(.A(new_n11493_), .B(new_n11481_), .Y(new_n11571_));
  NAND4X1  g11378(.A(\a[61] ), .B(\a[59] ), .C(\a[44] ), .D(\a[42] ), .Y(new_n11572_));
  NAND4X1  g11379(.A(\a[61] ), .B(\a[58] ), .C(\a[45] ), .D(\a[42] ), .Y(new_n11573_));
  AOI22X1  g11380(.A0(new_n11573_), .A1(new_n11572_), .B0(new_n6121_), .B1(new_n3918_), .Y(new_n11574_));
  NAND2X1  g11381(.A(\a[61] ), .B(\a[42] ), .Y(new_n11575_));
  AOI22X1  g11382(.A0(\a[59] ), .A1(\a[44] ), .B0(\a[58] ), .B1(\a[45] ), .Y(new_n11576_));
  AOI21X1  g11383(.A0(new_n6121_), .A1(new_n3918_), .B0(new_n11574_), .Y(new_n11577_));
  INVX1    g11384(.A(new_n11577_), .Y(new_n11578_));
  OAI22X1  g11385(.A0(new_n11578_), .A1(new_n11576_), .B0(new_n11575_), .B1(new_n11574_), .Y(new_n11579_));
  XOR2X1   g11386(.A(new_n11579_), .B(new_n11571_), .Y(new_n11580_));
  XOR2X1   g11387(.A(new_n11580_), .B(new_n11570_), .Y(new_n11581_));
  XOR2X1   g11388(.A(new_n11581_), .B(new_n11567_), .Y(new_n11582_));
  XOR2X1   g11389(.A(new_n11582_), .B(new_n11545_), .Y(new_n11583_));
  NOR2X1   g11390(.A(new_n11475_), .B(new_n11413_), .Y(new_n11584_));
  INVX1    g11391(.A(new_n11483_), .Y(new_n11585_));
  AOI21X1  g11392(.A0(new_n11585_), .A1(new_n11476_), .B0(new_n11584_), .Y(new_n11586_));
  NOR2X1   g11393(.A(new_n11437_), .B(new_n11423_), .Y(new_n11587_));
  AOI21X1  g11394(.A0(new_n11514_), .A1(new_n11407_), .B0(new_n11587_), .Y(new_n11588_));
  XOR2X1   g11395(.A(new_n11588_), .B(new_n11586_), .Y(new_n11589_));
  INVX1    g11396(.A(new_n11495_), .Y(new_n11590_));
  OR2X1    g11397(.A(new_n11503_), .B(new_n11590_), .Y(new_n11591_));
  OAI21X1  g11398(.A0(new_n11510_), .A1(new_n11504_), .B0(new_n11591_), .Y(new_n11592_));
  XOR2X1   g11399(.A(new_n11592_), .B(new_n11589_), .Y(new_n11593_));
  NOR2X1   g11400(.A(new_n11486_), .B(new_n11484_), .Y(new_n11594_));
  AOI21X1  g11401(.A0(new_n11511_), .A1(new_n11487_), .B0(new_n11594_), .Y(new_n11595_));
  NOR2X1   g11402(.A(new_n11518_), .B(new_n11516_), .Y(new_n11596_));
  AOI21X1  g11403(.A0(new_n11523_), .A1(new_n11519_), .B0(new_n11596_), .Y(new_n11597_));
  XOR2X1   g11404(.A(new_n11597_), .B(new_n11595_), .Y(new_n11598_));
  XOR2X1   g11405(.A(new_n11598_), .B(new_n11593_), .Y(new_n11599_));
  XOR2X1   g11406(.A(new_n11599_), .B(new_n11583_), .Y(new_n11600_));
  AND2X1   g11407(.A(new_n11512_), .B(new_n11473_), .Y(new_n11601_));
  AOI21X1  g11408(.A0(new_n11531_), .A1(new_n11513_), .B0(new_n11601_), .Y(new_n11602_));
  NOR2X1   g11409(.A(new_n11602_), .B(new_n11600_), .Y(new_n11603_));
  AND2X1   g11410(.A(new_n11602_), .B(new_n11600_), .Y(new_n11604_));
  OR2X1    g11411(.A(new_n11604_), .B(new_n11603_), .Y(new_n11605_));
  XOR2X1   g11412(.A(new_n11605_), .B(new_n11542_), .Y(\asquared[104] ));
  INVX1    g11413(.A(new_n11603_), .Y(new_n11607_));
  OAI21X1  g11414(.A0(new_n11604_), .A1(new_n11542_), .B0(new_n11607_), .Y(new_n11608_));
  XOR2X1   g11415(.A(new_n11581_), .B(new_n11566_), .Y(new_n11609_));
  AND2X1   g11416(.A(new_n11609_), .B(new_n11545_), .Y(new_n11610_));
  INVX1    g11417(.A(new_n11583_), .Y(new_n11611_));
  AOI21X1  g11418(.A0(new_n11599_), .A1(new_n11611_), .B0(new_n11610_), .Y(new_n11612_));
  NOR2X1   g11419(.A(new_n11597_), .B(new_n11595_), .Y(new_n11613_));
  AOI21X1  g11420(.A0(new_n11598_), .A1(new_n11593_), .B0(new_n11613_), .Y(new_n11614_));
  XOR2X1   g11421(.A(new_n11558_), .B(new_n11552_), .Y(new_n11615_));
  XOR2X1   g11422(.A(new_n11615_), .B(new_n11578_), .Y(new_n11616_));
  INVX1    g11423(.A(new_n11616_), .Y(new_n11617_));
  INVX1    g11424(.A(new_n11554_), .Y(new_n11618_));
  OR2X1    g11425(.A(new_n11560_), .B(new_n11618_), .Y(new_n11619_));
  OAI21X1  g11426(.A0(new_n11565_), .A1(new_n11561_), .B0(new_n11619_), .Y(new_n11620_));
  XOR2X1   g11427(.A(new_n11620_), .B(new_n11617_), .Y(new_n11621_));
  AOI22X1  g11428(.A0(\a[61] ), .A1(\a[43] ), .B0(\a[59] ), .B1(\a[45] ), .Y(new_n11622_));
  AOI22X1  g11429(.A0(new_n6428_), .A1(new_n4992_), .B0(new_n6427_), .B1(new_n3918_), .Y(new_n11623_));
  AOI21X1  g11430(.A0(new_n6020_), .A1(new_n7640_), .B0(new_n11623_), .Y(new_n11624_));
  AOI21X1  g11431(.A0(new_n6020_), .A1(new_n7640_), .B0(new_n11624_), .Y(new_n11625_));
  INVX1    g11432(.A(new_n11625_), .Y(new_n11626_));
  NAND2X1  g11433(.A(\a[60] ), .B(\a[44] ), .Y(new_n11627_));
  OAI22X1  g11434(.A0(new_n11627_), .A1(new_n11624_), .B0(new_n11626_), .B1(new_n11622_), .Y(new_n11628_));
  AND2X1   g11435(.A(new_n6119_), .B(new_n3893_), .Y(new_n11629_));
  NOR4X1   g11436(.A(new_n5379_), .B(new_n6022_), .C(new_n3926_), .D(new_n3460_), .Y(new_n11630_));
  OAI22X1  g11437(.A0(new_n11630_), .A1(new_n11629_), .B0(new_n11496_), .B1(new_n8297_), .Y(new_n11631_));
  NAND3X1  g11438(.A(new_n11631_), .B(\a[58] ), .C(\a[46] ), .Y(new_n11632_));
  OAI21X1  g11439(.A0(new_n11496_), .A1(new_n8297_), .B0(new_n11631_), .Y(new_n11633_));
  AOI22X1  g11440(.A0(\a[57] ), .A1(\a[47] ), .B0(\a[56] ), .B1(\a[48] ), .Y(new_n11634_));
  OAI21X1  g11441(.A0(new_n11634_), .A1(new_n11633_), .B0(new_n11632_), .Y(new_n11635_));
  XOR2X1   g11442(.A(new_n11635_), .B(new_n11628_), .Y(new_n11636_));
  INVX1    g11443(.A(new_n8136_), .Y(new_n11637_));
  AOI22X1  g11444(.A0(new_n8136_), .A1(new_n4904_), .B0(new_n5240_), .B1(new_n4321_), .Y(new_n11638_));
  AOI21X1  g11445(.A0(new_n5238_), .A1(new_n4484_), .B0(new_n11638_), .Y(new_n11639_));
  AOI21X1  g11446(.A0(new_n5238_), .A1(new_n4484_), .B0(new_n11639_), .Y(new_n11640_));
  INVX1    g11447(.A(new_n11640_), .Y(new_n11641_));
  AOI22X1  g11448(.A0(\a[54] ), .A1(\a[50] ), .B0(\a[53] ), .B1(\a[51] ), .Y(new_n11642_));
  OAI22X1  g11449(.A0(new_n11642_), .A1(new_n11641_), .B0(new_n11639_), .B1(new_n11637_), .Y(new_n11643_));
  INVX1    g11450(.A(new_n11643_), .Y(new_n11644_));
  XOR2X1   g11451(.A(new_n11644_), .B(new_n11636_), .Y(new_n11645_));
  XOR2X1   g11452(.A(new_n11645_), .B(new_n11621_), .Y(new_n11646_));
  XOR2X1   g11453(.A(new_n11646_), .B(new_n11614_), .Y(new_n11647_));
  AND2X1   g11454(.A(new_n11580_), .B(new_n11570_), .Y(new_n11648_));
  AOI21X1  g11455(.A0(new_n11581_), .A1(new_n11566_), .B0(new_n11648_), .Y(new_n11649_));
  NOR2X1   g11456(.A(new_n11588_), .B(new_n11586_), .Y(new_n11650_));
  AOI21X1  g11457(.A0(new_n11592_), .A1(new_n11589_), .B0(new_n11650_), .Y(new_n11651_));
  XOR2X1   g11458(.A(new_n11651_), .B(new_n11649_), .Y(new_n11652_));
  AND2X1   g11459(.A(new_n5048_), .B(new_n4321_), .Y(new_n11653_));
  OAI21X1  g11460(.A0(new_n11505_), .A1(new_n11653_), .B0(new_n11568_), .Y(new_n11654_));
  OAI21X1  g11461(.A0(new_n11569_), .A1(new_n11502_), .B0(new_n11654_), .Y(new_n11655_));
  INVX1    g11462(.A(new_n11563_), .Y(new_n11656_));
  AOI22X1  g11463(.A0(\a[63] ), .A1(\a[41] ), .B0(\a[62] ), .B1(\a[42] ), .Y(new_n11657_));
  AOI21X1  g11464(.A0(new_n6789_), .A1(new_n3607_), .B0(new_n11657_), .Y(new_n11658_));
  XOR2X1   g11465(.A(new_n11658_), .B(new_n11656_), .Y(new_n11659_));
  XOR2X1   g11466(.A(new_n11659_), .B(new_n11655_), .Y(new_n11660_));
  NAND2X1  g11467(.A(new_n11579_), .B(new_n11571_), .Y(new_n11661_));
  OAI21X1  g11468(.A0(new_n11493_), .A1(new_n11481_), .B0(new_n11661_), .Y(new_n11662_));
  XOR2X1   g11469(.A(new_n11662_), .B(new_n11660_), .Y(new_n11663_));
  XOR2X1   g11470(.A(new_n11663_), .B(new_n11652_), .Y(new_n11664_));
  XOR2X1   g11471(.A(new_n11664_), .B(new_n11647_), .Y(new_n11665_));
  XOR2X1   g11472(.A(new_n11665_), .B(new_n11612_), .Y(new_n11666_));
  XOR2X1   g11473(.A(new_n11666_), .B(new_n11608_), .Y(\asquared[105] ));
  XOR2X1   g11474(.A(new_n11641_), .B(new_n11633_), .Y(new_n11668_));
  XOR2X1   g11475(.A(new_n11668_), .B(new_n11625_), .Y(new_n11669_));
  AND2X1   g11476(.A(new_n11635_), .B(new_n11628_), .Y(new_n11670_));
  AOI21X1  g11477(.A0(new_n11643_), .A1(new_n11636_), .B0(new_n11670_), .Y(new_n11671_));
  XOR2X1   g11478(.A(new_n11671_), .B(new_n11669_), .Y(new_n11672_));
  AND2X1   g11479(.A(new_n11659_), .B(new_n11655_), .Y(new_n11673_));
  AOI21X1  g11480(.A0(new_n11662_), .A1(new_n11660_), .B0(new_n11673_), .Y(new_n11674_));
  XOR2X1   g11481(.A(new_n11674_), .B(new_n11672_), .Y(new_n11675_));
  NOR2X1   g11482(.A(new_n11651_), .B(new_n11649_), .Y(new_n11676_));
  AOI21X1  g11483(.A0(new_n11663_), .A1(new_n11652_), .B0(new_n11676_), .Y(new_n11677_));
  XOR2X1   g11484(.A(new_n11677_), .B(new_n11675_), .Y(new_n11678_));
  NAND2X1  g11485(.A(new_n11620_), .B(new_n11616_), .Y(new_n11679_));
  OAI21X1  g11486(.A0(new_n11645_), .A1(new_n11621_), .B0(new_n11679_), .Y(new_n11680_));
  AND2X1   g11487(.A(\a[53] ), .B(\a[43] ), .Y(new_n11681_));
  AOI21X1  g11488(.A0(new_n11681_), .A1(\a[62] ), .B0(new_n7336_), .Y(new_n11682_));
  AOI21X1  g11489(.A0(new_n11681_), .A1(\a[62] ), .B0(new_n5048_), .Y(new_n11683_));
  INVX1    g11490(.A(new_n11683_), .Y(new_n11684_));
  AOI21X1  g11491(.A0(\a[62] ), .A1(\a[43] ), .B0(\a[53] ), .Y(new_n11685_));
  OAI22X1  g11492(.A0(new_n11685_), .A1(new_n11684_), .B0(new_n11682_), .B1(new_n7336_), .Y(new_n11686_));
  INVX1    g11493(.A(new_n11686_), .Y(new_n11687_));
  NAND4X1  g11494(.A(\a[56] ), .B(\a[54] ), .C(\a[51] ), .D(\a[49] ), .Y(new_n11688_));
  NAND4X1  g11495(.A(\a[56] ), .B(\a[55] ), .C(\a[50] ), .D(\a[49] ), .Y(new_n11689_));
  AOI22X1  g11496(.A0(new_n11689_), .A1(new_n11688_), .B0(new_n5240_), .B1(new_n4484_), .Y(new_n11690_));
  NAND2X1  g11497(.A(\a[56] ), .B(\a[49] ), .Y(new_n11691_));
  AOI22X1  g11498(.A0(\a[55] ), .A1(\a[50] ), .B0(\a[54] ), .B1(\a[51] ), .Y(new_n11692_));
  AOI21X1  g11499(.A0(new_n5240_), .A1(new_n4484_), .B0(new_n11690_), .Y(new_n11693_));
  INVX1    g11500(.A(new_n11693_), .Y(new_n11694_));
  OAI22X1  g11501(.A0(new_n11694_), .A1(new_n11692_), .B0(new_n11691_), .B1(new_n11690_), .Y(new_n11695_));
  XOR2X1   g11502(.A(new_n11695_), .B(new_n11687_), .Y(new_n11696_));
  NOR2X1   g11503(.A(new_n11558_), .B(new_n11552_), .Y(new_n11697_));
  AOI21X1  g11504(.A0(new_n11615_), .A1(new_n11578_), .B0(new_n11697_), .Y(new_n11698_));
  XOR2X1   g11505(.A(new_n11698_), .B(new_n11696_), .Y(new_n11699_));
  NAND4X1  g11506(.A(\a[63] ), .B(\a[60] ), .C(\a[45] ), .D(\a[42] ), .Y(new_n11700_));
  NAND4X1  g11507(.A(\a[63] ), .B(\a[61] ), .C(\a[44] ), .D(\a[42] ), .Y(new_n11701_));
  AOI22X1  g11508(.A0(new_n11701_), .A1(new_n11700_), .B0(new_n6428_), .B1(new_n3918_), .Y(new_n11702_));
  AND2X1   g11509(.A(\a[63] ), .B(\a[42] ), .Y(new_n11703_));
  INVX1    g11510(.A(new_n11703_), .Y(new_n11704_));
  AOI21X1  g11511(.A0(new_n6428_), .A1(new_n3918_), .B0(new_n11702_), .Y(new_n11705_));
  INVX1    g11512(.A(new_n11705_), .Y(new_n11706_));
  AOI22X1  g11513(.A0(\a[61] ), .A1(\a[44] ), .B0(\a[60] ), .B1(\a[45] ), .Y(new_n11707_));
  OAI22X1  g11514(.A0(new_n11707_), .A1(new_n11706_), .B0(new_n11704_), .B1(new_n11702_), .Y(new_n11708_));
  AOI22X1  g11515(.A0(new_n11658_), .A1(new_n11656_), .B0(new_n6789_), .B1(new_n3607_), .Y(new_n11709_));
  XOR2X1   g11516(.A(new_n11709_), .B(new_n11708_), .Y(new_n11710_));
  OAI22X1  g11517(.A0(new_n6793_), .A1(new_n8296_), .B0(new_n8155_), .B1(new_n8299_), .Y(new_n11711_));
  OAI21X1  g11518(.A0(new_n8154_), .A1(new_n8297_), .B0(new_n11711_), .Y(new_n11712_));
  AND2X1   g11519(.A(\a[59] ), .B(\a[46] ), .Y(new_n11713_));
  AOI21X1  g11520(.A0(new_n6119_), .A1(new_n4272_), .B0(new_n11711_), .Y(new_n11714_));
  OAI22X1  g11521(.A0(new_n5379_), .A1(new_n4041_), .B0(new_n5441_), .B1(new_n3926_), .Y(new_n11715_));
  AOI22X1  g11522(.A0(new_n11715_), .A1(new_n11714_), .B0(new_n11713_), .B1(new_n11712_), .Y(new_n11716_));
  XOR2X1   g11523(.A(new_n11716_), .B(new_n11710_), .Y(new_n11717_));
  XOR2X1   g11524(.A(new_n11717_), .B(new_n11699_), .Y(new_n11718_));
  XOR2X1   g11525(.A(new_n11718_), .B(new_n11680_), .Y(new_n11719_));
  XOR2X1   g11526(.A(new_n11719_), .B(new_n11678_), .Y(new_n11720_));
  AND2X1   g11527(.A(new_n11598_), .B(new_n11593_), .Y(new_n11721_));
  OAI21X1  g11528(.A0(new_n11721_), .A1(new_n11613_), .B0(new_n11646_), .Y(new_n11722_));
  INVX1    g11529(.A(new_n11664_), .Y(new_n11723_));
  OAI21X1  g11530(.A0(new_n11723_), .A1(new_n11647_), .B0(new_n11722_), .Y(new_n11724_));
  NOR2X1   g11531(.A(new_n11724_), .B(new_n11720_), .Y(new_n11725_));
  AND2X1   g11532(.A(new_n11724_), .B(new_n11720_), .Y(new_n11726_));
  OR2X1    g11533(.A(new_n11726_), .B(new_n11725_), .Y(new_n11727_));
  NOR2X1   g11534(.A(new_n11665_), .B(new_n11612_), .Y(new_n11728_));
  AND2X1   g11535(.A(new_n11665_), .B(new_n11612_), .Y(new_n11729_));
  INVX1    g11536(.A(new_n11729_), .Y(new_n11730_));
  AOI21X1  g11537(.A0(new_n11730_), .A1(new_n11608_), .B0(new_n11728_), .Y(new_n11731_));
  XOR2X1   g11538(.A(new_n11731_), .B(new_n11727_), .Y(\asquared[106] ));
  NAND2X1  g11539(.A(new_n11719_), .B(new_n11678_), .Y(new_n11733_));
  OAI21X1  g11540(.A0(new_n11677_), .A1(new_n11675_), .B0(new_n11733_), .Y(new_n11734_));
  AND2X1   g11541(.A(new_n11671_), .B(new_n11669_), .Y(new_n11735_));
  OR2X1    g11542(.A(new_n11671_), .B(new_n11669_), .Y(new_n11736_));
  OAI21X1  g11543(.A0(new_n11674_), .A1(new_n11735_), .B0(new_n11736_), .Y(new_n11737_));
  NAND4X1  g11544(.A(\a[59] ), .B(\a[57] ), .C(\a[49] ), .D(\a[47] ), .Y(new_n11738_));
  NAND4X1  g11545(.A(\a[59] ), .B(\a[58] ), .C(\a[48] ), .D(\a[47] ), .Y(new_n11739_));
  AOI22X1  g11546(.A0(new_n11739_), .A1(new_n11738_), .B0(new_n6119_), .B1(new_n4274_), .Y(new_n11740_));
  AOI21X1  g11547(.A0(new_n6119_), .A1(new_n4274_), .B0(new_n11740_), .Y(new_n11741_));
  INVX1    g11548(.A(new_n11741_), .Y(new_n11742_));
  AOI22X1  g11549(.A0(\a[58] ), .A1(\a[48] ), .B0(\a[57] ), .B1(\a[49] ), .Y(new_n11743_));
  NAND2X1  g11550(.A(\a[59] ), .B(\a[47] ), .Y(new_n11744_));
  OAI22X1  g11551(.A0(new_n11744_), .A1(new_n11740_), .B0(new_n11743_), .B1(new_n11742_), .Y(new_n11745_));
  NAND4X1  g11552(.A(\a[56] ), .B(\a[54] ), .C(\a[52] ), .D(\a[50] ), .Y(new_n11746_));
  NAND4X1  g11553(.A(\a[56] ), .B(\a[55] ), .C(\a[51] ), .D(\a[50] ), .Y(new_n11747_));
  AOI22X1  g11554(.A0(new_n11747_), .A1(new_n11746_), .B0(new_n5240_), .B1(new_n7164_), .Y(new_n11748_));
  NAND2X1  g11555(.A(\a[56] ), .B(\a[50] ), .Y(new_n11749_));
  AOI21X1  g11556(.A0(new_n5240_), .A1(new_n7164_), .B0(new_n11748_), .Y(new_n11750_));
  INVX1    g11557(.A(new_n11750_), .Y(new_n11751_));
  AOI22X1  g11558(.A0(\a[55] ), .A1(\a[51] ), .B0(\a[54] ), .B1(\a[52] ), .Y(new_n11752_));
  OAI22X1  g11559(.A0(new_n11752_), .A1(new_n11751_), .B0(new_n11749_), .B1(new_n11748_), .Y(new_n11753_));
  XOR2X1   g11560(.A(new_n11753_), .B(new_n11745_), .Y(new_n11754_));
  AND2X1   g11561(.A(new_n11641_), .B(new_n11633_), .Y(new_n11755_));
  AOI21X1  g11562(.A0(new_n11668_), .A1(new_n11626_), .B0(new_n11755_), .Y(new_n11756_));
  XOR2X1   g11563(.A(new_n11756_), .B(new_n11754_), .Y(new_n11757_));
  XOR2X1   g11564(.A(new_n11714_), .B(new_n11705_), .Y(new_n11758_));
  INVX1    g11565(.A(new_n11758_), .Y(new_n11759_));
  INVX1    g11566(.A(new_n10045_), .Y(new_n11760_));
  NAND4X1  g11567(.A(\a[62] ), .B(\a[61] ), .C(\a[45] ), .D(\a[44] ), .Y(new_n11761_));
  NAND4X1  g11568(.A(\a[62] ), .B(\a[60] ), .C(\a[46] ), .D(\a[44] ), .Y(new_n11762_));
  AOI22X1  g11569(.A0(new_n11762_), .A1(new_n11761_), .B0(new_n6428_), .B1(new_n3809_), .Y(new_n11763_));
  NAND4X1  g11570(.A(\a[61] ), .B(\a[60] ), .C(\a[46] ), .D(\a[45] ), .Y(new_n11764_));
  NAND3X1  g11571(.A(new_n11762_), .B(new_n11761_), .C(new_n11764_), .Y(new_n11765_));
  AOI22X1  g11572(.A0(\a[61] ), .A1(\a[45] ), .B0(\a[60] ), .B1(\a[46] ), .Y(new_n11766_));
  OAI22X1  g11573(.A0(new_n11766_), .A1(new_n11765_), .B0(new_n11763_), .B1(new_n11760_), .Y(new_n11767_));
  XOR2X1   g11574(.A(new_n11767_), .B(new_n11759_), .Y(new_n11768_));
  NAND2X1  g11575(.A(new_n11768_), .B(new_n11757_), .Y(new_n11769_));
  OR2X1    g11576(.A(new_n11768_), .B(new_n11757_), .Y(new_n11770_));
  NAND3X1  g11577(.A(new_n11769_), .B(new_n11770_), .C(new_n11737_), .Y(new_n11771_));
  AND2X1   g11578(.A(new_n11771_), .B(new_n11770_), .Y(new_n11772_));
  AOI22X1  g11579(.A0(new_n11772_), .A1(new_n11769_), .B0(new_n11771_), .B1(new_n11737_), .Y(new_n11773_));
  AND2X1   g11580(.A(\a[63] ), .B(\a[43] ), .Y(new_n11774_));
  XOR2X1   g11581(.A(new_n11774_), .B(new_n11684_), .Y(new_n11775_));
  XOR2X1   g11582(.A(new_n11775_), .B(new_n11694_), .Y(new_n11776_));
  INVX1    g11583(.A(new_n11708_), .Y(new_n11777_));
  OR2X1    g11584(.A(new_n11716_), .B(new_n11710_), .Y(new_n11778_));
  OAI21X1  g11585(.A0(new_n11709_), .A1(new_n11777_), .B0(new_n11778_), .Y(new_n11779_));
  XOR2X1   g11586(.A(new_n11779_), .B(new_n11776_), .Y(new_n11780_));
  NAND2X1  g11587(.A(new_n11695_), .B(new_n11686_), .Y(new_n11781_));
  OAI21X1  g11588(.A0(new_n11698_), .A1(new_n11696_), .B0(new_n11781_), .Y(new_n11782_));
  XOR2X1   g11589(.A(new_n11782_), .B(new_n11780_), .Y(new_n11783_));
  AND2X1   g11590(.A(new_n11717_), .B(new_n11699_), .Y(new_n11784_));
  AOI21X1  g11591(.A0(new_n11718_), .A1(new_n11680_), .B0(new_n11784_), .Y(new_n11785_));
  XOR2X1   g11592(.A(new_n11785_), .B(new_n11783_), .Y(new_n11786_));
  XOR2X1   g11593(.A(new_n11786_), .B(new_n11773_), .Y(new_n11787_));
  AND2X1   g11594(.A(new_n11787_), .B(new_n11734_), .Y(new_n11788_));
  INVX1    g11595(.A(new_n11788_), .Y(new_n11789_));
  INVX1    g11596(.A(new_n11726_), .Y(new_n11790_));
  OAI21X1  g11597(.A0(new_n11731_), .A1(new_n11725_), .B0(new_n11790_), .Y(new_n11791_));
  NOR2X1   g11598(.A(new_n11787_), .B(new_n11734_), .Y(new_n11792_));
  INVX1    g11599(.A(new_n11792_), .Y(new_n11793_));
  AOI21X1  g11600(.A0(new_n11793_), .A1(new_n11789_), .B0(new_n11791_), .Y(new_n11794_));
  AND2X1   g11601(.A(new_n11793_), .B(new_n11791_), .Y(new_n11795_));
  AOI21X1  g11602(.A0(new_n11795_), .A1(new_n11789_), .B0(new_n11794_), .Y(\asquared[107] ));
  AOI21X1  g11603(.A0(new_n11793_), .A1(new_n11791_), .B0(new_n11788_), .Y(new_n11797_));
  INVX1    g11604(.A(new_n11783_), .Y(new_n11798_));
  OR2X1    g11605(.A(new_n11785_), .B(new_n11798_), .Y(new_n11799_));
  OAI21X1  g11606(.A0(new_n11786_), .A1(new_n11773_), .B0(new_n11799_), .Y(new_n11800_));
  AND2X1   g11607(.A(new_n11779_), .B(new_n11776_), .Y(new_n11801_));
  AOI21X1  g11608(.A0(new_n11782_), .A1(new_n11780_), .B0(new_n11801_), .Y(new_n11802_));
  XOR2X1   g11609(.A(new_n11765_), .B(new_n11742_), .Y(new_n11803_));
  INVX1    g11610(.A(new_n11803_), .Y(new_n11804_));
  NOR4X1   g11611(.A(new_n6549_), .B(new_n5379_), .C(new_n3915_), .D(new_n5268_), .Y(new_n11805_));
  NAND4X1  g11612(.A(\a[59] ), .B(\a[58] ), .C(\a[49] ), .D(\a[48] ), .Y(new_n11806_));
  NAND4X1  g11613(.A(\a[63] ), .B(\a[59] ), .C(\a[48] ), .D(\a[44] ), .Y(new_n11807_));
  AOI21X1  g11614(.A0(new_n11807_), .A1(new_n11806_), .B0(new_n11805_), .Y(new_n11808_));
  NAND2X1  g11615(.A(\a[59] ), .B(\a[48] ), .Y(new_n11809_));
  AOI22X1  g11616(.A0(\a[63] ), .A1(\a[44] ), .B0(\a[58] ), .B1(\a[49] ), .Y(new_n11810_));
  NOR2X1   g11617(.A(new_n11808_), .B(new_n11805_), .Y(new_n11811_));
  INVX1    g11618(.A(new_n11811_), .Y(new_n11812_));
  OAI22X1  g11619(.A0(new_n11812_), .A1(new_n11810_), .B0(new_n11809_), .B1(new_n11808_), .Y(new_n11813_));
  XOR2X1   g11620(.A(new_n11813_), .B(new_n11804_), .Y(new_n11814_));
  NOR3X1   g11621(.A(new_n10302_), .B(new_n4835_), .C(new_n5245_), .Y(new_n11815_));
  OAI21X1  g11622(.A0(new_n10302_), .A1(\a[53] ), .B0(\a[54] ), .Y(new_n11816_));
  OAI21X1  g11623(.A0(new_n10302_), .A1(\a[54] ), .B0(new_n11816_), .Y(new_n11817_));
  OAI21X1  g11624(.A0(new_n11815_), .A1(new_n5239_), .B0(new_n11817_), .Y(new_n11818_));
  NAND4X1  g11625(.A(\a[57] ), .B(\a[55] ), .C(\a[52] ), .D(\a[50] ), .Y(new_n11819_));
  NAND4X1  g11626(.A(\a[57] ), .B(\a[56] ), .C(\a[51] ), .D(\a[50] ), .Y(new_n11820_));
  AOI22X1  g11627(.A0(new_n11820_), .A1(new_n11819_), .B0(new_n6237_), .B1(new_n7164_), .Y(new_n11821_));
  NAND2X1  g11628(.A(\a[57] ), .B(\a[50] ), .Y(new_n11822_));
  NAND4X1  g11629(.A(\a[56] ), .B(\a[55] ), .C(\a[52] ), .D(\a[51] ), .Y(new_n11823_));
  NAND3X1  g11630(.A(new_n11820_), .B(new_n11819_), .C(new_n11823_), .Y(new_n11824_));
  AOI22X1  g11631(.A0(\a[56] ), .A1(\a[51] ), .B0(\a[55] ), .B1(\a[52] ), .Y(new_n11825_));
  OAI22X1  g11632(.A0(new_n11825_), .A1(new_n11824_), .B0(new_n11822_), .B1(new_n11821_), .Y(new_n11826_));
  XOR2X1   g11633(.A(new_n11826_), .B(new_n11818_), .Y(new_n11827_));
  NAND2X1  g11634(.A(\a[60] ), .B(\a[47] ), .Y(new_n11828_));
  NAND2X1  g11635(.A(\a[61] ), .B(\a[46] ), .Y(new_n11829_));
  AOI22X1  g11636(.A0(new_n11829_), .A1(new_n11828_), .B0(new_n6428_), .B1(new_n3893_), .Y(new_n11830_));
  XOR2X1   g11637(.A(new_n11830_), .B(new_n11750_), .Y(new_n11831_));
  XOR2X1   g11638(.A(new_n11831_), .B(new_n11827_), .Y(new_n11832_));
  XOR2X1   g11639(.A(new_n11832_), .B(new_n11814_), .Y(new_n11833_));
  XOR2X1   g11640(.A(new_n11833_), .B(new_n11802_), .Y(new_n11834_));
  NOR2X1   g11641(.A(new_n11714_), .B(new_n11705_), .Y(new_n11835_));
  AOI21X1  g11642(.A0(new_n11767_), .A1(new_n11758_), .B0(new_n11835_), .Y(new_n11836_));
  NAND2X1  g11643(.A(new_n11774_), .B(new_n11684_), .Y(new_n11837_));
  NOR2X1   g11644(.A(new_n11774_), .B(new_n11684_), .Y(new_n11838_));
  OAI21X1  g11645(.A0(new_n11838_), .A1(new_n11693_), .B0(new_n11837_), .Y(new_n11839_));
  XOR2X1   g11646(.A(new_n11839_), .B(new_n11836_), .Y(new_n11840_));
  AND2X1   g11647(.A(new_n11753_), .B(new_n11745_), .Y(new_n11841_));
  INVX1    g11648(.A(new_n11756_), .Y(new_n11842_));
  AOI21X1  g11649(.A0(new_n11842_), .A1(new_n11754_), .B0(new_n11841_), .Y(new_n11843_));
  XOR2X1   g11650(.A(new_n11843_), .B(new_n11840_), .Y(new_n11844_));
  XOR2X1   g11651(.A(new_n11844_), .B(new_n11772_), .Y(new_n11845_));
  XOR2X1   g11652(.A(new_n11845_), .B(new_n11834_), .Y(new_n11846_));
  NOR2X1   g11653(.A(new_n11846_), .B(new_n11800_), .Y(new_n11847_));
  AND2X1   g11654(.A(new_n11846_), .B(new_n11800_), .Y(new_n11848_));
  OR2X1    g11655(.A(new_n11848_), .B(new_n11847_), .Y(new_n11849_));
  XOR2X1   g11656(.A(new_n11849_), .B(new_n11797_), .Y(\asquared[108] ));
  INVX1    g11657(.A(new_n11772_), .Y(new_n11851_));
  NAND2X1  g11658(.A(new_n11844_), .B(new_n11851_), .Y(new_n11852_));
  OAI21X1  g11659(.A0(new_n11845_), .A1(new_n11834_), .B0(new_n11852_), .Y(new_n11853_));
  AND2X1   g11660(.A(new_n11765_), .B(new_n11742_), .Y(new_n11854_));
  AOI21X1  g11661(.A0(new_n11813_), .A1(new_n11803_), .B0(new_n11854_), .Y(new_n11855_));
  NAND4X1  g11662(.A(\a[57] ), .B(\a[55] ), .C(\a[53] ), .D(\a[51] ), .Y(new_n11856_));
  OAI21X1  g11663(.A0(new_n11496_), .A1(new_n7793_), .B0(new_n11856_), .Y(new_n11857_));
  OAI21X1  g11664(.A0(new_n8560_), .A1(new_n7336_), .B0(new_n11857_), .Y(new_n11858_));
  AOI21X1  g11665(.A0(new_n6237_), .A1(new_n5048_), .B0(new_n11857_), .Y(new_n11859_));
  OAI22X1  g11666(.A0(new_n6022_), .A1(new_n4354_), .B0(new_n4906_), .B1(new_n5245_), .Y(new_n11860_));
  AOI22X1  g11667(.A0(new_n11860_), .A1(new_n11859_), .B0(new_n11858_), .B1(new_n9550_), .Y(new_n11861_));
  XOR2X1   g11668(.A(new_n11861_), .B(new_n11855_), .Y(new_n11862_));
  NAND2X1  g11669(.A(new_n11826_), .B(new_n11818_), .Y(new_n11863_));
  INVX1    g11670(.A(new_n11827_), .Y(new_n11864_));
  OAI21X1  g11671(.A0(new_n11831_), .A1(new_n11864_), .B0(new_n11863_), .Y(new_n11865_));
  XOR2X1   g11672(.A(new_n11865_), .B(new_n11862_), .Y(new_n11866_));
  OR2X1    g11673(.A(new_n11832_), .B(new_n11814_), .Y(new_n11867_));
  AND2X1   g11674(.A(new_n11832_), .B(new_n11814_), .Y(new_n11868_));
  OAI21X1  g11675(.A0(new_n11868_), .A1(new_n11802_), .B0(new_n11867_), .Y(new_n11869_));
  XOR2X1   g11676(.A(new_n11869_), .B(new_n11866_), .Y(new_n11870_));
  XOR2X1   g11677(.A(new_n11824_), .B(new_n11816_), .Y(new_n11871_));
  XOR2X1   g11678(.A(new_n11871_), .B(new_n11811_), .Y(new_n11872_));
  AND2X1   g11679(.A(new_n11767_), .B(new_n11758_), .Y(new_n11873_));
  OAI21X1  g11680(.A0(new_n11873_), .A1(new_n11835_), .B0(new_n11839_), .Y(new_n11874_));
  OAI21X1  g11681(.A0(new_n11843_), .A1(new_n11840_), .B0(new_n11874_), .Y(new_n11875_));
  XOR2X1   g11682(.A(new_n11875_), .B(new_n11872_), .Y(new_n11876_));
  NAND4X1  g11683(.A(\a[63] ), .B(\a[61] ), .C(\a[47] ), .D(\a[45] ), .Y(new_n11877_));
  NAND4X1  g11684(.A(\a[63] ), .B(\a[62] ), .C(\a[46] ), .D(\a[45] ), .Y(new_n11878_));
  AOI22X1  g11685(.A0(new_n11878_), .A1(new_n11877_), .B0(new_n6556_), .B1(new_n3893_), .Y(new_n11879_));
  NOR3X1   g11686(.A(new_n11879_), .B(new_n6549_), .C(new_n3811_), .Y(new_n11880_));
  AOI21X1  g11687(.A0(new_n6556_), .A1(new_n3893_), .B0(new_n11879_), .Y(new_n11881_));
  AOI22X1  g11688(.A0(\a[62] ), .A1(\a[46] ), .B0(\a[61] ), .B1(\a[47] ), .Y(new_n11882_));
  INVX1    g11689(.A(new_n11882_), .Y(new_n11883_));
  AOI21X1  g11690(.A0(new_n11883_), .A1(new_n11881_), .B0(new_n11880_), .Y(new_n11884_));
  INVX1    g11691(.A(new_n11884_), .Y(new_n11885_));
  AOI22X1  g11692(.A0(new_n11830_), .A1(new_n11751_), .B0(new_n6428_), .B1(new_n3893_), .Y(new_n11886_));
  XOR2X1   g11693(.A(new_n11886_), .B(new_n11885_), .Y(new_n11887_));
  OAI22X1  g11694(.A0(new_n6796_), .A1(new_n8802_), .B0(new_n6794_), .B1(new_n4280_), .Y(new_n11888_));
  OAI21X1  g11695(.A0(new_n6793_), .A1(new_n7652_), .B0(new_n11888_), .Y(new_n11889_));
  AND2X1   g11696(.A(\a[60] ), .B(\a[48] ), .Y(new_n11890_));
  OAI22X1  g11697(.A0(new_n5617_), .A1(new_n3915_), .B0(new_n5379_), .B1(new_n4983_), .Y(new_n11891_));
  AOI21X1  g11698(.A0(new_n6121_), .A1(new_n4321_), .B0(new_n11888_), .Y(new_n11892_));
  AOI22X1  g11699(.A0(new_n11892_), .A1(new_n11891_), .B0(new_n11890_), .B1(new_n11889_), .Y(new_n11893_));
  XOR2X1   g11700(.A(new_n11893_), .B(new_n11887_), .Y(new_n11894_));
  XOR2X1   g11701(.A(new_n11894_), .B(new_n11876_), .Y(new_n11895_));
  XOR2X1   g11702(.A(new_n11895_), .B(new_n11870_), .Y(new_n11896_));
  AND2X1   g11703(.A(new_n11896_), .B(new_n11853_), .Y(new_n11897_));
  INVX1    g11704(.A(new_n11897_), .Y(new_n11898_));
  INVX1    g11705(.A(new_n11848_), .Y(new_n11899_));
  OAI21X1  g11706(.A0(new_n11847_), .A1(new_n11797_), .B0(new_n11899_), .Y(new_n11900_));
  NOR2X1   g11707(.A(new_n11896_), .B(new_n11853_), .Y(new_n11901_));
  INVX1    g11708(.A(new_n11901_), .Y(new_n11902_));
  AOI21X1  g11709(.A0(new_n11898_), .A1(new_n11902_), .B0(new_n11900_), .Y(new_n11903_));
  AND2X1   g11710(.A(new_n11902_), .B(new_n11900_), .Y(new_n11904_));
  AOI21X1  g11711(.A0(new_n11904_), .A1(new_n11898_), .B0(new_n11903_), .Y(\asquared[109] ));
  AOI21X1  g11712(.A0(new_n11902_), .A1(new_n11900_), .B0(new_n11897_), .Y(new_n11906_));
  AND2X1   g11713(.A(new_n10302_), .B(\a[54] ), .Y(new_n11907_));
  OAI21X1  g11714(.A0(new_n11815_), .A1(new_n11907_), .B0(new_n11824_), .Y(new_n11908_));
  OAI21X1  g11715(.A0(new_n11871_), .A1(new_n11811_), .B0(new_n11908_), .Y(new_n11909_));
  NOR3X1   g11716(.A(new_n10759_), .B(new_n4906_), .C(new_n4835_), .Y(new_n11910_));
  OAI21X1  g11717(.A0(new_n10759_), .A1(\a[54] ), .B0(\a[55] ), .Y(new_n11911_));
  OAI21X1  g11718(.A0(new_n10759_), .A1(\a[55] ), .B0(new_n11911_), .Y(new_n11912_));
  OAI21X1  g11719(.A0(new_n11910_), .A1(new_n5241_), .B0(new_n11912_), .Y(new_n11913_));
  XOR2X1   g11720(.A(new_n11913_), .B(new_n11909_), .Y(new_n11914_));
  OR2X1    g11721(.A(new_n11886_), .B(new_n11884_), .Y(new_n11915_));
  OAI21X1  g11722(.A0(new_n11893_), .A1(new_n11887_), .B0(new_n11915_), .Y(new_n11916_));
  XOR2X1   g11723(.A(new_n11916_), .B(new_n11914_), .Y(new_n11917_));
  INVX1    g11724(.A(new_n11917_), .Y(new_n11918_));
  AND2X1   g11725(.A(new_n11875_), .B(new_n11872_), .Y(new_n11919_));
  AOI21X1  g11726(.A0(new_n11894_), .A1(new_n11876_), .B0(new_n11919_), .Y(new_n11920_));
  XOR2X1   g11727(.A(new_n11920_), .B(new_n11918_), .Y(new_n11921_));
  INVX1    g11728(.A(new_n11921_), .Y(new_n11922_));
  AND2X1   g11729(.A(\a[63] ), .B(\a[46] ), .Y(new_n11923_));
  INVX1    g11730(.A(new_n11923_), .Y(new_n11924_));
  XOR2X1   g11731(.A(new_n11924_), .B(new_n11859_), .Y(new_n11925_));
  XOR2X1   g11732(.A(new_n11925_), .B(new_n11892_), .Y(new_n11926_));
  NOR2X1   g11733(.A(new_n11861_), .B(new_n11855_), .Y(new_n11927_));
  AOI21X1  g11734(.A0(new_n11865_), .A1(new_n11862_), .B0(new_n11927_), .Y(new_n11928_));
  XOR2X1   g11735(.A(new_n11928_), .B(new_n11926_), .Y(new_n11929_));
  NAND4X1  g11736(.A(\a[61] ), .B(\a[59] ), .C(\a[50] ), .D(\a[48] ), .Y(new_n11930_));
  NAND4X1  g11737(.A(\a[61] ), .B(\a[60] ), .C(\a[49] ), .D(\a[48] ), .Y(new_n11931_));
  AOI22X1  g11738(.A0(new_n11931_), .A1(new_n11930_), .B0(new_n6427_), .B1(new_n4321_), .Y(new_n11932_));
  AND2X1   g11739(.A(\a[61] ), .B(\a[48] ), .Y(new_n11933_));
  INVX1    g11740(.A(new_n11933_), .Y(new_n11934_));
  AOI21X1  g11741(.A0(new_n6427_), .A1(new_n4321_), .B0(new_n11932_), .Y(new_n11935_));
  INVX1    g11742(.A(new_n11935_), .Y(new_n11936_));
  AOI22X1  g11743(.A0(\a[60] ), .A1(\a[49] ), .B0(\a[59] ), .B1(\a[50] ), .Y(new_n11937_));
  OAI22X1  g11744(.A0(new_n11937_), .A1(new_n11936_), .B0(new_n11934_), .B1(new_n11932_), .Y(new_n11938_));
  XOR2X1   g11745(.A(new_n11938_), .B(new_n11881_), .Y(new_n11939_));
  NAND4X1  g11746(.A(\a[58] ), .B(\a[56] ), .C(\a[53] ), .D(\a[51] ), .Y(new_n11940_));
  OAI21X1  g11747(.A0(new_n8154_), .A1(new_n7793_), .B0(new_n11940_), .Y(new_n11941_));
  OAI21X1  g11748(.A0(new_n11496_), .A1(new_n7336_), .B0(new_n11941_), .Y(new_n11942_));
  AND2X1   g11749(.A(\a[58] ), .B(\a[51] ), .Y(new_n11943_));
  AOI21X1  g11750(.A0(new_n5554_), .A1(new_n5048_), .B0(new_n11941_), .Y(new_n11944_));
  OAI22X1  g11751(.A0(new_n5441_), .A1(new_n4354_), .B0(new_n6022_), .B1(new_n5245_), .Y(new_n11945_));
  AOI22X1  g11752(.A0(new_n11945_), .A1(new_n11944_), .B0(new_n11943_), .B1(new_n11942_), .Y(new_n11946_));
  XOR2X1   g11753(.A(new_n11946_), .B(new_n11939_), .Y(new_n11947_));
  XOR2X1   g11754(.A(new_n11947_), .B(new_n11929_), .Y(new_n11948_));
  XOR2X1   g11755(.A(new_n11948_), .B(new_n11922_), .Y(new_n11949_));
  AND2X1   g11756(.A(new_n11869_), .B(new_n11866_), .Y(new_n11950_));
  AOI21X1  g11757(.A0(new_n11895_), .A1(new_n11870_), .B0(new_n11950_), .Y(new_n11951_));
  NOR2X1   g11758(.A(new_n11951_), .B(new_n11949_), .Y(new_n11952_));
  AND2X1   g11759(.A(new_n11951_), .B(new_n11949_), .Y(new_n11953_));
  OR2X1    g11760(.A(new_n11953_), .B(new_n11952_), .Y(new_n11954_));
  XOR2X1   g11761(.A(new_n11954_), .B(new_n11906_), .Y(\asquared[110] ));
  NAND2X1  g11762(.A(new_n11948_), .B(new_n11921_), .Y(new_n11956_));
  OAI21X1  g11763(.A0(new_n11920_), .A1(new_n11918_), .B0(new_n11956_), .Y(new_n11957_));
  XOR2X1   g11764(.A(new_n11944_), .B(new_n11935_), .Y(new_n11958_));
  NAND4X1  g11765(.A(\a[61] ), .B(\a[59] ), .C(\a[51] ), .D(\a[49] ), .Y(new_n11959_));
  NAND4X1  g11766(.A(\a[61] ), .B(\a[60] ), .C(\a[50] ), .D(\a[49] ), .Y(new_n11960_));
  AOI22X1  g11767(.A0(new_n11960_), .A1(new_n11959_), .B0(new_n6427_), .B1(new_n4484_), .Y(new_n11961_));
  AND2X1   g11768(.A(\a[61] ), .B(\a[49] ), .Y(new_n11962_));
  INVX1    g11769(.A(new_n11962_), .Y(new_n11963_));
  AOI21X1  g11770(.A0(new_n6427_), .A1(new_n4484_), .B0(new_n11961_), .Y(new_n11964_));
  INVX1    g11771(.A(new_n11964_), .Y(new_n11965_));
  AOI22X1  g11772(.A0(\a[60] ), .A1(\a[50] ), .B0(\a[59] ), .B1(\a[51] ), .Y(new_n11966_));
  OAI22X1  g11773(.A0(new_n11966_), .A1(new_n11965_), .B0(new_n11963_), .B1(new_n11961_), .Y(new_n11967_));
  XOR2X1   g11774(.A(new_n11967_), .B(new_n11958_), .Y(new_n11968_));
  INVX1    g11775(.A(new_n11968_), .Y(new_n11969_));
  INVX1    g11776(.A(new_n11938_), .Y(new_n11970_));
  OR2X1    g11777(.A(new_n11946_), .B(new_n11939_), .Y(new_n11971_));
  OAI21X1  g11778(.A0(new_n11970_), .A1(new_n11881_), .B0(new_n11971_), .Y(new_n11972_));
  XOR2X1   g11779(.A(new_n11972_), .B(new_n11969_), .Y(new_n11973_));
  AND2X1   g11780(.A(new_n11913_), .B(new_n11909_), .Y(new_n11974_));
  AOI21X1  g11781(.A0(new_n11916_), .A1(new_n11914_), .B0(new_n11974_), .Y(new_n11975_));
  XOR2X1   g11782(.A(new_n11975_), .B(new_n11973_), .Y(new_n11976_));
  INVX1    g11783(.A(new_n11911_), .Y(new_n11977_));
  AOI22X1  g11784(.A0(\a[63] ), .A1(\a[47] ), .B0(\a[62] ), .B1(\a[48] ), .Y(new_n11978_));
  AOI21X1  g11785(.A0(new_n6789_), .A1(new_n4272_), .B0(new_n11978_), .Y(new_n11979_));
  XOR2X1   g11786(.A(new_n11979_), .B(new_n11977_), .Y(new_n11980_));
  AND2X1   g11787(.A(new_n6119_), .B(new_n5048_), .Y(new_n11981_));
  NOR4X1   g11788(.A(new_n5379_), .B(new_n6022_), .C(new_n4835_), .D(new_n4354_), .Y(new_n11982_));
  OAI22X1  g11789(.A0(new_n11982_), .A1(new_n11981_), .B0(new_n11496_), .B1(new_n5239_), .Y(new_n11983_));
  NAND3X1  g11790(.A(new_n11983_), .B(\a[58] ), .C(\a[52] ), .Y(new_n11984_));
  OAI21X1  g11791(.A0(new_n11496_), .A1(new_n5239_), .B0(new_n11983_), .Y(new_n11985_));
  AOI22X1  g11792(.A0(\a[57] ), .A1(\a[53] ), .B0(\a[56] ), .B1(\a[54] ), .Y(new_n11986_));
  OAI21X1  g11793(.A0(new_n11986_), .A1(new_n11985_), .B0(new_n11984_), .Y(new_n11987_));
  XOR2X1   g11794(.A(new_n11987_), .B(new_n11980_), .Y(new_n11988_));
  OR2X1    g11795(.A(new_n11924_), .B(new_n11859_), .Y(new_n11989_));
  AND2X1   g11796(.A(new_n11924_), .B(new_n11859_), .Y(new_n11990_));
  OAI21X1  g11797(.A0(new_n11990_), .A1(new_n11892_), .B0(new_n11989_), .Y(new_n11991_));
  XOR2X1   g11798(.A(new_n11991_), .B(new_n11988_), .Y(new_n11992_));
  NOR2X1   g11799(.A(new_n11928_), .B(new_n11926_), .Y(new_n11993_));
  AOI21X1  g11800(.A0(new_n11947_), .A1(new_n11929_), .B0(new_n11993_), .Y(new_n11994_));
  OR2X1    g11801(.A(new_n11994_), .B(new_n11992_), .Y(new_n11995_));
  INVX1    g11802(.A(new_n11992_), .Y(new_n11996_));
  XOR2X1   g11803(.A(new_n11994_), .B(new_n11996_), .Y(new_n11997_));
  AOI21X1  g11804(.A0(new_n11994_), .A1(new_n11992_), .B0(new_n11976_), .Y(new_n11998_));
  AOI22X1  g11805(.A0(new_n11998_), .A1(new_n11995_), .B0(new_n11997_), .B1(new_n11976_), .Y(new_n11999_));
  AND2X1   g11806(.A(new_n11999_), .B(new_n11957_), .Y(new_n12000_));
  INVX1    g11807(.A(new_n12000_), .Y(new_n12001_));
  INVX1    g11808(.A(new_n11952_), .Y(new_n12002_));
  OAI21X1  g11809(.A0(new_n11953_), .A1(new_n11906_), .B0(new_n12002_), .Y(new_n12003_));
  NOR2X1   g11810(.A(new_n11999_), .B(new_n11957_), .Y(new_n12004_));
  INVX1    g11811(.A(new_n12004_), .Y(new_n12005_));
  AOI21X1  g11812(.A0(new_n12001_), .A1(new_n12005_), .B0(new_n12003_), .Y(new_n12006_));
  AND2X1   g11813(.A(new_n12005_), .B(new_n12003_), .Y(new_n12007_));
  AOI21X1  g11814(.A0(new_n12007_), .A1(new_n12001_), .B0(new_n12006_), .Y(\asquared[111] ));
  AOI21X1  g11815(.A0(new_n12005_), .A1(new_n12003_), .B0(new_n12000_), .Y(new_n12009_));
  NOR2X1   g11816(.A(new_n11994_), .B(new_n11996_), .Y(new_n12010_));
  AOI21X1  g11817(.A0(new_n11997_), .A1(new_n11976_), .B0(new_n12010_), .Y(new_n12011_));
  XOR2X1   g11818(.A(new_n11985_), .B(new_n11965_), .Y(new_n12012_));
  AOI22X1  g11819(.A0(new_n11979_), .A1(new_n11977_), .B0(new_n6789_), .B1(new_n4272_), .Y(new_n12013_));
  INVX1    g11820(.A(new_n12013_), .Y(new_n12014_));
  XOR2X1   g11821(.A(new_n12014_), .B(new_n12012_), .Y(new_n12015_));
  INVX1    g11822(.A(new_n12015_), .Y(new_n12016_));
  NOR2X1   g11823(.A(new_n11944_), .B(new_n11935_), .Y(new_n12017_));
  AOI21X1  g11824(.A0(new_n11967_), .A1(new_n11958_), .B0(new_n12017_), .Y(new_n12018_));
  XOR2X1   g11825(.A(new_n12018_), .B(new_n12016_), .Y(new_n12019_));
  INVX1    g11826(.A(new_n12019_), .Y(new_n12020_));
  AND2X1   g11827(.A(new_n11987_), .B(new_n11980_), .Y(new_n12021_));
  AOI21X1  g11828(.A0(new_n11991_), .A1(new_n11988_), .B0(new_n12021_), .Y(new_n12022_));
  XOR2X1   g11829(.A(new_n12022_), .B(new_n12020_), .Y(new_n12023_));
  INVX1    g11830(.A(new_n12023_), .Y(new_n12024_));
  NAND4X1  g11831(.A(\a[63] ), .B(\a[60] ), .C(\a[51] ), .D(\a[48] ), .Y(new_n12025_));
  NAND4X1  g11832(.A(\a[63] ), .B(\a[61] ), .C(\a[50] ), .D(\a[48] ), .Y(new_n12026_));
  AOI22X1  g11833(.A0(new_n12026_), .A1(new_n12025_), .B0(new_n6428_), .B1(new_n4484_), .Y(new_n12027_));
  AOI21X1  g11834(.A0(new_n6428_), .A1(new_n4484_), .B0(new_n12027_), .Y(new_n12028_));
  INVX1    g11835(.A(new_n12028_), .Y(new_n12029_));
  AOI22X1  g11836(.A0(\a[61] ), .A1(\a[50] ), .B0(\a[60] ), .B1(\a[51] ), .Y(new_n12030_));
  NAND2X1  g11837(.A(\a[63] ), .B(\a[48] ), .Y(new_n12031_));
  OAI22X1  g11838(.A0(new_n12031_), .A1(new_n12027_), .B0(new_n12030_), .B1(new_n12029_), .Y(new_n12032_));
  AND2X1   g11839(.A(\a[62] ), .B(\a[56] ), .Y(new_n12033_));
  AOI21X1  g11840(.A0(new_n12033_), .A1(\a[49] ), .B0(new_n8560_), .Y(new_n12034_));
  AOI21X1  g11841(.A0(new_n12033_), .A1(\a[49] ), .B0(new_n6237_), .Y(new_n12035_));
  INVX1    g11842(.A(new_n12035_), .Y(new_n12036_));
  AOI21X1  g11843(.A0(\a[62] ), .A1(\a[49] ), .B0(\a[56] ), .Y(new_n12037_));
  OAI22X1  g11844(.A0(new_n12037_), .A1(new_n12036_), .B0(new_n12034_), .B1(new_n8560_), .Y(new_n12038_));
  INVX1    g11845(.A(new_n12038_), .Y(new_n12039_));
  XOR2X1   g11846(.A(new_n12039_), .B(new_n12032_), .Y(new_n12040_));
  OAI22X1  g11847(.A0(new_n7338_), .A1(new_n8155_), .B0(new_n6793_), .B1(new_n7336_), .Y(new_n12041_));
  OAI21X1  g11848(.A0(new_n8154_), .A1(new_n5239_), .B0(new_n12041_), .Y(new_n12042_));
  AND2X1   g11849(.A(\a[59] ), .B(\a[52] ), .Y(new_n12043_));
  OAI22X1  g11850(.A0(new_n5379_), .A1(new_n5245_), .B0(new_n5441_), .B1(new_n4835_), .Y(new_n12044_));
  AOI21X1  g11851(.A0(new_n6119_), .A1(new_n5238_), .B0(new_n12041_), .Y(new_n12045_));
  AOI22X1  g11852(.A0(new_n12045_), .A1(new_n12044_), .B0(new_n12043_), .B1(new_n12042_), .Y(new_n12046_));
  XOR2X1   g11853(.A(new_n12046_), .B(new_n12040_), .Y(new_n12047_));
  NAND2X1  g11854(.A(new_n11972_), .B(new_n11968_), .Y(new_n12048_));
  OAI21X1  g11855(.A0(new_n11975_), .A1(new_n11973_), .B0(new_n12048_), .Y(new_n12049_));
  XOR2X1   g11856(.A(new_n12049_), .B(new_n12047_), .Y(new_n12050_));
  XOR2X1   g11857(.A(new_n12050_), .B(new_n12024_), .Y(new_n12051_));
  NOR2X1   g11858(.A(new_n12051_), .B(new_n12011_), .Y(new_n12052_));
  AND2X1   g11859(.A(new_n12051_), .B(new_n12011_), .Y(new_n12053_));
  OR2X1    g11860(.A(new_n12053_), .B(new_n12052_), .Y(new_n12054_));
  XOR2X1   g11861(.A(new_n12054_), .B(new_n12009_), .Y(\asquared[112] ));
  AND2X1   g11862(.A(new_n12049_), .B(new_n12047_), .Y(new_n12056_));
  AOI21X1  g11863(.A0(new_n12050_), .A1(new_n12023_), .B0(new_n12056_), .Y(new_n12057_));
  OR2X1    g11864(.A(new_n12018_), .B(new_n12016_), .Y(new_n12058_));
  OAI21X1  g11865(.A0(new_n12022_), .A1(new_n12020_), .B0(new_n12058_), .Y(new_n12059_));
  AND2X1   g11866(.A(\a[63] ), .B(\a[60] ), .Y(new_n12060_));
  AOI22X1  g11867(.A0(new_n12060_), .A1(\a[52] ), .B0(new_n6688_), .B1(\a[51] ), .Y(new_n12061_));
  AND2X1   g11868(.A(new_n6428_), .B(new_n7164_), .Y(new_n12062_));
  NOR3X1   g11869(.A(new_n12062_), .B(new_n12061_), .C(new_n3915_), .Y(new_n12063_));
  AND2X1   g11870(.A(\a[63] ), .B(\a[49] ), .Y(new_n12064_));
  INVX1    g11871(.A(new_n12064_), .Y(new_n12065_));
  NOR2X1   g11872(.A(new_n12063_), .B(new_n12062_), .Y(new_n12066_));
  INVX1    g11873(.A(new_n12066_), .Y(new_n12067_));
  AOI22X1  g11874(.A0(\a[61] ), .A1(\a[51] ), .B0(\a[60] ), .B1(\a[52] ), .Y(new_n12068_));
  OAI22X1  g11875(.A0(new_n12068_), .A1(new_n12067_), .B0(new_n12065_), .B1(new_n12063_), .Y(new_n12069_));
  XOR2X1   g11876(.A(new_n12069_), .B(new_n12028_), .Y(new_n12070_));
  NAND4X1  g11877(.A(\a[59] ), .B(\a[58] ), .C(\a[54] ), .D(\a[53] ), .Y(new_n12071_));
  NAND4X1  g11878(.A(\a[59] ), .B(\a[57] ), .C(\a[55] ), .D(\a[53] ), .Y(new_n12072_));
  AOI22X1  g11879(.A0(new_n12072_), .A1(new_n12071_), .B0(new_n6119_), .B1(new_n5240_), .Y(new_n12073_));
  NOR3X1   g11880(.A(new_n12073_), .B(new_n5617_), .C(new_n5245_), .Y(new_n12074_));
  AOI21X1  g11881(.A0(new_n6119_), .A1(new_n5240_), .B0(new_n12073_), .Y(new_n12075_));
  OAI22X1  g11882(.A0(new_n5379_), .A1(new_n4835_), .B0(new_n5441_), .B1(new_n4906_), .Y(new_n12076_));
  AOI21X1  g11883(.A0(new_n12076_), .A1(new_n12075_), .B0(new_n12074_), .Y(new_n12077_));
  XOR2X1   g11884(.A(new_n12077_), .B(new_n12070_), .Y(new_n12078_));
  XOR2X1   g11885(.A(new_n12078_), .B(new_n12059_), .Y(new_n12079_));
  XOR2X1   g11886(.A(new_n12036_), .B(new_n11274_), .Y(new_n12080_));
  XOR2X1   g11887(.A(new_n12080_), .B(new_n12045_), .Y(new_n12081_));
  AND2X1   g11888(.A(new_n11985_), .B(new_n11965_), .Y(new_n12082_));
  AOI21X1  g11889(.A0(new_n12014_), .A1(new_n12012_), .B0(new_n12082_), .Y(new_n12083_));
  NAND2X1  g11890(.A(new_n12038_), .B(new_n12032_), .Y(new_n12084_));
  OAI21X1  g11891(.A0(new_n12046_), .A1(new_n12040_), .B0(new_n12084_), .Y(new_n12085_));
  XOR2X1   g11892(.A(new_n12085_), .B(new_n12083_), .Y(new_n12086_));
  XOR2X1   g11893(.A(new_n12086_), .B(new_n12081_), .Y(new_n12087_));
  XOR2X1   g11894(.A(new_n12087_), .B(new_n12079_), .Y(new_n12088_));
  INVX1    g11895(.A(new_n12088_), .Y(new_n12089_));
  NOR2X1   g11896(.A(new_n12089_), .B(new_n12057_), .Y(new_n12090_));
  INVX1    g11897(.A(new_n12090_), .Y(new_n12091_));
  INVX1    g11898(.A(new_n12052_), .Y(new_n12092_));
  OAI21X1  g11899(.A0(new_n12053_), .A1(new_n12009_), .B0(new_n12092_), .Y(new_n12093_));
  AND2X1   g11900(.A(new_n12089_), .B(new_n12057_), .Y(new_n12094_));
  INVX1    g11901(.A(new_n12094_), .Y(new_n12095_));
  AOI21X1  g11902(.A0(new_n12091_), .A1(new_n12095_), .B0(new_n12093_), .Y(new_n12096_));
  AND2X1   g11903(.A(new_n12095_), .B(new_n12093_), .Y(new_n12097_));
  AOI21X1  g11904(.A0(new_n12097_), .A1(new_n12091_), .B0(new_n12096_), .Y(\asquared[113] ));
  AOI21X1  g11905(.A0(new_n12095_), .A1(new_n12093_), .B0(new_n12090_), .Y(new_n12099_));
  AND2X1   g11906(.A(new_n12078_), .B(new_n12059_), .Y(new_n12100_));
  AND2X1   g11907(.A(new_n12087_), .B(new_n12079_), .Y(new_n12101_));
  NAND2X1  g11908(.A(\a[60] ), .B(\a[53] ), .Y(new_n12102_));
  NAND2X1  g11909(.A(\a[61] ), .B(\a[52] ), .Y(new_n12103_));
  AOI22X1  g11910(.A0(new_n12103_), .A1(new_n12102_), .B0(new_n6428_), .B1(new_n5048_), .Y(new_n12104_));
  XOR2X1   g11911(.A(new_n12104_), .B(new_n12075_), .Y(new_n12105_));
  OAI21X1  g11912(.A0(new_n8154_), .A1(new_n5239_), .B0(new_n12042_), .Y(new_n12106_));
  NOR3X1   g11913(.A(new_n12035_), .B(new_n6606_), .C(new_n4983_), .Y(new_n12107_));
  AOI21X1  g11914(.A0(new_n12080_), .A1(new_n12106_), .B0(new_n12107_), .Y(new_n12108_));
  XOR2X1   g11915(.A(new_n12108_), .B(new_n12105_), .Y(new_n12109_));
  NAND2X1  g11916(.A(new_n12069_), .B(new_n12029_), .Y(new_n12110_));
  OAI21X1  g11917(.A0(new_n12077_), .A1(new_n12070_), .B0(new_n12110_), .Y(new_n12111_));
  XOR2X1   g11918(.A(new_n12111_), .B(new_n12109_), .Y(new_n12112_));
  OR2X1    g11919(.A(new_n12046_), .B(new_n12040_), .Y(new_n12113_));
  AOI21X1  g11920(.A0(new_n12113_), .A1(new_n12084_), .B0(new_n12083_), .Y(new_n12114_));
  NOR2X1   g11921(.A(new_n12086_), .B(new_n12081_), .Y(new_n12115_));
  NOR2X1   g11922(.A(new_n12115_), .B(new_n12114_), .Y(new_n12116_));
  AOI22X1  g11923(.A0(\a[59] ), .A1(\a[54] ), .B0(\a[58] ), .B1(\a[55] ), .Y(new_n12117_));
  AND2X1   g11924(.A(\a[63] ), .B(\a[50] ), .Y(new_n12118_));
  AND2X1   g11925(.A(new_n6121_), .B(new_n5240_), .Y(new_n12119_));
  OAI21X1  g11926(.A0(new_n12117_), .A1(new_n12119_), .B0(new_n12118_), .Y(new_n12120_));
  NOR3X1   g11927(.A(new_n12117_), .B(new_n6549_), .C(new_n4983_), .Y(new_n12121_));
  OR2X1    g11928(.A(new_n12121_), .B(new_n12119_), .Y(new_n12122_));
  OAI21X1  g11929(.A0(new_n12122_), .A1(new_n12117_), .B0(new_n12120_), .Y(new_n12123_));
  XOR2X1   g11930(.A(new_n12123_), .B(new_n12066_), .Y(new_n12124_));
  INVX1    g11931(.A(new_n12124_), .Y(new_n12125_));
  NOR4X1   g11932(.A(new_n6606_), .B(new_n5441_), .C(new_n6022_), .D(new_n4349_), .Y(new_n12126_));
  AOI21X1  g11933(.A0(new_n9550_), .A1(\a[62] ), .B0(new_n5554_), .Y(new_n12127_));
  OAI21X1  g11934(.A0(new_n6606_), .A1(new_n4349_), .B0(new_n5441_), .Y(new_n12128_));
  AOI21X1  g11935(.A0(new_n12128_), .A1(new_n12127_), .B0(new_n12126_), .Y(new_n12129_));
  XOR2X1   g11936(.A(new_n12129_), .B(new_n12125_), .Y(new_n12130_));
  XOR2X1   g11937(.A(new_n12130_), .B(new_n12116_), .Y(new_n12131_));
  XOR2X1   g11938(.A(new_n12131_), .B(new_n12112_), .Y(new_n12132_));
  NOR3X1   g11939(.A(new_n12132_), .B(new_n12101_), .C(new_n12100_), .Y(new_n12133_));
  OR2X1    g11940(.A(new_n12101_), .B(new_n12100_), .Y(new_n12134_));
  AND2X1   g11941(.A(new_n12132_), .B(new_n12134_), .Y(new_n12135_));
  OR2X1    g11942(.A(new_n12135_), .B(new_n12133_), .Y(new_n12136_));
  XOR2X1   g11943(.A(new_n12136_), .B(new_n12099_), .Y(\asquared[114] ));
  NOR2X1   g11944(.A(new_n12130_), .B(new_n12116_), .Y(new_n12138_));
  AOI21X1  g11945(.A0(new_n12131_), .A1(new_n12112_), .B0(new_n12138_), .Y(new_n12139_));
  INVX1    g11946(.A(new_n12127_), .Y(new_n12140_));
  XOR2X1   g11947(.A(new_n12140_), .B(new_n12122_), .Y(new_n12141_));
  INVX1    g11948(.A(new_n12141_), .Y(new_n12142_));
  INVX1    g11949(.A(new_n12075_), .Y(new_n12143_));
  AOI22X1  g11950(.A0(new_n12104_), .A1(new_n12143_), .B0(new_n6428_), .B1(new_n5048_), .Y(new_n12144_));
  XOR2X1   g11951(.A(new_n12144_), .B(new_n12142_), .Y(new_n12145_));
  INVX1    g11952(.A(new_n12145_), .Y(new_n12146_));
  NOR2X1   g11953(.A(new_n12108_), .B(new_n12105_), .Y(new_n12147_));
  AOI21X1  g11954(.A0(new_n12111_), .A1(new_n12109_), .B0(new_n12147_), .Y(new_n12148_));
  XOR2X1   g11955(.A(new_n12148_), .B(new_n12146_), .Y(new_n12149_));
  AOI22X1  g11956(.A0(\a[62] ), .A1(\a[52] ), .B0(\a[61] ), .B1(\a[53] ), .Y(new_n12150_));
  NAND4X1  g11957(.A(\a[63] ), .B(\a[62] ), .C(\a[52] ), .D(\a[51] ), .Y(new_n12151_));
  NAND4X1  g11958(.A(\a[63] ), .B(\a[61] ), .C(\a[53] ), .D(\a[51] ), .Y(new_n12152_));
  AOI22X1  g11959(.A0(new_n12152_), .A1(new_n12151_), .B0(new_n6556_), .B1(new_n5048_), .Y(new_n12153_));
  AOI21X1  g11960(.A0(new_n6556_), .A1(new_n5048_), .B0(new_n12153_), .Y(new_n12154_));
  INVX1    g11961(.A(new_n12154_), .Y(new_n12155_));
  NAND2X1  g11962(.A(\a[63] ), .B(\a[51] ), .Y(new_n12156_));
  OAI22X1  g11963(.A0(new_n12156_), .A1(new_n12153_), .B0(new_n12155_), .B1(new_n12150_), .Y(new_n12157_));
  AOI22X1  g11964(.A0(new_n6795_), .A1(new_n5042_), .B0(new_n6427_), .B1(new_n5240_), .Y(new_n12158_));
  AOI21X1  g11965(.A0(new_n6237_), .A1(new_n6121_), .B0(new_n12158_), .Y(new_n12159_));
  AND2X1   g11966(.A(\a[60] ), .B(\a[54] ), .Y(new_n12160_));
  INVX1    g11967(.A(new_n12160_), .Y(new_n12161_));
  OAI22X1  g11968(.A0(new_n6796_), .A1(new_n8559_), .B0(new_n6794_), .B1(new_n5241_), .Y(new_n12162_));
  AOI21X1  g11969(.A0(new_n6237_), .A1(new_n6121_), .B0(new_n12162_), .Y(new_n12163_));
  INVX1    g11970(.A(new_n12163_), .Y(new_n12164_));
  AOI22X1  g11971(.A0(\a[59] ), .A1(\a[55] ), .B0(\a[58] ), .B1(\a[56] ), .Y(new_n12165_));
  OAI22X1  g11972(.A0(new_n12165_), .A1(new_n12164_), .B0(new_n12161_), .B1(new_n12159_), .Y(new_n12166_));
  INVX1    g11973(.A(new_n12166_), .Y(new_n12167_));
  XOR2X1   g11974(.A(new_n12167_), .B(new_n12157_), .Y(new_n12168_));
  NOR2X1   g11975(.A(new_n12129_), .B(new_n12124_), .Y(new_n12169_));
  AOI21X1  g11976(.A0(new_n12123_), .A1(new_n12067_), .B0(new_n12169_), .Y(new_n12170_));
  XOR2X1   g11977(.A(new_n12170_), .B(new_n12168_), .Y(new_n12171_));
  XOR2X1   g11978(.A(new_n12171_), .B(new_n12149_), .Y(new_n12172_));
  INVX1    g11979(.A(new_n12172_), .Y(new_n12173_));
  NOR2X1   g11980(.A(new_n12173_), .B(new_n12139_), .Y(new_n12174_));
  INVX1    g11981(.A(new_n12174_), .Y(new_n12175_));
  INVX1    g11982(.A(new_n12135_), .Y(new_n12176_));
  OAI21X1  g11983(.A0(new_n12133_), .A1(new_n12099_), .B0(new_n12176_), .Y(new_n12177_));
  NAND2X1  g11984(.A(new_n12173_), .B(new_n12139_), .Y(new_n12178_));
  AOI21X1  g11985(.A0(new_n12175_), .A1(new_n12178_), .B0(new_n12177_), .Y(new_n12179_));
  AND2X1   g11986(.A(new_n12178_), .B(new_n12177_), .Y(new_n12180_));
  AOI21X1  g11987(.A0(new_n12180_), .A1(new_n12175_), .B0(new_n12179_), .Y(\asquared[115] ));
  AOI21X1  g11988(.A0(new_n12178_), .A1(new_n12177_), .B0(new_n12174_), .Y(new_n12182_));
  NAND2X1  g11989(.A(new_n12171_), .B(new_n12149_), .Y(new_n12183_));
  OAI21X1  g11990(.A0(new_n12148_), .A1(new_n12146_), .B0(new_n12183_), .Y(new_n12184_));
  NAND3X1  g11991(.A(\a[62] ), .B(\a[58] ), .C(\a[53] ), .Y(new_n12185_));
  AND2X1   g11992(.A(new_n12185_), .B(new_n8154_), .Y(new_n12186_));
  INVX1    g11993(.A(new_n12186_), .Y(new_n12187_));
  AOI21X1  g11994(.A0(\a[62] ), .A1(\a[53] ), .B0(\a[58] ), .Y(new_n12188_));
  NAND4X1  g11995(.A(\a[62] ), .B(\a[58] ), .C(\a[57] ), .D(\a[53] ), .Y(new_n12189_));
  OAI21X1  g11996(.A0(new_n12188_), .A1(new_n12187_), .B0(new_n12189_), .Y(new_n12190_));
  NAND4X1  g11997(.A(\a[61] ), .B(\a[59] ), .C(\a[56] ), .D(\a[54] ), .Y(new_n12191_));
  NAND4X1  g11998(.A(\a[61] ), .B(\a[60] ), .C(\a[55] ), .D(\a[54] ), .Y(new_n12192_));
  AOI22X1  g11999(.A0(new_n12192_), .A1(new_n12191_), .B0(new_n6427_), .B1(new_n6237_), .Y(new_n12193_));
  NAND2X1  g12000(.A(\a[61] ), .B(\a[54] ), .Y(new_n12194_));
  AOI21X1  g12001(.A0(new_n6427_), .A1(new_n6237_), .B0(new_n12193_), .Y(new_n12195_));
  INVX1    g12002(.A(new_n12195_), .Y(new_n12196_));
  AOI22X1  g12003(.A0(\a[60] ), .A1(\a[55] ), .B0(\a[59] ), .B1(\a[56] ), .Y(new_n12197_));
  OAI22X1  g12004(.A0(new_n12197_), .A1(new_n12196_), .B0(new_n12194_), .B1(new_n12193_), .Y(new_n12198_));
  XOR2X1   g12005(.A(new_n12198_), .B(new_n12190_), .Y(new_n12199_));
  NAND2X1  g12006(.A(new_n12140_), .B(new_n12122_), .Y(new_n12200_));
  OAI21X1  g12007(.A0(new_n12144_), .A1(new_n12142_), .B0(new_n12200_), .Y(new_n12201_));
  XOR2X1   g12008(.A(new_n12201_), .B(new_n12199_), .Y(new_n12202_));
  NAND2X1  g12009(.A(\a[63] ), .B(\a[52] ), .Y(new_n12203_));
  XOR2X1   g12010(.A(new_n12203_), .B(new_n12164_), .Y(new_n12204_));
  XOR2X1   g12011(.A(new_n12204_), .B(new_n12154_), .Y(new_n12205_));
  NAND2X1  g12012(.A(new_n12166_), .B(new_n12157_), .Y(new_n12206_));
  OAI21X1  g12013(.A0(new_n12170_), .A1(new_n12168_), .B0(new_n12206_), .Y(new_n12207_));
  XOR2X1   g12014(.A(new_n12207_), .B(new_n12205_), .Y(new_n12208_));
  XOR2X1   g12015(.A(new_n12208_), .B(new_n12202_), .Y(new_n12209_));
  AND2X1   g12016(.A(new_n12209_), .B(new_n12184_), .Y(new_n12210_));
  NOR2X1   g12017(.A(new_n12209_), .B(new_n12184_), .Y(new_n12211_));
  OR2X1    g12018(.A(new_n12211_), .B(new_n12210_), .Y(new_n12212_));
  XOR2X1   g12019(.A(new_n12212_), .B(new_n12182_), .Y(\asquared[116] ));
  AND2X1   g12020(.A(new_n12198_), .B(new_n12190_), .Y(new_n12214_));
  AOI21X1  g12021(.A0(new_n12201_), .A1(new_n12199_), .B0(new_n12214_), .Y(new_n12215_));
  OR2X1    g12022(.A(new_n12203_), .B(new_n12163_), .Y(new_n12216_));
  OAI21X1  g12023(.A0(new_n12204_), .A1(new_n12154_), .B0(new_n12216_), .Y(new_n12217_));
  INVX1    g12024(.A(new_n12217_), .Y(new_n12218_));
  XOR2X1   g12025(.A(new_n12218_), .B(new_n12215_), .Y(new_n12219_));
  AND2X1   g12026(.A(\a[62] ), .B(\a[54] ), .Y(new_n12220_));
  AND2X1   g12027(.A(\a[63] ), .B(\a[53] ), .Y(new_n12221_));
  OAI22X1  g12028(.A0(new_n12221_), .A1(new_n12220_), .B0(new_n7972_), .B1(new_n5239_), .Y(new_n12222_));
  XOR2X1   g12029(.A(new_n12222_), .B(new_n12187_), .Y(new_n12223_));
  NAND4X1  g12030(.A(\a[61] ), .B(\a[59] ), .C(\a[57] ), .D(\a[55] ), .Y(new_n12224_));
  NAND4X1  g12031(.A(\a[61] ), .B(\a[60] ), .C(\a[56] ), .D(\a[55] ), .Y(new_n12225_));
  AOI22X1  g12032(.A0(new_n12225_), .A1(new_n12224_), .B0(new_n6427_), .B1(new_n5554_), .Y(new_n12226_));
  NAND2X1  g12033(.A(\a[61] ), .B(\a[55] ), .Y(new_n12227_));
  AOI21X1  g12034(.A0(new_n6427_), .A1(new_n5554_), .B0(new_n12226_), .Y(new_n12228_));
  INVX1    g12035(.A(new_n12228_), .Y(new_n12229_));
  AOI22X1  g12036(.A0(\a[60] ), .A1(\a[56] ), .B0(\a[59] ), .B1(\a[57] ), .Y(new_n12230_));
  OAI22X1  g12037(.A0(new_n12230_), .A1(new_n12229_), .B0(new_n12227_), .B1(new_n12226_), .Y(new_n12231_));
  AND2X1   g12038(.A(new_n12231_), .B(new_n12195_), .Y(new_n12232_));
  XOR2X1   g12039(.A(new_n12231_), .B(new_n12195_), .Y(new_n12233_));
  OAI21X1  g12040(.A0(new_n12231_), .A1(new_n12195_), .B0(new_n12223_), .Y(new_n12234_));
  OAI22X1  g12041(.A0(new_n12234_), .A1(new_n12232_), .B0(new_n12233_), .B1(new_n12223_), .Y(new_n12235_));
  XOR2X1   g12042(.A(new_n12235_), .B(new_n12219_), .Y(new_n12236_));
  AND2X1   g12043(.A(new_n12207_), .B(new_n12205_), .Y(new_n12237_));
  AOI21X1  g12044(.A0(new_n12208_), .A1(new_n12202_), .B0(new_n12237_), .Y(new_n12238_));
  NOR2X1   g12045(.A(new_n12238_), .B(new_n12236_), .Y(new_n12239_));
  INVX1    g12046(.A(new_n12239_), .Y(new_n12240_));
  INVX1    g12047(.A(new_n12210_), .Y(new_n12241_));
  OAI21X1  g12048(.A0(new_n12211_), .A1(new_n12182_), .B0(new_n12241_), .Y(new_n12242_));
  AND2X1   g12049(.A(new_n12238_), .B(new_n12236_), .Y(new_n12243_));
  INVX1    g12050(.A(new_n12243_), .Y(new_n12244_));
  AOI21X1  g12051(.A0(new_n12240_), .A1(new_n12244_), .B0(new_n12242_), .Y(new_n12245_));
  AND2X1   g12052(.A(new_n12244_), .B(new_n12242_), .Y(new_n12246_));
  AOI21X1  g12053(.A0(new_n12246_), .A1(new_n12240_), .B0(new_n12245_), .Y(\asquared[117] ));
  AOI21X1  g12054(.A0(new_n12244_), .A1(new_n12242_), .B0(new_n12239_), .Y(new_n12248_));
  NOR2X1   g12055(.A(new_n12218_), .B(new_n12215_), .Y(new_n12249_));
  INVX1    g12056(.A(new_n12235_), .Y(new_n12250_));
  AOI21X1  g12057(.A0(new_n12250_), .A1(new_n12219_), .B0(new_n12249_), .Y(new_n12251_));
  OAI22X1  g12058(.A0(new_n12222_), .A1(new_n12186_), .B0(new_n7972_), .B1(new_n5239_), .Y(new_n12252_));
  XOR2X1   g12059(.A(new_n12252_), .B(new_n12228_), .Y(new_n12253_));
  NAND4X1  g12060(.A(\a[63] ), .B(\a[60] ), .C(\a[57] ), .D(\a[54] ), .Y(new_n12254_));
  OAI21X1  g12061(.A0(new_n7973_), .A1(new_n8559_), .B0(new_n12254_), .Y(new_n12255_));
  OAI21X1  g12062(.A0(new_n6554_), .A1(new_n11496_), .B0(new_n12255_), .Y(new_n12256_));
  AND2X1   g12063(.A(\a[63] ), .B(\a[54] ), .Y(new_n12257_));
  OAI22X1  g12064(.A0(new_n6023_), .A1(new_n6022_), .B0(new_n5952_), .B1(new_n5441_), .Y(new_n12258_));
  AOI21X1  g12065(.A0(new_n6428_), .A1(new_n5554_), .B0(new_n12255_), .Y(new_n12259_));
  AOI22X1  g12066(.A0(new_n12259_), .A1(new_n12258_), .B0(new_n12257_), .B1(new_n12256_), .Y(new_n12260_));
  XOR2X1   g12067(.A(new_n12260_), .B(new_n12253_), .Y(new_n12261_));
  AND2X1   g12068(.A(new_n12231_), .B(new_n12196_), .Y(new_n12262_));
  INVX1    g12069(.A(new_n12262_), .Y(new_n12263_));
  OR2X1    g12070(.A(new_n12233_), .B(new_n12223_), .Y(new_n12264_));
  NAND2X1  g12071(.A(new_n12264_), .B(new_n12263_), .Y(new_n12265_));
  NAND4X1  g12072(.A(\a[62] ), .B(\a[59] ), .C(\a[58] ), .D(\a[55] ), .Y(new_n12266_));
  AND2X1   g12073(.A(\a[62] ), .B(\a[59] ), .Y(new_n12267_));
  AOI21X1  g12074(.A0(new_n12267_), .A1(\a[55] ), .B0(new_n6121_), .Y(new_n12268_));
  INVX1    g12075(.A(new_n12268_), .Y(new_n12269_));
  AOI21X1  g12076(.A0(\a[62] ), .A1(\a[55] ), .B0(\a[59] ), .Y(new_n12270_));
  OAI21X1  g12077(.A0(new_n12270_), .A1(new_n12269_), .B0(new_n12266_), .Y(new_n12271_));
  INVX1    g12078(.A(new_n12271_), .Y(new_n12272_));
  XOR2X1   g12079(.A(new_n12272_), .B(new_n12265_), .Y(new_n12273_));
  XOR2X1   g12080(.A(new_n12273_), .B(new_n12261_), .Y(new_n12274_));
  NOR2X1   g12081(.A(new_n12274_), .B(new_n12251_), .Y(new_n12275_));
  AND2X1   g12082(.A(new_n12274_), .B(new_n12251_), .Y(new_n12276_));
  OR2X1    g12083(.A(new_n12276_), .B(new_n12275_), .Y(new_n12277_));
  XOR2X1   g12084(.A(new_n12277_), .B(new_n12248_), .Y(\asquared[118] ));
  AND2X1   g12085(.A(\a[63] ), .B(\a[55] ), .Y(new_n12279_));
  XOR2X1   g12086(.A(new_n12279_), .B(new_n12269_), .Y(new_n12280_));
  INVX1    g12087(.A(new_n12280_), .Y(new_n12281_));
  XOR2X1   g12088(.A(new_n12281_), .B(new_n12259_), .Y(new_n12282_));
  INVX1    g12089(.A(new_n12282_), .Y(new_n12283_));
  AND2X1   g12090(.A(new_n12252_), .B(new_n12229_), .Y(new_n12284_));
  NOR2X1   g12091(.A(new_n12260_), .B(new_n12253_), .Y(new_n12285_));
  NOR2X1   g12092(.A(new_n12285_), .B(new_n12284_), .Y(new_n12286_));
  INVX1    g12093(.A(new_n12286_), .Y(new_n12287_));
  NAND4X1  g12094(.A(\a[62] ), .B(\a[60] ), .C(\a[58] ), .D(\a[56] ), .Y(new_n12288_));
  OAI21X1  g12095(.A0(new_n6557_), .A1(new_n11496_), .B0(new_n12288_), .Y(new_n12289_));
  OAI21X1  g12096(.A0(new_n6554_), .A1(new_n8154_), .B0(new_n12289_), .Y(new_n12290_));
  AOI21X1  g12097(.A0(new_n6428_), .A1(new_n6119_), .B0(new_n12289_), .Y(new_n12291_));
  OAI22X1  g12098(.A0(new_n6023_), .A1(new_n5441_), .B0(new_n5952_), .B1(new_n5379_), .Y(new_n12292_));
  AOI22X1  g12099(.A0(new_n12292_), .A1(new_n12291_), .B0(new_n12290_), .B1(new_n12033_), .Y(new_n12293_));
  XOR2X1   g12100(.A(new_n12293_), .B(new_n12287_), .Y(new_n12294_));
  XOR2X1   g12101(.A(new_n12294_), .B(new_n12283_), .Y(new_n12295_));
  INVX1    g12102(.A(new_n12295_), .Y(new_n12296_));
  AOI21X1  g12103(.A0(new_n12264_), .A1(new_n12263_), .B0(new_n12272_), .Y(new_n12297_));
  INVX1    g12104(.A(new_n12273_), .Y(new_n12298_));
  AOI21X1  g12105(.A0(new_n12298_), .A1(new_n12261_), .B0(new_n12297_), .Y(new_n12299_));
  XOR2X1   g12106(.A(new_n12299_), .B(new_n12296_), .Y(new_n12300_));
  INVX1    g12107(.A(new_n12275_), .Y(new_n12301_));
  OAI21X1  g12108(.A0(new_n12276_), .A1(new_n12248_), .B0(new_n12301_), .Y(new_n12302_));
  XOR2X1   g12109(.A(new_n12302_), .B(new_n12300_), .Y(\asquared[119] ));
  INVX1    g12110(.A(new_n12291_), .Y(new_n12304_));
  NAND2X1  g12111(.A(\a[61] ), .B(\a[58] ), .Y(new_n12305_));
  NAND2X1  g12112(.A(\a[63] ), .B(\a[56] ), .Y(new_n12306_));
  AOI22X1  g12113(.A0(new_n12306_), .A1(new_n12305_), .B0(new_n6688_), .B1(new_n5381_), .Y(new_n12307_));
  XOR2X1   g12114(.A(new_n12307_), .B(new_n12304_), .Y(new_n12308_));
  NAND4X1  g12115(.A(\a[62] ), .B(\a[60] ), .C(\a[59] ), .D(\a[57] ), .Y(new_n12309_));
  AOI21X1  g12116(.A0(new_n6191_), .A1(\a[57] ), .B0(new_n6427_), .Y(new_n12310_));
  INVX1    g12117(.A(new_n12310_), .Y(new_n12311_));
  AOI21X1  g12118(.A0(\a[62] ), .A1(\a[57] ), .B0(\a[60] ), .Y(new_n12312_));
  OAI21X1  g12119(.A0(new_n12312_), .A1(new_n12311_), .B0(new_n12309_), .Y(new_n12313_));
  XOR2X1   g12120(.A(new_n12313_), .B(new_n12308_), .Y(new_n12314_));
  NAND2X1  g12121(.A(new_n12279_), .B(new_n12269_), .Y(new_n12315_));
  OAI21X1  g12122(.A0(new_n12281_), .A1(new_n12259_), .B0(new_n12315_), .Y(new_n12316_));
  XOR2X1   g12123(.A(new_n12316_), .B(new_n12314_), .Y(new_n12317_));
  OR2X1    g12124(.A(new_n12293_), .B(new_n12286_), .Y(new_n12318_));
  OAI21X1  g12125(.A0(new_n12294_), .A1(new_n12283_), .B0(new_n12318_), .Y(new_n12319_));
  AND2X1   g12126(.A(new_n12319_), .B(new_n12317_), .Y(new_n12320_));
  NOR2X1   g12127(.A(new_n12319_), .B(new_n12317_), .Y(new_n12321_));
  OR2X1    g12128(.A(new_n12321_), .B(new_n12320_), .Y(new_n12322_));
  AND2X1   g12129(.A(new_n12299_), .B(new_n12296_), .Y(new_n12323_));
  INVX1    g12130(.A(new_n12323_), .Y(new_n12324_));
  NOR2X1   g12131(.A(new_n12299_), .B(new_n12296_), .Y(new_n12325_));
  AOI21X1  g12132(.A0(new_n12302_), .A1(new_n12324_), .B0(new_n12325_), .Y(new_n12326_));
  XOR2X1   g12133(.A(new_n12326_), .B(new_n12322_), .Y(\asquared[120] ));
  AND2X1   g12134(.A(new_n12313_), .B(new_n12308_), .Y(new_n12328_));
  AOI21X1  g12135(.A0(new_n12316_), .A1(new_n12314_), .B0(new_n12328_), .Y(new_n12329_));
  AOI22X1  g12136(.A0(new_n12307_), .A1(new_n12304_), .B0(new_n6688_), .B1(new_n5381_), .Y(new_n12330_));
  XOR2X1   g12137(.A(new_n12330_), .B(new_n12310_), .Y(new_n12331_));
  OAI22X1  g12138(.A0(new_n7973_), .A1(new_n8155_), .B0(new_n7972_), .B1(new_n8154_), .Y(new_n12332_));
  OAI21X1  g12139(.A0(new_n6557_), .A1(new_n6793_), .B0(new_n12332_), .Y(new_n12333_));
  AND2X1   g12140(.A(\a[63] ), .B(\a[57] ), .Y(new_n12334_));
  AOI21X1  g12141(.A0(new_n6556_), .A1(new_n6121_), .B0(new_n12332_), .Y(new_n12335_));
  OAI22X1  g12142(.A0(new_n6606_), .A1(new_n5379_), .B0(new_n6023_), .B1(new_n5617_), .Y(new_n12336_));
  AOI22X1  g12143(.A0(new_n12336_), .A1(new_n12335_), .B0(new_n12334_), .B1(new_n12333_), .Y(new_n12337_));
  XOR2X1   g12144(.A(new_n12337_), .B(new_n12331_), .Y(new_n12338_));
  NOR2X1   g12145(.A(new_n12338_), .B(new_n12329_), .Y(new_n12339_));
  INVX1    g12146(.A(new_n12339_), .Y(new_n12340_));
  INVX1    g12147(.A(new_n12320_), .Y(new_n12341_));
  OAI21X1  g12148(.A0(new_n12326_), .A1(new_n12321_), .B0(new_n12341_), .Y(new_n12342_));
  AND2X1   g12149(.A(new_n12338_), .B(new_n12329_), .Y(new_n12343_));
  INVX1    g12150(.A(new_n12343_), .Y(new_n12344_));
  AOI21X1  g12151(.A0(new_n12340_), .A1(new_n12344_), .B0(new_n12342_), .Y(new_n12345_));
  AND2X1   g12152(.A(new_n12344_), .B(new_n12342_), .Y(new_n12346_));
  AOI21X1  g12153(.A0(new_n12346_), .A1(new_n12340_), .B0(new_n12345_), .Y(\asquared[121] ));
  AND2X1   g12154(.A(\a[61] ), .B(new_n5952_), .Y(new_n12348_));
  XOR2X1   g12155(.A(new_n12348_), .B(new_n12267_), .Y(new_n12349_));
  AND2X1   g12156(.A(\a[63] ), .B(\a[58] ), .Y(new_n12350_));
  INVX1    g12157(.A(new_n12335_), .Y(new_n12351_));
  XOR2X1   g12158(.A(new_n12351_), .B(new_n12350_), .Y(new_n12352_));
  XOR2X1   g12159(.A(new_n12352_), .B(new_n12349_), .Y(new_n12353_));
  AND2X1   g12160(.A(new_n12330_), .B(new_n12310_), .Y(new_n12354_));
  OR2X1    g12161(.A(new_n12330_), .B(new_n12310_), .Y(new_n12355_));
  OAI21X1  g12162(.A0(new_n12337_), .A1(new_n12354_), .B0(new_n12355_), .Y(new_n12356_));
  NOR2X1   g12163(.A(new_n12356_), .B(new_n12353_), .Y(new_n12357_));
  AND2X1   g12164(.A(new_n12356_), .B(new_n12353_), .Y(new_n12358_));
  OR2X1    g12165(.A(new_n12358_), .B(new_n12357_), .Y(new_n12359_));
  AOI21X1  g12166(.A0(new_n12344_), .A1(new_n12342_), .B0(new_n12339_), .Y(new_n12360_));
  XOR2X1   g12167(.A(new_n12360_), .B(new_n12359_), .Y(\asquared[122] ));
  NAND2X1  g12168(.A(new_n12351_), .B(new_n12350_), .Y(new_n12362_));
  NAND2X1  g12169(.A(new_n12352_), .B(new_n12349_), .Y(new_n12363_));
  AOI22X1  g12170(.A0(\a[63] ), .A1(\a[59] ), .B0(\a[62] ), .B1(\a[60] ), .Y(new_n12364_));
  INVX1    g12171(.A(new_n12364_), .Y(new_n12365_));
  AND2X1   g12172(.A(new_n6789_), .B(new_n6427_), .Y(new_n12366_));
  OAI21X1  g12173(.A0(new_n12267_), .A1(\a[60] ), .B0(\a[61] ), .Y(new_n12367_));
  NOR3X1   g12174(.A(new_n12367_), .B(new_n12366_), .C(new_n12364_), .Y(new_n12368_));
  NOR2X1   g12175(.A(new_n12368_), .B(new_n12366_), .Y(new_n12369_));
  NOR2X1   g12176(.A(new_n12368_), .B(new_n12367_), .Y(new_n12370_));
  AOI21X1  g12177(.A0(new_n12369_), .A1(new_n12365_), .B0(new_n12370_), .Y(new_n12371_));
  AOI21X1  g12178(.A0(new_n12363_), .A1(new_n12362_), .B0(new_n12371_), .Y(new_n12372_));
  INVX1    g12179(.A(new_n12372_), .Y(new_n12373_));
  INVX1    g12180(.A(new_n12358_), .Y(new_n12374_));
  OAI21X1  g12181(.A0(new_n12360_), .A1(new_n12357_), .B0(new_n12374_), .Y(new_n12375_));
  NAND3X1  g12182(.A(new_n12371_), .B(new_n12363_), .C(new_n12362_), .Y(new_n12376_));
  AOI21X1  g12183(.A0(new_n12373_), .A1(new_n12376_), .B0(new_n12375_), .Y(new_n12377_));
  AND2X1   g12184(.A(new_n12376_), .B(new_n12375_), .Y(new_n12378_));
  AOI21X1  g12185(.A0(new_n12378_), .A1(new_n12373_), .B0(new_n12377_), .Y(\asquared[123] ));
  AND2X1   g12186(.A(\a[62] ), .B(new_n6023_), .Y(new_n12380_));
  XOR2X1   g12187(.A(new_n12380_), .B(new_n12060_), .Y(new_n12381_));
  XOR2X1   g12188(.A(new_n12381_), .B(new_n12369_), .Y(new_n12382_));
  AOI21X1  g12189(.A0(new_n12376_), .A1(new_n12375_), .B0(new_n12372_), .Y(new_n12383_));
  XOR2X1   g12190(.A(new_n12383_), .B(new_n12382_), .Y(\asquared[124] ));
  NOR3X1   g12191(.A(new_n12381_), .B(new_n12368_), .C(new_n12366_), .Y(new_n12385_));
  OAI21X1  g12192(.A0(new_n12368_), .A1(new_n12366_), .B0(new_n12381_), .Y(new_n12386_));
  OAI21X1  g12193(.A0(new_n12383_), .A1(new_n12385_), .B0(new_n12386_), .Y(new_n12387_));
  NOR4X1   g12194(.A(new_n6549_), .B(new_n6606_), .C(\a[61] ), .D(new_n5952_), .Y(new_n12388_));
  OR2X1    g12195(.A(new_n6688_), .B(new_n6556_), .Y(new_n12389_));
  NOR2X1   g12196(.A(new_n12389_), .B(new_n12388_), .Y(new_n12390_));
  AOI21X1  g12197(.A0(new_n6688_), .A1(\a[62] ), .B0(new_n12390_), .Y(new_n12391_));
  XOR2X1   g12198(.A(new_n12391_), .B(new_n12387_), .Y(\asquared[125] ));
  OR2X1    g12199(.A(new_n6549_), .B(\a[62] ), .Y(new_n12393_));
  INVX1    g12200(.A(new_n12390_), .Y(new_n12394_));
  AOI22X1  g12201(.A0(new_n12394_), .A1(new_n12387_), .B0(new_n6688_), .B1(\a[62] ), .Y(new_n12395_));
  XOR2X1   g12202(.A(new_n12395_), .B(new_n12393_), .Y(\asquared[126] ));
  AOI21X1  g12203(.A0(new_n12395_), .A1(new_n6606_), .B0(new_n6549_), .Y(\asquared[127] ));
  ZERO     g12204(.Y(\asquared[1] ));
  BUFX1    g12205(.A(\a[0] ), .Y(\asquared[0] ));
endmodule


