//Converted to Combinational , Module name: s298 , Timestamp: 2018-12-03T15:51:01.373071 
module s298 ( G0, G1, G2, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23, G117, G132, G66, G118, G133, G67, n19, n24, n29, n34, n39, n44, n49, n54, n59, n64, n69, n74, n79, n84 );
input G0, G1, G2, G10, G11, G12, G13, G14, G15, G16, G17, G18, G19, G20, G21, G22, G23;
output G117, G132, G66, G118, G133, G67, n19, n24, n29, n34, n39, n44, n49, n54, n59, n64, n69, n74, n79, n84;
wire n52, n53, n54_1, n55, n56, n58, n59_1, n60, n61, n62, n63, n65, n66, n67, n68, n69_1, n71, n72, n73, n74_1, n75, n76, n78, n79_1, n80, n81, n82, n84_1, n85, n86, n87, n88, n89, n90, n92, n93, n94, n95, n96, n97, n99, n100, n102, n103, n104, n105, n106, n108, n109, n110, n111, n113, n114, n115, n117, n118, n120, n121;
NOR2X1   g00(.A(G10), .B(G0), .Y(n19));
INVX1    g01(.A(G10), .Y(n52));
INVX1    g02(.A(G13), .Y(n53));
NOR3X1   g03(.A(n53), .B(G12), .C(n52), .Y(n54_1));
AOI21X1  g04(.A0(G11), .A1(G10), .B0(G0), .Y(n55));
OAI21X1  g05(.A0(G11), .A1(G10), .B0(n55), .Y(n56));
NOR2X1   g06(.A(n56), .B(n54_1), .Y(n24));
INVX1    g07(.A(G11), .Y(n58));
INVX1    g08(.A(G12), .Y(n59_1));
NOR3X1   g09(.A(n59_1), .B(n58), .C(n52), .Y(n60));
NOR2X1   g10(.A(G12), .B(G11), .Y(n61));
INVX1    g11(.A(G0), .Y(n62));
OAI21X1  g12(.A0(G12), .A1(G10), .B0(n62), .Y(n63));
NOR3X1   g13(.A(n63), .B(n61), .C(n60), .Y(n29));
NOR4X1   g14(.A(n59_1), .B(n58), .C(n52), .D(n53), .Y(n65));
NAND3X1  g15(.A(G12), .B(G11), .C(G10), .Y(n66));
AND2X1   g16(.A(n66), .B(n53), .Y(n67));
OR2X1    g17(.A(G12), .B(G11), .Y(n68));
OAI21X1  g18(.A0(n68), .A1(n52), .B0(n62), .Y(n69_1));
NOR3X1   g19(.A(n69_1), .B(n67), .C(n65), .Y(n34));
INVX1    g20(.A(G14), .Y(n71));
NOR4X1   g21(.A(n71), .B(n53), .C(n52), .D(n68), .Y(n72));
INVX1    g22(.A(G23), .Y(n73));
OAI21X1  g23(.A0(n73), .A1(n71), .B0(n62), .Y(n74_1));
NOR3X1   g24(.A(n68), .B(n53), .C(n52), .Y(n75));
NOR3X1   g25(.A(n75), .B(G23), .C(G14), .Y(n76));
NOR3X1   g26(.A(n76), .B(n74_1), .C(n72), .Y(n39));
NAND2X1  g27(.A(n59_1), .B(G11), .Y(n78));
INVX1    g28(.A(G22), .Y(n79_1));
NAND3X1  g29(.A(n79_1), .B(n71), .C(G13), .Y(n80));
NOR4X1   g30(.A(n79_1), .B(G14), .C(n53), .D(n68), .Y(n81));
OAI22X1  g31(.A0(n80), .A1(n78), .B0(G15), .B1(n81), .Y(n82));
NOR2X1   g32(.A(n82), .B(G0), .Y(n44));
INVX1    g33(.A(G15), .Y(n84_1));
NOR2X1   g34(.A(G12), .B(n58), .Y(n85));
NOR3X1   g35(.A(G22), .B(G14), .C(n53), .Y(n86));
NAND4X1  g36(.A(G22), .B(n71), .C(G13), .D(n61), .Y(n87));
AOI22X1  g37(.A0(n86), .A1(n85), .B0(n84_1), .B1(n87), .Y(n88));
OAI21X1  g38(.A0(n71), .A1(n59_1), .B0(n53), .Y(n89));
OAI21X1  g39(.A0(G16), .A1(n71), .B0(n89), .Y(n90));
NOR2X1   g40(.A(n90), .B(n88), .Y(n49));
NAND2X1  g41(.A(G14), .B(G12), .Y(n92));
NOR2X1   g42(.A(n92), .B(G17), .Y(n93));
AOI21X1  g43(.A0(G17), .A1(G14), .B0(n53), .Y(n94));
NOR3X1   g44(.A(n68), .B(n71), .C(G13), .Y(n95));
NOR3X1   g45(.A(G14), .B(n59_1), .C(n58), .Y(n96));
OR4X1    g46(.A(n95), .B(n94), .C(n93), .D(n96), .Y(n97));
NOR2X1   g47(.A(n97), .B(n88), .Y(n54));
NOR2X1   g48(.A(n92), .B(G18), .Y(n99));
AOI21X1  g49(.A0(G18), .A1(G14), .B0(n53), .Y(n100));
NOR4X1   g50(.A(n99), .B(n95), .C(n88), .D(n100), .Y(n59));
NOR4X1   g51(.A(G19), .B(n71), .C(n53), .D(n88), .Y(n102));
NAND3X1  g52(.A(G19), .B(G14), .C(G12), .Y(n103));
NAND2X1  g53(.A(n103), .B(n53), .Y(n104));
AOI21X1  g54(.A0(n61), .A1(G14), .B0(n104), .Y(n105));
MX2X1    g55(.A(G10), .B(n105), .S0(n82), .Y(n106));
NOR2X1   g56(.A(n106), .B(n102), .Y(n64));
NOR3X1   g57(.A(G13), .B(G12), .C(n58), .Y(n108));
NOR2X1   g58(.A(G20), .B(n53), .Y(n109));
OAI21X1  g59(.A0(G20), .A1(n59_1), .B0(G14), .Y(n110));
NOR3X1   g60(.A(n110), .B(n109), .C(n108), .Y(n111));
MX2X1    g61(.A(n52), .B(n111), .S0(n82), .Y(n69));
INVX1    g62(.A(G21), .Y(n113));
MX2X1    g63(.A(n58), .B(n113), .S0(G14), .Y(n114));
MX2X1    g64(.A(n59_1), .B(n71), .S0(G13), .Y(n115));
NOR3X1   g65(.A(n115), .B(n114), .C(n88), .Y(n74));
OR2X1    g66(.A(G22), .B(G2), .Y(n117));
AOI21X1  g67(.A0(G22), .A1(G2), .B0(G0), .Y(n118));
AND2X1   g68(.A(n118), .B(n117), .Y(n79));
OR2X1    g69(.A(G23), .B(G1), .Y(n120));
AOI21X1  g70(.A0(G23), .A1(G1), .B0(G0), .Y(n121));
AND2X1   g71(.A(n121), .B(n120), .Y(n84));
BUFX1    g72(.A(G18), .Y(G117));
BUFX1    g73(.A(G20), .Y(G132));
BUFX1    g74(.A(G16), .Y(G66));
BUFX1    g75(.A(G19), .Y(G118));
BUFX1    g76(.A(G21), .Y(G133));
BUFX1    g77(.A(G17), .Y(G67));
endmodule
