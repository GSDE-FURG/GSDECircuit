//Converted to Combinational , Module name: s400 , Timestamp: 2018-12-03T15:51:01.558102 
module s400 ( FM, TEST, CLR, TESTL, FML, OLATCH_Y2L, OLATCHVUC_6, OLATCHVUC_5, OLATCH_R1L, OLATCH_G2L, OLATCH_G1L, OLATCH_FEL, C3_Q3, C3_Q2, C3_Q1, C3_Q0, UC_16, UC_17, UC_18, UC_19, UC_8, UC_9, UC_10, UC_11, GRN2, YLW2, RED2, GRN1, YLW1, RED1, n19, n24, n29, n34, n39, n44, n49, n54, n59, n64, n69, n74, n79, n84, n89, n94, n99, n104, n109, n114, n119 );
input FM, TEST, CLR, TESTL, FML, OLATCH_Y2L, OLATCHVUC_6, OLATCHVUC_5, OLATCH_R1L, OLATCH_G2L, OLATCH_G1L, OLATCH_FEL, C3_Q3, C3_Q2, C3_Q1, C3_Q0, UC_16, UC_17, UC_18, UC_19, UC_8, UC_9, UC_10, UC_11;
output GRN2, YLW2, RED2, GRN1, YLW1, RED1, n19, n24, n29, n34, n39, n44, n49, n54, n59, n64, n69, n74, n79, n84, n89, n94, n99, n104, n109, n114, n119;
wire n74_1, n75, n77, n79_1, n80, n81, n83, n84_1, n85, n86, n87, n88, n89_1, n90, n91, n92, n93, n94_1, n95, n96, n97, n99_1, n100, n101, n103, n104_1, n106, n107, n109_1, n110, n111, n114_1, n115, n116, n117, n118, n119_1, n120, n121, n122, n123, n124, n125, n126, n127, n128, n130, n131, n132, n134, n135, n137, n139, n140, n141, n142, n143, n145, n146, n148, n149, n151, n153, n154, n155, n156, n158, n160;
INVX1    g00(.A(OLATCHVUC_5), .Y(RED2));
INVX1    g01(.A(OLATCHVUC_6), .Y(YLW1));
INVX1    g02(.A(CLR), .Y(n74_1));
OAI21X1  g03(.A0(TESTL), .A1(TEST), .B0(n74_1), .Y(n75));
AOI21X1  g04(.A0(TESTL), .A1(TEST), .B0(n75), .Y(n19));
OAI21X1  g05(.A0(FML), .A1(FM), .B0(n74_1), .Y(n77));
AOI21X1  g06(.A0(FML), .A1(FM), .B0(n77), .Y(n24));
INVX1    g07(.A(C3_Q1), .Y(n79_1));
INVX1    g08(.A(C3_Q0), .Y(n80));
OR2X1    g09(.A(C3_Q2), .B(CLR), .Y(n81));
NOR4X1   g10(.A(n80), .B(n79_1), .C(OLATCH_FEL), .D(n81), .Y(n29));
INVX1    g11(.A(UC_17), .Y(n83));
NAND2X1  g12(.A(OLATCH_FEL), .B(n74_1), .Y(n84_1));
NOR2X1   g13(.A(n80), .B(C3_Q1), .Y(n85));
INVX1    g14(.A(C3_Q2), .Y(n86));
NOR3X1   g15(.A(n86), .B(C3_Q3), .C(FML), .Y(n87));
AOI21X1  g16(.A0(n87), .A1(n85), .B0(n84_1), .Y(n88));
INVX1    g17(.A(FML), .Y(n89_1));
NAND2X1  g18(.A(C3_Q2), .B(n74_1), .Y(n90));
NOR4X1   g19(.A(C3_Q0), .B(C3_Q1), .C(n89_1), .D(n90), .Y(n91));
NOR2X1   g20(.A(n91), .B(n88), .Y(n92));
INVX1    g21(.A(C3_Q3), .Y(n93));
OR2X1    g22(.A(n81), .B(n93), .Y(n94_1));
NAND4X1  g23(.A(n93), .B(FML), .C(n74_1), .D(C3_Q2), .Y(n95));
OR2X1    g24(.A(C3_Q0), .B(C3_Q1), .Y(n96));
AOI21X1  g25(.A0(n95), .A1(n94_1), .B0(n96), .Y(n97));
OAI22X1  g26(.A0(n92), .A1(n83), .B0(n88), .B1(n97), .Y(n34));
NOR3X1   g27(.A(n96), .B(n93), .C(CLR), .Y(n99_1));
INVX1    g28(.A(OLATCH_FEL), .Y(n100));
AOI21X1  g29(.A0(n86), .A1(n100), .B0(CLR), .Y(n101));
OAI22X1  g30(.A0(n99_1), .A1(n101), .B0(n92), .B1(n83), .Y(n39));
NAND3X1  g31(.A(n86), .B(n93), .C(n100), .Y(n103));
NAND4X1  g32(.A(n79_1), .B(n86), .C(n100), .D(C3_Q0), .Y(n104_1));
NAND3X1  g33(.A(n104_1), .B(n103), .C(n74_1), .Y(n44));
NOR3X1   g34(.A(C3_Q0), .B(n93), .C(CLR), .Y(n106));
NOR3X1   g35(.A(n80), .B(n79_1), .C(CLR), .Y(n107));
NOR3X1   g36(.A(n107), .B(n106), .C(n101), .Y(n49));
NAND4X1  g37(.A(n79_1), .B(n93), .C(n89_1), .D(C3_Q0), .Y(n109_1));
AOI21X1  g38(.A0(C3_Q3), .A1(FML), .B0(n90), .Y(n110));
OAI21X1  g39(.A0(n96), .A1(n89_1), .B0(n110), .Y(n111));
AOI21X1  g40(.A0(n109_1), .A1(OLATCH_FEL), .B0(n111), .Y(n54));
OR2X1    g41(.A(n91), .B(n88), .Y(n59));
INVX1    g42(.A(TESTL), .Y(n114_1));
INVX1    g43(.A(UC_8), .Y(n115));
NOR3X1   g44(.A(UC_11), .B(UC_10), .C(UC_9), .Y(n116));
OAI21X1  g45(.A0(n116), .A1(n115), .B0(n114_1), .Y(n117));
INVX1    g46(.A(UC_16), .Y(n118));
NOR3X1   g47(.A(UC_19), .B(UC_18), .C(UC_17), .Y(n119_1));
NOR2X1   g48(.A(n119_1), .B(n118), .Y(n120));
NAND2X1  g49(.A(n120), .B(n117), .Y(n121));
NAND2X1  g50(.A(C3_Q0), .B(C3_Q1), .Y(n122));
NOR4X1   g51(.A(n121), .B(n86), .C(n93), .D(n122), .Y(n123));
AND2X1   g52(.A(n120), .B(n117), .Y(n124));
NOR2X1   g53(.A(n122), .B(n86), .Y(n125));
AOI21X1  g54(.A0(n125), .A1(n124), .B0(C3_Q3), .Y(n126));
OAI21X1  g55(.A0(n96), .A1(C3_Q2), .B0(C3_Q3), .Y(n127));
OAI21X1  g56(.A0(n127), .A1(n121), .B0(n74_1), .Y(n128));
NOR3X1   g57(.A(n128), .B(n126), .C(n123), .Y(n64));
NOR3X1   g58(.A(n122), .B(n121), .C(n86), .Y(n130));
INVX1    g59(.A(n122), .Y(n131));
AOI21X1  g60(.A0(n131), .A1(n124), .B0(C3_Q2), .Y(n132));
NOR3X1   g61(.A(n132), .B(n130), .C(n128), .Y(n69));
NOR3X1   g62(.A(n121), .B(n80), .C(n79_1), .Y(n134));
AOI21X1  g63(.A0(n124), .A1(C3_Q0), .B0(C3_Q1), .Y(n135));
NOR3X1   g64(.A(n135), .B(n134), .C(n128), .Y(n74));
XOR2X1   g65(.A(n121), .B(C3_Q0), .Y(n137));
NOR2X1   g66(.A(n137), .B(n128), .Y(n79));
AND2X1   g67(.A(UC_19), .B(UC_18), .Y(n139));
AND2X1   g68(.A(n139), .B(UC_17), .Y(n140));
AND2X1   g69(.A(n140), .B(n117), .Y(n141));
AOI21X1  g70(.A0(n120), .A1(n117), .B0(CLR), .Y(n142));
OAI21X1  g71(.A0(n141), .A1(UC_16), .B0(n142), .Y(n143));
AOI21X1  g72(.A0(n141), .A1(UC_16), .B0(n143), .Y(n84));
AND2X1   g73(.A(n139), .B(n117), .Y(n145));
OAI21X1  g74(.A0(n145), .A1(UC_17), .B0(n142), .Y(n146));
AOI21X1  g75(.A0(n145), .A1(UC_17), .B0(n146), .Y(n89));
AND2X1   g76(.A(n117), .B(UC_19), .Y(n148));
OAI21X1  g77(.A0(n148), .A1(UC_18), .B0(n142), .Y(n149));
AOI21X1  g78(.A0(n148), .A1(UC_18), .B0(n149), .Y(n94));
XOR2X1   g79(.A(n117), .B(UC_19), .Y(n151));
AND2X1   g80(.A(n151), .B(n142), .Y(n99));
NOR2X1   g81(.A(n116), .B(n115), .Y(n153));
AND2X1   g82(.A(UC_11), .B(UC_10), .Y(n154));
AND2X1   g83(.A(n154), .B(UC_9), .Y(n155));
XOR2X1   g84(.A(n155), .B(n115), .Y(n156));
NOR3X1   g85(.A(n156), .B(n153), .C(CLR), .Y(n104));
AOI21X1  g86(.A0(UC_11), .A1(UC_10), .B0(UC_9), .Y(n158));
NOR4X1   g87(.A(n155), .B(n153), .C(CLR), .D(n158), .Y(n109));
NOR2X1   g88(.A(UC_11), .B(UC_10), .Y(n160));
NOR4X1   g89(.A(n153), .B(n160), .C(CLR), .D(n154), .Y(n114));
NOR3X1   g90(.A(n153), .B(UC_11), .C(CLR), .Y(n119));
BUFX1    g91(.A(OLATCH_G2L), .Y(GRN2));
BUFX1    g92(.A(OLATCH_Y2L), .Y(YLW2));
BUFX1    g93(.A(OLATCH_G1L), .Y(GRN1));
BUFX1    g94(.A(OLATCH_R1L), .Y(RED1));
endmodule
