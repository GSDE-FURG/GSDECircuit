// Benchmark "top" written by ABC on Mon Sep 21 04:06:26 2020

module top ( 
    \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] ,
    \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] ,
    \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] ,
    \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] ,
    \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] ,
    \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] ,
    \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] ,
    \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] ,
    \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] ,
    \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] ,
    \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] ,
    \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] ,
    \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] ,
    \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] ,
    \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] ,
    \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] ,
    \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] ,
    \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] ,
    \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] ,
    \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] ,
    \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] ,
    \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] ,
    \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] ,
    \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] ,
    \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] ,
    \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] ,
    \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] ,
    \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] ,
    \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] ,
    \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] ,
    \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] ,
    \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] ,
    \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] ,
    \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] ,
    \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] ,
    \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] ,
    \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] ,
    \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] ,
    \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] ,
    \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] ,
    \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] ,
    \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] ,
    \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] ,
    \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] ,
    \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] ,
    \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] ,
    \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] ,
    \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] ,
    \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] ,
    \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] ,
    \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] ,
    \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] ,
    \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] ,
    \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] ,
    \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] ,
    \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] ,
    \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] ,
    \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] ,
    \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] ,
    \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] ,
    \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] ,
    \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] ,
    \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] ,
    \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] ,
    \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] ,
    \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] ,
    \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] ,
    \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] ,
    \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] ,
    \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] ,
    \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] ,
    \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] ,
    \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] ,
    \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] ,
    \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] ,
    \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] ,
    \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] ,
    \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] ,
    \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] ,
    \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] ,
    \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] ,
    \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] ,
    \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] ,
    \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] ,
    \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] ,
    \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] ,
    \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] ,
    \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] ,
    \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] ,
    \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] ,
    \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] ,
    \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] ,
    \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] ,
    \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] ,
    \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] ,
    \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] ,
    \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] ,
    \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] ,
    \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] ,
    \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] ,
    \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] ,
    \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] ,
    \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] ,
    \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] ,
    \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] ,
    \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] ,
    \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] ,
    \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] ,
    \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] ,
    \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] ,
    \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] ,
    \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] ,
    \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] ,
    \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] ,
    \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] ,
    \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] ,
    \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] ,
    \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] ,
    \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] ,
    \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] ,
    \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] ,
    \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] ,
    \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] ,
    \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] ,
    \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] ,
    \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] ,
    \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] ,
    \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] ,
    \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] ,
    \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] ,
    \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] ,
    \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] ,
    \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] ,
    \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] ,
    \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] ,
    \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] ,
    \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] ,
    \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] ,
    \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] ,
    \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] ,
    \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] ,
    \A[1000] ,
    maj  );
  input  \A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] ,
    \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] ,
    \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] ,
    \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] ,
    \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] ,
    \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] ,
    \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] ,
    \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] ,
    \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] ,
    \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] ,
    \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] ,
    \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] ,
    \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] ,
    \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] ,
    \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] ,
    \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] ,
    \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] ,
    \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] ,
    \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] ,
    \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] ,
    \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] ,
    \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] ,
    \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] ,
    \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] ,
    \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] ,
    \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] ,
    \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] ,
    \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] ,
    \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] ,
    \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] ,
    \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] ,
    \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] ,
    \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] ,
    \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] ,
    \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] ,
    \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] ,
    \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] ,
    \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] ,
    \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] ,
    \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] ,
    \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] ,
    \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] ,
    \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] ,
    \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] ,
    \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] ,
    \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] ,
    \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] ,
    \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] ,
    \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] ,
    \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] ,
    \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] ,
    \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] ,
    \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] ,
    \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] ,
    \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] ,
    \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] ,
    \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] ,
    \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] ,
    \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] ,
    \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] ,
    \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] ,
    \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] ,
    \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] ,
    \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] ,
    \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] ,
    \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] ,
    \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] ,
    \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] ,
    \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] ,
    \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] ,
    \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] ,
    \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] ,
    \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] ,
    \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] ,
    \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] ,
    \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] ,
    \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] ,
    \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] ,
    \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] ,
    \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] ,
    \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] ,
    \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] ,
    \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] ,
    \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] ,
    \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] ,
    \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] ,
    \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] ,
    \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] ,
    \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] ,
    \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] ,
    \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] ,
    \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] ,
    \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] ,
    \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] ,
    \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] ,
    \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] ,
    \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] ,
    \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] ,
    \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] ,
    \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] ,
    \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] ,
    \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] ,
    \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] ,
    \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] ,
    \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] ,
    \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] ,
    \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] ,
    \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] ,
    \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] ,
    \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] ,
    \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] ,
    \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] ,
    \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] ,
    \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] ,
    \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] ,
    \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] ,
    \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] ,
    \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] ,
    \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] ,
    \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] ,
    \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] ,
    \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] ,
    \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] ,
    \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] ,
    \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] ,
    \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] ,
    \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] ,
    \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] ,
    \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] ,
    \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] ,
    \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] ,
    \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] ,
    \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] ,
    \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] ,
    \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] ,
    \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] ,
    \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] ,
    \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] ,
    \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] ,
    \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] ,
    \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] ,
    \A[999] , \A[1000] ;
  output maj;
  wire new_n1003_, new_n1004_, new_n1005_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_, new_n1013_,
    new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_,
    new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_,
    new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_, new_n1031_,
    new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_, new_n1037_,
    new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_, new_n1043_,
    new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_, new_n1049_,
    new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_,
    new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_,
    new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_,
    new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_,
    new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_,
    new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_,
    new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_,
    new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_,
    new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_,
    new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_,
    new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_,
    new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_,
    new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_,
    new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_,
    new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_, new_n1229_,
    new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_, new_n1235_,
    new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_, new_n1241_,
    new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_, new_n1247_,
    new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_, new_n1253_,
    new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_, new_n1259_,
    new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_, new_n1265_,
    new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_, new_n1271_,
    new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_, new_n1277_,
    new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_, new_n1283_,
    new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_, new_n1289_,
    new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_, new_n1295_,
    new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_, new_n1301_,
    new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_, new_n1307_,
    new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_, new_n1313_,
    new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_, new_n1319_,
    new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_, new_n1325_,
    new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_, new_n1331_,
    new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_, new_n1337_,
    new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_, new_n1343_,
    new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_, new_n1349_,
    new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_, new_n1355_,
    new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_, new_n1361_,
    new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_, new_n1367_,
    new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_, new_n1373_,
    new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_, new_n1379_,
    new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_, new_n1385_,
    new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_, new_n1391_,
    new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_, new_n1397_,
    new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_, new_n1403_,
    new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_, new_n1409_,
    new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_, new_n1415_,
    new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_, new_n1421_,
    new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_, new_n1427_,
    new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_, new_n1433_,
    new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_, new_n1439_,
    new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_, new_n1445_,
    new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_, new_n1451_,
    new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_, new_n1457_,
    new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_, new_n1463_,
    new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_, new_n1469_,
    new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_, new_n1475_,
    new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_, new_n1481_,
    new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_, new_n1487_,
    new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_, new_n1493_,
    new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_, new_n1499_,
    new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_, new_n1505_,
    new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_, new_n1511_,
    new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_, new_n1517_,
    new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_, new_n1523_,
    new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_, new_n1529_,
    new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_, new_n1535_,
    new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_, new_n1541_,
    new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_, new_n1547_,
    new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_, new_n1553_,
    new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_, new_n1559_,
    new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_, new_n1565_,
    new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_, new_n1571_,
    new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_, new_n1577_,
    new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_, new_n1685_,
    new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_,
    new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_,
    new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_,
    new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_,
    new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_,
    new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_,
    new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_,
    new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_,
    new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_,
    new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_,
    new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_,
    new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_,
    new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_,
    new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_,
    new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_,
    new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_,
    new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_,
    new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_, new_n1793_,
    new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_, new_n1799_,
    new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_, new_n1805_,
    new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_, new_n1811_,
    new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_, new_n1817_,
    new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_, new_n1823_,
    new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_, new_n1829_,
    new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_, new_n1835_,
    new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_, new_n1841_,
    new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_, new_n1847_,
    new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_, new_n1853_,
    new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_, new_n1859_,
    new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_, new_n1865_,
    new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_, new_n1871_,
    new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_, new_n1877_,
    new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_, new_n1883_,
    new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_, new_n1889_,
    new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_, new_n1895_,
    new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_, new_n1901_,
    new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_, new_n1907_,
    new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_, new_n1913_,
    new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_, new_n1919_,
    new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_, new_n1925_,
    new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_, new_n1931_,
    new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_, new_n1937_,
    new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_, new_n1943_,
    new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_, new_n1949_,
    new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_, new_n1955_,
    new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_, new_n1961_,
    new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_, new_n1967_,
    new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_, new_n1973_,
    new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_, new_n1979_,
    new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_, new_n1985_,
    new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_, new_n1991_,
    new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_, new_n1997_,
    new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_, new_n2003_,
    new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_, new_n2009_,
    new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_, new_n2015_,
    new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_, new_n2021_,
    new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_, new_n2027_,
    new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_, new_n2033_,
    new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_, new_n2039_,
    new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_, new_n2045_,
    new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_, new_n2051_,
    new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_, new_n2057_,
    new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_, new_n2063_,
    new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_, new_n2069_,
    new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_, new_n2075_,
    new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_, new_n2081_,
    new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_, new_n2087_,
    new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_, new_n2093_,
    new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_, new_n2099_,
    new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_, new_n2105_,
    new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_, new_n2111_,
    new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_, new_n2117_,
    new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_, new_n2123_,
    new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_, new_n2129_,
    new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_, new_n2135_,
    new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_, new_n2141_,
    new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_, new_n2147_,
    new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_, new_n2153_,
    new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_, new_n2159_,
    new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_, new_n2165_,
    new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_, new_n2171_,
    new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_, new_n2177_,
    new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_, new_n2183_,
    new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_, new_n2189_,
    new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_, new_n2195_,
    new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_, new_n2201_,
    new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_, new_n2207_,
    new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_, new_n2213_,
    new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_, new_n2219_,
    new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_, new_n2225_,
    new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_, new_n2231_,
    new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_, new_n2237_,
    new_n2238_, new_n2239_, new_n2240_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2369_,
    new_n2370_, new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_,
    new_n2376_, new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_,
    new_n2382_, new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_,
    new_n2388_, new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_,
    new_n2394_, new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_,
    new_n2400_, new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_,
    new_n2406_, new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_,
    new_n2412_, new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_,
    new_n2418_, new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_,
    new_n2424_, new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_,
    new_n2430_, new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_,
    new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_,
    new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_,
    new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_,
    new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_,
    new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_,
    new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_,
    new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_,
    new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_,
    new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_,
    new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_,
    new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_,
    new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_,
    new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_, new_n2513_,
    new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_, new_n2519_,
    new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_, new_n2525_,
    new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_, new_n2531_,
    new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_, new_n2537_,
    new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_, new_n2543_,
    new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_, new_n2549_,
    new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_, new_n2555_,
    new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_, new_n2561_,
    new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_, new_n2567_,
    new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_, new_n2573_,
    new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_, new_n2579_,
    new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_, new_n2651_,
    new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_,
    new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_,
    new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_,
    new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_,
    new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_,
    new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_,
    new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_,
    new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_,
    new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_,
    new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2711_,
    new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_, new_n2717_,
    new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_, new_n2723_,
    new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_, new_n2729_,
    new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_, new_n2735_,
    new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_, new_n2741_,
    new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_, new_n2747_,
    new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_, new_n2753_,
    new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_, new_n2759_,
    new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_, new_n2765_,
    new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_, new_n2771_,
    new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_, new_n2777_,
    new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_, new_n2783_,
    new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_, new_n2789_,
    new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_, new_n2795_,
    new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_, new_n2801_,
    new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_, new_n2807_,
    new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_, new_n2813_,
    new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_, new_n2819_,
    new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_, new_n2825_,
    new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_, new_n2831_,
    new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_, new_n2837_,
    new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_, new_n2843_,
    new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_, new_n2849_,
    new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_, new_n2855_,
    new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_, new_n2861_,
    new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_, new_n2867_,
    new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_, new_n2873_,
    new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_, new_n2879_,
    new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_, new_n2885_,
    new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_, new_n2891_,
    new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_, new_n2897_,
    new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_, new_n2903_,
    new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_, new_n2909_,
    new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_, new_n2915_,
    new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_, new_n2921_,
    new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_, new_n2927_,
    new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_, new_n2933_,
    new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_, new_n2939_,
    new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_, new_n2945_,
    new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_, new_n2951_,
    new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_, new_n2957_,
    new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_, new_n2963_,
    new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_, new_n2969_,
    new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3300_, new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_,
    new_n3306_, new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_,
    new_n3312_, new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_,
    new_n3318_, new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_,
    new_n3324_, new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_,
    new_n3330_, new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_,
    new_n3336_, new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_,
    new_n3342_, new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_,
    new_n3348_, new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_,
    new_n3354_, new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_,
    new_n3360_, new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_,
    new_n3366_, new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_,
    new_n3372_, new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_,
    new_n3378_, new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_,
    new_n3384_, new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_,
    new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_,
    new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_,
    new_n3402_, new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_,
    new_n3414_, new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_,
    new_n3420_, new_n3421_, new_n3422_, new_n3423_, new_n3424_, new_n3425_,
    new_n3426_, new_n3427_, new_n3428_, new_n3429_, new_n3430_, new_n3431_,
    new_n3432_, new_n3433_, new_n3434_, new_n3435_, new_n3436_, new_n3437_,
    new_n3438_, new_n3439_, new_n3440_, new_n3441_, new_n3442_, new_n3443_,
    new_n3444_, new_n3445_, new_n3446_, new_n3447_, new_n3448_, new_n3449_,
    new_n3450_, new_n3451_, new_n3452_, new_n3453_, new_n3454_, new_n3455_,
    new_n3456_, new_n3457_, new_n3458_, new_n3459_, new_n3460_, new_n3461_,
    new_n3462_, new_n3463_, new_n3464_, new_n3465_, new_n3466_, new_n3467_,
    new_n3468_, new_n3469_, new_n3470_, new_n3471_, new_n3472_, new_n3473_,
    new_n3474_, new_n3475_, new_n3476_, new_n3477_, new_n3478_, new_n3479_,
    new_n3480_, new_n3481_, new_n3482_, new_n3483_, new_n3484_, new_n3485_,
    new_n3486_, new_n3487_, new_n3488_, new_n3489_, new_n3490_, new_n3491_,
    new_n3492_, new_n3493_, new_n3494_, new_n3495_, new_n3496_, new_n3497_,
    new_n3498_, new_n3499_, new_n3500_, new_n3501_, new_n3502_, new_n3503_,
    new_n3504_, new_n3505_, new_n3506_, new_n3507_, new_n3508_, new_n3509_,
    new_n3510_, new_n3511_, new_n3512_, new_n3513_, new_n3514_, new_n3515_,
    new_n3516_, new_n3517_, new_n3518_, new_n3519_, new_n3520_, new_n3521_,
    new_n3522_, new_n3523_, new_n3524_, new_n3525_, new_n3526_, new_n3527_,
    new_n3528_, new_n3529_, new_n3530_, new_n3531_, new_n3532_, new_n3533_,
    new_n3534_, new_n3535_, new_n3536_, new_n3537_, new_n3538_, new_n3539_,
    new_n3540_, new_n3541_, new_n3542_, new_n3543_, new_n3544_, new_n3545_,
    new_n3546_, new_n3547_, new_n3548_, new_n3549_, new_n3550_, new_n3551_,
    new_n3552_, new_n3553_, new_n3554_, new_n3555_, new_n3556_, new_n3557_,
    new_n3558_, new_n3559_, new_n3560_, new_n3561_, new_n3562_, new_n3563_,
    new_n3564_, new_n3565_, new_n3566_, new_n3567_, new_n3568_, new_n3569_,
    new_n3570_, new_n3571_, new_n3572_, new_n3573_, new_n3574_, new_n3575_,
    new_n3576_, new_n3577_, new_n3578_, new_n3579_, new_n3580_, new_n3581_,
    new_n3582_, new_n3583_, new_n3584_, new_n3585_, new_n3586_, new_n3587_,
    new_n3588_, new_n3589_, new_n3590_, new_n3591_, new_n3592_, new_n3593_,
    new_n3594_, new_n3595_, new_n3596_, new_n3597_, new_n3598_, new_n3599_,
    new_n3600_, new_n3601_, new_n3602_, new_n3603_, new_n3604_, new_n3605_,
    new_n3606_, new_n3607_, new_n3608_, new_n3609_, new_n3610_, new_n3611_,
    new_n3612_, new_n3613_, new_n3614_, new_n3615_, new_n3616_, new_n3617_,
    new_n3618_, new_n3619_, new_n3620_, new_n3621_, new_n3622_, new_n3623_,
    new_n3624_, new_n3625_, new_n3626_, new_n3627_, new_n3628_, new_n3629_,
    new_n3630_, new_n3631_, new_n3632_, new_n3633_, new_n3634_, new_n3635_,
    new_n3636_, new_n3637_, new_n3638_, new_n3639_, new_n3640_, new_n3641_,
    new_n3642_, new_n3643_, new_n3644_, new_n3645_, new_n3646_, new_n3647_,
    new_n3648_, new_n3649_, new_n3650_, new_n3651_, new_n3652_, new_n3653_,
    new_n3654_, new_n3655_, new_n3656_, new_n3657_, new_n3658_, new_n3659_,
    new_n3660_, new_n3661_, new_n3662_, new_n3663_, new_n3664_, new_n3665_,
    new_n3666_, new_n3667_, new_n3668_, new_n3669_, new_n3670_, new_n3671_,
    new_n3672_, new_n3673_, new_n3674_, new_n3675_, new_n3676_, new_n3677_,
    new_n3678_, new_n3679_, new_n3680_, new_n3681_, new_n3682_, new_n3683_,
    new_n3684_, new_n3685_, new_n3686_, new_n3687_, new_n3688_, new_n3689_,
    new_n3690_, new_n3691_, new_n3692_, new_n3693_, new_n3694_, new_n3695_,
    new_n3696_, new_n3697_, new_n3698_, new_n3699_, new_n3700_, new_n3701_,
    new_n3702_, new_n3703_, new_n3704_, new_n3705_, new_n3706_, new_n3707_,
    new_n3708_, new_n3709_, new_n3710_, new_n3711_, new_n3712_, new_n3713_,
    new_n3714_, new_n3715_, new_n3716_, new_n3717_, new_n3718_, new_n3719_,
    new_n3720_, new_n3721_, new_n3722_, new_n3723_, new_n3724_, new_n3725_,
    new_n3726_, new_n3727_, new_n3728_, new_n3729_, new_n3730_, new_n3731_,
    new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_, new_n3737_,
    new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_, new_n3743_,
    new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_, new_n3749_,
    new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_, new_n3755_,
    new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_, new_n3761_,
    new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_, new_n3767_,
    new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_, new_n3773_,
    new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_, new_n3779_,
    new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_, new_n3785_,
    new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_, new_n3791_,
    new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_, new_n3797_,
    new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_, new_n3803_,
    new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_, new_n3809_,
    new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_, new_n3815_,
    new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_, new_n3821_,
    new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_, new_n3827_,
    new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_, new_n3833_,
    new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_, new_n3839_,
    new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_, new_n3845_,
    new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_, new_n3851_,
    new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_, new_n3857_,
    new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_, new_n3863_,
    new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_, new_n3869_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_,
    new_n4158_, new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_,
    new_n4164_, new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_,
    new_n4170_, new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_,
    new_n4176_, new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_,
    new_n4182_, new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_,
    new_n4188_, new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_,
    new_n4194_, new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_,
    new_n4200_, new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_,
    new_n4206_, new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_,
    new_n4212_, new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_,
    new_n4218_, new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_,
    new_n4224_, new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_,
    new_n4230_, new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_,
    new_n4236_, new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_,
    new_n4242_, new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_,
    new_n4248_, new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_,
    new_n4254_, new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_,
    new_n4260_, new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_,
    new_n4266_, new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_,
    new_n4272_, new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_,
    new_n4278_, new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_,
    new_n4284_, new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_,
    new_n4290_, new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_,
    new_n4296_, new_n4297_, new_n4298_, new_n4299_, new_n4300_, new_n4301_,
    new_n4302_, new_n4303_, new_n4304_, new_n4305_, new_n4306_, new_n4307_,
    new_n4308_, new_n4309_, new_n4310_, new_n4311_, new_n4312_, new_n4313_,
    new_n4314_, new_n4315_, new_n4316_, new_n4317_, new_n4318_, new_n4319_,
    new_n4320_, new_n4321_, new_n4322_, new_n4323_, new_n4324_, new_n4325_,
    new_n4326_, new_n4327_, new_n4328_, new_n4329_, new_n4330_, new_n4331_,
    new_n4332_, new_n4333_, new_n4334_, new_n4335_, new_n4336_, new_n4337_,
    new_n4338_, new_n4339_, new_n4340_, new_n4341_, new_n4342_, new_n4343_,
    new_n4344_, new_n4345_, new_n4346_, new_n4347_, new_n4348_, new_n4349_,
    new_n4350_, new_n4351_, new_n4352_, new_n4353_, new_n4354_, new_n4355_,
    new_n4356_, new_n4357_, new_n4358_, new_n4359_, new_n4360_, new_n4361_,
    new_n4362_, new_n4363_, new_n4364_, new_n4365_, new_n4366_, new_n4367_,
    new_n4368_, new_n4369_, new_n4370_, new_n4371_, new_n4372_, new_n4373_,
    new_n4374_, new_n4375_, new_n4376_, new_n4377_, new_n4378_, new_n4379_,
    new_n4380_, new_n4381_, new_n4382_, new_n4383_, new_n4384_, new_n4385_,
    new_n4386_, new_n4387_, new_n4388_, new_n4389_, new_n4390_, new_n4391_,
    new_n4392_, new_n4393_, new_n4394_, new_n4395_, new_n4396_, new_n4397_,
    new_n4398_, new_n4399_, new_n4400_, new_n4401_, new_n4402_, new_n4403_,
    new_n4404_, new_n4405_, new_n4406_, new_n4407_, new_n4408_, new_n4409_,
    new_n4410_, new_n4411_, new_n4412_, new_n4413_, new_n4414_, new_n4415_,
    new_n4416_, new_n4417_, new_n4418_, new_n4419_, new_n4420_, new_n4421_,
    new_n4422_, new_n4423_, new_n4424_, new_n4425_, new_n4426_, new_n4427_,
    new_n4428_, new_n4429_, new_n4430_, new_n4431_, new_n4432_, new_n4433_,
    new_n4434_, new_n4435_, new_n4436_, new_n4437_, new_n4438_, new_n4439_,
    new_n4440_, new_n4441_, new_n4442_, new_n4443_, new_n4444_, new_n4445_,
    new_n4446_, new_n4447_, new_n4448_, new_n4449_, new_n4450_, new_n4451_,
    new_n4452_, new_n4453_, new_n4454_, new_n4455_, new_n4456_, new_n4457_,
    new_n4458_, new_n4459_, new_n4460_, new_n4461_, new_n4462_, new_n4463_,
    new_n4464_, new_n4465_, new_n4466_, new_n4467_, new_n4468_, new_n4469_,
    new_n4470_, new_n4471_, new_n4472_, new_n4473_, new_n4474_, new_n4475_,
    new_n4476_, new_n4477_, new_n4478_, new_n4479_, new_n4480_, new_n4481_,
    new_n4482_, new_n4483_, new_n4484_, new_n4485_, new_n4486_, new_n4487_,
    new_n4488_, new_n4489_, new_n4490_, new_n4491_, new_n4492_, new_n4493_,
    new_n4494_, new_n4495_, new_n4496_, new_n4497_, new_n4498_, new_n4499_,
    new_n4500_, new_n4501_, new_n4502_, new_n4503_, new_n4504_, new_n4505_,
    new_n4506_, new_n4507_, new_n4508_, new_n4509_, new_n4510_, new_n4511_,
    new_n4512_, new_n4513_, new_n4514_, new_n4515_, new_n4516_, new_n4517_,
    new_n4518_, new_n4519_, new_n4520_, new_n4521_, new_n4522_, new_n4523_,
    new_n4524_, new_n4525_, new_n4526_, new_n4527_, new_n4528_, new_n4529_,
    new_n4530_, new_n4531_, new_n4532_, new_n4533_, new_n4534_, new_n4535_,
    new_n4536_, new_n4537_, new_n4538_, new_n4539_, new_n4540_, new_n4541_,
    new_n4542_, new_n4543_, new_n4544_, new_n4545_, new_n4546_, new_n4547_,
    new_n4548_, new_n4549_, new_n4550_, new_n4551_, new_n4552_, new_n4553_,
    new_n4554_, new_n4555_, new_n4556_, new_n4557_, new_n4558_, new_n4559_,
    new_n4560_, new_n4561_, new_n4562_, new_n4563_, new_n4564_, new_n4565_,
    new_n4566_, new_n4567_, new_n4568_, new_n4569_, new_n4570_, new_n4571_,
    new_n4572_, new_n4573_, new_n4574_, new_n4575_, new_n4576_, new_n4577_,
    new_n4578_, new_n4579_, new_n4580_, new_n4581_, new_n4582_, new_n4583_,
    new_n4584_, new_n4585_, new_n4586_, new_n4587_, new_n4588_, new_n4589_,
    new_n4590_, new_n4591_, new_n4592_, new_n4593_, new_n4594_, new_n4595_,
    new_n4596_, new_n4597_, new_n4598_, new_n4599_, new_n4600_, new_n4601_,
    new_n4602_, new_n4603_, new_n4604_, new_n4605_, new_n4606_, new_n4607_,
    new_n4608_, new_n4609_, new_n4610_, new_n4611_, new_n4612_, new_n4613_,
    new_n4614_, new_n4615_, new_n4616_, new_n4617_, new_n4618_, new_n4619_,
    new_n4620_, new_n4621_, new_n4622_, new_n4623_, new_n4624_, new_n4625_,
    new_n4626_, new_n4627_, new_n4628_, new_n4629_, new_n4630_, new_n4631_,
    new_n4632_, new_n4633_, new_n4634_, new_n4635_, new_n4636_, new_n4637_,
    new_n4638_, new_n4639_, new_n4640_, new_n4641_, new_n4642_, new_n4643_,
    new_n4644_, new_n4645_, new_n4646_, new_n4647_, new_n4648_, new_n4649_,
    new_n4650_, new_n4651_, new_n4652_, new_n4653_, new_n4654_, new_n4655_,
    new_n4656_, new_n4657_, new_n4658_, new_n4659_, new_n4660_, new_n4661_,
    new_n4662_, new_n4663_, new_n4664_, new_n4665_, new_n4666_, new_n4667_,
    new_n4668_, new_n4669_, new_n4670_, new_n4671_, new_n4672_, new_n4673_,
    new_n4674_, new_n4675_, new_n4676_, new_n4677_, new_n4678_, new_n4679_,
    new_n4680_, new_n4681_, new_n4682_, new_n4683_, new_n4684_, new_n4685_,
    new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_, new_n4691_,
    new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_, new_n4697_,
    new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_, new_n4703_,
    new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_, new_n4709_,
    new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_, new_n4715_,
    new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_, new_n4721_,
    new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_, new_n4727_,
    new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_, new_n4733_,
    new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_, new_n4739_,
    new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_, new_n4745_,
    new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_, new_n4751_,
    new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_, new_n4757_,
    new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_, new_n4763_,
    new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_, new_n4769_,
    new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_, new_n4775_,
    new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_, new_n4781_,
    new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_, new_n4787_,
    new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_, new_n4793_,
    new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_, new_n4799_,
    new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_, new_n4805_,
    new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_, new_n4811_,
    new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_, new_n4817_,
    new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_, new_n4823_,
    new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_, new_n4829_,
    new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_, new_n4835_,
    new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_, new_n4841_,
    new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5045_,
    new_n5046_, new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_,
    new_n5052_, new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_,
    new_n5058_, new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_,
    new_n5064_, new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_,
    new_n5070_, new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_,
    new_n5076_, new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_,
    new_n5082_, new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_,
    new_n5088_, new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_,
    new_n5094_, new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_,
    new_n5100_, new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_,
    new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_,
    new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_,
    new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_,
    new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_,
    new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5309_,
    new_n5310_, new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_,
    new_n5316_, new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_,
    new_n5322_, new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_,
    new_n5328_, new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_,
    new_n5334_, new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_,
    new_n5340_, new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_,
    new_n5346_, new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_,
    new_n5352_, new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_,
    new_n5358_, new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_,
    new_n5364_, new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_,
    new_n5370_, new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_,
    new_n5376_, new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_,
    new_n5382_, new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_,
    new_n5388_, new_n5389_, new_n5390_, new_n5391_, new_n5392_, new_n5393_,
    new_n5394_, new_n5395_, new_n5396_, new_n5397_, new_n5398_, new_n5399_,
    new_n5400_, new_n5401_, new_n5402_, new_n5403_, new_n5404_, new_n5405_,
    new_n5406_, new_n5407_, new_n5408_, new_n5409_, new_n5410_, new_n5411_,
    new_n5412_, new_n5413_, new_n5414_, new_n5415_, new_n5416_, new_n5417_,
    new_n5418_, new_n5419_, new_n5420_, new_n5421_, new_n5422_, new_n5423_,
    new_n5424_, new_n5425_, new_n5426_, new_n5427_, new_n5428_, new_n5429_,
    new_n5430_, new_n5431_, new_n5432_, new_n5433_, new_n5434_, new_n5435_,
    new_n5436_, new_n5437_, new_n5438_, new_n5439_, new_n5440_, new_n5441_,
    new_n5442_, new_n5443_, new_n5444_, new_n5445_, new_n5446_, new_n5447_,
    new_n5448_, new_n5449_, new_n5450_, new_n5451_, new_n5452_, new_n5453_,
    new_n5454_, new_n5455_, new_n5456_, new_n5457_, new_n5458_, new_n5459_,
    new_n5460_, new_n5461_, new_n5462_, new_n5463_, new_n5464_, new_n5465_,
    new_n5466_, new_n5467_, new_n5468_, new_n5469_, new_n5470_, new_n5471_,
    new_n5472_, new_n5473_, new_n5474_, new_n5475_, new_n5476_, new_n5477_,
    new_n5478_, new_n5479_, new_n5480_, new_n5481_, new_n5482_, new_n5483_,
    new_n5484_, new_n5485_, new_n5486_, new_n5487_, new_n5488_, new_n5489_,
    new_n5490_, new_n5491_, new_n5492_, new_n5493_, new_n5494_, new_n5495_,
    new_n5496_, new_n5497_, new_n5498_, new_n5499_, new_n5500_, new_n5501_,
    new_n5502_, new_n5503_, new_n5504_, new_n5505_, new_n5506_, new_n5507_,
    new_n5508_, new_n5509_, new_n5510_, new_n5511_, new_n5512_, new_n5513_,
    new_n5514_, new_n5515_, new_n5516_, new_n5517_, new_n5518_, new_n5519_,
    new_n5520_, new_n5521_, new_n5522_, new_n5523_, new_n5524_, new_n5525_,
    new_n5526_, new_n5527_, new_n5528_, new_n5529_, new_n5530_, new_n5531_,
    new_n5532_, new_n5533_, new_n5534_, new_n5535_, new_n5536_, new_n5537_,
    new_n5538_, new_n5539_, new_n5540_, new_n5541_, new_n5542_, new_n5543_,
    new_n5544_, new_n5545_, new_n5546_, new_n5547_, new_n5548_, new_n5549_,
    new_n5550_, new_n5551_, new_n5552_, new_n5553_, new_n5554_, new_n5555_,
    new_n5556_, new_n5557_, new_n5558_, new_n5559_, new_n5560_, new_n5561_,
    new_n5562_, new_n5563_, new_n5564_, new_n5565_, new_n5566_, new_n5567_,
    new_n5568_, new_n5569_, new_n5570_, new_n5571_, new_n5572_, new_n5573_,
    new_n5574_, new_n5575_, new_n5576_, new_n5577_, new_n5578_, new_n5579_,
    new_n5580_, new_n5581_, new_n5582_, new_n5583_, new_n5584_, new_n5585_,
    new_n5586_, new_n5587_, new_n5588_, new_n5589_, new_n5590_, new_n5591_,
    new_n5592_, new_n5593_, new_n5594_, new_n5595_, new_n5596_, new_n5597_,
    new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_, new_n5603_,
    new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_, new_n5609_,
    new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_, new_n5615_,
    new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_, new_n5621_,
    new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_, new_n5627_,
    new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_, new_n5633_,
    new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_, new_n5639_,
    new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_, new_n5645_,
    new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_, new_n5651_,
    new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5656_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5716_, new_n5717_,
    new_n5718_, new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_,
    new_n5724_, new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_,
    new_n5730_, new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_,
    new_n5736_, new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_,
    new_n5742_, new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_,
    new_n5748_, new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_,
    new_n5754_, new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_,
    new_n5760_, new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_,
    new_n5766_, new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_,
    new_n5772_, new_n5773_, new_n5774_, new_n5775_, new_n5776_, new_n5777_,
    new_n5778_, new_n5779_, new_n5780_, new_n5781_, new_n5782_, new_n5783_,
    new_n5784_, new_n5785_, new_n5786_, new_n5787_, new_n5788_, new_n5789_,
    new_n5790_, new_n5791_, new_n5792_, new_n5793_, new_n5794_, new_n5795_,
    new_n5796_, new_n5797_, new_n5798_, new_n5799_, new_n5800_, new_n5801_,
    new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_, new_n5807_,
    new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_, new_n5813_,
    new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_, new_n5819_,
    new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_, new_n5825_,
    new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_, new_n5831_,
    new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_, new_n5837_,
    new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_, new_n5843_,
    new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_, new_n5849_,
    new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_, new_n5855_,
    new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_, new_n5861_,
    new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_, new_n5867_,
    new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_, new_n5873_,
    new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_, new_n5879_,
    new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_, new_n5885_,
    new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_, new_n5891_,
    new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_, new_n5897_,
    new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_, new_n5903_,
    new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_, new_n5909_,
    new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_, new_n5915_,
    new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_, new_n5921_,
    new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_, new_n5927_,
    new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_, new_n5933_,
    new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_, new_n5939_,
    new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_, new_n5945_,
    new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_, new_n5951_,
    new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_, new_n5957_,
    new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_, new_n5963_,
    new_n5964_, new_n5965_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_,
    new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6157_, new_n6158_, new_n6159_, new_n6160_, new_n6161_,
    new_n6162_, new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_,
    new_n6168_, new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_,
    new_n6174_, new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_,
    new_n6180_, new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_,
    new_n6186_, new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_,
    new_n6192_, new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_,
    new_n6198_, new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_,
    new_n6204_, new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_,
    new_n6210_, new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_,
    new_n6216_, new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_,
    new_n6222_, new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_,
    new_n6228_, new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_,
    new_n6234_, new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_,
    new_n6240_, new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_,
    new_n6246_, new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_,
    new_n6252_, new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_,
    new_n6258_, new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_,
    new_n6264_, new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_,
    new_n6270_, new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_,
    new_n6276_, new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_,
    new_n6282_, new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_,
    new_n6288_, new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_,
    new_n6294_, new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_,
    new_n6300_, new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_,
    new_n6306_, new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_,
    new_n6312_, new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_,
    new_n6318_, new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_,
    new_n6324_, new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_,
    new_n6330_, new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_,
    new_n6336_, new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_,
    new_n6342_, new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_,
    new_n6348_, new_n6349_, new_n6350_, new_n6351_, new_n6352_, new_n6353_,
    new_n6354_, new_n6355_, new_n6356_, new_n6357_, new_n6358_, new_n6359_,
    new_n6360_, new_n6361_, new_n6362_, new_n6363_, new_n6364_, new_n6365_,
    new_n6366_, new_n6367_, new_n6368_, new_n6369_, new_n6370_, new_n6371_,
    new_n6372_, new_n6373_, new_n6374_, new_n6375_, new_n6376_, new_n6377_,
    new_n6378_, new_n6379_, new_n6380_, new_n6381_, new_n6382_, new_n6383_,
    new_n6384_, new_n6385_, new_n6386_, new_n6387_, new_n6388_, new_n6389_,
    new_n6390_, new_n6391_, new_n6392_, new_n6393_, new_n6394_, new_n6395_,
    new_n6396_, new_n6397_, new_n6398_, new_n6399_, new_n6400_, new_n6401_,
    new_n6402_, new_n6403_, new_n6404_, new_n6405_, new_n6406_, new_n6407_,
    new_n6408_, new_n6409_, new_n6410_, new_n6411_, new_n6412_, new_n6413_,
    new_n6414_, new_n6415_, new_n6416_, new_n6417_, new_n6418_, new_n6419_,
    new_n6420_, new_n6421_, new_n6422_, new_n6423_, new_n6424_, new_n6425_,
    new_n6426_, new_n6427_, new_n6428_, new_n6429_, new_n6430_, new_n6431_,
    new_n6432_, new_n6433_, new_n6434_, new_n6435_, new_n6436_, new_n6437_,
    new_n6438_, new_n6439_, new_n6440_, new_n6441_, new_n6442_, new_n6443_,
    new_n6444_, new_n6445_, new_n6446_, new_n6447_, new_n6448_, new_n6449_,
    new_n6450_, new_n6451_, new_n6452_, new_n6453_, new_n6454_, new_n6455_,
    new_n6456_, new_n6457_, new_n6458_, new_n6459_, new_n6460_, new_n6461_,
    new_n6462_, new_n6463_, new_n6464_, new_n6465_, new_n6466_, new_n6467_,
    new_n6468_, new_n6469_, new_n6470_, new_n6471_, new_n6472_, new_n6473_,
    new_n6474_, new_n6475_, new_n6476_, new_n6477_, new_n6478_, new_n6479_,
    new_n6480_, new_n6481_, new_n6482_, new_n6483_, new_n6484_, new_n6485_,
    new_n6486_, new_n6487_, new_n6488_, new_n6489_, new_n6490_, new_n6491_,
    new_n6492_, new_n6493_, new_n6494_, new_n6495_, new_n6496_, new_n6497_,
    new_n6498_, new_n6499_, new_n6500_, new_n6501_, new_n6502_, new_n6503_,
    new_n6504_, new_n6505_, new_n6506_, new_n6507_, new_n6508_, new_n6509_,
    new_n6510_, new_n6511_, new_n6512_, new_n6513_, new_n6514_, new_n6515_,
    new_n6516_, new_n6517_, new_n6518_, new_n6519_, new_n6520_, new_n6521_,
    new_n6522_, new_n6523_, new_n6524_, new_n6525_, new_n6526_, new_n6527_,
    new_n6528_, new_n6529_, new_n6530_, new_n6531_, new_n6532_, new_n6533_,
    new_n6534_, new_n6535_, new_n6536_, new_n6537_, new_n6538_, new_n6539_,
    new_n6540_, new_n6541_, new_n6542_, new_n6543_, new_n6544_, new_n6545_,
    new_n6546_, new_n6547_, new_n6548_, new_n6549_, new_n6550_, new_n6551_,
    new_n6552_, new_n6553_, new_n6554_, new_n6555_, new_n6556_, new_n6557_,
    new_n6558_, new_n6559_, new_n6560_, new_n6561_, new_n6562_, new_n6563_,
    new_n6564_, new_n6565_, new_n6566_, new_n6567_, new_n6568_, new_n6569_,
    new_n6570_, new_n6571_, new_n6572_, new_n6573_, new_n6574_, new_n6575_,
    new_n6576_, new_n6577_, new_n6578_, new_n6579_, new_n6580_, new_n6581_,
    new_n6582_, new_n6583_, new_n6584_, new_n6585_, new_n6586_, new_n6587_,
    new_n6588_, new_n6589_, new_n6590_, new_n6591_, new_n6592_, new_n6593_,
    new_n6594_, new_n6595_, new_n6596_, new_n6597_, new_n6598_, new_n6599_,
    new_n6600_, new_n6601_, new_n6602_, new_n6603_, new_n6604_, new_n6605_,
    new_n6606_, new_n6607_, new_n6608_, new_n6609_, new_n6610_, new_n6611_,
    new_n6612_, new_n6613_, new_n6614_, new_n6615_, new_n6616_, new_n6617_,
    new_n6618_, new_n6619_, new_n6620_, new_n6621_, new_n6622_, new_n6623_,
    new_n6624_, new_n6625_, new_n6626_, new_n6627_, new_n6628_, new_n6629_,
    new_n6630_, new_n6631_, new_n6632_, new_n6633_, new_n6634_, new_n6635_,
    new_n6636_, new_n6637_, new_n6638_, new_n6639_, new_n6640_, new_n6641_,
    new_n6642_, new_n6643_, new_n6644_, new_n6645_, new_n6646_, new_n6647_,
    new_n6648_, new_n6649_, new_n6650_, new_n6651_, new_n6652_, new_n6653_,
    new_n6654_, new_n6655_, new_n6656_, new_n6657_, new_n6658_, new_n6659_,
    new_n6660_, new_n6661_, new_n6662_, new_n6663_, new_n6664_, new_n6665_,
    new_n6666_, new_n6667_, new_n6668_, new_n6669_, new_n6670_, new_n6671_,
    new_n6672_, new_n6673_, new_n6674_, new_n6675_, new_n6676_, new_n6677_,
    new_n6678_, new_n6679_, new_n6680_, new_n6681_, new_n6682_, new_n6683_,
    new_n6684_, new_n6685_, new_n6686_, new_n6687_, new_n6688_, new_n6689_,
    new_n6690_, new_n6691_, new_n6692_, new_n6693_, new_n6694_, new_n6695_,
    new_n6696_, new_n6697_, new_n6698_, new_n6699_, new_n6700_, new_n6701_,
    new_n6702_, new_n6703_, new_n6704_, new_n6705_, new_n6706_, new_n6707_,
    new_n6708_, new_n6709_, new_n6710_, new_n6711_, new_n6712_, new_n6713_,
    new_n6714_, new_n6715_, new_n6716_, new_n6717_, new_n6718_, new_n6719_,
    new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6724_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6771_, new_n6772_, new_n6773_,
    new_n6774_, new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_,
    new_n6780_, new_n6781_, new_n6782_, new_n6783_, new_n6784_, new_n6785_,
    new_n6786_, new_n6787_, new_n6788_, new_n6789_, new_n6790_, new_n6791_,
    new_n6792_, new_n6793_, new_n6794_, new_n6795_, new_n6796_, new_n6797_,
    new_n6798_, new_n6799_, new_n6800_, new_n6801_, new_n6802_, new_n6803_,
    new_n6804_, new_n6805_, new_n6806_, new_n6807_, new_n6808_, new_n6809_,
    new_n6810_, new_n6811_, new_n6812_, new_n6813_, new_n6814_, new_n6815_,
    new_n6816_, new_n6817_, new_n6818_, new_n6819_, new_n6820_, new_n6821_,
    new_n6822_, new_n6823_, new_n6824_, new_n6825_, new_n6826_, new_n6827_,
    new_n6828_, new_n6829_, new_n6830_, new_n6831_, new_n6832_, new_n6833_,
    new_n6834_, new_n6835_, new_n6836_, new_n6837_, new_n6838_, new_n6839_,
    new_n6840_, new_n6841_, new_n6842_, new_n6843_, new_n6844_, new_n6845_,
    new_n6846_, new_n6847_, new_n6848_, new_n6849_, new_n6850_, new_n6851_,
    new_n6852_, new_n6853_, new_n6854_, new_n6855_, new_n6856_, new_n6857_,
    new_n6858_, new_n6859_, new_n6860_, new_n6861_, new_n6862_, new_n6863_,
    new_n6864_, new_n6865_, new_n6866_, new_n6867_, new_n6868_, new_n6869_,
    new_n6870_, new_n6871_, new_n6872_, new_n6873_, new_n6874_, new_n6875_,
    new_n6876_, new_n6877_, new_n6878_, new_n6879_, new_n6880_, new_n6881_,
    new_n6882_, new_n6883_, new_n6884_, new_n6885_, new_n6886_, new_n6887_,
    new_n6888_, new_n6889_, new_n6890_, new_n6891_, new_n6892_, new_n6893_,
    new_n6894_, new_n6895_, new_n6896_, new_n6897_, new_n6898_, new_n6899_,
    new_n6900_, new_n6901_, new_n6902_, new_n6903_, new_n6904_, new_n6905_,
    new_n6906_, new_n6907_, new_n6908_, new_n6909_, new_n6910_, new_n6911_,
    new_n6912_, new_n6913_, new_n6914_, new_n6915_, new_n6916_, new_n6917_,
    new_n6918_, new_n6919_, new_n6920_, new_n6921_, new_n6922_, new_n6923_,
    new_n6924_, new_n6925_, new_n6926_, new_n6927_, new_n6928_, new_n6929_,
    new_n6930_, new_n6931_, new_n6932_, new_n6933_, new_n6934_, new_n6935_,
    new_n6936_, new_n6937_, new_n6938_, new_n6939_, new_n6940_, new_n6941_,
    new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_, new_n6947_,
    new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_, new_n6953_,
    new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_, new_n6959_,
    new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_, new_n6965_,
    new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_, new_n6971_,
    new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_, new_n6977_,
    new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_, new_n6983_,
    new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_, new_n6989_,
    new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_, new_n6995_,
    new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_, new_n7001_,
    new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_, new_n7007_,
    new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_, new_n7013_,
    new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_, new_n7019_,
    new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_, new_n7025_,
    new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_, new_n7031_,
    new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_, new_n7037_,
    new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_, new_n7043_,
    new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_, new_n7049_,
    new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_, new_n7055_,
    new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_, new_n7061_,
    new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_, new_n7067_,
    new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_, new_n7073_,
    new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_, new_n7079_,
    new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_, new_n7085_,
    new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_, new_n7091_,
    new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_, new_n7097_,
    new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_, new_n7103_,
    new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_, new_n7109_,
    new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_, new_n7115_,
    new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_, new_n7121_,
    new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_, new_n7127_,
    new_n7128_, new_n7129_, new_n7130_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_,
    new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_,
    new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_,
    new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_,
    new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_,
    new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_,
    new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_,
    new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_,
    new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_,
    new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_,
    new_n7350_, new_n7351_, new_n7352_, new_n7353_, new_n7354_, new_n7355_,
    new_n7356_, new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_,
    new_n7362_, new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_,
    new_n7368_, new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_,
    new_n7374_, new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_,
    new_n7380_, new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_,
    new_n7386_, new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_,
    new_n7392_, new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_,
    new_n7398_, new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_,
    new_n7404_, new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_,
    new_n7410_, new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_,
    new_n7416_, new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_,
    new_n7422_, new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_,
    new_n7428_, new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_,
    new_n7434_, new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_,
    new_n7440_, new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_,
    new_n7446_, new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_,
    new_n7452_, new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_,
    new_n7458_, new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_,
    new_n7464_, new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_,
    new_n7470_, new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_,
    new_n7476_, new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_,
    new_n7482_, new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_,
    new_n7488_, new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_,
    new_n7494_, new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_,
    new_n7500_, new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_,
    new_n7506_, new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_,
    new_n7512_, new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_,
    new_n7518_, new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_,
    new_n7524_, new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_,
    new_n7530_, new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_,
    new_n7536_, new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_,
    new_n7542_, new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_,
    new_n7548_, new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_,
    new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_,
    new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_,
    new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_, new_n7571_,
    new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_, new_n7577_,
    new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_, new_n7583_,
    new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_, new_n7589_,
    new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_, new_n7595_,
    new_n7596_, new_n7597_, new_n7598_, new_n7599_, new_n7600_, new_n7601_,
    new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_,
    new_n7608_, new_n7609_, new_n7610_, new_n7611_, new_n7612_, new_n7613_,
    new_n7614_, new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_,
    new_n7620_, new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_,
    new_n7626_, new_n7627_, new_n7628_, new_n7629_, new_n7630_, new_n7631_,
    new_n7632_, new_n7633_, new_n7634_, new_n7635_, new_n7636_, new_n7637_,
    new_n7638_, new_n7639_, new_n7640_, new_n7641_, new_n7642_, new_n7643_,
    new_n7644_, new_n7645_, new_n7646_, new_n7647_, new_n7648_, new_n7649_,
    new_n7650_, new_n7651_, new_n7652_, new_n7653_, new_n7654_, new_n7655_,
    new_n7656_, new_n7657_, new_n7658_, new_n7659_, new_n7660_, new_n7661_,
    new_n7662_, new_n7663_, new_n7664_, new_n7665_, new_n7666_, new_n7667_,
    new_n7668_, new_n7669_, new_n7670_, new_n7671_, new_n7672_, new_n7673_,
    new_n7674_, new_n7675_, new_n7676_, new_n7677_, new_n7678_, new_n7679_,
    new_n7680_, new_n7681_, new_n7682_, new_n7683_, new_n7684_, new_n7685_,
    new_n7686_, new_n7687_, new_n7688_, new_n7689_, new_n7690_, new_n7691_,
    new_n7692_, new_n7693_, new_n7694_, new_n7695_, new_n7696_, new_n7697_,
    new_n7698_, new_n7699_, new_n7700_, new_n7701_, new_n7702_, new_n7703_,
    new_n7704_, new_n7705_, new_n7706_, new_n7707_, new_n7708_, new_n7709_,
    new_n7710_, new_n7711_, new_n7712_, new_n7713_, new_n7714_, new_n7715_,
    new_n7716_, new_n7717_, new_n7718_, new_n7719_, new_n7720_, new_n7721_,
    new_n7722_, new_n7723_, new_n7724_, new_n7725_, new_n7726_, new_n7727_,
    new_n7728_, new_n7729_, new_n7730_, new_n7731_, new_n7732_, new_n7733_,
    new_n7734_, new_n7735_, new_n7736_, new_n7737_, new_n7738_, new_n7739_,
    new_n7740_, new_n7741_, new_n7742_, new_n7743_, new_n7744_, new_n7745_,
    new_n7746_, new_n7747_, new_n7748_, new_n7749_, new_n7750_, new_n7751_,
    new_n7752_, new_n7753_, new_n7754_, new_n7755_, new_n7756_, new_n7757_,
    new_n7758_, new_n7759_, new_n7760_, new_n7761_, new_n7762_, new_n7763_,
    new_n7764_, new_n7765_, new_n7766_, new_n7767_, new_n7768_, new_n7769_,
    new_n7770_, new_n7771_, new_n7772_, new_n7773_, new_n7774_, new_n7775_,
    new_n7776_, new_n7777_, new_n7778_, new_n7779_, new_n7780_, new_n7781_,
    new_n7782_, new_n7783_, new_n7784_, new_n7785_, new_n7786_, new_n7787_,
    new_n7788_, new_n7789_, new_n7790_, new_n7791_, new_n7792_, new_n7793_,
    new_n7794_, new_n7795_, new_n7796_, new_n7797_, new_n7798_, new_n7799_,
    new_n7800_, new_n7801_, new_n7802_, new_n7803_, new_n7804_, new_n7805_,
    new_n7806_, new_n7807_, new_n7808_, new_n7809_, new_n7810_, new_n7811_,
    new_n7812_, new_n7813_, new_n7814_, new_n7815_, new_n7816_, new_n7817_,
    new_n7818_, new_n7819_, new_n7820_, new_n7821_, new_n7822_, new_n7823_,
    new_n7824_, new_n7825_, new_n7826_, new_n7827_, new_n7828_, new_n7829_,
    new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_, new_n7835_,
    new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_, new_n7841_,
    new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_, new_n7847_,
    new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_, new_n7853_,
    new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_, new_n7859_,
    new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_, new_n7865_,
    new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_, new_n7871_,
    new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_, new_n7877_,
    new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_, new_n7883_,
    new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_, new_n7889_,
    new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_, new_n7895_,
    new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_, new_n7901_,
    new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_, new_n7907_,
    new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_, new_n7913_,
    new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_, new_n7919_,
    new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_, new_n7925_,
    new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_, new_n7931_,
    new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_, new_n7937_,
    new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_, new_n7943_,
    new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_, new_n7949_,
    new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_, new_n7955_,
    new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_, new_n7961_,
    new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_, new_n7967_,
    new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_, new_n7973_,
    new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_, new_n7979_,
    new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_, new_n7985_,
    new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_, new_n7991_,
    new_n7992_, new_n7993_, new_n7994_, new_n7995_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8115_, new_n8116_, new_n8117_,
    new_n8118_, new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_,
    new_n8124_, new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_,
    new_n8130_, new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_,
    new_n8136_, new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_,
    new_n8142_, new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_,
    new_n8148_, new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_,
    new_n8154_, new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_,
    new_n8160_, new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_,
    new_n8166_, new_n8167_, new_n8168_, new_n8169_, new_n8170_, new_n8171_,
    new_n8172_, new_n8173_, new_n8174_, new_n8175_, new_n8176_, new_n8177_,
    new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_, new_n8183_,
    new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_, new_n8189_,
    new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_, new_n8195_,
    new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_, new_n8201_,
    new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_, new_n8207_,
    new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_, new_n8213_,
    new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_,
    new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_,
    new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_, new_n8243_,
    new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_, new_n8249_,
    new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_, new_n8255_,
    new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_, new_n8261_,
    new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_, new_n8267_,
    new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_, new_n8273_,
    new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_, new_n8279_,
    new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_, new_n8285_,
    new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_, new_n8291_,
    new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_, new_n8297_,
    new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_, new_n8303_,
    new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_, new_n8309_,
    new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_, new_n8315_,
    new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_, new_n8321_,
    new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_, new_n8327_,
    new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_, new_n8333_,
    new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_, new_n8339_,
    new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_, new_n8345_,
    new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_, new_n8351_,
    new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_, new_n8357_,
    new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_, new_n8363_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8571_, new_n8572_, new_n8573_,
    new_n8574_, new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_,
    new_n8580_, new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_,
    new_n8586_, new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_,
    new_n8592_, new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_,
    new_n8598_, new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_,
    new_n8604_, new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_,
    new_n8610_, new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_,
    new_n8616_, new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_,
    new_n8622_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8942_, new_n8943_, new_n8944_, new_n8945_,
    new_n8946_, new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_,
    new_n8952_, new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_,
    new_n8958_, new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_,
    new_n8964_, new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_,
    new_n8970_, new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_,
    new_n8976_, new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_,
    new_n8982_, new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_,
    new_n8988_, new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_,
    new_n8994_, new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_,
    new_n9000_, new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_,
    new_n9006_, new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_,
    new_n9012_, new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_,
    new_n9018_, new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_,
    new_n9024_, new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_,
    new_n9030_, new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_,
    new_n9036_, new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_,
    new_n9042_, new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_,
    new_n9048_, new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_,
    new_n9054_, new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_,
    new_n9060_, new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_,
    new_n9066_, new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_,
    new_n9072_, new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_,
    new_n9078_, new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_,
    new_n9084_, new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_,
    new_n9090_, new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_,
    new_n9096_, new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_,
    new_n9102_, new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_,
    new_n9108_, new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_,
    new_n9114_, new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_,
    new_n9120_, new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_,
    new_n9126_, new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_,
    new_n9132_, new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_,
    new_n9138_, new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_,
    new_n9144_, new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_,
    new_n9150_, new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_,
    new_n9156_, new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_,
    new_n9162_, new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_,
    new_n9168_, new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_,
    new_n9174_, new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_,
    new_n9180_, new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_,
    new_n9186_, new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_,
    new_n9192_, new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_,
    new_n9198_, new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_,
    new_n9204_, new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_,
    new_n9210_, new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_,
    new_n9216_, new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_,
    new_n9222_, new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_,
    new_n9228_, new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_,
    new_n9234_, new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_,
    new_n9240_, new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_,
    new_n9246_, new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_,
    new_n9252_, new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_,
    new_n9258_, new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_,
    new_n9264_, new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_,
    new_n9270_, new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_,
    new_n9276_, new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_,
    new_n9282_, new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_,
    new_n9288_, new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_,
    new_n9294_, new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_,
    new_n9300_, new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_,
    new_n9306_, new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_,
    new_n9312_, new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_,
    new_n9318_, new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_,
    new_n9324_, new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_,
    new_n9330_, new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_,
    new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_,
    new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_,
    new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_,
    new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_,
    new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_,
    new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_,
    new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_,
    new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_,
    new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_,
    new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_,
    new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_,
    new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_,
    new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_,
    new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_,
    new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9425_,
    new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_, new_n9431_,
    new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_, new_n9437_,
    new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_, new_n9443_,
    new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_, new_n9449_,
    new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9455_,
    new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_, new_n9461_,
    new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_, new_n9467_,
    new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_, new_n9473_,
    new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_, new_n9479_,
    new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_, new_n9491_,
    new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9497_,
    new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_, new_n9503_,
    new_n9504_, new_n9505_, new_n9506_, new_n9507_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_,
    new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_,
    new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_,
    new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_,
    new_n9684_, new_n9685_, new_n9686_, new_n9687_, new_n9688_, new_n9689_,
    new_n9690_, new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_,
    new_n9696_, new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9702_, new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_,
    new_n9708_, new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_,
    new_n9714_, new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_,
    new_n9720_, new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_,
    new_n9726_, new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_,
    new_n9732_, new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_,
    new_n9738_, new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_,
    new_n9744_, new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_,
    new_n9750_, new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_,
    new_n9756_, new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_,
    new_n9762_, new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_,
    new_n9768_, new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_,
    new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_,
    new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_,
    new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_,
    new_n9792_, new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_,
    new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_,
    new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_,
    new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_,
    new_n9828_, new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_,
    new_n9834_, new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_,
    new_n9840_, new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_,
    new_n9846_, new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_,
    new_n9852_, new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_,
    new_n9858_, new_n9859_, new_n9860_, new_n9861_, new_n9862_, new_n9863_,
    new_n9864_, new_n9865_, new_n9866_, new_n9867_, new_n9868_, new_n9869_,
    new_n9870_, new_n9871_, new_n9872_, new_n9873_, new_n9874_, new_n9875_,
    new_n9876_, new_n9877_, new_n9878_, new_n9879_, new_n9880_, new_n9881_,
    new_n9882_, new_n9883_, new_n9884_, new_n9885_, new_n9886_, new_n9887_,
    new_n9888_, new_n9889_, new_n9890_, new_n9891_, new_n9892_, new_n9893_,
    new_n9894_, new_n9895_, new_n9896_, new_n9897_, new_n9898_, new_n9899_,
    new_n9900_, new_n9901_, new_n9902_, new_n9903_, new_n9904_, new_n9905_,
    new_n9906_, new_n9907_, new_n9908_, new_n9909_, new_n9910_, new_n9911_,
    new_n9912_, new_n9913_, new_n9914_, new_n9915_, new_n9916_, new_n9917_,
    new_n9918_, new_n9919_, new_n9920_, new_n9921_, new_n9922_, new_n9923_,
    new_n9924_, new_n9925_, new_n9926_, new_n9927_, new_n9928_, new_n9929_,
    new_n9930_, new_n9931_, new_n9932_, new_n9933_, new_n9934_, new_n9935_,
    new_n9936_, new_n9937_, new_n9938_, new_n9939_, new_n9940_, new_n9941_,
    new_n9942_, new_n9943_, new_n9944_, new_n9945_, new_n9946_, new_n9947_,
    new_n9948_, new_n9949_, new_n9950_, new_n9951_, new_n9952_, new_n9953_,
    new_n9954_, new_n9955_, new_n9956_, new_n9957_, new_n9958_, new_n9959_,
    new_n9960_, new_n9961_, new_n9962_, new_n9963_, new_n9964_, new_n9965_,
    new_n9966_, new_n9967_, new_n9968_, new_n9969_, new_n9970_, new_n9971_,
    new_n9972_, new_n9973_, new_n9974_, new_n9975_, new_n9976_, new_n9977_,
    new_n9978_, new_n9979_, new_n9980_, new_n9981_, new_n9982_, new_n9983_,
    new_n9984_, new_n9985_, new_n9986_, new_n9987_, new_n9988_, new_n9989_,
    new_n9990_, new_n9991_, new_n9992_, new_n9993_, new_n9994_, new_n9995_,
    new_n9996_, new_n9997_, new_n9998_, new_n9999_, new_n10000_,
    new_n10001_, new_n10002_, new_n10003_, new_n10004_, new_n10005_,
    new_n10006_, new_n10007_, new_n10008_, new_n10009_, new_n10010_,
    new_n10011_, new_n10012_, new_n10013_, new_n10014_, new_n10015_,
    new_n10016_, new_n10017_, new_n10018_, new_n10019_, new_n10020_,
    new_n10021_, new_n10022_, new_n10023_, new_n10024_, new_n10025_,
    new_n10026_, new_n10027_, new_n10028_, new_n10029_, new_n10030_,
    new_n10031_, new_n10032_, new_n10033_, new_n10034_, new_n10035_,
    new_n10036_, new_n10037_, new_n10038_, new_n10039_, new_n10040_,
    new_n10041_, new_n10042_, new_n10043_, new_n10044_, new_n10045_,
    new_n10046_, new_n10047_, new_n10048_, new_n10049_, new_n10050_,
    new_n10051_, new_n10052_, new_n10053_, new_n10054_, new_n10055_,
    new_n10056_, new_n10057_, new_n10058_, new_n10059_, new_n10060_,
    new_n10061_, new_n10062_, new_n10063_, new_n10064_, new_n10065_,
    new_n10066_, new_n10067_, new_n10068_, new_n10069_, new_n10070_,
    new_n10071_, new_n10072_, new_n10073_, new_n10074_, new_n10075_,
    new_n10076_, new_n10077_, new_n10078_, new_n10079_, new_n10080_,
    new_n10081_, new_n10082_, new_n10083_, new_n10084_, new_n10085_,
    new_n10086_, new_n10087_, new_n10088_, new_n10089_, new_n10090_,
    new_n10091_, new_n10092_, new_n10093_, new_n10094_, new_n10095_,
    new_n10096_, new_n10097_, new_n10098_, new_n10099_, new_n10100_,
    new_n10101_, new_n10102_, new_n10103_, new_n10104_, new_n10105_,
    new_n10106_, new_n10107_, new_n10108_, new_n10109_, new_n10110_,
    new_n10111_, new_n10112_, new_n10113_, new_n10114_, new_n10115_,
    new_n10116_, new_n10117_, new_n10118_, new_n10119_, new_n10120_,
    new_n10121_, new_n10122_, new_n10123_, new_n10124_, new_n10125_,
    new_n10126_, new_n10127_, new_n10128_, new_n10129_, new_n10130_,
    new_n10131_, new_n10132_, new_n10133_, new_n10134_, new_n10135_,
    new_n10136_, new_n10137_, new_n10138_, new_n10139_, new_n10140_,
    new_n10141_, new_n10142_, new_n10143_, new_n10144_, new_n10145_,
    new_n10146_, new_n10147_, new_n10148_, new_n10149_, new_n10150_,
    new_n10151_, new_n10152_, new_n10153_, new_n10154_, new_n10155_,
    new_n10156_, new_n10157_, new_n10158_, new_n10159_, new_n10160_,
    new_n10161_, new_n10162_, new_n10163_, new_n10164_, new_n10165_,
    new_n10166_, new_n10167_, new_n10168_, new_n10169_, new_n10170_,
    new_n10171_, new_n10172_, new_n10173_, new_n10174_, new_n10175_,
    new_n10176_, new_n10177_, new_n10178_, new_n10179_, new_n10180_,
    new_n10181_, new_n10182_, new_n10183_, new_n10184_, new_n10185_,
    new_n10186_, new_n10187_, new_n10188_, new_n10189_, new_n10190_,
    new_n10191_, new_n10192_, new_n10193_, new_n10194_, new_n10195_,
    new_n10196_, new_n10197_, new_n10198_, new_n10199_, new_n10200_,
    new_n10201_, new_n10202_, new_n10203_, new_n10204_, new_n10205_,
    new_n10206_, new_n10207_, new_n10208_, new_n10209_, new_n10210_,
    new_n10211_, new_n10212_, new_n10213_, new_n10214_, new_n10215_,
    new_n10216_, new_n10217_, new_n10218_, new_n10219_, new_n10220_,
    new_n10221_, new_n10222_, new_n10223_, new_n10224_, new_n10225_,
    new_n10226_, new_n10227_, new_n10228_, new_n10229_, new_n10230_,
    new_n10231_, new_n10232_, new_n10233_, new_n10234_, new_n10235_,
    new_n10236_, new_n10237_, new_n10238_, new_n10239_, new_n10240_,
    new_n10241_, new_n10242_, new_n10243_, new_n10244_, new_n10245_,
    new_n10246_, new_n10247_, new_n10248_, new_n10249_, new_n10250_,
    new_n10251_, new_n10252_, new_n10253_, new_n10254_, new_n10255_,
    new_n10256_, new_n10257_, new_n10258_, new_n10259_, new_n10260_,
    new_n10261_, new_n10262_, new_n10263_, new_n10264_, new_n10265_,
    new_n10266_, new_n10267_, new_n10268_, new_n10269_, new_n10270_,
    new_n10271_, new_n10272_, new_n10273_, new_n10274_, new_n10275_,
    new_n10276_, new_n10277_, new_n10278_, new_n10279_, new_n10280_,
    new_n10281_, new_n10282_, new_n10283_, new_n10284_, new_n10285_,
    new_n10286_, new_n10287_, new_n10288_, new_n10289_, new_n10290_,
    new_n10291_, new_n10292_, new_n10293_, new_n10294_, new_n10295_,
    new_n10296_, new_n10297_, new_n10298_, new_n10299_, new_n10300_,
    new_n10301_, new_n10302_, new_n10303_, new_n10304_, new_n10305_,
    new_n10306_, new_n10307_, new_n10308_, new_n10309_, new_n10310_,
    new_n10311_, new_n10312_, new_n10313_, new_n10314_, new_n10315_,
    new_n10316_, new_n10317_, new_n10318_, new_n10319_, new_n10320_,
    new_n10321_, new_n10322_, new_n10323_, new_n10324_, new_n10325_,
    new_n10326_, new_n10327_, new_n10328_, new_n10329_, new_n10330_,
    new_n10331_, new_n10332_, new_n10333_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10618_, new_n10619_, new_n10620_,
    new_n10621_, new_n10622_, new_n10623_, new_n10624_, new_n10625_,
    new_n10626_, new_n10627_, new_n10628_, new_n10629_, new_n10630_,
    new_n10631_, new_n10632_, new_n10633_, new_n10634_, new_n10635_,
    new_n10636_, new_n10637_, new_n10638_, new_n10639_, new_n10640_,
    new_n10641_, new_n10642_, new_n10643_, new_n10644_, new_n10645_,
    new_n10646_, new_n10647_, new_n10648_, new_n10649_, new_n10650_,
    new_n10651_, new_n10652_, new_n10653_, new_n10654_, new_n10655_,
    new_n10656_, new_n10657_, new_n10658_, new_n10659_, new_n10660_,
    new_n10661_, new_n10662_, new_n10663_, new_n10664_, new_n10665_,
    new_n10666_, new_n10667_, new_n10668_, new_n10669_, new_n10670_,
    new_n10671_, new_n10672_, new_n10673_, new_n10674_, new_n10675_,
    new_n10676_, new_n10677_, new_n10678_, new_n10679_, new_n10680_,
    new_n10681_, new_n10682_, new_n10683_, new_n10684_, new_n10685_,
    new_n10686_, new_n10687_, new_n10688_, new_n10689_, new_n10690_,
    new_n10691_, new_n10692_, new_n10693_, new_n10694_, new_n10695_,
    new_n10696_, new_n10697_, new_n10698_, new_n10699_, new_n10700_,
    new_n10701_, new_n10702_, new_n10703_, new_n10704_, new_n10705_,
    new_n10706_, new_n10707_, new_n10708_, new_n10709_, new_n10710_,
    new_n10711_, new_n10712_, new_n10713_, new_n10714_, new_n10715_,
    new_n10716_, new_n10717_, new_n10718_, new_n10719_, new_n10720_,
    new_n10721_, new_n10722_, new_n10723_, new_n10724_, new_n10725_,
    new_n10726_, new_n10727_, new_n10728_, new_n10729_, new_n10730_,
    new_n10731_, new_n10732_, new_n10733_, new_n10734_, new_n10735_,
    new_n10736_, new_n10737_, new_n10738_, new_n10739_, new_n10740_,
    new_n10741_, new_n10742_, new_n10743_, new_n10744_, new_n10745_,
    new_n10746_, new_n10747_, new_n10748_, new_n10749_, new_n10750_,
    new_n10751_, new_n10752_, new_n10753_, new_n10754_, new_n10755_,
    new_n10756_, new_n10757_, new_n10758_, new_n10759_, new_n10760_,
    new_n10761_, new_n10762_, new_n10763_, new_n10764_, new_n10765_,
    new_n10766_, new_n10767_, new_n10768_, new_n10769_, new_n10770_,
    new_n10771_, new_n10772_, new_n10773_, new_n10774_, new_n10775_,
    new_n10776_, new_n10777_, new_n10778_, new_n10779_, new_n10780_,
    new_n10781_, new_n10782_, new_n10783_, new_n10784_, new_n10785_,
    new_n10786_, new_n10787_, new_n10788_, new_n10789_, new_n10790_,
    new_n10791_, new_n10792_, new_n10793_, new_n10794_, new_n10795_,
    new_n10796_, new_n10797_, new_n10798_, new_n10799_, new_n10800_,
    new_n10801_, new_n10802_, new_n10803_, new_n10804_, new_n10805_,
    new_n10806_, new_n10807_, new_n10808_, new_n10809_, new_n10810_,
    new_n10811_, new_n10812_, new_n10813_, new_n10814_, new_n10815_,
    new_n10816_, new_n10817_, new_n10818_, new_n10819_, new_n10820_,
    new_n10821_, new_n10822_, new_n10823_, new_n10824_, new_n10825_,
    new_n10826_, new_n10827_, new_n10828_, new_n10829_, new_n10830_,
    new_n10831_, new_n10832_, new_n10833_, new_n10834_, new_n10835_,
    new_n10836_, new_n10837_, new_n10838_, new_n10839_, new_n10840_,
    new_n10841_, new_n10842_, new_n10843_, new_n10844_, new_n10845_,
    new_n10846_, new_n10847_, new_n10848_, new_n10849_, new_n10850_,
    new_n10851_, new_n10852_, new_n10853_, new_n10854_, new_n10855_,
    new_n10856_, new_n10857_, new_n10858_, new_n10859_, new_n10860_,
    new_n10861_, new_n10862_, new_n10863_, new_n10864_, new_n10865_,
    new_n10866_, new_n10867_, new_n10868_, new_n10869_, new_n10870_,
    new_n10871_, new_n10872_, new_n10873_, new_n10874_, new_n10875_,
    new_n10876_, new_n10877_, new_n10878_, new_n10879_, new_n10880_,
    new_n10881_, new_n10882_, new_n10883_, new_n10884_, new_n10885_,
    new_n10886_, new_n10887_, new_n10888_, new_n10889_, new_n10890_,
    new_n10891_, new_n10892_, new_n10893_, new_n10894_, new_n10895_,
    new_n10896_, new_n10897_, new_n10898_, new_n10899_, new_n10900_,
    new_n10901_, new_n10902_, new_n10903_, new_n10904_, new_n10905_,
    new_n10906_, new_n10907_, new_n10908_, new_n10909_, new_n10910_,
    new_n10911_, new_n10912_, new_n10913_, new_n10914_, new_n10915_,
    new_n10916_, new_n10917_, new_n10918_, new_n10919_, new_n10920_,
    new_n10921_, new_n10922_, new_n10923_, new_n10924_, new_n10925_,
    new_n10926_, new_n10927_, new_n10928_, new_n10929_, new_n10930_,
    new_n10931_, new_n10932_, new_n10933_, new_n10934_, new_n10935_,
    new_n10936_, new_n10937_, new_n10938_, new_n10939_, new_n10940_,
    new_n10941_, new_n10942_, new_n10943_, new_n10944_, new_n10945_,
    new_n10946_, new_n10947_, new_n10948_, new_n10949_, new_n10950_,
    new_n10951_, new_n10952_, new_n10953_, new_n10954_, new_n10955_,
    new_n10956_, new_n10957_, new_n10958_, new_n10959_, new_n10960_,
    new_n10961_, new_n10962_, new_n10963_, new_n10964_, new_n10965_,
    new_n10966_, new_n10967_, new_n10968_, new_n10969_, new_n10970_,
    new_n10971_, new_n10972_, new_n10973_, new_n10974_, new_n10975_,
    new_n10976_, new_n10977_, new_n10978_, new_n10979_, new_n10980_,
    new_n10981_, new_n10982_, new_n10983_, new_n10984_, new_n10985_,
    new_n10986_, new_n10987_, new_n10988_, new_n10989_, new_n10990_,
    new_n10991_, new_n10992_, new_n10993_, new_n10994_, new_n10995_,
    new_n10996_, new_n10997_, new_n10998_, new_n10999_, new_n11000_,
    new_n11001_, new_n11002_, new_n11003_, new_n11004_, new_n11005_,
    new_n11006_, new_n11007_, new_n11008_, new_n11009_, new_n11010_,
    new_n11011_, new_n11012_, new_n11013_, new_n11014_, new_n11015_,
    new_n11016_, new_n11017_, new_n11018_, new_n11019_, new_n11020_,
    new_n11021_, new_n11022_, new_n11023_, new_n11024_, new_n11025_,
    new_n11026_, new_n11027_, new_n11028_, new_n11029_, new_n11030_,
    new_n11031_, new_n11032_, new_n11033_, new_n11034_, new_n11035_,
    new_n11036_, new_n11037_, new_n11038_, new_n11039_, new_n11040_,
    new_n11041_, new_n11042_, new_n11043_, new_n11044_, new_n11045_,
    new_n11046_, new_n11047_, new_n11048_, new_n11049_, new_n11050_,
    new_n11051_, new_n11052_, new_n11053_, new_n11054_, new_n11055_,
    new_n11056_, new_n11057_, new_n11058_, new_n11059_, new_n11060_,
    new_n11061_, new_n11062_, new_n11063_, new_n11064_, new_n11065_,
    new_n11066_, new_n11067_, new_n11068_, new_n11069_, new_n11070_,
    new_n11071_, new_n11072_, new_n11073_, new_n11074_, new_n11075_,
    new_n11076_, new_n11077_, new_n11078_, new_n11079_, new_n11080_,
    new_n11081_, new_n11082_, new_n11083_, new_n11084_, new_n11085_,
    new_n11086_, new_n11087_, new_n11088_, new_n11089_, new_n11090_,
    new_n11091_, new_n11092_, new_n11093_, new_n11094_, new_n11095_,
    new_n11096_, new_n11097_, new_n11098_, new_n11099_, new_n11100_,
    new_n11101_, new_n11102_, new_n11103_, new_n11104_, new_n11105_,
    new_n11106_, new_n11107_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11297_, new_n11298_, new_n11299_, new_n11300_,
    new_n11301_, new_n11302_, new_n11303_, new_n11304_, new_n11305_,
    new_n11306_, new_n11307_, new_n11308_, new_n11309_, new_n11310_,
    new_n11311_, new_n11312_, new_n11313_, new_n11314_, new_n11315_,
    new_n11316_, new_n11317_, new_n11318_, new_n11319_, new_n11320_,
    new_n11321_, new_n11322_, new_n11323_, new_n11324_, new_n11325_,
    new_n11326_, new_n11327_, new_n11328_, new_n11329_, new_n11330_,
    new_n11331_, new_n11332_, new_n11333_, new_n11334_, new_n11335_,
    new_n11336_, new_n11337_, new_n11338_, new_n11339_, new_n11340_,
    new_n11341_, new_n11342_, new_n11343_, new_n11344_, new_n11345_,
    new_n11346_, new_n11347_, new_n11348_, new_n11349_, new_n11350_,
    new_n11351_, new_n11352_, new_n11353_, new_n11354_, new_n11355_,
    new_n11356_, new_n11357_, new_n11358_, new_n11359_, new_n11360_,
    new_n11361_, new_n11362_, new_n11363_, new_n11364_, new_n11365_,
    new_n11366_, new_n11367_, new_n11368_, new_n11369_, new_n11370_,
    new_n11371_, new_n11372_, new_n11373_, new_n11374_, new_n11375_,
    new_n11376_, new_n11377_, new_n11378_, new_n11379_, new_n11380_,
    new_n11381_, new_n11382_, new_n11383_, new_n11384_, new_n11385_,
    new_n11386_, new_n11387_, new_n11388_, new_n11389_, new_n11390_,
    new_n11391_, new_n11392_, new_n11393_, new_n11394_, new_n11395_,
    new_n11396_, new_n11397_, new_n11398_, new_n11399_, new_n11400_,
    new_n11401_, new_n11402_, new_n11403_, new_n11404_, new_n11405_,
    new_n11406_, new_n11407_, new_n11408_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11447_, new_n11448_, new_n11449_, new_n11450_,
    new_n11451_, new_n11452_, new_n11453_, new_n11454_, new_n11455_,
    new_n11456_, new_n11457_, new_n11458_, new_n11459_, new_n11460_,
    new_n11461_, new_n11462_, new_n11463_, new_n11464_, new_n11465_,
    new_n11466_, new_n11467_, new_n11468_, new_n11469_, new_n11470_,
    new_n11471_, new_n11472_, new_n11473_, new_n11474_, new_n11475_,
    new_n11476_, new_n11477_, new_n11478_, new_n11479_, new_n11480_,
    new_n11481_, new_n11482_, new_n11483_, new_n11484_, new_n11485_,
    new_n11486_, new_n11487_, new_n11488_, new_n11489_, new_n11490_,
    new_n11491_, new_n11492_, new_n11493_, new_n11494_, new_n11495_,
    new_n11496_, new_n11497_, new_n11498_, new_n11499_, new_n11500_,
    new_n11501_, new_n11502_, new_n11503_, new_n11504_, new_n11505_,
    new_n11506_, new_n11507_, new_n11508_, new_n11509_, new_n11510_,
    new_n11511_, new_n11512_, new_n11513_, new_n11514_, new_n11515_,
    new_n11516_, new_n11517_, new_n11518_, new_n11519_, new_n11520_,
    new_n11521_, new_n11522_, new_n11523_, new_n11524_, new_n11525_,
    new_n11526_, new_n11527_, new_n11528_, new_n11529_, new_n11530_,
    new_n11531_, new_n11532_, new_n11533_, new_n11534_, new_n11535_,
    new_n11536_, new_n11537_, new_n11538_, new_n11539_, new_n11540_,
    new_n11541_, new_n11542_, new_n11543_, new_n11544_, new_n11545_,
    new_n11546_, new_n11547_, new_n11548_, new_n11549_, new_n11550_,
    new_n11551_, new_n11552_, new_n11553_, new_n11554_, new_n11555_,
    new_n11556_, new_n11557_, new_n11558_, new_n11559_, new_n11560_,
    new_n11561_, new_n11562_, new_n11563_, new_n11564_, new_n11565_,
    new_n11566_, new_n11567_, new_n11568_, new_n11569_, new_n11570_,
    new_n11571_, new_n11572_, new_n11573_, new_n11574_, new_n11575_,
    new_n11576_, new_n11577_, new_n11578_, new_n11579_, new_n11580_,
    new_n11581_, new_n11582_, new_n11583_, new_n11584_, new_n11585_,
    new_n11586_, new_n11587_, new_n11588_, new_n11589_, new_n11590_,
    new_n11591_, new_n11592_, new_n11593_, new_n11594_, new_n11595_,
    new_n11596_, new_n11597_, new_n11598_, new_n11599_, new_n11600_,
    new_n11601_, new_n11602_, new_n11603_, new_n11604_, new_n11605_,
    new_n11606_, new_n11607_, new_n11608_, new_n11609_, new_n11610_,
    new_n11611_, new_n11612_, new_n11613_, new_n11614_, new_n11615_,
    new_n11616_, new_n11617_, new_n11618_, new_n11619_, new_n11620_,
    new_n11621_, new_n11622_, new_n11623_, new_n11624_, new_n11625_,
    new_n11626_, new_n11627_, new_n11628_, new_n11629_, new_n11630_,
    new_n11631_, new_n11632_, new_n11633_, new_n11634_, new_n11635_,
    new_n11636_, new_n11637_, new_n11638_, new_n11639_, new_n11640_,
    new_n11641_, new_n11642_, new_n11643_, new_n11644_, new_n11645_,
    new_n11646_, new_n11647_, new_n11648_, new_n11649_, new_n11650_,
    new_n11651_, new_n11652_, new_n11653_, new_n11654_, new_n11655_,
    new_n11656_, new_n11657_, new_n11658_, new_n11659_, new_n11660_,
    new_n11661_, new_n11662_, new_n11663_, new_n11664_, new_n11665_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11730_,
    new_n11731_, new_n11732_, new_n11733_, new_n11734_, new_n11735_,
    new_n11736_, new_n11737_, new_n11738_, new_n11739_, new_n11740_,
    new_n11741_, new_n11742_, new_n11743_, new_n11744_, new_n11745_,
    new_n11746_, new_n11747_, new_n11748_, new_n11749_, new_n11750_,
    new_n11751_, new_n11752_, new_n11753_, new_n11754_, new_n11755_,
    new_n11756_, new_n11757_, new_n11758_, new_n11759_, new_n11760_,
    new_n11761_, new_n11762_, new_n11763_, new_n11764_, new_n11765_,
    new_n11766_, new_n11767_, new_n11768_, new_n11769_, new_n11770_,
    new_n11771_, new_n11772_, new_n11773_, new_n11774_, new_n11775_,
    new_n11776_, new_n11777_, new_n11778_, new_n11779_, new_n11780_,
    new_n11781_, new_n11782_, new_n11783_, new_n11784_, new_n11785_,
    new_n11786_, new_n11787_, new_n11788_, new_n11789_, new_n11790_,
    new_n11791_, new_n11792_, new_n11793_, new_n11794_, new_n11795_,
    new_n11796_, new_n11797_, new_n11798_, new_n11799_, new_n11800_,
    new_n11801_, new_n11802_, new_n11803_, new_n11804_, new_n11805_,
    new_n11806_, new_n11807_, new_n11808_, new_n11809_, new_n11810_,
    new_n11811_, new_n11812_, new_n11813_, new_n11814_, new_n11815_,
    new_n11816_, new_n11817_, new_n11818_, new_n11819_, new_n11820_,
    new_n11821_, new_n11822_, new_n11823_, new_n11824_, new_n11825_,
    new_n11826_, new_n11827_, new_n11828_, new_n11829_, new_n11830_,
    new_n11831_, new_n11832_, new_n11833_, new_n11834_, new_n11835_,
    new_n11836_, new_n11837_, new_n11838_, new_n11839_, new_n11840_,
    new_n11841_, new_n11842_, new_n11843_, new_n11844_, new_n11845_,
    new_n11846_, new_n11847_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11976_, new_n11977_, new_n11978_, new_n11979_, new_n11980_,
    new_n11981_, new_n11982_, new_n11983_, new_n11984_, new_n11985_,
    new_n11986_, new_n11987_, new_n11988_, new_n11989_, new_n11990_,
    new_n11991_, new_n11992_, new_n11993_, new_n11994_, new_n11995_,
    new_n11996_, new_n11997_, new_n11998_, new_n11999_, new_n12000_,
    new_n12001_, new_n12002_, new_n12003_, new_n12004_, new_n12005_,
    new_n12006_, new_n12007_, new_n12008_, new_n12009_, new_n12010_,
    new_n12011_, new_n12012_, new_n12013_, new_n12014_, new_n12015_,
    new_n12016_, new_n12017_, new_n12018_, new_n12019_, new_n12020_,
    new_n12021_, new_n12022_, new_n12023_, new_n12024_, new_n12025_,
    new_n12026_, new_n12027_, new_n12028_, new_n12029_, new_n12030_,
    new_n12031_, new_n12032_, new_n12033_, new_n12034_, new_n12035_,
    new_n12036_, new_n12037_, new_n12038_, new_n12039_, new_n12040_,
    new_n12041_, new_n12042_, new_n12043_, new_n12044_, new_n12045_,
    new_n12046_, new_n12047_, new_n12048_, new_n12049_, new_n12050_,
    new_n12051_, new_n12052_, new_n12053_, new_n12054_, new_n12055_,
    new_n12056_, new_n12057_, new_n12058_, new_n12059_, new_n12060_,
    new_n12061_, new_n12062_, new_n12063_, new_n12064_, new_n12065_,
    new_n12066_, new_n12067_, new_n12068_, new_n12069_, new_n12070_,
    new_n12071_, new_n12072_, new_n12073_, new_n12074_, new_n12075_,
    new_n12076_, new_n12077_, new_n12078_, new_n12079_, new_n12080_,
    new_n12081_, new_n12082_, new_n12083_, new_n12084_, new_n12085_,
    new_n12086_, new_n12087_, new_n12088_, new_n12089_, new_n12090_,
    new_n12091_, new_n12092_, new_n12093_, new_n12094_, new_n12095_,
    new_n12096_, new_n12097_, new_n12098_, new_n12099_, new_n12100_,
    new_n12101_, new_n12102_, new_n12103_, new_n12104_, new_n12105_,
    new_n12106_, new_n12107_, new_n12108_, new_n12109_, new_n12110_,
    new_n12111_, new_n12112_, new_n12113_, new_n12114_, new_n12115_,
    new_n12116_, new_n12117_, new_n12118_, new_n12119_, new_n12120_,
    new_n12121_, new_n12122_, new_n12123_, new_n12124_, new_n12125_,
    new_n12126_, new_n12127_, new_n12128_, new_n12129_, new_n12130_,
    new_n12131_, new_n12132_, new_n12133_, new_n12134_, new_n12135_,
    new_n12136_, new_n12137_, new_n12138_, new_n12139_, new_n12140_,
    new_n12141_, new_n12142_, new_n12143_, new_n12144_, new_n12145_,
    new_n12146_, new_n12147_, new_n12148_, new_n12149_, new_n12150_,
    new_n12151_, new_n12152_, new_n12153_, new_n12154_, new_n12155_,
    new_n12156_, new_n12157_, new_n12158_, new_n12159_, new_n12160_,
    new_n12161_, new_n12162_, new_n12163_, new_n12164_, new_n12165_,
    new_n12166_, new_n12167_, new_n12168_, new_n12169_, new_n12170_,
    new_n12171_, new_n12172_, new_n12173_, new_n12174_, new_n12175_,
    new_n12176_, new_n12177_, new_n12178_, new_n12179_, new_n12180_,
    new_n12181_, new_n12182_, new_n12183_, new_n12184_, new_n12185_,
    new_n12186_, new_n12187_, new_n12188_, new_n12189_, new_n12190_,
    new_n12191_, new_n12192_, new_n12193_, new_n12194_, new_n12195_,
    new_n12196_, new_n12197_, new_n12198_, new_n12199_, new_n12200_,
    new_n12201_, new_n12202_, new_n12203_, new_n12204_, new_n12205_,
    new_n12206_, new_n12207_, new_n12208_, new_n12209_, new_n12210_,
    new_n12211_, new_n12212_, new_n12213_, new_n12214_, new_n12215_,
    new_n12216_, new_n12217_, new_n12218_, new_n12219_, new_n12220_,
    new_n12221_, new_n12222_, new_n12223_, new_n12224_, new_n12225_,
    new_n12226_, new_n12227_, new_n12228_, new_n12229_, new_n12230_,
    new_n12231_, new_n12232_, new_n12233_, new_n12234_, new_n12235_,
    new_n12236_, new_n12237_, new_n12238_, new_n12239_, new_n12240_,
    new_n12241_, new_n12242_, new_n12243_, new_n12244_, new_n12245_,
    new_n12246_, new_n12247_, new_n12248_, new_n12249_, new_n12250_,
    new_n12251_, new_n12252_, new_n12253_, new_n12254_, new_n12255_,
    new_n12256_, new_n12257_, new_n12258_, new_n12259_, new_n12260_,
    new_n12261_, new_n12262_, new_n12263_, new_n12264_, new_n12265_,
    new_n12266_, new_n12267_, new_n12268_, new_n12269_, new_n12270_,
    new_n12271_, new_n12272_, new_n12273_, new_n12274_, new_n12275_,
    new_n12276_, new_n12277_, new_n12278_, new_n12279_, new_n12280_,
    new_n12281_, new_n12282_, new_n12283_, new_n12284_, new_n12285_,
    new_n12286_, new_n12287_, new_n12288_, new_n12289_, new_n12290_,
    new_n12291_, new_n12292_, new_n12293_, new_n12294_, new_n12295_,
    new_n12296_, new_n12297_, new_n12298_, new_n12299_, new_n12300_,
    new_n12301_, new_n12302_, new_n12303_, new_n12304_, new_n12305_,
    new_n12306_, new_n12307_, new_n12308_, new_n12309_, new_n12310_,
    new_n12311_, new_n12312_, new_n12313_, new_n12314_, new_n12315_,
    new_n12316_, new_n12317_, new_n12318_, new_n12319_, new_n12320_,
    new_n12321_, new_n12322_, new_n12323_, new_n12324_, new_n12325_,
    new_n12326_, new_n12327_, new_n12328_, new_n12329_, new_n12330_,
    new_n12331_, new_n12332_, new_n12333_, new_n12334_, new_n12335_,
    new_n12336_, new_n12337_, new_n12338_, new_n12339_, new_n12340_,
    new_n12341_, new_n12342_, new_n12343_, new_n12344_, new_n12345_,
    new_n12346_, new_n12347_, new_n12348_, new_n12349_, new_n12350_,
    new_n12351_, new_n12352_, new_n12353_, new_n12354_, new_n12355_,
    new_n12356_, new_n12357_, new_n12358_, new_n12359_, new_n12360_,
    new_n12361_, new_n12362_, new_n12363_, new_n12364_, new_n12365_,
    new_n12366_, new_n12367_, new_n12368_, new_n12369_, new_n12370_,
    new_n12371_, new_n12372_, new_n12373_, new_n12374_, new_n12375_,
    new_n12376_, new_n12377_, new_n12378_, new_n12379_, new_n12380_,
    new_n12381_, new_n12382_, new_n12383_, new_n12384_, new_n12385_,
    new_n12386_, new_n12387_, new_n12388_, new_n12389_, new_n12390_,
    new_n12391_, new_n12392_, new_n12393_, new_n12394_, new_n12395_,
    new_n12396_, new_n12397_, new_n12398_, new_n12399_, new_n12400_,
    new_n12401_, new_n12402_, new_n12403_, new_n12404_, new_n12405_,
    new_n12406_, new_n12407_, new_n12408_, new_n12409_, new_n12410_,
    new_n12411_, new_n12412_, new_n12413_, new_n12414_, new_n12415_,
    new_n12416_, new_n12417_, new_n12418_, new_n12419_, new_n12420_,
    new_n12421_, new_n12422_, new_n12423_, new_n12424_, new_n12425_,
    new_n12426_, new_n12427_, new_n12428_, new_n12429_, new_n12430_,
    new_n12431_, new_n12432_, new_n12433_, new_n12434_, new_n12435_,
    new_n12436_, new_n12437_, new_n12438_, new_n12439_, new_n12440_,
    new_n12441_, new_n12442_, new_n12443_, new_n12444_, new_n12445_,
    new_n12446_, new_n12447_, new_n12448_, new_n12449_, new_n12450_,
    new_n12451_, new_n12452_, new_n12453_, new_n12454_, new_n12455_,
    new_n12456_, new_n12457_, new_n12458_, new_n12459_, new_n12460_,
    new_n12461_, new_n12462_, new_n12463_, new_n12464_, new_n12465_,
    new_n12466_, new_n12467_, new_n12468_, new_n12469_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12581_, new_n12582_, new_n12583_, new_n12584_, new_n12585_,
    new_n12586_, new_n12587_, new_n12588_, new_n12589_, new_n12590_,
    new_n12591_, new_n12592_, new_n12593_, new_n12594_, new_n12595_,
    new_n12596_, new_n12597_, new_n12598_, new_n12599_, new_n12600_,
    new_n12601_, new_n12602_, new_n12603_, new_n12604_, new_n12605_,
    new_n12606_, new_n12607_, new_n12608_, new_n12609_, new_n12610_,
    new_n12611_, new_n12612_, new_n12613_, new_n12614_, new_n12615_,
    new_n12616_, new_n12617_, new_n12618_, new_n12619_, new_n12620_,
    new_n12621_, new_n12622_, new_n12623_, new_n12624_, new_n12625_,
    new_n12626_, new_n12627_, new_n12628_, new_n12629_, new_n12630_,
    new_n12631_, new_n12632_, new_n12633_, new_n12634_, new_n12635_,
    new_n12636_, new_n12637_, new_n12638_, new_n12639_, new_n12640_,
    new_n12641_, new_n12642_, new_n12643_, new_n12644_, new_n12645_,
    new_n12646_, new_n12647_, new_n12648_, new_n12649_, new_n12650_,
    new_n12651_, new_n12652_, new_n12653_, new_n12654_, new_n12655_,
    new_n12656_, new_n12657_, new_n12658_, new_n12659_, new_n12660_,
    new_n12661_, new_n12662_, new_n12663_, new_n12664_, new_n12665_,
    new_n12666_, new_n12667_, new_n12668_, new_n12669_, new_n12670_,
    new_n12671_, new_n12672_, new_n12673_, new_n12674_, new_n12675_,
    new_n12676_, new_n12677_, new_n12678_, new_n12679_, new_n12680_,
    new_n12681_, new_n12682_, new_n12683_, new_n12684_, new_n12685_,
    new_n12686_, new_n12687_, new_n12688_, new_n12689_, new_n12690_,
    new_n12691_, new_n12692_, new_n12693_, new_n12694_, new_n12695_,
    new_n12696_, new_n12697_, new_n12698_, new_n12699_, new_n12700_,
    new_n12701_, new_n12702_, new_n12703_, new_n12704_, new_n12705_,
    new_n12706_, new_n12707_, new_n12708_, new_n12709_, new_n12710_,
    new_n12711_, new_n12712_, new_n12713_, new_n12714_, new_n12715_,
    new_n12716_, new_n12717_, new_n12718_, new_n12719_, new_n12720_,
    new_n12721_, new_n12722_, new_n12723_, new_n12724_, new_n12725_,
    new_n12726_, new_n12727_, new_n12728_, new_n12729_, new_n12730_,
    new_n12731_, new_n12732_, new_n12733_, new_n12734_, new_n12735_,
    new_n12736_, new_n12737_, new_n12738_, new_n12739_, new_n12740_,
    new_n12741_, new_n12742_, new_n12743_, new_n12744_, new_n12745_,
    new_n12746_, new_n12747_, new_n12748_, new_n12749_, new_n12750_,
    new_n12751_, new_n12752_, new_n12753_, new_n12754_, new_n12755_,
    new_n12756_, new_n12757_, new_n12758_, new_n12759_, new_n12760_,
    new_n12761_, new_n12762_, new_n12763_, new_n12764_, new_n12765_,
    new_n12766_, new_n12767_, new_n12768_, new_n12769_, new_n12770_,
    new_n12771_, new_n12772_, new_n12773_, new_n12774_, new_n12775_,
    new_n12776_, new_n12777_, new_n12778_, new_n12779_, new_n12780_,
    new_n12781_, new_n12782_, new_n12783_, new_n12784_, new_n12785_,
    new_n12786_, new_n12787_, new_n12788_, new_n12789_, new_n12790_,
    new_n12791_, new_n12792_, new_n12793_, new_n12794_, new_n12795_,
    new_n12796_, new_n12797_, new_n12798_, new_n12799_, new_n12800_,
    new_n12801_, new_n12802_, new_n12803_, new_n12804_, new_n12805_,
    new_n12806_, new_n12807_, new_n12808_, new_n12809_, new_n12810_,
    new_n12811_, new_n12812_, new_n12813_, new_n12814_, new_n12815_,
    new_n12816_, new_n12817_, new_n12818_, new_n12819_, new_n12820_,
    new_n12821_, new_n12822_, new_n12823_, new_n12824_, new_n12825_,
    new_n12826_, new_n12827_, new_n12828_, new_n12829_, new_n12830_,
    new_n12831_, new_n12832_, new_n12833_, new_n12834_, new_n12835_,
    new_n12836_, new_n12837_, new_n12838_, new_n12839_, new_n12840_,
    new_n12841_, new_n12842_, new_n12843_, new_n12844_, new_n12845_,
    new_n12846_, new_n12847_, new_n12848_, new_n12849_, new_n12850_,
    new_n12851_, new_n12852_, new_n12853_, new_n12854_, new_n12855_,
    new_n12856_, new_n12857_, new_n12858_, new_n12859_, new_n12860_,
    new_n12861_, new_n12862_, new_n12863_, new_n12864_, new_n12865_,
    new_n12866_, new_n12867_, new_n12868_, new_n12869_, new_n12870_,
    new_n12871_, new_n12872_, new_n12873_, new_n12874_, new_n12875_,
    new_n12876_, new_n12877_, new_n12878_, new_n12879_, new_n12880_,
    new_n12881_, new_n12882_, new_n12883_, new_n12884_, new_n12885_,
    new_n12886_, new_n12887_, new_n12888_, new_n12889_, new_n12890_,
    new_n12891_, new_n12892_, new_n12893_, new_n12894_, new_n12895_,
    new_n12896_, new_n12897_, new_n12898_, new_n12899_, new_n12900_,
    new_n12901_, new_n12902_, new_n12903_, new_n12904_, new_n12905_,
    new_n12906_, new_n12907_, new_n12908_, new_n12909_, new_n12910_,
    new_n12911_, new_n12912_, new_n12913_, new_n12914_, new_n12915_,
    new_n12916_, new_n12917_, new_n12918_, new_n12919_, new_n12920_,
    new_n12921_, new_n12922_, new_n12923_, new_n12924_, new_n12925_,
    new_n12926_, new_n12927_, new_n12928_, new_n12929_, new_n12930_,
    new_n12931_, new_n12932_, new_n12933_, new_n12934_, new_n12935_,
    new_n12936_, new_n12937_, new_n12938_, new_n12939_, new_n12940_,
    new_n12941_, new_n12942_, new_n12943_, new_n12944_, new_n12945_,
    new_n12946_, new_n12947_, new_n12948_, new_n12949_, new_n12950_,
    new_n12951_, new_n12952_, new_n12953_, new_n12954_, new_n12955_,
    new_n12956_, new_n12957_, new_n12958_, new_n12959_, new_n12960_,
    new_n12961_, new_n12962_, new_n12963_, new_n12964_, new_n12965_,
    new_n12966_, new_n12967_, new_n12968_, new_n12969_, new_n12970_,
    new_n12971_, new_n12972_, new_n12973_, new_n12974_, new_n12975_,
    new_n12976_, new_n12977_, new_n12978_, new_n12979_, new_n12980_,
    new_n12981_, new_n12982_, new_n12983_, new_n12984_, new_n12985_,
    new_n12986_, new_n12987_, new_n12988_, new_n12989_, new_n12990_,
    new_n12991_, new_n12992_, new_n12993_, new_n12994_, new_n12995_,
    new_n12996_, new_n12997_, new_n12998_, new_n12999_, new_n13000_,
    new_n13001_, new_n13002_, new_n13003_, new_n13004_, new_n13005_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13337_, new_n13338_, new_n13339_, new_n13340_, new_n13341_,
    new_n13342_, new_n13343_, new_n13344_, new_n13345_, new_n13346_,
    new_n13347_, new_n13348_, new_n13349_, new_n13352_, new_n13353_,
    new_n13354_, new_n13355_, new_n13356_, new_n13357_, new_n13358_;
  INVX1    g00000(.A(\A[716] ), .Y(new_n1003_));
  OR2X1    g00001(.A(new_n1003_), .B(\A[715] ), .Y(new_n1004_));
  INVX1    g00002(.A(\A[717] ), .Y(new_n1005_));
  AOI21X1  g00003(.A0(new_n1003_), .A1(\A[715] ), .B0(new_n1005_), .Y(new_n1006_));
  XOR2X1   g00004(.A(\A[716] ), .B(\A[715] ), .Y(new_n1007_));
  AND2X1   g00005(.A(new_n1007_), .B(new_n1005_), .Y(new_n1008_));
  AOI21X1  g00006(.A0(new_n1006_), .A1(new_n1004_), .B0(new_n1008_), .Y(new_n1009_));
  INVX1    g00007(.A(\A[720] ), .Y(new_n1010_));
  INVX1    g00008(.A(\A[719] ), .Y(new_n1011_));
  OR2X1    g00009(.A(new_n1011_), .B(\A[718] ), .Y(new_n1012_));
  AOI21X1  g00010(.A0(new_n1011_), .A1(\A[718] ), .B0(new_n1010_), .Y(new_n1013_));
  XOR2X1   g00011(.A(\A[719] ), .B(\A[718] ), .Y(new_n1014_));
  AOI22X1  g00012(.A0(new_n1014_), .A1(new_n1010_), .B0(new_n1013_), .B1(new_n1012_), .Y(new_n1015_));
  NOR2X1   g00013(.A(new_n1015_), .B(new_n1009_), .Y(new_n1016_));
  AND2X1   g00014(.A(\A[719] ), .B(\A[718] ), .Y(new_n1017_));
  AND2X1   g00015(.A(new_n1014_), .B(\A[720] ), .Y(new_n1018_));
  OR2X1    g00016(.A(new_n1018_), .B(new_n1017_), .Y(new_n1019_));
  AND2X1   g00017(.A(\A[716] ), .B(\A[715] ), .Y(new_n1020_));
  AOI21X1  g00018(.A0(new_n1007_), .A1(\A[717] ), .B0(new_n1020_), .Y(new_n1021_));
  XOR2X1   g00019(.A(new_n1021_), .B(new_n1019_), .Y(new_n1022_));
  XOR2X1   g00020(.A(new_n1022_), .B(new_n1016_), .Y(new_n1023_));
  XOR2X1   g00021(.A(new_n1015_), .B(new_n1009_), .Y(new_n1024_));
  OR2X1    g00022(.A(new_n1015_), .B(new_n1009_), .Y(new_n1025_));
  AOI21X1  g00023(.A0(new_n1014_), .A1(\A[720] ), .B0(new_n1017_), .Y(new_n1026_));
  OR2X1    g00024(.A(new_n1021_), .B(new_n1026_), .Y(new_n1027_));
  OAI21X1  g00025(.A0(new_n1022_), .A1(new_n1025_), .B0(new_n1027_), .Y(new_n1028_));
  AND2X1   g00026(.A(new_n1028_), .B(new_n1024_), .Y(new_n1029_));
  OR2X1    g00027(.A(new_n1029_), .B(new_n1023_), .Y(new_n1030_));
  AND2X1   g00028(.A(\A[725] ), .B(\A[724] ), .Y(new_n1031_));
  XOR2X1   g00029(.A(\A[725] ), .B(\A[724] ), .Y(new_n1032_));
  AOI21X1  g00030(.A0(new_n1032_), .A1(\A[726] ), .B0(new_n1031_), .Y(new_n1033_));
  AND2X1   g00031(.A(\A[722] ), .B(\A[721] ), .Y(new_n1034_));
  XOR2X1   g00032(.A(\A[722] ), .B(\A[721] ), .Y(new_n1035_));
  AOI21X1  g00033(.A0(new_n1035_), .A1(\A[723] ), .B0(new_n1034_), .Y(new_n1036_));
  INVX1    g00034(.A(\A[722] ), .Y(new_n1037_));
  OR2X1    g00035(.A(new_n1037_), .B(\A[721] ), .Y(new_n1038_));
  INVX1    g00036(.A(\A[723] ), .Y(new_n1039_));
  AOI21X1  g00037(.A0(new_n1037_), .A1(\A[721] ), .B0(new_n1039_), .Y(new_n1040_));
  AND2X1   g00038(.A(new_n1035_), .B(new_n1039_), .Y(new_n1041_));
  AOI21X1  g00039(.A0(new_n1040_), .A1(new_n1038_), .B0(new_n1041_), .Y(new_n1042_));
  INVX1    g00040(.A(\A[726] ), .Y(new_n1043_));
  INVX1    g00041(.A(\A[725] ), .Y(new_n1044_));
  OR2X1    g00042(.A(new_n1044_), .B(\A[724] ), .Y(new_n1045_));
  AOI21X1  g00043(.A0(new_n1044_), .A1(\A[724] ), .B0(new_n1043_), .Y(new_n1046_));
  AOI22X1  g00044(.A0(new_n1046_), .A1(new_n1045_), .B0(new_n1032_), .B1(new_n1043_), .Y(new_n1047_));
  OR4X1    g00045(.A(new_n1047_), .B(new_n1042_), .C(new_n1036_), .D(new_n1033_), .Y(new_n1048_));
  OR4X1    g00046(.A(new_n1021_), .B(new_n1026_), .C(new_n1015_), .D(new_n1009_), .Y(new_n1049_));
  XOR2X1   g00047(.A(new_n1047_), .B(new_n1042_), .Y(new_n1050_));
  NAND4X1  g00048(.A(new_n1050_), .B(new_n1049_), .C(new_n1048_), .D(new_n1024_), .Y(new_n1051_));
  XOR2X1   g00049(.A(new_n1036_), .B(new_n1033_), .Y(new_n1052_));
  NOR2X1   g00050(.A(new_n1047_), .B(new_n1042_), .Y(new_n1053_));
  NOR2X1   g00051(.A(new_n1036_), .B(new_n1033_), .Y(new_n1054_));
  AOI21X1  g00052(.A0(new_n1053_), .A1(new_n1052_), .B0(new_n1054_), .Y(new_n1055_));
  XOR2X1   g00053(.A(new_n1053_), .B(new_n1052_), .Y(new_n1056_));
  AND2X1   g00054(.A(new_n1040_), .B(new_n1038_), .Y(new_n1057_));
  OR2X1    g00055(.A(new_n1041_), .B(new_n1057_), .Y(new_n1058_));
  XOR2X1   g00056(.A(new_n1047_), .B(new_n1058_), .Y(new_n1059_));
  OAI21X1  g00057(.A0(new_n1059_), .A1(new_n1055_), .B0(new_n1056_), .Y(new_n1060_));
  XOR2X1   g00058(.A(new_n1060_), .B(new_n1051_), .Y(new_n1061_));
  AND2X1   g00059(.A(new_n1061_), .B(new_n1030_), .Y(new_n1062_));
  AND2X1   g00060(.A(new_n1006_), .B(new_n1004_), .Y(new_n1063_));
  OR2X1    g00061(.A(new_n1008_), .B(new_n1063_), .Y(new_n1064_));
  XOR2X1   g00062(.A(new_n1015_), .B(new_n1064_), .Y(new_n1065_));
  OR2X1    g00063(.A(new_n1047_), .B(new_n1042_), .Y(new_n1066_));
  XOR2X1   g00064(.A(new_n1066_), .B(new_n1052_), .Y(new_n1067_));
  NOR4X1   g00065(.A(new_n1021_), .B(new_n1026_), .C(new_n1015_), .D(new_n1009_), .Y(new_n1068_));
  NOR4X1   g00066(.A(new_n1059_), .B(new_n1068_), .C(new_n1067_), .D(new_n1065_), .Y(new_n1069_));
  AND2X1   g00067(.A(new_n1053_), .B(new_n1052_), .Y(new_n1070_));
  OAI22X1  g00068(.A0(new_n1050_), .A1(new_n1056_), .B0(new_n1054_), .B1(new_n1070_), .Y(new_n1071_));
  AOI22X1  g00069(.A0(new_n1071_), .A1(new_n1069_), .B0(new_n1060_), .B1(new_n1051_), .Y(new_n1072_));
  AND2X1   g00070(.A(new_n1050_), .B(new_n1048_), .Y(new_n1073_));
  XOR2X1   g00071(.A(new_n1015_), .B(new_n1064_), .Y(new_n1074_));
  XOR2X1   g00072(.A(new_n1074_), .B(new_n1073_), .Y(new_n1075_));
  INVX1    g00073(.A(\A[709] ), .Y(new_n1076_));
  OR2X1    g00074(.A(\A[710] ), .B(new_n1076_), .Y(new_n1077_));
  INVX1    g00075(.A(\A[711] ), .Y(new_n1078_));
  AOI21X1  g00076(.A0(\A[710] ), .A1(new_n1076_), .B0(new_n1078_), .Y(new_n1079_));
  AND2X1   g00077(.A(new_n1079_), .B(new_n1077_), .Y(new_n1080_));
  XOR2X1   g00078(.A(\A[710] ), .B(\A[709] ), .Y(new_n1081_));
  AND2X1   g00079(.A(new_n1081_), .B(new_n1078_), .Y(new_n1082_));
  OR2X1    g00080(.A(new_n1082_), .B(new_n1080_), .Y(new_n1083_));
  INVX1    g00081(.A(\A[714] ), .Y(new_n1084_));
  INVX1    g00082(.A(\A[712] ), .Y(new_n1085_));
  OR2X1    g00083(.A(\A[713] ), .B(new_n1085_), .Y(new_n1086_));
  AOI21X1  g00084(.A0(\A[713] ), .A1(new_n1085_), .B0(new_n1084_), .Y(new_n1087_));
  XOR2X1   g00085(.A(\A[713] ), .B(\A[712] ), .Y(new_n1088_));
  AOI22X1  g00086(.A0(new_n1088_), .A1(new_n1084_), .B0(new_n1087_), .B1(new_n1086_), .Y(new_n1089_));
  AND2X1   g00087(.A(\A[713] ), .B(\A[712] ), .Y(new_n1090_));
  AOI21X1  g00088(.A0(new_n1088_), .A1(\A[714] ), .B0(new_n1090_), .Y(new_n1091_));
  AND2X1   g00089(.A(\A[710] ), .B(\A[709] ), .Y(new_n1092_));
  AOI21X1  g00090(.A0(new_n1081_), .A1(\A[711] ), .B0(new_n1092_), .Y(new_n1093_));
  XOR2X1   g00091(.A(new_n1089_), .B(new_n1083_), .Y(new_n1094_));
  INVX1    g00092(.A(\A[703] ), .Y(new_n1095_));
  OR2X1    g00093(.A(\A[704] ), .B(new_n1095_), .Y(new_n1096_));
  INVX1    g00094(.A(\A[705] ), .Y(new_n1097_));
  AOI21X1  g00095(.A0(\A[704] ), .A1(new_n1095_), .B0(new_n1097_), .Y(new_n1098_));
  XOR2X1   g00096(.A(\A[704] ), .B(\A[703] ), .Y(new_n1099_));
  AND2X1   g00097(.A(new_n1099_), .B(new_n1097_), .Y(new_n1100_));
  AOI21X1  g00098(.A0(new_n1098_), .A1(new_n1096_), .B0(new_n1100_), .Y(new_n1101_));
  INVX1    g00099(.A(\A[708] ), .Y(new_n1102_));
  INVX1    g00100(.A(\A[706] ), .Y(new_n1103_));
  OR2X1    g00101(.A(\A[707] ), .B(new_n1103_), .Y(new_n1104_));
  AOI21X1  g00102(.A0(\A[707] ), .A1(new_n1103_), .B0(new_n1102_), .Y(new_n1105_));
  XOR2X1   g00103(.A(\A[707] ), .B(\A[706] ), .Y(new_n1106_));
  AOI22X1  g00104(.A0(new_n1106_), .A1(new_n1102_), .B0(new_n1105_), .B1(new_n1104_), .Y(new_n1107_));
  AND2X1   g00105(.A(\A[707] ), .B(\A[706] ), .Y(new_n1108_));
  AOI21X1  g00106(.A0(new_n1106_), .A1(\A[708] ), .B0(new_n1108_), .Y(new_n1109_));
  AND2X1   g00107(.A(\A[704] ), .B(\A[703] ), .Y(new_n1110_));
  AOI21X1  g00108(.A0(new_n1099_), .A1(\A[705] ), .B0(new_n1110_), .Y(new_n1111_));
  XOR2X1   g00109(.A(new_n1107_), .B(new_n1101_), .Y(new_n1112_));
  XOR2X1   g00110(.A(new_n1112_), .B(new_n1094_), .Y(new_n1113_));
  NOR2X1   g00111(.A(new_n1113_), .B(new_n1075_), .Y(new_n1114_));
  OAI21X1  g00112(.A0(new_n1072_), .A1(new_n1030_), .B0(new_n1114_), .Y(new_n1115_));
  NOR2X1   g00113(.A(new_n1072_), .B(new_n1030_), .Y(new_n1116_));
  OR2X1    g00114(.A(new_n1113_), .B(new_n1075_), .Y(new_n1117_));
  OAI21X1  g00115(.A0(new_n1116_), .A1(new_n1062_), .B0(new_n1117_), .Y(new_n1118_));
  OAI21X1  g00116(.A0(new_n1115_), .A1(new_n1062_), .B0(new_n1118_), .Y(new_n1119_));
  AND2X1   g00117(.A(new_n1098_), .B(new_n1096_), .Y(new_n1120_));
  OR2X1    g00118(.A(new_n1100_), .B(new_n1120_), .Y(new_n1121_));
  XOR2X1   g00119(.A(new_n1107_), .B(new_n1121_), .Y(new_n1122_));
  XOR2X1   g00120(.A(new_n1111_), .B(new_n1109_), .Y(new_n1123_));
  NOR2X1   g00121(.A(new_n1107_), .B(new_n1101_), .Y(new_n1124_));
  NOR2X1   g00122(.A(new_n1111_), .B(new_n1109_), .Y(new_n1125_));
  AOI21X1  g00123(.A0(new_n1124_), .A1(new_n1123_), .B0(new_n1125_), .Y(new_n1126_));
  XOR2X1   g00124(.A(new_n1124_), .B(new_n1123_), .Y(new_n1127_));
  OAI21X1  g00125(.A0(new_n1126_), .A1(new_n1122_), .B0(new_n1127_), .Y(new_n1128_));
  INVX1    g00126(.A(new_n1128_), .Y(new_n1129_));
  XOR2X1   g00127(.A(new_n1089_), .B(new_n1083_), .Y(new_n1130_));
  AOI21X1  g00128(.A0(new_n1079_), .A1(new_n1077_), .B0(new_n1082_), .Y(new_n1131_));
  NOR4X1   g00129(.A(new_n1093_), .B(new_n1091_), .C(new_n1089_), .D(new_n1131_), .Y(new_n1132_));
  NOR4X1   g00130(.A(new_n1111_), .B(new_n1109_), .C(new_n1107_), .D(new_n1101_), .Y(new_n1133_));
  OR4X1    g00131(.A(new_n1133_), .B(new_n1122_), .C(new_n1132_), .D(new_n1130_), .Y(new_n1134_));
  XOR2X1   g00132(.A(new_n1093_), .B(new_n1091_), .Y(new_n1135_));
  NOR2X1   g00133(.A(new_n1089_), .B(new_n1131_), .Y(new_n1136_));
  NOR2X1   g00134(.A(new_n1093_), .B(new_n1091_), .Y(new_n1137_));
  AOI21X1  g00135(.A0(new_n1136_), .A1(new_n1135_), .B0(new_n1137_), .Y(new_n1138_));
  XOR2X1   g00136(.A(new_n1136_), .B(new_n1135_), .Y(new_n1139_));
  OAI21X1  g00137(.A0(new_n1138_), .A1(new_n1130_), .B0(new_n1139_), .Y(new_n1140_));
  XOR2X1   g00138(.A(new_n1140_), .B(new_n1134_), .Y(new_n1141_));
  AND2X1   g00139(.A(new_n1141_), .B(new_n1128_), .Y(new_n1142_));
  AND2X1   g00140(.A(new_n1140_), .B(new_n1134_), .Y(new_n1143_));
  OR2X1    g00141(.A(new_n1089_), .B(new_n1131_), .Y(new_n1144_));
  XOR2X1   g00142(.A(new_n1144_), .B(new_n1135_), .Y(new_n1145_));
  OR4X1    g00143(.A(new_n1122_), .B(new_n1132_), .C(new_n1145_), .D(new_n1130_), .Y(new_n1146_));
  INVX1    g00144(.A(new_n1123_), .Y(new_n1147_));
  XOR2X1   g00145(.A(new_n1124_), .B(new_n1147_), .Y(new_n1148_));
  OAI22X1  g00146(.A0(new_n1148_), .A1(new_n1126_), .B0(new_n1138_), .B1(new_n1130_), .Y(new_n1149_));
  NOR2X1   g00147(.A(new_n1149_), .B(new_n1146_), .Y(new_n1150_));
  OR2X1    g00148(.A(new_n1150_), .B(new_n1143_), .Y(new_n1151_));
  AOI21X1  g00149(.A0(new_n1151_), .A1(new_n1129_), .B0(new_n1142_), .Y(new_n1152_));
  NAND2X1  g00150(.A(new_n1061_), .B(new_n1030_), .Y(new_n1153_));
  OR2X1    g00151(.A(new_n1072_), .B(new_n1030_), .Y(new_n1154_));
  NAND3X1  g00152(.A(new_n1117_), .B(new_n1154_), .C(new_n1153_), .Y(new_n1155_));
  OAI21X1  g00153(.A0(new_n1116_), .A1(new_n1062_), .B0(new_n1114_), .Y(new_n1156_));
  AOI21X1  g00154(.A0(new_n1156_), .A1(new_n1155_), .B0(new_n1152_), .Y(new_n1157_));
  AOI21X1  g00155(.A0(new_n1152_), .A1(new_n1119_), .B0(new_n1157_), .Y(new_n1158_));
  INVX1    g00156(.A(\A[728] ), .Y(new_n1159_));
  OR2X1    g00157(.A(new_n1159_), .B(\A[727] ), .Y(new_n1160_));
  INVX1    g00158(.A(\A[729] ), .Y(new_n1161_));
  AOI21X1  g00159(.A0(new_n1159_), .A1(\A[727] ), .B0(new_n1161_), .Y(new_n1162_));
  XOR2X1   g00160(.A(\A[728] ), .B(\A[727] ), .Y(new_n1163_));
  AND2X1   g00161(.A(new_n1163_), .B(new_n1161_), .Y(new_n1164_));
  AOI21X1  g00162(.A0(new_n1162_), .A1(new_n1160_), .B0(new_n1164_), .Y(new_n1165_));
  INVX1    g00163(.A(\A[732] ), .Y(new_n1166_));
  INVX1    g00164(.A(\A[731] ), .Y(new_n1167_));
  OR2X1    g00165(.A(new_n1167_), .B(\A[730] ), .Y(new_n1168_));
  AOI21X1  g00166(.A0(new_n1167_), .A1(\A[730] ), .B0(new_n1166_), .Y(new_n1169_));
  XOR2X1   g00167(.A(\A[731] ), .B(\A[730] ), .Y(new_n1170_));
  AOI22X1  g00168(.A0(new_n1170_), .A1(new_n1166_), .B0(new_n1169_), .B1(new_n1168_), .Y(new_n1171_));
  OR2X1    g00169(.A(new_n1171_), .B(new_n1165_), .Y(new_n1172_));
  AND2X1   g00170(.A(\A[731] ), .B(\A[730] ), .Y(new_n1173_));
  AND2X1   g00171(.A(new_n1170_), .B(\A[732] ), .Y(new_n1174_));
  OR2X1    g00172(.A(new_n1174_), .B(new_n1173_), .Y(new_n1175_));
  AND2X1   g00173(.A(\A[728] ), .B(\A[727] ), .Y(new_n1176_));
  AOI21X1  g00174(.A0(new_n1163_), .A1(\A[729] ), .B0(new_n1176_), .Y(new_n1177_));
  XOR2X1   g00175(.A(new_n1177_), .B(new_n1175_), .Y(new_n1178_));
  XOR2X1   g00176(.A(new_n1178_), .B(new_n1172_), .Y(new_n1179_));
  XOR2X1   g00177(.A(new_n1171_), .B(new_n1165_), .Y(new_n1180_));
  AOI21X1  g00178(.A0(new_n1170_), .A1(\A[732] ), .B0(new_n1173_), .Y(new_n1181_));
  OR2X1    g00179(.A(new_n1177_), .B(new_n1181_), .Y(new_n1182_));
  OAI21X1  g00180(.A0(new_n1178_), .A1(new_n1172_), .B0(new_n1182_), .Y(new_n1183_));
  NAND2X1  g00181(.A(new_n1183_), .B(new_n1180_), .Y(new_n1184_));
  NAND2X1  g00182(.A(new_n1184_), .B(new_n1179_), .Y(new_n1185_));
  AND2X1   g00183(.A(\A[737] ), .B(\A[736] ), .Y(new_n1186_));
  XOR2X1   g00184(.A(\A[737] ), .B(\A[736] ), .Y(new_n1187_));
  AOI21X1  g00185(.A0(new_n1187_), .A1(\A[738] ), .B0(new_n1186_), .Y(new_n1188_));
  AND2X1   g00186(.A(\A[734] ), .B(\A[733] ), .Y(new_n1189_));
  XOR2X1   g00187(.A(\A[734] ), .B(\A[733] ), .Y(new_n1190_));
  AOI21X1  g00188(.A0(new_n1190_), .A1(\A[735] ), .B0(new_n1189_), .Y(new_n1191_));
  INVX1    g00189(.A(\A[734] ), .Y(new_n1192_));
  OR2X1    g00190(.A(new_n1192_), .B(\A[733] ), .Y(new_n1193_));
  INVX1    g00191(.A(\A[735] ), .Y(new_n1194_));
  AOI21X1  g00192(.A0(new_n1192_), .A1(\A[733] ), .B0(new_n1194_), .Y(new_n1195_));
  AND2X1   g00193(.A(new_n1190_), .B(new_n1194_), .Y(new_n1196_));
  AOI21X1  g00194(.A0(new_n1195_), .A1(new_n1193_), .B0(new_n1196_), .Y(new_n1197_));
  INVX1    g00195(.A(\A[738] ), .Y(new_n1198_));
  INVX1    g00196(.A(\A[737] ), .Y(new_n1199_));
  OR2X1    g00197(.A(new_n1199_), .B(\A[736] ), .Y(new_n1200_));
  AOI21X1  g00198(.A0(new_n1199_), .A1(\A[736] ), .B0(new_n1198_), .Y(new_n1201_));
  AOI22X1  g00199(.A0(new_n1201_), .A1(new_n1200_), .B0(new_n1187_), .B1(new_n1198_), .Y(new_n1202_));
  OR4X1    g00200(.A(new_n1202_), .B(new_n1197_), .C(new_n1191_), .D(new_n1188_), .Y(new_n1203_));
  OR4X1    g00201(.A(new_n1177_), .B(new_n1181_), .C(new_n1171_), .D(new_n1165_), .Y(new_n1204_));
  XOR2X1   g00202(.A(new_n1202_), .B(new_n1197_), .Y(new_n1205_));
  NAND4X1  g00203(.A(new_n1205_), .B(new_n1204_), .C(new_n1203_), .D(new_n1180_), .Y(new_n1206_));
  XOR2X1   g00204(.A(new_n1191_), .B(new_n1188_), .Y(new_n1207_));
  NOR2X1   g00205(.A(new_n1202_), .B(new_n1197_), .Y(new_n1208_));
  NOR2X1   g00206(.A(new_n1191_), .B(new_n1188_), .Y(new_n1209_));
  AOI21X1  g00207(.A0(new_n1208_), .A1(new_n1207_), .B0(new_n1209_), .Y(new_n1210_));
  XOR2X1   g00208(.A(new_n1208_), .B(new_n1207_), .Y(new_n1211_));
  AND2X1   g00209(.A(new_n1195_), .B(new_n1193_), .Y(new_n1212_));
  OR2X1    g00210(.A(new_n1196_), .B(new_n1212_), .Y(new_n1213_));
  XOR2X1   g00211(.A(new_n1202_), .B(new_n1213_), .Y(new_n1214_));
  OAI21X1  g00212(.A0(new_n1214_), .A1(new_n1210_), .B0(new_n1211_), .Y(new_n1215_));
  XOR2X1   g00213(.A(new_n1215_), .B(new_n1206_), .Y(new_n1216_));
  INVX1    g00214(.A(new_n1206_), .Y(new_n1217_));
  OR2X1    g00215(.A(new_n1202_), .B(new_n1197_), .Y(new_n1218_));
  XOR2X1   g00216(.A(new_n1218_), .B(new_n1207_), .Y(new_n1219_));
  NOR2X1   g00217(.A(new_n1214_), .B(new_n1210_), .Y(new_n1220_));
  NOR2X1   g00218(.A(new_n1220_), .B(new_n1219_), .Y(new_n1221_));
  NOR4X1   g00219(.A(new_n1177_), .B(new_n1181_), .C(new_n1171_), .D(new_n1165_), .Y(new_n1222_));
  NAND2X1  g00220(.A(new_n1205_), .B(new_n1180_), .Y(new_n1223_));
  AOI21X1  g00221(.A0(new_n1214_), .A1(new_n1219_), .B0(new_n1210_), .Y(new_n1224_));
  OR4X1    g00222(.A(new_n1224_), .B(new_n1223_), .C(new_n1222_), .D(new_n1219_), .Y(new_n1225_));
  OAI21X1  g00223(.A0(new_n1221_), .A1(new_n1217_), .B0(new_n1225_), .Y(new_n1226_));
  MX2X1    g00224(.A(new_n1226_), .B(new_n1216_), .S0(new_n1185_), .Y(new_n1227_));
  INVX1    g00225(.A(\A[740] ), .Y(new_n1228_));
  OR2X1    g00226(.A(new_n1228_), .B(\A[739] ), .Y(new_n1229_));
  INVX1    g00227(.A(\A[741] ), .Y(new_n1230_));
  AOI21X1  g00228(.A0(new_n1228_), .A1(\A[739] ), .B0(new_n1230_), .Y(new_n1231_));
  XOR2X1   g00229(.A(\A[740] ), .B(\A[739] ), .Y(new_n1232_));
  AND2X1   g00230(.A(new_n1232_), .B(new_n1230_), .Y(new_n1233_));
  AOI21X1  g00231(.A0(new_n1231_), .A1(new_n1229_), .B0(new_n1233_), .Y(new_n1234_));
  INVX1    g00232(.A(\A[744] ), .Y(new_n1235_));
  INVX1    g00233(.A(\A[743] ), .Y(new_n1236_));
  OR2X1    g00234(.A(new_n1236_), .B(\A[742] ), .Y(new_n1237_));
  AOI21X1  g00235(.A0(new_n1236_), .A1(\A[742] ), .B0(new_n1235_), .Y(new_n1238_));
  XOR2X1   g00236(.A(\A[743] ), .B(\A[742] ), .Y(new_n1239_));
  AOI22X1  g00237(.A0(new_n1239_), .A1(new_n1235_), .B0(new_n1238_), .B1(new_n1237_), .Y(new_n1240_));
  NOR2X1   g00238(.A(new_n1240_), .B(new_n1234_), .Y(new_n1241_));
  AND2X1   g00239(.A(\A[743] ), .B(\A[742] ), .Y(new_n1242_));
  AND2X1   g00240(.A(new_n1239_), .B(\A[744] ), .Y(new_n1243_));
  OR2X1    g00241(.A(new_n1243_), .B(new_n1242_), .Y(new_n1244_));
  AND2X1   g00242(.A(\A[740] ), .B(\A[739] ), .Y(new_n1245_));
  AOI21X1  g00243(.A0(new_n1232_), .A1(\A[741] ), .B0(new_n1245_), .Y(new_n1246_));
  XOR2X1   g00244(.A(new_n1246_), .B(new_n1244_), .Y(new_n1247_));
  XOR2X1   g00245(.A(new_n1247_), .B(new_n1241_), .Y(new_n1248_));
  XOR2X1   g00246(.A(new_n1240_), .B(new_n1234_), .Y(new_n1249_));
  OR2X1    g00247(.A(new_n1240_), .B(new_n1234_), .Y(new_n1250_));
  AOI21X1  g00248(.A0(new_n1239_), .A1(\A[744] ), .B0(new_n1242_), .Y(new_n1251_));
  OR2X1    g00249(.A(new_n1246_), .B(new_n1251_), .Y(new_n1252_));
  OAI21X1  g00250(.A0(new_n1247_), .A1(new_n1250_), .B0(new_n1252_), .Y(new_n1253_));
  AND2X1   g00251(.A(new_n1253_), .B(new_n1249_), .Y(new_n1254_));
  OR2X1    g00252(.A(new_n1254_), .B(new_n1248_), .Y(new_n1255_));
  AND2X1   g00253(.A(\A[749] ), .B(\A[748] ), .Y(new_n1256_));
  XOR2X1   g00254(.A(\A[749] ), .B(\A[748] ), .Y(new_n1257_));
  AOI21X1  g00255(.A0(new_n1257_), .A1(\A[750] ), .B0(new_n1256_), .Y(new_n1258_));
  AND2X1   g00256(.A(\A[746] ), .B(\A[745] ), .Y(new_n1259_));
  XOR2X1   g00257(.A(\A[746] ), .B(\A[745] ), .Y(new_n1260_));
  AOI21X1  g00258(.A0(new_n1260_), .A1(\A[747] ), .B0(new_n1259_), .Y(new_n1261_));
  INVX1    g00259(.A(\A[746] ), .Y(new_n1262_));
  OR2X1    g00260(.A(new_n1262_), .B(\A[745] ), .Y(new_n1263_));
  INVX1    g00261(.A(\A[747] ), .Y(new_n1264_));
  AOI21X1  g00262(.A0(new_n1262_), .A1(\A[745] ), .B0(new_n1264_), .Y(new_n1265_));
  AND2X1   g00263(.A(new_n1260_), .B(new_n1264_), .Y(new_n1266_));
  AOI21X1  g00264(.A0(new_n1265_), .A1(new_n1263_), .B0(new_n1266_), .Y(new_n1267_));
  INVX1    g00265(.A(\A[750] ), .Y(new_n1268_));
  INVX1    g00266(.A(\A[749] ), .Y(new_n1269_));
  OR2X1    g00267(.A(new_n1269_), .B(\A[748] ), .Y(new_n1270_));
  AOI21X1  g00268(.A0(new_n1269_), .A1(\A[748] ), .B0(new_n1268_), .Y(new_n1271_));
  AOI22X1  g00269(.A0(new_n1271_), .A1(new_n1270_), .B0(new_n1257_), .B1(new_n1268_), .Y(new_n1272_));
  OR4X1    g00270(.A(new_n1272_), .B(new_n1267_), .C(new_n1261_), .D(new_n1258_), .Y(new_n1273_));
  OR4X1    g00271(.A(new_n1246_), .B(new_n1251_), .C(new_n1240_), .D(new_n1234_), .Y(new_n1274_));
  XOR2X1   g00272(.A(new_n1272_), .B(new_n1267_), .Y(new_n1275_));
  NAND4X1  g00273(.A(new_n1275_), .B(new_n1274_), .C(new_n1273_), .D(new_n1249_), .Y(new_n1276_));
  XOR2X1   g00274(.A(new_n1261_), .B(new_n1258_), .Y(new_n1277_));
  NOR2X1   g00275(.A(new_n1272_), .B(new_n1267_), .Y(new_n1278_));
  NOR2X1   g00276(.A(new_n1261_), .B(new_n1258_), .Y(new_n1279_));
  AOI21X1  g00277(.A0(new_n1278_), .A1(new_n1277_), .B0(new_n1279_), .Y(new_n1280_));
  XOR2X1   g00278(.A(new_n1278_), .B(new_n1277_), .Y(new_n1281_));
  AND2X1   g00279(.A(new_n1265_), .B(new_n1263_), .Y(new_n1282_));
  OR2X1    g00280(.A(new_n1266_), .B(new_n1282_), .Y(new_n1283_));
  XOR2X1   g00281(.A(new_n1272_), .B(new_n1283_), .Y(new_n1284_));
  OAI21X1  g00282(.A0(new_n1284_), .A1(new_n1280_), .B0(new_n1281_), .Y(new_n1285_));
  XOR2X1   g00283(.A(new_n1285_), .B(new_n1276_), .Y(new_n1286_));
  AND2X1   g00284(.A(new_n1286_), .B(new_n1255_), .Y(new_n1287_));
  AND2X1   g00285(.A(new_n1231_), .B(new_n1229_), .Y(new_n1288_));
  OR2X1    g00286(.A(new_n1233_), .B(new_n1288_), .Y(new_n1289_));
  XOR2X1   g00287(.A(new_n1240_), .B(new_n1289_), .Y(new_n1290_));
  OR2X1    g00288(.A(new_n1272_), .B(new_n1267_), .Y(new_n1291_));
  XOR2X1   g00289(.A(new_n1291_), .B(new_n1277_), .Y(new_n1292_));
  NOR4X1   g00290(.A(new_n1246_), .B(new_n1251_), .C(new_n1240_), .D(new_n1234_), .Y(new_n1293_));
  NOR4X1   g00291(.A(new_n1284_), .B(new_n1293_), .C(new_n1292_), .D(new_n1290_), .Y(new_n1294_));
  AND2X1   g00292(.A(new_n1278_), .B(new_n1277_), .Y(new_n1295_));
  OAI22X1  g00293(.A0(new_n1275_), .A1(new_n1281_), .B0(new_n1279_), .B1(new_n1295_), .Y(new_n1296_));
  AOI22X1  g00294(.A0(new_n1296_), .A1(new_n1294_), .B0(new_n1285_), .B1(new_n1276_), .Y(new_n1297_));
  NAND2X1  g00295(.A(new_n1275_), .B(new_n1273_), .Y(new_n1298_));
  XOR2X1   g00296(.A(new_n1240_), .B(new_n1234_), .Y(new_n1299_));
  XOR2X1   g00297(.A(new_n1299_), .B(new_n1298_), .Y(new_n1300_));
  NAND2X1  g00298(.A(new_n1205_), .B(new_n1203_), .Y(new_n1301_));
  XOR2X1   g00299(.A(new_n1171_), .B(new_n1165_), .Y(new_n1302_));
  XOR2X1   g00300(.A(new_n1302_), .B(new_n1301_), .Y(new_n1303_));
  NOR2X1   g00301(.A(new_n1303_), .B(new_n1300_), .Y(new_n1304_));
  OAI21X1  g00302(.A0(new_n1297_), .A1(new_n1255_), .B0(new_n1304_), .Y(new_n1305_));
  OR2X1    g00303(.A(new_n1305_), .B(new_n1287_), .Y(new_n1306_));
  NOR2X1   g00304(.A(new_n1297_), .B(new_n1255_), .Y(new_n1307_));
  OR2X1    g00305(.A(new_n1303_), .B(new_n1300_), .Y(new_n1308_));
  OAI21X1  g00306(.A0(new_n1307_), .A1(new_n1287_), .B0(new_n1308_), .Y(new_n1309_));
  AOI21X1  g00307(.A0(new_n1309_), .A1(new_n1306_), .B0(new_n1227_), .Y(new_n1310_));
  AND2X1   g00308(.A(new_n1184_), .B(new_n1179_), .Y(new_n1311_));
  AND2X1   g00309(.A(new_n1216_), .B(new_n1185_), .Y(new_n1312_));
  AOI21X1  g00310(.A0(new_n1226_), .A1(new_n1311_), .B0(new_n1312_), .Y(new_n1313_));
  OAI21X1  g00311(.A0(new_n1297_), .A1(new_n1255_), .B0(new_n1308_), .Y(new_n1314_));
  OR2X1    g00312(.A(new_n1314_), .B(new_n1287_), .Y(new_n1315_));
  OAI21X1  g00313(.A0(new_n1307_), .A1(new_n1287_), .B0(new_n1304_), .Y(new_n1316_));
  AOI21X1  g00314(.A0(new_n1316_), .A1(new_n1315_), .B0(new_n1313_), .Y(new_n1317_));
  XOR2X1   g00315(.A(new_n1303_), .B(new_n1300_), .Y(new_n1318_));
  INVX1    g00316(.A(new_n1318_), .Y(new_n1319_));
  INVX1    g00317(.A(new_n1113_), .Y(new_n1320_));
  XOR2X1   g00318(.A(new_n1320_), .B(new_n1075_), .Y(new_n1321_));
  OR2X1    g00319(.A(new_n1321_), .B(new_n1319_), .Y(new_n1322_));
  NOR3X1   g00320(.A(new_n1322_), .B(new_n1317_), .C(new_n1310_), .Y(new_n1323_));
  NOR2X1   g00321(.A(new_n1305_), .B(new_n1287_), .Y(new_n1324_));
  NAND2X1  g00322(.A(new_n1286_), .B(new_n1255_), .Y(new_n1325_));
  OR2X1    g00323(.A(new_n1297_), .B(new_n1255_), .Y(new_n1326_));
  AOI21X1  g00324(.A0(new_n1326_), .A1(new_n1325_), .B0(new_n1304_), .Y(new_n1327_));
  OAI21X1  g00325(.A0(new_n1327_), .A1(new_n1324_), .B0(new_n1313_), .Y(new_n1328_));
  NOR2X1   g00326(.A(new_n1314_), .B(new_n1287_), .Y(new_n1329_));
  AOI21X1  g00327(.A0(new_n1326_), .A1(new_n1325_), .B0(new_n1308_), .Y(new_n1330_));
  OAI21X1  g00328(.A0(new_n1330_), .A1(new_n1329_), .B0(new_n1227_), .Y(new_n1331_));
  NOR2X1   g00329(.A(new_n1321_), .B(new_n1319_), .Y(new_n1332_));
  AOI21X1  g00330(.A0(new_n1331_), .A1(new_n1328_), .B0(new_n1332_), .Y(new_n1333_));
  OAI21X1  g00331(.A0(new_n1333_), .A1(new_n1323_), .B0(new_n1158_), .Y(new_n1334_));
  NAND2X1  g00332(.A(new_n1156_), .B(new_n1155_), .Y(new_n1335_));
  MX2X1    g00333(.A(new_n1335_), .B(new_n1119_), .S0(new_n1152_), .Y(new_n1336_));
  NOR3X1   g00334(.A(new_n1332_), .B(new_n1317_), .C(new_n1310_), .Y(new_n1337_));
  AOI21X1  g00335(.A0(new_n1331_), .A1(new_n1328_), .B0(new_n1322_), .Y(new_n1338_));
  OAI21X1  g00336(.A0(new_n1338_), .A1(new_n1337_), .B0(new_n1336_), .Y(new_n1339_));
  XOR2X1   g00337(.A(new_n1321_), .B(new_n1318_), .Y(new_n1340_));
  INVX1    g00338(.A(\A[697] ), .Y(new_n1341_));
  OR2X1    g00339(.A(\A[698] ), .B(new_n1341_), .Y(new_n1342_));
  INVX1    g00340(.A(\A[699] ), .Y(new_n1343_));
  AOI21X1  g00341(.A0(\A[698] ), .A1(new_n1341_), .B0(new_n1343_), .Y(new_n1344_));
  XOR2X1   g00342(.A(\A[698] ), .B(\A[697] ), .Y(new_n1345_));
  AND2X1   g00343(.A(new_n1345_), .B(new_n1343_), .Y(new_n1346_));
  AOI21X1  g00344(.A0(new_n1344_), .A1(new_n1342_), .B0(new_n1346_), .Y(new_n1347_));
  INVX1    g00345(.A(\A[702] ), .Y(new_n1348_));
  INVX1    g00346(.A(\A[700] ), .Y(new_n1349_));
  OR2X1    g00347(.A(\A[701] ), .B(new_n1349_), .Y(new_n1350_));
  AOI21X1  g00348(.A0(\A[701] ), .A1(new_n1349_), .B0(new_n1348_), .Y(new_n1351_));
  XOR2X1   g00349(.A(\A[701] ), .B(\A[700] ), .Y(new_n1352_));
  AOI22X1  g00350(.A0(new_n1352_), .A1(new_n1348_), .B0(new_n1351_), .B1(new_n1350_), .Y(new_n1353_));
  AND2X1   g00351(.A(\A[701] ), .B(\A[700] ), .Y(new_n1354_));
  AOI21X1  g00352(.A0(new_n1352_), .A1(\A[702] ), .B0(new_n1354_), .Y(new_n1355_));
  AND2X1   g00353(.A(\A[698] ), .B(\A[697] ), .Y(new_n1356_));
  AOI21X1  g00354(.A0(new_n1345_), .A1(\A[699] ), .B0(new_n1356_), .Y(new_n1357_));
  XOR2X1   g00355(.A(new_n1353_), .B(new_n1347_), .Y(new_n1358_));
  INVX1    g00356(.A(\A[691] ), .Y(new_n1359_));
  OR2X1    g00357(.A(\A[692] ), .B(new_n1359_), .Y(new_n1360_));
  INVX1    g00358(.A(\A[693] ), .Y(new_n1361_));
  AOI21X1  g00359(.A0(\A[692] ), .A1(new_n1359_), .B0(new_n1361_), .Y(new_n1362_));
  XOR2X1   g00360(.A(\A[692] ), .B(\A[691] ), .Y(new_n1363_));
  AND2X1   g00361(.A(new_n1363_), .B(new_n1361_), .Y(new_n1364_));
  AOI21X1  g00362(.A0(new_n1362_), .A1(new_n1360_), .B0(new_n1364_), .Y(new_n1365_));
  INVX1    g00363(.A(\A[696] ), .Y(new_n1366_));
  INVX1    g00364(.A(\A[694] ), .Y(new_n1367_));
  OR2X1    g00365(.A(\A[695] ), .B(new_n1367_), .Y(new_n1368_));
  AOI21X1  g00366(.A0(\A[695] ), .A1(new_n1367_), .B0(new_n1366_), .Y(new_n1369_));
  XOR2X1   g00367(.A(\A[695] ), .B(\A[694] ), .Y(new_n1370_));
  AOI22X1  g00368(.A0(new_n1370_), .A1(new_n1366_), .B0(new_n1369_), .B1(new_n1368_), .Y(new_n1371_));
  AND2X1   g00369(.A(\A[695] ), .B(\A[694] ), .Y(new_n1372_));
  AOI21X1  g00370(.A0(new_n1370_), .A1(\A[696] ), .B0(new_n1372_), .Y(new_n1373_));
  AND2X1   g00371(.A(\A[692] ), .B(\A[691] ), .Y(new_n1374_));
  AOI21X1  g00372(.A0(new_n1363_), .A1(\A[693] ), .B0(new_n1374_), .Y(new_n1375_));
  XOR2X1   g00373(.A(new_n1371_), .B(new_n1365_), .Y(new_n1376_));
  XOR2X1   g00374(.A(new_n1376_), .B(new_n1358_), .Y(new_n1377_));
  INVX1    g00375(.A(\A[685] ), .Y(new_n1378_));
  OR2X1    g00376(.A(\A[686] ), .B(new_n1378_), .Y(new_n1379_));
  INVX1    g00377(.A(\A[687] ), .Y(new_n1380_));
  AOI21X1  g00378(.A0(\A[686] ), .A1(new_n1378_), .B0(new_n1380_), .Y(new_n1381_));
  AND2X1   g00379(.A(new_n1381_), .B(new_n1379_), .Y(new_n1382_));
  XOR2X1   g00380(.A(\A[686] ), .B(\A[685] ), .Y(new_n1383_));
  AND2X1   g00381(.A(new_n1383_), .B(new_n1380_), .Y(new_n1384_));
  OR2X1    g00382(.A(new_n1384_), .B(new_n1382_), .Y(new_n1385_));
  INVX1    g00383(.A(\A[690] ), .Y(new_n1386_));
  INVX1    g00384(.A(\A[688] ), .Y(new_n1387_));
  OR2X1    g00385(.A(\A[689] ), .B(new_n1387_), .Y(new_n1388_));
  AOI21X1  g00386(.A0(\A[689] ), .A1(new_n1387_), .B0(new_n1386_), .Y(new_n1389_));
  XOR2X1   g00387(.A(\A[689] ), .B(\A[688] ), .Y(new_n1390_));
  AOI22X1  g00388(.A0(new_n1390_), .A1(new_n1386_), .B0(new_n1389_), .B1(new_n1388_), .Y(new_n1391_));
  AND2X1   g00389(.A(\A[689] ), .B(\A[688] ), .Y(new_n1392_));
  AOI21X1  g00390(.A0(new_n1390_), .A1(\A[690] ), .B0(new_n1392_), .Y(new_n1393_));
  AND2X1   g00391(.A(\A[686] ), .B(\A[685] ), .Y(new_n1394_));
  AOI21X1  g00392(.A0(new_n1383_), .A1(\A[687] ), .B0(new_n1394_), .Y(new_n1395_));
  XOR2X1   g00393(.A(new_n1391_), .B(new_n1385_), .Y(new_n1396_));
  INVX1    g00394(.A(\A[679] ), .Y(new_n1397_));
  OR2X1    g00395(.A(\A[680] ), .B(new_n1397_), .Y(new_n1398_));
  INVX1    g00396(.A(\A[681] ), .Y(new_n1399_));
  AOI21X1  g00397(.A0(\A[680] ), .A1(new_n1397_), .B0(new_n1399_), .Y(new_n1400_));
  XOR2X1   g00398(.A(\A[680] ), .B(\A[679] ), .Y(new_n1401_));
  AND2X1   g00399(.A(new_n1401_), .B(new_n1399_), .Y(new_n1402_));
  AOI21X1  g00400(.A0(new_n1400_), .A1(new_n1398_), .B0(new_n1402_), .Y(new_n1403_));
  INVX1    g00401(.A(\A[684] ), .Y(new_n1404_));
  INVX1    g00402(.A(\A[682] ), .Y(new_n1405_));
  OR2X1    g00403(.A(\A[683] ), .B(new_n1405_), .Y(new_n1406_));
  AOI21X1  g00404(.A0(\A[683] ), .A1(new_n1405_), .B0(new_n1404_), .Y(new_n1407_));
  XOR2X1   g00405(.A(\A[683] ), .B(\A[682] ), .Y(new_n1408_));
  AOI22X1  g00406(.A0(new_n1408_), .A1(new_n1404_), .B0(new_n1407_), .B1(new_n1406_), .Y(new_n1409_));
  AND2X1   g00407(.A(\A[683] ), .B(\A[682] ), .Y(new_n1410_));
  AOI21X1  g00408(.A0(new_n1408_), .A1(\A[684] ), .B0(new_n1410_), .Y(new_n1411_));
  AND2X1   g00409(.A(\A[680] ), .B(\A[679] ), .Y(new_n1412_));
  AOI21X1  g00410(.A0(new_n1401_), .A1(\A[681] ), .B0(new_n1412_), .Y(new_n1413_));
  XOR2X1   g00411(.A(new_n1409_), .B(new_n1403_), .Y(new_n1414_));
  XOR2X1   g00412(.A(new_n1414_), .B(new_n1396_), .Y(new_n1415_));
  XOR2X1   g00413(.A(new_n1415_), .B(new_n1377_), .Y(new_n1416_));
  INVX1    g00414(.A(\A[673] ), .Y(new_n1417_));
  OR2X1    g00415(.A(\A[674] ), .B(new_n1417_), .Y(new_n1418_));
  INVX1    g00416(.A(\A[675] ), .Y(new_n1419_));
  AOI21X1  g00417(.A0(\A[674] ), .A1(new_n1417_), .B0(new_n1419_), .Y(new_n1420_));
  XOR2X1   g00418(.A(\A[674] ), .B(\A[673] ), .Y(new_n1421_));
  AND2X1   g00419(.A(new_n1421_), .B(new_n1419_), .Y(new_n1422_));
  AOI21X1  g00420(.A0(new_n1420_), .A1(new_n1418_), .B0(new_n1422_), .Y(new_n1423_));
  INVX1    g00421(.A(\A[678] ), .Y(new_n1424_));
  INVX1    g00422(.A(\A[676] ), .Y(new_n1425_));
  OR2X1    g00423(.A(\A[677] ), .B(new_n1425_), .Y(new_n1426_));
  AOI21X1  g00424(.A0(\A[677] ), .A1(new_n1425_), .B0(new_n1424_), .Y(new_n1427_));
  XOR2X1   g00425(.A(\A[677] ), .B(\A[676] ), .Y(new_n1428_));
  AOI22X1  g00426(.A0(new_n1428_), .A1(new_n1424_), .B0(new_n1427_), .B1(new_n1426_), .Y(new_n1429_));
  AND2X1   g00427(.A(\A[677] ), .B(\A[676] ), .Y(new_n1430_));
  AOI21X1  g00428(.A0(new_n1428_), .A1(\A[678] ), .B0(new_n1430_), .Y(new_n1431_));
  AND2X1   g00429(.A(\A[674] ), .B(\A[673] ), .Y(new_n1432_));
  AOI21X1  g00430(.A0(new_n1421_), .A1(\A[675] ), .B0(new_n1432_), .Y(new_n1433_));
  XOR2X1   g00431(.A(new_n1429_), .B(new_n1423_), .Y(new_n1434_));
  INVX1    g00432(.A(\A[667] ), .Y(new_n1435_));
  OR2X1    g00433(.A(\A[668] ), .B(new_n1435_), .Y(new_n1436_));
  INVX1    g00434(.A(\A[669] ), .Y(new_n1437_));
  AOI21X1  g00435(.A0(\A[668] ), .A1(new_n1435_), .B0(new_n1437_), .Y(new_n1438_));
  XOR2X1   g00436(.A(\A[668] ), .B(\A[667] ), .Y(new_n1439_));
  AND2X1   g00437(.A(new_n1439_), .B(new_n1437_), .Y(new_n1440_));
  AOI21X1  g00438(.A0(new_n1438_), .A1(new_n1436_), .B0(new_n1440_), .Y(new_n1441_));
  INVX1    g00439(.A(\A[672] ), .Y(new_n1442_));
  INVX1    g00440(.A(\A[670] ), .Y(new_n1443_));
  OR2X1    g00441(.A(\A[671] ), .B(new_n1443_), .Y(new_n1444_));
  AOI21X1  g00442(.A0(\A[671] ), .A1(new_n1443_), .B0(new_n1442_), .Y(new_n1445_));
  XOR2X1   g00443(.A(\A[671] ), .B(\A[670] ), .Y(new_n1446_));
  AOI22X1  g00444(.A0(new_n1446_), .A1(new_n1442_), .B0(new_n1445_), .B1(new_n1444_), .Y(new_n1447_));
  AND2X1   g00445(.A(\A[671] ), .B(\A[670] ), .Y(new_n1448_));
  AOI21X1  g00446(.A0(new_n1446_), .A1(\A[672] ), .B0(new_n1448_), .Y(new_n1449_));
  AND2X1   g00447(.A(\A[668] ), .B(\A[667] ), .Y(new_n1450_));
  AOI21X1  g00448(.A0(new_n1439_), .A1(\A[669] ), .B0(new_n1450_), .Y(new_n1451_));
  XOR2X1   g00449(.A(new_n1447_), .B(new_n1441_), .Y(new_n1452_));
  XOR2X1   g00450(.A(new_n1452_), .B(new_n1434_), .Y(new_n1453_));
  INVX1    g00451(.A(new_n1453_), .Y(new_n1454_));
  INVX1    g00452(.A(\A[661] ), .Y(new_n1455_));
  OR2X1    g00453(.A(\A[662] ), .B(new_n1455_), .Y(new_n1456_));
  INVX1    g00454(.A(\A[663] ), .Y(new_n1457_));
  AOI21X1  g00455(.A0(\A[662] ), .A1(new_n1455_), .B0(new_n1457_), .Y(new_n1458_));
  AND2X1   g00456(.A(new_n1458_), .B(new_n1456_), .Y(new_n1459_));
  XOR2X1   g00457(.A(\A[662] ), .B(\A[661] ), .Y(new_n1460_));
  AND2X1   g00458(.A(new_n1460_), .B(new_n1457_), .Y(new_n1461_));
  OR2X1    g00459(.A(new_n1461_), .B(new_n1459_), .Y(new_n1462_));
  INVX1    g00460(.A(\A[666] ), .Y(new_n1463_));
  INVX1    g00461(.A(\A[664] ), .Y(new_n1464_));
  OR2X1    g00462(.A(\A[665] ), .B(new_n1464_), .Y(new_n1465_));
  AOI21X1  g00463(.A0(\A[665] ), .A1(new_n1464_), .B0(new_n1463_), .Y(new_n1466_));
  XOR2X1   g00464(.A(\A[665] ), .B(\A[664] ), .Y(new_n1467_));
  AOI22X1  g00465(.A0(new_n1467_), .A1(new_n1463_), .B0(new_n1466_), .B1(new_n1465_), .Y(new_n1468_));
  AND2X1   g00466(.A(\A[665] ), .B(\A[664] ), .Y(new_n1469_));
  AOI21X1  g00467(.A0(new_n1467_), .A1(\A[666] ), .B0(new_n1469_), .Y(new_n1470_));
  AND2X1   g00468(.A(\A[662] ), .B(\A[661] ), .Y(new_n1471_));
  AOI21X1  g00469(.A0(new_n1460_), .A1(\A[663] ), .B0(new_n1471_), .Y(new_n1472_));
  XOR2X1   g00470(.A(new_n1468_), .B(new_n1462_), .Y(new_n1473_));
  INVX1    g00471(.A(\A[655] ), .Y(new_n1474_));
  OR2X1    g00472(.A(\A[656] ), .B(new_n1474_), .Y(new_n1475_));
  INVX1    g00473(.A(\A[657] ), .Y(new_n1476_));
  AOI21X1  g00474(.A0(\A[656] ), .A1(new_n1474_), .B0(new_n1476_), .Y(new_n1477_));
  XOR2X1   g00475(.A(\A[656] ), .B(\A[655] ), .Y(new_n1478_));
  AND2X1   g00476(.A(new_n1478_), .B(new_n1476_), .Y(new_n1479_));
  AOI21X1  g00477(.A0(new_n1477_), .A1(new_n1475_), .B0(new_n1479_), .Y(new_n1480_));
  INVX1    g00478(.A(\A[660] ), .Y(new_n1481_));
  INVX1    g00479(.A(\A[658] ), .Y(new_n1482_));
  OR2X1    g00480(.A(\A[659] ), .B(new_n1482_), .Y(new_n1483_));
  AOI21X1  g00481(.A0(\A[659] ), .A1(new_n1482_), .B0(new_n1481_), .Y(new_n1484_));
  XOR2X1   g00482(.A(\A[659] ), .B(\A[658] ), .Y(new_n1485_));
  AOI22X1  g00483(.A0(new_n1485_), .A1(new_n1481_), .B0(new_n1484_), .B1(new_n1483_), .Y(new_n1486_));
  AND2X1   g00484(.A(\A[659] ), .B(\A[658] ), .Y(new_n1487_));
  AOI21X1  g00485(.A0(new_n1485_), .A1(\A[660] ), .B0(new_n1487_), .Y(new_n1488_));
  AND2X1   g00486(.A(\A[656] ), .B(\A[655] ), .Y(new_n1489_));
  AOI21X1  g00487(.A0(new_n1478_), .A1(\A[657] ), .B0(new_n1489_), .Y(new_n1490_));
  XOR2X1   g00488(.A(new_n1486_), .B(new_n1480_), .Y(new_n1491_));
  XOR2X1   g00489(.A(new_n1491_), .B(new_n1473_), .Y(new_n1492_));
  XOR2X1   g00490(.A(new_n1492_), .B(new_n1454_), .Y(new_n1493_));
  XOR2X1   g00491(.A(new_n1493_), .B(new_n1416_), .Y(new_n1494_));
  NOR2X1   g00492(.A(new_n1494_), .B(new_n1340_), .Y(new_n1495_));
  NAND3X1  g00493(.A(new_n1495_), .B(new_n1339_), .C(new_n1334_), .Y(new_n1496_));
  NAND3X1  g00494(.A(new_n1332_), .B(new_n1331_), .C(new_n1328_), .Y(new_n1497_));
  OAI21X1  g00495(.A0(new_n1317_), .A1(new_n1310_), .B0(new_n1322_), .Y(new_n1498_));
  AOI21X1  g00496(.A0(new_n1498_), .A1(new_n1497_), .B0(new_n1336_), .Y(new_n1499_));
  NAND3X1  g00497(.A(new_n1322_), .B(new_n1331_), .C(new_n1328_), .Y(new_n1500_));
  OAI21X1  g00498(.A0(new_n1317_), .A1(new_n1310_), .B0(new_n1332_), .Y(new_n1501_));
  AOI21X1  g00499(.A0(new_n1501_), .A1(new_n1500_), .B0(new_n1158_), .Y(new_n1502_));
  INVX1    g00500(.A(new_n1495_), .Y(new_n1503_));
  OAI21X1  g00501(.A0(new_n1502_), .A1(new_n1499_), .B0(new_n1503_), .Y(new_n1504_));
  AND2X1   g00502(.A(new_n1504_), .B(new_n1496_), .Y(new_n1505_));
  AND2X1   g00503(.A(new_n1400_), .B(new_n1398_), .Y(new_n1506_));
  OR2X1    g00504(.A(new_n1402_), .B(new_n1506_), .Y(new_n1507_));
  XOR2X1   g00505(.A(new_n1409_), .B(new_n1507_), .Y(new_n1508_));
  XOR2X1   g00506(.A(new_n1413_), .B(new_n1411_), .Y(new_n1509_));
  NOR2X1   g00507(.A(new_n1409_), .B(new_n1403_), .Y(new_n1510_));
  NOR2X1   g00508(.A(new_n1413_), .B(new_n1411_), .Y(new_n1511_));
  AOI21X1  g00509(.A0(new_n1510_), .A1(new_n1509_), .B0(new_n1511_), .Y(new_n1512_));
  XOR2X1   g00510(.A(new_n1510_), .B(new_n1509_), .Y(new_n1513_));
  OAI21X1  g00511(.A0(new_n1512_), .A1(new_n1508_), .B0(new_n1513_), .Y(new_n1514_));
  INVX1    g00512(.A(new_n1514_), .Y(new_n1515_));
  XOR2X1   g00513(.A(new_n1391_), .B(new_n1385_), .Y(new_n1516_));
  AOI21X1  g00514(.A0(new_n1381_), .A1(new_n1379_), .B0(new_n1384_), .Y(new_n1517_));
  NOR4X1   g00515(.A(new_n1395_), .B(new_n1393_), .C(new_n1391_), .D(new_n1517_), .Y(new_n1518_));
  NOR4X1   g00516(.A(new_n1413_), .B(new_n1411_), .C(new_n1409_), .D(new_n1403_), .Y(new_n1519_));
  OR4X1    g00517(.A(new_n1519_), .B(new_n1508_), .C(new_n1518_), .D(new_n1516_), .Y(new_n1520_));
  XOR2X1   g00518(.A(new_n1395_), .B(new_n1393_), .Y(new_n1521_));
  NOR2X1   g00519(.A(new_n1391_), .B(new_n1517_), .Y(new_n1522_));
  NOR2X1   g00520(.A(new_n1395_), .B(new_n1393_), .Y(new_n1523_));
  AOI21X1  g00521(.A0(new_n1522_), .A1(new_n1521_), .B0(new_n1523_), .Y(new_n1524_));
  XOR2X1   g00522(.A(new_n1522_), .B(new_n1521_), .Y(new_n1525_));
  OAI21X1  g00523(.A0(new_n1524_), .A1(new_n1516_), .B0(new_n1525_), .Y(new_n1526_));
  XOR2X1   g00524(.A(new_n1526_), .B(new_n1520_), .Y(new_n1527_));
  AND2X1   g00525(.A(new_n1527_), .B(new_n1514_), .Y(new_n1528_));
  AND2X1   g00526(.A(new_n1526_), .B(new_n1520_), .Y(new_n1529_));
  OR2X1    g00527(.A(new_n1391_), .B(new_n1517_), .Y(new_n1530_));
  XOR2X1   g00528(.A(new_n1530_), .B(new_n1521_), .Y(new_n1531_));
  OR4X1    g00529(.A(new_n1508_), .B(new_n1518_), .C(new_n1531_), .D(new_n1516_), .Y(new_n1532_));
  OR4X1    g00530(.A(new_n1413_), .B(new_n1411_), .C(new_n1409_), .D(new_n1403_), .Y(new_n1533_));
  OAI21X1  g00531(.A0(new_n1524_), .A1(new_n1516_), .B0(new_n1533_), .Y(new_n1534_));
  NOR2X1   g00532(.A(new_n1534_), .B(new_n1532_), .Y(new_n1535_));
  OR2X1    g00533(.A(new_n1535_), .B(new_n1529_), .Y(new_n1536_));
  AOI21X1  g00534(.A0(new_n1536_), .A1(new_n1515_), .B0(new_n1528_), .Y(new_n1537_));
  AND2X1   g00535(.A(new_n1362_), .B(new_n1360_), .Y(new_n1538_));
  OR2X1    g00536(.A(new_n1364_), .B(new_n1538_), .Y(new_n1539_));
  XOR2X1   g00537(.A(new_n1371_), .B(new_n1539_), .Y(new_n1540_));
  XOR2X1   g00538(.A(new_n1375_), .B(new_n1373_), .Y(new_n1541_));
  NOR2X1   g00539(.A(new_n1371_), .B(new_n1365_), .Y(new_n1542_));
  NOR2X1   g00540(.A(new_n1375_), .B(new_n1373_), .Y(new_n1543_));
  AOI21X1  g00541(.A0(new_n1542_), .A1(new_n1541_), .B0(new_n1543_), .Y(new_n1544_));
  XOR2X1   g00542(.A(new_n1542_), .B(new_n1541_), .Y(new_n1545_));
  OAI21X1  g00543(.A0(new_n1544_), .A1(new_n1540_), .B0(new_n1545_), .Y(new_n1546_));
  AND2X1   g00544(.A(new_n1344_), .B(new_n1342_), .Y(new_n1547_));
  OR2X1    g00545(.A(new_n1346_), .B(new_n1547_), .Y(new_n1548_));
  XOR2X1   g00546(.A(new_n1353_), .B(new_n1548_), .Y(new_n1549_));
  NOR4X1   g00547(.A(new_n1357_), .B(new_n1355_), .C(new_n1353_), .D(new_n1347_), .Y(new_n1550_));
  NOR4X1   g00548(.A(new_n1375_), .B(new_n1373_), .C(new_n1371_), .D(new_n1365_), .Y(new_n1551_));
  OR4X1    g00549(.A(new_n1551_), .B(new_n1540_), .C(new_n1550_), .D(new_n1549_), .Y(new_n1552_));
  XOR2X1   g00550(.A(new_n1357_), .B(new_n1355_), .Y(new_n1553_));
  NOR2X1   g00551(.A(new_n1353_), .B(new_n1347_), .Y(new_n1554_));
  NOR2X1   g00552(.A(new_n1357_), .B(new_n1355_), .Y(new_n1555_));
  AOI21X1  g00553(.A0(new_n1554_), .A1(new_n1553_), .B0(new_n1555_), .Y(new_n1556_));
  XOR2X1   g00554(.A(new_n1554_), .B(new_n1553_), .Y(new_n1557_));
  OAI21X1  g00555(.A0(new_n1556_), .A1(new_n1549_), .B0(new_n1557_), .Y(new_n1558_));
  XOR2X1   g00556(.A(new_n1558_), .B(new_n1552_), .Y(new_n1559_));
  AND2X1   g00557(.A(new_n1559_), .B(new_n1546_), .Y(new_n1560_));
  NAND2X1  g00558(.A(new_n1558_), .B(new_n1552_), .Y(new_n1561_));
  OR2X1    g00559(.A(new_n1353_), .B(new_n1347_), .Y(new_n1562_));
  XOR2X1   g00560(.A(new_n1562_), .B(new_n1553_), .Y(new_n1563_));
  OR4X1    g00561(.A(new_n1540_), .B(new_n1550_), .C(new_n1563_), .D(new_n1549_), .Y(new_n1564_));
  AND2X1   g00562(.A(new_n1370_), .B(\A[696] ), .Y(new_n1565_));
  OR2X1    g00563(.A(new_n1565_), .B(new_n1372_), .Y(new_n1566_));
  XOR2X1   g00564(.A(new_n1375_), .B(new_n1566_), .Y(new_n1567_));
  XOR2X1   g00565(.A(new_n1542_), .B(new_n1567_), .Y(new_n1568_));
  OAI22X1  g00566(.A0(new_n1568_), .A1(new_n1544_), .B0(new_n1556_), .B1(new_n1549_), .Y(new_n1569_));
  OR2X1    g00567(.A(new_n1569_), .B(new_n1564_), .Y(new_n1570_));
  AOI21X1  g00568(.A0(new_n1570_), .A1(new_n1561_), .B0(new_n1546_), .Y(new_n1571_));
  INVX1    g00569(.A(new_n1377_), .Y(new_n1572_));
  OR2X1    g00570(.A(new_n1415_), .B(new_n1572_), .Y(new_n1573_));
  NOR3X1   g00571(.A(new_n1573_), .B(new_n1571_), .C(new_n1560_), .Y(new_n1574_));
  NAND2X1  g00572(.A(new_n1559_), .B(new_n1546_), .Y(new_n1575_));
  XOR2X1   g00573(.A(new_n1371_), .B(new_n1365_), .Y(new_n1576_));
  OR2X1    g00574(.A(new_n1371_), .B(new_n1365_), .Y(new_n1577_));
  OR2X1    g00575(.A(new_n1375_), .B(new_n1373_), .Y(new_n1578_));
  OAI21X1  g00576(.A0(new_n1577_), .A1(new_n1567_), .B0(new_n1578_), .Y(new_n1579_));
  AOI21X1  g00577(.A0(new_n1579_), .A1(new_n1576_), .B0(new_n1568_), .Y(new_n1580_));
  AND2X1   g00578(.A(new_n1558_), .B(new_n1552_), .Y(new_n1581_));
  NOR2X1   g00579(.A(new_n1569_), .B(new_n1564_), .Y(new_n1582_));
  OAI21X1  g00580(.A0(new_n1582_), .A1(new_n1581_), .B0(new_n1580_), .Y(new_n1583_));
  NOR2X1   g00581(.A(new_n1415_), .B(new_n1572_), .Y(new_n1584_));
  AOI21X1  g00582(.A0(new_n1583_), .A1(new_n1575_), .B0(new_n1584_), .Y(new_n1585_));
  OAI21X1  g00583(.A0(new_n1585_), .A1(new_n1574_), .B0(new_n1537_), .Y(new_n1586_));
  MX2X1    g00584(.A(new_n1536_), .B(new_n1527_), .S0(new_n1514_), .Y(new_n1587_));
  NOR3X1   g00585(.A(new_n1584_), .B(new_n1571_), .C(new_n1560_), .Y(new_n1588_));
  AOI21X1  g00586(.A0(new_n1583_), .A1(new_n1575_), .B0(new_n1573_), .Y(new_n1589_));
  OAI21X1  g00587(.A0(new_n1589_), .A1(new_n1588_), .B0(new_n1587_), .Y(new_n1590_));
  XOR2X1   g00588(.A(new_n1492_), .B(new_n1453_), .Y(new_n1591_));
  NOR2X1   g00589(.A(new_n1591_), .B(new_n1416_), .Y(new_n1592_));
  NAND3X1  g00590(.A(new_n1592_), .B(new_n1590_), .C(new_n1586_), .Y(new_n1593_));
  NAND3X1  g00591(.A(new_n1584_), .B(new_n1583_), .C(new_n1575_), .Y(new_n1594_));
  OAI21X1  g00592(.A0(new_n1571_), .A1(new_n1560_), .B0(new_n1573_), .Y(new_n1595_));
  AOI21X1  g00593(.A0(new_n1595_), .A1(new_n1594_), .B0(new_n1587_), .Y(new_n1596_));
  NAND3X1  g00594(.A(new_n1573_), .B(new_n1583_), .C(new_n1575_), .Y(new_n1597_));
  OAI21X1  g00595(.A0(new_n1571_), .A1(new_n1560_), .B0(new_n1584_), .Y(new_n1598_));
  AOI21X1  g00596(.A0(new_n1598_), .A1(new_n1597_), .B0(new_n1537_), .Y(new_n1599_));
  INVX1    g00597(.A(new_n1592_), .Y(new_n1600_));
  OAI21X1  g00598(.A0(new_n1599_), .A1(new_n1596_), .B0(new_n1600_), .Y(new_n1601_));
  AND2X1   g00599(.A(new_n1601_), .B(new_n1593_), .Y(new_n1602_));
  AND2X1   g00600(.A(new_n1438_), .B(new_n1436_), .Y(new_n1603_));
  OR2X1    g00601(.A(new_n1440_), .B(new_n1603_), .Y(new_n1604_));
  XOR2X1   g00602(.A(new_n1447_), .B(new_n1604_), .Y(new_n1605_));
  XOR2X1   g00603(.A(new_n1451_), .B(new_n1449_), .Y(new_n1606_));
  NOR2X1   g00604(.A(new_n1447_), .B(new_n1441_), .Y(new_n1607_));
  NOR2X1   g00605(.A(new_n1451_), .B(new_n1449_), .Y(new_n1608_));
  AOI21X1  g00606(.A0(new_n1607_), .A1(new_n1606_), .B0(new_n1608_), .Y(new_n1609_));
  XOR2X1   g00607(.A(new_n1607_), .B(new_n1606_), .Y(new_n1610_));
  OAI21X1  g00608(.A0(new_n1609_), .A1(new_n1605_), .B0(new_n1610_), .Y(new_n1611_));
  AND2X1   g00609(.A(new_n1420_), .B(new_n1418_), .Y(new_n1612_));
  OR2X1    g00610(.A(new_n1422_), .B(new_n1612_), .Y(new_n1613_));
  XOR2X1   g00611(.A(new_n1429_), .B(new_n1613_), .Y(new_n1614_));
  NOR4X1   g00612(.A(new_n1433_), .B(new_n1431_), .C(new_n1429_), .D(new_n1423_), .Y(new_n1615_));
  NOR4X1   g00613(.A(new_n1451_), .B(new_n1449_), .C(new_n1447_), .D(new_n1441_), .Y(new_n1616_));
  OR4X1    g00614(.A(new_n1616_), .B(new_n1605_), .C(new_n1615_), .D(new_n1614_), .Y(new_n1617_));
  XOR2X1   g00615(.A(new_n1433_), .B(new_n1431_), .Y(new_n1618_));
  NOR2X1   g00616(.A(new_n1429_), .B(new_n1423_), .Y(new_n1619_));
  NOR2X1   g00617(.A(new_n1433_), .B(new_n1431_), .Y(new_n1620_));
  AOI21X1  g00618(.A0(new_n1619_), .A1(new_n1618_), .B0(new_n1620_), .Y(new_n1621_));
  XOR2X1   g00619(.A(new_n1619_), .B(new_n1618_), .Y(new_n1622_));
  OAI21X1  g00620(.A0(new_n1621_), .A1(new_n1614_), .B0(new_n1622_), .Y(new_n1623_));
  XOR2X1   g00621(.A(new_n1623_), .B(new_n1617_), .Y(new_n1624_));
  NAND2X1  g00622(.A(new_n1624_), .B(new_n1611_), .Y(new_n1625_));
  XOR2X1   g00623(.A(new_n1447_), .B(new_n1441_), .Y(new_n1626_));
  AND2X1   g00624(.A(new_n1446_), .B(\A[672] ), .Y(new_n1627_));
  OR2X1    g00625(.A(new_n1627_), .B(new_n1448_), .Y(new_n1628_));
  XOR2X1   g00626(.A(new_n1451_), .B(new_n1628_), .Y(new_n1629_));
  OR2X1    g00627(.A(new_n1447_), .B(new_n1441_), .Y(new_n1630_));
  OR2X1    g00628(.A(new_n1451_), .B(new_n1449_), .Y(new_n1631_));
  OAI21X1  g00629(.A0(new_n1630_), .A1(new_n1629_), .B0(new_n1631_), .Y(new_n1632_));
  XOR2X1   g00630(.A(new_n1607_), .B(new_n1629_), .Y(new_n1633_));
  AOI21X1  g00631(.A0(new_n1632_), .A1(new_n1626_), .B0(new_n1633_), .Y(new_n1634_));
  AND2X1   g00632(.A(new_n1623_), .B(new_n1617_), .Y(new_n1635_));
  OR2X1    g00633(.A(new_n1429_), .B(new_n1423_), .Y(new_n1636_));
  XOR2X1   g00634(.A(new_n1636_), .B(new_n1618_), .Y(new_n1637_));
  OR4X1    g00635(.A(new_n1605_), .B(new_n1615_), .C(new_n1637_), .D(new_n1614_), .Y(new_n1638_));
  OAI22X1  g00636(.A0(new_n1633_), .A1(new_n1609_), .B0(new_n1621_), .B1(new_n1614_), .Y(new_n1639_));
  NOR2X1   g00637(.A(new_n1639_), .B(new_n1638_), .Y(new_n1640_));
  OAI21X1  g00638(.A0(new_n1640_), .A1(new_n1635_), .B0(new_n1634_), .Y(new_n1641_));
  NOR2X1   g00639(.A(new_n1492_), .B(new_n1454_), .Y(new_n1642_));
  NAND3X1  g00640(.A(new_n1642_), .B(new_n1641_), .C(new_n1625_), .Y(new_n1643_));
  AND2X1   g00641(.A(new_n1624_), .B(new_n1611_), .Y(new_n1644_));
  NAND2X1  g00642(.A(new_n1623_), .B(new_n1617_), .Y(new_n1645_));
  OR2X1    g00643(.A(new_n1639_), .B(new_n1638_), .Y(new_n1646_));
  AOI21X1  g00644(.A0(new_n1646_), .A1(new_n1645_), .B0(new_n1611_), .Y(new_n1647_));
  OR2X1    g00645(.A(new_n1492_), .B(new_n1454_), .Y(new_n1648_));
  OAI21X1  g00646(.A0(new_n1647_), .A1(new_n1644_), .B0(new_n1648_), .Y(new_n1649_));
  AND2X1   g00647(.A(new_n1477_), .B(new_n1475_), .Y(new_n1650_));
  OR2X1    g00648(.A(new_n1479_), .B(new_n1650_), .Y(new_n1651_));
  XOR2X1   g00649(.A(new_n1486_), .B(new_n1651_), .Y(new_n1652_));
  XOR2X1   g00650(.A(new_n1490_), .B(new_n1488_), .Y(new_n1653_));
  NOR2X1   g00651(.A(new_n1486_), .B(new_n1480_), .Y(new_n1654_));
  NOR2X1   g00652(.A(new_n1490_), .B(new_n1488_), .Y(new_n1655_));
  AOI21X1  g00653(.A0(new_n1654_), .A1(new_n1653_), .B0(new_n1655_), .Y(new_n1656_));
  XOR2X1   g00654(.A(new_n1654_), .B(new_n1653_), .Y(new_n1657_));
  OAI21X1  g00655(.A0(new_n1656_), .A1(new_n1652_), .B0(new_n1657_), .Y(new_n1658_));
  XOR2X1   g00656(.A(new_n1468_), .B(new_n1462_), .Y(new_n1659_));
  AOI21X1  g00657(.A0(new_n1458_), .A1(new_n1456_), .B0(new_n1461_), .Y(new_n1660_));
  NOR4X1   g00658(.A(new_n1472_), .B(new_n1470_), .C(new_n1468_), .D(new_n1660_), .Y(new_n1661_));
  NOR4X1   g00659(.A(new_n1490_), .B(new_n1488_), .C(new_n1486_), .D(new_n1480_), .Y(new_n1662_));
  OR4X1    g00660(.A(new_n1662_), .B(new_n1652_), .C(new_n1661_), .D(new_n1659_), .Y(new_n1663_));
  XOR2X1   g00661(.A(new_n1472_), .B(new_n1470_), .Y(new_n1664_));
  NOR2X1   g00662(.A(new_n1468_), .B(new_n1660_), .Y(new_n1665_));
  NOR2X1   g00663(.A(new_n1472_), .B(new_n1470_), .Y(new_n1666_));
  AOI21X1  g00664(.A0(new_n1665_), .A1(new_n1664_), .B0(new_n1666_), .Y(new_n1667_));
  XOR2X1   g00665(.A(new_n1665_), .B(new_n1664_), .Y(new_n1668_));
  OAI21X1  g00666(.A0(new_n1667_), .A1(new_n1659_), .B0(new_n1668_), .Y(new_n1669_));
  XOR2X1   g00667(.A(new_n1669_), .B(new_n1663_), .Y(new_n1670_));
  AND2X1   g00668(.A(new_n1669_), .B(new_n1663_), .Y(new_n1671_));
  OR2X1    g00669(.A(new_n1468_), .B(new_n1660_), .Y(new_n1672_));
  XOR2X1   g00670(.A(new_n1672_), .B(new_n1664_), .Y(new_n1673_));
  OR4X1    g00671(.A(new_n1652_), .B(new_n1661_), .C(new_n1673_), .D(new_n1659_), .Y(new_n1674_));
  OR4X1    g00672(.A(new_n1490_), .B(new_n1488_), .C(new_n1486_), .D(new_n1480_), .Y(new_n1675_));
  OAI21X1  g00673(.A0(new_n1667_), .A1(new_n1659_), .B0(new_n1675_), .Y(new_n1676_));
  NOR2X1   g00674(.A(new_n1676_), .B(new_n1674_), .Y(new_n1677_));
  OR2X1    g00675(.A(new_n1677_), .B(new_n1671_), .Y(new_n1678_));
  MX2X1    g00676(.A(new_n1678_), .B(new_n1670_), .S0(new_n1658_), .Y(new_n1679_));
  AOI21X1  g00677(.A0(new_n1649_), .A1(new_n1643_), .B0(new_n1679_), .Y(new_n1680_));
  INVX1    g00678(.A(new_n1658_), .Y(new_n1681_));
  AND2X1   g00679(.A(new_n1670_), .B(new_n1658_), .Y(new_n1682_));
  AOI21X1  g00680(.A0(new_n1678_), .A1(new_n1681_), .B0(new_n1682_), .Y(new_n1683_));
  NAND3X1  g00681(.A(new_n1648_), .B(new_n1641_), .C(new_n1625_), .Y(new_n1684_));
  OAI21X1  g00682(.A0(new_n1647_), .A1(new_n1644_), .B0(new_n1642_), .Y(new_n1685_));
  AOI21X1  g00683(.A0(new_n1685_), .A1(new_n1684_), .B0(new_n1683_), .Y(new_n1686_));
  OR2X1    g00684(.A(new_n1686_), .B(new_n1680_), .Y(new_n1687_));
  NOR3X1   g00685(.A(new_n1592_), .B(new_n1599_), .C(new_n1596_), .Y(new_n1688_));
  AOI21X1  g00686(.A0(new_n1590_), .A1(new_n1586_), .B0(new_n1600_), .Y(new_n1689_));
  OAI21X1  g00687(.A0(new_n1689_), .A1(new_n1688_), .B0(new_n1687_), .Y(new_n1690_));
  OAI21X1  g00688(.A0(new_n1687_), .A1(new_n1602_), .B0(new_n1690_), .Y(new_n1691_));
  NOR3X1   g00689(.A(new_n1495_), .B(new_n1502_), .C(new_n1499_), .Y(new_n1692_));
  AOI21X1  g00690(.A0(new_n1339_), .A1(new_n1334_), .B0(new_n1503_), .Y(new_n1693_));
  OAI21X1  g00691(.A0(new_n1693_), .A1(new_n1692_), .B0(new_n1691_), .Y(new_n1694_));
  OAI21X1  g00692(.A0(new_n1691_), .A1(new_n1505_), .B0(new_n1694_), .Y(new_n1695_));
  INVX1    g00693(.A(\A[776] ), .Y(new_n1696_));
  OR2X1    g00694(.A(new_n1696_), .B(\A[775] ), .Y(new_n1697_));
  INVX1    g00695(.A(\A[777] ), .Y(new_n1698_));
  AOI21X1  g00696(.A0(new_n1696_), .A1(\A[775] ), .B0(new_n1698_), .Y(new_n1699_));
  XOR2X1   g00697(.A(\A[776] ), .B(\A[775] ), .Y(new_n1700_));
  AND2X1   g00698(.A(new_n1700_), .B(new_n1698_), .Y(new_n1701_));
  AOI21X1  g00699(.A0(new_n1699_), .A1(new_n1697_), .B0(new_n1701_), .Y(new_n1702_));
  INVX1    g00700(.A(\A[780] ), .Y(new_n1703_));
  INVX1    g00701(.A(\A[779] ), .Y(new_n1704_));
  OR2X1    g00702(.A(new_n1704_), .B(\A[778] ), .Y(new_n1705_));
  AOI21X1  g00703(.A0(new_n1704_), .A1(\A[778] ), .B0(new_n1703_), .Y(new_n1706_));
  XOR2X1   g00704(.A(\A[779] ), .B(\A[778] ), .Y(new_n1707_));
  AOI22X1  g00705(.A0(new_n1707_), .A1(new_n1703_), .B0(new_n1706_), .B1(new_n1705_), .Y(new_n1708_));
  OR2X1    g00706(.A(new_n1708_), .B(new_n1702_), .Y(new_n1709_));
  AND2X1   g00707(.A(\A[779] ), .B(\A[778] ), .Y(new_n1710_));
  AND2X1   g00708(.A(new_n1707_), .B(\A[780] ), .Y(new_n1711_));
  OR2X1    g00709(.A(new_n1711_), .B(new_n1710_), .Y(new_n1712_));
  AND2X1   g00710(.A(\A[776] ), .B(\A[775] ), .Y(new_n1713_));
  AOI21X1  g00711(.A0(new_n1700_), .A1(\A[777] ), .B0(new_n1713_), .Y(new_n1714_));
  XOR2X1   g00712(.A(new_n1714_), .B(new_n1712_), .Y(new_n1715_));
  XOR2X1   g00713(.A(new_n1715_), .B(new_n1709_), .Y(new_n1716_));
  XOR2X1   g00714(.A(new_n1708_), .B(new_n1702_), .Y(new_n1717_));
  AOI21X1  g00715(.A0(new_n1707_), .A1(\A[780] ), .B0(new_n1710_), .Y(new_n1718_));
  OR2X1    g00716(.A(new_n1714_), .B(new_n1718_), .Y(new_n1719_));
  OAI21X1  g00717(.A0(new_n1715_), .A1(new_n1709_), .B0(new_n1719_), .Y(new_n1720_));
  NAND2X1  g00718(.A(new_n1720_), .B(new_n1717_), .Y(new_n1721_));
  AND2X1   g00719(.A(new_n1721_), .B(new_n1716_), .Y(new_n1722_));
  NAND2X1  g00720(.A(new_n1721_), .B(new_n1716_), .Y(new_n1723_));
  AND2X1   g00721(.A(\A[785] ), .B(\A[784] ), .Y(new_n1724_));
  XOR2X1   g00722(.A(\A[785] ), .B(\A[784] ), .Y(new_n1725_));
  AOI21X1  g00723(.A0(new_n1725_), .A1(\A[786] ), .B0(new_n1724_), .Y(new_n1726_));
  AND2X1   g00724(.A(\A[782] ), .B(\A[781] ), .Y(new_n1727_));
  XOR2X1   g00725(.A(\A[782] ), .B(\A[781] ), .Y(new_n1728_));
  AOI21X1  g00726(.A0(new_n1728_), .A1(\A[783] ), .B0(new_n1727_), .Y(new_n1729_));
  INVX1    g00727(.A(\A[782] ), .Y(new_n1730_));
  OR2X1    g00728(.A(new_n1730_), .B(\A[781] ), .Y(new_n1731_));
  INVX1    g00729(.A(\A[783] ), .Y(new_n1732_));
  AOI21X1  g00730(.A0(new_n1730_), .A1(\A[781] ), .B0(new_n1732_), .Y(new_n1733_));
  AND2X1   g00731(.A(new_n1728_), .B(new_n1732_), .Y(new_n1734_));
  AOI21X1  g00732(.A0(new_n1733_), .A1(new_n1731_), .B0(new_n1734_), .Y(new_n1735_));
  INVX1    g00733(.A(\A[786] ), .Y(new_n1736_));
  INVX1    g00734(.A(\A[785] ), .Y(new_n1737_));
  OR2X1    g00735(.A(new_n1737_), .B(\A[784] ), .Y(new_n1738_));
  AOI21X1  g00736(.A0(new_n1737_), .A1(\A[784] ), .B0(new_n1736_), .Y(new_n1739_));
  AOI22X1  g00737(.A0(new_n1739_), .A1(new_n1738_), .B0(new_n1725_), .B1(new_n1736_), .Y(new_n1740_));
  OR4X1    g00738(.A(new_n1740_), .B(new_n1735_), .C(new_n1729_), .D(new_n1726_), .Y(new_n1741_));
  OR4X1    g00739(.A(new_n1714_), .B(new_n1718_), .C(new_n1708_), .D(new_n1702_), .Y(new_n1742_));
  XOR2X1   g00740(.A(new_n1740_), .B(new_n1735_), .Y(new_n1743_));
  NAND4X1  g00741(.A(new_n1743_), .B(new_n1742_), .C(new_n1741_), .D(new_n1717_), .Y(new_n1744_));
  XOR2X1   g00742(.A(new_n1729_), .B(new_n1726_), .Y(new_n1745_));
  NOR2X1   g00743(.A(new_n1740_), .B(new_n1735_), .Y(new_n1746_));
  NOR2X1   g00744(.A(new_n1729_), .B(new_n1726_), .Y(new_n1747_));
  AOI21X1  g00745(.A0(new_n1746_), .A1(new_n1745_), .B0(new_n1747_), .Y(new_n1748_));
  XOR2X1   g00746(.A(new_n1746_), .B(new_n1745_), .Y(new_n1749_));
  AND2X1   g00747(.A(new_n1733_), .B(new_n1731_), .Y(new_n1750_));
  OR2X1    g00748(.A(new_n1734_), .B(new_n1750_), .Y(new_n1751_));
  XOR2X1   g00749(.A(new_n1740_), .B(new_n1751_), .Y(new_n1752_));
  OAI21X1  g00750(.A0(new_n1752_), .A1(new_n1748_), .B0(new_n1749_), .Y(new_n1753_));
  XOR2X1   g00751(.A(new_n1753_), .B(new_n1744_), .Y(new_n1754_));
  AND2X1   g00752(.A(new_n1754_), .B(new_n1723_), .Y(new_n1755_));
  INVX1    g00753(.A(new_n1744_), .Y(new_n1756_));
  OR2X1    g00754(.A(new_n1740_), .B(new_n1735_), .Y(new_n1757_));
  XOR2X1   g00755(.A(new_n1757_), .B(new_n1745_), .Y(new_n1758_));
  NOR2X1   g00756(.A(new_n1752_), .B(new_n1748_), .Y(new_n1759_));
  NOR2X1   g00757(.A(new_n1759_), .B(new_n1758_), .Y(new_n1760_));
  NOR4X1   g00758(.A(new_n1714_), .B(new_n1718_), .C(new_n1708_), .D(new_n1702_), .Y(new_n1761_));
  NAND2X1  g00759(.A(new_n1743_), .B(new_n1717_), .Y(new_n1762_));
  AOI21X1  g00760(.A0(new_n1752_), .A1(new_n1758_), .B0(new_n1748_), .Y(new_n1763_));
  OR4X1    g00761(.A(new_n1763_), .B(new_n1762_), .C(new_n1761_), .D(new_n1758_), .Y(new_n1764_));
  OAI21X1  g00762(.A0(new_n1760_), .A1(new_n1756_), .B0(new_n1764_), .Y(new_n1765_));
  AOI21X1  g00763(.A0(new_n1765_), .A1(new_n1722_), .B0(new_n1755_), .Y(new_n1766_));
  INVX1    g00764(.A(\A[788] ), .Y(new_n1767_));
  OR2X1    g00765(.A(new_n1767_), .B(\A[787] ), .Y(new_n1768_));
  INVX1    g00766(.A(\A[789] ), .Y(new_n1769_));
  AOI21X1  g00767(.A0(new_n1767_), .A1(\A[787] ), .B0(new_n1769_), .Y(new_n1770_));
  XOR2X1   g00768(.A(\A[788] ), .B(\A[787] ), .Y(new_n1771_));
  AND2X1   g00769(.A(new_n1771_), .B(new_n1769_), .Y(new_n1772_));
  AOI21X1  g00770(.A0(new_n1770_), .A1(new_n1768_), .B0(new_n1772_), .Y(new_n1773_));
  INVX1    g00771(.A(\A[792] ), .Y(new_n1774_));
  INVX1    g00772(.A(\A[791] ), .Y(new_n1775_));
  OR2X1    g00773(.A(new_n1775_), .B(\A[790] ), .Y(new_n1776_));
  AOI21X1  g00774(.A0(new_n1775_), .A1(\A[790] ), .B0(new_n1774_), .Y(new_n1777_));
  XOR2X1   g00775(.A(\A[791] ), .B(\A[790] ), .Y(new_n1778_));
  AOI22X1  g00776(.A0(new_n1778_), .A1(new_n1774_), .B0(new_n1777_), .B1(new_n1776_), .Y(new_n1779_));
  NOR2X1   g00777(.A(new_n1779_), .B(new_n1773_), .Y(new_n1780_));
  AND2X1   g00778(.A(\A[791] ), .B(\A[790] ), .Y(new_n1781_));
  AND2X1   g00779(.A(new_n1778_), .B(\A[792] ), .Y(new_n1782_));
  OR2X1    g00780(.A(new_n1782_), .B(new_n1781_), .Y(new_n1783_));
  AND2X1   g00781(.A(\A[788] ), .B(\A[787] ), .Y(new_n1784_));
  AOI21X1  g00782(.A0(new_n1771_), .A1(\A[789] ), .B0(new_n1784_), .Y(new_n1785_));
  XOR2X1   g00783(.A(new_n1785_), .B(new_n1783_), .Y(new_n1786_));
  XOR2X1   g00784(.A(new_n1786_), .B(new_n1780_), .Y(new_n1787_));
  XOR2X1   g00785(.A(new_n1779_), .B(new_n1773_), .Y(new_n1788_));
  OR2X1    g00786(.A(new_n1779_), .B(new_n1773_), .Y(new_n1789_));
  AOI21X1  g00787(.A0(new_n1778_), .A1(\A[792] ), .B0(new_n1781_), .Y(new_n1790_));
  OR2X1    g00788(.A(new_n1785_), .B(new_n1790_), .Y(new_n1791_));
  OAI21X1  g00789(.A0(new_n1786_), .A1(new_n1789_), .B0(new_n1791_), .Y(new_n1792_));
  AND2X1   g00790(.A(new_n1792_), .B(new_n1788_), .Y(new_n1793_));
  OR2X1    g00791(.A(new_n1793_), .B(new_n1787_), .Y(new_n1794_));
  AND2X1   g00792(.A(\A[797] ), .B(\A[796] ), .Y(new_n1795_));
  XOR2X1   g00793(.A(\A[797] ), .B(\A[796] ), .Y(new_n1796_));
  AOI21X1  g00794(.A0(new_n1796_), .A1(\A[798] ), .B0(new_n1795_), .Y(new_n1797_));
  AND2X1   g00795(.A(\A[794] ), .B(\A[793] ), .Y(new_n1798_));
  XOR2X1   g00796(.A(\A[794] ), .B(\A[793] ), .Y(new_n1799_));
  AOI21X1  g00797(.A0(new_n1799_), .A1(\A[795] ), .B0(new_n1798_), .Y(new_n1800_));
  INVX1    g00798(.A(\A[794] ), .Y(new_n1801_));
  OR2X1    g00799(.A(new_n1801_), .B(\A[793] ), .Y(new_n1802_));
  INVX1    g00800(.A(\A[795] ), .Y(new_n1803_));
  AOI21X1  g00801(.A0(new_n1801_), .A1(\A[793] ), .B0(new_n1803_), .Y(new_n1804_));
  AND2X1   g00802(.A(new_n1799_), .B(new_n1803_), .Y(new_n1805_));
  AOI21X1  g00803(.A0(new_n1804_), .A1(new_n1802_), .B0(new_n1805_), .Y(new_n1806_));
  INVX1    g00804(.A(\A[798] ), .Y(new_n1807_));
  INVX1    g00805(.A(\A[797] ), .Y(new_n1808_));
  OR2X1    g00806(.A(new_n1808_), .B(\A[796] ), .Y(new_n1809_));
  AOI21X1  g00807(.A0(new_n1808_), .A1(\A[796] ), .B0(new_n1807_), .Y(new_n1810_));
  AOI22X1  g00808(.A0(new_n1810_), .A1(new_n1809_), .B0(new_n1796_), .B1(new_n1807_), .Y(new_n1811_));
  OR4X1    g00809(.A(new_n1811_), .B(new_n1806_), .C(new_n1800_), .D(new_n1797_), .Y(new_n1812_));
  OR4X1    g00810(.A(new_n1785_), .B(new_n1790_), .C(new_n1779_), .D(new_n1773_), .Y(new_n1813_));
  XOR2X1   g00811(.A(new_n1811_), .B(new_n1806_), .Y(new_n1814_));
  NAND4X1  g00812(.A(new_n1814_), .B(new_n1813_), .C(new_n1812_), .D(new_n1788_), .Y(new_n1815_));
  XOR2X1   g00813(.A(new_n1800_), .B(new_n1797_), .Y(new_n1816_));
  NOR2X1   g00814(.A(new_n1811_), .B(new_n1806_), .Y(new_n1817_));
  NOR2X1   g00815(.A(new_n1800_), .B(new_n1797_), .Y(new_n1818_));
  AOI21X1  g00816(.A0(new_n1817_), .A1(new_n1816_), .B0(new_n1818_), .Y(new_n1819_));
  XOR2X1   g00817(.A(new_n1817_), .B(new_n1816_), .Y(new_n1820_));
  AND2X1   g00818(.A(new_n1804_), .B(new_n1802_), .Y(new_n1821_));
  OR2X1    g00819(.A(new_n1805_), .B(new_n1821_), .Y(new_n1822_));
  XOR2X1   g00820(.A(new_n1811_), .B(new_n1822_), .Y(new_n1823_));
  OAI21X1  g00821(.A0(new_n1823_), .A1(new_n1819_), .B0(new_n1820_), .Y(new_n1824_));
  XOR2X1   g00822(.A(new_n1824_), .B(new_n1815_), .Y(new_n1825_));
  AND2X1   g00823(.A(new_n1825_), .B(new_n1794_), .Y(new_n1826_));
  AND2X1   g00824(.A(new_n1770_), .B(new_n1768_), .Y(new_n1827_));
  OR2X1    g00825(.A(new_n1772_), .B(new_n1827_), .Y(new_n1828_));
  XOR2X1   g00826(.A(new_n1779_), .B(new_n1828_), .Y(new_n1829_));
  OR2X1    g00827(.A(new_n1811_), .B(new_n1806_), .Y(new_n1830_));
  XOR2X1   g00828(.A(new_n1830_), .B(new_n1816_), .Y(new_n1831_));
  NOR4X1   g00829(.A(new_n1785_), .B(new_n1790_), .C(new_n1779_), .D(new_n1773_), .Y(new_n1832_));
  NOR4X1   g00830(.A(new_n1823_), .B(new_n1832_), .C(new_n1831_), .D(new_n1829_), .Y(new_n1833_));
  AND2X1   g00831(.A(new_n1817_), .B(new_n1816_), .Y(new_n1834_));
  OAI22X1  g00832(.A0(new_n1814_), .A1(new_n1820_), .B0(new_n1818_), .B1(new_n1834_), .Y(new_n1835_));
  AOI22X1  g00833(.A0(new_n1835_), .A1(new_n1833_), .B0(new_n1824_), .B1(new_n1815_), .Y(new_n1836_));
  NAND2X1  g00834(.A(new_n1814_), .B(new_n1812_), .Y(new_n1837_));
  XOR2X1   g00835(.A(new_n1779_), .B(new_n1773_), .Y(new_n1838_));
  XOR2X1   g00836(.A(new_n1838_), .B(new_n1837_), .Y(new_n1839_));
  NAND2X1  g00837(.A(new_n1743_), .B(new_n1741_), .Y(new_n1840_));
  XOR2X1   g00838(.A(new_n1708_), .B(new_n1702_), .Y(new_n1841_));
  XOR2X1   g00839(.A(new_n1841_), .B(new_n1840_), .Y(new_n1842_));
  NOR2X1   g00840(.A(new_n1842_), .B(new_n1839_), .Y(new_n1843_));
  OAI21X1  g00841(.A0(new_n1836_), .A1(new_n1794_), .B0(new_n1843_), .Y(new_n1844_));
  NOR2X1   g00842(.A(new_n1844_), .B(new_n1826_), .Y(new_n1845_));
  NAND2X1  g00843(.A(new_n1825_), .B(new_n1794_), .Y(new_n1846_));
  OR2X1    g00844(.A(new_n1836_), .B(new_n1794_), .Y(new_n1847_));
  AOI21X1  g00845(.A0(new_n1847_), .A1(new_n1846_), .B0(new_n1843_), .Y(new_n1848_));
  OAI21X1  g00846(.A0(new_n1848_), .A1(new_n1845_), .B0(new_n1766_), .Y(new_n1849_));
  MX2X1    g00847(.A(new_n1765_), .B(new_n1754_), .S0(new_n1723_), .Y(new_n1850_));
  OR2X1    g00848(.A(new_n1842_), .B(new_n1839_), .Y(new_n1851_));
  OAI21X1  g00849(.A0(new_n1836_), .A1(new_n1794_), .B0(new_n1851_), .Y(new_n1852_));
  NOR2X1   g00850(.A(new_n1852_), .B(new_n1826_), .Y(new_n1853_));
  AOI21X1  g00851(.A0(new_n1847_), .A1(new_n1846_), .B0(new_n1851_), .Y(new_n1854_));
  OAI21X1  g00852(.A0(new_n1854_), .A1(new_n1853_), .B0(new_n1850_), .Y(new_n1855_));
  XOR2X1   g00853(.A(new_n1842_), .B(new_n1839_), .Y(new_n1856_));
  INVX1    g00854(.A(new_n1856_), .Y(new_n1857_));
  INVX1    g00855(.A(\A[769] ), .Y(new_n1858_));
  OR2X1    g00856(.A(\A[770] ), .B(new_n1858_), .Y(new_n1859_));
  INVX1    g00857(.A(\A[771] ), .Y(new_n1860_));
  AOI21X1  g00858(.A0(\A[770] ), .A1(new_n1858_), .B0(new_n1860_), .Y(new_n1861_));
  XOR2X1   g00859(.A(\A[770] ), .B(\A[769] ), .Y(new_n1862_));
  AND2X1   g00860(.A(new_n1862_), .B(new_n1860_), .Y(new_n1863_));
  AOI21X1  g00861(.A0(new_n1861_), .A1(new_n1859_), .B0(new_n1863_), .Y(new_n1864_));
  INVX1    g00862(.A(\A[774] ), .Y(new_n1865_));
  INVX1    g00863(.A(\A[772] ), .Y(new_n1866_));
  OR2X1    g00864(.A(\A[773] ), .B(new_n1866_), .Y(new_n1867_));
  AOI21X1  g00865(.A0(\A[773] ), .A1(new_n1866_), .B0(new_n1865_), .Y(new_n1868_));
  XOR2X1   g00866(.A(\A[773] ), .B(\A[772] ), .Y(new_n1869_));
  AOI22X1  g00867(.A0(new_n1869_), .A1(new_n1865_), .B0(new_n1868_), .B1(new_n1867_), .Y(new_n1870_));
  AND2X1   g00868(.A(\A[773] ), .B(\A[772] ), .Y(new_n1871_));
  AOI21X1  g00869(.A0(new_n1869_), .A1(\A[774] ), .B0(new_n1871_), .Y(new_n1872_));
  AND2X1   g00870(.A(\A[770] ), .B(\A[769] ), .Y(new_n1873_));
  AOI21X1  g00871(.A0(new_n1862_), .A1(\A[771] ), .B0(new_n1873_), .Y(new_n1874_));
  XOR2X1   g00872(.A(new_n1870_), .B(new_n1864_), .Y(new_n1875_));
  INVX1    g00873(.A(\A[763] ), .Y(new_n1876_));
  OR2X1    g00874(.A(\A[764] ), .B(new_n1876_), .Y(new_n1877_));
  INVX1    g00875(.A(\A[765] ), .Y(new_n1878_));
  AOI21X1  g00876(.A0(\A[764] ), .A1(new_n1876_), .B0(new_n1878_), .Y(new_n1879_));
  XOR2X1   g00877(.A(\A[764] ), .B(\A[763] ), .Y(new_n1880_));
  AND2X1   g00878(.A(new_n1880_), .B(new_n1878_), .Y(new_n1881_));
  AOI21X1  g00879(.A0(new_n1879_), .A1(new_n1877_), .B0(new_n1881_), .Y(new_n1882_));
  INVX1    g00880(.A(\A[768] ), .Y(new_n1883_));
  INVX1    g00881(.A(\A[766] ), .Y(new_n1884_));
  OR2X1    g00882(.A(\A[767] ), .B(new_n1884_), .Y(new_n1885_));
  AOI21X1  g00883(.A0(\A[767] ), .A1(new_n1884_), .B0(new_n1883_), .Y(new_n1886_));
  XOR2X1   g00884(.A(\A[767] ), .B(\A[766] ), .Y(new_n1887_));
  AOI22X1  g00885(.A0(new_n1887_), .A1(new_n1883_), .B0(new_n1886_), .B1(new_n1885_), .Y(new_n1888_));
  AND2X1   g00886(.A(\A[767] ), .B(\A[766] ), .Y(new_n1889_));
  AOI21X1  g00887(.A0(new_n1887_), .A1(\A[768] ), .B0(new_n1889_), .Y(new_n1890_));
  AND2X1   g00888(.A(\A[764] ), .B(\A[763] ), .Y(new_n1891_));
  AOI21X1  g00889(.A0(new_n1880_), .A1(\A[765] ), .B0(new_n1891_), .Y(new_n1892_));
  XOR2X1   g00890(.A(new_n1888_), .B(new_n1882_), .Y(new_n1893_));
  XOR2X1   g00891(.A(new_n1893_), .B(new_n1875_), .Y(new_n1894_));
  INVX1    g00892(.A(\A[757] ), .Y(new_n1895_));
  OR2X1    g00893(.A(\A[758] ), .B(new_n1895_), .Y(new_n1896_));
  INVX1    g00894(.A(\A[759] ), .Y(new_n1897_));
  AOI21X1  g00895(.A0(\A[758] ), .A1(new_n1895_), .B0(new_n1897_), .Y(new_n1898_));
  AND2X1   g00896(.A(new_n1898_), .B(new_n1896_), .Y(new_n1899_));
  XOR2X1   g00897(.A(\A[758] ), .B(\A[757] ), .Y(new_n1900_));
  AND2X1   g00898(.A(new_n1900_), .B(new_n1897_), .Y(new_n1901_));
  OR2X1    g00899(.A(new_n1901_), .B(new_n1899_), .Y(new_n1902_));
  INVX1    g00900(.A(\A[762] ), .Y(new_n1903_));
  INVX1    g00901(.A(\A[760] ), .Y(new_n1904_));
  OR2X1    g00902(.A(\A[761] ), .B(new_n1904_), .Y(new_n1905_));
  AOI21X1  g00903(.A0(\A[761] ), .A1(new_n1904_), .B0(new_n1903_), .Y(new_n1906_));
  XOR2X1   g00904(.A(\A[761] ), .B(\A[760] ), .Y(new_n1907_));
  AOI22X1  g00905(.A0(new_n1907_), .A1(new_n1903_), .B0(new_n1906_), .B1(new_n1905_), .Y(new_n1908_));
  AND2X1   g00906(.A(\A[761] ), .B(\A[760] ), .Y(new_n1909_));
  AOI21X1  g00907(.A0(new_n1907_), .A1(\A[762] ), .B0(new_n1909_), .Y(new_n1910_));
  AND2X1   g00908(.A(\A[758] ), .B(\A[757] ), .Y(new_n1911_));
  AOI21X1  g00909(.A0(new_n1900_), .A1(\A[759] ), .B0(new_n1911_), .Y(new_n1912_));
  XOR2X1   g00910(.A(new_n1908_), .B(new_n1902_), .Y(new_n1913_));
  INVX1    g00911(.A(\A[751] ), .Y(new_n1914_));
  OR2X1    g00912(.A(\A[752] ), .B(new_n1914_), .Y(new_n1915_));
  INVX1    g00913(.A(\A[753] ), .Y(new_n1916_));
  AOI21X1  g00914(.A0(\A[752] ), .A1(new_n1914_), .B0(new_n1916_), .Y(new_n1917_));
  XOR2X1   g00915(.A(\A[752] ), .B(\A[751] ), .Y(new_n1918_));
  AND2X1   g00916(.A(new_n1918_), .B(new_n1916_), .Y(new_n1919_));
  AOI21X1  g00917(.A0(new_n1917_), .A1(new_n1915_), .B0(new_n1919_), .Y(new_n1920_));
  INVX1    g00918(.A(\A[756] ), .Y(new_n1921_));
  INVX1    g00919(.A(\A[754] ), .Y(new_n1922_));
  OR2X1    g00920(.A(\A[755] ), .B(new_n1922_), .Y(new_n1923_));
  AOI21X1  g00921(.A0(\A[755] ), .A1(new_n1922_), .B0(new_n1921_), .Y(new_n1924_));
  XOR2X1   g00922(.A(\A[755] ), .B(\A[754] ), .Y(new_n1925_));
  AOI22X1  g00923(.A0(new_n1925_), .A1(new_n1921_), .B0(new_n1924_), .B1(new_n1923_), .Y(new_n1926_));
  AND2X1   g00924(.A(\A[755] ), .B(\A[754] ), .Y(new_n1927_));
  AOI21X1  g00925(.A0(new_n1925_), .A1(\A[756] ), .B0(new_n1927_), .Y(new_n1928_));
  AND2X1   g00926(.A(\A[752] ), .B(\A[751] ), .Y(new_n1929_));
  AOI21X1  g00927(.A0(new_n1918_), .A1(\A[753] ), .B0(new_n1929_), .Y(new_n1930_));
  XOR2X1   g00928(.A(new_n1926_), .B(new_n1920_), .Y(new_n1931_));
  XOR2X1   g00929(.A(new_n1931_), .B(new_n1913_), .Y(new_n1932_));
  XOR2X1   g00930(.A(new_n1932_), .B(new_n1894_), .Y(new_n1933_));
  NOR2X1   g00931(.A(new_n1933_), .B(new_n1857_), .Y(new_n1934_));
  NAND3X1  g00932(.A(new_n1934_), .B(new_n1855_), .C(new_n1849_), .Y(new_n1935_));
  OR2X1    g00933(.A(new_n1844_), .B(new_n1826_), .Y(new_n1936_));
  NOR2X1   g00934(.A(new_n1836_), .B(new_n1794_), .Y(new_n1937_));
  OAI21X1  g00935(.A0(new_n1937_), .A1(new_n1826_), .B0(new_n1851_), .Y(new_n1938_));
  AOI21X1  g00936(.A0(new_n1938_), .A1(new_n1936_), .B0(new_n1850_), .Y(new_n1939_));
  OR2X1    g00937(.A(new_n1852_), .B(new_n1826_), .Y(new_n1940_));
  OAI21X1  g00938(.A0(new_n1937_), .A1(new_n1826_), .B0(new_n1843_), .Y(new_n1941_));
  AOI21X1  g00939(.A0(new_n1941_), .A1(new_n1940_), .B0(new_n1766_), .Y(new_n1942_));
  OR2X1    g00940(.A(new_n1933_), .B(new_n1857_), .Y(new_n1943_));
  OAI21X1  g00941(.A0(new_n1942_), .A1(new_n1939_), .B0(new_n1943_), .Y(new_n1944_));
  AND2X1   g00942(.A(new_n1944_), .B(new_n1935_), .Y(new_n1945_));
  AND2X1   g00943(.A(new_n1879_), .B(new_n1877_), .Y(new_n1946_));
  OR2X1    g00944(.A(new_n1881_), .B(new_n1946_), .Y(new_n1947_));
  XOR2X1   g00945(.A(new_n1888_), .B(new_n1947_), .Y(new_n1948_));
  XOR2X1   g00946(.A(new_n1892_), .B(new_n1890_), .Y(new_n1949_));
  NOR2X1   g00947(.A(new_n1888_), .B(new_n1882_), .Y(new_n1950_));
  NOR2X1   g00948(.A(new_n1892_), .B(new_n1890_), .Y(new_n1951_));
  AOI21X1  g00949(.A0(new_n1950_), .A1(new_n1949_), .B0(new_n1951_), .Y(new_n1952_));
  XOR2X1   g00950(.A(new_n1950_), .B(new_n1949_), .Y(new_n1953_));
  OAI21X1  g00951(.A0(new_n1952_), .A1(new_n1948_), .B0(new_n1953_), .Y(new_n1954_));
  AND2X1   g00952(.A(new_n1861_), .B(new_n1859_), .Y(new_n1955_));
  OR2X1    g00953(.A(new_n1863_), .B(new_n1955_), .Y(new_n1956_));
  XOR2X1   g00954(.A(new_n1870_), .B(new_n1956_), .Y(new_n1957_));
  NOR4X1   g00955(.A(new_n1874_), .B(new_n1872_), .C(new_n1870_), .D(new_n1864_), .Y(new_n1958_));
  NOR4X1   g00956(.A(new_n1892_), .B(new_n1890_), .C(new_n1888_), .D(new_n1882_), .Y(new_n1959_));
  OR4X1    g00957(.A(new_n1959_), .B(new_n1948_), .C(new_n1958_), .D(new_n1957_), .Y(new_n1960_));
  XOR2X1   g00958(.A(new_n1874_), .B(new_n1872_), .Y(new_n1961_));
  NOR2X1   g00959(.A(new_n1870_), .B(new_n1864_), .Y(new_n1962_));
  NOR2X1   g00960(.A(new_n1874_), .B(new_n1872_), .Y(new_n1963_));
  AOI21X1  g00961(.A0(new_n1962_), .A1(new_n1961_), .B0(new_n1963_), .Y(new_n1964_));
  XOR2X1   g00962(.A(new_n1962_), .B(new_n1961_), .Y(new_n1965_));
  OAI21X1  g00963(.A0(new_n1964_), .A1(new_n1957_), .B0(new_n1965_), .Y(new_n1966_));
  XOR2X1   g00964(.A(new_n1966_), .B(new_n1960_), .Y(new_n1967_));
  NAND2X1  g00965(.A(new_n1967_), .B(new_n1954_), .Y(new_n1968_));
  XOR2X1   g00966(.A(new_n1888_), .B(new_n1882_), .Y(new_n1969_));
  AND2X1   g00967(.A(new_n1887_), .B(\A[768] ), .Y(new_n1970_));
  OR2X1    g00968(.A(new_n1970_), .B(new_n1889_), .Y(new_n1971_));
  XOR2X1   g00969(.A(new_n1892_), .B(new_n1971_), .Y(new_n1972_));
  OR2X1    g00970(.A(new_n1888_), .B(new_n1882_), .Y(new_n1973_));
  OR2X1    g00971(.A(new_n1892_), .B(new_n1890_), .Y(new_n1974_));
  OAI21X1  g00972(.A0(new_n1973_), .A1(new_n1972_), .B0(new_n1974_), .Y(new_n1975_));
  XOR2X1   g00973(.A(new_n1950_), .B(new_n1972_), .Y(new_n1976_));
  AOI21X1  g00974(.A0(new_n1975_), .A1(new_n1969_), .B0(new_n1976_), .Y(new_n1977_));
  AND2X1   g00975(.A(new_n1966_), .B(new_n1960_), .Y(new_n1978_));
  OR2X1    g00976(.A(new_n1870_), .B(new_n1864_), .Y(new_n1979_));
  XOR2X1   g00977(.A(new_n1979_), .B(new_n1961_), .Y(new_n1980_));
  OR4X1    g00978(.A(new_n1948_), .B(new_n1958_), .C(new_n1980_), .D(new_n1957_), .Y(new_n1981_));
  OAI22X1  g00979(.A0(new_n1976_), .A1(new_n1952_), .B0(new_n1964_), .B1(new_n1957_), .Y(new_n1982_));
  NOR2X1   g00980(.A(new_n1982_), .B(new_n1981_), .Y(new_n1983_));
  OAI21X1  g00981(.A0(new_n1983_), .A1(new_n1978_), .B0(new_n1977_), .Y(new_n1984_));
  INVX1    g00982(.A(new_n1894_), .Y(new_n1985_));
  NOR2X1   g00983(.A(new_n1932_), .B(new_n1985_), .Y(new_n1986_));
  NAND3X1  g00984(.A(new_n1986_), .B(new_n1984_), .C(new_n1968_), .Y(new_n1987_));
  AND2X1   g00985(.A(new_n1967_), .B(new_n1954_), .Y(new_n1988_));
  NAND2X1  g00986(.A(new_n1966_), .B(new_n1960_), .Y(new_n1989_));
  OR2X1    g00987(.A(new_n1982_), .B(new_n1981_), .Y(new_n1990_));
  AOI21X1  g00988(.A0(new_n1990_), .A1(new_n1989_), .B0(new_n1954_), .Y(new_n1991_));
  OR2X1    g00989(.A(new_n1932_), .B(new_n1985_), .Y(new_n1992_));
  OAI21X1  g00990(.A0(new_n1991_), .A1(new_n1988_), .B0(new_n1992_), .Y(new_n1993_));
  AND2X1   g00991(.A(new_n1917_), .B(new_n1915_), .Y(new_n1994_));
  OR2X1    g00992(.A(new_n1919_), .B(new_n1994_), .Y(new_n1995_));
  XOR2X1   g00993(.A(new_n1926_), .B(new_n1995_), .Y(new_n1996_));
  XOR2X1   g00994(.A(new_n1930_), .B(new_n1928_), .Y(new_n1997_));
  NOR2X1   g00995(.A(new_n1926_), .B(new_n1920_), .Y(new_n1998_));
  NOR2X1   g00996(.A(new_n1930_), .B(new_n1928_), .Y(new_n1999_));
  AOI21X1  g00997(.A0(new_n1998_), .A1(new_n1997_), .B0(new_n1999_), .Y(new_n2000_));
  XOR2X1   g00998(.A(new_n1998_), .B(new_n1997_), .Y(new_n2001_));
  OAI21X1  g00999(.A0(new_n2000_), .A1(new_n1996_), .B0(new_n2001_), .Y(new_n2002_));
  XOR2X1   g01000(.A(new_n1908_), .B(new_n1902_), .Y(new_n2003_));
  AOI21X1  g01001(.A0(new_n1898_), .A1(new_n1896_), .B0(new_n1901_), .Y(new_n2004_));
  NOR4X1   g01002(.A(new_n1912_), .B(new_n1910_), .C(new_n1908_), .D(new_n2004_), .Y(new_n2005_));
  NOR4X1   g01003(.A(new_n1930_), .B(new_n1928_), .C(new_n1926_), .D(new_n1920_), .Y(new_n2006_));
  OR4X1    g01004(.A(new_n2006_), .B(new_n1996_), .C(new_n2005_), .D(new_n2003_), .Y(new_n2007_));
  XOR2X1   g01005(.A(new_n1912_), .B(new_n1910_), .Y(new_n2008_));
  NOR2X1   g01006(.A(new_n1908_), .B(new_n2004_), .Y(new_n2009_));
  NOR2X1   g01007(.A(new_n1912_), .B(new_n1910_), .Y(new_n2010_));
  AOI21X1  g01008(.A0(new_n2009_), .A1(new_n2008_), .B0(new_n2010_), .Y(new_n2011_));
  XOR2X1   g01009(.A(new_n2009_), .B(new_n2008_), .Y(new_n2012_));
  OAI21X1  g01010(.A0(new_n2011_), .A1(new_n2003_), .B0(new_n2012_), .Y(new_n2013_));
  XOR2X1   g01011(.A(new_n2013_), .B(new_n2007_), .Y(new_n2014_));
  AND2X1   g01012(.A(new_n2013_), .B(new_n2007_), .Y(new_n2015_));
  OR2X1    g01013(.A(new_n1908_), .B(new_n2004_), .Y(new_n2016_));
  XOR2X1   g01014(.A(new_n2016_), .B(new_n2008_), .Y(new_n2017_));
  OR4X1    g01015(.A(new_n1996_), .B(new_n2005_), .C(new_n2017_), .D(new_n2003_), .Y(new_n2018_));
  AND2X1   g01016(.A(new_n1925_), .B(\A[756] ), .Y(new_n2019_));
  OR2X1    g01017(.A(new_n2019_), .B(new_n1927_), .Y(new_n2020_));
  XOR2X1   g01018(.A(new_n1930_), .B(new_n2020_), .Y(new_n2021_));
  XOR2X1   g01019(.A(new_n1998_), .B(new_n2021_), .Y(new_n2022_));
  OAI22X1  g01020(.A0(new_n2022_), .A1(new_n2000_), .B0(new_n2011_), .B1(new_n2003_), .Y(new_n2023_));
  NOR2X1   g01021(.A(new_n2023_), .B(new_n2018_), .Y(new_n2024_));
  OR2X1    g01022(.A(new_n2024_), .B(new_n2015_), .Y(new_n2025_));
  MX2X1    g01023(.A(new_n2025_), .B(new_n2014_), .S0(new_n2002_), .Y(new_n2026_));
  AOI21X1  g01024(.A0(new_n1993_), .A1(new_n1987_), .B0(new_n2026_), .Y(new_n2027_));
  INVX1    g01025(.A(new_n2002_), .Y(new_n2028_));
  AND2X1   g01026(.A(new_n2014_), .B(new_n2002_), .Y(new_n2029_));
  AOI21X1  g01027(.A0(new_n2025_), .A1(new_n2028_), .B0(new_n2029_), .Y(new_n2030_));
  NAND3X1  g01028(.A(new_n1992_), .B(new_n1984_), .C(new_n1968_), .Y(new_n2031_));
  OAI21X1  g01029(.A0(new_n1991_), .A1(new_n1988_), .B0(new_n1986_), .Y(new_n2032_));
  AOI21X1  g01030(.A0(new_n2032_), .A1(new_n2031_), .B0(new_n2030_), .Y(new_n2033_));
  NOR2X1   g01031(.A(new_n2033_), .B(new_n2027_), .Y(new_n2034_));
  NAND3X1  g01032(.A(new_n1943_), .B(new_n1855_), .C(new_n1849_), .Y(new_n2035_));
  OAI21X1  g01033(.A0(new_n1942_), .A1(new_n1939_), .B0(new_n1934_), .Y(new_n2036_));
  AND2X1   g01034(.A(new_n2036_), .B(new_n2035_), .Y(new_n2037_));
  MX2X1    g01035(.A(new_n2037_), .B(new_n1945_), .S0(new_n2034_), .Y(new_n2038_));
  INVX1    g01036(.A(\A[812] ), .Y(new_n2039_));
  OR2X1    g01037(.A(new_n2039_), .B(\A[811] ), .Y(new_n2040_));
  INVX1    g01038(.A(\A[813] ), .Y(new_n2041_));
  AOI21X1  g01039(.A0(new_n2039_), .A1(\A[811] ), .B0(new_n2041_), .Y(new_n2042_));
  XOR2X1   g01040(.A(\A[812] ), .B(\A[811] ), .Y(new_n2043_));
  AND2X1   g01041(.A(new_n2043_), .B(new_n2041_), .Y(new_n2044_));
  AOI21X1  g01042(.A0(new_n2042_), .A1(new_n2040_), .B0(new_n2044_), .Y(new_n2045_));
  INVX1    g01043(.A(\A[816] ), .Y(new_n2046_));
  INVX1    g01044(.A(\A[815] ), .Y(new_n2047_));
  OR2X1    g01045(.A(new_n2047_), .B(\A[814] ), .Y(new_n2048_));
  AOI21X1  g01046(.A0(new_n2047_), .A1(\A[814] ), .B0(new_n2046_), .Y(new_n2049_));
  XOR2X1   g01047(.A(\A[815] ), .B(\A[814] ), .Y(new_n2050_));
  AOI22X1  g01048(.A0(new_n2050_), .A1(new_n2046_), .B0(new_n2049_), .B1(new_n2048_), .Y(new_n2051_));
  NOR2X1   g01049(.A(new_n2051_), .B(new_n2045_), .Y(new_n2052_));
  AND2X1   g01050(.A(\A[815] ), .B(\A[814] ), .Y(new_n2053_));
  AND2X1   g01051(.A(new_n2050_), .B(\A[816] ), .Y(new_n2054_));
  OR2X1    g01052(.A(new_n2054_), .B(new_n2053_), .Y(new_n2055_));
  AND2X1   g01053(.A(\A[812] ), .B(\A[811] ), .Y(new_n2056_));
  AOI21X1  g01054(.A0(new_n2043_), .A1(\A[813] ), .B0(new_n2056_), .Y(new_n2057_));
  XOR2X1   g01055(.A(new_n2057_), .B(new_n2055_), .Y(new_n2058_));
  XOR2X1   g01056(.A(new_n2058_), .B(new_n2052_), .Y(new_n2059_));
  XOR2X1   g01057(.A(new_n2051_), .B(new_n2045_), .Y(new_n2060_));
  OR2X1    g01058(.A(new_n2051_), .B(new_n2045_), .Y(new_n2061_));
  AOI21X1  g01059(.A0(new_n2050_), .A1(\A[816] ), .B0(new_n2053_), .Y(new_n2062_));
  OR2X1    g01060(.A(new_n2057_), .B(new_n2062_), .Y(new_n2063_));
  OAI21X1  g01061(.A0(new_n2058_), .A1(new_n2061_), .B0(new_n2063_), .Y(new_n2064_));
  AND2X1   g01062(.A(new_n2064_), .B(new_n2060_), .Y(new_n2065_));
  OR2X1    g01063(.A(new_n2065_), .B(new_n2059_), .Y(new_n2066_));
  AND2X1   g01064(.A(\A[821] ), .B(\A[820] ), .Y(new_n2067_));
  XOR2X1   g01065(.A(\A[821] ), .B(\A[820] ), .Y(new_n2068_));
  AOI21X1  g01066(.A0(new_n2068_), .A1(\A[822] ), .B0(new_n2067_), .Y(new_n2069_));
  AND2X1   g01067(.A(\A[818] ), .B(\A[817] ), .Y(new_n2070_));
  XOR2X1   g01068(.A(\A[818] ), .B(\A[817] ), .Y(new_n2071_));
  AOI21X1  g01069(.A0(new_n2071_), .A1(\A[819] ), .B0(new_n2070_), .Y(new_n2072_));
  INVX1    g01070(.A(\A[818] ), .Y(new_n2073_));
  OR2X1    g01071(.A(new_n2073_), .B(\A[817] ), .Y(new_n2074_));
  INVX1    g01072(.A(\A[819] ), .Y(new_n2075_));
  AOI21X1  g01073(.A0(new_n2073_), .A1(\A[817] ), .B0(new_n2075_), .Y(new_n2076_));
  AND2X1   g01074(.A(new_n2071_), .B(new_n2075_), .Y(new_n2077_));
  AOI21X1  g01075(.A0(new_n2076_), .A1(new_n2074_), .B0(new_n2077_), .Y(new_n2078_));
  INVX1    g01076(.A(\A[822] ), .Y(new_n2079_));
  INVX1    g01077(.A(\A[821] ), .Y(new_n2080_));
  OR2X1    g01078(.A(new_n2080_), .B(\A[820] ), .Y(new_n2081_));
  AOI21X1  g01079(.A0(new_n2080_), .A1(\A[820] ), .B0(new_n2079_), .Y(new_n2082_));
  AOI22X1  g01080(.A0(new_n2082_), .A1(new_n2081_), .B0(new_n2068_), .B1(new_n2079_), .Y(new_n2083_));
  OR4X1    g01081(.A(new_n2083_), .B(new_n2078_), .C(new_n2072_), .D(new_n2069_), .Y(new_n2084_));
  OR4X1    g01082(.A(new_n2057_), .B(new_n2062_), .C(new_n2051_), .D(new_n2045_), .Y(new_n2085_));
  XOR2X1   g01083(.A(new_n2083_), .B(new_n2078_), .Y(new_n2086_));
  NAND4X1  g01084(.A(new_n2086_), .B(new_n2085_), .C(new_n2084_), .D(new_n2060_), .Y(new_n2087_));
  XOR2X1   g01085(.A(new_n2072_), .B(new_n2069_), .Y(new_n2088_));
  NOR2X1   g01086(.A(new_n2083_), .B(new_n2078_), .Y(new_n2089_));
  NOR2X1   g01087(.A(new_n2072_), .B(new_n2069_), .Y(new_n2090_));
  AOI21X1  g01088(.A0(new_n2089_), .A1(new_n2088_), .B0(new_n2090_), .Y(new_n2091_));
  XOR2X1   g01089(.A(new_n2089_), .B(new_n2088_), .Y(new_n2092_));
  AND2X1   g01090(.A(new_n2076_), .B(new_n2074_), .Y(new_n2093_));
  OR2X1    g01091(.A(new_n2077_), .B(new_n2093_), .Y(new_n2094_));
  XOR2X1   g01092(.A(new_n2083_), .B(new_n2094_), .Y(new_n2095_));
  OAI21X1  g01093(.A0(new_n2095_), .A1(new_n2091_), .B0(new_n2092_), .Y(new_n2096_));
  XOR2X1   g01094(.A(new_n2096_), .B(new_n2087_), .Y(new_n2097_));
  AND2X1   g01095(.A(new_n2097_), .B(new_n2066_), .Y(new_n2098_));
  AND2X1   g01096(.A(new_n2042_), .B(new_n2040_), .Y(new_n2099_));
  OR2X1    g01097(.A(new_n2044_), .B(new_n2099_), .Y(new_n2100_));
  XOR2X1   g01098(.A(new_n2051_), .B(new_n2100_), .Y(new_n2101_));
  OR2X1    g01099(.A(new_n2083_), .B(new_n2078_), .Y(new_n2102_));
  XOR2X1   g01100(.A(new_n2102_), .B(new_n2088_), .Y(new_n2103_));
  NOR4X1   g01101(.A(new_n2057_), .B(new_n2062_), .C(new_n2051_), .D(new_n2045_), .Y(new_n2104_));
  NOR4X1   g01102(.A(new_n2095_), .B(new_n2104_), .C(new_n2103_), .D(new_n2101_), .Y(new_n2105_));
  AND2X1   g01103(.A(new_n2089_), .B(new_n2088_), .Y(new_n2106_));
  OAI22X1  g01104(.A0(new_n2086_), .A1(new_n2092_), .B0(new_n2090_), .B1(new_n2106_), .Y(new_n2107_));
  AOI22X1  g01105(.A0(new_n2107_), .A1(new_n2105_), .B0(new_n2096_), .B1(new_n2087_), .Y(new_n2108_));
  AND2X1   g01106(.A(new_n2086_), .B(new_n2084_), .Y(new_n2109_));
  XOR2X1   g01107(.A(new_n2051_), .B(new_n2100_), .Y(new_n2110_));
  XOR2X1   g01108(.A(new_n2110_), .B(new_n2109_), .Y(new_n2111_));
  INVX1    g01109(.A(\A[805] ), .Y(new_n2112_));
  OR2X1    g01110(.A(\A[806] ), .B(new_n2112_), .Y(new_n2113_));
  INVX1    g01111(.A(\A[807] ), .Y(new_n2114_));
  AOI21X1  g01112(.A0(\A[806] ), .A1(new_n2112_), .B0(new_n2114_), .Y(new_n2115_));
  AND2X1   g01113(.A(new_n2115_), .B(new_n2113_), .Y(new_n2116_));
  XOR2X1   g01114(.A(\A[806] ), .B(\A[805] ), .Y(new_n2117_));
  AND2X1   g01115(.A(new_n2117_), .B(new_n2114_), .Y(new_n2118_));
  OR2X1    g01116(.A(new_n2118_), .B(new_n2116_), .Y(new_n2119_));
  INVX1    g01117(.A(\A[810] ), .Y(new_n2120_));
  INVX1    g01118(.A(\A[808] ), .Y(new_n2121_));
  OR2X1    g01119(.A(\A[809] ), .B(new_n2121_), .Y(new_n2122_));
  AOI21X1  g01120(.A0(\A[809] ), .A1(new_n2121_), .B0(new_n2120_), .Y(new_n2123_));
  XOR2X1   g01121(.A(\A[809] ), .B(\A[808] ), .Y(new_n2124_));
  AOI22X1  g01122(.A0(new_n2124_), .A1(new_n2120_), .B0(new_n2123_), .B1(new_n2122_), .Y(new_n2125_));
  AND2X1   g01123(.A(\A[809] ), .B(\A[808] ), .Y(new_n2126_));
  AOI21X1  g01124(.A0(new_n2124_), .A1(\A[810] ), .B0(new_n2126_), .Y(new_n2127_));
  AND2X1   g01125(.A(\A[806] ), .B(\A[805] ), .Y(new_n2128_));
  AOI21X1  g01126(.A0(new_n2117_), .A1(\A[807] ), .B0(new_n2128_), .Y(new_n2129_));
  XOR2X1   g01127(.A(new_n2125_), .B(new_n2119_), .Y(new_n2130_));
  INVX1    g01128(.A(\A[799] ), .Y(new_n2131_));
  OR2X1    g01129(.A(\A[800] ), .B(new_n2131_), .Y(new_n2132_));
  INVX1    g01130(.A(\A[801] ), .Y(new_n2133_));
  AOI21X1  g01131(.A0(\A[800] ), .A1(new_n2131_), .B0(new_n2133_), .Y(new_n2134_));
  XOR2X1   g01132(.A(\A[800] ), .B(\A[799] ), .Y(new_n2135_));
  AND2X1   g01133(.A(new_n2135_), .B(new_n2133_), .Y(new_n2136_));
  AOI21X1  g01134(.A0(new_n2134_), .A1(new_n2132_), .B0(new_n2136_), .Y(new_n2137_));
  INVX1    g01135(.A(\A[804] ), .Y(new_n2138_));
  INVX1    g01136(.A(\A[802] ), .Y(new_n2139_));
  OR2X1    g01137(.A(\A[803] ), .B(new_n2139_), .Y(new_n2140_));
  AOI21X1  g01138(.A0(\A[803] ), .A1(new_n2139_), .B0(new_n2138_), .Y(new_n2141_));
  XOR2X1   g01139(.A(\A[803] ), .B(\A[802] ), .Y(new_n2142_));
  AOI22X1  g01140(.A0(new_n2142_), .A1(new_n2138_), .B0(new_n2141_), .B1(new_n2140_), .Y(new_n2143_));
  AND2X1   g01141(.A(\A[803] ), .B(\A[802] ), .Y(new_n2144_));
  AOI21X1  g01142(.A0(new_n2142_), .A1(\A[804] ), .B0(new_n2144_), .Y(new_n2145_));
  AND2X1   g01143(.A(\A[800] ), .B(\A[799] ), .Y(new_n2146_));
  AOI21X1  g01144(.A0(new_n2135_), .A1(\A[801] ), .B0(new_n2146_), .Y(new_n2147_));
  XOR2X1   g01145(.A(new_n2143_), .B(new_n2137_), .Y(new_n2148_));
  XOR2X1   g01146(.A(new_n2148_), .B(new_n2130_), .Y(new_n2149_));
  NOR2X1   g01147(.A(new_n2149_), .B(new_n2111_), .Y(new_n2150_));
  OAI21X1  g01148(.A0(new_n2108_), .A1(new_n2066_), .B0(new_n2150_), .Y(new_n2151_));
  NOR2X1   g01149(.A(new_n2108_), .B(new_n2066_), .Y(new_n2152_));
  OR2X1    g01150(.A(new_n2149_), .B(new_n2111_), .Y(new_n2153_));
  OAI21X1  g01151(.A0(new_n2152_), .A1(new_n2098_), .B0(new_n2153_), .Y(new_n2154_));
  OAI21X1  g01152(.A0(new_n2151_), .A1(new_n2098_), .B0(new_n2154_), .Y(new_n2155_));
  AND2X1   g01153(.A(new_n2134_), .B(new_n2132_), .Y(new_n2156_));
  OR2X1    g01154(.A(new_n2136_), .B(new_n2156_), .Y(new_n2157_));
  XOR2X1   g01155(.A(new_n2143_), .B(new_n2157_), .Y(new_n2158_));
  XOR2X1   g01156(.A(new_n2147_), .B(new_n2145_), .Y(new_n2159_));
  NOR2X1   g01157(.A(new_n2143_), .B(new_n2137_), .Y(new_n2160_));
  NOR2X1   g01158(.A(new_n2147_), .B(new_n2145_), .Y(new_n2161_));
  AOI21X1  g01159(.A0(new_n2160_), .A1(new_n2159_), .B0(new_n2161_), .Y(new_n2162_));
  XOR2X1   g01160(.A(new_n2160_), .B(new_n2159_), .Y(new_n2163_));
  OAI21X1  g01161(.A0(new_n2162_), .A1(new_n2158_), .B0(new_n2163_), .Y(new_n2164_));
  INVX1    g01162(.A(new_n2164_), .Y(new_n2165_));
  XOR2X1   g01163(.A(new_n2125_), .B(new_n2119_), .Y(new_n2166_));
  AOI21X1  g01164(.A0(new_n2115_), .A1(new_n2113_), .B0(new_n2118_), .Y(new_n2167_));
  NOR4X1   g01165(.A(new_n2129_), .B(new_n2127_), .C(new_n2125_), .D(new_n2167_), .Y(new_n2168_));
  NOR4X1   g01166(.A(new_n2147_), .B(new_n2145_), .C(new_n2143_), .D(new_n2137_), .Y(new_n2169_));
  OR4X1    g01167(.A(new_n2169_), .B(new_n2158_), .C(new_n2168_), .D(new_n2166_), .Y(new_n2170_));
  XOR2X1   g01168(.A(new_n2129_), .B(new_n2127_), .Y(new_n2171_));
  NOR2X1   g01169(.A(new_n2125_), .B(new_n2167_), .Y(new_n2172_));
  NOR2X1   g01170(.A(new_n2129_), .B(new_n2127_), .Y(new_n2173_));
  AOI21X1  g01171(.A0(new_n2172_), .A1(new_n2171_), .B0(new_n2173_), .Y(new_n2174_));
  XOR2X1   g01172(.A(new_n2172_), .B(new_n2171_), .Y(new_n2175_));
  OAI21X1  g01173(.A0(new_n2174_), .A1(new_n2166_), .B0(new_n2175_), .Y(new_n2176_));
  XOR2X1   g01174(.A(new_n2176_), .B(new_n2170_), .Y(new_n2177_));
  AND2X1   g01175(.A(new_n2177_), .B(new_n2164_), .Y(new_n2178_));
  AND2X1   g01176(.A(new_n2176_), .B(new_n2170_), .Y(new_n2179_));
  OR2X1    g01177(.A(new_n2125_), .B(new_n2167_), .Y(new_n2180_));
  XOR2X1   g01178(.A(new_n2180_), .B(new_n2171_), .Y(new_n2181_));
  OR4X1    g01179(.A(new_n2158_), .B(new_n2168_), .C(new_n2181_), .D(new_n2166_), .Y(new_n2182_));
  INVX1    g01180(.A(new_n2159_), .Y(new_n2183_));
  XOR2X1   g01181(.A(new_n2160_), .B(new_n2183_), .Y(new_n2184_));
  OAI22X1  g01182(.A0(new_n2184_), .A1(new_n2162_), .B0(new_n2174_), .B1(new_n2166_), .Y(new_n2185_));
  NOR2X1   g01183(.A(new_n2185_), .B(new_n2182_), .Y(new_n2186_));
  OR2X1    g01184(.A(new_n2186_), .B(new_n2179_), .Y(new_n2187_));
  AOI21X1  g01185(.A0(new_n2187_), .A1(new_n2165_), .B0(new_n2178_), .Y(new_n2188_));
  NAND2X1  g01186(.A(new_n2097_), .B(new_n2066_), .Y(new_n2189_));
  OR2X1    g01187(.A(new_n2108_), .B(new_n2066_), .Y(new_n2190_));
  NAND3X1  g01188(.A(new_n2153_), .B(new_n2190_), .C(new_n2189_), .Y(new_n2191_));
  OAI21X1  g01189(.A0(new_n2152_), .A1(new_n2098_), .B0(new_n2150_), .Y(new_n2192_));
  NAND2X1  g01190(.A(new_n2192_), .B(new_n2191_), .Y(new_n2193_));
  MX2X1    g01191(.A(new_n2193_), .B(new_n2155_), .S0(new_n2188_), .Y(new_n2194_));
  INVX1    g01192(.A(\A[824] ), .Y(new_n2195_));
  OR2X1    g01193(.A(new_n2195_), .B(\A[823] ), .Y(new_n2196_));
  INVX1    g01194(.A(\A[825] ), .Y(new_n2197_));
  AOI21X1  g01195(.A0(new_n2195_), .A1(\A[823] ), .B0(new_n2197_), .Y(new_n2198_));
  XOR2X1   g01196(.A(\A[824] ), .B(\A[823] ), .Y(new_n2199_));
  AND2X1   g01197(.A(new_n2199_), .B(new_n2197_), .Y(new_n2200_));
  AOI21X1  g01198(.A0(new_n2198_), .A1(new_n2196_), .B0(new_n2200_), .Y(new_n2201_));
  INVX1    g01199(.A(\A[828] ), .Y(new_n2202_));
  INVX1    g01200(.A(\A[827] ), .Y(new_n2203_));
  OR2X1    g01201(.A(new_n2203_), .B(\A[826] ), .Y(new_n2204_));
  AOI21X1  g01202(.A0(new_n2203_), .A1(\A[826] ), .B0(new_n2202_), .Y(new_n2205_));
  XOR2X1   g01203(.A(\A[827] ), .B(\A[826] ), .Y(new_n2206_));
  AOI22X1  g01204(.A0(new_n2206_), .A1(new_n2202_), .B0(new_n2205_), .B1(new_n2204_), .Y(new_n2207_));
  OR2X1    g01205(.A(new_n2207_), .B(new_n2201_), .Y(new_n2208_));
  AND2X1   g01206(.A(\A[827] ), .B(\A[826] ), .Y(new_n2209_));
  AND2X1   g01207(.A(new_n2206_), .B(\A[828] ), .Y(new_n2210_));
  OR2X1    g01208(.A(new_n2210_), .B(new_n2209_), .Y(new_n2211_));
  AND2X1   g01209(.A(\A[824] ), .B(\A[823] ), .Y(new_n2212_));
  AOI21X1  g01210(.A0(new_n2199_), .A1(\A[825] ), .B0(new_n2212_), .Y(new_n2213_));
  XOR2X1   g01211(.A(new_n2213_), .B(new_n2211_), .Y(new_n2214_));
  XOR2X1   g01212(.A(new_n2214_), .B(new_n2208_), .Y(new_n2215_));
  XOR2X1   g01213(.A(new_n2207_), .B(new_n2201_), .Y(new_n2216_));
  AOI21X1  g01214(.A0(new_n2206_), .A1(\A[828] ), .B0(new_n2209_), .Y(new_n2217_));
  OR2X1    g01215(.A(new_n2213_), .B(new_n2217_), .Y(new_n2218_));
  OAI21X1  g01216(.A0(new_n2214_), .A1(new_n2208_), .B0(new_n2218_), .Y(new_n2219_));
  NAND2X1  g01217(.A(new_n2219_), .B(new_n2216_), .Y(new_n2220_));
  AND2X1   g01218(.A(new_n2220_), .B(new_n2215_), .Y(new_n2221_));
  NAND2X1  g01219(.A(new_n2220_), .B(new_n2215_), .Y(new_n2222_));
  AND2X1   g01220(.A(\A[833] ), .B(\A[832] ), .Y(new_n2223_));
  XOR2X1   g01221(.A(\A[833] ), .B(\A[832] ), .Y(new_n2224_));
  AOI21X1  g01222(.A0(new_n2224_), .A1(\A[834] ), .B0(new_n2223_), .Y(new_n2225_));
  AND2X1   g01223(.A(\A[830] ), .B(\A[829] ), .Y(new_n2226_));
  XOR2X1   g01224(.A(\A[830] ), .B(\A[829] ), .Y(new_n2227_));
  AOI21X1  g01225(.A0(new_n2227_), .A1(\A[831] ), .B0(new_n2226_), .Y(new_n2228_));
  INVX1    g01226(.A(\A[830] ), .Y(new_n2229_));
  OR2X1    g01227(.A(new_n2229_), .B(\A[829] ), .Y(new_n2230_));
  INVX1    g01228(.A(\A[831] ), .Y(new_n2231_));
  AOI21X1  g01229(.A0(new_n2229_), .A1(\A[829] ), .B0(new_n2231_), .Y(new_n2232_));
  AND2X1   g01230(.A(new_n2227_), .B(new_n2231_), .Y(new_n2233_));
  AOI21X1  g01231(.A0(new_n2232_), .A1(new_n2230_), .B0(new_n2233_), .Y(new_n2234_));
  INVX1    g01232(.A(\A[834] ), .Y(new_n2235_));
  INVX1    g01233(.A(\A[833] ), .Y(new_n2236_));
  OR2X1    g01234(.A(new_n2236_), .B(\A[832] ), .Y(new_n2237_));
  AOI21X1  g01235(.A0(new_n2236_), .A1(\A[832] ), .B0(new_n2235_), .Y(new_n2238_));
  AOI22X1  g01236(.A0(new_n2238_), .A1(new_n2237_), .B0(new_n2224_), .B1(new_n2235_), .Y(new_n2239_));
  OR4X1    g01237(.A(new_n2239_), .B(new_n2234_), .C(new_n2228_), .D(new_n2225_), .Y(new_n2240_));
  OR4X1    g01238(.A(new_n2213_), .B(new_n2217_), .C(new_n2207_), .D(new_n2201_), .Y(new_n2241_));
  XOR2X1   g01239(.A(new_n2239_), .B(new_n2234_), .Y(new_n2242_));
  NAND4X1  g01240(.A(new_n2242_), .B(new_n2241_), .C(new_n2240_), .D(new_n2216_), .Y(new_n2243_));
  XOR2X1   g01241(.A(new_n2228_), .B(new_n2225_), .Y(new_n2244_));
  NOR2X1   g01242(.A(new_n2239_), .B(new_n2234_), .Y(new_n2245_));
  NOR2X1   g01243(.A(new_n2228_), .B(new_n2225_), .Y(new_n2246_));
  AOI21X1  g01244(.A0(new_n2245_), .A1(new_n2244_), .B0(new_n2246_), .Y(new_n2247_));
  XOR2X1   g01245(.A(new_n2245_), .B(new_n2244_), .Y(new_n2248_));
  AND2X1   g01246(.A(new_n2232_), .B(new_n2230_), .Y(new_n2249_));
  OR2X1    g01247(.A(new_n2233_), .B(new_n2249_), .Y(new_n2250_));
  XOR2X1   g01248(.A(new_n2239_), .B(new_n2250_), .Y(new_n2251_));
  OAI21X1  g01249(.A0(new_n2251_), .A1(new_n2247_), .B0(new_n2248_), .Y(new_n2252_));
  XOR2X1   g01250(.A(new_n2252_), .B(new_n2243_), .Y(new_n2253_));
  AND2X1   g01251(.A(new_n2253_), .B(new_n2222_), .Y(new_n2254_));
  INVX1    g01252(.A(new_n2243_), .Y(new_n2255_));
  OR2X1    g01253(.A(new_n2239_), .B(new_n2234_), .Y(new_n2256_));
  XOR2X1   g01254(.A(new_n2256_), .B(new_n2244_), .Y(new_n2257_));
  NOR2X1   g01255(.A(new_n2251_), .B(new_n2247_), .Y(new_n2258_));
  NOR2X1   g01256(.A(new_n2258_), .B(new_n2257_), .Y(new_n2259_));
  NOR4X1   g01257(.A(new_n2213_), .B(new_n2217_), .C(new_n2207_), .D(new_n2201_), .Y(new_n2260_));
  NAND2X1  g01258(.A(new_n2242_), .B(new_n2216_), .Y(new_n2261_));
  AOI21X1  g01259(.A0(new_n2251_), .A1(new_n2257_), .B0(new_n2247_), .Y(new_n2262_));
  OR4X1    g01260(.A(new_n2262_), .B(new_n2261_), .C(new_n2260_), .D(new_n2257_), .Y(new_n2263_));
  OAI21X1  g01261(.A0(new_n2259_), .A1(new_n2255_), .B0(new_n2263_), .Y(new_n2264_));
  AOI21X1  g01262(.A0(new_n2264_), .A1(new_n2221_), .B0(new_n2254_), .Y(new_n2265_));
  INVX1    g01263(.A(\A[836] ), .Y(new_n2266_));
  OR2X1    g01264(.A(new_n2266_), .B(\A[835] ), .Y(new_n2267_));
  INVX1    g01265(.A(\A[837] ), .Y(new_n2268_));
  AOI21X1  g01266(.A0(new_n2266_), .A1(\A[835] ), .B0(new_n2268_), .Y(new_n2269_));
  XOR2X1   g01267(.A(\A[836] ), .B(\A[835] ), .Y(new_n2270_));
  AND2X1   g01268(.A(new_n2270_), .B(new_n2268_), .Y(new_n2271_));
  AOI21X1  g01269(.A0(new_n2269_), .A1(new_n2267_), .B0(new_n2271_), .Y(new_n2272_));
  INVX1    g01270(.A(\A[840] ), .Y(new_n2273_));
  INVX1    g01271(.A(\A[839] ), .Y(new_n2274_));
  OR2X1    g01272(.A(new_n2274_), .B(\A[838] ), .Y(new_n2275_));
  AOI21X1  g01273(.A0(new_n2274_), .A1(\A[838] ), .B0(new_n2273_), .Y(new_n2276_));
  XOR2X1   g01274(.A(\A[839] ), .B(\A[838] ), .Y(new_n2277_));
  AOI22X1  g01275(.A0(new_n2277_), .A1(new_n2273_), .B0(new_n2276_), .B1(new_n2275_), .Y(new_n2278_));
  NOR2X1   g01276(.A(new_n2278_), .B(new_n2272_), .Y(new_n2279_));
  AND2X1   g01277(.A(\A[839] ), .B(\A[838] ), .Y(new_n2280_));
  AND2X1   g01278(.A(new_n2277_), .B(\A[840] ), .Y(new_n2281_));
  OR2X1    g01279(.A(new_n2281_), .B(new_n2280_), .Y(new_n2282_));
  AND2X1   g01280(.A(\A[836] ), .B(\A[835] ), .Y(new_n2283_));
  AOI21X1  g01281(.A0(new_n2270_), .A1(\A[837] ), .B0(new_n2283_), .Y(new_n2284_));
  XOR2X1   g01282(.A(new_n2284_), .B(new_n2282_), .Y(new_n2285_));
  XOR2X1   g01283(.A(new_n2285_), .B(new_n2279_), .Y(new_n2286_));
  XOR2X1   g01284(.A(new_n2278_), .B(new_n2272_), .Y(new_n2287_));
  OR2X1    g01285(.A(new_n2278_), .B(new_n2272_), .Y(new_n2288_));
  AOI21X1  g01286(.A0(new_n2277_), .A1(\A[840] ), .B0(new_n2280_), .Y(new_n2289_));
  OR2X1    g01287(.A(new_n2284_), .B(new_n2289_), .Y(new_n2290_));
  OAI21X1  g01288(.A0(new_n2285_), .A1(new_n2288_), .B0(new_n2290_), .Y(new_n2291_));
  AND2X1   g01289(.A(new_n2291_), .B(new_n2287_), .Y(new_n2292_));
  OR2X1    g01290(.A(new_n2292_), .B(new_n2286_), .Y(new_n2293_));
  AND2X1   g01291(.A(\A[845] ), .B(\A[844] ), .Y(new_n2294_));
  XOR2X1   g01292(.A(\A[845] ), .B(\A[844] ), .Y(new_n2295_));
  AOI21X1  g01293(.A0(new_n2295_), .A1(\A[846] ), .B0(new_n2294_), .Y(new_n2296_));
  AND2X1   g01294(.A(\A[842] ), .B(\A[841] ), .Y(new_n2297_));
  XOR2X1   g01295(.A(\A[842] ), .B(\A[841] ), .Y(new_n2298_));
  AOI21X1  g01296(.A0(new_n2298_), .A1(\A[843] ), .B0(new_n2297_), .Y(new_n2299_));
  INVX1    g01297(.A(\A[842] ), .Y(new_n2300_));
  OR2X1    g01298(.A(new_n2300_), .B(\A[841] ), .Y(new_n2301_));
  INVX1    g01299(.A(\A[843] ), .Y(new_n2302_));
  AOI21X1  g01300(.A0(new_n2300_), .A1(\A[841] ), .B0(new_n2302_), .Y(new_n2303_));
  AND2X1   g01301(.A(new_n2298_), .B(new_n2302_), .Y(new_n2304_));
  AOI21X1  g01302(.A0(new_n2303_), .A1(new_n2301_), .B0(new_n2304_), .Y(new_n2305_));
  INVX1    g01303(.A(\A[846] ), .Y(new_n2306_));
  INVX1    g01304(.A(\A[845] ), .Y(new_n2307_));
  OR2X1    g01305(.A(new_n2307_), .B(\A[844] ), .Y(new_n2308_));
  AOI21X1  g01306(.A0(new_n2307_), .A1(\A[844] ), .B0(new_n2306_), .Y(new_n2309_));
  AOI22X1  g01307(.A0(new_n2309_), .A1(new_n2308_), .B0(new_n2295_), .B1(new_n2306_), .Y(new_n2310_));
  OR4X1    g01308(.A(new_n2310_), .B(new_n2305_), .C(new_n2299_), .D(new_n2296_), .Y(new_n2311_));
  OR4X1    g01309(.A(new_n2284_), .B(new_n2289_), .C(new_n2278_), .D(new_n2272_), .Y(new_n2312_));
  XOR2X1   g01310(.A(new_n2310_), .B(new_n2305_), .Y(new_n2313_));
  NAND4X1  g01311(.A(new_n2313_), .B(new_n2312_), .C(new_n2311_), .D(new_n2287_), .Y(new_n2314_));
  XOR2X1   g01312(.A(new_n2299_), .B(new_n2296_), .Y(new_n2315_));
  NOR2X1   g01313(.A(new_n2310_), .B(new_n2305_), .Y(new_n2316_));
  NOR2X1   g01314(.A(new_n2299_), .B(new_n2296_), .Y(new_n2317_));
  AOI21X1  g01315(.A0(new_n2316_), .A1(new_n2315_), .B0(new_n2317_), .Y(new_n2318_));
  XOR2X1   g01316(.A(new_n2316_), .B(new_n2315_), .Y(new_n2319_));
  AND2X1   g01317(.A(new_n2303_), .B(new_n2301_), .Y(new_n2320_));
  OR2X1    g01318(.A(new_n2304_), .B(new_n2320_), .Y(new_n2321_));
  XOR2X1   g01319(.A(new_n2310_), .B(new_n2321_), .Y(new_n2322_));
  OAI21X1  g01320(.A0(new_n2322_), .A1(new_n2318_), .B0(new_n2319_), .Y(new_n2323_));
  XOR2X1   g01321(.A(new_n2323_), .B(new_n2314_), .Y(new_n2324_));
  AND2X1   g01322(.A(new_n2324_), .B(new_n2293_), .Y(new_n2325_));
  AND2X1   g01323(.A(new_n2269_), .B(new_n2267_), .Y(new_n2326_));
  OR2X1    g01324(.A(new_n2271_), .B(new_n2326_), .Y(new_n2327_));
  XOR2X1   g01325(.A(new_n2278_), .B(new_n2327_), .Y(new_n2328_));
  OR2X1    g01326(.A(new_n2310_), .B(new_n2305_), .Y(new_n2329_));
  XOR2X1   g01327(.A(new_n2329_), .B(new_n2315_), .Y(new_n2330_));
  NOR4X1   g01328(.A(new_n2284_), .B(new_n2289_), .C(new_n2278_), .D(new_n2272_), .Y(new_n2331_));
  NOR4X1   g01329(.A(new_n2322_), .B(new_n2331_), .C(new_n2330_), .D(new_n2328_), .Y(new_n2332_));
  AND2X1   g01330(.A(new_n2316_), .B(new_n2315_), .Y(new_n2333_));
  OAI22X1  g01331(.A0(new_n2313_), .A1(new_n2319_), .B0(new_n2317_), .B1(new_n2333_), .Y(new_n2334_));
  AOI22X1  g01332(.A0(new_n2334_), .A1(new_n2332_), .B0(new_n2323_), .B1(new_n2314_), .Y(new_n2335_));
  NAND2X1  g01333(.A(new_n2313_), .B(new_n2311_), .Y(new_n2336_));
  XOR2X1   g01334(.A(new_n2278_), .B(new_n2272_), .Y(new_n2337_));
  XOR2X1   g01335(.A(new_n2337_), .B(new_n2336_), .Y(new_n2338_));
  NAND2X1  g01336(.A(new_n2242_), .B(new_n2240_), .Y(new_n2339_));
  XOR2X1   g01337(.A(new_n2207_), .B(new_n2201_), .Y(new_n2340_));
  XOR2X1   g01338(.A(new_n2340_), .B(new_n2339_), .Y(new_n2341_));
  NOR2X1   g01339(.A(new_n2341_), .B(new_n2338_), .Y(new_n2342_));
  OAI21X1  g01340(.A0(new_n2335_), .A1(new_n2293_), .B0(new_n2342_), .Y(new_n2343_));
  NOR2X1   g01341(.A(new_n2343_), .B(new_n2325_), .Y(new_n2344_));
  NAND2X1  g01342(.A(new_n2324_), .B(new_n2293_), .Y(new_n2345_));
  OR2X1    g01343(.A(new_n2335_), .B(new_n2293_), .Y(new_n2346_));
  AOI21X1  g01344(.A0(new_n2346_), .A1(new_n2345_), .B0(new_n2342_), .Y(new_n2347_));
  OAI21X1  g01345(.A0(new_n2347_), .A1(new_n2344_), .B0(new_n2265_), .Y(new_n2348_));
  MX2X1    g01346(.A(new_n2264_), .B(new_n2253_), .S0(new_n2222_), .Y(new_n2349_));
  OR2X1    g01347(.A(new_n2341_), .B(new_n2338_), .Y(new_n2350_));
  OAI21X1  g01348(.A0(new_n2335_), .A1(new_n2293_), .B0(new_n2350_), .Y(new_n2351_));
  NOR2X1   g01349(.A(new_n2351_), .B(new_n2325_), .Y(new_n2352_));
  AOI21X1  g01350(.A0(new_n2346_), .A1(new_n2345_), .B0(new_n2350_), .Y(new_n2353_));
  OAI21X1  g01351(.A0(new_n2353_), .A1(new_n2352_), .B0(new_n2349_), .Y(new_n2354_));
  XOR2X1   g01352(.A(new_n2341_), .B(new_n2338_), .Y(new_n2355_));
  INVX1    g01353(.A(new_n2355_), .Y(new_n2356_));
  INVX1    g01354(.A(new_n2149_), .Y(new_n2357_));
  XOR2X1   g01355(.A(new_n2357_), .B(new_n2111_), .Y(new_n2358_));
  NOR2X1   g01356(.A(new_n2358_), .B(new_n2356_), .Y(new_n2359_));
  NAND3X1  g01357(.A(new_n2359_), .B(new_n2354_), .C(new_n2348_), .Y(new_n2360_));
  OR2X1    g01358(.A(new_n2343_), .B(new_n2325_), .Y(new_n2361_));
  NOR2X1   g01359(.A(new_n2335_), .B(new_n2293_), .Y(new_n2362_));
  OAI21X1  g01360(.A0(new_n2362_), .A1(new_n2325_), .B0(new_n2350_), .Y(new_n2363_));
  AOI21X1  g01361(.A0(new_n2363_), .A1(new_n2361_), .B0(new_n2349_), .Y(new_n2364_));
  OR2X1    g01362(.A(new_n2351_), .B(new_n2325_), .Y(new_n2365_));
  OAI21X1  g01363(.A0(new_n2362_), .A1(new_n2325_), .B0(new_n2342_), .Y(new_n2366_));
  AOI21X1  g01364(.A0(new_n2366_), .A1(new_n2365_), .B0(new_n2265_), .Y(new_n2367_));
  OR2X1    g01365(.A(new_n2358_), .B(new_n2356_), .Y(new_n2368_));
  OAI21X1  g01366(.A0(new_n2367_), .A1(new_n2364_), .B0(new_n2368_), .Y(new_n2369_));
  AOI21X1  g01367(.A0(new_n2369_), .A1(new_n2360_), .B0(new_n2194_), .Y(new_n2370_));
  AOI21X1  g01368(.A0(new_n2192_), .A1(new_n2191_), .B0(new_n2188_), .Y(new_n2371_));
  AOI21X1  g01369(.A0(new_n2188_), .A1(new_n2155_), .B0(new_n2371_), .Y(new_n2372_));
  NAND3X1  g01370(.A(new_n2368_), .B(new_n2354_), .C(new_n2348_), .Y(new_n2373_));
  OAI21X1  g01371(.A0(new_n2367_), .A1(new_n2364_), .B0(new_n2359_), .Y(new_n2374_));
  AOI21X1  g01372(.A0(new_n2374_), .A1(new_n2373_), .B0(new_n2372_), .Y(new_n2375_));
  XOR2X1   g01373(.A(new_n2358_), .B(new_n2355_), .Y(new_n2376_));
  XOR2X1   g01374(.A(new_n1933_), .B(new_n1856_), .Y(new_n2377_));
  NOR2X1   g01375(.A(new_n2377_), .B(new_n2376_), .Y(new_n2378_));
  INVX1    g01376(.A(new_n2378_), .Y(new_n2379_));
  NOR3X1   g01377(.A(new_n2379_), .B(new_n2375_), .C(new_n2370_), .Y(new_n2380_));
  NOR3X1   g01378(.A(new_n2368_), .B(new_n2367_), .C(new_n2364_), .Y(new_n2381_));
  AOI21X1  g01379(.A0(new_n2354_), .A1(new_n2348_), .B0(new_n2359_), .Y(new_n2382_));
  OAI21X1  g01380(.A0(new_n2382_), .A1(new_n2381_), .B0(new_n2372_), .Y(new_n2383_));
  NOR3X1   g01381(.A(new_n2359_), .B(new_n2367_), .C(new_n2364_), .Y(new_n2384_));
  AOI21X1  g01382(.A0(new_n2354_), .A1(new_n2348_), .B0(new_n2368_), .Y(new_n2385_));
  OAI21X1  g01383(.A0(new_n2385_), .A1(new_n2384_), .B0(new_n2194_), .Y(new_n2386_));
  AOI21X1  g01384(.A0(new_n2386_), .A1(new_n2383_), .B0(new_n2378_), .Y(new_n2387_));
  OAI21X1  g01385(.A0(new_n2387_), .A1(new_n2380_), .B0(new_n2038_), .Y(new_n2388_));
  OR2X1    g01386(.A(new_n2033_), .B(new_n2027_), .Y(new_n2389_));
  NOR3X1   g01387(.A(new_n1934_), .B(new_n1942_), .C(new_n1939_), .Y(new_n2390_));
  AOI21X1  g01388(.A0(new_n1855_), .A1(new_n1849_), .B0(new_n1943_), .Y(new_n2391_));
  OAI21X1  g01389(.A0(new_n2391_), .A1(new_n2390_), .B0(new_n2389_), .Y(new_n2392_));
  OAI21X1  g01390(.A0(new_n2389_), .A1(new_n1945_), .B0(new_n2392_), .Y(new_n2393_));
  NOR3X1   g01391(.A(new_n2378_), .B(new_n2375_), .C(new_n2370_), .Y(new_n2394_));
  AOI21X1  g01392(.A0(new_n2386_), .A1(new_n2383_), .B0(new_n2379_), .Y(new_n2395_));
  OAI21X1  g01393(.A0(new_n2395_), .A1(new_n2394_), .B0(new_n2393_), .Y(new_n2396_));
  XOR2X1   g01394(.A(new_n1933_), .B(new_n1857_), .Y(new_n2397_));
  XOR2X1   g01395(.A(new_n2397_), .B(new_n2376_), .Y(new_n2398_));
  XOR2X1   g01396(.A(new_n1591_), .B(new_n1416_), .Y(new_n2399_));
  XOR2X1   g01397(.A(new_n2399_), .B(new_n1340_), .Y(new_n2400_));
  NOR2X1   g01398(.A(new_n2400_), .B(new_n2398_), .Y(new_n2401_));
  NAND3X1  g01399(.A(new_n2401_), .B(new_n2396_), .C(new_n2388_), .Y(new_n2402_));
  NAND3X1  g01400(.A(new_n2378_), .B(new_n2386_), .C(new_n2383_), .Y(new_n2403_));
  OAI21X1  g01401(.A0(new_n2375_), .A1(new_n2370_), .B0(new_n2379_), .Y(new_n2404_));
  AOI21X1  g01402(.A0(new_n2404_), .A1(new_n2403_), .B0(new_n2393_), .Y(new_n2405_));
  NAND3X1  g01403(.A(new_n2379_), .B(new_n2386_), .C(new_n2383_), .Y(new_n2406_));
  OAI21X1  g01404(.A0(new_n2375_), .A1(new_n2370_), .B0(new_n2378_), .Y(new_n2407_));
  AOI21X1  g01405(.A0(new_n2407_), .A1(new_n2406_), .B0(new_n2038_), .Y(new_n2408_));
  INVX1    g01406(.A(new_n2401_), .Y(new_n2409_));
  OAI21X1  g01407(.A0(new_n2408_), .A1(new_n2405_), .B0(new_n2409_), .Y(new_n2410_));
  AOI21X1  g01408(.A0(new_n2410_), .A1(new_n2402_), .B0(new_n1695_), .Y(new_n2411_));
  NOR2X1   g01409(.A(new_n1686_), .B(new_n1680_), .Y(new_n2412_));
  NAND3X1  g01410(.A(new_n1600_), .B(new_n1590_), .C(new_n1586_), .Y(new_n2413_));
  OAI21X1  g01411(.A0(new_n1599_), .A1(new_n1596_), .B0(new_n1592_), .Y(new_n2414_));
  AND2X1   g01412(.A(new_n2414_), .B(new_n2413_), .Y(new_n2415_));
  MX2X1    g01413(.A(new_n2415_), .B(new_n1602_), .S0(new_n2412_), .Y(new_n2416_));
  NAND3X1  g01414(.A(new_n1503_), .B(new_n1339_), .C(new_n1334_), .Y(new_n2417_));
  OAI21X1  g01415(.A0(new_n1502_), .A1(new_n1499_), .B0(new_n1495_), .Y(new_n2418_));
  AND2X1   g01416(.A(new_n2418_), .B(new_n2417_), .Y(new_n2419_));
  MX2X1    g01417(.A(new_n2419_), .B(new_n1505_), .S0(new_n2416_), .Y(new_n2420_));
  NAND3X1  g01418(.A(new_n2409_), .B(new_n2396_), .C(new_n2388_), .Y(new_n2421_));
  OAI21X1  g01419(.A0(new_n2408_), .A1(new_n2405_), .B0(new_n2401_), .Y(new_n2422_));
  AOI21X1  g01420(.A0(new_n2422_), .A1(new_n2421_), .B0(new_n2420_), .Y(new_n2423_));
  INVX1    g01421(.A(\A[469] ), .Y(new_n2424_));
  OR2X1    g01422(.A(\A[470] ), .B(new_n2424_), .Y(new_n2425_));
  INVX1    g01423(.A(\A[471] ), .Y(new_n2426_));
  AOI21X1  g01424(.A0(\A[470] ), .A1(new_n2424_), .B0(new_n2426_), .Y(new_n2427_));
  XOR2X1   g01425(.A(\A[470] ), .B(\A[469] ), .Y(new_n2428_));
  AND2X1   g01426(.A(new_n2428_), .B(new_n2426_), .Y(new_n2429_));
  AOI21X1  g01427(.A0(new_n2427_), .A1(new_n2425_), .B0(new_n2429_), .Y(new_n2430_));
  INVX1    g01428(.A(\A[474] ), .Y(new_n2431_));
  INVX1    g01429(.A(\A[472] ), .Y(new_n2432_));
  OR2X1    g01430(.A(\A[473] ), .B(new_n2432_), .Y(new_n2433_));
  AOI21X1  g01431(.A0(\A[473] ), .A1(new_n2432_), .B0(new_n2431_), .Y(new_n2434_));
  XOR2X1   g01432(.A(\A[473] ), .B(\A[472] ), .Y(new_n2435_));
  AOI22X1  g01433(.A0(new_n2435_), .A1(new_n2431_), .B0(new_n2434_), .B1(new_n2433_), .Y(new_n2436_));
  AND2X1   g01434(.A(\A[473] ), .B(\A[472] ), .Y(new_n2437_));
  AOI21X1  g01435(.A0(new_n2435_), .A1(\A[474] ), .B0(new_n2437_), .Y(new_n2438_));
  AND2X1   g01436(.A(\A[470] ), .B(\A[469] ), .Y(new_n2439_));
  AOI21X1  g01437(.A0(new_n2428_), .A1(\A[471] ), .B0(new_n2439_), .Y(new_n2440_));
  XOR2X1   g01438(.A(new_n2436_), .B(new_n2430_), .Y(new_n2441_));
  INVX1    g01439(.A(\A[466] ), .Y(new_n2442_));
  OR2X1    g01440(.A(\A[467] ), .B(new_n2442_), .Y(new_n2443_));
  INVX1    g01441(.A(\A[468] ), .Y(new_n2444_));
  AOI21X1  g01442(.A0(\A[467] ), .A1(new_n2442_), .B0(new_n2444_), .Y(new_n2445_));
  XOR2X1   g01443(.A(\A[467] ), .B(\A[466] ), .Y(new_n2446_));
  AND2X1   g01444(.A(new_n2446_), .B(new_n2444_), .Y(new_n2447_));
  AOI21X1  g01445(.A0(new_n2445_), .A1(new_n2443_), .B0(new_n2447_), .Y(new_n2448_));
  INVX1    g01446(.A(\A[465] ), .Y(new_n2449_));
  INVX1    g01447(.A(\A[463] ), .Y(new_n2450_));
  OR2X1    g01448(.A(\A[464] ), .B(new_n2450_), .Y(new_n2451_));
  AOI21X1  g01449(.A0(\A[464] ), .A1(new_n2450_), .B0(new_n2449_), .Y(new_n2452_));
  XOR2X1   g01450(.A(\A[464] ), .B(\A[463] ), .Y(new_n2453_));
  AOI22X1  g01451(.A0(new_n2453_), .A1(new_n2449_), .B0(new_n2452_), .B1(new_n2451_), .Y(new_n2454_));
  AND2X1   g01452(.A(\A[467] ), .B(\A[466] ), .Y(new_n2455_));
  AOI21X1  g01453(.A0(new_n2446_), .A1(\A[468] ), .B0(new_n2455_), .Y(new_n2456_));
  AND2X1   g01454(.A(\A[464] ), .B(\A[463] ), .Y(new_n2457_));
  AOI21X1  g01455(.A0(new_n2453_), .A1(\A[465] ), .B0(new_n2457_), .Y(new_n2458_));
  XOR2X1   g01456(.A(new_n2454_), .B(new_n2448_), .Y(new_n2459_));
  XOR2X1   g01457(.A(new_n2459_), .B(new_n2441_), .Y(new_n2460_));
  INVX1    g01458(.A(\A[481] ), .Y(new_n2461_));
  OR2X1    g01459(.A(\A[482] ), .B(new_n2461_), .Y(new_n2462_));
  INVX1    g01460(.A(\A[483] ), .Y(new_n2463_));
  AOI21X1  g01461(.A0(\A[482] ), .A1(new_n2461_), .B0(new_n2463_), .Y(new_n2464_));
  AND2X1   g01462(.A(new_n2464_), .B(new_n2462_), .Y(new_n2465_));
  XOR2X1   g01463(.A(\A[482] ), .B(\A[481] ), .Y(new_n2466_));
  AND2X1   g01464(.A(new_n2466_), .B(new_n2463_), .Y(new_n2467_));
  OR2X1    g01465(.A(new_n2467_), .B(new_n2465_), .Y(new_n2468_));
  INVX1    g01466(.A(\A[486] ), .Y(new_n2469_));
  INVX1    g01467(.A(\A[484] ), .Y(new_n2470_));
  OR2X1    g01468(.A(\A[485] ), .B(new_n2470_), .Y(new_n2471_));
  AOI21X1  g01469(.A0(\A[485] ), .A1(new_n2470_), .B0(new_n2469_), .Y(new_n2472_));
  XOR2X1   g01470(.A(\A[485] ), .B(\A[484] ), .Y(new_n2473_));
  AOI22X1  g01471(.A0(new_n2473_), .A1(new_n2469_), .B0(new_n2472_), .B1(new_n2471_), .Y(new_n2474_));
  AND2X1   g01472(.A(\A[485] ), .B(\A[484] ), .Y(new_n2475_));
  AOI21X1  g01473(.A0(new_n2473_), .A1(\A[486] ), .B0(new_n2475_), .Y(new_n2476_));
  AND2X1   g01474(.A(\A[482] ), .B(\A[481] ), .Y(new_n2477_));
  AOI21X1  g01475(.A0(new_n2466_), .A1(\A[483] ), .B0(new_n2477_), .Y(new_n2478_));
  XOR2X1   g01476(.A(new_n2474_), .B(new_n2468_), .Y(new_n2479_));
  INVX1    g01477(.A(\A[475] ), .Y(new_n2480_));
  OR2X1    g01478(.A(\A[476] ), .B(new_n2480_), .Y(new_n2481_));
  INVX1    g01479(.A(\A[477] ), .Y(new_n2482_));
  AOI21X1  g01480(.A0(\A[476] ), .A1(new_n2480_), .B0(new_n2482_), .Y(new_n2483_));
  XOR2X1   g01481(.A(\A[476] ), .B(\A[475] ), .Y(new_n2484_));
  AND2X1   g01482(.A(new_n2484_), .B(new_n2482_), .Y(new_n2485_));
  AOI21X1  g01483(.A0(new_n2483_), .A1(new_n2481_), .B0(new_n2485_), .Y(new_n2486_));
  INVX1    g01484(.A(\A[480] ), .Y(new_n2487_));
  INVX1    g01485(.A(\A[478] ), .Y(new_n2488_));
  OR2X1    g01486(.A(\A[479] ), .B(new_n2488_), .Y(new_n2489_));
  AOI21X1  g01487(.A0(\A[479] ), .A1(new_n2488_), .B0(new_n2487_), .Y(new_n2490_));
  XOR2X1   g01488(.A(\A[479] ), .B(\A[478] ), .Y(new_n2491_));
  AOI22X1  g01489(.A0(new_n2491_), .A1(new_n2487_), .B0(new_n2490_), .B1(new_n2489_), .Y(new_n2492_));
  AND2X1   g01490(.A(\A[479] ), .B(\A[478] ), .Y(new_n2493_));
  AOI21X1  g01491(.A0(new_n2491_), .A1(\A[480] ), .B0(new_n2493_), .Y(new_n2494_));
  AND2X1   g01492(.A(\A[476] ), .B(\A[475] ), .Y(new_n2495_));
  AOI21X1  g01493(.A0(new_n2484_), .A1(\A[477] ), .B0(new_n2495_), .Y(new_n2496_));
  XOR2X1   g01494(.A(new_n2492_), .B(new_n2486_), .Y(new_n2497_));
  XOR2X1   g01495(.A(new_n2497_), .B(new_n2479_), .Y(new_n2498_));
  XOR2X1   g01496(.A(new_n2498_), .B(new_n2460_), .Y(new_n2499_));
  INVX1    g01497(.A(\A[505] ), .Y(new_n2500_));
  OR2X1    g01498(.A(\A[506] ), .B(new_n2500_), .Y(new_n2501_));
  INVX1    g01499(.A(\A[507] ), .Y(new_n2502_));
  AOI21X1  g01500(.A0(\A[506] ), .A1(new_n2500_), .B0(new_n2502_), .Y(new_n2503_));
  XOR2X1   g01501(.A(\A[506] ), .B(\A[505] ), .Y(new_n2504_));
  AND2X1   g01502(.A(new_n2504_), .B(new_n2502_), .Y(new_n2505_));
  AOI21X1  g01503(.A0(new_n2503_), .A1(new_n2501_), .B0(new_n2505_), .Y(new_n2506_));
  INVX1    g01504(.A(\A[510] ), .Y(new_n2507_));
  INVX1    g01505(.A(\A[508] ), .Y(new_n2508_));
  OR2X1    g01506(.A(\A[509] ), .B(new_n2508_), .Y(new_n2509_));
  AOI21X1  g01507(.A0(\A[509] ), .A1(new_n2508_), .B0(new_n2507_), .Y(new_n2510_));
  XOR2X1   g01508(.A(\A[509] ), .B(\A[508] ), .Y(new_n2511_));
  AOI22X1  g01509(.A0(new_n2511_), .A1(new_n2507_), .B0(new_n2510_), .B1(new_n2509_), .Y(new_n2512_));
  AND2X1   g01510(.A(\A[509] ), .B(\A[508] ), .Y(new_n2513_));
  AOI21X1  g01511(.A0(new_n2511_), .A1(\A[510] ), .B0(new_n2513_), .Y(new_n2514_));
  AND2X1   g01512(.A(\A[506] ), .B(\A[505] ), .Y(new_n2515_));
  AOI21X1  g01513(.A0(new_n2504_), .A1(\A[507] ), .B0(new_n2515_), .Y(new_n2516_));
  XOR2X1   g01514(.A(new_n2512_), .B(new_n2506_), .Y(new_n2517_));
  INVX1    g01515(.A(\A[499] ), .Y(new_n2518_));
  OR2X1    g01516(.A(\A[500] ), .B(new_n2518_), .Y(new_n2519_));
  INVX1    g01517(.A(\A[501] ), .Y(new_n2520_));
  AOI21X1  g01518(.A0(\A[500] ), .A1(new_n2518_), .B0(new_n2520_), .Y(new_n2521_));
  XOR2X1   g01519(.A(\A[500] ), .B(\A[499] ), .Y(new_n2522_));
  AND2X1   g01520(.A(new_n2522_), .B(new_n2520_), .Y(new_n2523_));
  AOI21X1  g01521(.A0(new_n2521_), .A1(new_n2519_), .B0(new_n2523_), .Y(new_n2524_));
  INVX1    g01522(.A(\A[504] ), .Y(new_n2525_));
  INVX1    g01523(.A(\A[502] ), .Y(new_n2526_));
  OR2X1    g01524(.A(\A[503] ), .B(new_n2526_), .Y(new_n2527_));
  AOI21X1  g01525(.A0(\A[503] ), .A1(new_n2526_), .B0(new_n2525_), .Y(new_n2528_));
  XOR2X1   g01526(.A(\A[503] ), .B(\A[502] ), .Y(new_n2529_));
  AOI22X1  g01527(.A0(new_n2529_), .A1(new_n2525_), .B0(new_n2528_), .B1(new_n2527_), .Y(new_n2530_));
  AND2X1   g01528(.A(\A[503] ), .B(\A[502] ), .Y(new_n2531_));
  AOI21X1  g01529(.A0(new_n2529_), .A1(\A[504] ), .B0(new_n2531_), .Y(new_n2532_));
  AND2X1   g01530(.A(\A[500] ), .B(\A[499] ), .Y(new_n2533_));
  AOI21X1  g01531(.A0(new_n2522_), .A1(\A[501] ), .B0(new_n2533_), .Y(new_n2534_));
  XOR2X1   g01532(.A(new_n2530_), .B(new_n2524_), .Y(new_n2535_));
  XOR2X1   g01533(.A(new_n2535_), .B(new_n2517_), .Y(new_n2536_));
  INVX1    g01534(.A(new_n2536_), .Y(new_n2537_));
  INVX1    g01535(.A(\A[493] ), .Y(new_n2538_));
  OR2X1    g01536(.A(\A[494] ), .B(new_n2538_), .Y(new_n2539_));
  INVX1    g01537(.A(\A[495] ), .Y(new_n2540_));
  AOI21X1  g01538(.A0(\A[494] ), .A1(new_n2538_), .B0(new_n2540_), .Y(new_n2541_));
  AND2X1   g01539(.A(new_n2541_), .B(new_n2539_), .Y(new_n2542_));
  XOR2X1   g01540(.A(\A[494] ), .B(\A[493] ), .Y(new_n2543_));
  AND2X1   g01541(.A(new_n2543_), .B(new_n2540_), .Y(new_n2544_));
  OR2X1    g01542(.A(new_n2544_), .B(new_n2542_), .Y(new_n2545_));
  INVX1    g01543(.A(\A[498] ), .Y(new_n2546_));
  INVX1    g01544(.A(\A[496] ), .Y(new_n2547_));
  OR2X1    g01545(.A(\A[497] ), .B(new_n2547_), .Y(new_n2548_));
  AOI21X1  g01546(.A0(\A[497] ), .A1(new_n2547_), .B0(new_n2546_), .Y(new_n2549_));
  XOR2X1   g01547(.A(\A[497] ), .B(\A[496] ), .Y(new_n2550_));
  AOI22X1  g01548(.A0(new_n2550_), .A1(new_n2546_), .B0(new_n2549_), .B1(new_n2548_), .Y(new_n2551_));
  AND2X1   g01549(.A(\A[497] ), .B(\A[496] ), .Y(new_n2552_));
  AOI21X1  g01550(.A0(new_n2550_), .A1(\A[498] ), .B0(new_n2552_), .Y(new_n2553_));
  AND2X1   g01551(.A(\A[494] ), .B(\A[493] ), .Y(new_n2554_));
  AOI21X1  g01552(.A0(new_n2543_), .A1(\A[495] ), .B0(new_n2554_), .Y(new_n2555_));
  XOR2X1   g01553(.A(new_n2551_), .B(new_n2545_), .Y(new_n2556_));
  INVX1    g01554(.A(\A[487] ), .Y(new_n2557_));
  OR2X1    g01555(.A(\A[488] ), .B(new_n2557_), .Y(new_n2558_));
  INVX1    g01556(.A(\A[489] ), .Y(new_n2559_));
  AOI21X1  g01557(.A0(\A[488] ), .A1(new_n2557_), .B0(new_n2559_), .Y(new_n2560_));
  XOR2X1   g01558(.A(\A[488] ), .B(\A[487] ), .Y(new_n2561_));
  AND2X1   g01559(.A(new_n2561_), .B(new_n2559_), .Y(new_n2562_));
  AOI21X1  g01560(.A0(new_n2560_), .A1(new_n2558_), .B0(new_n2562_), .Y(new_n2563_));
  INVX1    g01561(.A(\A[492] ), .Y(new_n2564_));
  INVX1    g01562(.A(\A[490] ), .Y(new_n2565_));
  OR2X1    g01563(.A(\A[491] ), .B(new_n2565_), .Y(new_n2566_));
  AOI21X1  g01564(.A0(\A[491] ), .A1(new_n2565_), .B0(new_n2564_), .Y(new_n2567_));
  XOR2X1   g01565(.A(\A[491] ), .B(\A[490] ), .Y(new_n2568_));
  AOI22X1  g01566(.A0(new_n2568_), .A1(new_n2564_), .B0(new_n2567_), .B1(new_n2566_), .Y(new_n2569_));
  AND2X1   g01567(.A(\A[491] ), .B(\A[490] ), .Y(new_n2570_));
  AOI21X1  g01568(.A0(new_n2568_), .A1(\A[492] ), .B0(new_n2570_), .Y(new_n2571_));
  AND2X1   g01569(.A(\A[488] ), .B(\A[487] ), .Y(new_n2572_));
  AOI21X1  g01570(.A0(new_n2561_), .A1(\A[489] ), .B0(new_n2572_), .Y(new_n2573_));
  XOR2X1   g01571(.A(new_n2569_), .B(new_n2563_), .Y(new_n2574_));
  XOR2X1   g01572(.A(new_n2574_), .B(new_n2556_), .Y(new_n2575_));
  XOR2X1   g01573(.A(new_n2575_), .B(new_n2537_), .Y(new_n2576_));
  XOR2X1   g01574(.A(new_n2576_), .B(new_n2499_), .Y(new_n2577_));
  INVX1    g01575(.A(\A[553] ), .Y(new_n2578_));
  OR2X1    g01576(.A(\A[554] ), .B(new_n2578_), .Y(new_n2579_));
  INVX1    g01577(.A(\A[555] ), .Y(new_n2580_));
  AOI21X1  g01578(.A0(\A[554] ), .A1(new_n2578_), .B0(new_n2580_), .Y(new_n2581_));
  XOR2X1   g01579(.A(\A[554] ), .B(\A[553] ), .Y(new_n2582_));
  AND2X1   g01580(.A(new_n2582_), .B(new_n2580_), .Y(new_n2583_));
  AOI21X1  g01581(.A0(new_n2581_), .A1(new_n2579_), .B0(new_n2583_), .Y(new_n2584_));
  INVX1    g01582(.A(\A[558] ), .Y(new_n2585_));
  INVX1    g01583(.A(\A[556] ), .Y(new_n2586_));
  OR2X1    g01584(.A(\A[557] ), .B(new_n2586_), .Y(new_n2587_));
  AOI21X1  g01585(.A0(\A[557] ), .A1(new_n2586_), .B0(new_n2585_), .Y(new_n2588_));
  XOR2X1   g01586(.A(\A[557] ), .B(\A[556] ), .Y(new_n2589_));
  AOI22X1  g01587(.A0(new_n2589_), .A1(new_n2585_), .B0(new_n2588_), .B1(new_n2587_), .Y(new_n2590_));
  AND2X1   g01588(.A(\A[557] ), .B(\A[556] ), .Y(new_n2591_));
  AOI21X1  g01589(.A0(new_n2589_), .A1(\A[558] ), .B0(new_n2591_), .Y(new_n2592_));
  AND2X1   g01590(.A(\A[554] ), .B(\A[553] ), .Y(new_n2593_));
  AOI21X1  g01591(.A0(new_n2582_), .A1(\A[555] ), .B0(new_n2593_), .Y(new_n2594_));
  XOR2X1   g01592(.A(new_n2590_), .B(new_n2584_), .Y(new_n2595_));
  INVX1    g01593(.A(\A[547] ), .Y(new_n2596_));
  OR2X1    g01594(.A(\A[548] ), .B(new_n2596_), .Y(new_n2597_));
  INVX1    g01595(.A(\A[549] ), .Y(new_n2598_));
  AOI21X1  g01596(.A0(\A[548] ), .A1(new_n2596_), .B0(new_n2598_), .Y(new_n2599_));
  XOR2X1   g01597(.A(\A[548] ), .B(\A[547] ), .Y(new_n2600_));
  AND2X1   g01598(.A(new_n2600_), .B(new_n2598_), .Y(new_n2601_));
  AOI21X1  g01599(.A0(new_n2599_), .A1(new_n2597_), .B0(new_n2601_), .Y(new_n2602_));
  INVX1    g01600(.A(\A[552] ), .Y(new_n2603_));
  INVX1    g01601(.A(\A[550] ), .Y(new_n2604_));
  OR2X1    g01602(.A(\A[551] ), .B(new_n2604_), .Y(new_n2605_));
  AOI21X1  g01603(.A0(\A[551] ), .A1(new_n2604_), .B0(new_n2603_), .Y(new_n2606_));
  XOR2X1   g01604(.A(\A[551] ), .B(\A[550] ), .Y(new_n2607_));
  AOI22X1  g01605(.A0(new_n2607_), .A1(new_n2603_), .B0(new_n2606_), .B1(new_n2605_), .Y(new_n2608_));
  AND2X1   g01606(.A(\A[551] ), .B(\A[550] ), .Y(new_n2609_));
  AOI21X1  g01607(.A0(new_n2607_), .A1(\A[552] ), .B0(new_n2609_), .Y(new_n2610_));
  AND2X1   g01608(.A(\A[548] ), .B(\A[547] ), .Y(new_n2611_));
  AOI21X1  g01609(.A0(new_n2600_), .A1(\A[549] ), .B0(new_n2611_), .Y(new_n2612_));
  XOR2X1   g01610(.A(new_n2608_), .B(new_n2602_), .Y(new_n2613_));
  XOR2X1   g01611(.A(new_n2613_), .B(new_n2595_), .Y(new_n2614_));
  INVX1    g01612(.A(\A[541] ), .Y(new_n2615_));
  OR2X1    g01613(.A(\A[542] ), .B(new_n2615_), .Y(new_n2616_));
  INVX1    g01614(.A(\A[543] ), .Y(new_n2617_));
  AOI21X1  g01615(.A0(\A[542] ), .A1(new_n2615_), .B0(new_n2617_), .Y(new_n2618_));
  AND2X1   g01616(.A(new_n2618_), .B(new_n2616_), .Y(new_n2619_));
  XOR2X1   g01617(.A(\A[542] ), .B(\A[541] ), .Y(new_n2620_));
  AND2X1   g01618(.A(new_n2620_), .B(new_n2617_), .Y(new_n2621_));
  OR2X1    g01619(.A(new_n2621_), .B(new_n2619_), .Y(new_n2622_));
  INVX1    g01620(.A(\A[546] ), .Y(new_n2623_));
  INVX1    g01621(.A(\A[544] ), .Y(new_n2624_));
  OR2X1    g01622(.A(\A[545] ), .B(new_n2624_), .Y(new_n2625_));
  AOI21X1  g01623(.A0(\A[545] ), .A1(new_n2624_), .B0(new_n2623_), .Y(new_n2626_));
  XOR2X1   g01624(.A(\A[545] ), .B(\A[544] ), .Y(new_n2627_));
  AOI22X1  g01625(.A0(new_n2627_), .A1(new_n2623_), .B0(new_n2626_), .B1(new_n2625_), .Y(new_n2628_));
  AND2X1   g01626(.A(\A[545] ), .B(\A[544] ), .Y(new_n2629_));
  AOI21X1  g01627(.A0(new_n2627_), .A1(\A[546] ), .B0(new_n2629_), .Y(new_n2630_));
  AND2X1   g01628(.A(\A[542] ), .B(\A[541] ), .Y(new_n2631_));
  AOI21X1  g01629(.A0(new_n2620_), .A1(\A[543] ), .B0(new_n2631_), .Y(new_n2632_));
  XOR2X1   g01630(.A(new_n2628_), .B(new_n2622_), .Y(new_n2633_));
  INVX1    g01631(.A(\A[535] ), .Y(new_n2634_));
  OR2X1    g01632(.A(\A[536] ), .B(new_n2634_), .Y(new_n2635_));
  INVX1    g01633(.A(\A[537] ), .Y(new_n2636_));
  AOI21X1  g01634(.A0(\A[536] ), .A1(new_n2634_), .B0(new_n2636_), .Y(new_n2637_));
  XOR2X1   g01635(.A(\A[536] ), .B(\A[535] ), .Y(new_n2638_));
  AND2X1   g01636(.A(new_n2638_), .B(new_n2636_), .Y(new_n2639_));
  AOI21X1  g01637(.A0(new_n2637_), .A1(new_n2635_), .B0(new_n2639_), .Y(new_n2640_));
  INVX1    g01638(.A(\A[540] ), .Y(new_n2641_));
  INVX1    g01639(.A(\A[538] ), .Y(new_n2642_));
  OR2X1    g01640(.A(\A[539] ), .B(new_n2642_), .Y(new_n2643_));
  AOI21X1  g01641(.A0(\A[539] ), .A1(new_n2642_), .B0(new_n2641_), .Y(new_n2644_));
  XOR2X1   g01642(.A(\A[539] ), .B(\A[538] ), .Y(new_n2645_));
  AOI22X1  g01643(.A0(new_n2645_), .A1(new_n2641_), .B0(new_n2644_), .B1(new_n2643_), .Y(new_n2646_));
  AND2X1   g01644(.A(\A[539] ), .B(\A[538] ), .Y(new_n2647_));
  AOI21X1  g01645(.A0(new_n2645_), .A1(\A[540] ), .B0(new_n2647_), .Y(new_n2648_));
  AND2X1   g01646(.A(\A[536] ), .B(\A[535] ), .Y(new_n2649_));
  AOI21X1  g01647(.A0(new_n2638_), .A1(\A[537] ), .B0(new_n2649_), .Y(new_n2650_));
  XOR2X1   g01648(.A(new_n2646_), .B(new_n2640_), .Y(new_n2651_));
  XOR2X1   g01649(.A(new_n2651_), .B(new_n2633_), .Y(new_n2652_));
  XOR2X1   g01650(.A(new_n2652_), .B(new_n2614_), .Y(new_n2653_));
  INVX1    g01651(.A(\A[529] ), .Y(new_n2654_));
  OR2X1    g01652(.A(\A[530] ), .B(new_n2654_), .Y(new_n2655_));
  INVX1    g01653(.A(\A[531] ), .Y(new_n2656_));
  AOI21X1  g01654(.A0(\A[530] ), .A1(new_n2654_), .B0(new_n2656_), .Y(new_n2657_));
  XOR2X1   g01655(.A(\A[530] ), .B(\A[529] ), .Y(new_n2658_));
  AND2X1   g01656(.A(new_n2658_), .B(new_n2656_), .Y(new_n2659_));
  AOI21X1  g01657(.A0(new_n2657_), .A1(new_n2655_), .B0(new_n2659_), .Y(new_n2660_));
  INVX1    g01658(.A(\A[534] ), .Y(new_n2661_));
  INVX1    g01659(.A(\A[532] ), .Y(new_n2662_));
  OR2X1    g01660(.A(\A[533] ), .B(new_n2662_), .Y(new_n2663_));
  AOI21X1  g01661(.A0(\A[533] ), .A1(new_n2662_), .B0(new_n2661_), .Y(new_n2664_));
  XOR2X1   g01662(.A(\A[533] ), .B(\A[532] ), .Y(new_n2665_));
  AOI22X1  g01663(.A0(new_n2665_), .A1(new_n2661_), .B0(new_n2664_), .B1(new_n2663_), .Y(new_n2666_));
  AND2X1   g01664(.A(\A[533] ), .B(\A[532] ), .Y(new_n2667_));
  AOI21X1  g01665(.A0(new_n2665_), .A1(\A[534] ), .B0(new_n2667_), .Y(new_n2668_));
  AND2X1   g01666(.A(\A[530] ), .B(\A[529] ), .Y(new_n2669_));
  AOI21X1  g01667(.A0(new_n2658_), .A1(\A[531] ), .B0(new_n2669_), .Y(new_n2670_));
  XOR2X1   g01668(.A(new_n2666_), .B(new_n2660_), .Y(new_n2671_));
  INVX1    g01669(.A(\A[523] ), .Y(new_n2672_));
  OR2X1    g01670(.A(\A[524] ), .B(new_n2672_), .Y(new_n2673_));
  INVX1    g01671(.A(\A[525] ), .Y(new_n2674_));
  AOI21X1  g01672(.A0(\A[524] ), .A1(new_n2672_), .B0(new_n2674_), .Y(new_n2675_));
  XOR2X1   g01673(.A(\A[524] ), .B(\A[523] ), .Y(new_n2676_));
  AND2X1   g01674(.A(new_n2676_), .B(new_n2674_), .Y(new_n2677_));
  AOI21X1  g01675(.A0(new_n2675_), .A1(new_n2673_), .B0(new_n2677_), .Y(new_n2678_));
  INVX1    g01676(.A(\A[528] ), .Y(new_n2679_));
  INVX1    g01677(.A(\A[526] ), .Y(new_n2680_));
  OR2X1    g01678(.A(\A[527] ), .B(new_n2680_), .Y(new_n2681_));
  AOI21X1  g01679(.A0(\A[527] ), .A1(new_n2680_), .B0(new_n2679_), .Y(new_n2682_));
  XOR2X1   g01680(.A(\A[527] ), .B(\A[526] ), .Y(new_n2683_));
  AOI22X1  g01681(.A0(new_n2683_), .A1(new_n2679_), .B0(new_n2682_), .B1(new_n2681_), .Y(new_n2684_));
  AND2X1   g01682(.A(\A[527] ), .B(\A[526] ), .Y(new_n2685_));
  AOI21X1  g01683(.A0(new_n2683_), .A1(\A[528] ), .B0(new_n2685_), .Y(new_n2686_));
  AND2X1   g01684(.A(\A[524] ), .B(\A[523] ), .Y(new_n2687_));
  AOI21X1  g01685(.A0(new_n2676_), .A1(\A[525] ), .B0(new_n2687_), .Y(new_n2688_));
  XOR2X1   g01686(.A(new_n2684_), .B(new_n2678_), .Y(new_n2689_));
  XOR2X1   g01687(.A(new_n2689_), .B(new_n2671_), .Y(new_n2690_));
  INVX1    g01688(.A(new_n2690_), .Y(new_n2691_));
  INVX1    g01689(.A(\A[517] ), .Y(new_n2692_));
  OR2X1    g01690(.A(\A[518] ), .B(new_n2692_), .Y(new_n2693_));
  INVX1    g01691(.A(\A[519] ), .Y(new_n2694_));
  AOI21X1  g01692(.A0(\A[518] ), .A1(new_n2692_), .B0(new_n2694_), .Y(new_n2695_));
  AND2X1   g01693(.A(new_n2695_), .B(new_n2693_), .Y(new_n2696_));
  XOR2X1   g01694(.A(\A[518] ), .B(\A[517] ), .Y(new_n2697_));
  AND2X1   g01695(.A(new_n2697_), .B(new_n2694_), .Y(new_n2698_));
  OR2X1    g01696(.A(new_n2698_), .B(new_n2696_), .Y(new_n2699_));
  INVX1    g01697(.A(\A[522] ), .Y(new_n2700_));
  INVX1    g01698(.A(\A[520] ), .Y(new_n2701_));
  OR2X1    g01699(.A(\A[521] ), .B(new_n2701_), .Y(new_n2702_));
  AOI21X1  g01700(.A0(\A[521] ), .A1(new_n2701_), .B0(new_n2700_), .Y(new_n2703_));
  XOR2X1   g01701(.A(\A[521] ), .B(\A[520] ), .Y(new_n2704_));
  AOI22X1  g01702(.A0(new_n2704_), .A1(new_n2700_), .B0(new_n2703_), .B1(new_n2702_), .Y(new_n2705_));
  AND2X1   g01703(.A(\A[521] ), .B(\A[520] ), .Y(new_n2706_));
  AOI21X1  g01704(.A0(new_n2704_), .A1(\A[522] ), .B0(new_n2706_), .Y(new_n2707_));
  AND2X1   g01705(.A(\A[518] ), .B(\A[517] ), .Y(new_n2708_));
  AOI21X1  g01706(.A0(new_n2697_), .A1(\A[519] ), .B0(new_n2708_), .Y(new_n2709_));
  XOR2X1   g01707(.A(new_n2705_), .B(new_n2699_), .Y(new_n2710_));
  INVX1    g01708(.A(\A[511] ), .Y(new_n2711_));
  OR2X1    g01709(.A(\A[512] ), .B(new_n2711_), .Y(new_n2712_));
  INVX1    g01710(.A(\A[513] ), .Y(new_n2713_));
  AOI21X1  g01711(.A0(\A[512] ), .A1(new_n2711_), .B0(new_n2713_), .Y(new_n2714_));
  XOR2X1   g01712(.A(\A[512] ), .B(\A[511] ), .Y(new_n2715_));
  AND2X1   g01713(.A(new_n2715_), .B(new_n2713_), .Y(new_n2716_));
  AOI21X1  g01714(.A0(new_n2714_), .A1(new_n2712_), .B0(new_n2716_), .Y(new_n2717_));
  INVX1    g01715(.A(\A[516] ), .Y(new_n2718_));
  INVX1    g01716(.A(\A[514] ), .Y(new_n2719_));
  OR2X1    g01717(.A(\A[515] ), .B(new_n2719_), .Y(new_n2720_));
  AOI21X1  g01718(.A0(\A[515] ), .A1(new_n2719_), .B0(new_n2718_), .Y(new_n2721_));
  XOR2X1   g01719(.A(\A[515] ), .B(\A[514] ), .Y(new_n2722_));
  AOI22X1  g01720(.A0(new_n2722_), .A1(new_n2718_), .B0(new_n2721_), .B1(new_n2720_), .Y(new_n2723_));
  AND2X1   g01721(.A(\A[515] ), .B(\A[514] ), .Y(new_n2724_));
  AOI21X1  g01722(.A0(new_n2722_), .A1(\A[516] ), .B0(new_n2724_), .Y(new_n2725_));
  AND2X1   g01723(.A(\A[512] ), .B(\A[511] ), .Y(new_n2726_));
  AOI21X1  g01724(.A0(new_n2715_), .A1(\A[513] ), .B0(new_n2726_), .Y(new_n2727_));
  XOR2X1   g01725(.A(new_n2723_), .B(new_n2717_), .Y(new_n2728_));
  XOR2X1   g01726(.A(new_n2728_), .B(new_n2710_), .Y(new_n2729_));
  XOR2X1   g01727(.A(new_n2729_), .B(new_n2691_), .Y(new_n2730_));
  XOR2X1   g01728(.A(new_n2730_), .B(new_n2653_), .Y(new_n2731_));
  XOR2X1   g01729(.A(new_n2731_), .B(new_n2577_), .Y(new_n2732_));
  INVX1    g01730(.A(\A[649] ), .Y(new_n2733_));
  OR2X1    g01731(.A(\A[650] ), .B(new_n2733_), .Y(new_n2734_));
  INVX1    g01732(.A(\A[651] ), .Y(new_n2735_));
  AOI21X1  g01733(.A0(\A[650] ), .A1(new_n2733_), .B0(new_n2735_), .Y(new_n2736_));
  XOR2X1   g01734(.A(\A[650] ), .B(\A[649] ), .Y(new_n2737_));
  AND2X1   g01735(.A(new_n2737_), .B(new_n2735_), .Y(new_n2738_));
  AOI21X1  g01736(.A0(new_n2736_), .A1(new_n2734_), .B0(new_n2738_), .Y(new_n2739_));
  INVX1    g01737(.A(\A[654] ), .Y(new_n2740_));
  INVX1    g01738(.A(\A[652] ), .Y(new_n2741_));
  OR2X1    g01739(.A(\A[653] ), .B(new_n2741_), .Y(new_n2742_));
  AOI21X1  g01740(.A0(\A[653] ), .A1(new_n2741_), .B0(new_n2740_), .Y(new_n2743_));
  XOR2X1   g01741(.A(\A[653] ), .B(\A[652] ), .Y(new_n2744_));
  AOI22X1  g01742(.A0(new_n2744_), .A1(new_n2740_), .B0(new_n2743_), .B1(new_n2742_), .Y(new_n2745_));
  AND2X1   g01743(.A(\A[653] ), .B(\A[652] ), .Y(new_n2746_));
  AOI21X1  g01744(.A0(new_n2744_), .A1(\A[654] ), .B0(new_n2746_), .Y(new_n2747_));
  AND2X1   g01745(.A(\A[650] ), .B(\A[649] ), .Y(new_n2748_));
  AOI21X1  g01746(.A0(new_n2737_), .A1(\A[651] ), .B0(new_n2748_), .Y(new_n2749_));
  XOR2X1   g01747(.A(new_n2745_), .B(new_n2739_), .Y(new_n2750_));
  INVX1    g01748(.A(\A[643] ), .Y(new_n2751_));
  OR2X1    g01749(.A(\A[644] ), .B(new_n2751_), .Y(new_n2752_));
  INVX1    g01750(.A(\A[645] ), .Y(new_n2753_));
  AOI21X1  g01751(.A0(\A[644] ), .A1(new_n2751_), .B0(new_n2753_), .Y(new_n2754_));
  XOR2X1   g01752(.A(\A[644] ), .B(\A[643] ), .Y(new_n2755_));
  AND2X1   g01753(.A(new_n2755_), .B(new_n2753_), .Y(new_n2756_));
  AOI21X1  g01754(.A0(new_n2754_), .A1(new_n2752_), .B0(new_n2756_), .Y(new_n2757_));
  INVX1    g01755(.A(\A[648] ), .Y(new_n2758_));
  INVX1    g01756(.A(\A[646] ), .Y(new_n2759_));
  OR2X1    g01757(.A(\A[647] ), .B(new_n2759_), .Y(new_n2760_));
  AOI21X1  g01758(.A0(\A[647] ), .A1(new_n2759_), .B0(new_n2758_), .Y(new_n2761_));
  XOR2X1   g01759(.A(\A[647] ), .B(\A[646] ), .Y(new_n2762_));
  AOI22X1  g01760(.A0(new_n2762_), .A1(new_n2758_), .B0(new_n2761_), .B1(new_n2760_), .Y(new_n2763_));
  AND2X1   g01761(.A(\A[647] ), .B(\A[646] ), .Y(new_n2764_));
  AOI21X1  g01762(.A0(new_n2762_), .A1(\A[648] ), .B0(new_n2764_), .Y(new_n2765_));
  AND2X1   g01763(.A(\A[644] ), .B(\A[643] ), .Y(new_n2766_));
  AOI21X1  g01764(.A0(new_n2755_), .A1(\A[645] ), .B0(new_n2766_), .Y(new_n2767_));
  XOR2X1   g01765(.A(new_n2763_), .B(new_n2757_), .Y(new_n2768_));
  XOR2X1   g01766(.A(new_n2768_), .B(new_n2750_), .Y(new_n2769_));
  INVX1    g01767(.A(\A[637] ), .Y(new_n2770_));
  OR2X1    g01768(.A(\A[638] ), .B(new_n2770_), .Y(new_n2771_));
  INVX1    g01769(.A(\A[639] ), .Y(new_n2772_));
  AOI21X1  g01770(.A0(\A[638] ), .A1(new_n2770_), .B0(new_n2772_), .Y(new_n2773_));
  AND2X1   g01771(.A(new_n2773_), .B(new_n2771_), .Y(new_n2774_));
  XOR2X1   g01772(.A(\A[638] ), .B(\A[637] ), .Y(new_n2775_));
  AND2X1   g01773(.A(new_n2775_), .B(new_n2772_), .Y(new_n2776_));
  OR2X1    g01774(.A(new_n2776_), .B(new_n2774_), .Y(new_n2777_));
  INVX1    g01775(.A(\A[642] ), .Y(new_n2778_));
  INVX1    g01776(.A(\A[640] ), .Y(new_n2779_));
  OR2X1    g01777(.A(\A[641] ), .B(new_n2779_), .Y(new_n2780_));
  AOI21X1  g01778(.A0(\A[641] ), .A1(new_n2779_), .B0(new_n2778_), .Y(new_n2781_));
  XOR2X1   g01779(.A(\A[641] ), .B(\A[640] ), .Y(new_n2782_));
  AOI22X1  g01780(.A0(new_n2782_), .A1(new_n2778_), .B0(new_n2781_), .B1(new_n2780_), .Y(new_n2783_));
  AND2X1   g01781(.A(\A[641] ), .B(\A[640] ), .Y(new_n2784_));
  AOI21X1  g01782(.A0(new_n2782_), .A1(\A[642] ), .B0(new_n2784_), .Y(new_n2785_));
  AND2X1   g01783(.A(\A[638] ), .B(\A[637] ), .Y(new_n2786_));
  AOI21X1  g01784(.A0(new_n2775_), .A1(\A[639] ), .B0(new_n2786_), .Y(new_n2787_));
  XOR2X1   g01785(.A(new_n2783_), .B(new_n2777_), .Y(new_n2788_));
  INVX1    g01786(.A(\A[631] ), .Y(new_n2789_));
  OR2X1    g01787(.A(\A[632] ), .B(new_n2789_), .Y(new_n2790_));
  INVX1    g01788(.A(\A[633] ), .Y(new_n2791_));
  AOI21X1  g01789(.A0(\A[632] ), .A1(new_n2789_), .B0(new_n2791_), .Y(new_n2792_));
  XOR2X1   g01790(.A(\A[632] ), .B(\A[631] ), .Y(new_n2793_));
  AND2X1   g01791(.A(new_n2793_), .B(new_n2791_), .Y(new_n2794_));
  AOI21X1  g01792(.A0(new_n2792_), .A1(new_n2790_), .B0(new_n2794_), .Y(new_n2795_));
  INVX1    g01793(.A(\A[636] ), .Y(new_n2796_));
  INVX1    g01794(.A(\A[634] ), .Y(new_n2797_));
  OR2X1    g01795(.A(\A[635] ), .B(new_n2797_), .Y(new_n2798_));
  AOI21X1  g01796(.A0(\A[635] ), .A1(new_n2797_), .B0(new_n2796_), .Y(new_n2799_));
  XOR2X1   g01797(.A(\A[635] ), .B(\A[634] ), .Y(new_n2800_));
  AOI22X1  g01798(.A0(new_n2800_), .A1(new_n2796_), .B0(new_n2799_), .B1(new_n2798_), .Y(new_n2801_));
  AND2X1   g01799(.A(\A[635] ), .B(\A[634] ), .Y(new_n2802_));
  AOI21X1  g01800(.A0(new_n2800_), .A1(\A[636] ), .B0(new_n2802_), .Y(new_n2803_));
  AND2X1   g01801(.A(\A[632] ), .B(\A[631] ), .Y(new_n2804_));
  AOI21X1  g01802(.A0(new_n2793_), .A1(\A[633] ), .B0(new_n2804_), .Y(new_n2805_));
  XOR2X1   g01803(.A(new_n2801_), .B(new_n2795_), .Y(new_n2806_));
  XOR2X1   g01804(.A(new_n2806_), .B(new_n2788_), .Y(new_n2807_));
  XOR2X1   g01805(.A(new_n2807_), .B(new_n2769_), .Y(new_n2808_));
  INVX1    g01806(.A(\A[625] ), .Y(new_n2809_));
  OR2X1    g01807(.A(\A[626] ), .B(new_n2809_), .Y(new_n2810_));
  INVX1    g01808(.A(\A[627] ), .Y(new_n2811_));
  AOI21X1  g01809(.A0(\A[626] ), .A1(new_n2809_), .B0(new_n2811_), .Y(new_n2812_));
  XOR2X1   g01810(.A(\A[626] ), .B(\A[625] ), .Y(new_n2813_));
  AND2X1   g01811(.A(new_n2813_), .B(new_n2811_), .Y(new_n2814_));
  AOI21X1  g01812(.A0(new_n2812_), .A1(new_n2810_), .B0(new_n2814_), .Y(new_n2815_));
  INVX1    g01813(.A(\A[630] ), .Y(new_n2816_));
  INVX1    g01814(.A(\A[628] ), .Y(new_n2817_));
  OR2X1    g01815(.A(\A[629] ), .B(new_n2817_), .Y(new_n2818_));
  AOI21X1  g01816(.A0(\A[629] ), .A1(new_n2817_), .B0(new_n2816_), .Y(new_n2819_));
  XOR2X1   g01817(.A(\A[629] ), .B(\A[628] ), .Y(new_n2820_));
  AOI22X1  g01818(.A0(new_n2820_), .A1(new_n2816_), .B0(new_n2819_), .B1(new_n2818_), .Y(new_n2821_));
  AND2X1   g01819(.A(\A[629] ), .B(\A[628] ), .Y(new_n2822_));
  AOI21X1  g01820(.A0(new_n2820_), .A1(\A[630] ), .B0(new_n2822_), .Y(new_n2823_));
  AND2X1   g01821(.A(\A[626] ), .B(\A[625] ), .Y(new_n2824_));
  AOI21X1  g01822(.A0(new_n2813_), .A1(\A[627] ), .B0(new_n2824_), .Y(new_n2825_));
  XOR2X1   g01823(.A(new_n2821_), .B(new_n2815_), .Y(new_n2826_));
  INVX1    g01824(.A(\A[619] ), .Y(new_n2827_));
  OR2X1    g01825(.A(\A[620] ), .B(new_n2827_), .Y(new_n2828_));
  INVX1    g01826(.A(\A[621] ), .Y(new_n2829_));
  AOI21X1  g01827(.A0(\A[620] ), .A1(new_n2827_), .B0(new_n2829_), .Y(new_n2830_));
  XOR2X1   g01828(.A(\A[620] ), .B(\A[619] ), .Y(new_n2831_));
  AND2X1   g01829(.A(new_n2831_), .B(new_n2829_), .Y(new_n2832_));
  AOI21X1  g01830(.A0(new_n2830_), .A1(new_n2828_), .B0(new_n2832_), .Y(new_n2833_));
  INVX1    g01831(.A(\A[624] ), .Y(new_n2834_));
  INVX1    g01832(.A(\A[622] ), .Y(new_n2835_));
  OR2X1    g01833(.A(\A[623] ), .B(new_n2835_), .Y(new_n2836_));
  AOI21X1  g01834(.A0(\A[623] ), .A1(new_n2835_), .B0(new_n2834_), .Y(new_n2837_));
  XOR2X1   g01835(.A(\A[623] ), .B(\A[622] ), .Y(new_n2838_));
  AOI22X1  g01836(.A0(new_n2838_), .A1(new_n2834_), .B0(new_n2837_), .B1(new_n2836_), .Y(new_n2839_));
  AND2X1   g01837(.A(\A[623] ), .B(\A[622] ), .Y(new_n2840_));
  AOI21X1  g01838(.A0(new_n2838_), .A1(\A[624] ), .B0(new_n2840_), .Y(new_n2841_));
  AND2X1   g01839(.A(\A[620] ), .B(\A[619] ), .Y(new_n2842_));
  AOI21X1  g01840(.A0(new_n2831_), .A1(\A[621] ), .B0(new_n2842_), .Y(new_n2843_));
  XOR2X1   g01841(.A(new_n2839_), .B(new_n2833_), .Y(new_n2844_));
  XOR2X1   g01842(.A(new_n2844_), .B(new_n2826_), .Y(new_n2845_));
  INVX1    g01843(.A(\A[613] ), .Y(new_n2846_));
  OR2X1    g01844(.A(\A[614] ), .B(new_n2846_), .Y(new_n2847_));
  INVX1    g01845(.A(\A[615] ), .Y(new_n2848_));
  AOI21X1  g01846(.A0(\A[614] ), .A1(new_n2846_), .B0(new_n2848_), .Y(new_n2849_));
  AND2X1   g01847(.A(new_n2849_), .B(new_n2847_), .Y(new_n2850_));
  XOR2X1   g01848(.A(\A[614] ), .B(\A[613] ), .Y(new_n2851_));
  AND2X1   g01849(.A(new_n2851_), .B(new_n2848_), .Y(new_n2852_));
  OR2X1    g01850(.A(new_n2852_), .B(new_n2850_), .Y(new_n2853_));
  INVX1    g01851(.A(\A[618] ), .Y(new_n2854_));
  INVX1    g01852(.A(\A[616] ), .Y(new_n2855_));
  OR2X1    g01853(.A(\A[617] ), .B(new_n2855_), .Y(new_n2856_));
  AOI21X1  g01854(.A0(\A[617] ), .A1(new_n2855_), .B0(new_n2854_), .Y(new_n2857_));
  XOR2X1   g01855(.A(\A[617] ), .B(\A[616] ), .Y(new_n2858_));
  AOI22X1  g01856(.A0(new_n2858_), .A1(new_n2854_), .B0(new_n2857_), .B1(new_n2856_), .Y(new_n2859_));
  AND2X1   g01857(.A(\A[617] ), .B(\A[616] ), .Y(new_n2860_));
  AOI21X1  g01858(.A0(new_n2858_), .A1(\A[618] ), .B0(new_n2860_), .Y(new_n2861_));
  AND2X1   g01859(.A(\A[614] ), .B(\A[613] ), .Y(new_n2862_));
  AOI21X1  g01860(.A0(new_n2851_), .A1(\A[615] ), .B0(new_n2862_), .Y(new_n2863_));
  XOR2X1   g01861(.A(new_n2859_), .B(new_n2853_), .Y(new_n2864_));
  INVX1    g01862(.A(\A[607] ), .Y(new_n2865_));
  OR2X1    g01863(.A(\A[608] ), .B(new_n2865_), .Y(new_n2866_));
  INVX1    g01864(.A(\A[609] ), .Y(new_n2867_));
  AOI21X1  g01865(.A0(\A[608] ), .A1(new_n2865_), .B0(new_n2867_), .Y(new_n2868_));
  XOR2X1   g01866(.A(\A[608] ), .B(\A[607] ), .Y(new_n2869_));
  AND2X1   g01867(.A(new_n2869_), .B(new_n2867_), .Y(new_n2870_));
  AOI21X1  g01868(.A0(new_n2868_), .A1(new_n2866_), .B0(new_n2870_), .Y(new_n2871_));
  INVX1    g01869(.A(\A[612] ), .Y(new_n2872_));
  INVX1    g01870(.A(\A[610] ), .Y(new_n2873_));
  OR2X1    g01871(.A(\A[611] ), .B(new_n2873_), .Y(new_n2874_));
  AOI21X1  g01872(.A0(\A[611] ), .A1(new_n2873_), .B0(new_n2872_), .Y(new_n2875_));
  XOR2X1   g01873(.A(\A[611] ), .B(\A[610] ), .Y(new_n2876_));
  AOI22X1  g01874(.A0(new_n2876_), .A1(new_n2872_), .B0(new_n2875_), .B1(new_n2874_), .Y(new_n2877_));
  AND2X1   g01875(.A(\A[611] ), .B(\A[610] ), .Y(new_n2878_));
  AOI21X1  g01876(.A0(new_n2876_), .A1(\A[612] ), .B0(new_n2878_), .Y(new_n2879_));
  AND2X1   g01877(.A(\A[608] ), .B(\A[607] ), .Y(new_n2880_));
  AOI21X1  g01878(.A0(new_n2869_), .A1(\A[609] ), .B0(new_n2880_), .Y(new_n2881_));
  XOR2X1   g01879(.A(new_n2877_), .B(new_n2871_), .Y(new_n2882_));
  XOR2X1   g01880(.A(new_n2882_), .B(new_n2864_), .Y(new_n2883_));
  XOR2X1   g01881(.A(new_n2883_), .B(new_n2845_), .Y(new_n2884_));
  XOR2X1   g01882(.A(new_n2884_), .B(new_n2808_), .Y(new_n2885_));
  INVX1    g01883(.A(\A[601] ), .Y(new_n2886_));
  OR2X1    g01884(.A(\A[602] ), .B(new_n2886_), .Y(new_n2887_));
  INVX1    g01885(.A(\A[603] ), .Y(new_n2888_));
  AOI21X1  g01886(.A0(\A[602] ), .A1(new_n2886_), .B0(new_n2888_), .Y(new_n2889_));
  XOR2X1   g01887(.A(\A[602] ), .B(\A[601] ), .Y(new_n2890_));
  AND2X1   g01888(.A(new_n2890_), .B(new_n2888_), .Y(new_n2891_));
  AOI21X1  g01889(.A0(new_n2889_), .A1(new_n2887_), .B0(new_n2891_), .Y(new_n2892_));
  INVX1    g01890(.A(\A[606] ), .Y(new_n2893_));
  INVX1    g01891(.A(\A[604] ), .Y(new_n2894_));
  OR2X1    g01892(.A(\A[605] ), .B(new_n2894_), .Y(new_n2895_));
  AOI21X1  g01893(.A0(\A[605] ), .A1(new_n2894_), .B0(new_n2893_), .Y(new_n2896_));
  XOR2X1   g01894(.A(\A[605] ), .B(\A[604] ), .Y(new_n2897_));
  AOI22X1  g01895(.A0(new_n2897_), .A1(new_n2893_), .B0(new_n2896_), .B1(new_n2895_), .Y(new_n2898_));
  AND2X1   g01896(.A(\A[605] ), .B(\A[604] ), .Y(new_n2899_));
  AOI21X1  g01897(.A0(new_n2897_), .A1(\A[606] ), .B0(new_n2899_), .Y(new_n2900_));
  AND2X1   g01898(.A(\A[602] ), .B(\A[601] ), .Y(new_n2901_));
  AOI21X1  g01899(.A0(new_n2890_), .A1(\A[603] ), .B0(new_n2901_), .Y(new_n2902_));
  XOR2X1   g01900(.A(new_n2898_), .B(new_n2892_), .Y(new_n2903_));
  INVX1    g01901(.A(\A[595] ), .Y(new_n2904_));
  OR2X1    g01902(.A(\A[596] ), .B(new_n2904_), .Y(new_n2905_));
  INVX1    g01903(.A(\A[597] ), .Y(new_n2906_));
  AOI21X1  g01904(.A0(\A[596] ), .A1(new_n2904_), .B0(new_n2906_), .Y(new_n2907_));
  XOR2X1   g01905(.A(\A[596] ), .B(\A[595] ), .Y(new_n2908_));
  AND2X1   g01906(.A(new_n2908_), .B(new_n2906_), .Y(new_n2909_));
  AOI21X1  g01907(.A0(new_n2907_), .A1(new_n2905_), .B0(new_n2909_), .Y(new_n2910_));
  INVX1    g01908(.A(\A[600] ), .Y(new_n2911_));
  INVX1    g01909(.A(\A[598] ), .Y(new_n2912_));
  OR2X1    g01910(.A(\A[599] ), .B(new_n2912_), .Y(new_n2913_));
  AOI21X1  g01911(.A0(\A[599] ), .A1(new_n2912_), .B0(new_n2911_), .Y(new_n2914_));
  XOR2X1   g01912(.A(\A[599] ), .B(\A[598] ), .Y(new_n2915_));
  AOI22X1  g01913(.A0(new_n2915_), .A1(new_n2911_), .B0(new_n2914_), .B1(new_n2913_), .Y(new_n2916_));
  AND2X1   g01914(.A(\A[599] ), .B(\A[598] ), .Y(new_n2917_));
  AOI21X1  g01915(.A0(new_n2915_), .A1(\A[600] ), .B0(new_n2917_), .Y(new_n2918_));
  AND2X1   g01916(.A(\A[596] ), .B(\A[595] ), .Y(new_n2919_));
  AOI21X1  g01917(.A0(new_n2908_), .A1(\A[597] ), .B0(new_n2919_), .Y(new_n2920_));
  XOR2X1   g01918(.A(new_n2916_), .B(new_n2910_), .Y(new_n2921_));
  XOR2X1   g01919(.A(new_n2921_), .B(new_n2903_), .Y(new_n2922_));
  INVX1    g01920(.A(\A[589] ), .Y(new_n2923_));
  OR2X1    g01921(.A(\A[590] ), .B(new_n2923_), .Y(new_n2924_));
  INVX1    g01922(.A(\A[591] ), .Y(new_n2925_));
  AOI21X1  g01923(.A0(\A[590] ), .A1(new_n2923_), .B0(new_n2925_), .Y(new_n2926_));
  AND2X1   g01924(.A(new_n2926_), .B(new_n2924_), .Y(new_n2927_));
  XOR2X1   g01925(.A(\A[590] ), .B(\A[589] ), .Y(new_n2928_));
  AND2X1   g01926(.A(new_n2928_), .B(new_n2925_), .Y(new_n2929_));
  OR2X1    g01927(.A(new_n2929_), .B(new_n2927_), .Y(new_n2930_));
  INVX1    g01928(.A(\A[594] ), .Y(new_n2931_));
  INVX1    g01929(.A(\A[592] ), .Y(new_n2932_));
  OR2X1    g01930(.A(\A[593] ), .B(new_n2932_), .Y(new_n2933_));
  AOI21X1  g01931(.A0(\A[593] ), .A1(new_n2932_), .B0(new_n2931_), .Y(new_n2934_));
  XOR2X1   g01932(.A(\A[593] ), .B(\A[592] ), .Y(new_n2935_));
  AOI22X1  g01933(.A0(new_n2935_), .A1(new_n2931_), .B0(new_n2934_), .B1(new_n2933_), .Y(new_n2936_));
  AND2X1   g01934(.A(\A[593] ), .B(\A[592] ), .Y(new_n2937_));
  AOI21X1  g01935(.A0(new_n2935_), .A1(\A[594] ), .B0(new_n2937_), .Y(new_n2938_));
  AND2X1   g01936(.A(\A[590] ), .B(\A[589] ), .Y(new_n2939_));
  AOI21X1  g01937(.A0(new_n2928_), .A1(\A[591] ), .B0(new_n2939_), .Y(new_n2940_));
  XOR2X1   g01938(.A(new_n2936_), .B(new_n2930_), .Y(new_n2941_));
  INVX1    g01939(.A(\A[583] ), .Y(new_n2942_));
  OR2X1    g01940(.A(\A[584] ), .B(new_n2942_), .Y(new_n2943_));
  INVX1    g01941(.A(\A[585] ), .Y(new_n2944_));
  AOI21X1  g01942(.A0(\A[584] ), .A1(new_n2942_), .B0(new_n2944_), .Y(new_n2945_));
  XOR2X1   g01943(.A(\A[584] ), .B(\A[583] ), .Y(new_n2946_));
  AND2X1   g01944(.A(new_n2946_), .B(new_n2944_), .Y(new_n2947_));
  AOI21X1  g01945(.A0(new_n2945_), .A1(new_n2943_), .B0(new_n2947_), .Y(new_n2948_));
  INVX1    g01946(.A(\A[588] ), .Y(new_n2949_));
  INVX1    g01947(.A(\A[586] ), .Y(new_n2950_));
  OR2X1    g01948(.A(\A[587] ), .B(new_n2950_), .Y(new_n2951_));
  AOI21X1  g01949(.A0(\A[587] ), .A1(new_n2950_), .B0(new_n2949_), .Y(new_n2952_));
  XOR2X1   g01950(.A(\A[587] ), .B(\A[586] ), .Y(new_n2953_));
  AOI22X1  g01951(.A0(new_n2953_), .A1(new_n2949_), .B0(new_n2952_), .B1(new_n2951_), .Y(new_n2954_));
  AND2X1   g01952(.A(\A[587] ), .B(\A[586] ), .Y(new_n2955_));
  AOI21X1  g01953(.A0(new_n2953_), .A1(\A[588] ), .B0(new_n2955_), .Y(new_n2956_));
  AND2X1   g01954(.A(\A[584] ), .B(\A[583] ), .Y(new_n2957_));
  AOI21X1  g01955(.A0(new_n2946_), .A1(\A[585] ), .B0(new_n2957_), .Y(new_n2958_));
  XOR2X1   g01956(.A(new_n2954_), .B(new_n2948_), .Y(new_n2959_));
  XOR2X1   g01957(.A(new_n2959_), .B(new_n2941_), .Y(new_n2960_));
  XOR2X1   g01958(.A(new_n2960_), .B(new_n2922_), .Y(new_n2961_));
  INVX1    g01959(.A(\A[577] ), .Y(new_n2962_));
  OR2X1    g01960(.A(\A[578] ), .B(new_n2962_), .Y(new_n2963_));
  INVX1    g01961(.A(\A[579] ), .Y(new_n2964_));
  AOI21X1  g01962(.A0(\A[578] ), .A1(new_n2962_), .B0(new_n2964_), .Y(new_n2965_));
  XOR2X1   g01963(.A(\A[578] ), .B(\A[577] ), .Y(new_n2966_));
  AND2X1   g01964(.A(new_n2966_), .B(new_n2964_), .Y(new_n2967_));
  AOI21X1  g01965(.A0(new_n2965_), .A1(new_n2963_), .B0(new_n2967_), .Y(new_n2968_));
  INVX1    g01966(.A(\A[582] ), .Y(new_n2969_));
  INVX1    g01967(.A(\A[580] ), .Y(new_n2970_));
  OR2X1    g01968(.A(\A[581] ), .B(new_n2970_), .Y(new_n2971_));
  AOI21X1  g01969(.A0(\A[581] ), .A1(new_n2970_), .B0(new_n2969_), .Y(new_n2972_));
  XOR2X1   g01970(.A(\A[581] ), .B(\A[580] ), .Y(new_n2973_));
  AOI22X1  g01971(.A0(new_n2973_), .A1(new_n2969_), .B0(new_n2972_), .B1(new_n2971_), .Y(new_n2974_));
  AND2X1   g01972(.A(\A[581] ), .B(\A[580] ), .Y(new_n2975_));
  AOI21X1  g01973(.A0(new_n2973_), .A1(\A[582] ), .B0(new_n2975_), .Y(new_n2976_));
  AND2X1   g01974(.A(\A[578] ), .B(\A[577] ), .Y(new_n2977_));
  AOI21X1  g01975(.A0(new_n2966_), .A1(\A[579] ), .B0(new_n2977_), .Y(new_n2978_));
  XOR2X1   g01976(.A(new_n2974_), .B(new_n2968_), .Y(new_n2979_));
  INVX1    g01977(.A(\A[571] ), .Y(new_n2980_));
  OR2X1    g01978(.A(\A[572] ), .B(new_n2980_), .Y(new_n2981_));
  INVX1    g01979(.A(\A[573] ), .Y(new_n2982_));
  AOI21X1  g01980(.A0(\A[572] ), .A1(new_n2980_), .B0(new_n2982_), .Y(new_n2983_));
  XOR2X1   g01981(.A(\A[572] ), .B(\A[571] ), .Y(new_n2984_));
  AND2X1   g01982(.A(new_n2984_), .B(new_n2982_), .Y(new_n2985_));
  AOI21X1  g01983(.A0(new_n2983_), .A1(new_n2981_), .B0(new_n2985_), .Y(new_n2986_));
  INVX1    g01984(.A(\A[576] ), .Y(new_n2987_));
  INVX1    g01985(.A(\A[574] ), .Y(new_n2988_));
  OR2X1    g01986(.A(\A[575] ), .B(new_n2988_), .Y(new_n2989_));
  AOI21X1  g01987(.A0(\A[575] ), .A1(new_n2988_), .B0(new_n2987_), .Y(new_n2990_));
  XOR2X1   g01988(.A(\A[575] ), .B(\A[574] ), .Y(new_n2991_));
  AOI22X1  g01989(.A0(new_n2991_), .A1(new_n2987_), .B0(new_n2990_), .B1(new_n2989_), .Y(new_n2992_));
  AND2X1   g01990(.A(\A[575] ), .B(\A[574] ), .Y(new_n2993_));
  AOI21X1  g01991(.A0(new_n2991_), .A1(\A[576] ), .B0(new_n2993_), .Y(new_n2994_));
  AND2X1   g01992(.A(\A[572] ), .B(\A[571] ), .Y(new_n2995_));
  AOI21X1  g01993(.A0(new_n2984_), .A1(\A[573] ), .B0(new_n2995_), .Y(new_n2996_));
  XOR2X1   g01994(.A(new_n2992_), .B(new_n2986_), .Y(new_n2997_));
  XOR2X1   g01995(.A(new_n2997_), .B(new_n2979_), .Y(new_n2998_));
  INVX1    g01996(.A(new_n2998_), .Y(new_n2999_));
  INVX1    g01997(.A(\A[565] ), .Y(new_n3000_));
  OR2X1    g01998(.A(\A[566] ), .B(new_n3000_), .Y(new_n3001_));
  INVX1    g01999(.A(\A[567] ), .Y(new_n3002_));
  AOI21X1  g02000(.A0(\A[566] ), .A1(new_n3000_), .B0(new_n3002_), .Y(new_n3003_));
  AND2X1   g02001(.A(new_n3003_), .B(new_n3001_), .Y(new_n3004_));
  XOR2X1   g02002(.A(\A[566] ), .B(\A[565] ), .Y(new_n3005_));
  AND2X1   g02003(.A(new_n3005_), .B(new_n3002_), .Y(new_n3006_));
  OR2X1    g02004(.A(new_n3006_), .B(new_n3004_), .Y(new_n3007_));
  INVX1    g02005(.A(\A[570] ), .Y(new_n3008_));
  INVX1    g02006(.A(\A[568] ), .Y(new_n3009_));
  OR2X1    g02007(.A(\A[569] ), .B(new_n3009_), .Y(new_n3010_));
  AOI21X1  g02008(.A0(\A[569] ), .A1(new_n3009_), .B0(new_n3008_), .Y(new_n3011_));
  XOR2X1   g02009(.A(\A[569] ), .B(\A[568] ), .Y(new_n3012_));
  AOI22X1  g02010(.A0(new_n3012_), .A1(new_n3008_), .B0(new_n3011_), .B1(new_n3010_), .Y(new_n3013_));
  AND2X1   g02011(.A(\A[569] ), .B(\A[568] ), .Y(new_n3014_));
  AOI21X1  g02012(.A0(new_n3012_), .A1(\A[570] ), .B0(new_n3014_), .Y(new_n3015_));
  AND2X1   g02013(.A(\A[566] ), .B(\A[565] ), .Y(new_n3016_));
  AOI21X1  g02014(.A0(new_n3005_), .A1(\A[567] ), .B0(new_n3016_), .Y(new_n3017_));
  XOR2X1   g02015(.A(new_n3013_), .B(new_n3007_), .Y(new_n3018_));
  INVX1    g02016(.A(\A[559] ), .Y(new_n3019_));
  OR2X1    g02017(.A(\A[560] ), .B(new_n3019_), .Y(new_n3020_));
  INVX1    g02018(.A(\A[561] ), .Y(new_n3021_));
  AOI21X1  g02019(.A0(\A[560] ), .A1(new_n3019_), .B0(new_n3021_), .Y(new_n3022_));
  XOR2X1   g02020(.A(\A[560] ), .B(\A[559] ), .Y(new_n3023_));
  AND2X1   g02021(.A(new_n3023_), .B(new_n3021_), .Y(new_n3024_));
  AOI21X1  g02022(.A0(new_n3022_), .A1(new_n3020_), .B0(new_n3024_), .Y(new_n3025_));
  INVX1    g02023(.A(\A[564] ), .Y(new_n3026_));
  INVX1    g02024(.A(\A[562] ), .Y(new_n3027_));
  OR2X1    g02025(.A(\A[563] ), .B(new_n3027_), .Y(new_n3028_));
  AOI21X1  g02026(.A0(\A[563] ), .A1(new_n3027_), .B0(new_n3026_), .Y(new_n3029_));
  XOR2X1   g02027(.A(\A[563] ), .B(\A[562] ), .Y(new_n3030_));
  AOI22X1  g02028(.A0(new_n3030_), .A1(new_n3026_), .B0(new_n3029_), .B1(new_n3028_), .Y(new_n3031_));
  AND2X1   g02029(.A(\A[563] ), .B(\A[562] ), .Y(new_n3032_));
  AOI21X1  g02030(.A0(new_n3030_), .A1(\A[564] ), .B0(new_n3032_), .Y(new_n3033_));
  AND2X1   g02031(.A(\A[560] ), .B(\A[559] ), .Y(new_n3034_));
  AOI21X1  g02032(.A0(new_n3023_), .A1(\A[561] ), .B0(new_n3034_), .Y(new_n3035_));
  XOR2X1   g02033(.A(new_n3031_), .B(new_n3025_), .Y(new_n3036_));
  XOR2X1   g02034(.A(new_n3036_), .B(new_n3018_), .Y(new_n3037_));
  XOR2X1   g02035(.A(new_n3037_), .B(new_n2999_), .Y(new_n3038_));
  XOR2X1   g02036(.A(new_n3038_), .B(new_n2961_), .Y(new_n3039_));
  XOR2X1   g02037(.A(new_n3039_), .B(new_n2885_), .Y(new_n3040_));
  XOR2X1   g02038(.A(new_n3040_), .B(new_n2732_), .Y(new_n3041_));
  XOR2X1   g02039(.A(new_n2400_), .B(new_n2398_), .Y(new_n3042_));
  INVX1    g02040(.A(new_n3042_), .Y(new_n3043_));
  OR4X1    g02041(.A(new_n3043_), .B(new_n3041_), .C(new_n2423_), .D(new_n2411_), .Y(new_n3044_));
  OAI22X1  g02042(.A0(new_n3043_), .A1(new_n3041_), .B0(new_n2423_), .B1(new_n2411_), .Y(new_n3045_));
  NAND2X1  g02043(.A(new_n3045_), .B(new_n3044_), .Y(new_n3046_));
  AND2X1   g02044(.A(new_n2945_), .B(new_n2943_), .Y(new_n3047_));
  OR2X1    g02045(.A(new_n2947_), .B(new_n3047_), .Y(new_n3048_));
  XOR2X1   g02046(.A(new_n2954_), .B(new_n3048_), .Y(new_n3049_));
  XOR2X1   g02047(.A(new_n2958_), .B(new_n2956_), .Y(new_n3050_));
  NOR2X1   g02048(.A(new_n2954_), .B(new_n2948_), .Y(new_n3051_));
  NOR2X1   g02049(.A(new_n2958_), .B(new_n2956_), .Y(new_n3052_));
  AOI21X1  g02050(.A0(new_n3051_), .A1(new_n3050_), .B0(new_n3052_), .Y(new_n3053_));
  XOR2X1   g02051(.A(new_n3051_), .B(new_n3050_), .Y(new_n3054_));
  OAI21X1  g02052(.A0(new_n3053_), .A1(new_n3049_), .B0(new_n3054_), .Y(new_n3055_));
  INVX1    g02053(.A(new_n3055_), .Y(new_n3056_));
  XOR2X1   g02054(.A(new_n2936_), .B(new_n2930_), .Y(new_n3057_));
  AOI21X1  g02055(.A0(new_n2926_), .A1(new_n2924_), .B0(new_n2929_), .Y(new_n3058_));
  NOR4X1   g02056(.A(new_n2940_), .B(new_n2938_), .C(new_n2936_), .D(new_n3058_), .Y(new_n3059_));
  NOR4X1   g02057(.A(new_n2958_), .B(new_n2956_), .C(new_n2954_), .D(new_n2948_), .Y(new_n3060_));
  OR4X1    g02058(.A(new_n3060_), .B(new_n3049_), .C(new_n3059_), .D(new_n3057_), .Y(new_n3061_));
  XOR2X1   g02059(.A(new_n2940_), .B(new_n2938_), .Y(new_n3062_));
  NOR2X1   g02060(.A(new_n2936_), .B(new_n3058_), .Y(new_n3063_));
  NOR2X1   g02061(.A(new_n2940_), .B(new_n2938_), .Y(new_n3064_));
  AOI21X1  g02062(.A0(new_n3063_), .A1(new_n3062_), .B0(new_n3064_), .Y(new_n3065_));
  XOR2X1   g02063(.A(new_n3063_), .B(new_n3062_), .Y(new_n3066_));
  OAI21X1  g02064(.A0(new_n3065_), .A1(new_n3057_), .B0(new_n3066_), .Y(new_n3067_));
  XOR2X1   g02065(.A(new_n3067_), .B(new_n3061_), .Y(new_n3068_));
  AND2X1   g02066(.A(new_n3068_), .B(new_n3055_), .Y(new_n3069_));
  AND2X1   g02067(.A(new_n3067_), .B(new_n3061_), .Y(new_n3070_));
  OR2X1    g02068(.A(new_n2936_), .B(new_n3058_), .Y(new_n3071_));
  XOR2X1   g02069(.A(new_n3071_), .B(new_n3062_), .Y(new_n3072_));
  OR4X1    g02070(.A(new_n3049_), .B(new_n3059_), .C(new_n3072_), .D(new_n3057_), .Y(new_n3073_));
  OR4X1    g02071(.A(new_n2958_), .B(new_n2956_), .C(new_n2954_), .D(new_n2948_), .Y(new_n3074_));
  OAI21X1  g02072(.A0(new_n3065_), .A1(new_n3057_), .B0(new_n3074_), .Y(new_n3075_));
  NOR2X1   g02073(.A(new_n3075_), .B(new_n3073_), .Y(new_n3076_));
  OR2X1    g02074(.A(new_n3076_), .B(new_n3070_), .Y(new_n3077_));
  AOI21X1  g02075(.A0(new_n3077_), .A1(new_n3056_), .B0(new_n3069_), .Y(new_n3078_));
  AND2X1   g02076(.A(new_n2907_), .B(new_n2905_), .Y(new_n3079_));
  OR2X1    g02077(.A(new_n2909_), .B(new_n3079_), .Y(new_n3080_));
  XOR2X1   g02078(.A(new_n2916_), .B(new_n3080_), .Y(new_n3081_));
  XOR2X1   g02079(.A(new_n2920_), .B(new_n2918_), .Y(new_n3082_));
  NOR2X1   g02080(.A(new_n2916_), .B(new_n2910_), .Y(new_n3083_));
  NOR2X1   g02081(.A(new_n2920_), .B(new_n2918_), .Y(new_n3084_));
  AOI21X1  g02082(.A0(new_n3083_), .A1(new_n3082_), .B0(new_n3084_), .Y(new_n3085_));
  XOR2X1   g02083(.A(new_n3083_), .B(new_n3082_), .Y(new_n3086_));
  OAI21X1  g02084(.A0(new_n3085_), .A1(new_n3081_), .B0(new_n3086_), .Y(new_n3087_));
  AND2X1   g02085(.A(new_n2889_), .B(new_n2887_), .Y(new_n3088_));
  OR2X1    g02086(.A(new_n2891_), .B(new_n3088_), .Y(new_n3089_));
  XOR2X1   g02087(.A(new_n2898_), .B(new_n3089_), .Y(new_n3090_));
  NOR4X1   g02088(.A(new_n2902_), .B(new_n2900_), .C(new_n2898_), .D(new_n2892_), .Y(new_n3091_));
  NOR4X1   g02089(.A(new_n2920_), .B(new_n2918_), .C(new_n2916_), .D(new_n2910_), .Y(new_n3092_));
  OR4X1    g02090(.A(new_n3092_), .B(new_n3081_), .C(new_n3091_), .D(new_n3090_), .Y(new_n3093_));
  XOR2X1   g02091(.A(new_n2902_), .B(new_n2900_), .Y(new_n3094_));
  NOR2X1   g02092(.A(new_n2898_), .B(new_n2892_), .Y(new_n3095_));
  NOR2X1   g02093(.A(new_n2902_), .B(new_n2900_), .Y(new_n3096_));
  AOI21X1  g02094(.A0(new_n3095_), .A1(new_n3094_), .B0(new_n3096_), .Y(new_n3097_));
  XOR2X1   g02095(.A(new_n3095_), .B(new_n3094_), .Y(new_n3098_));
  OAI21X1  g02096(.A0(new_n3097_), .A1(new_n3090_), .B0(new_n3098_), .Y(new_n3099_));
  XOR2X1   g02097(.A(new_n3099_), .B(new_n3093_), .Y(new_n3100_));
  AND2X1   g02098(.A(new_n3100_), .B(new_n3087_), .Y(new_n3101_));
  NAND2X1  g02099(.A(new_n3099_), .B(new_n3093_), .Y(new_n3102_));
  OR2X1    g02100(.A(new_n2898_), .B(new_n2892_), .Y(new_n3103_));
  XOR2X1   g02101(.A(new_n3103_), .B(new_n3094_), .Y(new_n3104_));
  OR4X1    g02102(.A(new_n3081_), .B(new_n3091_), .C(new_n3104_), .D(new_n3090_), .Y(new_n3105_));
  AND2X1   g02103(.A(new_n2915_), .B(\A[600] ), .Y(new_n3106_));
  OR2X1    g02104(.A(new_n3106_), .B(new_n2917_), .Y(new_n3107_));
  XOR2X1   g02105(.A(new_n2920_), .B(new_n3107_), .Y(new_n3108_));
  XOR2X1   g02106(.A(new_n3083_), .B(new_n3108_), .Y(new_n3109_));
  OAI22X1  g02107(.A0(new_n3109_), .A1(new_n3085_), .B0(new_n3097_), .B1(new_n3090_), .Y(new_n3110_));
  OR2X1    g02108(.A(new_n3110_), .B(new_n3105_), .Y(new_n3111_));
  AOI21X1  g02109(.A0(new_n3111_), .A1(new_n3102_), .B0(new_n3087_), .Y(new_n3112_));
  INVX1    g02110(.A(new_n2922_), .Y(new_n3113_));
  OR2X1    g02111(.A(new_n2960_), .B(new_n3113_), .Y(new_n3114_));
  NOR3X1   g02112(.A(new_n3114_), .B(new_n3112_), .C(new_n3101_), .Y(new_n3115_));
  NAND2X1  g02113(.A(new_n3100_), .B(new_n3087_), .Y(new_n3116_));
  XOR2X1   g02114(.A(new_n2916_), .B(new_n2910_), .Y(new_n3117_));
  OR2X1    g02115(.A(new_n2916_), .B(new_n2910_), .Y(new_n3118_));
  OR2X1    g02116(.A(new_n2920_), .B(new_n2918_), .Y(new_n3119_));
  OAI21X1  g02117(.A0(new_n3118_), .A1(new_n3108_), .B0(new_n3119_), .Y(new_n3120_));
  AOI21X1  g02118(.A0(new_n3120_), .A1(new_n3117_), .B0(new_n3109_), .Y(new_n3121_));
  AND2X1   g02119(.A(new_n3099_), .B(new_n3093_), .Y(new_n3122_));
  NOR2X1   g02120(.A(new_n3110_), .B(new_n3105_), .Y(new_n3123_));
  OAI21X1  g02121(.A0(new_n3123_), .A1(new_n3122_), .B0(new_n3121_), .Y(new_n3124_));
  NOR2X1   g02122(.A(new_n2960_), .B(new_n3113_), .Y(new_n3125_));
  AOI21X1  g02123(.A0(new_n3124_), .A1(new_n3116_), .B0(new_n3125_), .Y(new_n3126_));
  OAI21X1  g02124(.A0(new_n3126_), .A1(new_n3115_), .B0(new_n3078_), .Y(new_n3127_));
  MX2X1    g02125(.A(new_n3077_), .B(new_n3068_), .S0(new_n3055_), .Y(new_n3128_));
  NOR3X1   g02126(.A(new_n3125_), .B(new_n3112_), .C(new_n3101_), .Y(new_n3129_));
  AOI21X1  g02127(.A0(new_n3124_), .A1(new_n3116_), .B0(new_n3114_), .Y(new_n3130_));
  OAI21X1  g02128(.A0(new_n3130_), .A1(new_n3129_), .B0(new_n3128_), .Y(new_n3131_));
  XOR2X1   g02129(.A(new_n3037_), .B(new_n2998_), .Y(new_n3132_));
  NOR2X1   g02130(.A(new_n3132_), .B(new_n2961_), .Y(new_n3133_));
  NAND3X1  g02131(.A(new_n3133_), .B(new_n3131_), .C(new_n3127_), .Y(new_n3134_));
  NAND3X1  g02132(.A(new_n3125_), .B(new_n3124_), .C(new_n3116_), .Y(new_n3135_));
  OAI21X1  g02133(.A0(new_n3112_), .A1(new_n3101_), .B0(new_n3114_), .Y(new_n3136_));
  AOI21X1  g02134(.A0(new_n3136_), .A1(new_n3135_), .B0(new_n3128_), .Y(new_n3137_));
  NAND3X1  g02135(.A(new_n3114_), .B(new_n3124_), .C(new_n3116_), .Y(new_n3138_));
  OAI21X1  g02136(.A0(new_n3112_), .A1(new_n3101_), .B0(new_n3125_), .Y(new_n3139_));
  AOI21X1  g02137(.A0(new_n3139_), .A1(new_n3138_), .B0(new_n3078_), .Y(new_n3140_));
  INVX1    g02138(.A(new_n3133_), .Y(new_n3141_));
  OAI21X1  g02139(.A0(new_n3140_), .A1(new_n3137_), .B0(new_n3141_), .Y(new_n3142_));
  AND2X1   g02140(.A(new_n3142_), .B(new_n3134_), .Y(new_n3143_));
  AND2X1   g02141(.A(new_n2983_), .B(new_n2981_), .Y(new_n3144_));
  OR2X1    g02142(.A(new_n2985_), .B(new_n3144_), .Y(new_n3145_));
  XOR2X1   g02143(.A(new_n2992_), .B(new_n3145_), .Y(new_n3146_));
  XOR2X1   g02144(.A(new_n2996_), .B(new_n2994_), .Y(new_n3147_));
  NOR2X1   g02145(.A(new_n2992_), .B(new_n2986_), .Y(new_n3148_));
  NOR2X1   g02146(.A(new_n2996_), .B(new_n2994_), .Y(new_n3149_));
  AOI21X1  g02147(.A0(new_n3148_), .A1(new_n3147_), .B0(new_n3149_), .Y(new_n3150_));
  XOR2X1   g02148(.A(new_n3148_), .B(new_n3147_), .Y(new_n3151_));
  OAI21X1  g02149(.A0(new_n3150_), .A1(new_n3146_), .B0(new_n3151_), .Y(new_n3152_));
  AND2X1   g02150(.A(new_n2965_), .B(new_n2963_), .Y(new_n3153_));
  OR2X1    g02151(.A(new_n2967_), .B(new_n3153_), .Y(new_n3154_));
  XOR2X1   g02152(.A(new_n2974_), .B(new_n3154_), .Y(new_n3155_));
  NOR4X1   g02153(.A(new_n2978_), .B(new_n2976_), .C(new_n2974_), .D(new_n2968_), .Y(new_n3156_));
  NOR4X1   g02154(.A(new_n2996_), .B(new_n2994_), .C(new_n2992_), .D(new_n2986_), .Y(new_n3157_));
  OR4X1    g02155(.A(new_n3157_), .B(new_n3146_), .C(new_n3156_), .D(new_n3155_), .Y(new_n3158_));
  XOR2X1   g02156(.A(new_n2978_), .B(new_n2976_), .Y(new_n3159_));
  NOR2X1   g02157(.A(new_n2974_), .B(new_n2968_), .Y(new_n3160_));
  NOR2X1   g02158(.A(new_n2978_), .B(new_n2976_), .Y(new_n3161_));
  AOI21X1  g02159(.A0(new_n3160_), .A1(new_n3159_), .B0(new_n3161_), .Y(new_n3162_));
  XOR2X1   g02160(.A(new_n3160_), .B(new_n3159_), .Y(new_n3163_));
  OAI21X1  g02161(.A0(new_n3162_), .A1(new_n3155_), .B0(new_n3163_), .Y(new_n3164_));
  XOR2X1   g02162(.A(new_n3164_), .B(new_n3158_), .Y(new_n3165_));
  NAND2X1  g02163(.A(new_n3165_), .B(new_n3152_), .Y(new_n3166_));
  XOR2X1   g02164(.A(new_n2992_), .B(new_n2986_), .Y(new_n3167_));
  AND2X1   g02165(.A(new_n2991_), .B(\A[576] ), .Y(new_n3168_));
  OR2X1    g02166(.A(new_n3168_), .B(new_n2993_), .Y(new_n3169_));
  XOR2X1   g02167(.A(new_n2996_), .B(new_n3169_), .Y(new_n3170_));
  OR2X1    g02168(.A(new_n2992_), .B(new_n2986_), .Y(new_n3171_));
  OR2X1    g02169(.A(new_n2996_), .B(new_n2994_), .Y(new_n3172_));
  OAI21X1  g02170(.A0(new_n3171_), .A1(new_n3170_), .B0(new_n3172_), .Y(new_n3173_));
  XOR2X1   g02171(.A(new_n3148_), .B(new_n3170_), .Y(new_n3174_));
  AOI21X1  g02172(.A0(new_n3173_), .A1(new_n3167_), .B0(new_n3174_), .Y(new_n3175_));
  AND2X1   g02173(.A(new_n3164_), .B(new_n3158_), .Y(new_n3176_));
  OR2X1    g02174(.A(new_n2974_), .B(new_n2968_), .Y(new_n3177_));
  XOR2X1   g02175(.A(new_n3177_), .B(new_n3159_), .Y(new_n3178_));
  OR4X1    g02176(.A(new_n3146_), .B(new_n3156_), .C(new_n3178_), .D(new_n3155_), .Y(new_n3179_));
  OAI22X1  g02177(.A0(new_n3174_), .A1(new_n3150_), .B0(new_n3162_), .B1(new_n3155_), .Y(new_n3180_));
  NOR2X1   g02178(.A(new_n3180_), .B(new_n3179_), .Y(new_n3181_));
  OAI21X1  g02179(.A0(new_n3181_), .A1(new_n3176_), .B0(new_n3175_), .Y(new_n3182_));
  NOR2X1   g02180(.A(new_n3037_), .B(new_n2999_), .Y(new_n3183_));
  NAND3X1  g02181(.A(new_n3183_), .B(new_n3182_), .C(new_n3166_), .Y(new_n3184_));
  AND2X1   g02182(.A(new_n3165_), .B(new_n3152_), .Y(new_n3185_));
  NAND2X1  g02183(.A(new_n3164_), .B(new_n3158_), .Y(new_n3186_));
  OR2X1    g02184(.A(new_n3180_), .B(new_n3179_), .Y(new_n3187_));
  AOI21X1  g02185(.A0(new_n3187_), .A1(new_n3186_), .B0(new_n3152_), .Y(new_n3188_));
  OR2X1    g02186(.A(new_n3037_), .B(new_n2999_), .Y(new_n3189_));
  OAI21X1  g02187(.A0(new_n3188_), .A1(new_n3185_), .B0(new_n3189_), .Y(new_n3190_));
  AND2X1   g02188(.A(new_n3022_), .B(new_n3020_), .Y(new_n3191_));
  OR2X1    g02189(.A(new_n3024_), .B(new_n3191_), .Y(new_n3192_));
  XOR2X1   g02190(.A(new_n3031_), .B(new_n3192_), .Y(new_n3193_));
  XOR2X1   g02191(.A(new_n3035_), .B(new_n3033_), .Y(new_n3194_));
  NOR2X1   g02192(.A(new_n3031_), .B(new_n3025_), .Y(new_n3195_));
  NOR2X1   g02193(.A(new_n3035_), .B(new_n3033_), .Y(new_n3196_));
  AOI21X1  g02194(.A0(new_n3195_), .A1(new_n3194_), .B0(new_n3196_), .Y(new_n3197_));
  XOR2X1   g02195(.A(new_n3195_), .B(new_n3194_), .Y(new_n3198_));
  OAI21X1  g02196(.A0(new_n3197_), .A1(new_n3193_), .B0(new_n3198_), .Y(new_n3199_));
  XOR2X1   g02197(.A(new_n3013_), .B(new_n3007_), .Y(new_n3200_));
  AOI21X1  g02198(.A0(new_n3003_), .A1(new_n3001_), .B0(new_n3006_), .Y(new_n3201_));
  NOR4X1   g02199(.A(new_n3017_), .B(new_n3015_), .C(new_n3013_), .D(new_n3201_), .Y(new_n3202_));
  NOR4X1   g02200(.A(new_n3035_), .B(new_n3033_), .C(new_n3031_), .D(new_n3025_), .Y(new_n3203_));
  OR4X1    g02201(.A(new_n3203_), .B(new_n3193_), .C(new_n3202_), .D(new_n3200_), .Y(new_n3204_));
  XOR2X1   g02202(.A(new_n3017_), .B(new_n3015_), .Y(new_n3205_));
  NOR2X1   g02203(.A(new_n3013_), .B(new_n3201_), .Y(new_n3206_));
  NOR2X1   g02204(.A(new_n3017_), .B(new_n3015_), .Y(new_n3207_));
  AOI21X1  g02205(.A0(new_n3206_), .A1(new_n3205_), .B0(new_n3207_), .Y(new_n3208_));
  XOR2X1   g02206(.A(new_n3206_), .B(new_n3205_), .Y(new_n3209_));
  OAI21X1  g02207(.A0(new_n3208_), .A1(new_n3200_), .B0(new_n3209_), .Y(new_n3210_));
  XOR2X1   g02208(.A(new_n3210_), .B(new_n3204_), .Y(new_n3211_));
  AND2X1   g02209(.A(new_n3210_), .B(new_n3204_), .Y(new_n3212_));
  OR2X1    g02210(.A(new_n3013_), .B(new_n3201_), .Y(new_n3213_));
  XOR2X1   g02211(.A(new_n3213_), .B(new_n3205_), .Y(new_n3214_));
  OR4X1    g02212(.A(new_n3193_), .B(new_n3202_), .C(new_n3214_), .D(new_n3200_), .Y(new_n3215_));
  OR4X1    g02213(.A(new_n3035_), .B(new_n3033_), .C(new_n3031_), .D(new_n3025_), .Y(new_n3216_));
  OAI21X1  g02214(.A0(new_n3208_), .A1(new_n3200_), .B0(new_n3216_), .Y(new_n3217_));
  NOR2X1   g02215(.A(new_n3217_), .B(new_n3215_), .Y(new_n3218_));
  OR2X1    g02216(.A(new_n3218_), .B(new_n3212_), .Y(new_n3219_));
  MX2X1    g02217(.A(new_n3219_), .B(new_n3211_), .S0(new_n3199_), .Y(new_n3220_));
  AOI21X1  g02218(.A0(new_n3190_), .A1(new_n3184_), .B0(new_n3220_), .Y(new_n3221_));
  INVX1    g02219(.A(new_n3199_), .Y(new_n3222_));
  AND2X1   g02220(.A(new_n3211_), .B(new_n3199_), .Y(new_n3223_));
  AOI21X1  g02221(.A0(new_n3219_), .A1(new_n3222_), .B0(new_n3223_), .Y(new_n3224_));
  NAND3X1  g02222(.A(new_n3189_), .B(new_n3182_), .C(new_n3166_), .Y(new_n3225_));
  OAI21X1  g02223(.A0(new_n3188_), .A1(new_n3185_), .B0(new_n3183_), .Y(new_n3226_));
  AOI21X1  g02224(.A0(new_n3226_), .A1(new_n3225_), .B0(new_n3224_), .Y(new_n3227_));
  NOR2X1   g02225(.A(new_n3227_), .B(new_n3221_), .Y(new_n3228_));
  NAND3X1  g02226(.A(new_n3141_), .B(new_n3131_), .C(new_n3127_), .Y(new_n3229_));
  OAI21X1  g02227(.A0(new_n3140_), .A1(new_n3137_), .B0(new_n3133_), .Y(new_n3230_));
  AND2X1   g02228(.A(new_n3230_), .B(new_n3229_), .Y(new_n3231_));
  MX2X1    g02229(.A(new_n3231_), .B(new_n3143_), .S0(new_n3228_), .Y(new_n3232_));
  AND2X1   g02230(.A(new_n2830_), .B(new_n2828_), .Y(new_n3233_));
  OR2X1    g02231(.A(new_n2832_), .B(new_n3233_), .Y(new_n3234_));
  XOR2X1   g02232(.A(new_n2839_), .B(new_n3234_), .Y(new_n3235_));
  XOR2X1   g02233(.A(new_n2843_), .B(new_n2841_), .Y(new_n3236_));
  NOR2X1   g02234(.A(new_n2839_), .B(new_n2833_), .Y(new_n3237_));
  NOR2X1   g02235(.A(new_n2843_), .B(new_n2841_), .Y(new_n3238_));
  AOI21X1  g02236(.A0(new_n3237_), .A1(new_n3236_), .B0(new_n3238_), .Y(new_n3239_));
  XOR2X1   g02237(.A(new_n3237_), .B(new_n3236_), .Y(new_n3240_));
  OAI21X1  g02238(.A0(new_n3239_), .A1(new_n3235_), .B0(new_n3240_), .Y(new_n3241_));
  AND2X1   g02239(.A(new_n2812_), .B(new_n2810_), .Y(new_n3242_));
  OR2X1    g02240(.A(new_n2814_), .B(new_n3242_), .Y(new_n3243_));
  XOR2X1   g02241(.A(new_n2821_), .B(new_n3243_), .Y(new_n3244_));
  NOR4X1   g02242(.A(new_n2825_), .B(new_n2823_), .C(new_n2821_), .D(new_n2815_), .Y(new_n3245_));
  NOR4X1   g02243(.A(new_n2843_), .B(new_n2841_), .C(new_n2839_), .D(new_n2833_), .Y(new_n3246_));
  OR4X1    g02244(.A(new_n3246_), .B(new_n3235_), .C(new_n3245_), .D(new_n3244_), .Y(new_n3247_));
  XOR2X1   g02245(.A(new_n2825_), .B(new_n2823_), .Y(new_n3248_));
  NOR2X1   g02246(.A(new_n2821_), .B(new_n2815_), .Y(new_n3249_));
  NOR2X1   g02247(.A(new_n2825_), .B(new_n2823_), .Y(new_n3250_));
  AOI21X1  g02248(.A0(new_n3249_), .A1(new_n3248_), .B0(new_n3250_), .Y(new_n3251_));
  XOR2X1   g02249(.A(new_n3249_), .B(new_n3248_), .Y(new_n3252_));
  OAI21X1  g02250(.A0(new_n3251_), .A1(new_n3244_), .B0(new_n3252_), .Y(new_n3253_));
  XOR2X1   g02251(.A(new_n3253_), .B(new_n3247_), .Y(new_n3254_));
  NAND2X1  g02252(.A(new_n3254_), .B(new_n3241_), .Y(new_n3255_));
  XOR2X1   g02253(.A(new_n2839_), .B(new_n2833_), .Y(new_n3256_));
  AND2X1   g02254(.A(new_n2838_), .B(\A[624] ), .Y(new_n3257_));
  OR2X1    g02255(.A(new_n3257_), .B(new_n2840_), .Y(new_n3258_));
  XOR2X1   g02256(.A(new_n2843_), .B(new_n3258_), .Y(new_n3259_));
  OR2X1    g02257(.A(new_n2839_), .B(new_n2833_), .Y(new_n3260_));
  OR2X1    g02258(.A(new_n2843_), .B(new_n2841_), .Y(new_n3261_));
  OAI21X1  g02259(.A0(new_n3260_), .A1(new_n3259_), .B0(new_n3261_), .Y(new_n3262_));
  XOR2X1   g02260(.A(new_n3237_), .B(new_n3259_), .Y(new_n3263_));
  AOI21X1  g02261(.A0(new_n3262_), .A1(new_n3256_), .B0(new_n3263_), .Y(new_n3264_));
  AND2X1   g02262(.A(new_n3253_), .B(new_n3247_), .Y(new_n3265_));
  OR2X1    g02263(.A(new_n2821_), .B(new_n2815_), .Y(new_n3266_));
  XOR2X1   g02264(.A(new_n3266_), .B(new_n3248_), .Y(new_n3267_));
  OR4X1    g02265(.A(new_n3235_), .B(new_n3245_), .C(new_n3267_), .D(new_n3244_), .Y(new_n3268_));
  OAI22X1  g02266(.A0(new_n3263_), .A1(new_n3239_), .B0(new_n3251_), .B1(new_n3244_), .Y(new_n3269_));
  NOR2X1   g02267(.A(new_n3269_), .B(new_n3268_), .Y(new_n3270_));
  OAI21X1  g02268(.A0(new_n3270_), .A1(new_n3265_), .B0(new_n3264_), .Y(new_n3271_));
  INVX1    g02269(.A(new_n2845_), .Y(new_n3272_));
  NOR2X1   g02270(.A(new_n2883_), .B(new_n3272_), .Y(new_n3273_));
  NAND3X1  g02271(.A(new_n3273_), .B(new_n3271_), .C(new_n3255_), .Y(new_n3274_));
  AND2X1   g02272(.A(new_n3254_), .B(new_n3241_), .Y(new_n3275_));
  NAND2X1  g02273(.A(new_n3253_), .B(new_n3247_), .Y(new_n3276_));
  OR2X1    g02274(.A(new_n3269_), .B(new_n3268_), .Y(new_n3277_));
  AOI21X1  g02275(.A0(new_n3277_), .A1(new_n3276_), .B0(new_n3241_), .Y(new_n3278_));
  OR2X1    g02276(.A(new_n2883_), .B(new_n3272_), .Y(new_n3279_));
  OAI21X1  g02277(.A0(new_n3278_), .A1(new_n3275_), .B0(new_n3279_), .Y(new_n3280_));
  AND2X1   g02278(.A(new_n2868_), .B(new_n2866_), .Y(new_n3281_));
  OR2X1    g02279(.A(new_n2870_), .B(new_n3281_), .Y(new_n3282_));
  XOR2X1   g02280(.A(new_n2877_), .B(new_n3282_), .Y(new_n3283_));
  XOR2X1   g02281(.A(new_n2881_), .B(new_n2879_), .Y(new_n3284_));
  NOR2X1   g02282(.A(new_n2877_), .B(new_n2871_), .Y(new_n3285_));
  NOR2X1   g02283(.A(new_n2881_), .B(new_n2879_), .Y(new_n3286_));
  AOI21X1  g02284(.A0(new_n3285_), .A1(new_n3284_), .B0(new_n3286_), .Y(new_n3287_));
  XOR2X1   g02285(.A(new_n3285_), .B(new_n3284_), .Y(new_n3288_));
  OAI21X1  g02286(.A0(new_n3287_), .A1(new_n3283_), .B0(new_n3288_), .Y(new_n3289_));
  XOR2X1   g02287(.A(new_n2859_), .B(new_n2853_), .Y(new_n3290_));
  AOI21X1  g02288(.A0(new_n2849_), .A1(new_n2847_), .B0(new_n2852_), .Y(new_n3291_));
  NOR4X1   g02289(.A(new_n2863_), .B(new_n2861_), .C(new_n2859_), .D(new_n3291_), .Y(new_n3292_));
  NOR4X1   g02290(.A(new_n2881_), .B(new_n2879_), .C(new_n2877_), .D(new_n2871_), .Y(new_n3293_));
  OR4X1    g02291(.A(new_n3293_), .B(new_n3283_), .C(new_n3292_), .D(new_n3290_), .Y(new_n3294_));
  XOR2X1   g02292(.A(new_n2863_), .B(new_n2861_), .Y(new_n3295_));
  NOR2X1   g02293(.A(new_n2859_), .B(new_n3291_), .Y(new_n3296_));
  NOR2X1   g02294(.A(new_n2863_), .B(new_n2861_), .Y(new_n3297_));
  AOI21X1  g02295(.A0(new_n3296_), .A1(new_n3295_), .B0(new_n3297_), .Y(new_n3298_));
  XOR2X1   g02296(.A(new_n3296_), .B(new_n3295_), .Y(new_n3299_));
  OAI21X1  g02297(.A0(new_n3298_), .A1(new_n3290_), .B0(new_n3299_), .Y(new_n3300_));
  XOR2X1   g02298(.A(new_n3300_), .B(new_n3294_), .Y(new_n3301_));
  AND2X1   g02299(.A(new_n3300_), .B(new_n3294_), .Y(new_n3302_));
  OR2X1    g02300(.A(new_n2859_), .B(new_n3291_), .Y(new_n3303_));
  XOR2X1   g02301(.A(new_n3303_), .B(new_n3295_), .Y(new_n3304_));
  OR4X1    g02302(.A(new_n3283_), .B(new_n3292_), .C(new_n3304_), .D(new_n3290_), .Y(new_n3305_));
  OR4X1    g02303(.A(new_n2881_), .B(new_n2879_), .C(new_n2877_), .D(new_n2871_), .Y(new_n3306_));
  OAI21X1  g02304(.A0(new_n3298_), .A1(new_n3290_), .B0(new_n3306_), .Y(new_n3307_));
  NOR2X1   g02305(.A(new_n3307_), .B(new_n3305_), .Y(new_n3308_));
  OR2X1    g02306(.A(new_n3308_), .B(new_n3302_), .Y(new_n3309_));
  MX2X1    g02307(.A(new_n3309_), .B(new_n3301_), .S0(new_n3289_), .Y(new_n3310_));
  AOI21X1  g02308(.A0(new_n3280_), .A1(new_n3274_), .B0(new_n3310_), .Y(new_n3311_));
  INVX1    g02309(.A(new_n3289_), .Y(new_n3312_));
  AND2X1   g02310(.A(new_n3301_), .B(new_n3289_), .Y(new_n3313_));
  AOI21X1  g02311(.A0(new_n3309_), .A1(new_n3312_), .B0(new_n3313_), .Y(new_n3314_));
  NAND3X1  g02312(.A(new_n3279_), .B(new_n3271_), .C(new_n3255_), .Y(new_n3315_));
  OAI21X1  g02313(.A0(new_n3278_), .A1(new_n3275_), .B0(new_n3273_), .Y(new_n3316_));
  AOI21X1  g02314(.A0(new_n3316_), .A1(new_n3315_), .B0(new_n3314_), .Y(new_n3317_));
  OR2X1    g02315(.A(new_n3317_), .B(new_n3311_), .Y(new_n3318_));
  AND2X1   g02316(.A(new_n2792_), .B(new_n2790_), .Y(new_n3319_));
  OR2X1    g02317(.A(new_n2794_), .B(new_n3319_), .Y(new_n3320_));
  XOR2X1   g02318(.A(new_n2801_), .B(new_n3320_), .Y(new_n3321_));
  XOR2X1   g02319(.A(new_n2805_), .B(new_n2803_), .Y(new_n3322_));
  NOR2X1   g02320(.A(new_n2801_), .B(new_n2795_), .Y(new_n3323_));
  NOR2X1   g02321(.A(new_n2805_), .B(new_n2803_), .Y(new_n3324_));
  AOI21X1  g02322(.A0(new_n3323_), .A1(new_n3322_), .B0(new_n3324_), .Y(new_n3325_));
  XOR2X1   g02323(.A(new_n3323_), .B(new_n3322_), .Y(new_n3326_));
  OAI21X1  g02324(.A0(new_n3325_), .A1(new_n3321_), .B0(new_n3326_), .Y(new_n3327_));
  INVX1    g02325(.A(new_n3327_), .Y(new_n3328_));
  XOR2X1   g02326(.A(new_n2783_), .B(new_n2777_), .Y(new_n3329_));
  AOI21X1  g02327(.A0(new_n2773_), .A1(new_n2771_), .B0(new_n2776_), .Y(new_n3330_));
  NOR4X1   g02328(.A(new_n2787_), .B(new_n2785_), .C(new_n2783_), .D(new_n3330_), .Y(new_n3331_));
  NOR4X1   g02329(.A(new_n2805_), .B(new_n2803_), .C(new_n2801_), .D(new_n2795_), .Y(new_n3332_));
  OR4X1    g02330(.A(new_n3332_), .B(new_n3321_), .C(new_n3331_), .D(new_n3329_), .Y(new_n3333_));
  XOR2X1   g02331(.A(new_n2787_), .B(new_n2785_), .Y(new_n3334_));
  NOR2X1   g02332(.A(new_n2783_), .B(new_n3330_), .Y(new_n3335_));
  NOR2X1   g02333(.A(new_n2787_), .B(new_n2785_), .Y(new_n3336_));
  AOI21X1  g02334(.A0(new_n3335_), .A1(new_n3334_), .B0(new_n3336_), .Y(new_n3337_));
  XOR2X1   g02335(.A(new_n3335_), .B(new_n3334_), .Y(new_n3338_));
  OAI21X1  g02336(.A0(new_n3337_), .A1(new_n3329_), .B0(new_n3338_), .Y(new_n3339_));
  XOR2X1   g02337(.A(new_n3339_), .B(new_n3333_), .Y(new_n3340_));
  AND2X1   g02338(.A(new_n3340_), .B(new_n3327_), .Y(new_n3341_));
  AND2X1   g02339(.A(new_n3339_), .B(new_n3333_), .Y(new_n3342_));
  OR2X1    g02340(.A(new_n2783_), .B(new_n3330_), .Y(new_n3343_));
  XOR2X1   g02341(.A(new_n3343_), .B(new_n3334_), .Y(new_n3344_));
  OR4X1    g02342(.A(new_n3321_), .B(new_n3331_), .C(new_n3344_), .D(new_n3329_), .Y(new_n3345_));
  OR4X1    g02343(.A(new_n2805_), .B(new_n2803_), .C(new_n2801_), .D(new_n2795_), .Y(new_n3346_));
  OAI21X1  g02344(.A0(new_n3337_), .A1(new_n3329_), .B0(new_n3346_), .Y(new_n3347_));
  NOR2X1   g02345(.A(new_n3347_), .B(new_n3345_), .Y(new_n3348_));
  OR2X1    g02346(.A(new_n3348_), .B(new_n3342_), .Y(new_n3349_));
  AOI21X1  g02347(.A0(new_n3349_), .A1(new_n3328_), .B0(new_n3341_), .Y(new_n3350_));
  AND2X1   g02348(.A(new_n2754_), .B(new_n2752_), .Y(new_n3351_));
  OR2X1    g02349(.A(new_n2756_), .B(new_n3351_), .Y(new_n3352_));
  XOR2X1   g02350(.A(new_n2763_), .B(new_n3352_), .Y(new_n3353_));
  XOR2X1   g02351(.A(new_n2767_), .B(new_n2765_), .Y(new_n3354_));
  NOR2X1   g02352(.A(new_n2763_), .B(new_n2757_), .Y(new_n3355_));
  NOR2X1   g02353(.A(new_n2767_), .B(new_n2765_), .Y(new_n3356_));
  AOI21X1  g02354(.A0(new_n3355_), .A1(new_n3354_), .B0(new_n3356_), .Y(new_n3357_));
  XOR2X1   g02355(.A(new_n3355_), .B(new_n3354_), .Y(new_n3358_));
  OAI21X1  g02356(.A0(new_n3357_), .A1(new_n3353_), .B0(new_n3358_), .Y(new_n3359_));
  AND2X1   g02357(.A(new_n2736_), .B(new_n2734_), .Y(new_n3360_));
  OR2X1    g02358(.A(new_n2738_), .B(new_n3360_), .Y(new_n3361_));
  XOR2X1   g02359(.A(new_n2745_), .B(new_n3361_), .Y(new_n3362_));
  NOR4X1   g02360(.A(new_n2749_), .B(new_n2747_), .C(new_n2745_), .D(new_n2739_), .Y(new_n3363_));
  NOR4X1   g02361(.A(new_n2767_), .B(new_n2765_), .C(new_n2763_), .D(new_n2757_), .Y(new_n3364_));
  OR4X1    g02362(.A(new_n3364_), .B(new_n3353_), .C(new_n3363_), .D(new_n3362_), .Y(new_n3365_));
  XOR2X1   g02363(.A(new_n2749_), .B(new_n2747_), .Y(new_n3366_));
  NOR2X1   g02364(.A(new_n2745_), .B(new_n2739_), .Y(new_n3367_));
  NOR2X1   g02365(.A(new_n2749_), .B(new_n2747_), .Y(new_n3368_));
  AOI21X1  g02366(.A0(new_n3367_), .A1(new_n3366_), .B0(new_n3368_), .Y(new_n3369_));
  XOR2X1   g02367(.A(new_n3367_), .B(new_n3366_), .Y(new_n3370_));
  OAI21X1  g02368(.A0(new_n3369_), .A1(new_n3362_), .B0(new_n3370_), .Y(new_n3371_));
  XOR2X1   g02369(.A(new_n3371_), .B(new_n3365_), .Y(new_n3372_));
  AND2X1   g02370(.A(new_n3372_), .B(new_n3359_), .Y(new_n3373_));
  NAND2X1  g02371(.A(new_n3371_), .B(new_n3365_), .Y(new_n3374_));
  OR2X1    g02372(.A(new_n2745_), .B(new_n2739_), .Y(new_n3375_));
  XOR2X1   g02373(.A(new_n3375_), .B(new_n3366_), .Y(new_n3376_));
  OR4X1    g02374(.A(new_n3353_), .B(new_n3363_), .C(new_n3376_), .D(new_n3362_), .Y(new_n3377_));
  AND2X1   g02375(.A(new_n2762_), .B(\A[648] ), .Y(new_n3378_));
  OR2X1    g02376(.A(new_n3378_), .B(new_n2764_), .Y(new_n3379_));
  XOR2X1   g02377(.A(new_n2767_), .B(new_n3379_), .Y(new_n3380_));
  XOR2X1   g02378(.A(new_n3355_), .B(new_n3380_), .Y(new_n3381_));
  OAI22X1  g02379(.A0(new_n3381_), .A1(new_n3357_), .B0(new_n3369_), .B1(new_n3362_), .Y(new_n3382_));
  OR2X1    g02380(.A(new_n3382_), .B(new_n3377_), .Y(new_n3383_));
  AOI21X1  g02381(.A0(new_n3383_), .A1(new_n3374_), .B0(new_n3359_), .Y(new_n3384_));
  INVX1    g02382(.A(new_n2769_), .Y(new_n3385_));
  OR2X1    g02383(.A(new_n2807_), .B(new_n3385_), .Y(new_n3386_));
  NOR3X1   g02384(.A(new_n3386_), .B(new_n3384_), .C(new_n3373_), .Y(new_n3387_));
  NAND2X1  g02385(.A(new_n3372_), .B(new_n3359_), .Y(new_n3388_));
  XOR2X1   g02386(.A(new_n2763_), .B(new_n2757_), .Y(new_n3389_));
  OR2X1    g02387(.A(new_n2763_), .B(new_n2757_), .Y(new_n3390_));
  OR2X1    g02388(.A(new_n2767_), .B(new_n2765_), .Y(new_n3391_));
  OAI21X1  g02389(.A0(new_n3390_), .A1(new_n3380_), .B0(new_n3391_), .Y(new_n3392_));
  AOI21X1  g02390(.A0(new_n3392_), .A1(new_n3389_), .B0(new_n3381_), .Y(new_n3393_));
  AND2X1   g02391(.A(new_n3371_), .B(new_n3365_), .Y(new_n3394_));
  NOR2X1   g02392(.A(new_n3382_), .B(new_n3377_), .Y(new_n3395_));
  OAI21X1  g02393(.A0(new_n3395_), .A1(new_n3394_), .B0(new_n3393_), .Y(new_n3396_));
  NOR2X1   g02394(.A(new_n2807_), .B(new_n3385_), .Y(new_n3397_));
  AOI21X1  g02395(.A0(new_n3396_), .A1(new_n3388_), .B0(new_n3397_), .Y(new_n3398_));
  OAI21X1  g02396(.A0(new_n3398_), .A1(new_n3387_), .B0(new_n3350_), .Y(new_n3399_));
  MX2X1    g02397(.A(new_n3349_), .B(new_n3340_), .S0(new_n3327_), .Y(new_n3400_));
  NOR3X1   g02398(.A(new_n3397_), .B(new_n3384_), .C(new_n3373_), .Y(new_n3401_));
  AOI21X1  g02399(.A0(new_n3396_), .A1(new_n3388_), .B0(new_n3386_), .Y(new_n3402_));
  OAI21X1  g02400(.A0(new_n3402_), .A1(new_n3401_), .B0(new_n3400_), .Y(new_n3403_));
  NOR2X1   g02401(.A(new_n2884_), .B(new_n2808_), .Y(new_n3404_));
  NAND3X1  g02402(.A(new_n3404_), .B(new_n3403_), .C(new_n3399_), .Y(new_n3405_));
  NAND3X1  g02403(.A(new_n3397_), .B(new_n3396_), .C(new_n3388_), .Y(new_n3406_));
  OAI21X1  g02404(.A0(new_n3384_), .A1(new_n3373_), .B0(new_n3386_), .Y(new_n3407_));
  AOI21X1  g02405(.A0(new_n3407_), .A1(new_n3406_), .B0(new_n3400_), .Y(new_n3408_));
  NAND3X1  g02406(.A(new_n3386_), .B(new_n3396_), .C(new_n3388_), .Y(new_n3409_));
  OAI21X1  g02407(.A0(new_n3384_), .A1(new_n3373_), .B0(new_n3397_), .Y(new_n3410_));
  AOI21X1  g02408(.A0(new_n3410_), .A1(new_n3409_), .B0(new_n3350_), .Y(new_n3411_));
  INVX1    g02409(.A(new_n3404_), .Y(new_n3412_));
  OAI21X1  g02410(.A0(new_n3411_), .A1(new_n3408_), .B0(new_n3412_), .Y(new_n3413_));
  AOI21X1  g02411(.A0(new_n3413_), .A1(new_n3405_), .B0(new_n3318_), .Y(new_n3414_));
  NOR2X1   g02412(.A(new_n3317_), .B(new_n3311_), .Y(new_n3415_));
  NAND3X1  g02413(.A(new_n3412_), .B(new_n3403_), .C(new_n3399_), .Y(new_n3416_));
  OAI21X1  g02414(.A0(new_n3411_), .A1(new_n3408_), .B0(new_n3404_), .Y(new_n3417_));
  AOI21X1  g02415(.A0(new_n3417_), .A1(new_n3416_), .B0(new_n3415_), .Y(new_n3418_));
  INVX1    g02416(.A(new_n2885_), .Y(new_n3419_));
  NOR2X1   g02417(.A(new_n3039_), .B(new_n3419_), .Y(new_n3420_));
  INVX1    g02418(.A(new_n3420_), .Y(new_n3421_));
  NOR3X1   g02419(.A(new_n3421_), .B(new_n3418_), .C(new_n3414_), .Y(new_n3422_));
  NOR3X1   g02420(.A(new_n3412_), .B(new_n3411_), .C(new_n3408_), .Y(new_n3423_));
  AOI21X1  g02421(.A0(new_n3403_), .A1(new_n3399_), .B0(new_n3404_), .Y(new_n3424_));
  OAI21X1  g02422(.A0(new_n3424_), .A1(new_n3423_), .B0(new_n3415_), .Y(new_n3425_));
  NOR3X1   g02423(.A(new_n3404_), .B(new_n3411_), .C(new_n3408_), .Y(new_n3426_));
  AOI21X1  g02424(.A0(new_n3403_), .A1(new_n3399_), .B0(new_n3412_), .Y(new_n3427_));
  OAI21X1  g02425(.A0(new_n3427_), .A1(new_n3426_), .B0(new_n3318_), .Y(new_n3428_));
  AOI21X1  g02426(.A0(new_n3428_), .A1(new_n3425_), .B0(new_n3420_), .Y(new_n3429_));
  OAI21X1  g02427(.A0(new_n3429_), .A1(new_n3422_), .B0(new_n3232_), .Y(new_n3430_));
  OR2X1    g02428(.A(new_n3227_), .B(new_n3221_), .Y(new_n3431_));
  NOR3X1   g02429(.A(new_n3133_), .B(new_n3140_), .C(new_n3137_), .Y(new_n3432_));
  AOI21X1  g02430(.A0(new_n3131_), .A1(new_n3127_), .B0(new_n3141_), .Y(new_n3433_));
  OAI21X1  g02431(.A0(new_n3433_), .A1(new_n3432_), .B0(new_n3431_), .Y(new_n3434_));
  OAI21X1  g02432(.A0(new_n3431_), .A1(new_n3143_), .B0(new_n3434_), .Y(new_n3435_));
  NOR3X1   g02433(.A(new_n3420_), .B(new_n3418_), .C(new_n3414_), .Y(new_n3436_));
  AOI21X1  g02434(.A0(new_n3428_), .A1(new_n3425_), .B0(new_n3421_), .Y(new_n3437_));
  OAI21X1  g02435(.A0(new_n3437_), .A1(new_n3436_), .B0(new_n3435_), .Y(new_n3438_));
  INVX1    g02436(.A(new_n3040_), .Y(new_n3439_));
  AND2X1   g02437(.A(new_n3439_), .B(new_n2732_), .Y(new_n3440_));
  NAND3X1  g02438(.A(new_n3440_), .B(new_n3438_), .C(new_n3430_), .Y(new_n3441_));
  NAND3X1  g02439(.A(new_n3420_), .B(new_n3428_), .C(new_n3425_), .Y(new_n3442_));
  OAI21X1  g02440(.A0(new_n3418_), .A1(new_n3414_), .B0(new_n3421_), .Y(new_n3443_));
  AOI21X1  g02441(.A0(new_n3443_), .A1(new_n3442_), .B0(new_n3435_), .Y(new_n3444_));
  NAND3X1  g02442(.A(new_n3421_), .B(new_n3428_), .C(new_n3425_), .Y(new_n3445_));
  OAI21X1  g02443(.A0(new_n3418_), .A1(new_n3414_), .B0(new_n3420_), .Y(new_n3446_));
  AOI21X1  g02444(.A0(new_n3446_), .A1(new_n3445_), .B0(new_n3232_), .Y(new_n3447_));
  INVX1    g02445(.A(new_n3440_), .Y(new_n3448_));
  OAI21X1  g02446(.A0(new_n3447_), .A1(new_n3444_), .B0(new_n3448_), .Y(new_n3449_));
  AND2X1   g02447(.A(new_n3449_), .B(new_n3441_), .Y(new_n3450_));
  AND2X1   g02448(.A(new_n2675_), .B(new_n2673_), .Y(new_n3451_));
  OR2X1    g02449(.A(new_n2677_), .B(new_n3451_), .Y(new_n3452_));
  XOR2X1   g02450(.A(new_n2684_), .B(new_n3452_), .Y(new_n3453_));
  XOR2X1   g02451(.A(new_n2688_), .B(new_n2686_), .Y(new_n3454_));
  NOR2X1   g02452(.A(new_n2684_), .B(new_n2678_), .Y(new_n3455_));
  NOR2X1   g02453(.A(new_n2688_), .B(new_n2686_), .Y(new_n3456_));
  AOI21X1  g02454(.A0(new_n3455_), .A1(new_n3454_), .B0(new_n3456_), .Y(new_n3457_));
  XOR2X1   g02455(.A(new_n3455_), .B(new_n3454_), .Y(new_n3458_));
  OAI21X1  g02456(.A0(new_n3457_), .A1(new_n3453_), .B0(new_n3458_), .Y(new_n3459_));
  AND2X1   g02457(.A(new_n2657_), .B(new_n2655_), .Y(new_n3460_));
  OR2X1    g02458(.A(new_n2659_), .B(new_n3460_), .Y(new_n3461_));
  XOR2X1   g02459(.A(new_n2666_), .B(new_n3461_), .Y(new_n3462_));
  NOR4X1   g02460(.A(new_n2670_), .B(new_n2668_), .C(new_n2666_), .D(new_n2660_), .Y(new_n3463_));
  NOR4X1   g02461(.A(new_n2688_), .B(new_n2686_), .C(new_n2684_), .D(new_n2678_), .Y(new_n3464_));
  OR4X1    g02462(.A(new_n3464_), .B(new_n3453_), .C(new_n3463_), .D(new_n3462_), .Y(new_n3465_));
  XOR2X1   g02463(.A(new_n2670_), .B(new_n2668_), .Y(new_n3466_));
  NOR2X1   g02464(.A(new_n2666_), .B(new_n2660_), .Y(new_n3467_));
  NOR2X1   g02465(.A(new_n2670_), .B(new_n2668_), .Y(new_n3468_));
  AOI21X1  g02466(.A0(new_n3467_), .A1(new_n3466_), .B0(new_n3468_), .Y(new_n3469_));
  XOR2X1   g02467(.A(new_n3467_), .B(new_n3466_), .Y(new_n3470_));
  OAI21X1  g02468(.A0(new_n3469_), .A1(new_n3462_), .B0(new_n3470_), .Y(new_n3471_));
  XOR2X1   g02469(.A(new_n3471_), .B(new_n3465_), .Y(new_n3472_));
  NAND2X1  g02470(.A(new_n3472_), .B(new_n3459_), .Y(new_n3473_));
  XOR2X1   g02471(.A(new_n2684_), .B(new_n2678_), .Y(new_n3474_));
  AND2X1   g02472(.A(new_n2683_), .B(\A[528] ), .Y(new_n3475_));
  OR2X1    g02473(.A(new_n3475_), .B(new_n2685_), .Y(new_n3476_));
  XOR2X1   g02474(.A(new_n2688_), .B(new_n3476_), .Y(new_n3477_));
  OR2X1    g02475(.A(new_n2684_), .B(new_n2678_), .Y(new_n3478_));
  OR2X1    g02476(.A(new_n2688_), .B(new_n2686_), .Y(new_n3479_));
  OAI21X1  g02477(.A0(new_n3478_), .A1(new_n3477_), .B0(new_n3479_), .Y(new_n3480_));
  XOR2X1   g02478(.A(new_n3455_), .B(new_n3477_), .Y(new_n3481_));
  AOI21X1  g02479(.A0(new_n3480_), .A1(new_n3474_), .B0(new_n3481_), .Y(new_n3482_));
  AND2X1   g02480(.A(new_n3471_), .B(new_n3465_), .Y(new_n3483_));
  OR2X1    g02481(.A(new_n2666_), .B(new_n2660_), .Y(new_n3484_));
  XOR2X1   g02482(.A(new_n3484_), .B(new_n3466_), .Y(new_n3485_));
  OR4X1    g02483(.A(new_n3453_), .B(new_n3463_), .C(new_n3485_), .D(new_n3462_), .Y(new_n3486_));
  OAI22X1  g02484(.A0(new_n3481_), .A1(new_n3457_), .B0(new_n3469_), .B1(new_n3462_), .Y(new_n3487_));
  NOR2X1   g02485(.A(new_n3487_), .B(new_n3486_), .Y(new_n3488_));
  OAI21X1  g02486(.A0(new_n3488_), .A1(new_n3483_), .B0(new_n3482_), .Y(new_n3489_));
  NOR2X1   g02487(.A(new_n2729_), .B(new_n2691_), .Y(new_n3490_));
  NAND3X1  g02488(.A(new_n3490_), .B(new_n3489_), .C(new_n3473_), .Y(new_n3491_));
  AND2X1   g02489(.A(new_n3472_), .B(new_n3459_), .Y(new_n3492_));
  NAND2X1  g02490(.A(new_n3471_), .B(new_n3465_), .Y(new_n3493_));
  OR2X1    g02491(.A(new_n3487_), .B(new_n3486_), .Y(new_n3494_));
  AOI21X1  g02492(.A0(new_n3494_), .A1(new_n3493_), .B0(new_n3459_), .Y(new_n3495_));
  OR2X1    g02493(.A(new_n2729_), .B(new_n2691_), .Y(new_n3496_));
  OAI21X1  g02494(.A0(new_n3495_), .A1(new_n3492_), .B0(new_n3496_), .Y(new_n3497_));
  AND2X1   g02495(.A(new_n2714_), .B(new_n2712_), .Y(new_n3498_));
  OR2X1    g02496(.A(new_n2716_), .B(new_n3498_), .Y(new_n3499_));
  XOR2X1   g02497(.A(new_n2723_), .B(new_n3499_), .Y(new_n3500_));
  XOR2X1   g02498(.A(new_n2727_), .B(new_n2725_), .Y(new_n3501_));
  NOR2X1   g02499(.A(new_n2723_), .B(new_n2717_), .Y(new_n3502_));
  NOR2X1   g02500(.A(new_n2727_), .B(new_n2725_), .Y(new_n3503_));
  AOI21X1  g02501(.A0(new_n3502_), .A1(new_n3501_), .B0(new_n3503_), .Y(new_n3504_));
  XOR2X1   g02502(.A(new_n3502_), .B(new_n3501_), .Y(new_n3505_));
  OAI21X1  g02503(.A0(new_n3504_), .A1(new_n3500_), .B0(new_n3505_), .Y(new_n3506_));
  XOR2X1   g02504(.A(new_n2705_), .B(new_n2699_), .Y(new_n3507_));
  AOI21X1  g02505(.A0(new_n2695_), .A1(new_n2693_), .B0(new_n2698_), .Y(new_n3508_));
  NOR4X1   g02506(.A(new_n2709_), .B(new_n2707_), .C(new_n2705_), .D(new_n3508_), .Y(new_n3509_));
  NOR4X1   g02507(.A(new_n2727_), .B(new_n2725_), .C(new_n2723_), .D(new_n2717_), .Y(new_n3510_));
  OR4X1    g02508(.A(new_n3510_), .B(new_n3500_), .C(new_n3509_), .D(new_n3507_), .Y(new_n3511_));
  XOR2X1   g02509(.A(new_n2709_), .B(new_n2707_), .Y(new_n3512_));
  NOR2X1   g02510(.A(new_n2705_), .B(new_n3508_), .Y(new_n3513_));
  NOR2X1   g02511(.A(new_n2709_), .B(new_n2707_), .Y(new_n3514_));
  AOI21X1  g02512(.A0(new_n3513_), .A1(new_n3512_), .B0(new_n3514_), .Y(new_n3515_));
  XOR2X1   g02513(.A(new_n3513_), .B(new_n3512_), .Y(new_n3516_));
  OAI21X1  g02514(.A0(new_n3515_), .A1(new_n3507_), .B0(new_n3516_), .Y(new_n3517_));
  XOR2X1   g02515(.A(new_n3517_), .B(new_n3511_), .Y(new_n3518_));
  AND2X1   g02516(.A(new_n3517_), .B(new_n3511_), .Y(new_n3519_));
  OR2X1    g02517(.A(new_n2705_), .B(new_n3508_), .Y(new_n3520_));
  XOR2X1   g02518(.A(new_n3520_), .B(new_n3512_), .Y(new_n3521_));
  OR4X1    g02519(.A(new_n3500_), .B(new_n3509_), .C(new_n3521_), .D(new_n3507_), .Y(new_n3522_));
  OR4X1    g02520(.A(new_n2727_), .B(new_n2725_), .C(new_n2723_), .D(new_n2717_), .Y(new_n3523_));
  OAI21X1  g02521(.A0(new_n3515_), .A1(new_n3507_), .B0(new_n3523_), .Y(new_n3524_));
  NOR2X1   g02522(.A(new_n3524_), .B(new_n3522_), .Y(new_n3525_));
  OR2X1    g02523(.A(new_n3525_), .B(new_n3519_), .Y(new_n3526_));
  MX2X1    g02524(.A(new_n3526_), .B(new_n3518_), .S0(new_n3506_), .Y(new_n3527_));
  AOI21X1  g02525(.A0(new_n3497_), .A1(new_n3491_), .B0(new_n3527_), .Y(new_n3528_));
  INVX1    g02526(.A(new_n3506_), .Y(new_n3529_));
  AND2X1   g02527(.A(new_n3518_), .B(new_n3506_), .Y(new_n3530_));
  AOI21X1  g02528(.A0(new_n3526_), .A1(new_n3529_), .B0(new_n3530_), .Y(new_n3531_));
  NAND3X1  g02529(.A(new_n3496_), .B(new_n3489_), .C(new_n3473_), .Y(new_n3532_));
  OAI21X1  g02530(.A0(new_n3495_), .A1(new_n3492_), .B0(new_n3490_), .Y(new_n3533_));
  AOI21X1  g02531(.A0(new_n3533_), .A1(new_n3532_), .B0(new_n3531_), .Y(new_n3534_));
  NOR2X1   g02532(.A(new_n3534_), .B(new_n3528_), .Y(new_n3535_));
  AND2X1   g02533(.A(new_n2637_), .B(new_n2635_), .Y(new_n3536_));
  OR2X1    g02534(.A(new_n2639_), .B(new_n3536_), .Y(new_n3537_));
  XOR2X1   g02535(.A(new_n2646_), .B(new_n3537_), .Y(new_n3538_));
  XOR2X1   g02536(.A(new_n2650_), .B(new_n2648_), .Y(new_n3539_));
  NOR2X1   g02537(.A(new_n2646_), .B(new_n2640_), .Y(new_n3540_));
  NOR2X1   g02538(.A(new_n2650_), .B(new_n2648_), .Y(new_n3541_));
  AOI21X1  g02539(.A0(new_n3540_), .A1(new_n3539_), .B0(new_n3541_), .Y(new_n3542_));
  XOR2X1   g02540(.A(new_n3540_), .B(new_n3539_), .Y(new_n3543_));
  OAI21X1  g02541(.A0(new_n3542_), .A1(new_n3538_), .B0(new_n3543_), .Y(new_n3544_));
  XOR2X1   g02542(.A(new_n2628_), .B(new_n2622_), .Y(new_n3545_));
  AOI21X1  g02543(.A0(new_n2618_), .A1(new_n2616_), .B0(new_n2621_), .Y(new_n3546_));
  NOR4X1   g02544(.A(new_n2632_), .B(new_n2630_), .C(new_n2628_), .D(new_n3546_), .Y(new_n3547_));
  NOR4X1   g02545(.A(new_n2650_), .B(new_n2648_), .C(new_n2646_), .D(new_n2640_), .Y(new_n3548_));
  OR4X1    g02546(.A(new_n3548_), .B(new_n3538_), .C(new_n3547_), .D(new_n3545_), .Y(new_n3549_));
  XOR2X1   g02547(.A(new_n2632_), .B(new_n2630_), .Y(new_n3550_));
  NOR2X1   g02548(.A(new_n2628_), .B(new_n3546_), .Y(new_n3551_));
  NOR2X1   g02549(.A(new_n2632_), .B(new_n2630_), .Y(new_n3552_));
  AOI21X1  g02550(.A0(new_n3551_), .A1(new_n3550_), .B0(new_n3552_), .Y(new_n3553_));
  XOR2X1   g02551(.A(new_n3551_), .B(new_n3550_), .Y(new_n3554_));
  OAI21X1  g02552(.A0(new_n3553_), .A1(new_n3545_), .B0(new_n3554_), .Y(new_n3555_));
  XOR2X1   g02553(.A(new_n3555_), .B(new_n3549_), .Y(new_n3556_));
  AND2X1   g02554(.A(new_n3555_), .B(new_n3549_), .Y(new_n3557_));
  OR2X1    g02555(.A(new_n2628_), .B(new_n3546_), .Y(new_n3558_));
  XOR2X1   g02556(.A(new_n3558_), .B(new_n3550_), .Y(new_n3559_));
  OR4X1    g02557(.A(new_n3538_), .B(new_n3547_), .C(new_n3559_), .D(new_n3545_), .Y(new_n3560_));
  OR4X1    g02558(.A(new_n2650_), .B(new_n2648_), .C(new_n2646_), .D(new_n2640_), .Y(new_n3561_));
  OAI21X1  g02559(.A0(new_n3553_), .A1(new_n3545_), .B0(new_n3561_), .Y(new_n3562_));
  NOR2X1   g02560(.A(new_n3562_), .B(new_n3560_), .Y(new_n3563_));
  OR2X1    g02561(.A(new_n3563_), .B(new_n3557_), .Y(new_n3564_));
  MX2X1    g02562(.A(new_n3564_), .B(new_n3556_), .S0(new_n3544_), .Y(new_n3565_));
  AND2X1   g02563(.A(new_n2599_), .B(new_n2597_), .Y(new_n3566_));
  OR2X1    g02564(.A(new_n2601_), .B(new_n3566_), .Y(new_n3567_));
  XOR2X1   g02565(.A(new_n2608_), .B(new_n3567_), .Y(new_n3568_));
  XOR2X1   g02566(.A(new_n2612_), .B(new_n2610_), .Y(new_n3569_));
  NOR2X1   g02567(.A(new_n2608_), .B(new_n2602_), .Y(new_n3570_));
  NOR2X1   g02568(.A(new_n2612_), .B(new_n2610_), .Y(new_n3571_));
  AOI21X1  g02569(.A0(new_n3570_), .A1(new_n3569_), .B0(new_n3571_), .Y(new_n3572_));
  XOR2X1   g02570(.A(new_n3570_), .B(new_n3569_), .Y(new_n3573_));
  OAI21X1  g02571(.A0(new_n3572_), .A1(new_n3568_), .B0(new_n3573_), .Y(new_n3574_));
  AND2X1   g02572(.A(new_n2581_), .B(new_n2579_), .Y(new_n3575_));
  OR2X1    g02573(.A(new_n2583_), .B(new_n3575_), .Y(new_n3576_));
  XOR2X1   g02574(.A(new_n2590_), .B(new_n3576_), .Y(new_n3577_));
  NOR4X1   g02575(.A(new_n2594_), .B(new_n2592_), .C(new_n2590_), .D(new_n2584_), .Y(new_n3578_));
  NOR4X1   g02576(.A(new_n2612_), .B(new_n2610_), .C(new_n2608_), .D(new_n2602_), .Y(new_n3579_));
  OR4X1    g02577(.A(new_n3579_), .B(new_n3568_), .C(new_n3578_), .D(new_n3577_), .Y(new_n3580_));
  XOR2X1   g02578(.A(new_n2594_), .B(new_n2592_), .Y(new_n3581_));
  NOR2X1   g02579(.A(new_n2590_), .B(new_n2584_), .Y(new_n3582_));
  NOR2X1   g02580(.A(new_n2594_), .B(new_n2592_), .Y(new_n3583_));
  AOI21X1  g02581(.A0(new_n3582_), .A1(new_n3581_), .B0(new_n3583_), .Y(new_n3584_));
  XOR2X1   g02582(.A(new_n3582_), .B(new_n3581_), .Y(new_n3585_));
  OAI21X1  g02583(.A0(new_n3584_), .A1(new_n3577_), .B0(new_n3585_), .Y(new_n3586_));
  XOR2X1   g02584(.A(new_n3586_), .B(new_n3580_), .Y(new_n3587_));
  NAND2X1  g02585(.A(new_n3587_), .B(new_n3574_), .Y(new_n3588_));
  XOR2X1   g02586(.A(new_n2608_), .B(new_n2602_), .Y(new_n3589_));
  AND2X1   g02587(.A(new_n2607_), .B(\A[552] ), .Y(new_n3590_));
  OR2X1    g02588(.A(new_n3590_), .B(new_n2609_), .Y(new_n3591_));
  XOR2X1   g02589(.A(new_n2612_), .B(new_n3591_), .Y(new_n3592_));
  OR2X1    g02590(.A(new_n2608_), .B(new_n2602_), .Y(new_n3593_));
  OR2X1    g02591(.A(new_n2612_), .B(new_n2610_), .Y(new_n3594_));
  OAI21X1  g02592(.A0(new_n3593_), .A1(new_n3592_), .B0(new_n3594_), .Y(new_n3595_));
  XOR2X1   g02593(.A(new_n3570_), .B(new_n3592_), .Y(new_n3596_));
  AOI21X1  g02594(.A0(new_n3595_), .A1(new_n3589_), .B0(new_n3596_), .Y(new_n3597_));
  AND2X1   g02595(.A(new_n3586_), .B(new_n3580_), .Y(new_n3598_));
  OR2X1    g02596(.A(new_n2590_), .B(new_n2584_), .Y(new_n3599_));
  XOR2X1   g02597(.A(new_n3599_), .B(new_n3581_), .Y(new_n3600_));
  OR4X1    g02598(.A(new_n3568_), .B(new_n3578_), .C(new_n3600_), .D(new_n3577_), .Y(new_n3601_));
  OAI22X1  g02599(.A0(new_n3596_), .A1(new_n3572_), .B0(new_n3584_), .B1(new_n3577_), .Y(new_n3602_));
  NOR2X1   g02600(.A(new_n3602_), .B(new_n3601_), .Y(new_n3603_));
  OAI21X1  g02601(.A0(new_n3603_), .A1(new_n3598_), .B0(new_n3597_), .Y(new_n3604_));
  INVX1    g02602(.A(new_n2614_), .Y(new_n3605_));
  NOR2X1   g02603(.A(new_n2652_), .B(new_n3605_), .Y(new_n3606_));
  NAND3X1  g02604(.A(new_n3606_), .B(new_n3604_), .C(new_n3588_), .Y(new_n3607_));
  AND2X1   g02605(.A(new_n3587_), .B(new_n3574_), .Y(new_n3608_));
  NAND2X1  g02606(.A(new_n3586_), .B(new_n3580_), .Y(new_n3609_));
  OR2X1    g02607(.A(new_n3602_), .B(new_n3601_), .Y(new_n3610_));
  AOI21X1  g02608(.A0(new_n3610_), .A1(new_n3609_), .B0(new_n3574_), .Y(new_n3611_));
  OR2X1    g02609(.A(new_n2652_), .B(new_n3605_), .Y(new_n3612_));
  OAI21X1  g02610(.A0(new_n3611_), .A1(new_n3608_), .B0(new_n3612_), .Y(new_n3613_));
  AOI21X1  g02611(.A0(new_n3613_), .A1(new_n3607_), .B0(new_n3565_), .Y(new_n3614_));
  INVX1    g02612(.A(new_n3544_), .Y(new_n3615_));
  AND2X1   g02613(.A(new_n3556_), .B(new_n3544_), .Y(new_n3616_));
  AOI21X1  g02614(.A0(new_n3564_), .A1(new_n3615_), .B0(new_n3616_), .Y(new_n3617_));
  NAND3X1  g02615(.A(new_n3612_), .B(new_n3604_), .C(new_n3588_), .Y(new_n3618_));
  OAI21X1  g02616(.A0(new_n3611_), .A1(new_n3608_), .B0(new_n3606_), .Y(new_n3619_));
  AOI21X1  g02617(.A0(new_n3619_), .A1(new_n3618_), .B0(new_n3617_), .Y(new_n3620_));
  XOR2X1   g02618(.A(new_n2729_), .B(new_n2690_), .Y(new_n3621_));
  NOR2X1   g02619(.A(new_n3621_), .B(new_n2653_), .Y(new_n3622_));
  INVX1    g02620(.A(new_n3622_), .Y(new_n3623_));
  NOR3X1   g02621(.A(new_n3623_), .B(new_n3620_), .C(new_n3614_), .Y(new_n3624_));
  NOR3X1   g02622(.A(new_n3612_), .B(new_n3611_), .C(new_n3608_), .Y(new_n3625_));
  AOI21X1  g02623(.A0(new_n3604_), .A1(new_n3588_), .B0(new_n3606_), .Y(new_n3626_));
  OAI21X1  g02624(.A0(new_n3626_), .A1(new_n3625_), .B0(new_n3617_), .Y(new_n3627_));
  NOR3X1   g02625(.A(new_n3606_), .B(new_n3611_), .C(new_n3608_), .Y(new_n3628_));
  AOI21X1  g02626(.A0(new_n3604_), .A1(new_n3588_), .B0(new_n3612_), .Y(new_n3629_));
  OAI21X1  g02627(.A0(new_n3629_), .A1(new_n3628_), .B0(new_n3565_), .Y(new_n3630_));
  AOI21X1  g02628(.A0(new_n3630_), .A1(new_n3627_), .B0(new_n3622_), .Y(new_n3631_));
  OAI21X1  g02629(.A0(new_n3631_), .A1(new_n3624_), .B0(new_n3535_), .Y(new_n3632_));
  OR2X1    g02630(.A(new_n3534_), .B(new_n3528_), .Y(new_n3633_));
  NOR3X1   g02631(.A(new_n3622_), .B(new_n3620_), .C(new_n3614_), .Y(new_n3634_));
  AOI21X1  g02632(.A0(new_n3630_), .A1(new_n3627_), .B0(new_n3623_), .Y(new_n3635_));
  OAI21X1  g02633(.A0(new_n3635_), .A1(new_n3634_), .B0(new_n3633_), .Y(new_n3636_));
  NOR2X1   g02634(.A(new_n2731_), .B(new_n2577_), .Y(new_n3637_));
  NAND3X1  g02635(.A(new_n3637_), .B(new_n3636_), .C(new_n3632_), .Y(new_n3638_));
  NAND3X1  g02636(.A(new_n3622_), .B(new_n3630_), .C(new_n3627_), .Y(new_n3639_));
  OAI21X1  g02637(.A0(new_n3620_), .A1(new_n3614_), .B0(new_n3623_), .Y(new_n3640_));
  AOI21X1  g02638(.A0(new_n3640_), .A1(new_n3639_), .B0(new_n3633_), .Y(new_n3641_));
  NAND3X1  g02639(.A(new_n3623_), .B(new_n3630_), .C(new_n3627_), .Y(new_n3642_));
  OAI21X1  g02640(.A0(new_n3620_), .A1(new_n3614_), .B0(new_n3622_), .Y(new_n3643_));
  AOI21X1  g02641(.A0(new_n3643_), .A1(new_n3642_), .B0(new_n3535_), .Y(new_n3644_));
  INVX1    g02642(.A(new_n3637_), .Y(new_n3645_));
  OAI21X1  g02643(.A0(new_n3644_), .A1(new_n3641_), .B0(new_n3645_), .Y(new_n3646_));
  AND2X1   g02644(.A(new_n3646_), .B(new_n3638_), .Y(new_n3647_));
  AND2X1   g02645(.A(new_n2560_), .B(new_n2558_), .Y(new_n3648_));
  OR2X1    g02646(.A(new_n2562_), .B(new_n3648_), .Y(new_n3649_));
  XOR2X1   g02647(.A(new_n2569_), .B(new_n3649_), .Y(new_n3650_));
  XOR2X1   g02648(.A(new_n2573_), .B(new_n2571_), .Y(new_n3651_));
  NOR2X1   g02649(.A(new_n2569_), .B(new_n2563_), .Y(new_n3652_));
  NOR2X1   g02650(.A(new_n2573_), .B(new_n2571_), .Y(new_n3653_));
  AOI21X1  g02651(.A0(new_n3652_), .A1(new_n3651_), .B0(new_n3653_), .Y(new_n3654_));
  XOR2X1   g02652(.A(new_n3652_), .B(new_n3651_), .Y(new_n3655_));
  OAI21X1  g02653(.A0(new_n3654_), .A1(new_n3650_), .B0(new_n3655_), .Y(new_n3656_));
  INVX1    g02654(.A(new_n3656_), .Y(new_n3657_));
  XOR2X1   g02655(.A(new_n2551_), .B(new_n2545_), .Y(new_n3658_));
  AOI21X1  g02656(.A0(new_n2541_), .A1(new_n2539_), .B0(new_n2544_), .Y(new_n3659_));
  NOR4X1   g02657(.A(new_n2555_), .B(new_n2553_), .C(new_n2551_), .D(new_n3659_), .Y(new_n3660_));
  NOR4X1   g02658(.A(new_n2573_), .B(new_n2571_), .C(new_n2569_), .D(new_n2563_), .Y(new_n3661_));
  OR4X1    g02659(.A(new_n3661_), .B(new_n3650_), .C(new_n3660_), .D(new_n3658_), .Y(new_n3662_));
  XOR2X1   g02660(.A(new_n2555_), .B(new_n2553_), .Y(new_n3663_));
  NOR2X1   g02661(.A(new_n2551_), .B(new_n3659_), .Y(new_n3664_));
  NOR2X1   g02662(.A(new_n2555_), .B(new_n2553_), .Y(new_n3665_));
  AOI21X1  g02663(.A0(new_n3664_), .A1(new_n3663_), .B0(new_n3665_), .Y(new_n3666_));
  XOR2X1   g02664(.A(new_n3664_), .B(new_n3663_), .Y(new_n3667_));
  OAI21X1  g02665(.A0(new_n3666_), .A1(new_n3658_), .B0(new_n3667_), .Y(new_n3668_));
  XOR2X1   g02666(.A(new_n3668_), .B(new_n3662_), .Y(new_n3669_));
  AND2X1   g02667(.A(new_n3669_), .B(new_n3656_), .Y(new_n3670_));
  AND2X1   g02668(.A(new_n3668_), .B(new_n3662_), .Y(new_n3671_));
  OR2X1    g02669(.A(new_n2551_), .B(new_n3659_), .Y(new_n3672_));
  XOR2X1   g02670(.A(new_n3672_), .B(new_n3663_), .Y(new_n3673_));
  OR4X1    g02671(.A(new_n3650_), .B(new_n3660_), .C(new_n3673_), .D(new_n3658_), .Y(new_n3674_));
  OR4X1    g02672(.A(new_n2573_), .B(new_n2571_), .C(new_n2569_), .D(new_n2563_), .Y(new_n3675_));
  OAI21X1  g02673(.A0(new_n3666_), .A1(new_n3658_), .B0(new_n3675_), .Y(new_n3676_));
  NOR2X1   g02674(.A(new_n3676_), .B(new_n3674_), .Y(new_n3677_));
  OR2X1    g02675(.A(new_n3677_), .B(new_n3671_), .Y(new_n3678_));
  AOI21X1  g02676(.A0(new_n3678_), .A1(new_n3657_), .B0(new_n3670_), .Y(new_n3679_));
  AND2X1   g02677(.A(new_n2521_), .B(new_n2519_), .Y(new_n3680_));
  OR2X1    g02678(.A(new_n2523_), .B(new_n3680_), .Y(new_n3681_));
  XOR2X1   g02679(.A(new_n2530_), .B(new_n3681_), .Y(new_n3682_));
  XOR2X1   g02680(.A(new_n2534_), .B(new_n2532_), .Y(new_n3683_));
  NOR2X1   g02681(.A(new_n2530_), .B(new_n2524_), .Y(new_n3684_));
  NOR2X1   g02682(.A(new_n2534_), .B(new_n2532_), .Y(new_n3685_));
  AOI21X1  g02683(.A0(new_n3684_), .A1(new_n3683_), .B0(new_n3685_), .Y(new_n3686_));
  XOR2X1   g02684(.A(new_n3684_), .B(new_n3683_), .Y(new_n3687_));
  OAI21X1  g02685(.A0(new_n3686_), .A1(new_n3682_), .B0(new_n3687_), .Y(new_n3688_));
  AND2X1   g02686(.A(new_n2503_), .B(new_n2501_), .Y(new_n3689_));
  OR2X1    g02687(.A(new_n2505_), .B(new_n3689_), .Y(new_n3690_));
  XOR2X1   g02688(.A(new_n2512_), .B(new_n3690_), .Y(new_n3691_));
  NOR4X1   g02689(.A(new_n2516_), .B(new_n2514_), .C(new_n2512_), .D(new_n2506_), .Y(new_n3692_));
  NOR4X1   g02690(.A(new_n2534_), .B(new_n2532_), .C(new_n2530_), .D(new_n2524_), .Y(new_n3693_));
  OR4X1    g02691(.A(new_n3693_), .B(new_n3682_), .C(new_n3692_), .D(new_n3691_), .Y(new_n3694_));
  XOR2X1   g02692(.A(new_n2516_), .B(new_n2514_), .Y(new_n3695_));
  NOR2X1   g02693(.A(new_n2512_), .B(new_n2506_), .Y(new_n3696_));
  NOR2X1   g02694(.A(new_n2516_), .B(new_n2514_), .Y(new_n3697_));
  AOI21X1  g02695(.A0(new_n3696_), .A1(new_n3695_), .B0(new_n3697_), .Y(new_n3698_));
  XOR2X1   g02696(.A(new_n3696_), .B(new_n3695_), .Y(new_n3699_));
  OAI21X1  g02697(.A0(new_n3698_), .A1(new_n3691_), .B0(new_n3699_), .Y(new_n3700_));
  XOR2X1   g02698(.A(new_n3700_), .B(new_n3694_), .Y(new_n3701_));
  AND2X1   g02699(.A(new_n3701_), .B(new_n3688_), .Y(new_n3702_));
  NAND2X1  g02700(.A(new_n3700_), .B(new_n3694_), .Y(new_n3703_));
  OR2X1    g02701(.A(new_n2512_), .B(new_n2506_), .Y(new_n3704_));
  XOR2X1   g02702(.A(new_n3704_), .B(new_n3695_), .Y(new_n3705_));
  OR4X1    g02703(.A(new_n3682_), .B(new_n3692_), .C(new_n3705_), .D(new_n3691_), .Y(new_n3706_));
  AND2X1   g02704(.A(new_n2529_), .B(\A[504] ), .Y(new_n3707_));
  OR2X1    g02705(.A(new_n3707_), .B(new_n2531_), .Y(new_n3708_));
  XOR2X1   g02706(.A(new_n2534_), .B(new_n3708_), .Y(new_n3709_));
  XOR2X1   g02707(.A(new_n3684_), .B(new_n3709_), .Y(new_n3710_));
  OAI22X1  g02708(.A0(new_n3710_), .A1(new_n3686_), .B0(new_n3698_), .B1(new_n3691_), .Y(new_n3711_));
  OR2X1    g02709(.A(new_n3711_), .B(new_n3706_), .Y(new_n3712_));
  AOI21X1  g02710(.A0(new_n3712_), .A1(new_n3703_), .B0(new_n3688_), .Y(new_n3713_));
  OR2X1    g02711(.A(new_n2575_), .B(new_n2537_), .Y(new_n3714_));
  NOR3X1   g02712(.A(new_n3714_), .B(new_n3713_), .C(new_n3702_), .Y(new_n3715_));
  NAND2X1  g02713(.A(new_n3701_), .B(new_n3688_), .Y(new_n3716_));
  XOR2X1   g02714(.A(new_n2530_), .B(new_n2524_), .Y(new_n3717_));
  OR2X1    g02715(.A(new_n2530_), .B(new_n2524_), .Y(new_n3718_));
  OR2X1    g02716(.A(new_n2534_), .B(new_n2532_), .Y(new_n3719_));
  OAI21X1  g02717(.A0(new_n3718_), .A1(new_n3709_), .B0(new_n3719_), .Y(new_n3720_));
  AOI21X1  g02718(.A0(new_n3720_), .A1(new_n3717_), .B0(new_n3710_), .Y(new_n3721_));
  AND2X1   g02719(.A(new_n3700_), .B(new_n3694_), .Y(new_n3722_));
  NOR2X1   g02720(.A(new_n3711_), .B(new_n3706_), .Y(new_n3723_));
  OAI21X1  g02721(.A0(new_n3723_), .A1(new_n3722_), .B0(new_n3721_), .Y(new_n3724_));
  NOR2X1   g02722(.A(new_n2575_), .B(new_n2537_), .Y(new_n3725_));
  AOI21X1  g02723(.A0(new_n3724_), .A1(new_n3716_), .B0(new_n3725_), .Y(new_n3726_));
  OAI21X1  g02724(.A0(new_n3726_), .A1(new_n3715_), .B0(new_n3679_), .Y(new_n3727_));
  MX2X1    g02725(.A(new_n3678_), .B(new_n3669_), .S0(new_n3656_), .Y(new_n3728_));
  NOR3X1   g02726(.A(new_n3725_), .B(new_n3713_), .C(new_n3702_), .Y(new_n3729_));
  AOI21X1  g02727(.A0(new_n3724_), .A1(new_n3716_), .B0(new_n3714_), .Y(new_n3730_));
  OAI21X1  g02728(.A0(new_n3730_), .A1(new_n3729_), .B0(new_n3728_), .Y(new_n3731_));
  XOR2X1   g02729(.A(new_n2575_), .B(new_n2536_), .Y(new_n3732_));
  NOR2X1   g02730(.A(new_n3732_), .B(new_n2499_), .Y(new_n3733_));
  NAND3X1  g02731(.A(new_n3733_), .B(new_n3731_), .C(new_n3727_), .Y(new_n3734_));
  NAND3X1  g02732(.A(new_n3725_), .B(new_n3724_), .C(new_n3716_), .Y(new_n3735_));
  OAI21X1  g02733(.A0(new_n3713_), .A1(new_n3702_), .B0(new_n3714_), .Y(new_n3736_));
  AOI21X1  g02734(.A0(new_n3736_), .A1(new_n3735_), .B0(new_n3728_), .Y(new_n3737_));
  NAND3X1  g02735(.A(new_n3714_), .B(new_n3724_), .C(new_n3716_), .Y(new_n3738_));
  OAI21X1  g02736(.A0(new_n3713_), .A1(new_n3702_), .B0(new_n3725_), .Y(new_n3739_));
  AOI21X1  g02737(.A0(new_n3739_), .A1(new_n3738_), .B0(new_n3679_), .Y(new_n3740_));
  INVX1    g02738(.A(new_n3733_), .Y(new_n3741_));
  OAI21X1  g02739(.A0(new_n3740_), .A1(new_n3737_), .B0(new_n3741_), .Y(new_n3742_));
  AND2X1   g02740(.A(new_n3742_), .B(new_n3734_), .Y(new_n3743_));
  AND2X1   g02741(.A(new_n2483_), .B(new_n2481_), .Y(new_n3744_));
  OR2X1    g02742(.A(new_n2485_), .B(new_n3744_), .Y(new_n3745_));
  XOR2X1   g02743(.A(new_n2492_), .B(new_n3745_), .Y(new_n3746_));
  XOR2X1   g02744(.A(new_n2496_), .B(new_n2494_), .Y(new_n3747_));
  NOR2X1   g02745(.A(new_n2492_), .B(new_n2486_), .Y(new_n3748_));
  NOR2X1   g02746(.A(new_n2496_), .B(new_n2494_), .Y(new_n3749_));
  AOI21X1  g02747(.A0(new_n3748_), .A1(new_n3747_), .B0(new_n3749_), .Y(new_n3750_));
  XOR2X1   g02748(.A(new_n3748_), .B(new_n3747_), .Y(new_n3751_));
  OAI21X1  g02749(.A0(new_n3750_), .A1(new_n3746_), .B0(new_n3751_), .Y(new_n3752_));
  XOR2X1   g02750(.A(new_n2474_), .B(new_n2468_), .Y(new_n3753_));
  AOI21X1  g02751(.A0(new_n2464_), .A1(new_n2462_), .B0(new_n2467_), .Y(new_n3754_));
  NOR4X1   g02752(.A(new_n2478_), .B(new_n2476_), .C(new_n2474_), .D(new_n3754_), .Y(new_n3755_));
  NOR4X1   g02753(.A(new_n2496_), .B(new_n2494_), .C(new_n2492_), .D(new_n2486_), .Y(new_n3756_));
  OR4X1    g02754(.A(new_n3756_), .B(new_n3746_), .C(new_n3755_), .D(new_n3753_), .Y(new_n3757_));
  XOR2X1   g02755(.A(new_n2478_), .B(new_n2476_), .Y(new_n3758_));
  NOR2X1   g02756(.A(new_n2474_), .B(new_n3754_), .Y(new_n3759_));
  NOR2X1   g02757(.A(new_n2478_), .B(new_n2476_), .Y(new_n3760_));
  AOI21X1  g02758(.A0(new_n3759_), .A1(new_n3758_), .B0(new_n3760_), .Y(new_n3761_));
  XOR2X1   g02759(.A(new_n3759_), .B(new_n3758_), .Y(new_n3762_));
  OAI21X1  g02760(.A0(new_n3761_), .A1(new_n3753_), .B0(new_n3762_), .Y(new_n3763_));
  XOR2X1   g02761(.A(new_n3763_), .B(new_n3757_), .Y(new_n3764_));
  NAND2X1  g02762(.A(new_n3764_), .B(new_n3752_), .Y(new_n3765_));
  XOR2X1   g02763(.A(new_n2492_), .B(new_n2486_), .Y(new_n3766_));
  AND2X1   g02764(.A(new_n3748_), .B(new_n3747_), .Y(new_n3767_));
  OR2X1    g02765(.A(new_n3749_), .B(new_n3767_), .Y(new_n3768_));
  OR2X1    g02766(.A(new_n2492_), .B(new_n2486_), .Y(new_n3769_));
  XOR2X1   g02767(.A(new_n3769_), .B(new_n3747_), .Y(new_n3770_));
  AOI21X1  g02768(.A0(new_n3768_), .A1(new_n3766_), .B0(new_n3770_), .Y(new_n3771_));
  AND2X1   g02769(.A(new_n3763_), .B(new_n3757_), .Y(new_n3772_));
  OR2X1    g02770(.A(new_n2474_), .B(new_n3754_), .Y(new_n3773_));
  XOR2X1   g02771(.A(new_n3773_), .B(new_n3758_), .Y(new_n3774_));
  OR4X1    g02772(.A(new_n3746_), .B(new_n3755_), .C(new_n3774_), .D(new_n3753_), .Y(new_n3775_));
  OAI22X1  g02773(.A0(new_n3770_), .A1(new_n3750_), .B0(new_n3761_), .B1(new_n3753_), .Y(new_n3776_));
  NOR2X1   g02774(.A(new_n3776_), .B(new_n3775_), .Y(new_n3777_));
  OAI21X1  g02775(.A0(new_n3777_), .A1(new_n3772_), .B0(new_n3771_), .Y(new_n3778_));
  INVX1    g02776(.A(new_n2460_), .Y(new_n3779_));
  NOR2X1   g02777(.A(new_n2498_), .B(new_n3779_), .Y(new_n3780_));
  NAND3X1  g02778(.A(new_n3780_), .B(new_n3778_), .C(new_n3765_), .Y(new_n3781_));
  AND2X1   g02779(.A(new_n3764_), .B(new_n3752_), .Y(new_n3782_));
  NAND2X1  g02780(.A(new_n3763_), .B(new_n3757_), .Y(new_n3783_));
  OR2X1    g02781(.A(new_n3776_), .B(new_n3775_), .Y(new_n3784_));
  AOI21X1  g02782(.A0(new_n3784_), .A1(new_n3783_), .B0(new_n3752_), .Y(new_n3785_));
  OR2X1    g02783(.A(new_n2498_), .B(new_n3779_), .Y(new_n3786_));
  OAI21X1  g02784(.A0(new_n3785_), .A1(new_n3782_), .B0(new_n3786_), .Y(new_n3787_));
  OR2X1    g02785(.A(new_n2454_), .B(new_n2448_), .Y(new_n3788_));
  AND2X1   g02786(.A(new_n2446_), .B(\A[468] ), .Y(new_n3789_));
  OR2X1    g02787(.A(new_n3789_), .B(new_n2455_), .Y(new_n3790_));
  XOR2X1   g02788(.A(new_n2458_), .B(new_n3790_), .Y(new_n3791_));
  XOR2X1   g02789(.A(new_n3791_), .B(new_n3788_), .Y(new_n3792_));
  XOR2X1   g02790(.A(new_n2454_), .B(new_n2448_), .Y(new_n3793_));
  OR2X1    g02791(.A(new_n2458_), .B(new_n2456_), .Y(new_n3794_));
  OAI21X1  g02792(.A0(new_n3791_), .A1(new_n3788_), .B0(new_n3794_), .Y(new_n3795_));
  NAND2X1  g02793(.A(new_n3795_), .B(new_n3793_), .Y(new_n3796_));
  NAND2X1  g02794(.A(new_n3796_), .B(new_n3792_), .Y(new_n3797_));
  AND2X1   g02795(.A(new_n2427_), .B(new_n2425_), .Y(new_n3798_));
  OR2X1    g02796(.A(new_n2429_), .B(new_n3798_), .Y(new_n3799_));
  XOR2X1   g02797(.A(new_n2436_), .B(new_n3799_), .Y(new_n3800_));
  NOR4X1   g02798(.A(new_n2440_), .B(new_n2438_), .C(new_n2436_), .D(new_n2430_), .Y(new_n3801_));
  AND2X1   g02799(.A(new_n2445_), .B(new_n2443_), .Y(new_n3802_));
  OR2X1    g02800(.A(new_n2447_), .B(new_n3802_), .Y(new_n3803_));
  XOR2X1   g02801(.A(new_n2454_), .B(new_n3803_), .Y(new_n3804_));
  NOR4X1   g02802(.A(new_n2458_), .B(new_n2456_), .C(new_n2454_), .D(new_n2448_), .Y(new_n3805_));
  OR4X1    g02803(.A(new_n3805_), .B(new_n3804_), .C(new_n3801_), .D(new_n3800_), .Y(new_n3806_));
  XOR2X1   g02804(.A(new_n2440_), .B(new_n2438_), .Y(new_n3807_));
  NOR2X1   g02805(.A(new_n2436_), .B(new_n2430_), .Y(new_n3808_));
  NOR2X1   g02806(.A(new_n2440_), .B(new_n2438_), .Y(new_n3809_));
  AOI21X1  g02807(.A0(new_n3808_), .A1(new_n3807_), .B0(new_n3809_), .Y(new_n3810_));
  XOR2X1   g02808(.A(new_n3808_), .B(new_n3807_), .Y(new_n3811_));
  OAI21X1  g02809(.A0(new_n3810_), .A1(new_n3800_), .B0(new_n3811_), .Y(new_n3812_));
  XOR2X1   g02810(.A(new_n3812_), .B(new_n3806_), .Y(new_n3813_));
  NOR4X1   g02811(.A(new_n3805_), .B(new_n3804_), .C(new_n3801_), .D(new_n3800_), .Y(new_n3814_));
  OR2X1    g02812(.A(new_n2436_), .B(new_n2430_), .Y(new_n3815_));
  XOR2X1   g02813(.A(new_n3815_), .B(new_n3807_), .Y(new_n3816_));
  NOR2X1   g02814(.A(new_n3810_), .B(new_n3800_), .Y(new_n3817_));
  NOR2X1   g02815(.A(new_n3817_), .B(new_n3816_), .Y(new_n3818_));
  OR4X1    g02816(.A(new_n3804_), .B(new_n3801_), .C(new_n3816_), .D(new_n3800_), .Y(new_n3819_));
  OR2X1    g02817(.A(new_n3817_), .B(new_n3805_), .Y(new_n3820_));
  OAI22X1  g02818(.A0(new_n3820_), .A1(new_n3819_), .B0(new_n3818_), .B1(new_n3814_), .Y(new_n3821_));
  MX2X1    g02819(.A(new_n3821_), .B(new_n3813_), .S0(new_n3797_), .Y(new_n3822_));
  AOI21X1  g02820(.A0(new_n3787_), .A1(new_n3781_), .B0(new_n3822_), .Y(new_n3823_));
  AND2X1   g02821(.A(new_n3796_), .B(new_n3792_), .Y(new_n3824_));
  AND2X1   g02822(.A(new_n3813_), .B(new_n3797_), .Y(new_n3825_));
  AOI21X1  g02823(.A0(new_n3821_), .A1(new_n3824_), .B0(new_n3825_), .Y(new_n3826_));
  NAND3X1  g02824(.A(new_n3786_), .B(new_n3778_), .C(new_n3765_), .Y(new_n3827_));
  OAI21X1  g02825(.A0(new_n3785_), .A1(new_n3782_), .B0(new_n3780_), .Y(new_n3828_));
  AOI21X1  g02826(.A0(new_n3828_), .A1(new_n3827_), .B0(new_n3826_), .Y(new_n3829_));
  NOR2X1   g02827(.A(new_n3829_), .B(new_n3823_), .Y(new_n3830_));
  NAND3X1  g02828(.A(new_n3741_), .B(new_n3731_), .C(new_n3727_), .Y(new_n3831_));
  OAI21X1  g02829(.A0(new_n3740_), .A1(new_n3737_), .B0(new_n3733_), .Y(new_n3832_));
  AND2X1   g02830(.A(new_n3832_), .B(new_n3831_), .Y(new_n3833_));
  MX2X1    g02831(.A(new_n3833_), .B(new_n3743_), .S0(new_n3830_), .Y(new_n3834_));
  NAND3X1  g02832(.A(new_n3645_), .B(new_n3636_), .C(new_n3632_), .Y(new_n3835_));
  OAI21X1  g02833(.A0(new_n3644_), .A1(new_n3641_), .B0(new_n3637_), .Y(new_n3836_));
  AND2X1   g02834(.A(new_n3836_), .B(new_n3835_), .Y(new_n3837_));
  MX2X1    g02835(.A(new_n3837_), .B(new_n3647_), .S0(new_n3834_), .Y(new_n3838_));
  NAND3X1  g02836(.A(new_n3448_), .B(new_n3438_), .C(new_n3430_), .Y(new_n3839_));
  OAI21X1  g02837(.A0(new_n3447_), .A1(new_n3444_), .B0(new_n3440_), .Y(new_n3840_));
  AND2X1   g02838(.A(new_n3840_), .B(new_n3839_), .Y(new_n3841_));
  MX2X1    g02839(.A(new_n3841_), .B(new_n3450_), .S0(new_n3838_), .Y(new_n3842_));
  INVX1    g02840(.A(new_n3041_), .Y(new_n3843_));
  AND2X1   g02841(.A(new_n3042_), .B(new_n3843_), .Y(new_n3844_));
  OR2X1    g02842(.A(new_n3844_), .B(new_n2423_), .Y(new_n3845_));
  OAI21X1  g02843(.A0(new_n2423_), .A1(new_n2411_), .B0(new_n3844_), .Y(new_n3846_));
  OAI21X1  g02844(.A0(new_n3845_), .A1(new_n2411_), .B0(new_n3846_), .Y(new_n3847_));
  MX2X1    g02845(.A(new_n3847_), .B(new_n3046_), .S0(new_n3842_), .Y(new_n3848_));
  INVX1    g02846(.A(new_n3848_), .Y(new_n3849_));
  INVX1    g02847(.A(\A[968] ), .Y(new_n3850_));
  OR2X1    g02848(.A(new_n3850_), .B(\A[967] ), .Y(new_n3851_));
  INVX1    g02849(.A(\A[969] ), .Y(new_n3852_));
  AOI21X1  g02850(.A0(new_n3850_), .A1(\A[967] ), .B0(new_n3852_), .Y(new_n3853_));
  XOR2X1   g02851(.A(\A[968] ), .B(\A[967] ), .Y(new_n3854_));
  AND2X1   g02852(.A(new_n3854_), .B(new_n3852_), .Y(new_n3855_));
  AOI21X1  g02853(.A0(new_n3853_), .A1(new_n3851_), .B0(new_n3855_), .Y(new_n3856_));
  INVX1    g02854(.A(\A[972] ), .Y(new_n3857_));
  INVX1    g02855(.A(\A[971] ), .Y(new_n3858_));
  OR2X1    g02856(.A(new_n3858_), .B(\A[970] ), .Y(new_n3859_));
  AOI21X1  g02857(.A0(new_n3858_), .A1(\A[970] ), .B0(new_n3857_), .Y(new_n3860_));
  XOR2X1   g02858(.A(\A[971] ), .B(\A[970] ), .Y(new_n3861_));
  AOI22X1  g02859(.A0(new_n3861_), .A1(new_n3857_), .B0(new_n3860_), .B1(new_n3859_), .Y(new_n3862_));
  NOR2X1   g02860(.A(new_n3862_), .B(new_n3856_), .Y(new_n3863_));
  AND2X1   g02861(.A(\A[971] ), .B(\A[970] ), .Y(new_n3864_));
  AND2X1   g02862(.A(new_n3861_), .B(\A[972] ), .Y(new_n3865_));
  OR2X1    g02863(.A(new_n3865_), .B(new_n3864_), .Y(new_n3866_));
  AND2X1   g02864(.A(\A[968] ), .B(\A[967] ), .Y(new_n3867_));
  AOI21X1  g02865(.A0(new_n3854_), .A1(\A[969] ), .B0(new_n3867_), .Y(new_n3868_));
  XOR2X1   g02866(.A(new_n3868_), .B(new_n3866_), .Y(new_n3869_));
  XOR2X1   g02867(.A(new_n3869_), .B(new_n3863_), .Y(new_n3870_));
  XOR2X1   g02868(.A(new_n3862_), .B(new_n3856_), .Y(new_n3871_));
  OR2X1    g02869(.A(new_n3862_), .B(new_n3856_), .Y(new_n3872_));
  AOI21X1  g02870(.A0(new_n3861_), .A1(\A[972] ), .B0(new_n3864_), .Y(new_n3873_));
  OR2X1    g02871(.A(new_n3868_), .B(new_n3873_), .Y(new_n3874_));
  OAI21X1  g02872(.A0(new_n3869_), .A1(new_n3872_), .B0(new_n3874_), .Y(new_n3875_));
  AND2X1   g02873(.A(new_n3875_), .B(new_n3871_), .Y(new_n3876_));
  OR2X1    g02874(.A(new_n3876_), .B(new_n3870_), .Y(new_n3877_));
  AND2X1   g02875(.A(\A[977] ), .B(\A[976] ), .Y(new_n3878_));
  XOR2X1   g02876(.A(\A[977] ), .B(\A[976] ), .Y(new_n3879_));
  AOI21X1  g02877(.A0(new_n3879_), .A1(\A[978] ), .B0(new_n3878_), .Y(new_n3880_));
  AND2X1   g02878(.A(\A[974] ), .B(\A[973] ), .Y(new_n3881_));
  XOR2X1   g02879(.A(\A[974] ), .B(\A[973] ), .Y(new_n3882_));
  AOI21X1  g02880(.A0(new_n3882_), .A1(\A[975] ), .B0(new_n3881_), .Y(new_n3883_));
  INVX1    g02881(.A(\A[974] ), .Y(new_n3884_));
  OR2X1    g02882(.A(new_n3884_), .B(\A[973] ), .Y(new_n3885_));
  INVX1    g02883(.A(\A[975] ), .Y(new_n3886_));
  AOI21X1  g02884(.A0(new_n3884_), .A1(\A[973] ), .B0(new_n3886_), .Y(new_n3887_));
  AND2X1   g02885(.A(new_n3882_), .B(new_n3886_), .Y(new_n3888_));
  AOI21X1  g02886(.A0(new_n3887_), .A1(new_n3885_), .B0(new_n3888_), .Y(new_n3889_));
  INVX1    g02887(.A(\A[978] ), .Y(new_n3890_));
  INVX1    g02888(.A(\A[977] ), .Y(new_n3891_));
  OR2X1    g02889(.A(new_n3891_), .B(\A[976] ), .Y(new_n3892_));
  AOI21X1  g02890(.A0(new_n3891_), .A1(\A[976] ), .B0(new_n3890_), .Y(new_n3893_));
  AOI22X1  g02891(.A0(new_n3893_), .A1(new_n3892_), .B0(new_n3879_), .B1(new_n3890_), .Y(new_n3894_));
  OR4X1    g02892(.A(new_n3894_), .B(new_n3889_), .C(new_n3883_), .D(new_n3880_), .Y(new_n3895_));
  OR4X1    g02893(.A(new_n3868_), .B(new_n3873_), .C(new_n3862_), .D(new_n3856_), .Y(new_n3896_));
  XOR2X1   g02894(.A(new_n3894_), .B(new_n3889_), .Y(new_n3897_));
  NAND4X1  g02895(.A(new_n3897_), .B(new_n3896_), .C(new_n3895_), .D(new_n3871_), .Y(new_n3898_));
  XOR2X1   g02896(.A(new_n3883_), .B(new_n3880_), .Y(new_n3899_));
  NOR2X1   g02897(.A(new_n3894_), .B(new_n3889_), .Y(new_n3900_));
  NOR2X1   g02898(.A(new_n3883_), .B(new_n3880_), .Y(new_n3901_));
  AOI21X1  g02899(.A0(new_n3900_), .A1(new_n3899_), .B0(new_n3901_), .Y(new_n3902_));
  XOR2X1   g02900(.A(new_n3900_), .B(new_n3899_), .Y(new_n3903_));
  AND2X1   g02901(.A(new_n3887_), .B(new_n3885_), .Y(new_n3904_));
  OR2X1    g02902(.A(new_n3888_), .B(new_n3904_), .Y(new_n3905_));
  XOR2X1   g02903(.A(new_n3894_), .B(new_n3905_), .Y(new_n3906_));
  OAI21X1  g02904(.A0(new_n3906_), .A1(new_n3902_), .B0(new_n3903_), .Y(new_n3907_));
  XOR2X1   g02905(.A(new_n3907_), .B(new_n3898_), .Y(new_n3908_));
  INVX1    g02906(.A(new_n3898_), .Y(new_n3909_));
  OR2X1    g02907(.A(new_n3894_), .B(new_n3889_), .Y(new_n3910_));
  XOR2X1   g02908(.A(new_n3910_), .B(new_n3899_), .Y(new_n3911_));
  NOR2X1   g02909(.A(new_n3906_), .B(new_n3902_), .Y(new_n3912_));
  NOR2X1   g02910(.A(new_n3912_), .B(new_n3911_), .Y(new_n3913_));
  NOR4X1   g02911(.A(new_n3868_), .B(new_n3873_), .C(new_n3862_), .D(new_n3856_), .Y(new_n3914_));
  NAND2X1  g02912(.A(new_n3897_), .B(new_n3871_), .Y(new_n3915_));
  AOI21X1  g02913(.A0(new_n3906_), .A1(new_n3911_), .B0(new_n3902_), .Y(new_n3916_));
  OR4X1    g02914(.A(new_n3916_), .B(new_n3915_), .C(new_n3914_), .D(new_n3911_), .Y(new_n3917_));
  OAI21X1  g02915(.A0(new_n3913_), .A1(new_n3909_), .B0(new_n3917_), .Y(new_n3918_));
  MX2X1    g02916(.A(new_n3918_), .B(new_n3908_), .S0(new_n3877_), .Y(new_n3919_));
  INVX1    g02917(.A(\A[980] ), .Y(new_n3920_));
  OR2X1    g02918(.A(new_n3920_), .B(\A[979] ), .Y(new_n3921_));
  INVX1    g02919(.A(\A[981] ), .Y(new_n3922_));
  AOI21X1  g02920(.A0(new_n3920_), .A1(\A[979] ), .B0(new_n3922_), .Y(new_n3923_));
  XOR2X1   g02921(.A(\A[980] ), .B(\A[979] ), .Y(new_n3924_));
  AND2X1   g02922(.A(new_n3924_), .B(new_n3922_), .Y(new_n3925_));
  AOI21X1  g02923(.A0(new_n3923_), .A1(new_n3921_), .B0(new_n3925_), .Y(new_n3926_));
  INVX1    g02924(.A(\A[984] ), .Y(new_n3927_));
  INVX1    g02925(.A(\A[983] ), .Y(new_n3928_));
  OR2X1    g02926(.A(new_n3928_), .B(\A[982] ), .Y(new_n3929_));
  AOI21X1  g02927(.A0(new_n3928_), .A1(\A[982] ), .B0(new_n3927_), .Y(new_n3930_));
  XOR2X1   g02928(.A(\A[983] ), .B(\A[982] ), .Y(new_n3931_));
  AOI22X1  g02929(.A0(new_n3931_), .A1(new_n3927_), .B0(new_n3930_), .B1(new_n3929_), .Y(new_n3932_));
  NOR2X1   g02930(.A(new_n3932_), .B(new_n3926_), .Y(new_n3933_));
  AND2X1   g02931(.A(\A[983] ), .B(\A[982] ), .Y(new_n3934_));
  AND2X1   g02932(.A(new_n3931_), .B(\A[984] ), .Y(new_n3935_));
  OR2X1    g02933(.A(new_n3935_), .B(new_n3934_), .Y(new_n3936_));
  AND2X1   g02934(.A(\A[980] ), .B(\A[979] ), .Y(new_n3937_));
  AOI21X1  g02935(.A0(new_n3924_), .A1(\A[981] ), .B0(new_n3937_), .Y(new_n3938_));
  XOR2X1   g02936(.A(new_n3938_), .B(new_n3936_), .Y(new_n3939_));
  XOR2X1   g02937(.A(new_n3939_), .B(new_n3933_), .Y(new_n3940_));
  XOR2X1   g02938(.A(new_n3932_), .B(new_n3926_), .Y(new_n3941_));
  OR2X1    g02939(.A(new_n3932_), .B(new_n3926_), .Y(new_n3942_));
  AOI21X1  g02940(.A0(new_n3931_), .A1(\A[984] ), .B0(new_n3934_), .Y(new_n3943_));
  OR2X1    g02941(.A(new_n3938_), .B(new_n3943_), .Y(new_n3944_));
  OAI21X1  g02942(.A0(new_n3939_), .A1(new_n3942_), .B0(new_n3944_), .Y(new_n3945_));
  AND2X1   g02943(.A(new_n3945_), .B(new_n3941_), .Y(new_n3946_));
  OR2X1    g02944(.A(new_n3946_), .B(new_n3940_), .Y(new_n3947_));
  AND2X1   g02945(.A(new_n3923_), .B(new_n3921_), .Y(new_n3948_));
  OR2X1    g02946(.A(new_n3925_), .B(new_n3948_), .Y(new_n3949_));
  XOR2X1   g02947(.A(new_n3932_), .B(new_n3949_), .Y(new_n3950_));
  AND2X1   g02948(.A(\A[989] ), .B(\A[988] ), .Y(new_n3951_));
  XOR2X1   g02949(.A(\A[989] ), .B(\A[988] ), .Y(new_n3952_));
  AOI21X1  g02950(.A0(new_n3952_), .A1(\A[990] ), .B0(new_n3951_), .Y(new_n3953_));
  AND2X1   g02951(.A(\A[986] ), .B(\A[985] ), .Y(new_n3954_));
  XOR2X1   g02952(.A(\A[986] ), .B(\A[985] ), .Y(new_n3955_));
  AOI21X1  g02953(.A0(new_n3955_), .A1(\A[987] ), .B0(new_n3954_), .Y(new_n3956_));
  INVX1    g02954(.A(\A[986] ), .Y(new_n3957_));
  OR2X1    g02955(.A(new_n3957_), .B(\A[985] ), .Y(new_n3958_));
  INVX1    g02956(.A(\A[987] ), .Y(new_n3959_));
  AOI21X1  g02957(.A0(new_n3957_), .A1(\A[985] ), .B0(new_n3959_), .Y(new_n3960_));
  AND2X1   g02958(.A(new_n3955_), .B(new_n3959_), .Y(new_n3961_));
  AOI21X1  g02959(.A0(new_n3960_), .A1(new_n3958_), .B0(new_n3961_), .Y(new_n3962_));
  INVX1    g02960(.A(\A[990] ), .Y(new_n3963_));
  INVX1    g02961(.A(\A[989] ), .Y(new_n3964_));
  OR2X1    g02962(.A(new_n3964_), .B(\A[988] ), .Y(new_n3965_));
  AOI21X1  g02963(.A0(new_n3964_), .A1(\A[988] ), .B0(new_n3963_), .Y(new_n3966_));
  AOI22X1  g02964(.A0(new_n3966_), .A1(new_n3965_), .B0(new_n3952_), .B1(new_n3963_), .Y(new_n3967_));
  NOR4X1   g02965(.A(new_n3967_), .B(new_n3962_), .C(new_n3956_), .D(new_n3953_), .Y(new_n3968_));
  NOR4X1   g02966(.A(new_n3938_), .B(new_n3943_), .C(new_n3932_), .D(new_n3926_), .Y(new_n3969_));
  AND2X1   g02967(.A(new_n3960_), .B(new_n3958_), .Y(new_n3970_));
  OR2X1    g02968(.A(new_n3961_), .B(new_n3970_), .Y(new_n3971_));
  XOR2X1   g02969(.A(new_n3967_), .B(new_n3971_), .Y(new_n3972_));
  OR4X1    g02970(.A(new_n3972_), .B(new_n3969_), .C(new_n3968_), .D(new_n3950_), .Y(new_n3973_));
  XOR2X1   g02971(.A(new_n3956_), .B(new_n3953_), .Y(new_n3974_));
  NOR2X1   g02972(.A(new_n3967_), .B(new_n3962_), .Y(new_n3975_));
  NOR2X1   g02973(.A(new_n3956_), .B(new_n3953_), .Y(new_n3976_));
  AOI21X1  g02974(.A0(new_n3975_), .A1(new_n3974_), .B0(new_n3976_), .Y(new_n3977_));
  XOR2X1   g02975(.A(new_n3975_), .B(new_n3974_), .Y(new_n3978_));
  OAI21X1  g02976(.A0(new_n3972_), .A1(new_n3977_), .B0(new_n3978_), .Y(new_n3979_));
  XOR2X1   g02977(.A(new_n3979_), .B(new_n3973_), .Y(new_n3980_));
  NAND2X1  g02978(.A(new_n3980_), .B(new_n3947_), .Y(new_n3981_));
  OR2X1    g02979(.A(new_n3967_), .B(new_n3962_), .Y(new_n3982_));
  XOR2X1   g02980(.A(new_n3982_), .B(new_n3974_), .Y(new_n3983_));
  NOR4X1   g02981(.A(new_n3972_), .B(new_n3969_), .C(new_n3983_), .D(new_n3950_), .Y(new_n3984_));
  AND2X1   g02982(.A(new_n3975_), .B(new_n3974_), .Y(new_n3985_));
  XOR2X1   g02983(.A(new_n3967_), .B(new_n3962_), .Y(new_n3986_));
  OAI22X1  g02984(.A0(new_n3986_), .A1(new_n3978_), .B0(new_n3976_), .B1(new_n3985_), .Y(new_n3987_));
  AOI22X1  g02985(.A0(new_n3987_), .A1(new_n3984_), .B0(new_n3979_), .B1(new_n3973_), .Y(new_n3988_));
  OR2X1    g02986(.A(new_n3988_), .B(new_n3947_), .Y(new_n3989_));
  OR2X1    g02987(.A(new_n3972_), .B(new_n3968_), .Y(new_n3990_));
  XOR2X1   g02988(.A(new_n3932_), .B(new_n3926_), .Y(new_n3991_));
  XOR2X1   g02989(.A(new_n3991_), .B(new_n3990_), .Y(new_n3992_));
  NAND2X1  g02990(.A(new_n3897_), .B(new_n3895_), .Y(new_n3993_));
  XOR2X1   g02991(.A(new_n3862_), .B(new_n3856_), .Y(new_n3994_));
  XOR2X1   g02992(.A(new_n3994_), .B(new_n3993_), .Y(new_n3995_));
  NOR2X1   g02993(.A(new_n3995_), .B(new_n3992_), .Y(new_n3996_));
  NAND3X1  g02994(.A(new_n3996_), .B(new_n3989_), .C(new_n3981_), .Y(new_n3997_));
  AND2X1   g02995(.A(new_n3980_), .B(new_n3947_), .Y(new_n3998_));
  NOR2X1   g02996(.A(new_n3988_), .B(new_n3947_), .Y(new_n3999_));
  OR2X1    g02997(.A(new_n3995_), .B(new_n3992_), .Y(new_n4000_));
  OAI21X1  g02998(.A0(new_n3999_), .A1(new_n3998_), .B0(new_n4000_), .Y(new_n4001_));
  AOI21X1  g02999(.A0(new_n4001_), .A1(new_n3997_), .B0(new_n3919_), .Y(new_n4002_));
  AOI21X1  g03000(.A0(new_n3875_), .A1(new_n3871_), .B0(new_n3870_), .Y(new_n4003_));
  AND2X1   g03001(.A(new_n3908_), .B(new_n3877_), .Y(new_n4004_));
  AOI21X1  g03002(.A0(new_n3918_), .A1(new_n4003_), .B0(new_n4004_), .Y(new_n4005_));
  NAND3X1  g03003(.A(new_n4000_), .B(new_n3989_), .C(new_n3981_), .Y(new_n4006_));
  OAI21X1  g03004(.A0(new_n3999_), .A1(new_n3998_), .B0(new_n3996_), .Y(new_n4007_));
  AOI21X1  g03005(.A0(new_n4007_), .A1(new_n4006_), .B0(new_n4005_), .Y(new_n4008_));
  NOR2X1   g03006(.A(new_n3972_), .B(new_n3968_), .Y(new_n4009_));
  XOR2X1   g03007(.A(new_n3991_), .B(new_n4009_), .Y(new_n4010_));
  XOR2X1   g03008(.A(new_n3995_), .B(new_n4010_), .Y(new_n4011_));
  INVX1    g03009(.A(\A[961] ), .Y(new_n4012_));
  OR2X1    g03010(.A(\A[962] ), .B(new_n4012_), .Y(new_n4013_));
  INVX1    g03011(.A(\A[963] ), .Y(new_n4014_));
  AOI21X1  g03012(.A0(\A[962] ), .A1(new_n4012_), .B0(new_n4014_), .Y(new_n4015_));
  XOR2X1   g03013(.A(\A[962] ), .B(\A[961] ), .Y(new_n4016_));
  AND2X1   g03014(.A(new_n4016_), .B(new_n4014_), .Y(new_n4017_));
  AOI21X1  g03015(.A0(new_n4015_), .A1(new_n4013_), .B0(new_n4017_), .Y(new_n4018_));
  INVX1    g03016(.A(\A[966] ), .Y(new_n4019_));
  INVX1    g03017(.A(\A[964] ), .Y(new_n4020_));
  OR2X1    g03018(.A(\A[965] ), .B(new_n4020_), .Y(new_n4021_));
  AOI21X1  g03019(.A0(\A[965] ), .A1(new_n4020_), .B0(new_n4019_), .Y(new_n4022_));
  XOR2X1   g03020(.A(\A[965] ), .B(\A[964] ), .Y(new_n4023_));
  AOI22X1  g03021(.A0(new_n4023_), .A1(new_n4019_), .B0(new_n4022_), .B1(new_n4021_), .Y(new_n4024_));
  AND2X1   g03022(.A(\A[965] ), .B(\A[964] ), .Y(new_n4025_));
  AOI21X1  g03023(.A0(new_n4023_), .A1(\A[966] ), .B0(new_n4025_), .Y(new_n4026_));
  AND2X1   g03024(.A(\A[962] ), .B(\A[961] ), .Y(new_n4027_));
  AOI21X1  g03025(.A0(new_n4016_), .A1(\A[963] ), .B0(new_n4027_), .Y(new_n4028_));
  XOR2X1   g03026(.A(new_n4024_), .B(new_n4018_), .Y(new_n4029_));
  INVX1    g03027(.A(\A[955] ), .Y(new_n4030_));
  OR2X1    g03028(.A(\A[956] ), .B(new_n4030_), .Y(new_n4031_));
  INVX1    g03029(.A(\A[957] ), .Y(new_n4032_));
  AOI21X1  g03030(.A0(\A[956] ), .A1(new_n4030_), .B0(new_n4032_), .Y(new_n4033_));
  XOR2X1   g03031(.A(\A[956] ), .B(\A[955] ), .Y(new_n4034_));
  AND2X1   g03032(.A(new_n4034_), .B(new_n4032_), .Y(new_n4035_));
  AOI21X1  g03033(.A0(new_n4033_), .A1(new_n4031_), .B0(new_n4035_), .Y(new_n4036_));
  INVX1    g03034(.A(\A[960] ), .Y(new_n4037_));
  INVX1    g03035(.A(\A[958] ), .Y(new_n4038_));
  OR2X1    g03036(.A(\A[959] ), .B(new_n4038_), .Y(new_n4039_));
  AOI21X1  g03037(.A0(\A[959] ), .A1(new_n4038_), .B0(new_n4037_), .Y(new_n4040_));
  XOR2X1   g03038(.A(\A[959] ), .B(\A[958] ), .Y(new_n4041_));
  AOI22X1  g03039(.A0(new_n4041_), .A1(new_n4037_), .B0(new_n4040_), .B1(new_n4039_), .Y(new_n4042_));
  AND2X1   g03040(.A(\A[959] ), .B(\A[958] ), .Y(new_n4043_));
  AOI21X1  g03041(.A0(new_n4041_), .A1(\A[960] ), .B0(new_n4043_), .Y(new_n4044_));
  AND2X1   g03042(.A(\A[956] ), .B(\A[955] ), .Y(new_n4045_));
  AOI21X1  g03043(.A0(new_n4034_), .A1(\A[957] ), .B0(new_n4045_), .Y(new_n4046_));
  XOR2X1   g03044(.A(new_n4042_), .B(new_n4036_), .Y(new_n4047_));
  XOR2X1   g03045(.A(new_n4047_), .B(new_n4029_), .Y(new_n4048_));
  INVX1    g03046(.A(\A[949] ), .Y(new_n4049_));
  OR2X1    g03047(.A(\A[950] ), .B(new_n4049_), .Y(new_n4050_));
  INVX1    g03048(.A(\A[951] ), .Y(new_n4051_));
  AOI21X1  g03049(.A0(\A[950] ), .A1(new_n4049_), .B0(new_n4051_), .Y(new_n4052_));
  AND2X1   g03050(.A(new_n4052_), .B(new_n4050_), .Y(new_n4053_));
  XOR2X1   g03051(.A(\A[950] ), .B(\A[949] ), .Y(new_n4054_));
  AND2X1   g03052(.A(new_n4054_), .B(new_n4051_), .Y(new_n4055_));
  OR2X1    g03053(.A(new_n4055_), .B(new_n4053_), .Y(new_n4056_));
  INVX1    g03054(.A(\A[954] ), .Y(new_n4057_));
  INVX1    g03055(.A(\A[952] ), .Y(new_n4058_));
  OR2X1    g03056(.A(\A[953] ), .B(new_n4058_), .Y(new_n4059_));
  AOI21X1  g03057(.A0(\A[953] ), .A1(new_n4058_), .B0(new_n4057_), .Y(new_n4060_));
  XOR2X1   g03058(.A(\A[953] ), .B(\A[952] ), .Y(new_n4061_));
  AOI22X1  g03059(.A0(new_n4061_), .A1(new_n4057_), .B0(new_n4060_), .B1(new_n4059_), .Y(new_n4062_));
  AND2X1   g03060(.A(\A[953] ), .B(\A[952] ), .Y(new_n4063_));
  AOI21X1  g03061(.A0(new_n4061_), .A1(\A[954] ), .B0(new_n4063_), .Y(new_n4064_));
  AND2X1   g03062(.A(\A[950] ), .B(\A[949] ), .Y(new_n4065_));
  AOI21X1  g03063(.A0(new_n4054_), .A1(\A[951] ), .B0(new_n4065_), .Y(new_n4066_));
  XOR2X1   g03064(.A(new_n4062_), .B(new_n4056_), .Y(new_n4067_));
  INVX1    g03065(.A(\A[943] ), .Y(new_n4068_));
  OR2X1    g03066(.A(\A[944] ), .B(new_n4068_), .Y(new_n4069_));
  INVX1    g03067(.A(\A[945] ), .Y(new_n4070_));
  AOI21X1  g03068(.A0(\A[944] ), .A1(new_n4068_), .B0(new_n4070_), .Y(new_n4071_));
  XOR2X1   g03069(.A(\A[944] ), .B(\A[943] ), .Y(new_n4072_));
  AND2X1   g03070(.A(new_n4072_), .B(new_n4070_), .Y(new_n4073_));
  AOI21X1  g03071(.A0(new_n4071_), .A1(new_n4069_), .B0(new_n4073_), .Y(new_n4074_));
  INVX1    g03072(.A(\A[948] ), .Y(new_n4075_));
  INVX1    g03073(.A(\A[946] ), .Y(new_n4076_));
  OR2X1    g03074(.A(\A[947] ), .B(new_n4076_), .Y(new_n4077_));
  AOI21X1  g03075(.A0(\A[947] ), .A1(new_n4076_), .B0(new_n4075_), .Y(new_n4078_));
  XOR2X1   g03076(.A(\A[947] ), .B(\A[946] ), .Y(new_n4079_));
  AOI22X1  g03077(.A0(new_n4079_), .A1(new_n4075_), .B0(new_n4078_), .B1(new_n4077_), .Y(new_n4080_));
  AND2X1   g03078(.A(\A[947] ), .B(\A[946] ), .Y(new_n4081_));
  AOI21X1  g03079(.A0(new_n4079_), .A1(\A[948] ), .B0(new_n4081_), .Y(new_n4082_));
  AND2X1   g03080(.A(\A[944] ), .B(\A[943] ), .Y(new_n4083_));
  AOI21X1  g03081(.A0(new_n4072_), .A1(\A[945] ), .B0(new_n4083_), .Y(new_n4084_));
  XOR2X1   g03082(.A(new_n4080_), .B(new_n4074_), .Y(new_n4085_));
  XOR2X1   g03083(.A(new_n4085_), .B(new_n4067_), .Y(new_n4086_));
  XOR2X1   g03084(.A(new_n4086_), .B(new_n4048_), .Y(new_n4087_));
  OR4X1    g03085(.A(new_n4087_), .B(new_n4011_), .C(new_n4008_), .D(new_n4002_), .Y(new_n4088_));
  OAI22X1  g03086(.A0(new_n4087_), .A1(new_n4011_), .B0(new_n4008_), .B1(new_n4002_), .Y(new_n4089_));
  AND2X1   g03087(.A(new_n4089_), .B(new_n4088_), .Y(new_n4090_));
  AND2X1   g03088(.A(new_n4033_), .B(new_n4031_), .Y(new_n4091_));
  OR2X1    g03089(.A(new_n4035_), .B(new_n4091_), .Y(new_n4092_));
  XOR2X1   g03090(.A(new_n4042_), .B(new_n4092_), .Y(new_n4093_));
  XOR2X1   g03091(.A(new_n4046_), .B(new_n4044_), .Y(new_n4094_));
  NOR2X1   g03092(.A(new_n4042_), .B(new_n4036_), .Y(new_n4095_));
  NOR2X1   g03093(.A(new_n4046_), .B(new_n4044_), .Y(new_n4096_));
  AOI21X1  g03094(.A0(new_n4095_), .A1(new_n4094_), .B0(new_n4096_), .Y(new_n4097_));
  XOR2X1   g03095(.A(new_n4095_), .B(new_n4094_), .Y(new_n4098_));
  OAI21X1  g03096(.A0(new_n4097_), .A1(new_n4093_), .B0(new_n4098_), .Y(new_n4099_));
  AND2X1   g03097(.A(new_n4015_), .B(new_n4013_), .Y(new_n4100_));
  OR2X1    g03098(.A(new_n4017_), .B(new_n4100_), .Y(new_n4101_));
  XOR2X1   g03099(.A(new_n4024_), .B(new_n4101_), .Y(new_n4102_));
  NOR4X1   g03100(.A(new_n4028_), .B(new_n4026_), .C(new_n4024_), .D(new_n4018_), .Y(new_n4103_));
  NOR4X1   g03101(.A(new_n4046_), .B(new_n4044_), .C(new_n4042_), .D(new_n4036_), .Y(new_n4104_));
  OR4X1    g03102(.A(new_n4104_), .B(new_n4093_), .C(new_n4103_), .D(new_n4102_), .Y(new_n4105_));
  XOR2X1   g03103(.A(new_n4028_), .B(new_n4026_), .Y(new_n4106_));
  NOR2X1   g03104(.A(new_n4024_), .B(new_n4018_), .Y(new_n4107_));
  NOR2X1   g03105(.A(new_n4028_), .B(new_n4026_), .Y(new_n4108_));
  AOI21X1  g03106(.A0(new_n4107_), .A1(new_n4106_), .B0(new_n4108_), .Y(new_n4109_));
  XOR2X1   g03107(.A(new_n4107_), .B(new_n4106_), .Y(new_n4110_));
  OAI21X1  g03108(.A0(new_n4109_), .A1(new_n4102_), .B0(new_n4110_), .Y(new_n4111_));
  XOR2X1   g03109(.A(new_n4111_), .B(new_n4105_), .Y(new_n4112_));
  NAND2X1  g03110(.A(new_n4112_), .B(new_n4099_), .Y(new_n4113_));
  XOR2X1   g03111(.A(new_n4042_), .B(new_n4036_), .Y(new_n4114_));
  AND2X1   g03112(.A(new_n4041_), .B(\A[960] ), .Y(new_n4115_));
  OR2X1    g03113(.A(new_n4115_), .B(new_n4043_), .Y(new_n4116_));
  XOR2X1   g03114(.A(new_n4046_), .B(new_n4116_), .Y(new_n4117_));
  OR2X1    g03115(.A(new_n4042_), .B(new_n4036_), .Y(new_n4118_));
  OR2X1    g03116(.A(new_n4046_), .B(new_n4044_), .Y(new_n4119_));
  OAI21X1  g03117(.A0(new_n4118_), .A1(new_n4117_), .B0(new_n4119_), .Y(new_n4120_));
  XOR2X1   g03118(.A(new_n4095_), .B(new_n4117_), .Y(new_n4121_));
  AOI21X1  g03119(.A0(new_n4120_), .A1(new_n4114_), .B0(new_n4121_), .Y(new_n4122_));
  AND2X1   g03120(.A(new_n4111_), .B(new_n4105_), .Y(new_n4123_));
  OR2X1    g03121(.A(new_n4024_), .B(new_n4018_), .Y(new_n4124_));
  XOR2X1   g03122(.A(new_n4124_), .B(new_n4106_), .Y(new_n4125_));
  OR4X1    g03123(.A(new_n4093_), .B(new_n4103_), .C(new_n4125_), .D(new_n4102_), .Y(new_n4126_));
  OAI22X1  g03124(.A0(new_n4121_), .A1(new_n4097_), .B0(new_n4109_), .B1(new_n4102_), .Y(new_n4127_));
  NOR2X1   g03125(.A(new_n4127_), .B(new_n4126_), .Y(new_n4128_));
  OAI21X1  g03126(.A0(new_n4128_), .A1(new_n4123_), .B0(new_n4122_), .Y(new_n4129_));
  INVX1    g03127(.A(new_n4048_), .Y(new_n4130_));
  NOR2X1   g03128(.A(new_n4086_), .B(new_n4130_), .Y(new_n4131_));
  NAND3X1  g03129(.A(new_n4131_), .B(new_n4129_), .C(new_n4113_), .Y(new_n4132_));
  AND2X1   g03130(.A(new_n4112_), .B(new_n4099_), .Y(new_n4133_));
  NAND2X1  g03131(.A(new_n4111_), .B(new_n4105_), .Y(new_n4134_));
  OR2X1    g03132(.A(new_n4127_), .B(new_n4126_), .Y(new_n4135_));
  AOI21X1  g03133(.A0(new_n4135_), .A1(new_n4134_), .B0(new_n4099_), .Y(new_n4136_));
  OR2X1    g03134(.A(new_n4086_), .B(new_n4130_), .Y(new_n4137_));
  OAI21X1  g03135(.A0(new_n4136_), .A1(new_n4133_), .B0(new_n4137_), .Y(new_n4138_));
  AND2X1   g03136(.A(new_n4071_), .B(new_n4069_), .Y(new_n4139_));
  OR2X1    g03137(.A(new_n4073_), .B(new_n4139_), .Y(new_n4140_));
  XOR2X1   g03138(.A(new_n4080_), .B(new_n4140_), .Y(new_n4141_));
  XOR2X1   g03139(.A(new_n4084_), .B(new_n4082_), .Y(new_n4142_));
  NOR2X1   g03140(.A(new_n4080_), .B(new_n4074_), .Y(new_n4143_));
  NOR2X1   g03141(.A(new_n4084_), .B(new_n4082_), .Y(new_n4144_));
  AOI21X1  g03142(.A0(new_n4143_), .A1(new_n4142_), .B0(new_n4144_), .Y(new_n4145_));
  XOR2X1   g03143(.A(new_n4143_), .B(new_n4142_), .Y(new_n4146_));
  OAI21X1  g03144(.A0(new_n4145_), .A1(new_n4141_), .B0(new_n4146_), .Y(new_n4147_));
  XOR2X1   g03145(.A(new_n4062_), .B(new_n4056_), .Y(new_n4148_));
  AOI21X1  g03146(.A0(new_n4052_), .A1(new_n4050_), .B0(new_n4055_), .Y(new_n4149_));
  NOR4X1   g03147(.A(new_n4066_), .B(new_n4064_), .C(new_n4062_), .D(new_n4149_), .Y(new_n4150_));
  NOR4X1   g03148(.A(new_n4084_), .B(new_n4082_), .C(new_n4080_), .D(new_n4074_), .Y(new_n4151_));
  OR4X1    g03149(.A(new_n4151_), .B(new_n4141_), .C(new_n4150_), .D(new_n4148_), .Y(new_n4152_));
  XOR2X1   g03150(.A(new_n4066_), .B(new_n4064_), .Y(new_n4153_));
  NOR2X1   g03151(.A(new_n4062_), .B(new_n4149_), .Y(new_n4154_));
  NOR2X1   g03152(.A(new_n4066_), .B(new_n4064_), .Y(new_n4155_));
  AOI21X1  g03153(.A0(new_n4154_), .A1(new_n4153_), .B0(new_n4155_), .Y(new_n4156_));
  XOR2X1   g03154(.A(new_n4154_), .B(new_n4153_), .Y(new_n4157_));
  OAI21X1  g03155(.A0(new_n4156_), .A1(new_n4148_), .B0(new_n4157_), .Y(new_n4158_));
  XOR2X1   g03156(.A(new_n4158_), .B(new_n4152_), .Y(new_n4159_));
  AND2X1   g03157(.A(new_n4158_), .B(new_n4152_), .Y(new_n4160_));
  OR2X1    g03158(.A(new_n4062_), .B(new_n4149_), .Y(new_n4161_));
  XOR2X1   g03159(.A(new_n4161_), .B(new_n4153_), .Y(new_n4162_));
  OR4X1    g03160(.A(new_n4141_), .B(new_n4150_), .C(new_n4162_), .D(new_n4148_), .Y(new_n4163_));
  AND2X1   g03161(.A(new_n4079_), .B(\A[948] ), .Y(new_n4164_));
  OR2X1    g03162(.A(new_n4164_), .B(new_n4081_), .Y(new_n4165_));
  XOR2X1   g03163(.A(new_n4084_), .B(new_n4165_), .Y(new_n4166_));
  XOR2X1   g03164(.A(new_n4143_), .B(new_n4166_), .Y(new_n4167_));
  OAI22X1  g03165(.A0(new_n4167_), .A1(new_n4145_), .B0(new_n4156_), .B1(new_n4148_), .Y(new_n4168_));
  NOR2X1   g03166(.A(new_n4168_), .B(new_n4163_), .Y(new_n4169_));
  OR2X1    g03167(.A(new_n4169_), .B(new_n4160_), .Y(new_n4170_));
  MX2X1    g03168(.A(new_n4170_), .B(new_n4159_), .S0(new_n4147_), .Y(new_n4171_));
  AOI21X1  g03169(.A0(new_n4138_), .A1(new_n4132_), .B0(new_n4171_), .Y(new_n4172_));
  INVX1    g03170(.A(new_n4147_), .Y(new_n4173_));
  AND2X1   g03171(.A(new_n4159_), .B(new_n4147_), .Y(new_n4174_));
  AOI21X1  g03172(.A0(new_n4170_), .A1(new_n4173_), .B0(new_n4174_), .Y(new_n4175_));
  NAND3X1  g03173(.A(new_n4137_), .B(new_n4129_), .C(new_n4113_), .Y(new_n4176_));
  OAI21X1  g03174(.A0(new_n4136_), .A1(new_n4133_), .B0(new_n4131_), .Y(new_n4177_));
  AOI21X1  g03175(.A0(new_n4177_), .A1(new_n4176_), .B0(new_n4175_), .Y(new_n4178_));
  NOR2X1   g03176(.A(new_n4178_), .B(new_n4172_), .Y(new_n4179_));
  INVX1    g03177(.A(new_n4179_), .Y(new_n4180_));
  NOR2X1   g03178(.A(new_n4087_), .B(new_n4011_), .Y(new_n4181_));
  OR2X1    g03179(.A(new_n4008_), .B(new_n4002_), .Y(new_n4182_));
  NOR3X1   g03180(.A(new_n4181_), .B(new_n4008_), .C(new_n4002_), .Y(new_n4183_));
  AOI21X1  g03181(.A0(new_n4182_), .A1(new_n4181_), .B0(new_n4183_), .Y(new_n4184_));
  OR2X1    g03182(.A(new_n4184_), .B(new_n4179_), .Y(new_n4185_));
  OAI21X1  g03183(.A0(new_n4180_), .A1(new_n4090_), .B0(new_n4185_), .Y(new_n4186_));
  INVX1    g03184(.A(\A[9] ), .Y(new_n4187_));
  INVX1    g03185(.A(\A[8] ), .Y(new_n4188_));
  OR2X1    g03186(.A(new_n4188_), .B(\A[7] ), .Y(new_n4189_));
  AOI21X1  g03187(.A0(new_n4188_), .A1(\A[7] ), .B0(new_n4187_), .Y(new_n4190_));
  XOR2X1   g03188(.A(\A[8] ), .B(\A[7] ), .Y(new_n4191_));
  AOI22X1  g03189(.A0(new_n4191_), .A1(new_n4187_), .B0(new_n4190_), .B1(new_n4189_), .Y(new_n4192_));
  INVX1    g03190(.A(\A[12] ), .Y(new_n4193_));
  INVX1    g03191(.A(\A[11] ), .Y(new_n4194_));
  OR2X1    g03192(.A(new_n4194_), .B(\A[10] ), .Y(new_n4195_));
  AOI21X1  g03193(.A0(new_n4194_), .A1(\A[10] ), .B0(new_n4193_), .Y(new_n4196_));
  XOR2X1   g03194(.A(\A[11] ), .B(\A[10] ), .Y(new_n4197_));
  AOI22X1  g03195(.A0(new_n4197_), .A1(new_n4193_), .B0(new_n4196_), .B1(new_n4195_), .Y(new_n4198_));
  NOR2X1   g03196(.A(new_n4198_), .B(new_n4192_), .Y(new_n4199_));
  AND2X1   g03197(.A(\A[11] ), .B(\A[10] ), .Y(new_n4200_));
  AND2X1   g03198(.A(new_n4197_), .B(\A[12] ), .Y(new_n4201_));
  OR2X1    g03199(.A(new_n4201_), .B(new_n4200_), .Y(new_n4202_));
  AND2X1   g03200(.A(\A[8] ), .B(\A[7] ), .Y(new_n4203_));
  AOI21X1  g03201(.A0(new_n4191_), .A1(\A[9] ), .B0(new_n4203_), .Y(new_n4204_));
  XOR2X1   g03202(.A(new_n4204_), .B(new_n4202_), .Y(new_n4205_));
  XOR2X1   g03203(.A(new_n4205_), .B(new_n4199_), .Y(new_n4206_));
  XOR2X1   g03204(.A(new_n4198_), .B(new_n4192_), .Y(new_n4207_));
  OR2X1    g03205(.A(new_n4198_), .B(new_n4192_), .Y(new_n4208_));
  AOI21X1  g03206(.A0(new_n4197_), .A1(\A[12] ), .B0(new_n4200_), .Y(new_n4209_));
  OR2X1    g03207(.A(new_n4204_), .B(new_n4209_), .Y(new_n4210_));
  OAI21X1  g03208(.A0(new_n4205_), .A1(new_n4208_), .B0(new_n4210_), .Y(new_n4211_));
  AOI21X1  g03209(.A0(new_n4211_), .A1(new_n4207_), .B0(new_n4206_), .Y(new_n4212_));
  INVX1    g03210(.A(\A[7] ), .Y(new_n4213_));
  AND2X1   g03211(.A(\A[8] ), .B(new_n4213_), .Y(new_n4214_));
  OAI21X1  g03212(.A0(\A[8] ), .A1(new_n4213_), .B0(\A[9] ), .Y(new_n4215_));
  NAND2X1  g03213(.A(new_n4191_), .B(new_n4187_), .Y(new_n4216_));
  OAI21X1  g03214(.A0(new_n4215_), .A1(new_n4214_), .B0(new_n4216_), .Y(new_n4217_));
  XOR2X1   g03215(.A(new_n4198_), .B(new_n4217_), .Y(new_n4218_));
  AND2X1   g03216(.A(\A[17] ), .B(\A[16] ), .Y(new_n4219_));
  XOR2X1   g03217(.A(\A[17] ), .B(\A[16] ), .Y(new_n4220_));
  AOI21X1  g03218(.A0(new_n4220_), .A1(\A[18] ), .B0(new_n4219_), .Y(new_n4221_));
  AND2X1   g03219(.A(\A[14] ), .B(\A[13] ), .Y(new_n4222_));
  XOR2X1   g03220(.A(\A[14] ), .B(\A[13] ), .Y(new_n4223_));
  AOI21X1  g03221(.A0(new_n4223_), .A1(\A[15] ), .B0(new_n4222_), .Y(new_n4224_));
  INVX1    g03222(.A(\A[15] ), .Y(new_n4225_));
  INVX1    g03223(.A(\A[14] ), .Y(new_n4226_));
  OR2X1    g03224(.A(new_n4226_), .B(\A[13] ), .Y(new_n4227_));
  AOI21X1  g03225(.A0(new_n4226_), .A1(\A[13] ), .B0(new_n4225_), .Y(new_n4228_));
  AOI22X1  g03226(.A0(new_n4228_), .A1(new_n4227_), .B0(new_n4223_), .B1(new_n4225_), .Y(new_n4229_));
  INVX1    g03227(.A(\A[18] ), .Y(new_n4230_));
  INVX1    g03228(.A(\A[17] ), .Y(new_n4231_));
  OR2X1    g03229(.A(new_n4231_), .B(\A[16] ), .Y(new_n4232_));
  AOI21X1  g03230(.A0(new_n4231_), .A1(\A[16] ), .B0(new_n4230_), .Y(new_n4233_));
  AOI22X1  g03231(.A0(new_n4233_), .A1(new_n4232_), .B0(new_n4220_), .B1(new_n4230_), .Y(new_n4234_));
  NOR4X1   g03232(.A(new_n4234_), .B(new_n4229_), .C(new_n4224_), .D(new_n4221_), .Y(new_n4235_));
  NOR4X1   g03233(.A(new_n4204_), .B(new_n4209_), .C(new_n4198_), .D(new_n4192_), .Y(new_n4236_));
  INVX1    g03234(.A(\A[13] ), .Y(new_n4237_));
  AND2X1   g03235(.A(\A[14] ), .B(new_n4237_), .Y(new_n4238_));
  OAI21X1  g03236(.A0(\A[14] ), .A1(new_n4237_), .B0(\A[15] ), .Y(new_n4239_));
  NAND2X1  g03237(.A(new_n4223_), .B(new_n4225_), .Y(new_n4240_));
  OAI21X1  g03238(.A0(new_n4239_), .A1(new_n4238_), .B0(new_n4240_), .Y(new_n4241_));
  XOR2X1   g03239(.A(new_n4234_), .B(new_n4241_), .Y(new_n4242_));
  OR4X1    g03240(.A(new_n4242_), .B(new_n4236_), .C(new_n4235_), .D(new_n4218_), .Y(new_n4243_));
  AND2X1   g03241(.A(new_n4220_), .B(\A[18] ), .Y(new_n4244_));
  OR2X1    g03242(.A(new_n4244_), .B(new_n4219_), .Y(new_n4245_));
  XOR2X1   g03243(.A(new_n4224_), .B(new_n4245_), .Y(new_n4246_));
  OR2X1    g03244(.A(new_n4234_), .B(new_n4229_), .Y(new_n4247_));
  OR2X1    g03245(.A(new_n4224_), .B(new_n4221_), .Y(new_n4248_));
  OAI21X1  g03246(.A0(new_n4247_), .A1(new_n4246_), .B0(new_n4248_), .Y(new_n4249_));
  NOR2X1   g03247(.A(new_n4234_), .B(new_n4229_), .Y(new_n4250_));
  XOR2X1   g03248(.A(new_n4250_), .B(new_n4246_), .Y(new_n4251_));
  XOR2X1   g03249(.A(new_n4234_), .B(new_n4229_), .Y(new_n4252_));
  AOI21X1  g03250(.A0(new_n4252_), .A1(new_n4249_), .B0(new_n4251_), .Y(new_n4253_));
  XOR2X1   g03251(.A(new_n4253_), .B(new_n4243_), .Y(new_n4254_));
  XOR2X1   g03252(.A(new_n4205_), .B(new_n4208_), .Y(new_n4255_));
  XOR2X1   g03253(.A(new_n4204_), .B(new_n4209_), .Y(new_n4256_));
  NOR2X1   g03254(.A(new_n4204_), .B(new_n4209_), .Y(new_n4257_));
  AOI21X1  g03255(.A0(new_n4256_), .A1(new_n4199_), .B0(new_n4257_), .Y(new_n4258_));
  OAI21X1  g03256(.A0(new_n4258_), .A1(new_n4218_), .B0(new_n4255_), .Y(new_n4259_));
  XOR2X1   g03257(.A(new_n4224_), .B(new_n4221_), .Y(new_n4260_));
  NOR2X1   g03258(.A(new_n4224_), .B(new_n4221_), .Y(new_n4261_));
  AOI21X1  g03259(.A0(new_n4250_), .A1(new_n4260_), .B0(new_n4261_), .Y(new_n4262_));
  XOR2X1   g03260(.A(new_n4250_), .B(new_n4260_), .Y(new_n4263_));
  OAI21X1  g03261(.A0(new_n4242_), .A1(new_n4262_), .B0(new_n4263_), .Y(new_n4264_));
  NOR4X1   g03262(.A(new_n4242_), .B(new_n4236_), .C(new_n4251_), .D(new_n4218_), .Y(new_n4265_));
  OAI21X1  g03263(.A0(new_n4252_), .A1(new_n4263_), .B0(new_n4249_), .Y(new_n4266_));
  AOI22X1  g03264(.A0(new_n4266_), .A1(new_n4265_), .B0(new_n4264_), .B1(new_n4243_), .Y(new_n4267_));
  OR2X1    g03265(.A(new_n4267_), .B(new_n4259_), .Y(new_n4268_));
  OAI21X1  g03266(.A0(new_n4254_), .A1(new_n4212_), .B0(new_n4268_), .Y(new_n4269_));
  INVX1    g03267(.A(\A[21] ), .Y(new_n4270_));
  INVX1    g03268(.A(\A[20] ), .Y(new_n4271_));
  OR2X1    g03269(.A(new_n4271_), .B(\A[19] ), .Y(new_n4272_));
  AOI21X1  g03270(.A0(new_n4271_), .A1(\A[19] ), .B0(new_n4270_), .Y(new_n4273_));
  XOR2X1   g03271(.A(\A[20] ), .B(\A[19] ), .Y(new_n4274_));
  AOI22X1  g03272(.A0(new_n4274_), .A1(new_n4270_), .B0(new_n4273_), .B1(new_n4272_), .Y(new_n4275_));
  INVX1    g03273(.A(\A[24] ), .Y(new_n4276_));
  INVX1    g03274(.A(\A[23] ), .Y(new_n4277_));
  OR2X1    g03275(.A(new_n4277_), .B(\A[22] ), .Y(new_n4278_));
  AOI21X1  g03276(.A0(new_n4277_), .A1(\A[22] ), .B0(new_n4276_), .Y(new_n4279_));
  XOR2X1   g03277(.A(\A[23] ), .B(\A[22] ), .Y(new_n4280_));
  AOI22X1  g03278(.A0(new_n4280_), .A1(new_n4276_), .B0(new_n4279_), .B1(new_n4278_), .Y(new_n4281_));
  OR2X1    g03279(.A(new_n4281_), .B(new_n4275_), .Y(new_n4282_));
  AND2X1   g03280(.A(\A[23] ), .B(\A[22] ), .Y(new_n4283_));
  AND2X1   g03281(.A(new_n4280_), .B(\A[24] ), .Y(new_n4284_));
  OR2X1    g03282(.A(new_n4284_), .B(new_n4283_), .Y(new_n4285_));
  AND2X1   g03283(.A(\A[20] ), .B(\A[19] ), .Y(new_n4286_));
  AOI21X1  g03284(.A0(new_n4274_), .A1(\A[21] ), .B0(new_n4286_), .Y(new_n4287_));
  XOR2X1   g03285(.A(new_n4287_), .B(new_n4285_), .Y(new_n4288_));
  XOR2X1   g03286(.A(new_n4288_), .B(new_n4282_), .Y(new_n4289_));
  INVX1    g03287(.A(\A[19] ), .Y(new_n4290_));
  AND2X1   g03288(.A(\A[20] ), .B(new_n4290_), .Y(new_n4291_));
  OAI21X1  g03289(.A0(\A[20] ), .A1(new_n4290_), .B0(\A[21] ), .Y(new_n4292_));
  NAND2X1  g03290(.A(new_n4274_), .B(new_n4270_), .Y(new_n4293_));
  OAI21X1  g03291(.A0(new_n4292_), .A1(new_n4291_), .B0(new_n4293_), .Y(new_n4294_));
  XOR2X1   g03292(.A(new_n4281_), .B(new_n4294_), .Y(new_n4295_));
  NOR2X1   g03293(.A(new_n4281_), .B(new_n4275_), .Y(new_n4296_));
  AOI21X1  g03294(.A0(new_n4280_), .A1(\A[24] ), .B0(new_n4283_), .Y(new_n4297_));
  XOR2X1   g03295(.A(new_n4287_), .B(new_n4297_), .Y(new_n4298_));
  NOR2X1   g03296(.A(new_n4287_), .B(new_n4297_), .Y(new_n4299_));
  AOI21X1  g03297(.A0(new_n4298_), .A1(new_n4296_), .B0(new_n4299_), .Y(new_n4300_));
  OAI21X1  g03298(.A0(new_n4300_), .A1(new_n4295_), .B0(new_n4289_), .Y(new_n4301_));
  AND2X1   g03299(.A(\A[29] ), .B(\A[28] ), .Y(new_n4302_));
  XOR2X1   g03300(.A(\A[29] ), .B(\A[28] ), .Y(new_n4303_));
  AOI21X1  g03301(.A0(new_n4303_), .A1(\A[30] ), .B0(new_n4302_), .Y(new_n4304_));
  AND2X1   g03302(.A(\A[26] ), .B(\A[25] ), .Y(new_n4305_));
  XOR2X1   g03303(.A(\A[26] ), .B(\A[25] ), .Y(new_n4306_));
  AOI21X1  g03304(.A0(new_n4306_), .A1(\A[27] ), .B0(new_n4305_), .Y(new_n4307_));
  INVX1    g03305(.A(\A[27] ), .Y(new_n4308_));
  INVX1    g03306(.A(\A[26] ), .Y(new_n4309_));
  OR2X1    g03307(.A(new_n4309_), .B(\A[25] ), .Y(new_n4310_));
  AOI21X1  g03308(.A0(new_n4309_), .A1(\A[25] ), .B0(new_n4308_), .Y(new_n4311_));
  AOI22X1  g03309(.A0(new_n4311_), .A1(new_n4310_), .B0(new_n4306_), .B1(new_n4308_), .Y(new_n4312_));
  INVX1    g03310(.A(\A[30] ), .Y(new_n4313_));
  INVX1    g03311(.A(\A[29] ), .Y(new_n4314_));
  OR2X1    g03312(.A(new_n4314_), .B(\A[28] ), .Y(new_n4315_));
  AOI21X1  g03313(.A0(new_n4314_), .A1(\A[28] ), .B0(new_n4313_), .Y(new_n4316_));
  AOI22X1  g03314(.A0(new_n4316_), .A1(new_n4315_), .B0(new_n4303_), .B1(new_n4313_), .Y(new_n4317_));
  NOR4X1   g03315(.A(new_n4317_), .B(new_n4312_), .C(new_n4307_), .D(new_n4304_), .Y(new_n4318_));
  NOR4X1   g03316(.A(new_n4287_), .B(new_n4297_), .C(new_n4281_), .D(new_n4275_), .Y(new_n4319_));
  INVX1    g03317(.A(\A[25] ), .Y(new_n4320_));
  AND2X1   g03318(.A(\A[26] ), .B(new_n4320_), .Y(new_n4321_));
  OAI21X1  g03319(.A0(\A[26] ), .A1(new_n4320_), .B0(\A[27] ), .Y(new_n4322_));
  NAND2X1  g03320(.A(new_n4306_), .B(new_n4308_), .Y(new_n4323_));
  OAI21X1  g03321(.A0(new_n4322_), .A1(new_n4321_), .B0(new_n4323_), .Y(new_n4324_));
  XOR2X1   g03322(.A(new_n4317_), .B(new_n4324_), .Y(new_n4325_));
  OR4X1    g03323(.A(new_n4325_), .B(new_n4319_), .C(new_n4318_), .D(new_n4295_), .Y(new_n4326_));
  XOR2X1   g03324(.A(new_n4307_), .B(new_n4304_), .Y(new_n4327_));
  NOR2X1   g03325(.A(new_n4317_), .B(new_n4312_), .Y(new_n4328_));
  NOR2X1   g03326(.A(new_n4307_), .B(new_n4304_), .Y(new_n4329_));
  AOI21X1  g03327(.A0(new_n4328_), .A1(new_n4327_), .B0(new_n4329_), .Y(new_n4330_));
  XOR2X1   g03328(.A(new_n4328_), .B(new_n4327_), .Y(new_n4331_));
  OAI21X1  g03329(.A0(new_n4325_), .A1(new_n4330_), .B0(new_n4331_), .Y(new_n4332_));
  XOR2X1   g03330(.A(new_n4332_), .B(new_n4326_), .Y(new_n4333_));
  NAND2X1  g03331(.A(new_n4333_), .B(new_n4301_), .Y(new_n4334_));
  OR2X1    g03332(.A(new_n4325_), .B(new_n4318_), .Y(new_n4335_));
  XOR2X1   g03333(.A(new_n4281_), .B(new_n4275_), .Y(new_n4336_));
  XOR2X1   g03334(.A(new_n4336_), .B(new_n4335_), .Y(new_n4337_));
  OR2X1    g03335(.A(new_n4242_), .B(new_n4235_), .Y(new_n4338_));
  XOR2X1   g03336(.A(new_n4198_), .B(new_n4192_), .Y(new_n4339_));
  XOR2X1   g03337(.A(new_n4339_), .B(new_n4338_), .Y(new_n4340_));
  OR2X1    g03338(.A(new_n4340_), .B(new_n4337_), .Y(new_n4341_));
  XOR2X1   g03339(.A(new_n4288_), .B(new_n4296_), .Y(new_n4342_));
  XOR2X1   g03340(.A(new_n4281_), .B(new_n4275_), .Y(new_n4343_));
  OR2X1    g03341(.A(new_n4287_), .B(new_n4297_), .Y(new_n4344_));
  OAI21X1  g03342(.A0(new_n4288_), .A1(new_n4282_), .B0(new_n4344_), .Y(new_n4345_));
  AOI21X1  g03343(.A0(new_n4345_), .A1(new_n4343_), .B0(new_n4342_), .Y(new_n4346_));
  NOR4X1   g03344(.A(new_n4325_), .B(new_n4319_), .C(new_n4318_), .D(new_n4295_), .Y(new_n4347_));
  AND2X1   g03345(.A(new_n4303_), .B(\A[30] ), .Y(new_n4348_));
  OR2X1    g03346(.A(new_n4348_), .B(new_n4302_), .Y(new_n4349_));
  XOR2X1   g03347(.A(new_n4307_), .B(new_n4349_), .Y(new_n4350_));
  OR2X1    g03348(.A(new_n4317_), .B(new_n4312_), .Y(new_n4351_));
  OR2X1    g03349(.A(new_n4307_), .B(new_n4304_), .Y(new_n4352_));
  OAI21X1  g03350(.A0(new_n4351_), .A1(new_n4350_), .B0(new_n4352_), .Y(new_n4353_));
  XOR2X1   g03351(.A(new_n4328_), .B(new_n4350_), .Y(new_n4354_));
  XOR2X1   g03352(.A(new_n4317_), .B(new_n4312_), .Y(new_n4355_));
  AOI21X1  g03353(.A0(new_n4355_), .A1(new_n4353_), .B0(new_n4354_), .Y(new_n4356_));
  OR4X1    g03354(.A(new_n4325_), .B(new_n4319_), .C(new_n4354_), .D(new_n4295_), .Y(new_n4357_));
  AOI21X1  g03355(.A0(new_n4325_), .A1(new_n4354_), .B0(new_n4330_), .Y(new_n4358_));
  OAI22X1  g03356(.A0(new_n4358_), .A1(new_n4357_), .B0(new_n4356_), .B1(new_n4347_), .Y(new_n4359_));
  AOI21X1  g03357(.A0(new_n4359_), .A1(new_n4346_), .B0(new_n4341_), .Y(new_n4360_));
  MX2X1    g03358(.A(new_n4359_), .B(new_n4333_), .S0(new_n4301_), .Y(new_n4361_));
  AOI22X1  g03359(.A0(new_n4361_), .A1(new_n4341_), .B0(new_n4360_), .B1(new_n4334_), .Y(new_n4362_));
  OR2X1    g03360(.A(new_n4362_), .B(new_n4269_), .Y(new_n4363_));
  XOR2X1   g03361(.A(new_n4340_), .B(new_n4337_), .Y(new_n4364_));
  INVX1    g03362(.A(\A[991] ), .Y(new_n4365_));
  OR2X1    g03363(.A(\A[992] ), .B(new_n4365_), .Y(new_n4366_));
  INVX1    g03364(.A(\A[993] ), .Y(new_n4367_));
  AOI21X1  g03365(.A0(\A[992] ), .A1(new_n4365_), .B0(new_n4367_), .Y(new_n4368_));
  XOR2X1   g03366(.A(\A[992] ), .B(\A[991] ), .Y(new_n4369_));
  AND2X1   g03367(.A(new_n4369_), .B(new_n4367_), .Y(new_n4370_));
  AOI21X1  g03368(.A0(new_n4368_), .A1(new_n4366_), .B0(new_n4370_), .Y(new_n4371_));
  INVX1    g03369(.A(\A[996] ), .Y(new_n4372_));
  INVX1    g03370(.A(\A[994] ), .Y(new_n4373_));
  OR2X1    g03371(.A(\A[995] ), .B(new_n4373_), .Y(new_n4374_));
  AOI21X1  g03372(.A0(\A[995] ), .A1(new_n4373_), .B0(new_n4372_), .Y(new_n4375_));
  XOR2X1   g03373(.A(\A[995] ), .B(\A[994] ), .Y(new_n4376_));
  AOI22X1  g03374(.A0(new_n4376_), .A1(new_n4372_), .B0(new_n4375_), .B1(new_n4374_), .Y(new_n4377_));
  AND2X1   g03375(.A(\A[995] ), .B(\A[994] ), .Y(new_n4378_));
  AOI21X1  g03376(.A0(new_n4376_), .A1(\A[996] ), .B0(new_n4378_), .Y(new_n4379_));
  AND2X1   g03377(.A(\A[992] ), .B(\A[991] ), .Y(new_n4380_));
  AOI21X1  g03378(.A0(new_n4369_), .A1(\A[993] ), .B0(new_n4380_), .Y(new_n4381_));
  XOR2X1   g03379(.A(new_n4377_), .B(new_n4371_), .Y(new_n4382_));
  INVX1    g03380(.A(\A[6] ), .Y(new_n4383_));
  INVX1    g03381(.A(\A[1] ), .Y(new_n4384_));
  AND2X1   g03382(.A(new_n4384_), .B(\A[0] ), .Y(new_n4385_));
  INVX1    g03383(.A(\A[2] ), .Y(new_n4386_));
  XOR2X1   g03384(.A(\A[1] ), .B(\A[0] ), .Y(new_n4387_));
  NAND2X1  g03385(.A(new_n4387_), .B(new_n4386_), .Y(new_n4388_));
  OAI21X1  g03386(.A0(new_n4384_), .A1(\A[0] ), .B0(\A[2] ), .Y(new_n4389_));
  OAI21X1  g03387(.A0(new_n4389_), .A1(new_n4385_), .B0(new_n4388_), .Y(new_n4390_));
  NAND2X1  g03388(.A(new_n4390_), .B(new_n4383_), .Y(new_n4391_));
  INVX1    g03389(.A(\A[3] ), .Y(new_n4392_));
  AND2X1   g03390(.A(\A[4] ), .B(new_n4392_), .Y(new_n4393_));
  OAI21X1  g03391(.A0(\A[4] ), .A1(new_n4392_), .B0(\A[5] ), .Y(new_n4394_));
  XOR2X1   g03392(.A(\A[4] ), .B(new_n4392_), .Y(new_n4395_));
  OAI22X1  g03393(.A0(new_n4395_), .A1(\A[5] ), .B0(new_n4394_), .B1(new_n4393_), .Y(new_n4396_));
  AOI21X1  g03394(.A0(new_n4387_), .A1(new_n4386_), .B0(new_n4383_), .Y(new_n4397_));
  OAI21X1  g03395(.A0(new_n4389_), .A1(new_n4385_), .B0(new_n4397_), .Y(new_n4398_));
  AND2X1   g03396(.A(new_n4398_), .B(new_n4396_), .Y(new_n4399_));
  AND2X1   g03397(.A(new_n4399_), .B(new_n4391_), .Y(new_n4400_));
  INVX1    g03398(.A(\A[997] ), .Y(new_n4401_));
  OR2X1    g03399(.A(\A[998] ), .B(new_n4401_), .Y(new_n4402_));
  INVX1    g03400(.A(\A[999] ), .Y(new_n4403_));
  AOI21X1  g03401(.A0(\A[998] ), .A1(new_n4401_), .B0(new_n4403_), .Y(new_n4404_));
  AND2X1   g03402(.A(new_n4404_), .B(new_n4402_), .Y(new_n4405_));
  XOR2X1   g03403(.A(\A[998] ), .B(\A[997] ), .Y(new_n4406_));
  AND2X1   g03404(.A(new_n4406_), .B(new_n4403_), .Y(new_n4407_));
  OR2X1    g03405(.A(new_n4407_), .B(new_n4405_), .Y(new_n4408_));
  OR2X1    g03406(.A(new_n4389_), .B(new_n4385_), .Y(new_n4409_));
  AOI22X1  g03407(.A0(new_n4397_), .A1(new_n4409_), .B0(new_n4390_), .B1(new_n4383_), .Y(new_n4410_));
  OAI21X1  g03408(.A0(new_n4410_), .A1(new_n4396_), .B0(new_n4408_), .Y(new_n4411_));
  OR2X1    g03409(.A(new_n4394_), .B(new_n4393_), .Y(new_n4412_));
  OR2X1    g03410(.A(new_n4395_), .B(\A[5] ), .Y(new_n4413_));
  AND2X1   g03411(.A(new_n4413_), .B(new_n4412_), .Y(new_n4414_));
  INVX1    g03412(.A(\A[0] ), .Y(new_n4415_));
  OR2X1    g03413(.A(\A[1] ), .B(new_n4415_), .Y(new_n4416_));
  AOI21X1  g03414(.A0(\A[1] ), .A1(new_n4415_), .B0(new_n4386_), .Y(new_n4417_));
  AOI22X1  g03415(.A0(new_n4417_), .A1(new_n4416_), .B0(new_n4387_), .B1(new_n4386_), .Y(new_n4418_));
  OAI21X1  g03416(.A0(new_n4418_), .A1(\A[6] ), .B0(new_n4398_), .Y(new_n4419_));
  AOI22X1  g03417(.A0(new_n4419_), .A1(new_n4414_), .B0(new_n4399_), .B1(new_n4391_), .Y(new_n4420_));
  OAI22X1  g03418(.A0(new_n4420_), .A1(new_n4408_), .B0(new_n4411_), .B1(new_n4400_), .Y(new_n4421_));
  XOR2X1   g03419(.A(new_n4421_), .B(new_n4382_), .Y(new_n4422_));
  NAND2X1  g03420(.A(new_n4422_), .B(new_n4364_), .Y(new_n4423_));
  AND2X1   g03421(.A(new_n4333_), .B(new_n4301_), .Y(new_n4424_));
  XOR2X1   g03422(.A(new_n4356_), .B(new_n4326_), .Y(new_n4425_));
  NOR4X1   g03423(.A(new_n4325_), .B(new_n4319_), .C(new_n4354_), .D(new_n4295_), .Y(new_n4426_));
  OAI21X1  g03424(.A0(new_n4355_), .A1(new_n4331_), .B0(new_n4353_), .Y(new_n4427_));
  AOI22X1  g03425(.A0(new_n4427_), .A1(new_n4426_), .B0(new_n4332_), .B1(new_n4326_), .Y(new_n4428_));
  MX2X1    g03426(.A(new_n4428_), .B(new_n4425_), .S0(new_n4301_), .Y(new_n4429_));
  OAI21X1  g03427(.A0(new_n4428_), .A1(new_n4301_), .B0(new_n4341_), .Y(new_n4430_));
  OAI22X1  g03428(.A0(new_n4430_), .A1(new_n4424_), .B0(new_n4429_), .B1(new_n4341_), .Y(new_n4431_));
  AOI21X1  g03429(.A0(new_n4431_), .A1(new_n4269_), .B0(new_n4423_), .Y(new_n4432_));
  NOR2X1   g03430(.A(new_n4340_), .B(new_n4337_), .Y(new_n4433_));
  OAI21X1  g03431(.A0(new_n4428_), .A1(new_n4301_), .B0(new_n4433_), .Y(new_n4434_));
  OAI22X1  g03432(.A0(new_n4429_), .A1(new_n4433_), .B0(new_n4434_), .B1(new_n4424_), .Y(new_n4435_));
  MX2X1    g03433(.A(new_n4435_), .B(new_n4431_), .S0(new_n4269_), .Y(new_n4436_));
  AOI22X1  g03434(.A0(new_n4436_), .A1(new_n4423_), .B0(new_n4432_), .B1(new_n4363_), .Y(new_n4437_));
  INVX1    g03435(.A(new_n4371_), .Y(new_n4438_));
  XOR2X1   g03436(.A(new_n4377_), .B(new_n4438_), .Y(new_n4439_));
  XOR2X1   g03437(.A(new_n4381_), .B(new_n4379_), .Y(new_n4440_));
  NOR2X1   g03438(.A(new_n4377_), .B(new_n4371_), .Y(new_n4441_));
  NOR2X1   g03439(.A(new_n4381_), .B(new_n4379_), .Y(new_n4442_));
  AOI21X1  g03440(.A0(new_n4441_), .A1(new_n4440_), .B0(new_n4442_), .Y(new_n4443_));
  XOR2X1   g03441(.A(new_n4441_), .B(new_n4440_), .Y(new_n4444_));
  OAI21X1  g03442(.A0(new_n4443_), .A1(new_n4439_), .B0(new_n4444_), .Y(new_n4445_));
  AND2X1   g03443(.A(\A[998] ), .B(\A[997] ), .Y(new_n4446_));
  AOI21X1  g03444(.A0(new_n4406_), .A1(\A[999] ), .B0(new_n4446_), .Y(new_n4447_));
  INVX1    g03445(.A(new_n4447_), .Y(new_n4448_));
  XOR2X1   g03446(.A(\A[4] ), .B(\A[3] ), .Y(new_n4449_));
  AND2X1   g03447(.A(\A[4] ), .B(\A[3] ), .Y(new_n4450_));
  AOI21X1  g03448(.A0(new_n4449_), .A1(\A[5] ), .B0(new_n4450_), .Y(new_n4451_));
  AND2X1   g03449(.A(\A[1] ), .B(\A[0] ), .Y(new_n4452_));
  AOI21X1  g03450(.A0(new_n4387_), .A1(\A[2] ), .B0(new_n4452_), .Y(new_n4453_));
  XOR2X1   g03451(.A(new_n4453_), .B(new_n4451_), .Y(new_n4454_));
  INVX1    g03452(.A(new_n4454_), .Y(new_n4455_));
  AOI21X1  g03453(.A0(new_n4390_), .A1(\A[6] ), .B0(new_n4454_), .Y(new_n4456_));
  OAI21X1  g03454(.A0(new_n4410_), .A1(new_n4414_), .B0(new_n4456_), .Y(new_n4457_));
  AOI22X1  g03455(.A0(new_n4419_), .A1(new_n4396_), .B0(new_n4390_), .B1(\A[6] ), .Y(new_n4458_));
  OAI21X1  g03456(.A0(new_n4458_), .A1(new_n4455_), .B0(new_n4457_), .Y(new_n4459_));
  AOI21X1  g03457(.A0(new_n4404_), .A1(new_n4402_), .B0(new_n4407_), .Y(new_n4460_));
  NOR2X1   g03458(.A(new_n4420_), .B(new_n4460_), .Y(new_n4461_));
  XOR2X1   g03459(.A(new_n4461_), .B(new_n4459_), .Y(new_n4462_));
  AND2X1   g03460(.A(new_n4462_), .B(new_n4448_), .Y(new_n4463_));
  AND2X1   g03461(.A(new_n4421_), .B(new_n4382_), .Y(new_n4464_));
  OR2X1    g03462(.A(new_n4420_), .B(new_n4460_), .Y(new_n4465_));
  AND2X1   g03463(.A(new_n4465_), .B(new_n4459_), .Y(new_n4466_));
  OAI21X1  g03464(.A0(new_n4465_), .A1(new_n4459_), .B0(new_n4447_), .Y(new_n4467_));
  OAI21X1  g03465(.A0(new_n4467_), .A1(new_n4466_), .B0(new_n4464_), .Y(new_n4468_));
  NAND2X1  g03466(.A(new_n4465_), .B(new_n4459_), .Y(new_n4469_));
  NAND2X1  g03467(.A(new_n4419_), .B(new_n4396_), .Y(new_n4470_));
  OAI22X1  g03468(.A0(new_n4410_), .A1(new_n4414_), .B0(new_n4418_), .B1(new_n4383_), .Y(new_n4471_));
  AOI22X1  g03469(.A0(new_n4471_), .A1(new_n4454_), .B0(new_n4456_), .B1(new_n4470_), .Y(new_n4472_));
  AOI21X1  g03470(.A0(new_n4461_), .A1(new_n4472_), .B0(new_n4448_), .Y(new_n4473_));
  AOI22X1  g03471(.A0(new_n4473_), .A1(new_n4469_), .B0(new_n4462_), .B1(new_n4448_), .Y(new_n4474_));
  OAI22X1  g03472(.A0(new_n4474_), .A1(new_n4464_), .B0(new_n4468_), .B1(new_n4463_), .Y(new_n4475_));
  NAND2X1  g03473(.A(new_n4421_), .B(new_n4382_), .Y(new_n4476_));
  OAI21X1  g03474(.A0(new_n4467_), .A1(new_n4466_), .B0(new_n4476_), .Y(new_n4477_));
  OAI22X1  g03475(.A0(new_n4477_), .A1(new_n4463_), .B0(new_n4474_), .B1(new_n4476_), .Y(new_n4478_));
  MX2X1    g03476(.A(new_n4478_), .B(new_n4475_), .S0(new_n4445_), .Y(new_n4479_));
  AND2X1   g03477(.A(new_n4422_), .B(new_n4364_), .Y(new_n4480_));
  AOI21X1  g03478(.A0(new_n4431_), .A1(new_n4269_), .B0(new_n4480_), .Y(new_n4481_));
  AOI22X1  g03479(.A0(new_n4481_), .A1(new_n4363_), .B0(new_n4436_), .B1(new_n4480_), .Y(new_n4482_));
  MX2X1    g03480(.A(new_n4437_), .B(new_n4482_), .S0(new_n4479_), .Y(new_n4483_));
  INVX1    g03481(.A(\A[45] ), .Y(new_n4484_));
  INVX1    g03482(.A(\A[44] ), .Y(new_n4485_));
  OR2X1    g03483(.A(new_n4485_), .B(\A[43] ), .Y(new_n4486_));
  AOI21X1  g03484(.A0(new_n4485_), .A1(\A[43] ), .B0(new_n4484_), .Y(new_n4487_));
  XOR2X1   g03485(.A(\A[44] ), .B(\A[43] ), .Y(new_n4488_));
  AOI22X1  g03486(.A0(new_n4488_), .A1(new_n4484_), .B0(new_n4487_), .B1(new_n4486_), .Y(new_n4489_));
  INVX1    g03487(.A(\A[48] ), .Y(new_n4490_));
  INVX1    g03488(.A(\A[47] ), .Y(new_n4491_));
  OR2X1    g03489(.A(new_n4491_), .B(\A[46] ), .Y(new_n4492_));
  AOI21X1  g03490(.A0(new_n4491_), .A1(\A[46] ), .B0(new_n4490_), .Y(new_n4493_));
  XOR2X1   g03491(.A(\A[47] ), .B(\A[46] ), .Y(new_n4494_));
  AOI22X1  g03492(.A0(new_n4494_), .A1(new_n4490_), .B0(new_n4493_), .B1(new_n4492_), .Y(new_n4495_));
  OR2X1    g03493(.A(new_n4495_), .B(new_n4489_), .Y(new_n4496_));
  AND2X1   g03494(.A(\A[47] ), .B(\A[46] ), .Y(new_n4497_));
  AND2X1   g03495(.A(new_n4494_), .B(\A[48] ), .Y(new_n4498_));
  OR2X1    g03496(.A(new_n4498_), .B(new_n4497_), .Y(new_n4499_));
  AND2X1   g03497(.A(\A[44] ), .B(\A[43] ), .Y(new_n4500_));
  AOI21X1  g03498(.A0(new_n4488_), .A1(\A[45] ), .B0(new_n4500_), .Y(new_n4501_));
  XOR2X1   g03499(.A(new_n4501_), .B(new_n4499_), .Y(new_n4502_));
  XOR2X1   g03500(.A(new_n4502_), .B(new_n4496_), .Y(new_n4503_));
  INVX1    g03501(.A(\A[43] ), .Y(new_n4504_));
  AND2X1   g03502(.A(\A[44] ), .B(new_n4504_), .Y(new_n4505_));
  OAI21X1  g03503(.A0(\A[44] ), .A1(new_n4504_), .B0(\A[45] ), .Y(new_n4506_));
  NAND2X1  g03504(.A(new_n4488_), .B(new_n4484_), .Y(new_n4507_));
  OAI21X1  g03505(.A0(new_n4506_), .A1(new_n4505_), .B0(new_n4507_), .Y(new_n4508_));
  XOR2X1   g03506(.A(new_n4495_), .B(new_n4508_), .Y(new_n4509_));
  NOR2X1   g03507(.A(new_n4495_), .B(new_n4489_), .Y(new_n4510_));
  AOI21X1  g03508(.A0(new_n4494_), .A1(\A[48] ), .B0(new_n4497_), .Y(new_n4511_));
  XOR2X1   g03509(.A(new_n4501_), .B(new_n4511_), .Y(new_n4512_));
  NOR2X1   g03510(.A(new_n4501_), .B(new_n4511_), .Y(new_n4513_));
  AOI21X1  g03511(.A0(new_n4512_), .A1(new_n4510_), .B0(new_n4513_), .Y(new_n4514_));
  OAI21X1  g03512(.A0(new_n4514_), .A1(new_n4509_), .B0(new_n4503_), .Y(new_n4515_));
  AND2X1   g03513(.A(\A[53] ), .B(\A[52] ), .Y(new_n4516_));
  XOR2X1   g03514(.A(\A[53] ), .B(\A[52] ), .Y(new_n4517_));
  AOI21X1  g03515(.A0(new_n4517_), .A1(\A[54] ), .B0(new_n4516_), .Y(new_n4518_));
  AND2X1   g03516(.A(\A[50] ), .B(\A[49] ), .Y(new_n4519_));
  XOR2X1   g03517(.A(\A[50] ), .B(\A[49] ), .Y(new_n4520_));
  AOI21X1  g03518(.A0(new_n4520_), .A1(\A[51] ), .B0(new_n4519_), .Y(new_n4521_));
  INVX1    g03519(.A(\A[51] ), .Y(new_n4522_));
  INVX1    g03520(.A(\A[50] ), .Y(new_n4523_));
  OR2X1    g03521(.A(new_n4523_), .B(\A[49] ), .Y(new_n4524_));
  AOI21X1  g03522(.A0(new_n4523_), .A1(\A[49] ), .B0(new_n4522_), .Y(new_n4525_));
  AOI22X1  g03523(.A0(new_n4525_), .A1(new_n4524_), .B0(new_n4520_), .B1(new_n4522_), .Y(new_n4526_));
  INVX1    g03524(.A(\A[54] ), .Y(new_n4527_));
  INVX1    g03525(.A(\A[53] ), .Y(new_n4528_));
  OR2X1    g03526(.A(new_n4528_), .B(\A[52] ), .Y(new_n4529_));
  AOI21X1  g03527(.A0(new_n4528_), .A1(\A[52] ), .B0(new_n4527_), .Y(new_n4530_));
  AOI22X1  g03528(.A0(new_n4530_), .A1(new_n4529_), .B0(new_n4517_), .B1(new_n4527_), .Y(new_n4531_));
  NOR4X1   g03529(.A(new_n4531_), .B(new_n4526_), .C(new_n4521_), .D(new_n4518_), .Y(new_n4532_));
  NOR4X1   g03530(.A(new_n4501_), .B(new_n4511_), .C(new_n4495_), .D(new_n4489_), .Y(new_n4533_));
  INVX1    g03531(.A(\A[49] ), .Y(new_n4534_));
  AND2X1   g03532(.A(\A[50] ), .B(new_n4534_), .Y(new_n4535_));
  OAI21X1  g03533(.A0(\A[50] ), .A1(new_n4534_), .B0(\A[51] ), .Y(new_n4536_));
  NAND2X1  g03534(.A(new_n4520_), .B(new_n4522_), .Y(new_n4537_));
  OAI21X1  g03535(.A0(new_n4536_), .A1(new_n4535_), .B0(new_n4537_), .Y(new_n4538_));
  XOR2X1   g03536(.A(new_n4531_), .B(new_n4538_), .Y(new_n4539_));
  OR4X1    g03537(.A(new_n4539_), .B(new_n4533_), .C(new_n4532_), .D(new_n4509_), .Y(new_n4540_));
  XOR2X1   g03538(.A(new_n4521_), .B(new_n4518_), .Y(new_n4541_));
  NOR2X1   g03539(.A(new_n4531_), .B(new_n4526_), .Y(new_n4542_));
  NOR2X1   g03540(.A(new_n4521_), .B(new_n4518_), .Y(new_n4543_));
  AOI21X1  g03541(.A0(new_n4542_), .A1(new_n4541_), .B0(new_n4543_), .Y(new_n4544_));
  XOR2X1   g03542(.A(new_n4542_), .B(new_n4541_), .Y(new_n4545_));
  OAI21X1  g03543(.A0(new_n4539_), .A1(new_n4544_), .B0(new_n4545_), .Y(new_n4546_));
  XOR2X1   g03544(.A(new_n4546_), .B(new_n4540_), .Y(new_n4547_));
  NAND2X1  g03545(.A(new_n4547_), .B(new_n4515_), .Y(new_n4548_));
  XOR2X1   g03546(.A(new_n4495_), .B(new_n4489_), .Y(new_n4549_));
  OAI21X1  g03547(.A0(new_n4539_), .A1(new_n4532_), .B0(new_n4549_), .Y(new_n4550_));
  OR4X1    g03548(.A(new_n4531_), .B(new_n4526_), .C(new_n4521_), .D(new_n4518_), .Y(new_n4551_));
  XOR2X1   g03549(.A(new_n4531_), .B(new_n4526_), .Y(new_n4552_));
  XOR2X1   g03550(.A(new_n4495_), .B(new_n4508_), .Y(new_n4553_));
  NAND3X1  g03551(.A(new_n4553_), .B(new_n4552_), .C(new_n4551_), .Y(new_n4554_));
  AND2X1   g03552(.A(new_n4554_), .B(new_n4550_), .Y(new_n4555_));
  INVX1    g03553(.A(\A[38] ), .Y(new_n4556_));
  AND2X1   g03554(.A(new_n4556_), .B(\A[37] ), .Y(new_n4557_));
  OAI21X1  g03555(.A0(new_n4556_), .A1(\A[37] ), .B0(\A[39] ), .Y(new_n4558_));
  INVX1    g03556(.A(\A[39] ), .Y(new_n4559_));
  XOR2X1   g03557(.A(\A[38] ), .B(\A[37] ), .Y(new_n4560_));
  NAND2X1  g03558(.A(new_n4560_), .B(new_n4559_), .Y(new_n4561_));
  OAI21X1  g03559(.A0(new_n4558_), .A1(new_n4557_), .B0(new_n4561_), .Y(new_n4562_));
  INVX1    g03560(.A(\A[42] ), .Y(new_n4563_));
  INVX1    g03561(.A(\A[40] ), .Y(new_n4564_));
  OR2X1    g03562(.A(\A[41] ), .B(new_n4564_), .Y(new_n4565_));
  AOI21X1  g03563(.A0(\A[41] ), .A1(new_n4564_), .B0(new_n4563_), .Y(new_n4566_));
  XOR2X1   g03564(.A(\A[41] ), .B(\A[40] ), .Y(new_n4567_));
  AOI22X1  g03565(.A0(new_n4567_), .A1(new_n4563_), .B0(new_n4566_), .B1(new_n4565_), .Y(new_n4568_));
  AND2X1   g03566(.A(\A[41] ), .B(\A[40] ), .Y(new_n4569_));
  AOI21X1  g03567(.A0(new_n4567_), .A1(\A[42] ), .B0(new_n4569_), .Y(new_n4570_));
  AND2X1   g03568(.A(\A[38] ), .B(\A[37] ), .Y(new_n4571_));
  AOI21X1  g03569(.A0(new_n4560_), .A1(\A[39] ), .B0(new_n4571_), .Y(new_n4572_));
  XOR2X1   g03570(.A(new_n4568_), .B(new_n4562_), .Y(new_n4573_));
  INVX1    g03571(.A(\A[33] ), .Y(new_n4574_));
  INVX1    g03572(.A(\A[31] ), .Y(new_n4575_));
  OR2X1    g03573(.A(\A[32] ), .B(new_n4575_), .Y(new_n4576_));
  AOI21X1  g03574(.A0(\A[32] ), .A1(new_n4575_), .B0(new_n4574_), .Y(new_n4577_));
  XOR2X1   g03575(.A(\A[32] ), .B(\A[31] ), .Y(new_n4578_));
  AOI22X1  g03576(.A0(new_n4578_), .A1(new_n4574_), .B0(new_n4577_), .B1(new_n4576_), .Y(new_n4579_));
  INVX1    g03577(.A(\A[36] ), .Y(new_n4580_));
  INVX1    g03578(.A(\A[34] ), .Y(new_n4581_));
  OR2X1    g03579(.A(\A[35] ), .B(new_n4581_), .Y(new_n4582_));
  AOI21X1  g03580(.A0(\A[35] ), .A1(new_n4581_), .B0(new_n4580_), .Y(new_n4583_));
  XOR2X1   g03581(.A(\A[35] ), .B(\A[34] ), .Y(new_n4584_));
  AOI22X1  g03582(.A0(new_n4584_), .A1(new_n4580_), .B0(new_n4583_), .B1(new_n4582_), .Y(new_n4585_));
  AND2X1   g03583(.A(\A[35] ), .B(\A[34] ), .Y(new_n4586_));
  AOI21X1  g03584(.A0(new_n4584_), .A1(\A[36] ), .B0(new_n4586_), .Y(new_n4587_));
  AND2X1   g03585(.A(\A[32] ), .B(\A[31] ), .Y(new_n4588_));
  AOI21X1  g03586(.A0(new_n4578_), .A1(\A[33] ), .B0(new_n4588_), .Y(new_n4589_));
  XOR2X1   g03587(.A(new_n4585_), .B(new_n4579_), .Y(new_n4590_));
  XOR2X1   g03588(.A(new_n4590_), .B(new_n4573_), .Y(new_n4591_));
  OR2X1    g03589(.A(new_n4591_), .B(new_n4555_), .Y(new_n4592_));
  XOR2X1   g03590(.A(new_n4502_), .B(new_n4510_), .Y(new_n4593_));
  XOR2X1   g03591(.A(new_n4495_), .B(new_n4489_), .Y(new_n4594_));
  OR2X1    g03592(.A(new_n4501_), .B(new_n4511_), .Y(new_n4595_));
  OAI21X1  g03593(.A0(new_n4502_), .A1(new_n4496_), .B0(new_n4595_), .Y(new_n4596_));
  AOI21X1  g03594(.A0(new_n4596_), .A1(new_n4594_), .B0(new_n4593_), .Y(new_n4597_));
  NOR4X1   g03595(.A(new_n4539_), .B(new_n4533_), .C(new_n4532_), .D(new_n4509_), .Y(new_n4598_));
  AND2X1   g03596(.A(new_n4517_), .B(\A[54] ), .Y(new_n4599_));
  OR2X1    g03597(.A(new_n4599_), .B(new_n4516_), .Y(new_n4600_));
  XOR2X1   g03598(.A(new_n4521_), .B(new_n4600_), .Y(new_n4601_));
  OR2X1    g03599(.A(new_n4531_), .B(new_n4526_), .Y(new_n4602_));
  OR2X1    g03600(.A(new_n4521_), .B(new_n4518_), .Y(new_n4603_));
  OAI21X1  g03601(.A0(new_n4602_), .A1(new_n4601_), .B0(new_n4603_), .Y(new_n4604_));
  XOR2X1   g03602(.A(new_n4542_), .B(new_n4601_), .Y(new_n4605_));
  AOI21X1  g03603(.A0(new_n4552_), .A1(new_n4604_), .B0(new_n4605_), .Y(new_n4606_));
  OR4X1    g03604(.A(new_n4539_), .B(new_n4533_), .C(new_n4605_), .D(new_n4509_), .Y(new_n4607_));
  AOI21X1  g03605(.A0(new_n4539_), .A1(new_n4605_), .B0(new_n4544_), .Y(new_n4608_));
  OAI22X1  g03606(.A0(new_n4608_), .A1(new_n4607_), .B0(new_n4606_), .B1(new_n4598_), .Y(new_n4609_));
  AOI21X1  g03607(.A0(new_n4609_), .A1(new_n4597_), .B0(new_n4592_), .Y(new_n4610_));
  MX2X1    g03608(.A(new_n4609_), .B(new_n4547_), .S0(new_n4515_), .Y(new_n4611_));
  AOI22X1  g03609(.A0(new_n4611_), .A1(new_n4592_), .B0(new_n4610_), .B1(new_n4548_), .Y(new_n4612_));
  INVX1    g03610(.A(\A[32] ), .Y(new_n4613_));
  AND2X1   g03611(.A(new_n4613_), .B(\A[31] ), .Y(new_n4614_));
  OAI21X1  g03612(.A0(new_n4613_), .A1(\A[31] ), .B0(\A[33] ), .Y(new_n4615_));
  NAND2X1  g03613(.A(new_n4578_), .B(new_n4574_), .Y(new_n4616_));
  OAI21X1  g03614(.A0(new_n4615_), .A1(new_n4614_), .B0(new_n4616_), .Y(new_n4617_));
  XOR2X1   g03615(.A(new_n4585_), .B(new_n4617_), .Y(new_n4618_));
  XOR2X1   g03616(.A(new_n4589_), .B(new_n4587_), .Y(new_n4619_));
  NOR2X1   g03617(.A(new_n4585_), .B(new_n4579_), .Y(new_n4620_));
  NOR2X1   g03618(.A(new_n4589_), .B(new_n4587_), .Y(new_n4621_));
  AOI21X1  g03619(.A0(new_n4620_), .A1(new_n4619_), .B0(new_n4621_), .Y(new_n4622_));
  XOR2X1   g03620(.A(new_n4620_), .B(new_n4619_), .Y(new_n4623_));
  OAI21X1  g03621(.A0(new_n4622_), .A1(new_n4618_), .B0(new_n4623_), .Y(new_n4624_));
  XOR2X1   g03622(.A(new_n4568_), .B(new_n4562_), .Y(new_n4625_));
  INVX1    g03623(.A(\A[37] ), .Y(new_n4626_));
  OR2X1    g03624(.A(\A[38] ), .B(new_n4626_), .Y(new_n4627_));
  AOI21X1  g03625(.A0(\A[38] ), .A1(new_n4626_), .B0(new_n4559_), .Y(new_n4628_));
  AOI22X1  g03626(.A0(new_n4560_), .A1(new_n4559_), .B0(new_n4628_), .B1(new_n4627_), .Y(new_n4629_));
  NOR4X1   g03627(.A(new_n4572_), .B(new_n4570_), .C(new_n4568_), .D(new_n4629_), .Y(new_n4630_));
  NOR4X1   g03628(.A(new_n4589_), .B(new_n4587_), .C(new_n4585_), .D(new_n4579_), .Y(new_n4631_));
  OR4X1    g03629(.A(new_n4631_), .B(new_n4618_), .C(new_n4630_), .D(new_n4625_), .Y(new_n4632_));
  XOR2X1   g03630(.A(new_n4568_), .B(new_n4629_), .Y(new_n4633_));
  AND2X1   g03631(.A(new_n4567_), .B(\A[42] ), .Y(new_n4634_));
  OR2X1    g03632(.A(new_n4634_), .B(new_n4569_), .Y(new_n4635_));
  XOR2X1   g03633(.A(new_n4572_), .B(new_n4635_), .Y(new_n4636_));
  OR2X1    g03634(.A(new_n4568_), .B(new_n4629_), .Y(new_n4637_));
  OR2X1    g03635(.A(new_n4572_), .B(new_n4570_), .Y(new_n4638_));
  OAI21X1  g03636(.A0(new_n4637_), .A1(new_n4636_), .B0(new_n4638_), .Y(new_n4639_));
  NOR2X1   g03637(.A(new_n4568_), .B(new_n4629_), .Y(new_n4640_));
  XOR2X1   g03638(.A(new_n4640_), .B(new_n4636_), .Y(new_n4641_));
  AOI21X1  g03639(.A0(new_n4639_), .A1(new_n4633_), .B0(new_n4641_), .Y(new_n4642_));
  XOR2X1   g03640(.A(new_n4642_), .B(new_n4632_), .Y(new_n4643_));
  XOR2X1   g03641(.A(new_n4572_), .B(new_n4570_), .Y(new_n4644_));
  NOR2X1   g03642(.A(new_n4572_), .B(new_n4570_), .Y(new_n4645_));
  AOI21X1  g03643(.A0(new_n4640_), .A1(new_n4644_), .B0(new_n4645_), .Y(new_n4646_));
  XOR2X1   g03644(.A(new_n4640_), .B(new_n4644_), .Y(new_n4647_));
  OAI21X1  g03645(.A0(new_n4646_), .A1(new_n4625_), .B0(new_n4647_), .Y(new_n4648_));
  NOR4X1   g03646(.A(new_n4618_), .B(new_n4641_), .C(new_n4639_), .D(new_n4625_), .Y(new_n4649_));
  AOI21X1  g03647(.A0(new_n4639_), .A1(new_n4633_), .B0(new_n4631_), .Y(new_n4650_));
  AOI22X1  g03648(.A0(new_n4650_), .A1(new_n4649_), .B0(new_n4648_), .B1(new_n4632_), .Y(new_n4651_));
  MX2X1    g03649(.A(new_n4651_), .B(new_n4643_), .S0(new_n4624_), .Y(new_n4652_));
  AOI21X1  g03650(.A0(new_n4554_), .A1(new_n4550_), .B0(new_n4591_), .Y(new_n4653_));
  AOI21X1  g03651(.A0(new_n4609_), .A1(new_n4597_), .B0(new_n4653_), .Y(new_n4654_));
  AOI22X1  g03652(.A0(new_n4654_), .A1(new_n4548_), .B0(new_n4611_), .B1(new_n4653_), .Y(new_n4655_));
  MX2X1    g03653(.A(new_n4655_), .B(new_n4612_), .S0(new_n4652_), .Y(new_n4656_));
  INVX1    g03654(.A(\A[57] ), .Y(new_n4657_));
  INVX1    g03655(.A(\A[56] ), .Y(new_n4658_));
  OR2X1    g03656(.A(new_n4658_), .B(\A[55] ), .Y(new_n4659_));
  AOI21X1  g03657(.A0(new_n4658_), .A1(\A[55] ), .B0(new_n4657_), .Y(new_n4660_));
  XOR2X1   g03658(.A(\A[56] ), .B(\A[55] ), .Y(new_n4661_));
  AOI22X1  g03659(.A0(new_n4661_), .A1(new_n4657_), .B0(new_n4660_), .B1(new_n4659_), .Y(new_n4662_));
  INVX1    g03660(.A(\A[60] ), .Y(new_n4663_));
  INVX1    g03661(.A(\A[59] ), .Y(new_n4664_));
  OR2X1    g03662(.A(new_n4664_), .B(\A[58] ), .Y(new_n4665_));
  AOI21X1  g03663(.A0(new_n4664_), .A1(\A[58] ), .B0(new_n4663_), .Y(new_n4666_));
  XOR2X1   g03664(.A(\A[59] ), .B(\A[58] ), .Y(new_n4667_));
  AOI22X1  g03665(.A0(new_n4667_), .A1(new_n4663_), .B0(new_n4666_), .B1(new_n4665_), .Y(new_n4668_));
  OR2X1    g03666(.A(new_n4668_), .B(new_n4662_), .Y(new_n4669_));
  AND2X1   g03667(.A(\A[59] ), .B(\A[58] ), .Y(new_n4670_));
  AND2X1   g03668(.A(new_n4667_), .B(\A[60] ), .Y(new_n4671_));
  OR2X1    g03669(.A(new_n4671_), .B(new_n4670_), .Y(new_n4672_));
  AND2X1   g03670(.A(\A[56] ), .B(\A[55] ), .Y(new_n4673_));
  AOI21X1  g03671(.A0(new_n4661_), .A1(\A[57] ), .B0(new_n4673_), .Y(new_n4674_));
  XOR2X1   g03672(.A(new_n4674_), .B(new_n4672_), .Y(new_n4675_));
  XOR2X1   g03673(.A(new_n4675_), .B(new_n4669_), .Y(new_n4676_));
  INVX1    g03674(.A(\A[55] ), .Y(new_n4677_));
  AND2X1   g03675(.A(\A[56] ), .B(new_n4677_), .Y(new_n4678_));
  OAI21X1  g03676(.A0(\A[56] ), .A1(new_n4677_), .B0(\A[57] ), .Y(new_n4679_));
  NAND2X1  g03677(.A(new_n4661_), .B(new_n4657_), .Y(new_n4680_));
  OAI21X1  g03678(.A0(new_n4679_), .A1(new_n4678_), .B0(new_n4680_), .Y(new_n4681_));
  XOR2X1   g03679(.A(new_n4668_), .B(new_n4681_), .Y(new_n4682_));
  NOR2X1   g03680(.A(new_n4668_), .B(new_n4662_), .Y(new_n4683_));
  AOI21X1  g03681(.A0(new_n4667_), .A1(\A[60] ), .B0(new_n4670_), .Y(new_n4684_));
  XOR2X1   g03682(.A(new_n4674_), .B(new_n4684_), .Y(new_n4685_));
  NOR2X1   g03683(.A(new_n4674_), .B(new_n4684_), .Y(new_n4686_));
  AOI21X1  g03684(.A0(new_n4685_), .A1(new_n4683_), .B0(new_n4686_), .Y(new_n4687_));
  OAI21X1  g03685(.A0(new_n4687_), .A1(new_n4682_), .B0(new_n4676_), .Y(new_n4688_));
  AND2X1   g03686(.A(\A[65] ), .B(\A[64] ), .Y(new_n4689_));
  XOR2X1   g03687(.A(\A[65] ), .B(\A[64] ), .Y(new_n4690_));
  AOI21X1  g03688(.A0(new_n4690_), .A1(\A[66] ), .B0(new_n4689_), .Y(new_n4691_));
  AND2X1   g03689(.A(\A[62] ), .B(\A[61] ), .Y(new_n4692_));
  XOR2X1   g03690(.A(\A[62] ), .B(\A[61] ), .Y(new_n4693_));
  AOI21X1  g03691(.A0(new_n4693_), .A1(\A[63] ), .B0(new_n4692_), .Y(new_n4694_));
  INVX1    g03692(.A(\A[63] ), .Y(new_n4695_));
  INVX1    g03693(.A(\A[62] ), .Y(new_n4696_));
  OR2X1    g03694(.A(new_n4696_), .B(\A[61] ), .Y(new_n4697_));
  AOI21X1  g03695(.A0(new_n4696_), .A1(\A[61] ), .B0(new_n4695_), .Y(new_n4698_));
  AOI22X1  g03696(.A0(new_n4698_), .A1(new_n4697_), .B0(new_n4693_), .B1(new_n4695_), .Y(new_n4699_));
  INVX1    g03697(.A(\A[66] ), .Y(new_n4700_));
  INVX1    g03698(.A(\A[65] ), .Y(new_n4701_));
  OR2X1    g03699(.A(new_n4701_), .B(\A[64] ), .Y(new_n4702_));
  AOI21X1  g03700(.A0(new_n4701_), .A1(\A[64] ), .B0(new_n4700_), .Y(new_n4703_));
  AOI22X1  g03701(.A0(new_n4703_), .A1(new_n4702_), .B0(new_n4690_), .B1(new_n4700_), .Y(new_n4704_));
  NOR4X1   g03702(.A(new_n4704_), .B(new_n4699_), .C(new_n4694_), .D(new_n4691_), .Y(new_n4705_));
  NOR4X1   g03703(.A(new_n4674_), .B(new_n4684_), .C(new_n4668_), .D(new_n4662_), .Y(new_n4706_));
  INVX1    g03704(.A(\A[61] ), .Y(new_n4707_));
  AND2X1   g03705(.A(\A[62] ), .B(new_n4707_), .Y(new_n4708_));
  OAI21X1  g03706(.A0(\A[62] ), .A1(new_n4707_), .B0(\A[63] ), .Y(new_n4709_));
  NAND2X1  g03707(.A(new_n4693_), .B(new_n4695_), .Y(new_n4710_));
  OAI21X1  g03708(.A0(new_n4709_), .A1(new_n4708_), .B0(new_n4710_), .Y(new_n4711_));
  XOR2X1   g03709(.A(new_n4704_), .B(new_n4711_), .Y(new_n4712_));
  OR4X1    g03710(.A(new_n4712_), .B(new_n4706_), .C(new_n4705_), .D(new_n4682_), .Y(new_n4713_));
  AND2X1   g03711(.A(new_n4690_), .B(\A[66] ), .Y(new_n4714_));
  OR2X1    g03712(.A(new_n4714_), .B(new_n4689_), .Y(new_n4715_));
  XOR2X1   g03713(.A(new_n4694_), .B(new_n4715_), .Y(new_n4716_));
  OR2X1    g03714(.A(new_n4704_), .B(new_n4699_), .Y(new_n4717_));
  OR2X1    g03715(.A(new_n4694_), .B(new_n4691_), .Y(new_n4718_));
  OAI21X1  g03716(.A0(new_n4717_), .A1(new_n4716_), .B0(new_n4718_), .Y(new_n4719_));
  NOR2X1   g03717(.A(new_n4704_), .B(new_n4699_), .Y(new_n4720_));
  XOR2X1   g03718(.A(new_n4720_), .B(new_n4716_), .Y(new_n4721_));
  XOR2X1   g03719(.A(new_n4704_), .B(new_n4699_), .Y(new_n4722_));
  AOI21X1  g03720(.A0(new_n4722_), .A1(new_n4719_), .B0(new_n4721_), .Y(new_n4723_));
  XOR2X1   g03721(.A(new_n4723_), .B(new_n4713_), .Y(new_n4724_));
  XOR2X1   g03722(.A(new_n4694_), .B(new_n4691_), .Y(new_n4725_));
  NOR2X1   g03723(.A(new_n4694_), .B(new_n4691_), .Y(new_n4726_));
  AOI21X1  g03724(.A0(new_n4720_), .A1(new_n4725_), .B0(new_n4726_), .Y(new_n4727_));
  XOR2X1   g03725(.A(new_n4720_), .B(new_n4725_), .Y(new_n4728_));
  OAI21X1  g03726(.A0(new_n4712_), .A1(new_n4727_), .B0(new_n4728_), .Y(new_n4729_));
  NOR4X1   g03727(.A(new_n4712_), .B(new_n4706_), .C(new_n4721_), .D(new_n4682_), .Y(new_n4730_));
  OAI21X1  g03728(.A0(new_n4722_), .A1(new_n4728_), .B0(new_n4719_), .Y(new_n4731_));
  AOI22X1  g03729(.A0(new_n4731_), .A1(new_n4730_), .B0(new_n4729_), .B1(new_n4713_), .Y(new_n4732_));
  MX2X1    g03730(.A(new_n4732_), .B(new_n4724_), .S0(new_n4688_), .Y(new_n4733_));
  INVX1    g03731(.A(\A[69] ), .Y(new_n4734_));
  INVX1    g03732(.A(\A[68] ), .Y(new_n4735_));
  OR2X1    g03733(.A(new_n4735_), .B(\A[67] ), .Y(new_n4736_));
  AOI21X1  g03734(.A0(new_n4735_), .A1(\A[67] ), .B0(new_n4734_), .Y(new_n4737_));
  XOR2X1   g03735(.A(\A[68] ), .B(\A[67] ), .Y(new_n4738_));
  AOI22X1  g03736(.A0(new_n4738_), .A1(new_n4734_), .B0(new_n4737_), .B1(new_n4736_), .Y(new_n4739_));
  INVX1    g03737(.A(\A[72] ), .Y(new_n4740_));
  INVX1    g03738(.A(\A[71] ), .Y(new_n4741_));
  OR2X1    g03739(.A(new_n4741_), .B(\A[70] ), .Y(new_n4742_));
  AOI21X1  g03740(.A0(new_n4741_), .A1(\A[70] ), .B0(new_n4740_), .Y(new_n4743_));
  XOR2X1   g03741(.A(\A[71] ), .B(\A[70] ), .Y(new_n4744_));
  AOI22X1  g03742(.A0(new_n4744_), .A1(new_n4740_), .B0(new_n4743_), .B1(new_n4742_), .Y(new_n4745_));
  OR2X1    g03743(.A(new_n4745_), .B(new_n4739_), .Y(new_n4746_));
  AND2X1   g03744(.A(\A[71] ), .B(\A[70] ), .Y(new_n4747_));
  AND2X1   g03745(.A(new_n4744_), .B(\A[72] ), .Y(new_n4748_));
  OR2X1    g03746(.A(new_n4748_), .B(new_n4747_), .Y(new_n4749_));
  AND2X1   g03747(.A(\A[68] ), .B(\A[67] ), .Y(new_n4750_));
  AOI21X1  g03748(.A0(new_n4738_), .A1(\A[69] ), .B0(new_n4750_), .Y(new_n4751_));
  XOR2X1   g03749(.A(new_n4751_), .B(new_n4749_), .Y(new_n4752_));
  XOR2X1   g03750(.A(new_n4752_), .B(new_n4746_), .Y(new_n4753_));
  INVX1    g03751(.A(\A[67] ), .Y(new_n4754_));
  AND2X1   g03752(.A(\A[68] ), .B(new_n4754_), .Y(new_n4755_));
  OAI21X1  g03753(.A0(\A[68] ), .A1(new_n4754_), .B0(\A[69] ), .Y(new_n4756_));
  NAND2X1  g03754(.A(new_n4738_), .B(new_n4734_), .Y(new_n4757_));
  OAI21X1  g03755(.A0(new_n4756_), .A1(new_n4755_), .B0(new_n4757_), .Y(new_n4758_));
  XOR2X1   g03756(.A(new_n4745_), .B(new_n4758_), .Y(new_n4759_));
  NOR2X1   g03757(.A(new_n4745_), .B(new_n4739_), .Y(new_n4760_));
  AOI21X1  g03758(.A0(new_n4744_), .A1(\A[72] ), .B0(new_n4747_), .Y(new_n4761_));
  XOR2X1   g03759(.A(new_n4751_), .B(new_n4761_), .Y(new_n4762_));
  NOR2X1   g03760(.A(new_n4751_), .B(new_n4761_), .Y(new_n4763_));
  AOI21X1  g03761(.A0(new_n4762_), .A1(new_n4760_), .B0(new_n4763_), .Y(new_n4764_));
  OAI21X1  g03762(.A0(new_n4764_), .A1(new_n4759_), .B0(new_n4753_), .Y(new_n4765_));
  AND2X1   g03763(.A(\A[77] ), .B(\A[76] ), .Y(new_n4766_));
  XOR2X1   g03764(.A(\A[77] ), .B(\A[76] ), .Y(new_n4767_));
  AOI21X1  g03765(.A0(new_n4767_), .A1(\A[78] ), .B0(new_n4766_), .Y(new_n4768_));
  AND2X1   g03766(.A(\A[74] ), .B(\A[73] ), .Y(new_n4769_));
  XOR2X1   g03767(.A(\A[74] ), .B(\A[73] ), .Y(new_n4770_));
  AOI21X1  g03768(.A0(new_n4770_), .A1(\A[75] ), .B0(new_n4769_), .Y(new_n4771_));
  INVX1    g03769(.A(\A[75] ), .Y(new_n4772_));
  INVX1    g03770(.A(\A[74] ), .Y(new_n4773_));
  OR2X1    g03771(.A(new_n4773_), .B(\A[73] ), .Y(new_n4774_));
  AOI21X1  g03772(.A0(new_n4773_), .A1(\A[73] ), .B0(new_n4772_), .Y(new_n4775_));
  AOI22X1  g03773(.A0(new_n4775_), .A1(new_n4774_), .B0(new_n4770_), .B1(new_n4772_), .Y(new_n4776_));
  INVX1    g03774(.A(\A[78] ), .Y(new_n4777_));
  INVX1    g03775(.A(\A[77] ), .Y(new_n4778_));
  OR2X1    g03776(.A(new_n4778_), .B(\A[76] ), .Y(new_n4779_));
  AOI21X1  g03777(.A0(new_n4778_), .A1(\A[76] ), .B0(new_n4777_), .Y(new_n4780_));
  AOI22X1  g03778(.A0(new_n4780_), .A1(new_n4779_), .B0(new_n4767_), .B1(new_n4777_), .Y(new_n4781_));
  NOR4X1   g03779(.A(new_n4781_), .B(new_n4776_), .C(new_n4771_), .D(new_n4768_), .Y(new_n4782_));
  NOR4X1   g03780(.A(new_n4751_), .B(new_n4761_), .C(new_n4745_), .D(new_n4739_), .Y(new_n4783_));
  INVX1    g03781(.A(\A[73] ), .Y(new_n4784_));
  AND2X1   g03782(.A(\A[74] ), .B(new_n4784_), .Y(new_n4785_));
  OAI21X1  g03783(.A0(\A[74] ), .A1(new_n4784_), .B0(\A[75] ), .Y(new_n4786_));
  NAND2X1  g03784(.A(new_n4770_), .B(new_n4772_), .Y(new_n4787_));
  OAI21X1  g03785(.A0(new_n4786_), .A1(new_n4785_), .B0(new_n4787_), .Y(new_n4788_));
  XOR2X1   g03786(.A(new_n4781_), .B(new_n4788_), .Y(new_n4789_));
  OR4X1    g03787(.A(new_n4789_), .B(new_n4783_), .C(new_n4782_), .D(new_n4759_), .Y(new_n4790_));
  XOR2X1   g03788(.A(new_n4771_), .B(new_n4768_), .Y(new_n4791_));
  NOR2X1   g03789(.A(new_n4781_), .B(new_n4776_), .Y(new_n4792_));
  NOR2X1   g03790(.A(new_n4771_), .B(new_n4768_), .Y(new_n4793_));
  AOI21X1  g03791(.A0(new_n4792_), .A1(new_n4791_), .B0(new_n4793_), .Y(new_n4794_));
  XOR2X1   g03792(.A(new_n4792_), .B(new_n4791_), .Y(new_n4795_));
  OAI21X1  g03793(.A0(new_n4789_), .A1(new_n4794_), .B0(new_n4795_), .Y(new_n4796_));
  XOR2X1   g03794(.A(new_n4796_), .B(new_n4790_), .Y(new_n4797_));
  AND2X1   g03795(.A(new_n4797_), .B(new_n4765_), .Y(new_n4798_));
  OR2X1    g03796(.A(new_n4789_), .B(new_n4782_), .Y(new_n4799_));
  XOR2X1   g03797(.A(new_n4745_), .B(new_n4739_), .Y(new_n4800_));
  XOR2X1   g03798(.A(new_n4800_), .B(new_n4799_), .Y(new_n4801_));
  OR2X1    g03799(.A(new_n4712_), .B(new_n4705_), .Y(new_n4802_));
  XOR2X1   g03800(.A(new_n4668_), .B(new_n4662_), .Y(new_n4803_));
  XOR2X1   g03801(.A(new_n4803_), .B(new_n4802_), .Y(new_n4804_));
  NOR2X1   g03802(.A(new_n4804_), .B(new_n4801_), .Y(new_n4805_));
  AND2X1   g03803(.A(new_n4767_), .B(\A[78] ), .Y(new_n4806_));
  OR2X1    g03804(.A(new_n4806_), .B(new_n4766_), .Y(new_n4807_));
  XOR2X1   g03805(.A(new_n4771_), .B(new_n4807_), .Y(new_n4808_));
  XOR2X1   g03806(.A(new_n4792_), .B(new_n4808_), .Y(new_n4809_));
  NOR4X1   g03807(.A(new_n4789_), .B(new_n4783_), .C(new_n4809_), .D(new_n4759_), .Y(new_n4810_));
  OR2X1    g03808(.A(new_n4781_), .B(new_n4776_), .Y(new_n4811_));
  OR2X1    g03809(.A(new_n4771_), .B(new_n4768_), .Y(new_n4812_));
  OAI21X1  g03810(.A0(new_n4811_), .A1(new_n4808_), .B0(new_n4812_), .Y(new_n4813_));
  XOR2X1   g03811(.A(new_n4781_), .B(new_n4776_), .Y(new_n4814_));
  OAI21X1  g03812(.A0(new_n4814_), .A1(new_n4795_), .B0(new_n4813_), .Y(new_n4815_));
  AOI22X1  g03813(.A0(new_n4815_), .A1(new_n4810_), .B0(new_n4796_), .B1(new_n4790_), .Y(new_n4816_));
  OAI21X1  g03814(.A0(new_n4816_), .A1(new_n4765_), .B0(new_n4805_), .Y(new_n4817_));
  AOI21X1  g03815(.A0(new_n4814_), .A1(new_n4813_), .B0(new_n4809_), .Y(new_n4818_));
  XOR2X1   g03816(.A(new_n4818_), .B(new_n4790_), .Y(new_n4819_));
  MX2X1    g03817(.A(new_n4816_), .B(new_n4819_), .S0(new_n4765_), .Y(new_n4820_));
  OAI22X1  g03818(.A0(new_n4820_), .A1(new_n4805_), .B0(new_n4817_), .B1(new_n4798_), .Y(new_n4821_));
  AND2X1   g03819(.A(new_n4821_), .B(new_n4733_), .Y(new_n4822_));
  XOR2X1   g03820(.A(new_n4745_), .B(new_n4758_), .Y(new_n4823_));
  XOR2X1   g03821(.A(new_n4823_), .B(new_n4799_), .Y(new_n4824_));
  XOR2X1   g03822(.A(new_n4804_), .B(new_n4824_), .Y(new_n4825_));
  INVX1    g03823(.A(new_n4591_), .Y(new_n4826_));
  XOR2X1   g03824(.A(new_n4826_), .B(new_n4555_), .Y(new_n4827_));
  NOR2X1   g03825(.A(new_n4827_), .B(new_n4825_), .Y(new_n4828_));
  NAND2X1  g03826(.A(new_n4797_), .B(new_n4765_), .Y(new_n4829_));
  NOR4X1   g03827(.A(new_n4789_), .B(new_n4783_), .C(new_n4782_), .D(new_n4759_), .Y(new_n4830_));
  OR4X1    g03828(.A(new_n4789_), .B(new_n4783_), .C(new_n4809_), .D(new_n4759_), .Y(new_n4831_));
  AOI21X1  g03829(.A0(new_n4789_), .A1(new_n4809_), .B0(new_n4794_), .Y(new_n4832_));
  OAI22X1  g03830(.A0(new_n4832_), .A1(new_n4831_), .B0(new_n4818_), .B1(new_n4830_), .Y(new_n4833_));
  MX2X1    g03831(.A(new_n4833_), .B(new_n4797_), .S0(new_n4765_), .Y(new_n4834_));
  XOR2X1   g03832(.A(new_n4752_), .B(new_n4760_), .Y(new_n4835_));
  XOR2X1   g03833(.A(new_n4745_), .B(new_n4739_), .Y(new_n4836_));
  OR2X1    g03834(.A(new_n4751_), .B(new_n4761_), .Y(new_n4837_));
  OAI21X1  g03835(.A0(new_n4752_), .A1(new_n4746_), .B0(new_n4837_), .Y(new_n4838_));
  AOI21X1  g03836(.A0(new_n4838_), .A1(new_n4836_), .B0(new_n4835_), .Y(new_n4839_));
  AOI21X1  g03837(.A0(new_n4833_), .A1(new_n4839_), .B0(new_n4805_), .Y(new_n4840_));
  AOI22X1  g03838(.A0(new_n4840_), .A1(new_n4829_), .B0(new_n4834_), .B1(new_n4805_), .Y(new_n4841_));
  OAI21X1  g03839(.A0(new_n4841_), .A1(new_n4733_), .B0(new_n4828_), .Y(new_n4842_));
  NOR4X1   g03840(.A(new_n4712_), .B(new_n4706_), .C(new_n4705_), .D(new_n4682_), .Y(new_n4843_));
  XOR2X1   g03841(.A(new_n4723_), .B(new_n4843_), .Y(new_n4844_));
  OR4X1    g03842(.A(new_n4712_), .B(new_n4706_), .C(new_n4721_), .D(new_n4682_), .Y(new_n4845_));
  AOI21X1  g03843(.A0(new_n4712_), .A1(new_n4721_), .B0(new_n4727_), .Y(new_n4846_));
  OAI22X1  g03844(.A0(new_n4846_), .A1(new_n4845_), .B0(new_n4723_), .B1(new_n4843_), .Y(new_n4847_));
  MX2X1    g03845(.A(new_n4847_), .B(new_n4844_), .S0(new_n4688_), .Y(new_n4848_));
  OR2X1    g03846(.A(new_n4804_), .B(new_n4801_), .Y(new_n4849_));
  AOI21X1  g03847(.A0(new_n4833_), .A1(new_n4839_), .B0(new_n4849_), .Y(new_n4850_));
  AOI22X1  g03848(.A0(new_n4834_), .A1(new_n4849_), .B0(new_n4850_), .B1(new_n4829_), .Y(new_n4851_));
  MX2X1    g03849(.A(new_n4851_), .B(new_n4841_), .S0(new_n4848_), .Y(new_n4852_));
  OAI22X1  g03850(.A0(new_n4852_), .A1(new_n4828_), .B0(new_n4842_), .B1(new_n4822_), .Y(new_n4853_));
  AND2X1   g03851(.A(new_n4853_), .B(new_n4656_), .Y(new_n4854_));
  XOR2X1   g03852(.A(new_n4827_), .B(new_n4825_), .Y(new_n4855_));
  INVX1    g03853(.A(new_n4855_), .Y(new_n4856_));
  INVX1    g03854(.A(new_n4382_), .Y(new_n4857_));
  XOR2X1   g03855(.A(new_n4421_), .B(new_n4857_), .Y(new_n4858_));
  XOR2X1   g03856(.A(new_n4281_), .B(new_n4294_), .Y(new_n4859_));
  XOR2X1   g03857(.A(new_n4859_), .B(new_n4335_), .Y(new_n4860_));
  AND2X1   g03858(.A(new_n4340_), .B(new_n4860_), .Y(new_n4861_));
  NOR2X1   g03859(.A(new_n4340_), .B(new_n4860_), .Y(new_n4862_));
  NOR3X1   g03860(.A(new_n4858_), .B(new_n4862_), .C(new_n4861_), .Y(new_n4863_));
  AOI21X1  g03861(.A0(new_n4858_), .A1(new_n4364_), .B0(new_n4863_), .Y(new_n4864_));
  NOR2X1   g03862(.A(new_n4864_), .B(new_n4856_), .Y(new_n4865_));
  OR2X1    g03863(.A(new_n4851_), .B(new_n4848_), .Y(new_n4866_));
  OAI21X1  g03864(.A0(new_n4816_), .A1(new_n4765_), .B0(new_n4849_), .Y(new_n4867_));
  OAI22X1  g03865(.A0(new_n4867_), .A1(new_n4798_), .B0(new_n4820_), .B1(new_n4849_), .Y(new_n4868_));
  MX2X1    g03866(.A(new_n4821_), .B(new_n4868_), .S0(new_n4848_), .Y(new_n4869_));
  AOI21X1  g03867(.A0(new_n4868_), .A1(new_n4848_), .B0(new_n4828_), .Y(new_n4870_));
  AOI22X1  g03868(.A0(new_n4870_), .A1(new_n4866_), .B0(new_n4869_), .B1(new_n4828_), .Y(new_n4871_));
  OAI21X1  g03869(.A0(new_n4871_), .A1(new_n4656_), .B0(new_n4865_), .Y(new_n4872_));
  OR2X1    g03870(.A(new_n4827_), .B(new_n4825_), .Y(new_n4873_));
  AOI21X1  g03871(.A0(new_n4868_), .A1(new_n4848_), .B0(new_n4873_), .Y(new_n4874_));
  AOI22X1  g03872(.A0(new_n4869_), .A1(new_n4873_), .B0(new_n4874_), .B1(new_n4866_), .Y(new_n4875_));
  MX2X1    g03873(.A(new_n4871_), .B(new_n4875_), .S0(new_n4656_), .Y(new_n4876_));
  OAI22X1  g03874(.A0(new_n4876_), .A1(new_n4865_), .B0(new_n4872_), .B1(new_n4854_), .Y(new_n4877_));
  AND2X1   g03875(.A(new_n4877_), .B(new_n4483_), .Y(new_n4878_));
  MX2X1    g03876(.A(new_n4267_), .B(new_n4254_), .S0(new_n4259_), .Y(new_n4879_));
  AND2X1   g03877(.A(new_n4435_), .B(new_n4879_), .Y(new_n4880_));
  AOI21X1  g03878(.A0(new_n4359_), .A1(new_n4346_), .B0(new_n4433_), .Y(new_n4881_));
  AOI22X1  g03879(.A0(new_n4881_), .A1(new_n4334_), .B0(new_n4361_), .B1(new_n4433_), .Y(new_n4882_));
  OAI21X1  g03880(.A0(new_n4882_), .A1(new_n4879_), .B0(new_n4480_), .Y(new_n4883_));
  MX2X1    g03881(.A(new_n4362_), .B(new_n4882_), .S0(new_n4269_), .Y(new_n4884_));
  OAI22X1  g03882(.A0(new_n4884_), .A1(new_n4480_), .B0(new_n4883_), .B1(new_n4880_), .Y(new_n4885_));
  OAI21X1  g03883(.A0(new_n4882_), .A1(new_n4879_), .B0(new_n4423_), .Y(new_n4886_));
  OAI22X1  g03884(.A0(new_n4886_), .A1(new_n4880_), .B0(new_n4884_), .B1(new_n4423_), .Y(new_n4887_));
  MX2X1    g03885(.A(new_n4885_), .B(new_n4887_), .S0(new_n4479_), .Y(new_n4888_));
  OR2X1    g03886(.A(new_n4864_), .B(new_n4856_), .Y(new_n4889_));
  OAI21X1  g03887(.A0(new_n4871_), .A1(new_n4656_), .B0(new_n4889_), .Y(new_n4890_));
  OAI22X1  g03888(.A0(new_n4890_), .A1(new_n4854_), .B0(new_n4876_), .B1(new_n4889_), .Y(new_n4891_));
  AND2X1   g03889(.A(new_n4891_), .B(new_n4888_), .Y(new_n4892_));
  XOR2X1   g03890(.A(new_n4864_), .B(new_n4855_), .Y(new_n4893_));
  XOR2X1   g03891(.A(new_n4087_), .B(new_n4011_), .Y(new_n4894_));
  INVX1    g03892(.A(new_n4894_), .Y(new_n4895_));
  OR4X1    g03893(.A(new_n4895_), .B(new_n4893_), .C(new_n4892_), .D(new_n4878_), .Y(new_n4896_));
  NOR2X1   g03894(.A(new_n4895_), .B(new_n4893_), .Y(new_n4897_));
  AND2X1   g03895(.A(new_n4547_), .B(new_n4515_), .Y(new_n4898_));
  NOR4X1   g03896(.A(new_n4539_), .B(new_n4533_), .C(new_n4605_), .D(new_n4509_), .Y(new_n4899_));
  OAI21X1  g03897(.A0(new_n4552_), .A1(new_n4545_), .B0(new_n4604_), .Y(new_n4900_));
  AOI22X1  g03898(.A0(new_n4900_), .A1(new_n4899_), .B0(new_n4546_), .B1(new_n4540_), .Y(new_n4901_));
  OAI21X1  g03899(.A0(new_n4901_), .A1(new_n4515_), .B0(new_n4653_), .Y(new_n4902_));
  XOR2X1   g03900(.A(new_n4606_), .B(new_n4540_), .Y(new_n4903_));
  MX2X1    g03901(.A(new_n4901_), .B(new_n4903_), .S0(new_n4515_), .Y(new_n4904_));
  OAI22X1  g03902(.A0(new_n4904_), .A1(new_n4653_), .B0(new_n4902_), .B1(new_n4898_), .Y(new_n4905_));
  OAI21X1  g03903(.A0(new_n4901_), .A1(new_n4515_), .B0(new_n4592_), .Y(new_n4906_));
  OAI22X1  g03904(.A0(new_n4906_), .A1(new_n4898_), .B0(new_n4904_), .B1(new_n4592_), .Y(new_n4907_));
  MX2X1    g03905(.A(new_n4907_), .B(new_n4905_), .S0(new_n4652_), .Y(new_n4908_));
  OR2X1    g03906(.A(new_n4875_), .B(new_n4908_), .Y(new_n4909_));
  OAI21X1  g03907(.A0(new_n4841_), .A1(new_n4733_), .B0(new_n4873_), .Y(new_n4910_));
  OAI22X1  g03908(.A0(new_n4910_), .A1(new_n4822_), .B0(new_n4852_), .B1(new_n4873_), .Y(new_n4911_));
  AOI21X1  g03909(.A0(new_n4911_), .A1(new_n4908_), .B0(new_n4889_), .Y(new_n4912_));
  MX2X1    g03910(.A(new_n4911_), .B(new_n4853_), .S0(new_n4656_), .Y(new_n4913_));
  AOI22X1  g03911(.A0(new_n4913_), .A1(new_n4889_), .B0(new_n4912_), .B1(new_n4909_), .Y(new_n4914_));
  AOI21X1  g03912(.A0(new_n4911_), .A1(new_n4908_), .B0(new_n4865_), .Y(new_n4915_));
  AOI22X1  g03913(.A0(new_n4915_), .A1(new_n4909_), .B0(new_n4913_), .B1(new_n4865_), .Y(new_n4916_));
  MX2X1    g03914(.A(new_n4916_), .B(new_n4914_), .S0(new_n4483_), .Y(new_n4917_));
  OR2X1    g03915(.A(new_n4917_), .B(new_n4897_), .Y(new_n4918_));
  AOI21X1  g03916(.A0(new_n4918_), .A1(new_n4896_), .B0(new_n4186_), .Y(new_n4919_));
  INVX1    g03917(.A(new_n4897_), .Y(new_n4920_));
  OAI21X1  g03918(.A0(new_n4916_), .A1(new_n4483_), .B0(new_n4920_), .Y(new_n4921_));
  OAI22X1  g03919(.A0(new_n4921_), .A1(new_n4878_), .B0(new_n4917_), .B1(new_n4920_), .Y(new_n4922_));
  AND2X1   g03920(.A(new_n4922_), .B(new_n4186_), .Y(new_n4923_));
  OR2X1    g03921(.A(new_n4894_), .B(new_n4893_), .Y(new_n4924_));
  AOI21X1  g03922(.A0(new_n4864_), .A1(new_n4855_), .B0(new_n4895_), .Y(new_n4925_));
  OAI21X1  g03923(.A0(new_n4864_), .A1(new_n4855_), .B0(new_n4925_), .Y(new_n4926_));
  NAND2X1  g03924(.A(new_n4926_), .B(new_n4924_), .Y(new_n4927_));
  INVX1    g03925(.A(\A[937] ), .Y(new_n4928_));
  OR2X1    g03926(.A(\A[938] ), .B(new_n4928_), .Y(new_n4929_));
  INVX1    g03927(.A(\A[939] ), .Y(new_n4930_));
  AOI21X1  g03928(.A0(\A[938] ), .A1(new_n4928_), .B0(new_n4930_), .Y(new_n4931_));
  XOR2X1   g03929(.A(\A[938] ), .B(\A[937] ), .Y(new_n4932_));
  AND2X1   g03930(.A(new_n4932_), .B(new_n4930_), .Y(new_n4933_));
  AOI21X1  g03931(.A0(new_n4931_), .A1(new_n4929_), .B0(new_n4933_), .Y(new_n4934_));
  INVX1    g03932(.A(\A[942] ), .Y(new_n4935_));
  INVX1    g03933(.A(\A[940] ), .Y(new_n4936_));
  OR2X1    g03934(.A(\A[941] ), .B(new_n4936_), .Y(new_n4937_));
  AOI21X1  g03935(.A0(\A[941] ), .A1(new_n4936_), .B0(new_n4935_), .Y(new_n4938_));
  XOR2X1   g03936(.A(\A[941] ), .B(\A[940] ), .Y(new_n4939_));
  AOI22X1  g03937(.A0(new_n4939_), .A1(new_n4935_), .B0(new_n4938_), .B1(new_n4937_), .Y(new_n4940_));
  AND2X1   g03938(.A(\A[941] ), .B(\A[940] ), .Y(new_n4941_));
  AOI21X1  g03939(.A0(new_n4939_), .A1(\A[942] ), .B0(new_n4941_), .Y(new_n4942_));
  AND2X1   g03940(.A(\A[938] ), .B(\A[937] ), .Y(new_n4943_));
  AOI21X1  g03941(.A0(new_n4932_), .A1(\A[939] ), .B0(new_n4943_), .Y(new_n4944_));
  XOR2X1   g03942(.A(new_n4940_), .B(new_n4934_), .Y(new_n4945_));
  INVX1    g03943(.A(\A[931] ), .Y(new_n4946_));
  OR2X1    g03944(.A(\A[932] ), .B(new_n4946_), .Y(new_n4947_));
  INVX1    g03945(.A(\A[933] ), .Y(new_n4948_));
  AOI21X1  g03946(.A0(\A[932] ), .A1(new_n4946_), .B0(new_n4948_), .Y(new_n4949_));
  XOR2X1   g03947(.A(\A[932] ), .B(\A[931] ), .Y(new_n4950_));
  AND2X1   g03948(.A(new_n4950_), .B(new_n4948_), .Y(new_n4951_));
  AOI21X1  g03949(.A0(new_n4949_), .A1(new_n4947_), .B0(new_n4951_), .Y(new_n4952_));
  INVX1    g03950(.A(\A[936] ), .Y(new_n4953_));
  INVX1    g03951(.A(\A[934] ), .Y(new_n4954_));
  OR2X1    g03952(.A(\A[935] ), .B(new_n4954_), .Y(new_n4955_));
  AOI21X1  g03953(.A0(\A[935] ), .A1(new_n4954_), .B0(new_n4953_), .Y(new_n4956_));
  XOR2X1   g03954(.A(\A[935] ), .B(\A[934] ), .Y(new_n4957_));
  AOI22X1  g03955(.A0(new_n4957_), .A1(new_n4953_), .B0(new_n4956_), .B1(new_n4955_), .Y(new_n4958_));
  AND2X1   g03956(.A(\A[935] ), .B(\A[934] ), .Y(new_n4959_));
  AOI21X1  g03957(.A0(new_n4957_), .A1(\A[936] ), .B0(new_n4959_), .Y(new_n4960_));
  AND2X1   g03958(.A(\A[932] ), .B(\A[931] ), .Y(new_n4961_));
  AOI21X1  g03959(.A0(new_n4950_), .A1(\A[933] ), .B0(new_n4961_), .Y(new_n4962_));
  XOR2X1   g03960(.A(new_n4958_), .B(new_n4952_), .Y(new_n4963_));
  XOR2X1   g03961(.A(new_n4963_), .B(new_n4945_), .Y(new_n4964_));
  INVX1    g03962(.A(\A[925] ), .Y(new_n4965_));
  OR2X1    g03963(.A(\A[926] ), .B(new_n4965_), .Y(new_n4966_));
  INVX1    g03964(.A(\A[927] ), .Y(new_n4967_));
  AOI21X1  g03965(.A0(\A[926] ), .A1(new_n4965_), .B0(new_n4967_), .Y(new_n4968_));
  AND2X1   g03966(.A(new_n4968_), .B(new_n4966_), .Y(new_n4969_));
  XOR2X1   g03967(.A(\A[926] ), .B(\A[925] ), .Y(new_n4970_));
  AND2X1   g03968(.A(new_n4970_), .B(new_n4967_), .Y(new_n4971_));
  OR2X1    g03969(.A(new_n4971_), .B(new_n4969_), .Y(new_n4972_));
  INVX1    g03970(.A(\A[930] ), .Y(new_n4973_));
  INVX1    g03971(.A(\A[928] ), .Y(new_n4974_));
  OR2X1    g03972(.A(\A[929] ), .B(new_n4974_), .Y(new_n4975_));
  AOI21X1  g03973(.A0(\A[929] ), .A1(new_n4974_), .B0(new_n4973_), .Y(new_n4976_));
  XOR2X1   g03974(.A(\A[929] ), .B(\A[928] ), .Y(new_n4977_));
  AOI22X1  g03975(.A0(new_n4977_), .A1(new_n4973_), .B0(new_n4976_), .B1(new_n4975_), .Y(new_n4978_));
  AND2X1   g03976(.A(\A[929] ), .B(\A[928] ), .Y(new_n4979_));
  AOI21X1  g03977(.A0(new_n4977_), .A1(\A[930] ), .B0(new_n4979_), .Y(new_n4980_));
  AND2X1   g03978(.A(\A[926] ), .B(\A[925] ), .Y(new_n4981_));
  AOI21X1  g03979(.A0(new_n4970_), .A1(\A[927] ), .B0(new_n4981_), .Y(new_n4982_));
  XOR2X1   g03980(.A(new_n4978_), .B(new_n4972_), .Y(new_n4983_));
  INVX1    g03981(.A(\A[919] ), .Y(new_n4984_));
  OR2X1    g03982(.A(\A[920] ), .B(new_n4984_), .Y(new_n4985_));
  INVX1    g03983(.A(\A[921] ), .Y(new_n4986_));
  AOI21X1  g03984(.A0(\A[920] ), .A1(new_n4984_), .B0(new_n4986_), .Y(new_n4987_));
  XOR2X1   g03985(.A(\A[920] ), .B(\A[919] ), .Y(new_n4988_));
  AND2X1   g03986(.A(new_n4988_), .B(new_n4986_), .Y(new_n4989_));
  AOI21X1  g03987(.A0(new_n4987_), .A1(new_n4985_), .B0(new_n4989_), .Y(new_n4990_));
  INVX1    g03988(.A(\A[924] ), .Y(new_n4991_));
  INVX1    g03989(.A(\A[922] ), .Y(new_n4992_));
  OR2X1    g03990(.A(\A[923] ), .B(new_n4992_), .Y(new_n4993_));
  AOI21X1  g03991(.A0(\A[923] ), .A1(new_n4992_), .B0(new_n4991_), .Y(new_n4994_));
  XOR2X1   g03992(.A(\A[923] ), .B(\A[922] ), .Y(new_n4995_));
  AOI22X1  g03993(.A0(new_n4995_), .A1(new_n4991_), .B0(new_n4994_), .B1(new_n4993_), .Y(new_n4996_));
  AND2X1   g03994(.A(\A[923] ), .B(\A[922] ), .Y(new_n4997_));
  AOI21X1  g03995(.A0(new_n4995_), .A1(\A[924] ), .B0(new_n4997_), .Y(new_n4998_));
  AND2X1   g03996(.A(\A[920] ), .B(\A[919] ), .Y(new_n4999_));
  AOI21X1  g03997(.A0(new_n4988_), .A1(\A[921] ), .B0(new_n4999_), .Y(new_n5000_));
  XOR2X1   g03998(.A(new_n4996_), .B(new_n4990_), .Y(new_n5001_));
  XOR2X1   g03999(.A(new_n5001_), .B(new_n4983_), .Y(new_n5002_));
  XOR2X1   g04000(.A(new_n5002_), .B(new_n4964_), .Y(new_n5003_));
  INVX1    g04001(.A(\A[913] ), .Y(new_n5004_));
  OR2X1    g04002(.A(\A[914] ), .B(new_n5004_), .Y(new_n5005_));
  INVX1    g04003(.A(\A[915] ), .Y(new_n5006_));
  AOI21X1  g04004(.A0(\A[914] ), .A1(new_n5004_), .B0(new_n5006_), .Y(new_n5007_));
  XOR2X1   g04005(.A(\A[914] ), .B(\A[913] ), .Y(new_n5008_));
  AND2X1   g04006(.A(new_n5008_), .B(new_n5006_), .Y(new_n5009_));
  AOI21X1  g04007(.A0(new_n5007_), .A1(new_n5005_), .B0(new_n5009_), .Y(new_n5010_));
  INVX1    g04008(.A(\A[918] ), .Y(new_n5011_));
  INVX1    g04009(.A(\A[916] ), .Y(new_n5012_));
  OR2X1    g04010(.A(\A[917] ), .B(new_n5012_), .Y(new_n5013_));
  AOI21X1  g04011(.A0(\A[917] ), .A1(new_n5012_), .B0(new_n5011_), .Y(new_n5014_));
  XOR2X1   g04012(.A(\A[917] ), .B(\A[916] ), .Y(new_n5015_));
  AOI22X1  g04013(.A0(new_n5015_), .A1(new_n5011_), .B0(new_n5014_), .B1(new_n5013_), .Y(new_n5016_));
  AND2X1   g04014(.A(\A[917] ), .B(\A[916] ), .Y(new_n5017_));
  AOI21X1  g04015(.A0(new_n5015_), .A1(\A[918] ), .B0(new_n5017_), .Y(new_n5018_));
  AND2X1   g04016(.A(\A[914] ), .B(\A[913] ), .Y(new_n5019_));
  AOI21X1  g04017(.A0(new_n5008_), .A1(\A[915] ), .B0(new_n5019_), .Y(new_n5020_));
  XOR2X1   g04018(.A(new_n5016_), .B(new_n5010_), .Y(new_n5021_));
  INVX1    g04019(.A(\A[907] ), .Y(new_n5022_));
  OR2X1    g04020(.A(\A[908] ), .B(new_n5022_), .Y(new_n5023_));
  INVX1    g04021(.A(\A[909] ), .Y(new_n5024_));
  AOI21X1  g04022(.A0(\A[908] ), .A1(new_n5022_), .B0(new_n5024_), .Y(new_n5025_));
  XOR2X1   g04023(.A(\A[908] ), .B(\A[907] ), .Y(new_n5026_));
  AND2X1   g04024(.A(new_n5026_), .B(new_n5024_), .Y(new_n5027_));
  AOI21X1  g04025(.A0(new_n5025_), .A1(new_n5023_), .B0(new_n5027_), .Y(new_n5028_));
  INVX1    g04026(.A(\A[912] ), .Y(new_n5029_));
  INVX1    g04027(.A(\A[910] ), .Y(new_n5030_));
  OR2X1    g04028(.A(\A[911] ), .B(new_n5030_), .Y(new_n5031_));
  AOI21X1  g04029(.A0(\A[911] ), .A1(new_n5030_), .B0(new_n5029_), .Y(new_n5032_));
  XOR2X1   g04030(.A(\A[911] ), .B(\A[910] ), .Y(new_n5033_));
  AOI22X1  g04031(.A0(new_n5033_), .A1(new_n5029_), .B0(new_n5032_), .B1(new_n5031_), .Y(new_n5034_));
  AND2X1   g04032(.A(\A[911] ), .B(\A[910] ), .Y(new_n5035_));
  AOI21X1  g04033(.A0(new_n5033_), .A1(\A[912] ), .B0(new_n5035_), .Y(new_n5036_));
  AND2X1   g04034(.A(\A[908] ), .B(\A[907] ), .Y(new_n5037_));
  AOI21X1  g04035(.A0(new_n5026_), .A1(\A[909] ), .B0(new_n5037_), .Y(new_n5038_));
  XOR2X1   g04036(.A(new_n5034_), .B(new_n5028_), .Y(new_n5039_));
  XOR2X1   g04037(.A(new_n5039_), .B(new_n5021_), .Y(new_n5040_));
  INVX1    g04038(.A(new_n5040_), .Y(new_n5041_));
  INVX1    g04039(.A(\A[901] ), .Y(new_n5042_));
  OR2X1    g04040(.A(\A[902] ), .B(new_n5042_), .Y(new_n5043_));
  INVX1    g04041(.A(\A[903] ), .Y(new_n5044_));
  AOI21X1  g04042(.A0(\A[902] ), .A1(new_n5042_), .B0(new_n5044_), .Y(new_n5045_));
  AND2X1   g04043(.A(new_n5045_), .B(new_n5043_), .Y(new_n5046_));
  XOR2X1   g04044(.A(\A[902] ), .B(\A[901] ), .Y(new_n5047_));
  AND2X1   g04045(.A(new_n5047_), .B(new_n5044_), .Y(new_n5048_));
  OR2X1    g04046(.A(new_n5048_), .B(new_n5046_), .Y(new_n5049_));
  INVX1    g04047(.A(\A[906] ), .Y(new_n5050_));
  INVX1    g04048(.A(\A[904] ), .Y(new_n5051_));
  OR2X1    g04049(.A(\A[905] ), .B(new_n5051_), .Y(new_n5052_));
  AOI21X1  g04050(.A0(\A[905] ), .A1(new_n5051_), .B0(new_n5050_), .Y(new_n5053_));
  XOR2X1   g04051(.A(\A[905] ), .B(\A[904] ), .Y(new_n5054_));
  AOI22X1  g04052(.A0(new_n5054_), .A1(new_n5050_), .B0(new_n5053_), .B1(new_n5052_), .Y(new_n5055_));
  AND2X1   g04053(.A(\A[905] ), .B(\A[904] ), .Y(new_n5056_));
  AOI21X1  g04054(.A0(new_n5054_), .A1(\A[906] ), .B0(new_n5056_), .Y(new_n5057_));
  AND2X1   g04055(.A(\A[902] ), .B(\A[901] ), .Y(new_n5058_));
  AOI21X1  g04056(.A0(new_n5047_), .A1(\A[903] ), .B0(new_n5058_), .Y(new_n5059_));
  XOR2X1   g04057(.A(new_n5055_), .B(new_n5049_), .Y(new_n5060_));
  INVX1    g04058(.A(\A[895] ), .Y(new_n5061_));
  OR2X1    g04059(.A(\A[896] ), .B(new_n5061_), .Y(new_n5062_));
  INVX1    g04060(.A(\A[897] ), .Y(new_n5063_));
  AOI21X1  g04061(.A0(\A[896] ), .A1(new_n5061_), .B0(new_n5063_), .Y(new_n5064_));
  XOR2X1   g04062(.A(\A[896] ), .B(\A[895] ), .Y(new_n5065_));
  AND2X1   g04063(.A(new_n5065_), .B(new_n5063_), .Y(new_n5066_));
  AOI21X1  g04064(.A0(new_n5064_), .A1(new_n5062_), .B0(new_n5066_), .Y(new_n5067_));
  INVX1    g04065(.A(\A[900] ), .Y(new_n5068_));
  INVX1    g04066(.A(\A[898] ), .Y(new_n5069_));
  OR2X1    g04067(.A(\A[899] ), .B(new_n5069_), .Y(new_n5070_));
  AOI21X1  g04068(.A0(\A[899] ), .A1(new_n5069_), .B0(new_n5068_), .Y(new_n5071_));
  XOR2X1   g04069(.A(\A[899] ), .B(\A[898] ), .Y(new_n5072_));
  AOI22X1  g04070(.A0(new_n5072_), .A1(new_n5068_), .B0(new_n5071_), .B1(new_n5070_), .Y(new_n5073_));
  AND2X1   g04071(.A(\A[899] ), .B(\A[898] ), .Y(new_n5074_));
  AOI21X1  g04072(.A0(new_n5072_), .A1(\A[900] ), .B0(new_n5074_), .Y(new_n5075_));
  AND2X1   g04073(.A(\A[896] ), .B(\A[895] ), .Y(new_n5076_));
  AOI21X1  g04074(.A0(new_n5065_), .A1(\A[897] ), .B0(new_n5076_), .Y(new_n5077_));
  XOR2X1   g04075(.A(new_n5073_), .B(new_n5067_), .Y(new_n5078_));
  XOR2X1   g04076(.A(new_n5078_), .B(new_n5060_), .Y(new_n5079_));
  XOR2X1   g04077(.A(new_n5079_), .B(new_n5041_), .Y(new_n5080_));
  XOR2X1   g04078(.A(new_n5080_), .B(new_n5003_), .Y(new_n5081_));
  INVX1    g04079(.A(\A[889] ), .Y(new_n5082_));
  OR2X1    g04080(.A(\A[890] ), .B(new_n5082_), .Y(new_n5083_));
  INVX1    g04081(.A(\A[891] ), .Y(new_n5084_));
  AOI21X1  g04082(.A0(\A[890] ), .A1(new_n5082_), .B0(new_n5084_), .Y(new_n5085_));
  XOR2X1   g04083(.A(\A[890] ), .B(\A[889] ), .Y(new_n5086_));
  AND2X1   g04084(.A(new_n5086_), .B(new_n5084_), .Y(new_n5087_));
  AOI21X1  g04085(.A0(new_n5085_), .A1(new_n5083_), .B0(new_n5087_), .Y(new_n5088_));
  INVX1    g04086(.A(\A[894] ), .Y(new_n5089_));
  INVX1    g04087(.A(\A[892] ), .Y(new_n5090_));
  OR2X1    g04088(.A(\A[893] ), .B(new_n5090_), .Y(new_n5091_));
  AOI21X1  g04089(.A0(\A[893] ), .A1(new_n5090_), .B0(new_n5089_), .Y(new_n5092_));
  XOR2X1   g04090(.A(\A[893] ), .B(\A[892] ), .Y(new_n5093_));
  AOI22X1  g04091(.A0(new_n5093_), .A1(new_n5089_), .B0(new_n5092_), .B1(new_n5091_), .Y(new_n5094_));
  AND2X1   g04092(.A(\A[893] ), .B(\A[892] ), .Y(new_n5095_));
  AOI21X1  g04093(.A0(new_n5093_), .A1(\A[894] ), .B0(new_n5095_), .Y(new_n5096_));
  AND2X1   g04094(.A(\A[890] ), .B(\A[889] ), .Y(new_n5097_));
  AOI21X1  g04095(.A0(new_n5086_), .A1(\A[891] ), .B0(new_n5097_), .Y(new_n5098_));
  XOR2X1   g04096(.A(new_n5094_), .B(new_n5088_), .Y(new_n5099_));
  INVX1    g04097(.A(\A[883] ), .Y(new_n5100_));
  OR2X1    g04098(.A(\A[884] ), .B(new_n5100_), .Y(new_n5101_));
  INVX1    g04099(.A(\A[885] ), .Y(new_n5102_));
  AOI21X1  g04100(.A0(\A[884] ), .A1(new_n5100_), .B0(new_n5102_), .Y(new_n5103_));
  XOR2X1   g04101(.A(\A[884] ), .B(\A[883] ), .Y(new_n5104_));
  AND2X1   g04102(.A(new_n5104_), .B(new_n5102_), .Y(new_n5105_));
  AOI21X1  g04103(.A0(new_n5103_), .A1(new_n5101_), .B0(new_n5105_), .Y(new_n5106_));
  INVX1    g04104(.A(\A[888] ), .Y(new_n5107_));
  INVX1    g04105(.A(\A[886] ), .Y(new_n5108_));
  OR2X1    g04106(.A(\A[887] ), .B(new_n5108_), .Y(new_n5109_));
  AOI21X1  g04107(.A0(\A[887] ), .A1(new_n5108_), .B0(new_n5107_), .Y(new_n5110_));
  XOR2X1   g04108(.A(\A[887] ), .B(\A[886] ), .Y(new_n5111_));
  AOI22X1  g04109(.A0(new_n5111_), .A1(new_n5107_), .B0(new_n5110_), .B1(new_n5109_), .Y(new_n5112_));
  AND2X1   g04110(.A(\A[887] ), .B(\A[886] ), .Y(new_n5113_));
  AOI21X1  g04111(.A0(new_n5111_), .A1(\A[888] ), .B0(new_n5113_), .Y(new_n5114_));
  AND2X1   g04112(.A(\A[884] ), .B(\A[883] ), .Y(new_n5115_));
  AOI21X1  g04113(.A0(new_n5104_), .A1(\A[885] ), .B0(new_n5115_), .Y(new_n5116_));
  XOR2X1   g04114(.A(new_n5112_), .B(new_n5106_), .Y(new_n5117_));
  XOR2X1   g04115(.A(new_n5117_), .B(new_n5099_), .Y(new_n5118_));
  INVX1    g04116(.A(\A[877] ), .Y(new_n5119_));
  OR2X1    g04117(.A(\A[878] ), .B(new_n5119_), .Y(new_n5120_));
  INVX1    g04118(.A(\A[879] ), .Y(new_n5121_));
  AOI21X1  g04119(.A0(\A[878] ), .A1(new_n5119_), .B0(new_n5121_), .Y(new_n5122_));
  AND2X1   g04120(.A(new_n5122_), .B(new_n5120_), .Y(new_n5123_));
  XOR2X1   g04121(.A(\A[878] ), .B(\A[877] ), .Y(new_n5124_));
  AND2X1   g04122(.A(new_n5124_), .B(new_n5121_), .Y(new_n5125_));
  OR2X1    g04123(.A(new_n5125_), .B(new_n5123_), .Y(new_n5126_));
  INVX1    g04124(.A(\A[882] ), .Y(new_n5127_));
  INVX1    g04125(.A(\A[880] ), .Y(new_n5128_));
  OR2X1    g04126(.A(\A[881] ), .B(new_n5128_), .Y(new_n5129_));
  AOI21X1  g04127(.A0(\A[881] ), .A1(new_n5128_), .B0(new_n5127_), .Y(new_n5130_));
  XOR2X1   g04128(.A(\A[881] ), .B(\A[880] ), .Y(new_n5131_));
  AOI22X1  g04129(.A0(new_n5131_), .A1(new_n5127_), .B0(new_n5130_), .B1(new_n5129_), .Y(new_n5132_));
  AND2X1   g04130(.A(\A[881] ), .B(\A[880] ), .Y(new_n5133_));
  AOI21X1  g04131(.A0(new_n5131_), .A1(\A[882] ), .B0(new_n5133_), .Y(new_n5134_));
  AND2X1   g04132(.A(\A[878] ), .B(\A[877] ), .Y(new_n5135_));
  AOI21X1  g04133(.A0(new_n5124_), .A1(\A[879] ), .B0(new_n5135_), .Y(new_n5136_));
  XOR2X1   g04134(.A(new_n5132_), .B(new_n5126_), .Y(new_n5137_));
  INVX1    g04135(.A(\A[871] ), .Y(new_n5138_));
  OR2X1    g04136(.A(\A[872] ), .B(new_n5138_), .Y(new_n5139_));
  INVX1    g04137(.A(\A[873] ), .Y(new_n5140_));
  AOI21X1  g04138(.A0(\A[872] ), .A1(new_n5138_), .B0(new_n5140_), .Y(new_n5141_));
  XOR2X1   g04139(.A(\A[872] ), .B(\A[871] ), .Y(new_n5142_));
  AND2X1   g04140(.A(new_n5142_), .B(new_n5140_), .Y(new_n5143_));
  AOI21X1  g04141(.A0(new_n5141_), .A1(new_n5139_), .B0(new_n5143_), .Y(new_n5144_));
  INVX1    g04142(.A(\A[876] ), .Y(new_n5145_));
  INVX1    g04143(.A(\A[874] ), .Y(new_n5146_));
  OR2X1    g04144(.A(\A[875] ), .B(new_n5146_), .Y(new_n5147_));
  AOI21X1  g04145(.A0(\A[875] ), .A1(new_n5146_), .B0(new_n5145_), .Y(new_n5148_));
  XOR2X1   g04146(.A(\A[875] ), .B(\A[874] ), .Y(new_n5149_));
  AOI22X1  g04147(.A0(new_n5149_), .A1(new_n5145_), .B0(new_n5148_), .B1(new_n5147_), .Y(new_n5150_));
  AND2X1   g04148(.A(\A[875] ), .B(\A[874] ), .Y(new_n5151_));
  AOI21X1  g04149(.A0(new_n5149_), .A1(\A[876] ), .B0(new_n5151_), .Y(new_n5152_));
  AND2X1   g04150(.A(\A[872] ), .B(\A[871] ), .Y(new_n5153_));
  AOI21X1  g04151(.A0(new_n5142_), .A1(\A[873] ), .B0(new_n5153_), .Y(new_n5154_));
  XOR2X1   g04152(.A(new_n5150_), .B(new_n5144_), .Y(new_n5155_));
  XOR2X1   g04153(.A(new_n5155_), .B(new_n5137_), .Y(new_n5156_));
  XOR2X1   g04154(.A(new_n5156_), .B(new_n5118_), .Y(new_n5157_));
  INVX1    g04155(.A(\A[865] ), .Y(new_n5158_));
  OR2X1    g04156(.A(\A[866] ), .B(new_n5158_), .Y(new_n5159_));
  INVX1    g04157(.A(\A[867] ), .Y(new_n5160_));
  AOI21X1  g04158(.A0(\A[866] ), .A1(new_n5158_), .B0(new_n5160_), .Y(new_n5161_));
  XOR2X1   g04159(.A(\A[866] ), .B(\A[865] ), .Y(new_n5162_));
  AND2X1   g04160(.A(new_n5162_), .B(new_n5160_), .Y(new_n5163_));
  AOI21X1  g04161(.A0(new_n5161_), .A1(new_n5159_), .B0(new_n5163_), .Y(new_n5164_));
  INVX1    g04162(.A(\A[870] ), .Y(new_n5165_));
  INVX1    g04163(.A(\A[868] ), .Y(new_n5166_));
  OR2X1    g04164(.A(\A[869] ), .B(new_n5166_), .Y(new_n5167_));
  AOI21X1  g04165(.A0(\A[869] ), .A1(new_n5166_), .B0(new_n5165_), .Y(new_n5168_));
  XOR2X1   g04166(.A(\A[869] ), .B(\A[868] ), .Y(new_n5169_));
  AOI22X1  g04167(.A0(new_n5169_), .A1(new_n5165_), .B0(new_n5168_), .B1(new_n5167_), .Y(new_n5170_));
  AND2X1   g04168(.A(\A[869] ), .B(\A[868] ), .Y(new_n5171_));
  AOI21X1  g04169(.A0(new_n5169_), .A1(\A[870] ), .B0(new_n5171_), .Y(new_n5172_));
  AND2X1   g04170(.A(\A[866] ), .B(\A[865] ), .Y(new_n5173_));
  AOI21X1  g04171(.A0(new_n5162_), .A1(\A[867] ), .B0(new_n5173_), .Y(new_n5174_));
  XOR2X1   g04172(.A(new_n5170_), .B(new_n5164_), .Y(new_n5175_));
  INVX1    g04173(.A(\A[859] ), .Y(new_n5176_));
  OR2X1    g04174(.A(\A[860] ), .B(new_n5176_), .Y(new_n5177_));
  INVX1    g04175(.A(\A[861] ), .Y(new_n5178_));
  AOI21X1  g04176(.A0(\A[860] ), .A1(new_n5176_), .B0(new_n5178_), .Y(new_n5179_));
  XOR2X1   g04177(.A(\A[860] ), .B(\A[859] ), .Y(new_n5180_));
  AND2X1   g04178(.A(new_n5180_), .B(new_n5178_), .Y(new_n5181_));
  AOI21X1  g04179(.A0(new_n5179_), .A1(new_n5177_), .B0(new_n5181_), .Y(new_n5182_));
  INVX1    g04180(.A(\A[864] ), .Y(new_n5183_));
  INVX1    g04181(.A(\A[862] ), .Y(new_n5184_));
  OR2X1    g04182(.A(\A[863] ), .B(new_n5184_), .Y(new_n5185_));
  AOI21X1  g04183(.A0(\A[863] ), .A1(new_n5184_), .B0(new_n5183_), .Y(new_n5186_));
  XOR2X1   g04184(.A(\A[863] ), .B(\A[862] ), .Y(new_n5187_));
  AOI22X1  g04185(.A0(new_n5187_), .A1(new_n5183_), .B0(new_n5186_), .B1(new_n5185_), .Y(new_n5188_));
  AND2X1   g04186(.A(\A[863] ), .B(\A[862] ), .Y(new_n5189_));
  AOI21X1  g04187(.A0(new_n5187_), .A1(\A[864] ), .B0(new_n5189_), .Y(new_n5190_));
  AND2X1   g04188(.A(\A[860] ), .B(\A[859] ), .Y(new_n5191_));
  AOI21X1  g04189(.A0(new_n5180_), .A1(\A[861] ), .B0(new_n5191_), .Y(new_n5192_));
  XOR2X1   g04190(.A(new_n5188_), .B(new_n5182_), .Y(new_n5193_));
  XOR2X1   g04191(.A(new_n5193_), .B(new_n5175_), .Y(new_n5194_));
  INVX1    g04192(.A(new_n5194_), .Y(new_n5195_));
  INVX1    g04193(.A(\A[853] ), .Y(new_n5196_));
  OR2X1    g04194(.A(\A[854] ), .B(new_n5196_), .Y(new_n5197_));
  INVX1    g04195(.A(\A[855] ), .Y(new_n5198_));
  AOI21X1  g04196(.A0(\A[854] ), .A1(new_n5196_), .B0(new_n5198_), .Y(new_n5199_));
  AND2X1   g04197(.A(new_n5199_), .B(new_n5197_), .Y(new_n5200_));
  XOR2X1   g04198(.A(\A[854] ), .B(\A[853] ), .Y(new_n5201_));
  AND2X1   g04199(.A(new_n5201_), .B(new_n5198_), .Y(new_n5202_));
  OR2X1    g04200(.A(new_n5202_), .B(new_n5200_), .Y(new_n5203_));
  INVX1    g04201(.A(\A[858] ), .Y(new_n5204_));
  INVX1    g04202(.A(\A[856] ), .Y(new_n5205_));
  OR2X1    g04203(.A(\A[857] ), .B(new_n5205_), .Y(new_n5206_));
  AOI21X1  g04204(.A0(\A[857] ), .A1(new_n5205_), .B0(new_n5204_), .Y(new_n5207_));
  XOR2X1   g04205(.A(\A[857] ), .B(\A[856] ), .Y(new_n5208_));
  AOI22X1  g04206(.A0(new_n5208_), .A1(new_n5204_), .B0(new_n5207_), .B1(new_n5206_), .Y(new_n5209_));
  AND2X1   g04207(.A(\A[857] ), .B(\A[856] ), .Y(new_n5210_));
  AOI21X1  g04208(.A0(new_n5208_), .A1(\A[858] ), .B0(new_n5210_), .Y(new_n5211_));
  AND2X1   g04209(.A(\A[854] ), .B(\A[853] ), .Y(new_n5212_));
  AOI21X1  g04210(.A0(new_n5201_), .A1(\A[855] ), .B0(new_n5212_), .Y(new_n5213_));
  XOR2X1   g04211(.A(new_n5209_), .B(new_n5203_), .Y(new_n5214_));
  INVX1    g04212(.A(\A[847] ), .Y(new_n5215_));
  OR2X1    g04213(.A(\A[848] ), .B(new_n5215_), .Y(new_n5216_));
  INVX1    g04214(.A(\A[849] ), .Y(new_n5217_));
  AOI21X1  g04215(.A0(\A[848] ), .A1(new_n5215_), .B0(new_n5217_), .Y(new_n5218_));
  XOR2X1   g04216(.A(\A[848] ), .B(\A[847] ), .Y(new_n5219_));
  AND2X1   g04217(.A(new_n5219_), .B(new_n5217_), .Y(new_n5220_));
  AOI21X1  g04218(.A0(new_n5218_), .A1(new_n5216_), .B0(new_n5220_), .Y(new_n5221_));
  INVX1    g04219(.A(\A[852] ), .Y(new_n5222_));
  INVX1    g04220(.A(\A[850] ), .Y(new_n5223_));
  OR2X1    g04221(.A(\A[851] ), .B(new_n5223_), .Y(new_n5224_));
  AOI21X1  g04222(.A0(\A[851] ), .A1(new_n5223_), .B0(new_n5222_), .Y(new_n5225_));
  XOR2X1   g04223(.A(\A[851] ), .B(\A[850] ), .Y(new_n5226_));
  AOI22X1  g04224(.A0(new_n5226_), .A1(new_n5222_), .B0(new_n5225_), .B1(new_n5224_), .Y(new_n5227_));
  AND2X1   g04225(.A(\A[851] ), .B(\A[850] ), .Y(new_n5228_));
  AOI21X1  g04226(.A0(new_n5226_), .A1(\A[852] ), .B0(new_n5228_), .Y(new_n5229_));
  AND2X1   g04227(.A(\A[848] ), .B(\A[847] ), .Y(new_n5230_));
  AOI21X1  g04228(.A0(new_n5219_), .A1(\A[849] ), .B0(new_n5230_), .Y(new_n5231_));
  XOR2X1   g04229(.A(new_n5227_), .B(new_n5221_), .Y(new_n5232_));
  XOR2X1   g04230(.A(new_n5232_), .B(new_n5214_), .Y(new_n5233_));
  XOR2X1   g04231(.A(new_n5233_), .B(new_n5195_), .Y(new_n5234_));
  XOR2X1   g04232(.A(new_n5234_), .B(new_n5157_), .Y(new_n5235_));
  XOR2X1   g04233(.A(new_n5235_), .B(new_n5081_), .Y(new_n5236_));
  NAND2X1  g04234(.A(new_n5236_), .B(new_n4927_), .Y(new_n5237_));
  NOR3X1   g04235(.A(new_n5237_), .B(new_n4923_), .C(new_n4919_), .Y(new_n5238_));
  MX2X1    g04236(.A(new_n4184_), .B(new_n4090_), .S0(new_n4179_), .Y(new_n5239_));
  NOR3X1   g04237(.A(new_n4920_), .B(new_n4892_), .C(new_n4878_), .Y(new_n5240_));
  MX2X1    g04238(.A(new_n4891_), .B(new_n4877_), .S0(new_n4483_), .Y(new_n5241_));
  AND2X1   g04239(.A(new_n5241_), .B(new_n4920_), .Y(new_n5242_));
  OAI21X1  g04240(.A0(new_n5242_), .A1(new_n5240_), .B0(new_n5239_), .Y(new_n5243_));
  OR2X1    g04241(.A(new_n4914_), .B(new_n4888_), .Y(new_n5244_));
  AOI21X1  g04242(.A0(new_n4891_), .A1(new_n4888_), .B0(new_n4897_), .Y(new_n5245_));
  AOI22X1  g04243(.A0(new_n5245_), .A1(new_n5244_), .B0(new_n5241_), .B1(new_n4897_), .Y(new_n5246_));
  OR2X1    g04244(.A(new_n5246_), .B(new_n5239_), .Y(new_n5247_));
  AND2X1   g04245(.A(new_n5236_), .B(new_n4927_), .Y(new_n5248_));
  AOI21X1  g04246(.A0(new_n5247_), .A1(new_n5243_), .B0(new_n5248_), .Y(new_n5249_));
  AND2X1   g04247(.A(new_n5141_), .B(new_n5139_), .Y(new_n5250_));
  OR2X1    g04248(.A(new_n5143_), .B(new_n5250_), .Y(new_n5251_));
  XOR2X1   g04249(.A(new_n5150_), .B(new_n5251_), .Y(new_n5252_));
  XOR2X1   g04250(.A(new_n5154_), .B(new_n5152_), .Y(new_n5253_));
  NOR2X1   g04251(.A(new_n5150_), .B(new_n5144_), .Y(new_n5254_));
  NOR2X1   g04252(.A(new_n5154_), .B(new_n5152_), .Y(new_n5255_));
  AOI21X1  g04253(.A0(new_n5254_), .A1(new_n5253_), .B0(new_n5255_), .Y(new_n5256_));
  XOR2X1   g04254(.A(new_n5254_), .B(new_n5253_), .Y(new_n5257_));
  OAI21X1  g04255(.A0(new_n5256_), .A1(new_n5252_), .B0(new_n5257_), .Y(new_n5258_));
  INVX1    g04256(.A(new_n5258_), .Y(new_n5259_));
  XOR2X1   g04257(.A(new_n5132_), .B(new_n5126_), .Y(new_n5260_));
  AOI21X1  g04258(.A0(new_n5122_), .A1(new_n5120_), .B0(new_n5125_), .Y(new_n5261_));
  NOR4X1   g04259(.A(new_n5136_), .B(new_n5134_), .C(new_n5132_), .D(new_n5261_), .Y(new_n5262_));
  NOR4X1   g04260(.A(new_n5154_), .B(new_n5152_), .C(new_n5150_), .D(new_n5144_), .Y(new_n5263_));
  OR4X1    g04261(.A(new_n5263_), .B(new_n5252_), .C(new_n5262_), .D(new_n5260_), .Y(new_n5264_));
  XOR2X1   g04262(.A(new_n5136_), .B(new_n5134_), .Y(new_n5265_));
  NOR2X1   g04263(.A(new_n5132_), .B(new_n5261_), .Y(new_n5266_));
  NOR2X1   g04264(.A(new_n5136_), .B(new_n5134_), .Y(new_n5267_));
  AOI21X1  g04265(.A0(new_n5266_), .A1(new_n5265_), .B0(new_n5267_), .Y(new_n5268_));
  XOR2X1   g04266(.A(new_n5266_), .B(new_n5265_), .Y(new_n5269_));
  OAI21X1  g04267(.A0(new_n5268_), .A1(new_n5260_), .B0(new_n5269_), .Y(new_n5270_));
  XOR2X1   g04268(.A(new_n5270_), .B(new_n5264_), .Y(new_n5271_));
  AND2X1   g04269(.A(new_n5271_), .B(new_n5258_), .Y(new_n5272_));
  AND2X1   g04270(.A(new_n5270_), .B(new_n5264_), .Y(new_n5273_));
  OR2X1    g04271(.A(new_n5132_), .B(new_n5261_), .Y(new_n5274_));
  XOR2X1   g04272(.A(new_n5274_), .B(new_n5265_), .Y(new_n5275_));
  OR4X1    g04273(.A(new_n5252_), .B(new_n5262_), .C(new_n5275_), .D(new_n5260_), .Y(new_n5276_));
  OR4X1    g04274(.A(new_n5154_), .B(new_n5152_), .C(new_n5150_), .D(new_n5144_), .Y(new_n5277_));
  OAI21X1  g04275(.A0(new_n5268_), .A1(new_n5260_), .B0(new_n5277_), .Y(new_n5278_));
  NOR2X1   g04276(.A(new_n5278_), .B(new_n5276_), .Y(new_n5279_));
  OR2X1    g04277(.A(new_n5279_), .B(new_n5273_), .Y(new_n5280_));
  AOI21X1  g04278(.A0(new_n5280_), .A1(new_n5259_), .B0(new_n5272_), .Y(new_n5281_));
  AND2X1   g04279(.A(new_n5103_), .B(new_n5101_), .Y(new_n5282_));
  OR2X1    g04280(.A(new_n5105_), .B(new_n5282_), .Y(new_n5283_));
  XOR2X1   g04281(.A(new_n5112_), .B(new_n5283_), .Y(new_n5284_));
  XOR2X1   g04282(.A(new_n5116_), .B(new_n5114_), .Y(new_n5285_));
  NOR2X1   g04283(.A(new_n5112_), .B(new_n5106_), .Y(new_n5286_));
  NOR2X1   g04284(.A(new_n5116_), .B(new_n5114_), .Y(new_n5287_));
  AOI21X1  g04285(.A0(new_n5286_), .A1(new_n5285_), .B0(new_n5287_), .Y(new_n5288_));
  XOR2X1   g04286(.A(new_n5286_), .B(new_n5285_), .Y(new_n5289_));
  OAI21X1  g04287(.A0(new_n5288_), .A1(new_n5284_), .B0(new_n5289_), .Y(new_n5290_));
  AND2X1   g04288(.A(new_n5085_), .B(new_n5083_), .Y(new_n5291_));
  OR2X1    g04289(.A(new_n5087_), .B(new_n5291_), .Y(new_n5292_));
  XOR2X1   g04290(.A(new_n5094_), .B(new_n5292_), .Y(new_n5293_));
  NOR4X1   g04291(.A(new_n5098_), .B(new_n5096_), .C(new_n5094_), .D(new_n5088_), .Y(new_n5294_));
  NOR4X1   g04292(.A(new_n5116_), .B(new_n5114_), .C(new_n5112_), .D(new_n5106_), .Y(new_n5295_));
  OR4X1    g04293(.A(new_n5295_), .B(new_n5284_), .C(new_n5294_), .D(new_n5293_), .Y(new_n5296_));
  XOR2X1   g04294(.A(new_n5098_), .B(new_n5096_), .Y(new_n5297_));
  NOR2X1   g04295(.A(new_n5094_), .B(new_n5088_), .Y(new_n5298_));
  NOR2X1   g04296(.A(new_n5098_), .B(new_n5096_), .Y(new_n5299_));
  AOI21X1  g04297(.A0(new_n5298_), .A1(new_n5297_), .B0(new_n5299_), .Y(new_n5300_));
  XOR2X1   g04298(.A(new_n5298_), .B(new_n5297_), .Y(new_n5301_));
  OAI21X1  g04299(.A0(new_n5300_), .A1(new_n5293_), .B0(new_n5301_), .Y(new_n5302_));
  XOR2X1   g04300(.A(new_n5302_), .B(new_n5296_), .Y(new_n5303_));
  AND2X1   g04301(.A(new_n5303_), .B(new_n5290_), .Y(new_n5304_));
  NAND2X1  g04302(.A(new_n5302_), .B(new_n5296_), .Y(new_n5305_));
  OR2X1    g04303(.A(new_n5094_), .B(new_n5088_), .Y(new_n5306_));
  XOR2X1   g04304(.A(new_n5306_), .B(new_n5297_), .Y(new_n5307_));
  OR4X1    g04305(.A(new_n5284_), .B(new_n5294_), .C(new_n5307_), .D(new_n5293_), .Y(new_n5308_));
  AND2X1   g04306(.A(new_n5111_), .B(\A[888] ), .Y(new_n5309_));
  OR2X1    g04307(.A(new_n5309_), .B(new_n5113_), .Y(new_n5310_));
  XOR2X1   g04308(.A(new_n5116_), .B(new_n5310_), .Y(new_n5311_));
  XOR2X1   g04309(.A(new_n5286_), .B(new_n5311_), .Y(new_n5312_));
  OAI22X1  g04310(.A0(new_n5312_), .A1(new_n5288_), .B0(new_n5300_), .B1(new_n5293_), .Y(new_n5313_));
  OR2X1    g04311(.A(new_n5313_), .B(new_n5308_), .Y(new_n5314_));
  AOI21X1  g04312(.A0(new_n5314_), .A1(new_n5305_), .B0(new_n5290_), .Y(new_n5315_));
  INVX1    g04313(.A(new_n5118_), .Y(new_n5316_));
  OR2X1    g04314(.A(new_n5156_), .B(new_n5316_), .Y(new_n5317_));
  NOR3X1   g04315(.A(new_n5317_), .B(new_n5315_), .C(new_n5304_), .Y(new_n5318_));
  NAND2X1  g04316(.A(new_n5303_), .B(new_n5290_), .Y(new_n5319_));
  XOR2X1   g04317(.A(new_n5112_), .B(new_n5106_), .Y(new_n5320_));
  OR2X1    g04318(.A(new_n5112_), .B(new_n5106_), .Y(new_n5321_));
  OR2X1    g04319(.A(new_n5116_), .B(new_n5114_), .Y(new_n5322_));
  OAI21X1  g04320(.A0(new_n5321_), .A1(new_n5311_), .B0(new_n5322_), .Y(new_n5323_));
  AOI21X1  g04321(.A0(new_n5323_), .A1(new_n5320_), .B0(new_n5312_), .Y(new_n5324_));
  AND2X1   g04322(.A(new_n5302_), .B(new_n5296_), .Y(new_n5325_));
  NOR2X1   g04323(.A(new_n5313_), .B(new_n5308_), .Y(new_n5326_));
  OAI21X1  g04324(.A0(new_n5326_), .A1(new_n5325_), .B0(new_n5324_), .Y(new_n5327_));
  NOR2X1   g04325(.A(new_n5156_), .B(new_n5316_), .Y(new_n5328_));
  AOI21X1  g04326(.A0(new_n5327_), .A1(new_n5319_), .B0(new_n5328_), .Y(new_n5329_));
  OAI21X1  g04327(.A0(new_n5329_), .A1(new_n5318_), .B0(new_n5281_), .Y(new_n5330_));
  MX2X1    g04328(.A(new_n5280_), .B(new_n5271_), .S0(new_n5258_), .Y(new_n5331_));
  NOR3X1   g04329(.A(new_n5328_), .B(new_n5315_), .C(new_n5304_), .Y(new_n5332_));
  AOI21X1  g04330(.A0(new_n5327_), .A1(new_n5319_), .B0(new_n5317_), .Y(new_n5333_));
  OAI21X1  g04331(.A0(new_n5333_), .A1(new_n5332_), .B0(new_n5331_), .Y(new_n5334_));
  XOR2X1   g04332(.A(new_n5233_), .B(new_n5194_), .Y(new_n5335_));
  NOR2X1   g04333(.A(new_n5335_), .B(new_n5157_), .Y(new_n5336_));
  NAND3X1  g04334(.A(new_n5336_), .B(new_n5334_), .C(new_n5330_), .Y(new_n5337_));
  NAND3X1  g04335(.A(new_n5328_), .B(new_n5327_), .C(new_n5319_), .Y(new_n5338_));
  OAI21X1  g04336(.A0(new_n5315_), .A1(new_n5304_), .B0(new_n5317_), .Y(new_n5339_));
  AOI21X1  g04337(.A0(new_n5339_), .A1(new_n5338_), .B0(new_n5331_), .Y(new_n5340_));
  NAND3X1  g04338(.A(new_n5317_), .B(new_n5327_), .C(new_n5319_), .Y(new_n5341_));
  OAI21X1  g04339(.A0(new_n5315_), .A1(new_n5304_), .B0(new_n5328_), .Y(new_n5342_));
  AOI21X1  g04340(.A0(new_n5342_), .A1(new_n5341_), .B0(new_n5281_), .Y(new_n5343_));
  INVX1    g04341(.A(new_n5336_), .Y(new_n5344_));
  OAI21X1  g04342(.A0(new_n5343_), .A1(new_n5340_), .B0(new_n5344_), .Y(new_n5345_));
  AND2X1   g04343(.A(new_n5345_), .B(new_n5337_), .Y(new_n5346_));
  AND2X1   g04344(.A(new_n5179_), .B(new_n5177_), .Y(new_n5347_));
  OR2X1    g04345(.A(new_n5181_), .B(new_n5347_), .Y(new_n5348_));
  XOR2X1   g04346(.A(new_n5188_), .B(new_n5348_), .Y(new_n5349_));
  XOR2X1   g04347(.A(new_n5192_), .B(new_n5190_), .Y(new_n5350_));
  NOR2X1   g04348(.A(new_n5188_), .B(new_n5182_), .Y(new_n5351_));
  NOR2X1   g04349(.A(new_n5192_), .B(new_n5190_), .Y(new_n5352_));
  AOI21X1  g04350(.A0(new_n5351_), .A1(new_n5350_), .B0(new_n5352_), .Y(new_n5353_));
  XOR2X1   g04351(.A(new_n5351_), .B(new_n5350_), .Y(new_n5354_));
  OAI21X1  g04352(.A0(new_n5353_), .A1(new_n5349_), .B0(new_n5354_), .Y(new_n5355_));
  AND2X1   g04353(.A(new_n5161_), .B(new_n5159_), .Y(new_n5356_));
  OR2X1    g04354(.A(new_n5163_), .B(new_n5356_), .Y(new_n5357_));
  XOR2X1   g04355(.A(new_n5170_), .B(new_n5357_), .Y(new_n5358_));
  NOR4X1   g04356(.A(new_n5174_), .B(new_n5172_), .C(new_n5170_), .D(new_n5164_), .Y(new_n5359_));
  NOR4X1   g04357(.A(new_n5192_), .B(new_n5190_), .C(new_n5188_), .D(new_n5182_), .Y(new_n5360_));
  OR4X1    g04358(.A(new_n5360_), .B(new_n5349_), .C(new_n5359_), .D(new_n5358_), .Y(new_n5361_));
  XOR2X1   g04359(.A(new_n5174_), .B(new_n5172_), .Y(new_n5362_));
  NOR2X1   g04360(.A(new_n5170_), .B(new_n5164_), .Y(new_n5363_));
  NOR2X1   g04361(.A(new_n5174_), .B(new_n5172_), .Y(new_n5364_));
  AOI21X1  g04362(.A0(new_n5363_), .A1(new_n5362_), .B0(new_n5364_), .Y(new_n5365_));
  XOR2X1   g04363(.A(new_n5363_), .B(new_n5362_), .Y(new_n5366_));
  OAI21X1  g04364(.A0(new_n5365_), .A1(new_n5358_), .B0(new_n5366_), .Y(new_n5367_));
  XOR2X1   g04365(.A(new_n5367_), .B(new_n5361_), .Y(new_n5368_));
  NAND2X1  g04366(.A(new_n5368_), .B(new_n5355_), .Y(new_n5369_));
  XOR2X1   g04367(.A(new_n5188_), .B(new_n5182_), .Y(new_n5370_));
  AND2X1   g04368(.A(new_n5187_), .B(\A[864] ), .Y(new_n5371_));
  OR2X1    g04369(.A(new_n5371_), .B(new_n5189_), .Y(new_n5372_));
  XOR2X1   g04370(.A(new_n5192_), .B(new_n5372_), .Y(new_n5373_));
  OR2X1    g04371(.A(new_n5188_), .B(new_n5182_), .Y(new_n5374_));
  OR2X1    g04372(.A(new_n5192_), .B(new_n5190_), .Y(new_n5375_));
  OAI21X1  g04373(.A0(new_n5374_), .A1(new_n5373_), .B0(new_n5375_), .Y(new_n5376_));
  XOR2X1   g04374(.A(new_n5351_), .B(new_n5373_), .Y(new_n5377_));
  AOI21X1  g04375(.A0(new_n5376_), .A1(new_n5370_), .B0(new_n5377_), .Y(new_n5378_));
  AND2X1   g04376(.A(new_n5367_), .B(new_n5361_), .Y(new_n5379_));
  OR2X1    g04377(.A(new_n5170_), .B(new_n5164_), .Y(new_n5380_));
  XOR2X1   g04378(.A(new_n5380_), .B(new_n5362_), .Y(new_n5381_));
  OR4X1    g04379(.A(new_n5349_), .B(new_n5359_), .C(new_n5381_), .D(new_n5358_), .Y(new_n5382_));
  OAI22X1  g04380(.A0(new_n5377_), .A1(new_n5353_), .B0(new_n5365_), .B1(new_n5358_), .Y(new_n5383_));
  NOR2X1   g04381(.A(new_n5383_), .B(new_n5382_), .Y(new_n5384_));
  OAI21X1  g04382(.A0(new_n5384_), .A1(new_n5379_), .B0(new_n5378_), .Y(new_n5385_));
  NOR2X1   g04383(.A(new_n5233_), .B(new_n5195_), .Y(new_n5386_));
  NAND3X1  g04384(.A(new_n5386_), .B(new_n5385_), .C(new_n5369_), .Y(new_n5387_));
  AND2X1   g04385(.A(new_n5368_), .B(new_n5355_), .Y(new_n5388_));
  NAND2X1  g04386(.A(new_n5367_), .B(new_n5361_), .Y(new_n5389_));
  OR2X1    g04387(.A(new_n5383_), .B(new_n5382_), .Y(new_n5390_));
  AOI21X1  g04388(.A0(new_n5390_), .A1(new_n5389_), .B0(new_n5355_), .Y(new_n5391_));
  OR2X1    g04389(.A(new_n5233_), .B(new_n5195_), .Y(new_n5392_));
  OAI21X1  g04390(.A0(new_n5391_), .A1(new_n5388_), .B0(new_n5392_), .Y(new_n5393_));
  AND2X1   g04391(.A(new_n5218_), .B(new_n5216_), .Y(new_n5394_));
  OR2X1    g04392(.A(new_n5220_), .B(new_n5394_), .Y(new_n5395_));
  XOR2X1   g04393(.A(new_n5227_), .B(new_n5395_), .Y(new_n5396_));
  XOR2X1   g04394(.A(new_n5231_), .B(new_n5229_), .Y(new_n5397_));
  NOR2X1   g04395(.A(new_n5227_), .B(new_n5221_), .Y(new_n5398_));
  NOR2X1   g04396(.A(new_n5231_), .B(new_n5229_), .Y(new_n5399_));
  AOI21X1  g04397(.A0(new_n5398_), .A1(new_n5397_), .B0(new_n5399_), .Y(new_n5400_));
  XOR2X1   g04398(.A(new_n5398_), .B(new_n5397_), .Y(new_n5401_));
  OAI21X1  g04399(.A0(new_n5400_), .A1(new_n5396_), .B0(new_n5401_), .Y(new_n5402_));
  XOR2X1   g04400(.A(new_n5209_), .B(new_n5203_), .Y(new_n5403_));
  AOI21X1  g04401(.A0(new_n5199_), .A1(new_n5197_), .B0(new_n5202_), .Y(new_n5404_));
  NOR4X1   g04402(.A(new_n5213_), .B(new_n5211_), .C(new_n5209_), .D(new_n5404_), .Y(new_n5405_));
  NOR4X1   g04403(.A(new_n5231_), .B(new_n5229_), .C(new_n5227_), .D(new_n5221_), .Y(new_n5406_));
  OR4X1    g04404(.A(new_n5406_), .B(new_n5396_), .C(new_n5405_), .D(new_n5403_), .Y(new_n5407_));
  XOR2X1   g04405(.A(new_n5213_), .B(new_n5211_), .Y(new_n5408_));
  NOR2X1   g04406(.A(new_n5209_), .B(new_n5404_), .Y(new_n5409_));
  NOR2X1   g04407(.A(new_n5213_), .B(new_n5211_), .Y(new_n5410_));
  AOI21X1  g04408(.A0(new_n5409_), .A1(new_n5408_), .B0(new_n5410_), .Y(new_n5411_));
  XOR2X1   g04409(.A(new_n5409_), .B(new_n5408_), .Y(new_n5412_));
  OAI21X1  g04410(.A0(new_n5411_), .A1(new_n5403_), .B0(new_n5412_), .Y(new_n5413_));
  XOR2X1   g04411(.A(new_n5413_), .B(new_n5407_), .Y(new_n5414_));
  AND2X1   g04412(.A(new_n5413_), .B(new_n5407_), .Y(new_n5415_));
  OR2X1    g04413(.A(new_n5209_), .B(new_n5404_), .Y(new_n5416_));
  XOR2X1   g04414(.A(new_n5416_), .B(new_n5408_), .Y(new_n5417_));
  OR4X1    g04415(.A(new_n5396_), .B(new_n5405_), .C(new_n5417_), .D(new_n5403_), .Y(new_n5418_));
  OR4X1    g04416(.A(new_n5231_), .B(new_n5229_), .C(new_n5227_), .D(new_n5221_), .Y(new_n5419_));
  OAI21X1  g04417(.A0(new_n5411_), .A1(new_n5403_), .B0(new_n5419_), .Y(new_n5420_));
  NOR2X1   g04418(.A(new_n5420_), .B(new_n5418_), .Y(new_n5421_));
  OR2X1    g04419(.A(new_n5421_), .B(new_n5415_), .Y(new_n5422_));
  MX2X1    g04420(.A(new_n5422_), .B(new_n5414_), .S0(new_n5402_), .Y(new_n5423_));
  AOI21X1  g04421(.A0(new_n5393_), .A1(new_n5387_), .B0(new_n5423_), .Y(new_n5424_));
  INVX1    g04422(.A(new_n5402_), .Y(new_n5425_));
  AND2X1   g04423(.A(new_n5414_), .B(new_n5402_), .Y(new_n5426_));
  AOI21X1  g04424(.A0(new_n5422_), .A1(new_n5425_), .B0(new_n5426_), .Y(new_n5427_));
  NAND3X1  g04425(.A(new_n5392_), .B(new_n5385_), .C(new_n5369_), .Y(new_n5428_));
  OAI21X1  g04426(.A0(new_n5391_), .A1(new_n5388_), .B0(new_n5386_), .Y(new_n5429_));
  AOI21X1  g04427(.A0(new_n5429_), .A1(new_n5428_), .B0(new_n5427_), .Y(new_n5430_));
  OR2X1    g04428(.A(new_n5430_), .B(new_n5424_), .Y(new_n5431_));
  NOR3X1   g04429(.A(new_n5336_), .B(new_n5343_), .C(new_n5340_), .Y(new_n5432_));
  AOI21X1  g04430(.A0(new_n5334_), .A1(new_n5330_), .B0(new_n5344_), .Y(new_n5433_));
  OAI21X1  g04431(.A0(new_n5433_), .A1(new_n5432_), .B0(new_n5431_), .Y(new_n5434_));
  OAI21X1  g04432(.A0(new_n5431_), .A1(new_n5346_), .B0(new_n5434_), .Y(new_n5435_));
  AND2X1   g04433(.A(new_n5025_), .B(new_n5023_), .Y(new_n5436_));
  OR2X1    g04434(.A(new_n5027_), .B(new_n5436_), .Y(new_n5437_));
  XOR2X1   g04435(.A(new_n5034_), .B(new_n5437_), .Y(new_n5438_));
  XOR2X1   g04436(.A(new_n5038_), .B(new_n5036_), .Y(new_n5439_));
  NOR2X1   g04437(.A(new_n5034_), .B(new_n5028_), .Y(new_n5440_));
  NOR2X1   g04438(.A(new_n5038_), .B(new_n5036_), .Y(new_n5441_));
  AOI21X1  g04439(.A0(new_n5440_), .A1(new_n5439_), .B0(new_n5441_), .Y(new_n5442_));
  XOR2X1   g04440(.A(new_n5440_), .B(new_n5439_), .Y(new_n5443_));
  OAI21X1  g04441(.A0(new_n5442_), .A1(new_n5438_), .B0(new_n5443_), .Y(new_n5444_));
  AND2X1   g04442(.A(new_n5007_), .B(new_n5005_), .Y(new_n5445_));
  OR2X1    g04443(.A(new_n5009_), .B(new_n5445_), .Y(new_n5446_));
  XOR2X1   g04444(.A(new_n5016_), .B(new_n5446_), .Y(new_n5447_));
  NOR4X1   g04445(.A(new_n5020_), .B(new_n5018_), .C(new_n5016_), .D(new_n5010_), .Y(new_n5448_));
  NOR4X1   g04446(.A(new_n5038_), .B(new_n5036_), .C(new_n5034_), .D(new_n5028_), .Y(new_n5449_));
  OR4X1    g04447(.A(new_n5449_), .B(new_n5438_), .C(new_n5448_), .D(new_n5447_), .Y(new_n5450_));
  XOR2X1   g04448(.A(new_n5020_), .B(new_n5018_), .Y(new_n5451_));
  NOR2X1   g04449(.A(new_n5016_), .B(new_n5010_), .Y(new_n5452_));
  NOR2X1   g04450(.A(new_n5020_), .B(new_n5018_), .Y(new_n5453_));
  AOI21X1  g04451(.A0(new_n5452_), .A1(new_n5451_), .B0(new_n5453_), .Y(new_n5454_));
  XOR2X1   g04452(.A(new_n5452_), .B(new_n5451_), .Y(new_n5455_));
  OAI21X1  g04453(.A0(new_n5454_), .A1(new_n5447_), .B0(new_n5455_), .Y(new_n5456_));
  XOR2X1   g04454(.A(new_n5456_), .B(new_n5450_), .Y(new_n5457_));
  NAND2X1  g04455(.A(new_n5457_), .B(new_n5444_), .Y(new_n5458_));
  XOR2X1   g04456(.A(new_n5034_), .B(new_n5028_), .Y(new_n5459_));
  AND2X1   g04457(.A(new_n5033_), .B(\A[912] ), .Y(new_n5460_));
  OR2X1    g04458(.A(new_n5460_), .B(new_n5035_), .Y(new_n5461_));
  XOR2X1   g04459(.A(new_n5038_), .B(new_n5461_), .Y(new_n5462_));
  OR2X1    g04460(.A(new_n5034_), .B(new_n5028_), .Y(new_n5463_));
  OR2X1    g04461(.A(new_n5038_), .B(new_n5036_), .Y(new_n5464_));
  OAI21X1  g04462(.A0(new_n5463_), .A1(new_n5462_), .B0(new_n5464_), .Y(new_n5465_));
  XOR2X1   g04463(.A(new_n5440_), .B(new_n5462_), .Y(new_n5466_));
  AOI21X1  g04464(.A0(new_n5465_), .A1(new_n5459_), .B0(new_n5466_), .Y(new_n5467_));
  AND2X1   g04465(.A(new_n5456_), .B(new_n5450_), .Y(new_n5468_));
  OR2X1    g04466(.A(new_n5016_), .B(new_n5010_), .Y(new_n5469_));
  XOR2X1   g04467(.A(new_n5469_), .B(new_n5451_), .Y(new_n5470_));
  OR4X1    g04468(.A(new_n5438_), .B(new_n5448_), .C(new_n5470_), .D(new_n5447_), .Y(new_n5471_));
  OAI22X1  g04469(.A0(new_n5466_), .A1(new_n5442_), .B0(new_n5454_), .B1(new_n5447_), .Y(new_n5472_));
  NOR2X1   g04470(.A(new_n5472_), .B(new_n5471_), .Y(new_n5473_));
  OAI21X1  g04471(.A0(new_n5473_), .A1(new_n5468_), .B0(new_n5467_), .Y(new_n5474_));
  NOR2X1   g04472(.A(new_n5079_), .B(new_n5041_), .Y(new_n5475_));
  NAND3X1  g04473(.A(new_n5475_), .B(new_n5474_), .C(new_n5458_), .Y(new_n5476_));
  AND2X1   g04474(.A(new_n5457_), .B(new_n5444_), .Y(new_n5477_));
  NAND2X1  g04475(.A(new_n5456_), .B(new_n5450_), .Y(new_n5478_));
  OR2X1    g04476(.A(new_n5472_), .B(new_n5471_), .Y(new_n5479_));
  AOI21X1  g04477(.A0(new_n5479_), .A1(new_n5478_), .B0(new_n5444_), .Y(new_n5480_));
  OR2X1    g04478(.A(new_n5079_), .B(new_n5041_), .Y(new_n5481_));
  OAI21X1  g04479(.A0(new_n5480_), .A1(new_n5477_), .B0(new_n5481_), .Y(new_n5482_));
  AND2X1   g04480(.A(new_n5064_), .B(new_n5062_), .Y(new_n5483_));
  OR2X1    g04481(.A(new_n5066_), .B(new_n5483_), .Y(new_n5484_));
  XOR2X1   g04482(.A(new_n5073_), .B(new_n5484_), .Y(new_n5485_));
  XOR2X1   g04483(.A(new_n5077_), .B(new_n5075_), .Y(new_n5486_));
  NOR2X1   g04484(.A(new_n5073_), .B(new_n5067_), .Y(new_n5487_));
  NOR2X1   g04485(.A(new_n5077_), .B(new_n5075_), .Y(new_n5488_));
  AOI21X1  g04486(.A0(new_n5487_), .A1(new_n5486_), .B0(new_n5488_), .Y(new_n5489_));
  XOR2X1   g04487(.A(new_n5487_), .B(new_n5486_), .Y(new_n5490_));
  OAI21X1  g04488(.A0(new_n5489_), .A1(new_n5485_), .B0(new_n5490_), .Y(new_n5491_));
  XOR2X1   g04489(.A(new_n5055_), .B(new_n5049_), .Y(new_n5492_));
  AOI21X1  g04490(.A0(new_n5045_), .A1(new_n5043_), .B0(new_n5048_), .Y(new_n5493_));
  NOR4X1   g04491(.A(new_n5059_), .B(new_n5057_), .C(new_n5055_), .D(new_n5493_), .Y(new_n5494_));
  NOR4X1   g04492(.A(new_n5077_), .B(new_n5075_), .C(new_n5073_), .D(new_n5067_), .Y(new_n5495_));
  OR4X1    g04493(.A(new_n5495_), .B(new_n5485_), .C(new_n5494_), .D(new_n5492_), .Y(new_n5496_));
  XOR2X1   g04494(.A(new_n5059_), .B(new_n5057_), .Y(new_n5497_));
  NOR2X1   g04495(.A(new_n5055_), .B(new_n5493_), .Y(new_n5498_));
  NOR2X1   g04496(.A(new_n5059_), .B(new_n5057_), .Y(new_n5499_));
  AOI21X1  g04497(.A0(new_n5498_), .A1(new_n5497_), .B0(new_n5499_), .Y(new_n5500_));
  XOR2X1   g04498(.A(new_n5498_), .B(new_n5497_), .Y(new_n5501_));
  OAI21X1  g04499(.A0(new_n5500_), .A1(new_n5492_), .B0(new_n5501_), .Y(new_n5502_));
  XOR2X1   g04500(.A(new_n5502_), .B(new_n5496_), .Y(new_n5503_));
  AND2X1   g04501(.A(new_n5502_), .B(new_n5496_), .Y(new_n5504_));
  OR2X1    g04502(.A(new_n5055_), .B(new_n5493_), .Y(new_n5505_));
  XOR2X1   g04503(.A(new_n5505_), .B(new_n5497_), .Y(new_n5506_));
  OR4X1    g04504(.A(new_n5485_), .B(new_n5494_), .C(new_n5506_), .D(new_n5492_), .Y(new_n5507_));
  OR4X1    g04505(.A(new_n5077_), .B(new_n5075_), .C(new_n5073_), .D(new_n5067_), .Y(new_n5508_));
  OAI21X1  g04506(.A0(new_n5500_), .A1(new_n5492_), .B0(new_n5508_), .Y(new_n5509_));
  NOR2X1   g04507(.A(new_n5509_), .B(new_n5507_), .Y(new_n5510_));
  OR2X1    g04508(.A(new_n5510_), .B(new_n5504_), .Y(new_n5511_));
  MX2X1    g04509(.A(new_n5511_), .B(new_n5503_), .S0(new_n5491_), .Y(new_n5512_));
  AOI21X1  g04510(.A0(new_n5482_), .A1(new_n5476_), .B0(new_n5512_), .Y(new_n5513_));
  INVX1    g04511(.A(new_n5491_), .Y(new_n5514_));
  AND2X1   g04512(.A(new_n5503_), .B(new_n5491_), .Y(new_n5515_));
  AOI21X1  g04513(.A0(new_n5511_), .A1(new_n5514_), .B0(new_n5515_), .Y(new_n5516_));
  NAND3X1  g04514(.A(new_n5481_), .B(new_n5474_), .C(new_n5458_), .Y(new_n5517_));
  OAI21X1  g04515(.A0(new_n5480_), .A1(new_n5477_), .B0(new_n5475_), .Y(new_n5518_));
  AOI21X1  g04516(.A0(new_n5518_), .A1(new_n5517_), .B0(new_n5516_), .Y(new_n5519_));
  OR2X1    g04517(.A(new_n5519_), .B(new_n5513_), .Y(new_n5520_));
  AND2X1   g04518(.A(new_n4987_), .B(new_n4985_), .Y(new_n5521_));
  OR2X1    g04519(.A(new_n4989_), .B(new_n5521_), .Y(new_n5522_));
  XOR2X1   g04520(.A(new_n4996_), .B(new_n5522_), .Y(new_n5523_));
  XOR2X1   g04521(.A(new_n5000_), .B(new_n4998_), .Y(new_n5524_));
  NOR2X1   g04522(.A(new_n4996_), .B(new_n4990_), .Y(new_n5525_));
  NOR2X1   g04523(.A(new_n5000_), .B(new_n4998_), .Y(new_n5526_));
  AOI21X1  g04524(.A0(new_n5525_), .A1(new_n5524_), .B0(new_n5526_), .Y(new_n5527_));
  XOR2X1   g04525(.A(new_n5525_), .B(new_n5524_), .Y(new_n5528_));
  OAI21X1  g04526(.A0(new_n5527_), .A1(new_n5523_), .B0(new_n5528_), .Y(new_n5529_));
  INVX1    g04527(.A(new_n5529_), .Y(new_n5530_));
  XOR2X1   g04528(.A(new_n4978_), .B(new_n4972_), .Y(new_n5531_));
  AOI21X1  g04529(.A0(new_n4968_), .A1(new_n4966_), .B0(new_n4971_), .Y(new_n5532_));
  NOR4X1   g04530(.A(new_n4982_), .B(new_n4980_), .C(new_n4978_), .D(new_n5532_), .Y(new_n5533_));
  NOR4X1   g04531(.A(new_n5000_), .B(new_n4998_), .C(new_n4996_), .D(new_n4990_), .Y(new_n5534_));
  OR4X1    g04532(.A(new_n5534_), .B(new_n5523_), .C(new_n5533_), .D(new_n5531_), .Y(new_n5535_));
  XOR2X1   g04533(.A(new_n4982_), .B(new_n4980_), .Y(new_n5536_));
  NOR2X1   g04534(.A(new_n4978_), .B(new_n5532_), .Y(new_n5537_));
  NOR2X1   g04535(.A(new_n4982_), .B(new_n4980_), .Y(new_n5538_));
  AOI21X1  g04536(.A0(new_n5537_), .A1(new_n5536_), .B0(new_n5538_), .Y(new_n5539_));
  XOR2X1   g04537(.A(new_n5537_), .B(new_n5536_), .Y(new_n5540_));
  OAI21X1  g04538(.A0(new_n5539_), .A1(new_n5531_), .B0(new_n5540_), .Y(new_n5541_));
  XOR2X1   g04539(.A(new_n5541_), .B(new_n5535_), .Y(new_n5542_));
  AND2X1   g04540(.A(new_n5542_), .B(new_n5529_), .Y(new_n5543_));
  AND2X1   g04541(.A(new_n5541_), .B(new_n5535_), .Y(new_n5544_));
  OR2X1    g04542(.A(new_n4978_), .B(new_n5532_), .Y(new_n5545_));
  XOR2X1   g04543(.A(new_n5545_), .B(new_n5536_), .Y(new_n5546_));
  OR4X1    g04544(.A(new_n5523_), .B(new_n5533_), .C(new_n5546_), .D(new_n5531_), .Y(new_n5547_));
  OR4X1    g04545(.A(new_n5000_), .B(new_n4998_), .C(new_n4996_), .D(new_n4990_), .Y(new_n5548_));
  OAI21X1  g04546(.A0(new_n5539_), .A1(new_n5531_), .B0(new_n5548_), .Y(new_n5549_));
  NOR2X1   g04547(.A(new_n5549_), .B(new_n5547_), .Y(new_n5550_));
  OR2X1    g04548(.A(new_n5550_), .B(new_n5544_), .Y(new_n5551_));
  AOI21X1  g04549(.A0(new_n5551_), .A1(new_n5530_), .B0(new_n5543_), .Y(new_n5552_));
  AND2X1   g04550(.A(new_n4949_), .B(new_n4947_), .Y(new_n5553_));
  OR2X1    g04551(.A(new_n4951_), .B(new_n5553_), .Y(new_n5554_));
  XOR2X1   g04552(.A(new_n4958_), .B(new_n5554_), .Y(new_n5555_));
  XOR2X1   g04553(.A(new_n4962_), .B(new_n4960_), .Y(new_n5556_));
  NOR2X1   g04554(.A(new_n4958_), .B(new_n4952_), .Y(new_n5557_));
  NOR2X1   g04555(.A(new_n4962_), .B(new_n4960_), .Y(new_n5558_));
  AOI21X1  g04556(.A0(new_n5557_), .A1(new_n5556_), .B0(new_n5558_), .Y(new_n5559_));
  XOR2X1   g04557(.A(new_n5557_), .B(new_n5556_), .Y(new_n5560_));
  OAI21X1  g04558(.A0(new_n5559_), .A1(new_n5555_), .B0(new_n5560_), .Y(new_n5561_));
  AND2X1   g04559(.A(new_n4931_), .B(new_n4929_), .Y(new_n5562_));
  OR2X1    g04560(.A(new_n4933_), .B(new_n5562_), .Y(new_n5563_));
  XOR2X1   g04561(.A(new_n4940_), .B(new_n5563_), .Y(new_n5564_));
  NOR4X1   g04562(.A(new_n4944_), .B(new_n4942_), .C(new_n4940_), .D(new_n4934_), .Y(new_n5565_));
  NOR4X1   g04563(.A(new_n4962_), .B(new_n4960_), .C(new_n4958_), .D(new_n4952_), .Y(new_n5566_));
  OR4X1    g04564(.A(new_n5566_), .B(new_n5555_), .C(new_n5565_), .D(new_n5564_), .Y(new_n5567_));
  XOR2X1   g04565(.A(new_n4944_), .B(new_n4942_), .Y(new_n5568_));
  NOR2X1   g04566(.A(new_n4940_), .B(new_n4934_), .Y(new_n5569_));
  NOR2X1   g04567(.A(new_n4944_), .B(new_n4942_), .Y(new_n5570_));
  AOI21X1  g04568(.A0(new_n5569_), .A1(new_n5568_), .B0(new_n5570_), .Y(new_n5571_));
  XOR2X1   g04569(.A(new_n5569_), .B(new_n5568_), .Y(new_n5572_));
  OAI21X1  g04570(.A0(new_n5571_), .A1(new_n5564_), .B0(new_n5572_), .Y(new_n5573_));
  XOR2X1   g04571(.A(new_n5573_), .B(new_n5567_), .Y(new_n5574_));
  AND2X1   g04572(.A(new_n5574_), .B(new_n5561_), .Y(new_n5575_));
  NAND2X1  g04573(.A(new_n5573_), .B(new_n5567_), .Y(new_n5576_));
  OR2X1    g04574(.A(new_n4940_), .B(new_n4934_), .Y(new_n5577_));
  XOR2X1   g04575(.A(new_n5577_), .B(new_n5568_), .Y(new_n5578_));
  OR4X1    g04576(.A(new_n5555_), .B(new_n5565_), .C(new_n5578_), .D(new_n5564_), .Y(new_n5579_));
  AND2X1   g04577(.A(new_n4957_), .B(\A[936] ), .Y(new_n5580_));
  OR2X1    g04578(.A(new_n5580_), .B(new_n4959_), .Y(new_n5581_));
  XOR2X1   g04579(.A(new_n4962_), .B(new_n5581_), .Y(new_n5582_));
  XOR2X1   g04580(.A(new_n5557_), .B(new_n5582_), .Y(new_n5583_));
  OAI22X1  g04581(.A0(new_n5583_), .A1(new_n5559_), .B0(new_n5571_), .B1(new_n5564_), .Y(new_n5584_));
  OR2X1    g04582(.A(new_n5584_), .B(new_n5579_), .Y(new_n5585_));
  AOI21X1  g04583(.A0(new_n5585_), .A1(new_n5576_), .B0(new_n5561_), .Y(new_n5586_));
  INVX1    g04584(.A(new_n4964_), .Y(new_n5587_));
  OR2X1    g04585(.A(new_n5002_), .B(new_n5587_), .Y(new_n5588_));
  NOR3X1   g04586(.A(new_n5588_), .B(new_n5586_), .C(new_n5575_), .Y(new_n5589_));
  NAND2X1  g04587(.A(new_n5574_), .B(new_n5561_), .Y(new_n5590_));
  XOR2X1   g04588(.A(new_n4958_), .B(new_n4952_), .Y(new_n5591_));
  OR2X1    g04589(.A(new_n4958_), .B(new_n4952_), .Y(new_n5592_));
  OR2X1    g04590(.A(new_n4962_), .B(new_n4960_), .Y(new_n5593_));
  OAI21X1  g04591(.A0(new_n5592_), .A1(new_n5582_), .B0(new_n5593_), .Y(new_n5594_));
  AOI21X1  g04592(.A0(new_n5594_), .A1(new_n5591_), .B0(new_n5583_), .Y(new_n5595_));
  AND2X1   g04593(.A(new_n5573_), .B(new_n5567_), .Y(new_n5596_));
  NOR2X1   g04594(.A(new_n5584_), .B(new_n5579_), .Y(new_n5597_));
  OAI21X1  g04595(.A0(new_n5597_), .A1(new_n5596_), .B0(new_n5595_), .Y(new_n5598_));
  NOR2X1   g04596(.A(new_n5002_), .B(new_n5587_), .Y(new_n5599_));
  AOI21X1  g04597(.A0(new_n5598_), .A1(new_n5590_), .B0(new_n5599_), .Y(new_n5600_));
  OAI21X1  g04598(.A0(new_n5600_), .A1(new_n5589_), .B0(new_n5552_), .Y(new_n5601_));
  MX2X1    g04599(.A(new_n5551_), .B(new_n5542_), .S0(new_n5529_), .Y(new_n5602_));
  NOR3X1   g04600(.A(new_n5599_), .B(new_n5586_), .C(new_n5575_), .Y(new_n5603_));
  AOI21X1  g04601(.A0(new_n5598_), .A1(new_n5590_), .B0(new_n5588_), .Y(new_n5604_));
  OAI21X1  g04602(.A0(new_n5604_), .A1(new_n5603_), .B0(new_n5602_), .Y(new_n5605_));
  XOR2X1   g04603(.A(new_n5079_), .B(new_n5040_), .Y(new_n5606_));
  NOR2X1   g04604(.A(new_n5606_), .B(new_n5003_), .Y(new_n5607_));
  NAND3X1  g04605(.A(new_n5607_), .B(new_n5605_), .C(new_n5601_), .Y(new_n5608_));
  NAND3X1  g04606(.A(new_n5599_), .B(new_n5598_), .C(new_n5590_), .Y(new_n5609_));
  OAI21X1  g04607(.A0(new_n5586_), .A1(new_n5575_), .B0(new_n5588_), .Y(new_n5610_));
  AOI21X1  g04608(.A0(new_n5610_), .A1(new_n5609_), .B0(new_n5602_), .Y(new_n5611_));
  NAND3X1  g04609(.A(new_n5588_), .B(new_n5598_), .C(new_n5590_), .Y(new_n5612_));
  OAI21X1  g04610(.A0(new_n5586_), .A1(new_n5575_), .B0(new_n5599_), .Y(new_n5613_));
  AOI21X1  g04611(.A0(new_n5613_), .A1(new_n5612_), .B0(new_n5552_), .Y(new_n5614_));
  INVX1    g04612(.A(new_n5607_), .Y(new_n5615_));
  OAI21X1  g04613(.A0(new_n5614_), .A1(new_n5611_), .B0(new_n5615_), .Y(new_n5616_));
  AOI21X1  g04614(.A0(new_n5616_), .A1(new_n5608_), .B0(new_n5520_), .Y(new_n5617_));
  NOR2X1   g04615(.A(new_n5519_), .B(new_n5513_), .Y(new_n5618_));
  NAND3X1  g04616(.A(new_n5615_), .B(new_n5605_), .C(new_n5601_), .Y(new_n5619_));
  OAI21X1  g04617(.A0(new_n5614_), .A1(new_n5611_), .B0(new_n5607_), .Y(new_n5620_));
  AOI21X1  g04618(.A0(new_n5620_), .A1(new_n5619_), .B0(new_n5618_), .Y(new_n5621_));
  OR4X1    g04619(.A(new_n5621_), .B(new_n5617_), .C(new_n5235_), .D(new_n5081_), .Y(new_n5622_));
  OAI22X1  g04620(.A0(new_n5621_), .A1(new_n5617_), .B0(new_n5235_), .B1(new_n5081_), .Y(new_n5623_));
  AOI21X1  g04621(.A0(new_n5623_), .A1(new_n5622_), .B0(new_n5435_), .Y(new_n5624_));
  NOR2X1   g04622(.A(new_n5235_), .B(new_n5081_), .Y(new_n5625_));
  OR2X1    g04623(.A(new_n5625_), .B(new_n5621_), .Y(new_n5626_));
  OAI21X1  g04624(.A0(new_n5621_), .A1(new_n5617_), .B0(new_n5625_), .Y(new_n5627_));
  OAI21X1  g04625(.A0(new_n5626_), .A1(new_n5617_), .B0(new_n5627_), .Y(new_n5628_));
  AOI21X1  g04626(.A0(new_n5628_), .A1(new_n5435_), .B0(new_n5624_), .Y(new_n5629_));
  OAI21X1  g04627(.A0(new_n5249_), .A1(new_n5238_), .B0(new_n5629_), .Y(new_n5630_));
  NAND2X1  g04628(.A(new_n5623_), .B(new_n5622_), .Y(new_n5631_));
  NOR2X1   g04629(.A(new_n5430_), .B(new_n5424_), .Y(new_n5632_));
  NAND3X1  g04630(.A(new_n5344_), .B(new_n5334_), .C(new_n5330_), .Y(new_n5633_));
  OAI21X1  g04631(.A0(new_n5343_), .A1(new_n5340_), .B0(new_n5336_), .Y(new_n5634_));
  AND2X1   g04632(.A(new_n5634_), .B(new_n5633_), .Y(new_n5635_));
  MX2X1    g04633(.A(new_n5635_), .B(new_n5346_), .S0(new_n5632_), .Y(new_n5636_));
  MX2X1    g04634(.A(new_n5628_), .B(new_n5631_), .S0(new_n5636_), .Y(new_n5637_));
  AOI21X1  g04635(.A0(new_n4922_), .A1(new_n4186_), .B0(new_n5248_), .Y(new_n5638_));
  AND2X1   g04636(.A(new_n5638_), .B(new_n5243_), .Y(new_n5639_));
  AOI21X1  g04637(.A0(new_n5247_), .A1(new_n5243_), .B0(new_n5237_), .Y(new_n5640_));
  OAI21X1  g04638(.A0(new_n5640_), .A1(new_n5639_), .B0(new_n5637_), .Y(new_n5641_));
  NAND2X1  g04639(.A(new_n5641_), .B(new_n5630_), .Y(new_n5642_));
  INVX1    g04640(.A(\A[201] ), .Y(new_n5643_));
  INVX1    g04641(.A(\A[200] ), .Y(new_n5644_));
  OR2X1    g04642(.A(new_n5644_), .B(\A[199] ), .Y(new_n5645_));
  AOI21X1  g04643(.A0(new_n5644_), .A1(\A[199] ), .B0(new_n5643_), .Y(new_n5646_));
  XOR2X1   g04644(.A(\A[200] ), .B(\A[199] ), .Y(new_n5647_));
  AOI22X1  g04645(.A0(new_n5647_), .A1(new_n5643_), .B0(new_n5646_), .B1(new_n5645_), .Y(new_n5648_));
  INVX1    g04646(.A(\A[204] ), .Y(new_n5649_));
  INVX1    g04647(.A(\A[203] ), .Y(new_n5650_));
  OR2X1    g04648(.A(new_n5650_), .B(\A[202] ), .Y(new_n5651_));
  AOI21X1  g04649(.A0(new_n5650_), .A1(\A[202] ), .B0(new_n5649_), .Y(new_n5652_));
  XOR2X1   g04650(.A(\A[203] ), .B(\A[202] ), .Y(new_n5653_));
  AOI22X1  g04651(.A0(new_n5653_), .A1(new_n5649_), .B0(new_n5652_), .B1(new_n5651_), .Y(new_n5654_));
  OR2X1    g04652(.A(new_n5654_), .B(new_n5648_), .Y(new_n5655_));
  AND2X1   g04653(.A(\A[203] ), .B(\A[202] ), .Y(new_n5656_));
  AND2X1   g04654(.A(new_n5653_), .B(\A[204] ), .Y(new_n5657_));
  OR2X1    g04655(.A(new_n5657_), .B(new_n5656_), .Y(new_n5658_));
  AND2X1   g04656(.A(\A[200] ), .B(\A[199] ), .Y(new_n5659_));
  AOI21X1  g04657(.A0(new_n5647_), .A1(\A[201] ), .B0(new_n5659_), .Y(new_n5660_));
  XOR2X1   g04658(.A(new_n5660_), .B(new_n5658_), .Y(new_n5661_));
  XOR2X1   g04659(.A(new_n5661_), .B(new_n5655_), .Y(new_n5662_));
  INVX1    g04660(.A(\A[199] ), .Y(new_n5663_));
  AND2X1   g04661(.A(\A[200] ), .B(new_n5663_), .Y(new_n5664_));
  OAI21X1  g04662(.A0(\A[200] ), .A1(new_n5663_), .B0(\A[201] ), .Y(new_n5665_));
  NAND2X1  g04663(.A(new_n5647_), .B(new_n5643_), .Y(new_n5666_));
  OAI21X1  g04664(.A0(new_n5665_), .A1(new_n5664_), .B0(new_n5666_), .Y(new_n5667_));
  XOR2X1   g04665(.A(new_n5654_), .B(new_n5667_), .Y(new_n5668_));
  NOR2X1   g04666(.A(new_n5654_), .B(new_n5648_), .Y(new_n5669_));
  AOI21X1  g04667(.A0(new_n5653_), .A1(\A[204] ), .B0(new_n5656_), .Y(new_n5670_));
  XOR2X1   g04668(.A(new_n5660_), .B(new_n5670_), .Y(new_n5671_));
  NOR2X1   g04669(.A(new_n5660_), .B(new_n5670_), .Y(new_n5672_));
  AOI21X1  g04670(.A0(new_n5671_), .A1(new_n5669_), .B0(new_n5672_), .Y(new_n5673_));
  OAI21X1  g04671(.A0(new_n5673_), .A1(new_n5668_), .B0(new_n5662_), .Y(new_n5674_));
  AND2X1   g04672(.A(\A[209] ), .B(\A[208] ), .Y(new_n5675_));
  XOR2X1   g04673(.A(\A[209] ), .B(\A[208] ), .Y(new_n5676_));
  AOI21X1  g04674(.A0(new_n5676_), .A1(\A[210] ), .B0(new_n5675_), .Y(new_n5677_));
  AND2X1   g04675(.A(\A[206] ), .B(\A[205] ), .Y(new_n5678_));
  XOR2X1   g04676(.A(\A[206] ), .B(\A[205] ), .Y(new_n5679_));
  AOI21X1  g04677(.A0(new_n5679_), .A1(\A[207] ), .B0(new_n5678_), .Y(new_n5680_));
  INVX1    g04678(.A(\A[207] ), .Y(new_n5681_));
  INVX1    g04679(.A(\A[206] ), .Y(new_n5682_));
  OR2X1    g04680(.A(new_n5682_), .B(\A[205] ), .Y(new_n5683_));
  AOI21X1  g04681(.A0(new_n5682_), .A1(\A[205] ), .B0(new_n5681_), .Y(new_n5684_));
  AOI22X1  g04682(.A0(new_n5684_), .A1(new_n5683_), .B0(new_n5679_), .B1(new_n5681_), .Y(new_n5685_));
  INVX1    g04683(.A(\A[210] ), .Y(new_n5686_));
  INVX1    g04684(.A(\A[209] ), .Y(new_n5687_));
  OR2X1    g04685(.A(new_n5687_), .B(\A[208] ), .Y(new_n5688_));
  AOI21X1  g04686(.A0(new_n5687_), .A1(\A[208] ), .B0(new_n5686_), .Y(new_n5689_));
  AOI22X1  g04687(.A0(new_n5689_), .A1(new_n5688_), .B0(new_n5676_), .B1(new_n5686_), .Y(new_n5690_));
  NOR4X1   g04688(.A(new_n5690_), .B(new_n5685_), .C(new_n5680_), .D(new_n5677_), .Y(new_n5691_));
  NOR4X1   g04689(.A(new_n5660_), .B(new_n5670_), .C(new_n5654_), .D(new_n5648_), .Y(new_n5692_));
  INVX1    g04690(.A(\A[205] ), .Y(new_n5693_));
  AND2X1   g04691(.A(\A[206] ), .B(new_n5693_), .Y(new_n5694_));
  OAI21X1  g04692(.A0(\A[206] ), .A1(new_n5693_), .B0(\A[207] ), .Y(new_n5695_));
  NAND2X1  g04693(.A(new_n5679_), .B(new_n5681_), .Y(new_n5696_));
  OAI21X1  g04694(.A0(new_n5695_), .A1(new_n5694_), .B0(new_n5696_), .Y(new_n5697_));
  XOR2X1   g04695(.A(new_n5690_), .B(new_n5697_), .Y(new_n5698_));
  OR4X1    g04696(.A(new_n5698_), .B(new_n5692_), .C(new_n5691_), .D(new_n5668_), .Y(new_n5699_));
  AND2X1   g04697(.A(new_n5676_), .B(\A[210] ), .Y(new_n5700_));
  OR2X1    g04698(.A(new_n5700_), .B(new_n5675_), .Y(new_n5701_));
  XOR2X1   g04699(.A(new_n5680_), .B(new_n5701_), .Y(new_n5702_));
  OR2X1    g04700(.A(new_n5690_), .B(new_n5685_), .Y(new_n5703_));
  OR2X1    g04701(.A(new_n5680_), .B(new_n5677_), .Y(new_n5704_));
  OAI21X1  g04702(.A0(new_n5703_), .A1(new_n5702_), .B0(new_n5704_), .Y(new_n5705_));
  NOR2X1   g04703(.A(new_n5690_), .B(new_n5685_), .Y(new_n5706_));
  XOR2X1   g04704(.A(new_n5706_), .B(new_n5702_), .Y(new_n5707_));
  XOR2X1   g04705(.A(new_n5690_), .B(new_n5685_), .Y(new_n5708_));
  AOI21X1  g04706(.A0(new_n5708_), .A1(new_n5705_), .B0(new_n5707_), .Y(new_n5709_));
  XOR2X1   g04707(.A(new_n5709_), .B(new_n5699_), .Y(new_n5710_));
  XOR2X1   g04708(.A(new_n5680_), .B(new_n5677_), .Y(new_n5711_));
  NOR2X1   g04709(.A(new_n5680_), .B(new_n5677_), .Y(new_n5712_));
  AOI21X1  g04710(.A0(new_n5706_), .A1(new_n5711_), .B0(new_n5712_), .Y(new_n5713_));
  XOR2X1   g04711(.A(new_n5706_), .B(new_n5711_), .Y(new_n5714_));
  OAI21X1  g04712(.A0(new_n5698_), .A1(new_n5713_), .B0(new_n5714_), .Y(new_n5715_));
  NOR4X1   g04713(.A(new_n5698_), .B(new_n5692_), .C(new_n5707_), .D(new_n5668_), .Y(new_n5716_));
  OAI21X1  g04714(.A0(new_n5708_), .A1(new_n5714_), .B0(new_n5705_), .Y(new_n5717_));
  AOI22X1  g04715(.A0(new_n5717_), .A1(new_n5716_), .B0(new_n5715_), .B1(new_n5699_), .Y(new_n5718_));
  MX2X1    g04716(.A(new_n5718_), .B(new_n5710_), .S0(new_n5674_), .Y(new_n5719_));
  INVX1    g04717(.A(\A[213] ), .Y(new_n5720_));
  INVX1    g04718(.A(\A[212] ), .Y(new_n5721_));
  OR2X1    g04719(.A(new_n5721_), .B(\A[211] ), .Y(new_n5722_));
  AOI21X1  g04720(.A0(new_n5721_), .A1(\A[211] ), .B0(new_n5720_), .Y(new_n5723_));
  XOR2X1   g04721(.A(\A[212] ), .B(\A[211] ), .Y(new_n5724_));
  AOI22X1  g04722(.A0(new_n5724_), .A1(new_n5720_), .B0(new_n5723_), .B1(new_n5722_), .Y(new_n5725_));
  INVX1    g04723(.A(\A[216] ), .Y(new_n5726_));
  INVX1    g04724(.A(\A[215] ), .Y(new_n5727_));
  OR2X1    g04725(.A(new_n5727_), .B(\A[214] ), .Y(new_n5728_));
  AOI21X1  g04726(.A0(new_n5727_), .A1(\A[214] ), .B0(new_n5726_), .Y(new_n5729_));
  XOR2X1   g04727(.A(\A[215] ), .B(\A[214] ), .Y(new_n5730_));
  AOI22X1  g04728(.A0(new_n5730_), .A1(new_n5726_), .B0(new_n5729_), .B1(new_n5728_), .Y(new_n5731_));
  OR2X1    g04729(.A(new_n5731_), .B(new_n5725_), .Y(new_n5732_));
  AND2X1   g04730(.A(\A[215] ), .B(\A[214] ), .Y(new_n5733_));
  AND2X1   g04731(.A(new_n5730_), .B(\A[216] ), .Y(new_n5734_));
  OR2X1    g04732(.A(new_n5734_), .B(new_n5733_), .Y(new_n5735_));
  AND2X1   g04733(.A(\A[212] ), .B(\A[211] ), .Y(new_n5736_));
  AOI21X1  g04734(.A0(new_n5724_), .A1(\A[213] ), .B0(new_n5736_), .Y(new_n5737_));
  XOR2X1   g04735(.A(new_n5737_), .B(new_n5735_), .Y(new_n5738_));
  XOR2X1   g04736(.A(new_n5738_), .B(new_n5732_), .Y(new_n5739_));
  INVX1    g04737(.A(\A[211] ), .Y(new_n5740_));
  AND2X1   g04738(.A(\A[212] ), .B(new_n5740_), .Y(new_n5741_));
  OAI21X1  g04739(.A0(\A[212] ), .A1(new_n5740_), .B0(\A[213] ), .Y(new_n5742_));
  NAND2X1  g04740(.A(new_n5724_), .B(new_n5720_), .Y(new_n5743_));
  OAI21X1  g04741(.A0(new_n5742_), .A1(new_n5741_), .B0(new_n5743_), .Y(new_n5744_));
  XOR2X1   g04742(.A(new_n5731_), .B(new_n5744_), .Y(new_n5745_));
  NOR2X1   g04743(.A(new_n5731_), .B(new_n5725_), .Y(new_n5746_));
  AOI21X1  g04744(.A0(new_n5730_), .A1(\A[216] ), .B0(new_n5733_), .Y(new_n5747_));
  XOR2X1   g04745(.A(new_n5737_), .B(new_n5747_), .Y(new_n5748_));
  NOR2X1   g04746(.A(new_n5737_), .B(new_n5747_), .Y(new_n5749_));
  AOI21X1  g04747(.A0(new_n5748_), .A1(new_n5746_), .B0(new_n5749_), .Y(new_n5750_));
  OAI21X1  g04748(.A0(new_n5750_), .A1(new_n5745_), .B0(new_n5739_), .Y(new_n5751_));
  AND2X1   g04749(.A(\A[221] ), .B(\A[220] ), .Y(new_n5752_));
  XOR2X1   g04750(.A(\A[221] ), .B(\A[220] ), .Y(new_n5753_));
  AOI21X1  g04751(.A0(new_n5753_), .A1(\A[222] ), .B0(new_n5752_), .Y(new_n5754_));
  AND2X1   g04752(.A(\A[218] ), .B(\A[217] ), .Y(new_n5755_));
  XOR2X1   g04753(.A(\A[218] ), .B(\A[217] ), .Y(new_n5756_));
  AOI21X1  g04754(.A0(new_n5756_), .A1(\A[219] ), .B0(new_n5755_), .Y(new_n5757_));
  INVX1    g04755(.A(\A[219] ), .Y(new_n5758_));
  INVX1    g04756(.A(\A[218] ), .Y(new_n5759_));
  OR2X1    g04757(.A(new_n5759_), .B(\A[217] ), .Y(new_n5760_));
  AOI21X1  g04758(.A0(new_n5759_), .A1(\A[217] ), .B0(new_n5758_), .Y(new_n5761_));
  AOI22X1  g04759(.A0(new_n5761_), .A1(new_n5760_), .B0(new_n5756_), .B1(new_n5758_), .Y(new_n5762_));
  INVX1    g04760(.A(\A[222] ), .Y(new_n5763_));
  INVX1    g04761(.A(\A[221] ), .Y(new_n5764_));
  OR2X1    g04762(.A(new_n5764_), .B(\A[220] ), .Y(new_n5765_));
  AOI21X1  g04763(.A0(new_n5764_), .A1(\A[220] ), .B0(new_n5763_), .Y(new_n5766_));
  AOI22X1  g04764(.A0(new_n5766_), .A1(new_n5765_), .B0(new_n5753_), .B1(new_n5763_), .Y(new_n5767_));
  NOR4X1   g04765(.A(new_n5767_), .B(new_n5762_), .C(new_n5757_), .D(new_n5754_), .Y(new_n5768_));
  NOR4X1   g04766(.A(new_n5737_), .B(new_n5747_), .C(new_n5731_), .D(new_n5725_), .Y(new_n5769_));
  INVX1    g04767(.A(\A[217] ), .Y(new_n5770_));
  AND2X1   g04768(.A(\A[218] ), .B(new_n5770_), .Y(new_n5771_));
  OAI21X1  g04769(.A0(\A[218] ), .A1(new_n5770_), .B0(\A[219] ), .Y(new_n5772_));
  NAND2X1  g04770(.A(new_n5756_), .B(new_n5758_), .Y(new_n5773_));
  OAI21X1  g04771(.A0(new_n5772_), .A1(new_n5771_), .B0(new_n5773_), .Y(new_n5774_));
  XOR2X1   g04772(.A(new_n5767_), .B(new_n5774_), .Y(new_n5775_));
  OR4X1    g04773(.A(new_n5775_), .B(new_n5769_), .C(new_n5768_), .D(new_n5745_), .Y(new_n5776_));
  XOR2X1   g04774(.A(new_n5757_), .B(new_n5754_), .Y(new_n5777_));
  NOR2X1   g04775(.A(new_n5767_), .B(new_n5762_), .Y(new_n5778_));
  NOR2X1   g04776(.A(new_n5757_), .B(new_n5754_), .Y(new_n5779_));
  AOI21X1  g04777(.A0(new_n5778_), .A1(new_n5777_), .B0(new_n5779_), .Y(new_n5780_));
  XOR2X1   g04778(.A(new_n5778_), .B(new_n5777_), .Y(new_n5781_));
  OAI21X1  g04779(.A0(new_n5775_), .A1(new_n5780_), .B0(new_n5781_), .Y(new_n5782_));
  XOR2X1   g04780(.A(new_n5782_), .B(new_n5776_), .Y(new_n5783_));
  AND2X1   g04781(.A(new_n5783_), .B(new_n5751_), .Y(new_n5784_));
  OR2X1    g04782(.A(new_n5775_), .B(new_n5768_), .Y(new_n5785_));
  XOR2X1   g04783(.A(new_n5731_), .B(new_n5725_), .Y(new_n5786_));
  XOR2X1   g04784(.A(new_n5786_), .B(new_n5785_), .Y(new_n5787_));
  OR2X1    g04785(.A(new_n5698_), .B(new_n5691_), .Y(new_n5788_));
  XOR2X1   g04786(.A(new_n5654_), .B(new_n5648_), .Y(new_n5789_));
  XOR2X1   g04787(.A(new_n5789_), .B(new_n5788_), .Y(new_n5790_));
  NOR2X1   g04788(.A(new_n5790_), .B(new_n5787_), .Y(new_n5791_));
  AND2X1   g04789(.A(new_n5753_), .B(\A[222] ), .Y(new_n5792_));
  OR2X1    g04790(.A(new_n5792_), .B(new_n5752_), .Y(new_n5793_));
  XOR2X1   g04791(.A(new_n5757_), .B(new_n5793_), .Y(new_n5794_));
  XOR2X1   g04792(.A(new_n5778_), .B(new_n5794_), .Y(new_n5795_));
  NOR4X1   g04793(.A(new_n5775_), .B(new_n5769_), .C(new_n5795_), .D(new_n5745_), .Y(new_n5796_));
  OR2X1    g04794(.A(new_n5767_), .B(new_n5762_), .Y(new_n5797_));
  OR2X1    g04795(.A(new_n5757_), .B(new_n5754_), .Y(new_n5798_));
  OAI21X1  g04796(.A0(new_n5797_), .A1(new_n5794_), .B0(new_n5798_), .Y(new_n5799_));
  XOR2X1   g04797(.A(new_n5767_), .B(new_n5762_), .Y(new_n5800_));
  OAI21X1  g04798(.A0(new_n5800_), .A1(new_n5781_), .B0(new_n5799_), .Y(new_n5801_));
  AOI22X1  g04799(.A0(new_n5801_), .A1(new_n5796_), .B0(new_n5782_), .B1(new_n5776_), .Y(new_n5802_));
  OAI21X1  g04800(.A0(new_n5802_), .A1(new_n5751_), .B0(new_n5791_), .Y(new_n5803_));
  AOI21X1  g04801(.A0(new_n5800_), .A1(new_n5799_), .B0(new_n5795_), .Y(new_n5804_));
  XOR2X1   g04802(.A(new_n5804_), .B(new_n5776_), .Y(new_n5805_));
  MX2X1    g04803(.A(new_n5802_), .B(new_n5805_), .S0(new_n5751_), .Y(new_n5806_));
  OAI22X1  g04804(.A0(new_n5806_), .A1(new_n5791_), .B0(new_n5803_), .B1(new_n5784_), .Y(new_n5807_));
  AND2X1   g04805(.A(new_n5807_), .B(new_n5719_), .Y(new_n5808_));
  XOR2X1   g04806(.A(new_n5731_), .B(new_n5744_), .Y(new_n5809_));
  XOR2X1   g04807(.A(new_n5809_), .B(new_n5785_), .Y(new_n5810_));
  XOR2X1   g04808(.A(new_n5790_), .B(new_n5810_), .Y(new_n5811_));
  INVX1    g04809(.A(\A[194] ), .Y(new_n5812_));
  AND2X1   g04810(.A(new_n5812_), .B(\A[193] ), .Y(new_n5813_));
  OAI21X1  g04811(.A0(new_n5812_), .A1(\A[193] ), .B0(\A[195] ), .Y(new_n5814_));
  INVX1    g04812(.A(\A[195] ), .Y(new_n5815_));
  XOR2X1   g04813(.A(\A[194] ), .B(\A[193] ), .Y(new_n5816_));
  NAND2X1  g04814(.A(new_n5816_), .B(new_n5815_), .Y(new_n5817_));
  OAI21X1  g04815(.A0(new_n5814_), .A1(new_n5813_), .B0(new_n5817_), .Y(new_n5818_));
  INVX1    g04816(.A(\A[198] ), .Y(new_n5819_));
  INVX1    g04817(.A(\A[196] ), .Y(new_n5820_));
  OR2X1    g04818(.A(\A[197] ), .B(new_n5820_), .Y(new_n5821_));
  AOI21X1  g04819(.A0(\A[197] ), .A1(new_n5820_), .B0(new_n5819_), .Y(new_n5822_));
  XOR2X1   g04820(.A(\A[197] ), .B(\A[196] ), .Y(new_n5823_));
  AOI22X1  g04821(.A0(new_n5823_), .A1(new_n5819_), .B0(new_n5822_), .B1(new_n5821_), .Y(new_n5824_));
  AND2X1   g04822(.A(\A[197] ), .B(\A[196] ), .Y(new_n5825_));
  AOI21X1  g04823(.A0(new_n5823_), .A1(\A[198] ), .B0(new_n5825_), .Y(new_n5826_));
  AND2X1   g04824(.A(\A[194] ), .B(\A[193] ), .Y(new_n5827_));
  AOI21X1  g04825(.A0(new_n5816_), .A1(\A[195] ), .B0(new_n5827_), .Y(new_n5828_));
  XOR2X1   g04826(.A(new_n5824_), .B(new_n5818_), .Y(new_n5829_));
  INVX1    g04827(.A(\A[189] ), .Y(new_n5830_));
  INVX1    g04828(.A(\A[187] ), .Y(new_n5831_));
  OR2X1    g04829(.A(\A[188] ), .B(new_n5831_), .Y(new_n5832_));
  AOI21X1  g04830(.A0(\A[188] ), .A1(new_n5831_), .B0(new_n5830_), .Y(new_n5833_));
  XOR2X1   g04831(.A(\A[188] ), .B(\A[187] ), .Y(new_n5834_));
  AOI22X1  g04832(.A0(new_n5834_), .A1(new_n5830_), .B0(new_n5833_), .B1(new_n5832_), .Y(new_n5835_));
  INVX1    g04833(.A(\A[192] ), .Y(new_n5836_));
  INVX1    g04834(.A(\A[190] ), .Y(new_n5837_));
  OR2X1    g04835(.A(\A[191] ), .B(new_n5837_), .Y(new_n5838_));
  AOI21X1  g04836(.A0(\A[191] ), .A1(new_n5837_), .B0(new_n5836_), .Y(new_n5839_));
  XOR2X1   g04837(.A(\A[191] ), .B(\A[190] ), .Y(new_n5840_));
  AOI22X1  g04838(.A0(new_n5840_), .A1(new_n5836_), .B0(new_n5839_), .B1(new_n5838_), .Y(new_n5841_));
  AND2X1   g04839(.A(\A[191] ), .B(\A[190] ), .Y(new_n5842_));
  AOI21X1  g04840(.A0(new_n5840_), .A1(\A[192] ), .B0(new_n5842_), .Y(new_n5843_));
  AND2X1   g04841(.A(\A[188] ), .B(\A[187] ), .Y(new_n5844_));
  AOI21X1  g04842(.A0(new_n5834_), .A1(\A[189] ), .B0(new_n5844_), .Y(new_n5845_));
  XOR2X1   g04843(.A(new_n5841_), .B(new_n5835_), .Y(new_n5846_));
  XOR2X1   g04844(.A(new_n5846_), .B(new_n5829_), .Y(new_n5847_));
  INVX1    g04845(.A(new_n5847_), .Y(new_n5848_));
  INVX1    g04846(.A(\A[182] ), .Y(new_n5849_));
  AND2X1   g04847(.A(new_n5849_), .B(\A[181] ), .Y(new_n5850_));
  OAI21X1  g04848(.A0(new_n5849_), .A1(\A[181] ), .B0(\A[183] ), .Y(new_n5851_));
  INVX1    g04849(.A(\A[183] ), .Y(new_n5852_));
  XOR2X1   g04850(.A(\A[182] ), .B(\A[181] ), .Y(new_n5853_));
  NAND2X1  g04851(.A(new_n5853_), .B(new_n5852_), .Y(new_n5854_));
  OAI21X1  g04852(.A0(new_n5851_), .A1(new_n5850_), .B0(new_n5854_), .Y(new_n5855_));
  INVX1    g04853(.A(\A[186] ), .Y(new_n5856_));
  INVX1    g04854(.A(\A[184] ), .Y(new_n5857_));
  OR2X1    g04855(.A(\A[185] ), .B(new_n5857_), .Y(new_n5858_));
  AOI21X1  g04856(.A0(\A[185] ), .A1(new_n5857_), .B0(new_n5856_), .Y(new_n5859_));
  XOR2X1   g04857(.A(\A[185] ), .B(\A[184] ), .Y(new_n5860_));
  AOI22X1  g04858(.A0(new_n5860_), .A1(new_n5856_), .B0(new_n5859_), .B1(new_n5858_), .Y(new_n5861_));
  AND2X1   g04859(.A(\A[185] ), .B(\A[184] ), .Y(new_n5862_));
  AOI21X1  g04860(.A0(new_n5860_), .A1(\A[186] ), .B0(new_n5862_), .Y(new_n5863_));
  AND2X1   g04861(.A(\A[182] ), .B(\A[181] ), .Y(new_n5864_));
  AOI21X1  g04862(.A0(new_n5853_), .A1(\A[183] ), .B0(new_n5864_), .Y(new_n5865_));
  XOR2X1   g04863(.A(new_n5861_), .B(new_n5855_), .Y(new_n5866_));
  INVX1    g04864(.A(\A[177] ), .Y(new_n5867_));
  INVX1    g04865(.A(\A[175] ), .Y(new_n5868_));
  OR2X1    g04866(.A(\A[176] ), .B(new_n5868_), .Y(new_n5869_));
  AOI21X1  g04867(.A0(\A[176] ), .A1(new_n5868_), .B0(new_n5867_), .Y(new_n5870_));
  XOR2X1   g04868(.A(\A[176] ), .B(\A[175] ), .Y(new_n5871_));
  AOI22X1  g04869(.A0(new_n5871_), .A1(new_n5867_), .B0(new_n5870_), .B1(new_n5869_), .Y(new_n5872_));
  INVX1    g04870(.A(\A[180] ), .Y(new_n5873_));
  INVX1    g04871(.A(\A[178] ), .Y(new_n5874_));
  OR2X1    g04872(.A(\A[179] ), .B(new_n5874_), .Y(new_n5875_));
  AOI21X1  g04873(.A0(\A[179] ), .A1(new_n5874_), .B0(new_n5873_), .Y(new_n5876_));
  XOR2X1   g04874(.A(\A[179] ), .B(\A[178] ), .Y(new_n5877_));
  AOI22X1  g04875(.A0(new_n5877_), .A1(new_n5873_), .B0(new_n5876_), .B1(new_n5875_), .Y(new_n5878_));
  AND2X1   g04876(.A(\A[179] ), .B(\A[178] ), .Y(new_n5879_));
  AOI21X1  g04877(.A0(new_n5877_), .A1(\A[180] ), .B0(new_n5879_), .Y(new_n5880_));
  AND2X1   g04878(.A(\A[176] ), .B(\A[175] ), .Y(new_n5881_));
  AOI21X1  g04879(.A0(new_n5871_), .A1(\A[177] ), .B0(new_n5881_), .Y(new_n5882_));
  XOR2X1   g04880(.A(new_n5878_), .B(new_n5872_), .Y(new_n5883_));
  XOR2X1   g04881(.A(new_n5883_), .B(new_n5866_), .Y(new_n5884_));
  XOR2X1   g04882(.A(new_n5884_), .B(new_n5848_), .Y(new_n5885_));
  NOR2X1   g04883(.A(new_n5885_), .B(new_n5811_), .Y(new_n5886_));
  NAND2X1  g04884(.A(new_n5783_), .B(new_n5751_), .Y(new_n5887_));
  NOR4X1   g04885(.A(new_n5775_), .B(new_n5769_), .C(new_n5768_), .D(new_n5745_), .Y(new_n5888_));
  OR4X1    g04886(.A(new_n5775_), .B(new_n5769_), .C(new_n5795_), .D(new_n5745_), .Y(new_n5889_));
  AOI21X1  g04887(.A0(new_n5775_), .A1(new_n5795_), .B0(new_n5780_), .Y(new_n5890_));
  OAI22X1  g04888(.A0(new_n5890_), .A1(new_n5889_), .B0(new_n5804_), .B1(new_n5888_), .Y(new_n5891_));
  MX2X1    g04889(.A(new_n5891_), .B(new_n5783_), .S0(new_n5751_), .Y(new_n5892_));
  XOR2X1   g04890(.A(new_n5738_), .B(new_n5746_), .Y(new_n5893_));
  XOR2X1   g04891(.A(new_n5731_), .B(new_n5725_), .Y(new_n5894_));
  OR2X1    g04892(.A(new_n5737_), .B(new_n5747_), .Y(new_n5895_));
  OAI21X1  g04893(.A0(new_n5738_), .A1(new_n5732_), .B0(new_n5895_), .Y(new_n5896_));
  AOI21X1  g04894(.A0(new_n5896_), .A1(new_n5894_), .B0(new_n5893_), .Y(new_n5897_));
  AOI21X1  g04895(.A0(new_n5891_), .A1(new_n5897_), .B0(new_n5791_), .Y(new_n5898_));
  AOI22X1  g04896(.A0(new_n5898_), .A1(new_n5887_), .B0(new_n5892_), .B1(new_n5791_), .Y(new_n5899_));
  OAI21X1  g04897(.A0(new_n5899_), .A1(new_n5719_), .B0(new_n5886_), .Y(new_n5900_));
  NOR4X1   g04898(.A(new_n5698_), .B(new_n5692_), .C(new_n5691_), .D(new_n5668_), .Y(new_n5901_));
  XOR2X1   g04899(.A(new_n5709_), .B(new_n5901_), .Y(new_n5902_));
  OR4X1    g04900(.A(new_n5698_), .B(new_n5692_), .C(new_n5707_), .D(new_n5668_), .Y(new_n5903_));
  AOI21X1  g04901(.A0(new_n5698_), .A1(new_n5707_), .B0(new_n5713_), .Y(new_n5904_));
  OAI22X1  g04902(.A0(new_n5904_), .A1(new_n5903_), .B0(new_n5709_), .B1(new_n5901_), .Y(new_n5905_));
  MX2X1    g04903(.A(new_n5905_), .B(new_n5902_), .S0(new_n5674_), .Y(new_n5906_));
  OR2X1    g04904(.A(new_n5790_), .B(new_n5787_), .Y(new_n5907_));
  AOI21X1  g04905(.A0(new_n5891_), .A1(new_n5897_), .B0(new_n5907_), .Y(new_n5908_));
  AOI22X1  g04906(.A0(new_n5892_), .A1(new_n5907_), .B0(new_n5908_), .B1(new_n5887_), .Y(new_n5909_));
  MX2X1    g04907(.A(new_n5909_), .B(new_n5899_), .S0(new_n5906_), .Y(new_n5910_));
  OAI22X1  g04908(.A0(new_n5910_), .A1(new_n5886_), .B0(new_n5900_), .B1(new_n5808_), .Y(new_n5911_));
  INVX1    g04909(.A(\A[188] ), .Y(new_n5912_));
  AND2X1   g04910(.A(new_n5912_), .B(\A[187] ), .Y(new_n5913_));
  OAI21X1  g04911(.A0(new_n5912_), .A1(\A[187] ), .B0(\A[189] ), .Y(new_n5914_));
  NAND2X1  g04912(.A(new_n5834_), .B(new_n5830_), .Y(new_n5915_));
  OAI21X1  g04913(.A0(new_n5914_), .A1(new_n5913_), .B0(new_n5915_), .Y(new_n5916_));
  XOR2X1   g04914(.A(new_n5841_), .B(new_n5916_), .Y(new_n5917_));
  XOR2X1   g04915(.A(new_n5845_), .B(new_n5843_), .Y(new_n5918_));
  NOR2X1   g04916(.A(new_n5841_), .B(new_n5835_), .Y(new_n5919_));
  NOR2X1   g04917(.A(new_n5845_), .B(new_n5843_), .Y(new_n5920_));
  AOI21X1  g04918(.A0(new_n5919_), .A1(new_n5918_), .B0(new_n5920_), .Y(new_n5921_));
  XOR2X1   g04919(.A(new_n5919_), .B(new_n5918_), .Y(new_n5922_));
  OAI21X1  g04920(.A0(new_n5921_), .A1(new_n5917_), .B0(new_n5922_), .Y(new_n5923_));
  XOR2X1   g04921(.A(new_n5824_), .B(new_n5818_), .Y(new_n5924_));
  INVX1    g04922(.A(\A[193] ), .Y(new_n5925_));
  OR2X1    g04923(.A(\A[194] ), .B(new_n5925_), .Y(new_n5926_));
  AOI21X1  g04924(.A0(\A[194] ), .A1(new_n5925_), .B0(new_n5815_), .Y(new_n5927_));
  AOI22X1  g04925(.A0(new_n5816_), .A1(new_n5815_), .B0(new_n5927_), .B1(new_n5926_), .Y(new_n5928_));
  NOR4X1   g04926(.A(new_n5828_), .B(new_n5826_), .C(new_n5824_), .D(new_n5928_), .Y(new_n5929_));
  NOR4X1   g04927(.A(new_n5845_), .B(new_n5843_), .C(new_n5841_), .D(new_n5835_), .Y(new_n5930_));
  OR4X1    g04928(.A(new_n5930_), .B(new_n5917_), .C(new_n5929_), .D(new_n5924_), .Y(new_n5931_));
  XOR2X1   g04929(.A(new_n5828_), .B(new_n5826_), .Y(new_n5932_));
  NOR2X1   g04930(.A(new_n5824_), .B(new_n5928_), .Y(new_n5933_));
  NOR2X1   g04931(.A(new_n5828_), .B(new_n5826_), .Y(new_n5934_));
  AOI21X1  g04932(.A0(new_n5933_), .A1(new_n5932_), .B0(new_n5934_), .Y(new_n5935_));
  XOR2X1   g04933(.A(new_n5933_), .B(new_n5932_), .Y(new_n5936_));
  OAI21X1  g04934(.A0(new_n5935_), .A1(new_n5924_), .B0(new_n5936_), .Y(new_n5937_));
  XOR2X1   g04935(.A(new_n5937_), .B(new_n5931_), .Y(new_n5938_));
  NAND2X1  g04936(.A(new_n5938_), .B(new_n5923_), .Y(new_n5939_));
  OR2X1    g04937(.A(new_n5884_), .B(new_n5847_), .Y(new_n5940_));
  XOR2X1   g04938(.A(new_n5841_), .B(new_n5835_), .Y(new_n5941_));
  AND2X1   g04939(.A(new_n5840_), .B(\A[192] ), .Y(new_n5942_));
  OR2X1    g04940(.A(new_n5942_), .B(new_n5842_), .Y(new_n5943_));
  XOR2X1   g04941(.A(new_n5845_), .B(new_n5943_), .Y(new_n5944_));
  OR2X1    g04942(.A(new_n5841_), .B(new_n5835_), .Y(new_n5945_));
  OR2X1    g04943(.A(new_n5845_), .B(new_n5843_), .Y(new_n5946_));
  OAI21X1  g04944(.A0(new_n5945_), .A1(new_n5944_), .B0(new_n5946_), .Y(new_n5947_));
  XOR2X1   g04945(.A(new_n5919_), .B(new_n5944_), .Y(new_n5948_));
  AOI21X1  g04946(.A0(new_n5947_), .A1(new_n5941_), .B0(new_n5948_), .Y(new_n5949_));
  NOR4X1   g04947(.A(new_n5930_), .B(new_n5917_), .C(new_n5929_), .D(new_n5924_), .Y(new_n5950_));
  XOR2X1   g04948(.A(new_n5824_), .B(new_n5928_), .Y(new_n5951_));
  AND2X1   g04949(.A(new_n5823_), .B(\A[198] ), .Y(new_n5952_));
  OR2X1    g04950(.A(new_n5952_), .B(new_n5825_), .Y(new_n5953_));
  XOR2X1   g04951(.A(new_n5828_), .B(new_n5953_), .Y(new_n5954_));
  OR2X1    g04952(.A(new_n5824_), .B(new_n5928_), .Y(new_n5955_));
  OR2X1    g04953(.A(new_n5828_), .B(new_n5826_), .Y(new_n5956_));
  OAI21X1  g04954(.A0(new_n5955_), .A1(new_n5954_), .B0(new_n5956_), .Y(new_n5957_));
  XOR2X1   g04955(.A(new_n5955_), .B(new_n5932_), .Y(new_n5958_));
  AOI21X1  g04956(.A0(new_n5957_), .A1(new_n5951_), .B0(new_n5958_), .Y(new_n5959_));
  OR4X1    g04957(.A(new_n5917_), .B(new_n5929_), .C(new_n5958_), .D(new_n5924_), .Y(new_n5960_));
  OAI22X1  g04958(.A0(new_n5948_), .A1(new_n5921_), .B0(new_n5935_), .B1(new_n5924_), .Y(new_n5961_));
  OAI22X1  g04959(.A0(new_n5961_), .A1(new_n5960_), .B0(new_n5959_), .B1(new_n5950_), .Y(new_n5962_));
  AOI21X1  g04960(.A0(new_n5962_), .A1(new_n5949_), .B0(new_n5940_), .Y(new_n5963_));
  MX2X1    g04961(.A(new_n5962_), .B(new_n5938_), .S0(new_n5923_), .Y(new_n5964_));
  AOI22X1  g04962(.A0(new_n5964_), .A1(new_n5940_), .B0(new_n5963_), .B1(new_n5939_), .Y(new_n5965_));
  INVX1    g04963(.A(\A[176] ), .Y(new_n5966_));
  AND2X1   g04964(.A(new_n5966_), .B(\A[175] ), .Y(new_n5967_));
  OAI21X1  g04965(.A0(new_n5966_), .A1(\A[175] ), .B0(\A[177] ), .Y(new_n5968_));
  NAND2X1  g04966(.A(new_n5871_), .B(new_n5867_), .Y(new_n5969_));
  OAI21X1  g04967(.A0(new_n5968_), .A1(new_n5967_), .B0(new_n5969_), .Y(new_n5970_));
  XOR2X1   g04968(.A(new_n5878_), .B(new_n5970_), .Y(new_n5971_));
  XOR2X1   g04969(.A(new_n5882_), .B(new_n5880_), .Y(new_n5972_));
  NOR2X1   g04970(.A(new_n5878_), .B(new_n5872_), .Y(new_n5973_));
  NOR2X1   g04971(.A(new_n5882_), .B(new_n5880_), .Y(new_n5974_));
  AOI21X1  g04972(.A0(new_n5973_), .A1(new_n5972_), .B0(new_n5974_), .Y(new_n5975_));
  XOR2X1   g04973(.A(new_n5973_), .B(new_n5972_), .Y(new_n5976_));
  OAI21X1  g04974(.A0(new_n5975_), .A1(new_n5971_), .B0(new_n5976_), .Y(new_n5977_));
  XOR2X1   g04975(.A(new_n5861_), .B(new_n5855_), .Y(new_n5978_));
  INVX1    g04976(.A(\A[181] ), .Y(new_n5979_));
  OR2X1    g04977(.A(\A[182] ), .B(new_n5979_), .Y(new_n5980_));
  AOI21X1  g04978(.A0(\A[182] ), .A1(new_n5979_), .B0(new_n5852_), .Y(new_n5981_));
  AOI22X1  g04979(.A0(new_n5853_), .A1(new_n5852_), .B0(new_n5981_), .B1(new_n5980_), .Y(new_n5982_));
  NOR4X1   g04980(.A(new_n5865_), .B(new_n5863_), .C(new_n5861_), .D(new_n5982_), .Y(new_n5983_));
  NOR4X1   g04981(.A(new_n5882_), .B(new_n5880_), .C(new_n5878_), .D(new_n5872_), .Y(new_n5984_));
  OR4X1    g04982(.A(new_n5984_), .B(new_n5971_), .C(new_n5983_), .D(new_n5978_), .Y(new_n5985_));
  XOR2X1   g04983(.A(new_n5861_), .B(new_n5982_), .Y(new_n5986_));
  AND2X1   g04984(.A(new_n5860_), .B(\A[186] ), .Y(new_n5987_));
  OR2X1    g04985(.A(new_n5987_), .B(new_n5862_), .Y(new_n5988_));
  XOR2X1   g04986(.A(new_n5865_), .B(new_n5988_), .Y(new_n5989_));
  OR2X1    g04987(.A(new_n5861_), .B(new_n5982_), .Y(new_n5990_));
  OR2X1    g04988(.A(new_n5865_), .B(new_n5863_), .Y(new_n5991_));
  OAI21X1  g04989(.A0(new_n5990_), .A1(new_n5989_), .B0(new_n5991_), .Y(new_n5992_));
  NOR2X1   g04990(.A(new_n5861_), .B(new_n5982_), .Y(new_n5993_));
  XOR2X1   g04991(.A(new_n5993_), .B(new_n5989_), .Y(new_n5994_));
  AOI21X1  g04992(.A0(new_n5992_), .A1(new_n5986_), .B0(new_n5994_), .Y(new_n5995_));
  XOR2X1   g04993(.A(new_n5995_), .B(new_n5985_), .Y(new_n5996_));
  XOR2X1   g04994(.A(new_n5865_), .B(new_n5863_), .Y(new_n5997_));
  NOR2X1   g04995(.A(new_n5865_), .B(new_n5863_), .Y(new_n5998_));
  AOI21X1  g04996(.A0(new_n5993_), .A1(new_n5997_), .B0(new_n5998_), .Y(new_n5999_));
  XOR2X1   g04997(.A(new_n5993_), .B(new_n5997_), .Y(new_n6000_));
  OAI21X1  g04998(.A0(new_n5999_), .A1(new_n5978_), .B0(new_n6000_), .Y(new_n6001_));
  NOR4X1   g04999(.A(new_n5971_), .B(new_n5994_), .C(new_n5992_), .D(new_n5978_), .Y(new_n6002_));
  AOI21X1  g05000(.A0(new_n5992_), .A1(new_n5986_), .B0(new_n5984_), .Y(new_n6003_));
  AOI22X1  g05001(.A0(new_n6003_), .A1(new_n6002_), .B0(new_n6001_), .B1(new_n5985_), .Y(new_n6004_));
  MX2X1    g05002(.A(new_n6004_), .B(new_n5996_), .S0(new_n5977_), .Y(new_n6005_));
  NOR2X1   g05003(.A(new_n5884_), .B(new_n5847_), .Y(new_n6006_));
  AOI21X1  g05004(.A0(new_n5962_), .A1(new_n5949_), .B0(new_n6006_), .Y(new_n6007_));
  AOI22X1  g05005(.A0(new_n6007_), .A1(new_n5939_), .B0(new_n5964_), .B1(new_n6006_), .Y(new_n6008_));
  MX2X1    g05006(.A(new_n6008_), .B(new_n5965_), .S0(new_n6005_), .Y(new_n6009_));
  OR2X1    g05007(.A(new_n5885_), .B(new_n5811_), .Y(new_n6010_));
  OAI21X1  g05008(.A0(new_n5899_), .A1(new_n5719_), .B0(new_n6010_), .Y(new_n6011_));
  OAI22X1  g05009(.A0(new_n6011_), .A1(new_n5808_), .B0(new_n5910_), .B1(new_n6010_), .Y(new_n6012_));
  MX2X1    g05010(.A(new_n6012_), .B(new_n5911_), .S0(new_n6009_), .Y(new_n6013_));
  INVX1    g05011(.A(\A[237] ), .Y(new_n6014_));
  INVX1    g05012(.A(\A[236] ), .Y(new_n6015_));
  OR2X1    g05013(.A(new_n6015_), .B(\A[235] ), .Y(new_n6016_));
  AOI21X1  g05014(.A0(new_n6015_), .A1(\A[235] ), .B0(new_n6014_), .Y(new_n6017_));
  XOR2X1   g05015(.A(\A[236] ), .B(\A[235] ), .Y(new_n6018_));
  AOI22X1  g05016(.A0(new_n6018_), .A1(new_n6014_), .B0(new_n6017_), .B1(new_n6016_), .Y(new_n6019_));
  INVX1    g05017(.A(\A[240] ), .Y(new_n6020_));
  INVX1    g05018(.A(\A[239] ), .Y(new_n6021_));
  OR2X1    g05019(.A(new_n6021_), .B(\A[238] ), .Y(new_n6022_));
  AOI21X1  g05020(.A0(new_n6021_), .A1(\A[238] ), .B0(new_n6020_), .Y(new_n6023_));
  XOR2X1   g05021(.A(\A[239] ), .B(\A[238] ), .Y(new_n6024_));
  AOI22X1  g05022(.A0(new_n6024_), .A1(new_n6020_), .B0(new_n6023_), .B1(new_n6022_), .Y(new_n6025_));
  OR2X1    g05023(.A(new_n6025_), .B(new_n6019_), .Y(new_n6026_));
  AND2X1   g05024(.A(\A[239] ), .B(\A[238] ), .Y(new_n6027_));
  AND2X1   g05025(.A(new_n6024_), .B(\A[240] ), .Y(new_n6028_));
  OR2X1    g05026(.A(new_n6028_), .B(new_n6027_), .Y(new_n6029_));
  AND2X1   g05027(.A(\A[236] ), .B(\A[235] ), .Y(new_n6030_));
  AOI21X1  g05028(.A0(new_n6018_), .A1(\A[237] ), .B0(new_n6030_), .Y(new_n6031_));
  XOR2X1   g05029(.A(new_n6031_), .B(new_n6029_), .Y(new_n6032_));
  XOR2X1   g05030(.A(new_n6032_), .B(new_n6026_), .Y(new_n6033_));
  INVX1    g05031(.A(\A[235] ), .Y(new_n6034_));
  AND2X1   g05032(.A(\A[236] ), .B(new_n6034_), .Y(new_n6035_));
  OAI21X1  g05033(.A0(\A[236] ), .A1(new_n6034_), .B0(\A[237] ), .Y(new_n6036_));
  NAND2X1  g05034(.A(new_n6018_), .B(new_n6014_), .Y(new_n6037_));
  OAI21X1  g05035(.A0(new_n6036_), .A1(new_n6035_), .B0(new_n6037_), .Y(new_n6038_));
  XOR2X1   g05036(.A(new_n6025_), .B(new_n6038_), .Y(new_n6039_));
  NOR2X1   g05037(.A(new_n6025_), .B(new_n6019_), .Y(new_n6040_));
  AOI21X1  g05038(.A0(new_n6024_), .A1(\A[240] ), .B0(new_n6027_), .Y(new_n6041_));
  XOR2X1   g05039(.A(new_n6031_), .B(new_n6041_), .Y(new_n6042_));
  NOR2X1   g05040(.A(new_n6031_), .B(new_n6041_), .Y(new_n6043_));
  AOI21X1  g05041(.A0(new_n6042_), .A1(new_n6040_), .B0(new_n6043_), .Y(new_n6044_));
  OAI21X1  g05042(.A0(new_n6044_), .A1(new_n6039_), .B0(new_n6033_), .Y(new_n6045_));
  AND2X1   g05043(.A(\A[245] ), .B(\A[244] ), .Y(new_n6046_));
  XOR2X1   g05044(.A(\A[245] ), .B(\A[244] ), .Y(new_n6047_));
  AOI21X1  g05045(.A0(new_n6047_), .A1(\A[246] ), .B0(new_n6046_), .Y(new_n6048_));
  AND2X1   g05046(.A(\A[242] ), .B(\A[241] ), .Y(new_n6049_));
  XOR2X1   g05047(.A(\A[242] ), .B(\A[241] ), .Y(new_n6050_));
  AOI21X1  g05048(.A0(new_n6050_), .A1(\A[243] ), .B0(new_n6049_), .Y(new_n6051_));
  INVX1    g05049(.A(\A[243] ), .Y(new_n6052_));
  INVX1    g05050(.A(\A[242] ), .Y(new_n6053_));
  OR2X1    g05051(.A(new_n6053_), .B(\A[241] ), .Y(new_n6054_));
  AOI21X1  g05052(.A0(new_n6053_), .A1(\A[241] ), .B0(new_n6052_), .Y(new_n6055_));
  AOI22X1  g05053(.A0(new_n6055_), .A1(new_n6054_), .B0(new_n6050_), .B1(new_n6052_), .Y(new_n6056_));
  INVX1    g05054(.A(\A[246] ), .Y(new_n6057_));
  INVX1    g05055(.A(\A[245] ), .Y(new_n6058_));
  OR2X1    g05056(.A(new_n6058_), .B(\A[244] ), .Y(new_n6059_));
  AOI21X1  g05057(.A0(new_n6058_), .A1(\A[244] ), .B0(new_n6057_), .Y(new_n6060_));
  AOI22X1  g05058(.A0(new_n6060_), .A1(new_n6059_), .B0(new_n6047_), .B1(new_n6057_), .Y(new_n6061_));
  NOR4X1   g05059(.A(new_n6061_), .B(new_n6056_), .C(new_n6051_), .D(new_n6048_), .Y(new_n6062_));
  NOR4X1   g05060(.A(new_n6031_), .B(new_n6041_), .C(new_n6025_), .D(new_n6019_), .Y(new_n6063_));
  INVX1    g05061(.A(\A[241] ), .Y(new_n6064_));
  AND2X1   g05062(.A(\A[242] ), .B(new_n6064_), .Y(new_n6065_));
  OAI21X1  g05063(.A0(\A[242] ), .A1(new_n6064_), .B0(\A[243] ), .Y(new_n6066_));
  NAND2X1  g05064(.A(new_n6050_), .B(new_n6052_), .Y(new_n6067_));
  OAI21X1  g05065(.A0(new_n6066_), .A1(new_n6065_), .B0(new_n6067_), .Y(new_n6068_));
  XOR2X1   g05066(.A(new_n6061_), .B(new_n6068_), .Y(new_n6069_));
  OR4X1    g05067(.A(new_n6069_), .B(new_n6063_), .C(new_n6062_), .D(new_n6039_), .Y(new_n6070_));
  XOR2X1   g05068(.A(new_n6051_), .B(new_n6048_), .Y(new_n6071_));
  NOR2X1   g05069(.A(new_n6061_), .B(new_n6056_), .Y(new_n6072_));
  NOR2X1   g05070(.A(new_n6051_), .B(new_n6048_), .Y(new_n6073_));
  AOI21X1  g05071(.A0(new_n6072_), .A1(new_n6071_), .B0(new_n6073_), .Y(new_n6074_));
  XOR2X1   g05072(.A(new_n6072_), .B(new_n6071_), .Y(new_n6075_));
  OAI21X1  g05073(.A0(new_n6069_), .A1(new_n6074_), .B0(new_n6075_), .Y(new_n6076_));
  XOR2X1   g05074(.A(new_n6076_), .B(new_n6070_), .Y(new_n6077_));
  AND2X1   g05075(.A(new_n6077_), .B(new_n6045_), .Y(new_n6078_));
  XOR2X1   g05076(.A(new_n6025_), .B(new_n6019_), .Y(new_n6079_));
  OAI21X1  g05077(.A0(new_n6069_), .A1(new_n6062_), .B0(new_n6079_), .Y(new_n6080_));
  OR4X1    g05078(.A(new_n6061_), .B(new_n6056_), .C(new_n6051_), .D(new_n6048_), .Y(new_n6081_));
  XOR2X1   g05079(.A(new_n6061_), .B(new_n6056_), .Y(new_n6082_));
  XOR2X1   g05080(.A(new_n6025_), .B(new_n6038_), .Y(new_n6083_));
  NAND3X1  g05081(.A(new_n6083_), .B(new_n6082_), .C(new_n6081_), .Y(new_n6084_));
  INVX1    g05082(.A(\A[230] ), .Y(new_n6085_));
  AND2X1   g05083(.A(new_n6085_), .B(\A[229] ), .Y(new_n6086_));
  OAI21X1  g05084(.A0(new_n6085_), .A1(\A[229] ), .B0(\A[231] ), .Y(new_n6087_));
  INVX1    g05085(.A(\A[231] ), .Y(new_n6088_));
  XOR2X1   g05086(.A(\A[230] ), .B(\A[229] ), .Y(new_n6089_));
  NAND2X1  g05087(.A(new_n6089_), .B(new_n6088_), .Y(new_n6090_));
  OAI21X1  g05088(.A0(new_n6087_), .A1(new_n6086_), .B0(new_n6090_), .Y(new_n6091_));
  INVX1    g05089(.A(\A[234] ), .Y(new_n6092_));
  INVX1    g05090(.A(\A[232] ), .Y(new_n6093_));
  OR2X1    g05091(.A(\A[233] ), .B(new_n6093_), .Y(new_n6094_));
  AOI21X1  g05092(.A0(\A[233] ), .A1(new_n6093_), .B0(new_n6092_), .Y(new_n6095_));
  XOR2X1   g05093(.A(\A[233] ), .B(\A[232] ), .Y(new_n6096_));
  AOI22X1  g05094(.A0(new_n6096_), .A1(new_n6092_), .B0(new_n6095_), .B1(new_n6094_), .Y(new_n6097_));
  AND2X1   g05095(.A(\A[233] ), .B(\A[232] ), .Y(new_n6098_));
  AOI21X1  g05096(.A0(new_n6096_), .A1(\A[234] ), .B0(new_n6098_), .Y(new_n6099_));
  AND2X1   g05097(.A(\A[230] ), .B(\A[229] ), .Y(new_n6100_));
  AOI21X1  g05098(.A0(new_n6089_), .A1(\A[231] ), .B0(new_n6100_), .Y(new_n6101_));
  XOR2X1   g05099(.A(new_n6097_), .B(new_n6091_), .Y(new_n6102_));
  INVX1    g05100(.A(\A[225] ), .Y(new_n6103_));
  INVX1    g05101(.A(\A[223] ), .Y(new_n6104_));
  OR2X1    g05102(.A(\A[224] ), .B(new_n6104_), .Y(new_n6105_));
  AOI21X1  g05103(.A0(\A[224] ), .A1(new_n6104_), .B0(new_n6103_), .Y(new_n6106_));
  XOR2X1   g05104(.A(\A[224] ), .B(\A[223] ), .Y(new_n6107_));
  AOI22X1  g05105(.A0(new_n6107_), .A1(new_n6103_), .B0(new_n6106_), .B1(new_n6105_), .Y(new_n6108_));
  INVX1    g05106(.A(\A[228] ), .Y(new_n6109_));
  INVX1    g05107(.A(\A[226] ), .Y(new_n6110_));
  OR2X1    g05108(.A(\A[227] ), .B(new_n6110_), .Y(new_n6111_));
  AOI21X1  g05109(.A0(\A[227] ), .A1(new_n6110_), .B0(new_n6109_), .Y(new_n6112_));
  XOR2X1   g05110(.A(\A[227] ), .B(\A[226] ), .Y(new_n6113_));
  AOI22X1  g05111(.A0(new_n6113_), .A1(new_n6109_), .B0(new_n6112_), .B1(new_n6111_), .Y(new_n6114_));
  AND2X1   g05112(.A(\A[227] ), .B(\A[226] ), .Y(new_n6115_));
  AOI21X1  g05113(.A0(new_n6113_), .A1(\A[228] ), .B0(new_n6115_), .Y(new_n6116_));
  AND2X1   g05114(.A(\A[224] ), .B(\A[223] ), .Y(new_n6117_));
  AOI21X1  g05115(.A0(new_n6107_), .A1(\A[225] ), .B0(new_n6117_), .Y(new_n6118_));
  XOR2X1   g05116(.A(new_n6114_), .B(new_n6108_), .Y(new_n6119_));
  XOR2X1   g05117(.A(new_n6119_), .B(new_n6102_), .Y(new_n6120_));
  AOI21X1  g05118(.A0(new_n6084_), .A1(new_n6080_), .B0(new_n6120_), .Y(new_n6121_));
  AND2X1   g05119(.A(new_n6047_), .B(\A[246] ), .Y(new_n6122_));
  OR2X1    g05120(.A(new_n6122_), .B(new_n6046_), .Y(new_n6123_));
  XOR2X1   g05121(.A(new_n6051_), .B(new_n6123_), .Y(new_n6124_));
  XOR2X1   g05122(.A(new_n6072_), .B(new_n6124_), .Y(new_n6125_));
  NOR4X1   g05123(.A(new_n6069_), .B(new_n6063_), .C(new_n6125_), .D(new_n6039_), .Y(new_n6126_));
  OR2X1    g05124(.A(new_n6061_), .B(new_n6056_), .Y(new_n6127_));
  OR2X1    g05125(.A(new_n6051_), .B(new_n6048_), .Y(new_n6128_));
  OAI21X1  g05126(.A0(new_n6127_), .A1(new_n6124_), .B0(new_n6128_), .Y(new_n6129_));
  OAI21X1  g05127(.A0(new_n6082_), .A1(new_n6075_), .B0(new_n6129_), .Y(new_n6130_));
  AOI22X1  g05128(.A0(new_n6130_), .A1(new_n6126_), .B0(new_n6076_), .B1(new_n6070_), .Y(new_n6131_));
  OAI21X1  g05129(.A0(new_n6131_), .A1(new_n6045_), .B0(new_n6121_), .Y(new_n6132_));
  AOI21X1  g05130(.A0(new_n6082_), .A1(new_n6129_), .B0(new_n6125_), .Y(new_n6133_));
  XOR2X1   g05131(.A(new_n6133_), .B(new_n6070_), .Y(new_n6134_));
  MX2X1    g05132(.A(new_n6131_), .B(new_n6134_), .S0(new_n6045_), .Y(new_n6135_));
  OAI22X1  g05133(.A0(new_n6135_), .A1(new_n6121_), .B0(new_n6132_), .B1(new_n6078_), .Y(new_n6136_));
  INVX1    g05134(.A(\A[224] ), .Y(new_n6137_));
  AND2X1   g05135(.A(new_n6137_), .B(\A[223] ), .Y(new_n6138_));
  OAI21X1  g05136(.A0(new_n6137_), .A1(\A[223] ), .B0(\A[225] ), .Y(new_n6139_));
  NAND2X1  g05137(.A(new_n6107_), .B(new_n6103_), .Y(new_n6140_));
  OAI21X1  g05138(.A0(new_n6139_), .A1(new_n6138_), .B0(new_n6140_), .Y(new_n6141_));
  XOR2X1   g05139(.A(new_n6114_), .B(new_n6141_), .Y(new_n6142_));
  XOR2X1   g05140(.A(new_n6118_), .B(new_n6116_), .Y(new_n6143_));
  NOR2X1   g05141(.A(new_n6114_), .B(new_n6108_), .Y(new_n6144_));
  NOR2X1   g05142(.A(new_n6118_), .B(new_n6116_), .Y(new_n6145_));
  AOI21X1  g05143(.A0(new_n6144_), .A1(new_n6143_), .B0(new_n6145_), .Y(new_n6146_));
  XOR2X1   g05144(.A(new_n6144_), .B(new_n6143_), .Y(new_n6147_));
  OAI21X1  g05145(.A0(new_n6146_), .A1(new_n6142_), .B0(new_n6147_), .Y(new_n6148_));
  XOR2X1   g05146(.A(new_n6097_), .B(new_n6091_), .Y(new_n6149_));
  INVX1    g05147(.A(\A[229] ), .Y(new_n6150_));
  OR2X1    g05148(.A(\A[230] ), .B(new_n6150_), .Y(new_n6151_));
  AOI21X1  g05149(.A0(\A[230] ), .A1(new_n6150_), .B0(new_n6088_), .Y(new_n6152_));
  AOI22X1  g05150(.A0(new_n6089_), .A1(new_n6088_), .B0(new_n6152_), .B1(new_n6151_), .Y(new_n6153_));
  NOR4X1   g05151(.A(new_n6101_), .B(new_n6099_), .C(new_n6097_), .D(new_n6153_), .Y(new_n6154_));
  NOR4X1   g05152(.A(new_n6118_), .B(new_n6116_), .C(new_n6114_), .D(new_n6108_), .Y(new_n6155_));
  OR4X1    g05153(.A(new_n6155_), .B(new_n6142_), .C(new_n6154_), .D(new_n6149_), .Y(new_n6156_));
  XOR2X1   g05154(.A(new_n6097_), .B(new_n6153_), .Y(new_n6157_));
  AND2X1   g05155(.A(new_n6096_), .B(\A[234] ), .Y(new_n6158_));
  OR2X1    g05156(.A(new_n6158_), .B(new_n6098_), .Y(new_n6159_));
  XOR2X1   g05157(.A(new_n6101_), .B(new_n6159_), .Y(new_n6160_));
  OR2X1    g05158(.A(new_n6097_), .B(new_n6153_), .Y(new_n6161_));
  OR2X1    g05159(.A(new_n6101_), .B(new_n6099_), .Y(new_n6162_));
  OAI21X1  g05160(.A0(new_n6161_), .A1(new_n6160_), .B0(new_n6162_), .Y(new_n6163_));
  NOR2X1   g05161(.A(new_n6097_), .B(new_n6153_), .Y(new_n6164_));
  XOR2X1   g05162(.A(new_n6164_), .B(new_n6160_), .Y(new_n6165_));
  AOI21X1  g05163(.A0(new_n6163_), .A1(new_n6157_), .B0(new_n6165_), .Y(new_n6166_));
  XOR2X1   g05164(.A(new_n6166_), .B(new_n6156_), .Y(new_n6167_));
  XOR2X1   g05165(.A(new_n6101_), .B(new_n6099_), .Y(new_n6168_));
  NOR2X1   g05166(.A(new_n6101_), .B(new_n6099_), .Y(new_n6169_));
  AOI21X1  g05167(.A0(new_n6164_), .A1(new_n6168_), .B0(new_n6169_), .Y(new_n6170_));
  XOR2X1   g05168(.A(new_n6164_), .B(new_n6168_), .Y(new_n6171_));
  OAI21X1  g05169(.A0(new_n6170_), .A1(new_n6149_), .B0(new_n6171_), .Y(new_n6172_));
  NOR4X1   g05170(.A(new_n6142_), .B(new_n6165_), .C(new_n6163_), .D(new_n6149_), .Y(new_n6173_));
  AOI21X1  g05171(.A0(new_n6163_), .A1(new_n6157_), .B0(new_n6155_), .Y(new_n6174_));
  AOI22X1  g05172(.A0(new_n6174_), .A1(new_n6173_), .B0(new_n6172_), .B1(new_n6156_), .Y(new_n6175_));
  MX2X1    g05173(.A(new_n6175_), .B(new_n6167_), .S0(new_n6148_), .Y(new_n6176_));
  AND2X1   g05174(.A(new_n6084_), .B(new_n6080_), .Y(new_n6177_));
  OR2X1    g05175(.A(new_n6120_), .B(new_n6177_), .Y(new_n6178_));
  OAI21X1  g05176(.A0(new_n6131_), .A1(new_n6045_), .B0(new_n6178_), .Y(new_n6179_));
  OAI22X1  g05177(.A0(new_n6179_), .A1(new_n6078_), .B0(new_n6135_), .B1(new_n6178_), .Y(new_n6180_));
  MX2X1    g05178(.A(new_n6180_), .B(new_n6136_), .S0(new_n6176_), .Y(new_n6181_));
  INVX1    g05179(.A(\A[249] ), .Y(new_n6182_));
  INVX1    g05180(.A(\A[248] ), .Y(new_n6183_));
  OR2X1    g05181(.A(new_n6183_), .B(\A[247] ), .Y(new_n6184_));
  AOI21X1  g05182(.A0(new_n6183_), .A1(\A[247] ), .B0(new_n6182_), .Y(new_n6185_));
  XOR2X1   g05183(.A(\A[248] ), .B(\A[247] ), .Y(new_n6186_));
  AOI22X1  g05184(.A0(new_n6186_), .A1(new_n6182_), .B0(new_n6185_), .B1(new_n6184_), .Y(new_n6187_));
  INVX1    g05185(.A(\A[252] ), .Y(new_n6188_));
  INVX1    g05186(.A(\A[251] ), .Y(new_n6189_));
  OR2X1    g05187(.A(new_n6189_), .B(\A[250] ), .Y(new_n6190_));
  AOI21X1  g05188(.A0(new_n6189_), .A1(\A[250] ), .B0(new_n6188_), .Y(new_n6191_));
  XOR2X1   g05189(.A(\A[251] ), .B(\A[250] ), .Y(new_n6192_));
  AOI22X1  g05190(.A0(new_n6192_), .A1(new_n6188_), .B0(new_n6191_), .B1(new_n6190_), .Y(new_n6193_));
  OR2X1    g05191(.A(new_n6193_), .B(new_n6187_), .Y(new_n6194_));
  AND2X1   g05192(.A(\A[251] ), .B(\A[250] ), .Y(new_n6195_));
  AND2X1   g05193(.A(new_n6192_), .B(\A[252] ), .Y(new_n6196_));
  OR2X1    g05194(.A(new_n6196_), .B(new_n6195_), .Y(new_n6197_));
  AND2X1   g05195(.A(\A[248] ), .B(\A[247] ), .Y(new_n6198_));
  AOI21X1  g05196(.A0(new_n6186_), .A1(\A[249] ), .B0(new_n6198_), .Y(new_n6199_));
  XOR2X1   g05197(.A(new_n6199_), .B(new_n6197_), .Y(new_n6200_));
  XOR2X1   g05198(.A(new_n6200_), .B(new_n6194_), .Y(new_n6201_));
  INVX1    g05199(.A(\A[247] ), .Y(new_n6202_));
  AND2X1   g05200(.A(\A[248] ), .B(new_n6202_), .Y(new_n6203_));
  OAI21X1  g05201(.A0(\A[248] ), .A1(new_n6202_), .B0(\A[249] ), .Y(new_n6204_));
  NAND2X1  g05202(.A(new_n6186_), .B(new_n6182_), .Y(new_n6205_));
  OAI21X1  g05203(.A0(new_n6204_), .A1(new_n6203_), .B0(new_n6205_), .Y(new_n6206_));
  XOR2X1   g05204(.A(new_n6193_), .B(new_n6206_), .Y(new_n6207_));
  NOR2X1   g05205(.A(new_n6193_), .B(new_n6187_), .Y(new_n6208_));
  AOI21X1  g05206(.A0(new_n6192_), .A1(\A[252] ), .B0(new_n6195_), .Y(new_n6209_));
  XOR2X1   g05207(.A(new_n6199_), .B(new_n6209_), .Y(new_n6210_));
  NOR2X1   g05208(.A(new_n6199_), .B(new_n6209_), .Y(new_n6211_));
  AOI21X1  g05209(.A0(new_n6210_), .A1(new_n6208_), .B0(new_n6211_), .Y(new_n6212_));
  OAI21X1  g05210(.A0(new_n6212_), .A1(new_n6207_), .B0(new_n6201_), .Y(new_n6213_));
  AND2X1   g05211(.A(\A[257] ), .B(\A[256] ), .Y(new_n6214_));
  XOR2X1   g05212(.A(\A[257] ), .B(\A[256] ), .Y(new_n6215_));
  AOI21X1  g05213(.A0(new_n6215_), .A1(\A[258] ), .B0(new_n6214_), .Y(new_n6216_));
  AND2X1   g05214(.A(\A[254] ), .B(\A[253] ), .Y(new_n6217_));
  XOR2X1   g05215(.A(\A[254] ), .B(\A[253] ), .Y(new_n6218_));
  AOI21X1  g05216(.A0(new_n6218_), .A1(\A[255] ), .B0(new_n6217_), .Y(new_n6219_));
  INVX1    g05217(.A(\A[255] ), .Y(new_n6220_));
  INVX1    g05218(.A(\A[254] ), .Y(new_n6221_));
  OR2X1    g05219(.A(new_n6221_), .B(\A[253] ), .Y(new_n6222_));
  AOI21X1  g05220(.A0(new_n6221_), .A1(\A[253] ), .B0(new_n6220_), .Y(new_n6223_));
  AOI22X1  g05221(.A0(new_n6223_), .A1(new_n6222_), .B0(new_n6218_), .B1(new_n6220_), .Y(new_n6224_));
  INVX1    g05222(.A(\A[258] ), .Y(new_n6225_));
  INVX1    g05223(.A(\A[257] ), .Y(new_n6226_));
  OR2X1    g05224(.A(new_n6226_), .B(\A[256] ), .Y(new_n6227_));
  AOI21X1  g05225(.A0(new_n6226_), .A1(\A[256] ), .B0(new_n6225_), .Y(new_n6228_));
  AOI22X1  g05226(.A0(new_n6228_), .A1(new_n6227_), .B0(new_n6215_), .B1(new_n6225_), .Y(new_n6229_));
  NOR4X1   g05227(.A(new_n6229_), .B(new_n6224_), .C(new_n6219_), .D(new_n6216_), .Y(new_n6230_));
  NOR4X1   g05228(.A(new_n6199_), .B(new_n6209_), .C(new_n6193_), .D(new_n6187_), .Y(new_n6231_));
  INVX1    g05229(.A(\A[253] ), .Y(new_n6232_));
  AND2X1   g05230(.A(\A[254] ), .B(new_n6232_), .Y(new_n6233_));
  OAI21X1  g05231(.A0(\A[254] ), .A1(new_n6232_), .B0(\A[255] ), .Y(new_n6234_));
  NAND2X1  g05232(.A(new_n6218_), .B(new_n6220_), .Y(new_n6235_));
  OAI21X1  g05233(.A0(new_n6234_), .A1(new_n6233_), .B0(new_n6235_), .Y(new_n6236_));
  XOR2X1   g05234(.A(new_n6229_), .B(new_n6236_), .Y(new_n6237_));
  NOR4X1   g05235(.A(new_n6237_), .B(new_n6231_), .C(new_n6230_), .D(new_n6207_), .Y(new_n6238_));
  AND2X1   g05236(.A(new_n6215_), .B(\A[258] ), .Y(new_n6239_));
  OR2X1    g05237(.A(new_n6239_), .B(new_n6214_), .Y(new_n6240_));
  XOR2X1   g05238(.A(new_n6219_), .B(new_n6240_), .Y(new_n6241_));
  OR2X1    g05239(.A(new_n6229_), .B(new_n6224_), .Y(new_n6242_));
  OR2X1    g05240(.A(new_n6219_), .B(new_n6216_), .Y(new_n6243_));
  OAI21X1  g05241(.A0(new_n6242_), .A1(new_n6241_), .B0(new_n6243_), .Y(new_n6244_));
  NOR2X1   g05242(.A(new_n6229_), .B(new_n6224_), .Y(new_n6245_));
  XOR2X1   g05243(.A(new_n6245_), .B(new_n6241_), .Y(new_n6246_));
  XOR2X1   g05244(.A(new_n6229_), .B(new_n6224_), .Y(new_n6247_));
  AOI21X1  g05245(.A0(new_n6247_), .A1(new_n6244_), .B0(new_n6246_), .Y(new_n6248_));
  XOR2X1   g05246(.A(new_n6248_), .B(new_n6238_), .Y(new_n6249_));
  OR4X1    g05247(.A(new_n6237_), .B(new_n6231_), .C(new_n6246_), .D(new_n6207_), .Y(new_n6250_));
  XOR2X1   g05248(.A(new_n6219_), .B(new_n6216_), .Y(new_n6251_));
  NOR2X1   g05249(.A(new_n6219_), .B(new_n6216_), .Y(new_n6252_));
  AOI21X1  g05250(.A0(new_n6245_), .A1(new_n6251_), .B0(new_n6252_), .Y(new_n6253_));
  AOI21X1  g05251(.A0(new_n6237_), .A1(new_n6246_), .B0(new_n6253_), .Y(new_n6254_));
  OAI22X1  g05252(.A0(new_n6254_), .A1(new_n6250_), .B0(new_n6248_), .B1(new_n6238_), .Y(new_n6255_));
  MX2X1    g05253(.A(new_n6255_), .B(new_n6249_), .S0(new_n6213_), .Y(new_n6256_));
  INVX1    g05254(.A(\A[261] ), .Y(new_n6257_));
  INVX1    g05255(.A(\A[260] ), .Y(new_n6258_));
  OR2X1    g05256(.A(new_n6258_), .B(\A[259] ), .Y(new_n6259_));
  AOI21X1  g05257(.A0(new_n6258_), .A1(\A[259] ), .B0(new_n6257_), .Y(new_n6260_));
  XOR2X1   g05258(.A(\A[260] ), .B(\A[259] ), .Y(new_n6261_));
  AOI22X1  g05259(.A0(new_n6261_), .A1(new_n6257_), .B0(new_n6260_), .B1(new_n6259_), .Y(new_n6262_));
  INVX1    g05260(.A(\A[264] ), .Y(new_n6263_));
  INVX1    g05261(.A(\A[263] ), .Y(new_n6264_));
  OR2X1    g05262(.A(new_n6264_), .B(\A[262] ), .Y(new_n6265_));
  AOI21X1  g05263(.A0(new_n6264_), .A1(\A[262] ), .B0(new_n6263_), .Y(new_n6266_));
  XOR2X1   g05264(.A(\A[263] ), .B(\A[262] ), .Y(new_n6267_));
  AOI22X1  g05265(.A0(new_n6267_), .A1(new_n6263_), .B0(new_n6266_), .B1(new_n6265_), .Y(new_n6268_));
  OR2X1    g05266(.A(new_n6268_), .B(new_n6262_), .Y(new_n6269_));
  AND2X1   g05267(.A(\A[263] ), .B(\A[262] ), .Y(new_n6270_));
  AND2X1   g05268(.A(new_n6267_), .B(\A[264] ), .Y(new_n6271_));
  OR2X1    g05269(.A(new_n6271_), .B(new_n6270_), .Y(new_n6272_));
  AND2X1   g05270(.A(\A[260] ), .B(\A[259] ), .Y(new_n6273_));
  AOI21X1  g05271(.A0(new_n6261_), .A1(\A[261] ), .B0(new_n6273_), .Y(new_n6274_));
  XOR2X1   g05272(.A(new_n6274_), .B(new_n6272_), .Y(new_n6275_));
  XOR2X1   g05273(.A(new_n6275_), .B(new_n6269_), .Y(new_n6276_));
  INVX1    g05274(.A(\A[259] ), .Y(new_n6277_));
  AND2X1   g05275(.A(\A[260] ), .B(new_n6277_), .Y(new_n6278_));
  OAI21X1  g05276(.A0(\A[260] ), .A1(new_n6277_), .B0(\A[261] ), .Y(new_n6279_));
  NAND2X1  g05277(.A(new_n6261_), .B(new_n6257_), .Y(new_n6280_));
  OAI21X1  g05278(.A0(new_n6279_), .A1(new_n6278_), .B0(new_n6280_), .Y(new_n6281_));
  XOR2X1   g05279(.A(new_n6268_), .B(new_n6281_), .Y(new_n6282_));
  NOR2X1   g05280(.A(new_n6268_), .B(new_n6262_), .Y(new_n6283_));
  AOI21X1  g05281(.A0(new_n6267_), .A1(\A[264] ), .B0(new_n6270_), .Y(new_n6284_));
  XOR2X1   g05282(.A(new_n6274_), .B(new_n6284_), .Y(new_n6285_));
  NOR2X1   g05283(.A(new_n6274_), .B(new_n6284_), .Y(new_n6286_));
  AOI21X1  g05284(.A0(new_n6285_), .A1(new_n6283_), .B0(new_n6286_), .Y(new_n6287_));
  OAI21X1  g05285(.A0(new_n6287_), .A1(new_n6282_), .B0(new_n6276_), .Y(new_n6288_));
  AND2X1   g05286(.A(\A[269] ), .B(\A[268] ), .Y(new_n6289_));
  XOR2X1   g05287(.A(\A[269] ), .B(\A[268] ), .Y(new_n6290_));
  AOI21X1  g05288(.A0(new_n6290_), .A1(\A[270] ), .B0(new_n6289_), .Y(new_n6291_));
  AND2X1   g05289(.A(\A[266] ), .B(\A[265] ), .Y(new_n6292_));
  XOR2X1   g05290(.A(\A[266] ), .B(\A[265] ), .Y(new_n6293_));
  AOI21X1  g05291(.A0(new_n6293_), .A1(\A[267] ), .B0(new_n6292_), .Y(new_n6294_));
  INVX1    g05292(.A(\A[267] ), .Y(new_n6295_));
  INVX1    g05293(.A(\A[266] ), .Y(new_n6296_));
  OR2X1    g05294(.A(new_n6296_), .B(\A[265] ), .Y(new_n6297_));
  AOI21X1  g05295(.A0(new_n6296_), .A1(\A[265] ), .B0(new_n6295_), .Y(new_n6298_));
  AOI22X1  g05296(.A0(new_n6298_), .A1(new_n6297_), .B0(new_n6293_), .B1(new_n6295_), .Y(new_n6299_));
  INVX1    g05297(.A(\A[270] ), .Y(new_n6300_));
  INVX1    g05298(.A(\A[269] ), .Y(new_n6301_));
  OR2X1    g05299(.A(new_n6301_), .B(\A[268] ), .Y(new_n6302_));
  AOI21X1  g05300(.A0(new_n6301_), .A1(\A[268] ), .B0(new_n6300_), .Y(new_n6303_));
  AOI22X1  g05301(.A0(new_n6303_), .A1(new_n6302_), .B0(new_n6290_), .B1(new_n6300_), .Y(new_n6304_));
  NOR4X1   g05302(.A(new_n6304_), .B(new_n6299_), .C(new_n6294_), .D(new_n6291_), .Y(new_n6305_));
  NOR4X1   g05303(.A(new_n6274_), .B(new_n6284_), .C(new_n6268_), .D(new_n6262_), .Y(new_n6306_));
  INVX1    g05304(.A(\A[265] ), .Y(new_n6307_));
  AND2X1   g05305(.A(\A[266] ), .B(new_n6307_), .Y(new_n6308_));
  OAI21X1  g05306(.A0(\A[266] ), .A1(new_n6307_), .B0(\A[267] ), .Y(new_n6309_));
  NAND2X1  g05307(.A(new_n6293_), .B(new_n6295_), .Y(new_n6310_));
  OAI21X1  g05308(.A0(new_n6309_), .A1(new_n6308_), .B0(new_n6310_), .Y(new_n6311_));
  XOR2X1   g05309(.A(new_n6304_), .B(new_n6311_), .Y(new_n6312_));
  OR4X1    g05310(.A(new_n6312_), .B(new_n6306_), .C(new_n6305_), .D(new_n6282_), .Y(new_n6313_));
  XOR2X1   g05311(.A(new_n6294_), .B(new_n6291_), .Y(new_n6314_));
  NOR2X1   g05312(.A(new_n6304_), .B(new_n6299_), .Y(new_n6315_));
  NOR2X1   g05313(.A(new_n6294_), .B(new_n6291_), .Y(new_n6316_));
  AOI21X1  g05314(.A0(new_n6315_), .A1(new_n6314_), .B0(new_n6316_), .Y(new_n6317_));
  XOR2X1   g05315(.A(new_n6315_), .B(new_n6314_), .Y(new_n6318_));
  OAI21X1  g05316(.A0(new_n6312_), .A1(new_n6317_), .B0(new_n6318_), .Y(new_n6319_));
  XOR2X1   g05317(.A(new_n6319_), .B(new_n6313_), .Y(new_n6320_));
  NAND2X1  g05318(.A(new_n6320_), .B(new_n6288_), .Y(new_n6321_));
  OR2X1    g05319(.A(new_n6312_), .B(new_n6305_), .Y(new_n6322_));
  XOR2X1   g05320(.A(new_n6268_), .B(new_n6262_), .Y(new_n6323_));
  XOR2X1   g05321(.A(new_n6323_), .B(new_n6322_), .Y(new_n6324_));
  OR2X1    g05322(.A(new_n6237_), .B(new_n6230_), .Y(new_n6325_));
  XOR2X1   g05323(.A(new_n6193_), .B(new_n6187_), .Y(new_n6326_));
  XOR2X1   g05324(.A(new_n6326_), .B(new_n6325_), .Y(new_n6327_));
  OR2X1    g05325(.A(new_n6327_), .B(new_n6324_), .Y(new_n6328_));
  XOR2X1   g05326(.A(new_n6275_), .B(new_n6283_), .Y(new_n6329_));
  XOR2X1   g05327(.A(new_n6268_), .B(new_n6262_), .Y(new_n6330_));
  OR2X1    g05328(.A(new_n6274_), .B(new_n6284_), .Y(new_n6331_));
  OAI21X1  g05329(.A0(new_n6275_), .A1(new_n6269_), .B0(new_n6331_), .Y(new_n6332_));
  AOI21X1  g05330(.A0(new_n6332_), .A1(new_n6330_), .B0(new_n6329_), .Y(new_n6333_));
  NOR4X1   g05331(.A(new_n6312_), .B(new_n6306_), .C(new_n6305_), .D(new_n6282_), .Y(new_n6334_));
  AND2X1   g05332(.A(new_n6290_), .B(\A[270] ), .Y(new_n6335_));
  OR2X1    g05333(.A(new_n6335_), .B(new_n6289_), .Y(new_n6336_));
  XOR2X1   g05334(.A(new_n6294_), .B(new_n6336_), .Y(new_n6337_));
  OR2X1    g05335(.A(new_n6304_), .B(new_n6299_), .Y(new_n6338_));
  OR2X1    g05336(.A(new_n6294_), .B(new_n6291_), .Y(new_n6339_));
  OAI21X1  g05337(.A0(new_n6338_), .A1(new_n6337_), .B0(new_n6339_), .Y(new_n6340_));
  XOR2X1   g05338(.A(new_n6315_), .B(new_n6337_), .Y(new_n6341_));
  XOR2X1   g05339(.A(new_n6304_), .B(new_n6299_), .Y(new_n6342_));
  AOI21X1  g05340(.A0(new_n6342_), .A1(new_n6340_), .B0(new_n6341_), .Y(new_n6343_));
  OR4X1    g05341(.A(new_n6312_), .B(new_n6306_), .C(new_n6341_), .D(new_n6282_), .Y(new_n6344_));
  AOI21X1  g05342(.A0(new_n6312_), .A1(new_n6341_), .B0(new_n6317_), .Y(new_n6345_));
  OAI22X1  g05343(.A0(new_n6345_), .A1(new_n6344_), .B0(new_n6343_), .B1(new_n6334_), .Y(new_n6346_));
  AOI21X1  g05344(.A0(new_n6346_), .A1(new_n6333_), .B0(new_n6328_), .Y(new_n6347_));
  MX2X1    g05345(.A(new_n6346_), .B(new_n6320_), .S0(new_n6288_), .Y(new_n6348_));
  AOI22X1  g05346(.A0(new_n6348_), .A1(new_n6328_), .B0(new_n6347_), .B1(new_n6321_), .Y(new_n6349_));
  OR2X1    g05347(.A(new_n6349_), .B(new_n6256_), .Y(new_n6350_));
  XOR2X1   g05348(.A(new_n6268_), .B(new_n6281_), .Y(new_n6351_));
  XOR2X1   g05349(.A(new_n6351_), .B(new_n6322_), .Y(new_n6352_));
  XOR2X1   g05350(.A(new_n6327_), .B(new_n6352_), .Y(new_n6353_));
  INVX1    g05351(.A(new_n6120_), .Y(new_n6354_));
  XOR2X1   g05352(.A(new_n6354_), .B(new_n6177_), .Y(new_n6355_));
  OR2X1    g05353(.A(new_n6355_), .B(new_n6353_), .Y(new_n6356_));
  AND2X1   g05354(.A(new_n6320_), .B(new_n6288_), .Y(new_n6357_));
  XOR2X1   g05355(.A(new_n6343_), .B(new_n6313_), .Y(new_n6358_));
  NOR4X1   g05356(.A(new_n6312_), .B(new_n6306_), .C(new_n6341_), .D(new_n6282_), .Y(new_n6359_));
  OAI21X1  g05357(.A0(new_n6342_), .A1(new_n6318_), .B0(new_n6340_), .Y(new_n6360_));
  AOI22X1  g05358(.A0(new_n6360_), .A1(new_n6359_), .B0(new_n6319_), .B1(new_n6313_), .Y(new_n6361_));
  MX2X1    g05359(.A(new_n6361_), .B(new_n6358_), .S0(new_n6288_), .Y(new_n6362_));
  OAI21X1  g05360(.A0(new_n6361_), .A1(new_n6288_), .B0(new_n6328_), .Y(new_n6363_));
  OAI22X1  g05361(.A0(new_n6363_), .A1(new_n6357_), .B0(new_n6362_), .B1(new_n6328_), .Y(new_n6364_));
  AOI21X1  g05362(.A0(new_n6364_), .A1(new_n6256_), .B0(new_n6356_), .Y(new_n6365_));
  NOR2X1   g05363(.A(new_n6327_), .B(new_n6324_), .Y(new_n6366_));
  OAI21X1  g05364(.A0(new_n6361_), .A1(new_n6288_), .B0(new_n6366_), .Y(new_n6367_));
  OAI22X1  g05365(.A0(new_n6362_), .A1(new_n6366_), .B0(new_n6367_), .B1(new_n6357_), .Y(new_n6368_));
  MX2X1    g05366(.A(new_n6368_), .B(new_n6364_), .S0(new_n6256_), .Y(new_n6369_));
  AOI22X1  g05367(.A0(new_n6369_), .A1(new_n6356_), .B0(new_n6365_), .B1(new_n6350_), .Y(new_n6370_));
  OR2X1    g05368(.A(new_n6370_), .B(new_n6181_), .Y(new_n6371_));
  XOR2X1   g05369(.A(new_n6355_), .B(new_n6353_), .Y(new_n6372_));
  INVX1    g05370(.A(new_n6372_), .Y(new_n6373_));
  XOR2X1   g05371(.A(new_n5884_), .B(new_n5847_), .Y(new_n6374_));
  XOR2X1   g05372(.A(new_n6374_), .B(new_n5811_), .Y(new_n6375_));
  OR2X1    g05373(.A(new_n6375_), .B(new_n6373_), .Y(new_n6376_));
  OR4X1    g05374(.A(new_n6237_), .B(new_n6231_), .C(new_n6230_), .D(new_n6207_), .Y(new_n6377_));
  XOR2X1   g05375(.A(new_n6248_), .B(new_n6377_), .Y(new_n6378_));
  XOR2X1   g05376(.A(new_n6245_), .B(new_n6251_), .Y(new_n6379_));
  OAI21X1  g05377(.A0(new_n6237_), .A1(new_n6253_), .B0(new_n6379_), .Y(new_n6380_));
  NOR4X1   g05378(.A(new_n6237_), .B(new_n6231_), .C(new_n6246_), .D(new_n6207_), .Y(new_n6381_));
  OAI21X1  g05379(.A0(new_n6247_), .A1(new_n6379_), .B0(new_n6244_), .Y(new_n6382_));
  AOI22X1  g05380(.A0(new_n6382_), .A1(new_n6381_), .B0(new_n6380_), .B1(new_n6377_), .Y(new_n6383_));
  MX2X1    g05381(.A(new_n6383_), .B(new_n6378_), .S0(new_n6213_), .Y(new_n6384_));
  AND2X1   g05382(.A(new_n6368_), .B(new_n6384_), .Y(new_n6385_));
  AOI21X1  g05383(.A0(new_n6346_), .A1(new_n6333_), .B0(new_n6366_), .Y(new_n6386_));
  AOI22X1  g05384(.A0(new_n6386_), .A1(new_n6321_), .B0(new_n6348_), .B1(new_n6366_), .Y(new_n6387_));
  MX2X1    g05385(.A(new_n6349_), .B(new_n6387_), .S0(new_n6256_), .Y(new_n6388_));
  OAI21X1  g05386(.A0(new_n6387_), .A1(new_n6384_), .B0(new_n6356_), .Y(new_n6389_));
  OAI22X1  g05387(.A0(new_n6389_), .A1(new_n6385_), .B0(new_n6388_), .B1(new_n6356_), .Y(new_n6390_));
  AOI21X1  g05388(.A0(new_n6390_), .A1(new_n6181_), .B0(new_n6376_), .Y(new_n6391_));
  NAND2X1  g05389(.A(new_n6077_), .B(new_n6045_), .Y(new_n6392_));
  XOR2X1   g05390(.A(new_n6032_), .B(new_n6040_), .Y(new_n6393_));
  XOR2X1   g05391(.A(new_n6025_), .B(new_n6019_), .Y(new_n6394_));
  OR2X1    g05392(.A(new_n6031_), .B(new_n6041_), .Y(new_n6395_));
  OAI21X1  g05393(.A0(new_n6032_), .A1(new_n6026_), .B0(new_n6395_), .Y(new_n6396_));
  AOI21X1  g05394(.A0(new_n6396_), .A1(new_n6394_), .B0(new_n6393_), .Y(new_n6397_));
  NOR4X1   g05395(.A(new_n6069_), .B(new_n6063_), .C(new_n6062_), .D(new_n6039_), .Y(new_n6398_));
  OR4X1    g05396(.A(new_n6069_), .B(new_n6063_), .C(new_n6125_), .D(new_n6039_), .Y(new_n6399_));
  AOI21X1  g05397(.A0(new_n6069_), .A1(new_n6125_), .B0(new_n6074_), .Y(new_n6400_));
  OAI22X1  g05398(.A0(new_n6400_), .A1(new_n6399_), .B0(new_n6133_), .B1(new_n6398_), .Y(new_n6401_));
  AOI21X1  g05399(.A0(new_n6401_), .A1(new_n6397_), .B0(new_n6178_), .Y(new_n6402_));
  MX2X1    g05400(.A(new_n6401_), .B(new_n6077_), .S0(new_n6045_), .Y(new_n6403_));
  AOI22X1  g05401(.A0(new_n6403_), .A1(new_n6178_), .B0(new_n6402_), .B1(new_n6392_), .Y(new_n6404_));
  AOI21X1  g05402(.A0(new_n6401_), .A1(new_n6397_), .B0(new_n6121_), .Y(new_n6405_));
  AOI22X1  g05403(.A0(new_n6405_), .A1(new_n6392_), .B0(new_n6403_), .B1(new_n6121_), .Y(new_n6406_));
  MX2X1    g05404(.A(new_n6406_), .B(new_n6404_), .S0(new_n6176_), .Y(new_n6407_));
  NOR2X1   g05405(.A(new_n6355_), .B(new_n6353_), .Y(new_n6408_));
  OAI21X1  g05406(.A0(new_n6387_), .A1(new_n6384_), .B0(new_n6408_), .Y(new_n6409_));
  OAI22X1  g05407(.A0(new_n6388_), .A1(new_n6408_), .B0(new_n6409_), .B1(new_n6385_), .Y(new_n6410_));
  MX2X1    g05408(.A(new_n6390_), .B(new_n6410_), .S0(new_n6407_), .Y(new_n6411_));
  AOI22X1  g05409(.A0(new_n6411_), .A1(new_n6376_), .B0(new_n6391_), .B1(new_n6371_), .Y(new_n6412_));
  OR2X1    g05410(.A(new_n6412_), .B(new_n6013_), .Y(new_n6413_));
  XOR2X1   g05411(.A(new_n6375_), .B(new_n6372_), .Y(new_n6414_));
  INVX1    g05412(.A(\A[170] ), .Y(new_n6415_));
  AND2X1   g05413(.A(new_n6415_), .B(\A[169] ), .Y(new_n6416_));
  OAI21X1  g05414(.A0(new_n6415_), .A1(\A[169] ), .B0(\A[171] ), .Y(new_n6417_));
  INVX1    g05415(.A(\A[171] ), .Y(new_n6418_));
  XOR2X1   g05416(.A(\A[170] ), .B(\A[169] ), .Y(new_n6419_));
  NAND2X1  g05417(.A(new_n6419_), .B(new_n6418_), .Y(new_n6420_));
  OAI21X1  g05418(.A0(new_n6417_), .A1(new_n6416_), .B0(new_n6420_), .Y(new_n6421_));
  INVX1    g05419(.A(\A[174] ), .Y(new_n6422_));
  INVX1    g05420(.A(\A[172] ), .Y(new_n6423_));
  OR2X1    g05421(.A(\A[173] ), .B(new_n6423_), .Y(new_n6424_));
  AOI21X1  g05422(.A0(\A[173] ), .A1(new_n6423_), .B0(new_n6422_), .Y(new_n6425_));
  XOR2X1   g05423(.A(\A[173] ), .B(\A[172] ), .Y(new_n6426_));
  AOI22X1  g05424(.A0(new_n6426_), .A1(new_n6422_), .B0(new_n6425_), .B1(new_n6424_), .Y(new_n6427_));
  AND2X1   g05425(.A(\A[173] ), .B(\A[172] ), .Y(new_n6428_));
  AOI21X1  g05426(.A0(new_n6426_), .A1(\A[174] ), .B0(new_n6428_), .Y(new_n6429_));
  AND2X1   g05427(.A(\A[170] ), .B(\A[169] ), .Y(new_n6430_));
  AOI21X1  g05428(.A0(new_n6419_), .A1(\A[171] ), .B0(new_n6430_), .Y(new_n6431_));
  XOR2X1   g05429(.A(new_n6427_), .B(new_n6421_), .Y(new_n6432_));
  INVX1    g05430(.A(\A[165] ), .Y(new_n6433_));
  INVX1    g05431(.A(\A[163] ), .Y(new_n6434_));
  OR2X1    g05432(.A(\A[164] ), .B(new_n6434_), .Y(new_n6435_));
  AOI21X1  g05433(.A0(\A[164] ), .A1(new_n6434_), .B0(new_n6433_), .Y(new_n6436_));
  XOR2X1   g05434(.A(\A[164] ), .B(\A[163] ), .Y(new_n6437_));
  AOI22X1  g05435(.A0(new_n6437_), .A1(new_n6433_), .B0(new_n6436_), .B1(new_n6435_), .Y(new_n6438_));
  INVX1    g05436(.A(\A[168] ), .Y(new_n6439_));
  INVX1    g05437(.A(\A[166] ), .Y(new_n6440_));
  OR2X1    g05438(.A(\A[167] ), .B(new_n6440_), .Y(new_n6441_));
  AOI21X1  g05439(.A0(\A[167] ), .A1(new_n6440_), .B0(new_n6439_), .Y(new_n6442_));
  XOR2X1   g05440(.A(\A[167] ), .B(\A[166] ), .Y(new_n6443_));
  AOI22X1  g05441(.A0(new_n6443_), .A1(new_n6439_), .B0(new_n6442_), .B1(new_n6441_), .Y(new_n6444_));
  AND2X1   g05442(.A(\A[167] ), .B(\A[166] ), .Y(new_n6445_));
  AOI21X1  g05443(.A0(new_n6443_), .A1(\A[168] ), .B0(new_n6445_), .Y(new_n6446_));
  AND2X1   g05444(.A(\A[164] ), .B(\A[163] ), .Y(new_n6447_));
  AOI21X1  g05445(.A0(new_n6437_), .A1(\A[165] ), .B0(new_n6447_), .Y(new_n6448_));
  XOR2X1   g05446(.A(new_n6444_), .B(new_n6438_), .Y(new_n6449_));
  XOR2X1   g05447(.A(new_n6449_), .B(new_n6432_), .Y(new_n6450_));
  INVX1    g05448(.A(\A[158] ), .Y(new_n6451_));
  AND2X1   g05449(.A(new_n6451_), .B(\A[157] ), .Y(new_n6452_));
  OAI21X1  g05450(.A0(new_n6451_), .A1(\A[157] ), .B0(\A[159] ), .Y(new_n6453_));
  INVX1    g05451(.A(\A[159] ), .Y(new_n6454_));
  XOR2X1   g05452(.A(\A[158] ), .B(\A[157] ), .Y(new_n6455_));
  NAND2X1  g05453(.A(new_n6455_), .B(new_n6454_), .Y(new_n6456_));
  OAI21X1  g05454(.A0(new_n6453_), .A1(new_n6452_), .B0(new_n6456_), .Y(new_n6457_));
  INVX1    g05455(.A(\A[162] ), .Y(new_n6458_));
  INVX1    g05456(.A(\A[160] ), .Y(new_n6459_));
  OR2X1    g05457(.A(\A[161] ), .B(new_n6459_), .Y(new_n6460_));
  AOI21X1  g05458(.A0(\A[161] ), .A1(new_n6459_), .B0(new_n6458_), .Y(new_n6461_));
  XOR2X1   g05459(.A(\A[161] ), .B(\A[160] ), .Y(new_n6462_));
  AOI22X1  g05460(.A0(new_n6462_), .A1(new_n6458_), .B0(new_n6461_), .B1(new_n6460_), .Y(new_n6463_));
  AND2X1   g05461(.A(\A[161] ), .B(\A[160] ), .Y(new_n6464_));
  AOI21X1  g05462(.A0(new_n6462_), .A1(\A[162] ), .B0(new_n6464_), .Y(new_n6465_));
  AND2X1   g05463(.A(\A[158] ), .B(\A[157] ), .Y(new_n6466_));
  AOI21X1  g05464(.A0(new_n6455_), .A1(\A[159] ), .B0(new_n6466_), .Y(new_n6467_));
  XOR2X1   g05465(.A(new_n6463_), .B(new_n6457_), .Y(new_n6468_));
  INVX1    g05466(.A(\A[153] ), .Y(new_n6469_));
  INVX1    g05467(.A(\A[151] ), .Y(new_n6470_));
  OR2X1    g05468(.A(\A[152] ), .B(new_n6470_), .Y(new_n6471_));
  AOI21X1  g05469(.A0(\A[152] ), .A1(new_n6470_), .B0(new_n6469_), .Y(new_n6472_));
  XOR2X1   g05470(.A(\A[152] ), .B(\A[151] ), .Y(new_n6473_));
  AOI22X1  g05471(.A0(new_n6473_), .A1(new_n6469_), .B0(new_n6472_), .B1(new_n6471_), .Y(new_n6474_));
  INVX1    g05472(.A(\A[156] ), .Y(new_n6475_));
  INVX1    g05473(.A(\A[154] ), .Y(new_n6476_));
  OR2X1    g05474(.A(\A[155] ), .B(new_n6476_), .Y(new_n6477_));
  AOI21X1  g05475(.A0(\A[155] ), .A1(new_n6476_), .B0(new_n6475_), .Y(new_n6478_));
  XOR2X1   g05476(.A(\A[155] ), .B(\A[154] ), .Y(new_n6479_));
  AOI22X1  g05477(.A0(new_n6479_), .A1(new_n6475_), .B0(new_n6478_), .B1(new_n6477_), .Y(new_n6480_));
  AND2X1   g05478(.A(\A[155] ), .B(\A[154] ), .Y(new_n6481_));
  AOI21X1  g05479(.A0(new_n6479_), .A1(\A[156] ), .B0(new_n6481_), .Y(new_n6482_));
  AND2X1   g05480(.A(\A[152] ), .B(\A[151] ), .Y(new_n6483_));
  AOI21X1  g05481(.A0(new_n6473_), .A1(\A[153] ), .B0(new_n6483_), .Y(new_n6484_));
  XOR2X1   g05482(.A(new_n6480_), .B(new_n6474_), .Y(new_n6485_));
  XOR2X1   g05483(.A(new_n6485_), .B(new_n6468_), .Y(new_n6486_));
  XOR2X1   g05484(.A(new_n6486_), .B(new_n6450_), .Y(new_n6487_));
  INVX1    g05485(.A(\A[146] ), .Y(new_n6488_));
  AND2X1   g05486(.A(new_n6488_), .B(\A[145] ), .Y(new_n6489_));
  OAI21X1  g05487(.A0(new_n6488_), .A1(\A[145] ), .B0(\A[147] ), .Y(new_n6490_));
  INVX1    g05488(.A(\A[147] ), .Y(new_n6491_));
  XOR2X1   g05489(.A(\A[146] ), .B(\A[145] ), .Y(new_n6492_));
  NAND2X1  g05490(.A(new_n6492_), .B(new_n6491_), .Y(new_n6493_));
  OAI21X1  g05491(.A0(new_n6490_), .A1(new_n6489_), .B0(new_n6493_), .Y(new_n6494_));
  INVX1    g05492(.A(\A[150] ), .Y(new_n6495_));
  INVX1    g05493(.A(\A[148] ), .Y(new_n6496_));
  OR2X1    g05494(.A(\A[149] ), .B(new_n6496_), .Y(new_n6497_));
  AOI21X1  g05495(.A0(\A[149] ), .A1(new_n6496_), .B0(new_n6495_), .Y(new_n6498_));
  XOR2X1   g05496(.A(\A[149] ), .B(\A[148] ), .Y(new_n6499_));
  AOI22X1  g05497(.A0(new_n6499_), .A1(new_n6495_), .B0(new_n6498_), .B1(new_n6497_), .Y(new_n6500_));
  AND2X1   g05498(.A(\A[149] ), .B(\A[148] ), .Y(new_n6501_));
  AOI21X1  g05499(.A0(new_n6499_), .A1(\A[150] ), .B0(new_n6501_), .Y(new_n6502_));
  AND2X1   g05500(.A(\A[146] ), .B(\A[145] ), .Y(new_n6503_));
  AOI21X1  g05501(.A0(new_n6492_), .A1(\A[147] ), .B0(new_n6503_), .Y(new_n6504_));
  XOR2X1   g05502(.A(new_n6500_), .B(new_n6494_), .Y(new_n6505_));
  INVX1    g05503(.A(\A[141] ), .Y(new_n6506_));
  INVX1    g05504(.A(\A[139] ), .Y(new_n6507_));
  OR2X1    g05505(.A(\A[140] ), .B(new_n6507_), .Y(new_n6508_));
  AOI21X1  g05506(.A0(\A[140] ), .A1(new_n6507_), .B0(new_n6506_), .Y(new_n6509_));
  XOR2X1   g05507(.A(\A[140] ), .B(\A[139] ), .Y(new_n6510_));
  AOI22X1  g05508(.A0(new_n6510_), .A1(new_n6506_), .B0(new_n6509_), .B1(new_n6508_), .Y(new_n6511_));
  INVX1    g05509(.A(\A[144] ), .Y(new_n6512_));
  INVX1    g05510(.A(\A[142] ), .Y(new_n6513_));
  OR2X1    g05511(.A(\A[143] ), .B(new_n6513_), .Y(new_n6514_));
  AOI21X1  g05512(.A0(\A[143] ), .A1(new_n6513_), .B0(new_n6512_), .Y(new_n6515_));
  XOR2X1   g05513(.A(\A[143] ), .B(\A[142] ), .Y(new_n6516_));
  AOI22X1  g05514(.A0(new_n6516_), .A1(new_n6512_), .B0(new_n6515_), .B1(new_n6514_), .Y(new_n6517_));
  AND2X1   g05515(.A(\A[143] ), .B(\A[142] ), .Y(new_n6518_));
  AOI21X1  g05516(.A0(new_n6516_), .A1(\A[144] ), .B0(new_n6518_), .Y(new_n6519_));
  AND2X1   g05517(.A(\A[140] ), .B(\A[139] ), .Y(new_n6520_));
  AOI21X1  g05518(.A0(new_n6510_), .A1(\A[141] ), .B0(new_n6520_), .Y(new_n6521_));
  XOR2X1   g05519(.A(new_n6517_), .B(new_n6511_), .Y(new_n6522_));
  XOR2X1   g05520(.A(new_n6522_), .B(new_n6505_), .Y(new_n6523_));
  INVX1    g05521(.A(new_n6523_), .Y(new_n6524_));
  INVX1    g05522(.A(\A[134] ), .Y(new_n6525_));
  AND2X1   g05523(.A(new_n6525_), .B(\A[133] ), .Y(new_n6526_));
  OAI21X1  g05524(.A0(new_n6525_), .A1(\A[133] ), .B0(\A[135] ), .Y(new_n6527_));
  INVX1    g05525(.A(\A[135] ), .Y(new_n6528_));
  XOR2X1   g05526(.A(\A[134] ), .B(\A[133] ), .Y(new_n6529_));
  NAND2X1  g05527(.A(new_n6529_), .B(new_n6528_), .Y(new_n6530_));
  OAI21X1  g05528(.A0(new_n6527_), .A1(new_n6526_), .B0(new_n6530_), .Y(new_n6531_));
  INVX1    g05529(.A(\A[138] ), .Y(new_n6532_));
  INVX1    g05530(.A(\A[136] ), .Y(new_n6533_));
  OR2X1    g05531(.A(\A[137] ), .B(new_n6533_), .Y(new_n6534_));
  AOI21X1  g05532(.A0(\A[137] ), .A1(new_n6533_), .B0(new_n6532_), .Y(new_n6535_));
  XOR2X1   g05533(.A(\A[137] ), .B(\A[136] ), .Y(new_n6536_));
  AOI22X1  g05534(.A0(new_n6536_), .A1(new_n6532_), .B0(new_n6535_), .B1(new_n6534_), .Y(new_n6537_));
  AND2X1   g05535(.A(\A[137] ), .B(\A[136] ), .Y(new_n6538_));
  AOI21X1  g05536(.A0(new_n6536_), .A1(\A[138] ), .B0(new_n6538_), .Y(new_n6539_));
  AND2X1   g05537(.A(\A[134] ), .B(\A[133] ), .Y(new_n6540_));
  AOI21X1  g05538(.A0(new_n6529_), .A1(\A[135] ), .B0(new_n6540_), .Y(new_n6541_));
  XOR2X1   g05539(.A(new_n6537_), .B(new_n6531_), .Y(new_n6542_));
  INVX1    g05540(.A(\A[129] ), .Y(new_n6543_));
  INVX1    g05541(.A(\A[127] ), .Y(new_n6544_));
  OR2X1    g05542(.A(\A[128] ), .B(new_n6544_), .Y(new_n6545_));
  AOI21X1  g05543(.A0(\A[128] ), .A1(new_n6544_), .B0(new_n6543_), .Y(new_n6546_));
  XOR2X1   g05544(.A(\A[128] ), .B(\A[127] ), .Y(new_n6547_));
  AOI22X1  g05545(.A0(new_n6547_), .A1(new_n6543_), .B0(new_n6546_), .B1(new_n6545_), .Y(new_n6548_));
  INVX1    g05546(.A(\A[132] ), .Y(new_n6549_));
  INVX1    g05547(.A(\A[130] ), .Y(new_n6550_));
  OR2X1    g05548(.A(\A[131] ), .B(new_n6550_), .Y(new_n6551_));
  AOI21X1  g05549(.A0(\A[131] ), .A1(new_n6550_), .B0(new_n6549_), .Y(new_n6552_));
  XOR2X1   g05550(.A(\A[131] ), .B(\A[130] ), .Y(new_n6553_));
  AOI22X1  g05551(.A0(new_n6553_), .A1(new_n6549_), .B0(new_n6552_), .B1(new_n6551_), .Y(new_n6554_));
  AND2X1   g05552(.A(\A[131] ), .B(\A[130] ), .Y(new_n6555_));
  AOI21X1  g05553(.A0(new_n6553_), .A1(\A[132] ), .B0(new_n6555_), .Y(new_n6556_));
  AND2X1   g05554(.A(\A[128] ), .B(\A[127] ), .Y(new_n6557_));
  AOI21X1  g05555(.A0(new_n6547_), .A1(\A[129] ), .B0(new_n6557_), .Y(new_n6558_));
  XOR2X1   g05556(.A(new_n6554_), .B(new_n6548_), .Y(new_n6559_));
  XOR2X1   g05557(.A(new_n6559_), .B(new_n6542_), .Y(new_n6560_));
  XOR2X1   g05558(.A(new_n6560_), .B(new_n6524_), .Y(new_n6561_));
  XOR2X1   g05559(.A(new_n6561_), .B(new_n6487_), .Y(new_n6562_));
  INVX1    g05560(.A(\A[122] ), .Y(new_n6563_));
  AND2X1   g05561(.A(new_n6563_), .B(\A[121] ), .Y(new_n6564_));
  OAI21X1  g05562(.A0(new_n6563_), .A1(\A[121] ), .B0(\A[123] ), .Y(new_n6565_));
  INVX1    g05563(.A(\A[123] ), .Y(new_n6566_));
  XOR2X1   g05564(.A(\A[122] ), .B(\A[121] ), .Y(new_n6567_));
  NAND2X1  g05565(.A(new_n6567_), .B(new_n6566_), .Y(new_n6568_));
  OAI21X1  g05566(.A0(new_n6565_), .A1(new_n6564_), .B0(new_n6568_), .Y(new_n6569_));
  INVX1    g05567(.A(\A[126] ), .Y(new_n6570_));
  INVX1    g05568(.A(\A[124] ), .Y(new_n6571_));
  OR2X1    g05569(.A(\A[125] ), .B(new_n6571_), .Y(new_n6572_));
  AOI21X1  g05570(.A0(\A[125] ), .A1(new_n6571_), .B0(new_n6570_), .Y(new_n6573_));
  XOR2X1   g05571(.A(\A[125] ), .B(\A[124] ), .Y(new_n6574_));
  AOI22X1  g05572(.A0(new_n6574_), .A1(new_n6570_), .B0(new_n6573_), .B1(new_n6572_), .Y(new_n6575_));
  AND2X1   g05573(.A(\A[125] ), .B(\A[124] ), .Y(new_n6576_));
  AOI21X1  g05574(.A0(new_n6574_), .A1(\A[126] ), .B0(new_n6576_), .Y(new_n6577_));
  AND2X1   g05575(.A(\A[122] ), .B(\A[121] ), .Y(new_n6578_));
  AOI21X1  g05576(.A0(new_n6567_), .A1(\A[123] ), .B0(new_n6578_), .Y(new_n6579_));
  XOR2X1   g05577(.A(new_n6575_), .B(new_n6569_), .Y(new_n6580_));
  INVX1    g05578(.A(\A[117] ), .Y(new_n6581_));
  INVX1    g05579(.A(\A[115] ), .Y(new_n6582_));
  OR2X1    g05580(.A(\A[116] ), .B(new_n6582_), .Y(new_n6583_));
  AOI21X1  g05581(.A0(\A[116] ), .A1(new_n6582_), .B0(new_n6581_), .Y(new_n6584_));
  XOR2X1   g05582(.A(\A[116] ), .B(\A[115] ), .Y(new_n6585_));
  AOI22X1  g05583(.A0(new_n6585_), .A1(new_n6581_), .B0(new_n6584_), .B1(new_n6583_), .Y(new_n6586_));
  INVX1    g05584(.A(\A[120] ), .Y(new_n6587_));
  INVX1    g05585(.A(\A[118] ), .Y(new_n6588_));
  OR2X1    g05586(.A(\A[119] ), .B(new_n6588_), .Y(new_n6589_));
  AOI21X1  g05587(.A0(\A[119] ), .A1(new_n6588_), .B0(new_n6587_), .Y(new_n6590_));
  XOR2X1   g05588(.A(\A[119] ), .B(\A[118] ), .Y(new_n6591_));
  AOI22X1  g05589(.A0(new_n6591_), .A1(new_n6587_), .B0(new_n6590_), .B1(new_n6589_), .Y(new_n6592_));
  AND2X1   g05590(.A(\A[119] ), .B(\A[118] ), .Y(new_n6593_));
  AOI21X1  g05591(.A0(new_n6591_), .A1(\A[120] ), .B0(new_n6593_), .Y(new_n6594_));
  AND2X1   g05592(.A(\A[116] ), .B(\A[115] ), .Y(new_n6595_));
  AOI21X1  g05593(.A0(new_n6585_), .A1(\A[117] ), .B0(new_n6595_), .Y(new_n6596_));
  XOR2X1   g05594(.A(new_n6592_), .B(new_n6586_), .Y(new_n6597_));
  XOR2X1   g05595(.A(new_n6597_), .B(new_n6580_), .Y(new_n6598_));
  INVX1    g05596(.A(\A[110] ), .Y(new_n6599_));
  AND2X1   g05597(.A(new_n6599_), .B(\A[109] ), .Y(new_n6600_));
  OAI21X1  g05598(.A0(new_n6599_), .A1(\A[109] ), .B0(\A[111] ), .Y(new_n6601_));
  INVX1    g05599(.A(\A[111] ), .Y(new_n6602_));
  XOR2X1   g05600(.A(\A[110] ), .B(\A[109] ), .Y(new_n6603_));
  NAND2X1  g05601(.A(new_n6603_), .B(new_n6602_), .Y(new_n6604_));
  OAI21X1  g05602(.A0(new_n6601_), .A1(new_n6600_), .B0(new_n6604_), .Y(new_n6605_));
  INVX1    g05603(.A(\A[114] ), .Y(new_n6606_));
  INVX1    g05604(.A(\A[112] ), .Y(new_n6607_));
  OR2X1    g05605(.A(\A[113] ), .B(new_n6607_), .Y(new_n6608_));
  AOI21X1  g05606(.A0(\A[113] ), .A1(new_n6607_), .B0(new_n6606_), .Y(new_n6609_));
  XOR2X1   g05607(.A(\A[113] ), .B(\A[112] ), .Y(new_n6610_));
  AOI22X1  g05608(.A0(new_n6610_), .A1(new_n6606_), .B0(new_n6609_), .B1(new_n6608_), .Y(new_n6611_));
  AND2X1   g05609(.A(\A[113] ), .B(\A[112] ), .Y(new_n6612_));
  AOI21X1  g05610(.A0(new_n6610_), .A1(\A[114] ), .B0(new_n6612_), .Y(new_n6613_));
  AND2X1   g05611(.A(\A[110] ), .B(\A[109] ), .Y(new_n6614_));
  AOI21X1  g05612(.A0(new_n6603_), .A1(\A[111] ), .B0(new_n6614_), .Y(new_n6615_));
  XOR2X1   g05613(.A(new_n6611_), .B(new_n6605_), .Y(new_n6616_));
  INVX1    g05614(.A(\A[105] ), .Y(new_n6617_));
  INVX1    g05615(.A(\A[103] ), .Y(new_n6618_));
  OR2X1    g05616(.A(\A[104] ), .B(new_n6618_), .Y(new_n6619_));
  AOI21X1  g05617(.A0(\A[104] ), .A1(new_n6618_), .B0(new_n6617_), .Y(new_n6620_));
  XOR2X1   g05618(.A(\A[104] ), .B(\A[103] ), .Y(new_n6621_));
  AOI22X1  g05619(.A0(new_n6621_), .A1(new_n6617_), .B0(new_n6620_), .B1(new_n6619_), .Y(new_n6622_));
  INVX1    g05620(.A(\A[108] ), .Y(new_n6623_));
  INVX1    g05621(.A(\A[106] ), .Y(new_n6624_));
  OR2X1    g05622(.A(\A[107] ), .B(new_n6624_), .Y(new_n6625_));
  AOI21X1  g05623(.A0(\A[107] ), .A1(new_n6624_), .B0(new_n6623_), .Y(new_n6626_));
  XOR2X1   g05624(.A(\A[107] ), .B(\A[106] ), .Y(new_n6627_));
  AOI22X1  g05625(.A0(new_n6627_), .A1(new_n6623_), .B0(new_n6626_), .B1(new_n6625_), .Y(new_n6628_));
  AND2X1   g05626(.A(\A[107] ), .B(\A[106] ), .Y(new_n6629_));
  AOI21X1  g05627(.A0(new_n6627_), .A1(\A[108] ), .B0(new_n6629_), .Y(new_n6630_));
  AND2X1   g05628(.A(\A[104] ), .B(\A[103] ), .Y(new_n6631_));
  AOI21X1  g05629(.A0(new_n6621_), .A1(\A[105] ), .B0(new_n6631_), .Y(new_n6632_));
  XOR2X1   g05630(.A(new_n6628_), .B(new_n6622_), .Y(new_n6633_));
  XOR2X1   g05631(.A(new_n6633_), .B(new_n6616_), .Y(new_n6634_));
  XOR2X1   g05632(.A(new_n6634_), .B(new_n6598_), .Y(new_n6635_));
  INVX1    g05633(.A(new_n6635_), .Y(new_n6636_));
  INVX1    g05634(.A(\A[98] ), .Y(new_n6637_));
  AND2X1   g05635(.A(new_n6637_), .B(\A[97] ), .Y(new_n6638_));
  OAI21X1  g05636(.A0(new_n6637_), .A1(\A[97] ), .B0(\A[99] ), .Y(new_n6639_));
  INVX1    g05637(.A(\A[99] ), .Y(new_n6640_));
  XOR2X1   g05638(.A(\A[98] ), .B(\A[97] ), .Y(new_n6641_));
  NAND2X1  g05639(.A(new_n6641_), .B(new_n6640_), .Y(new_n6642_));
  OAI21X1  g05640(.A0(new_n6639_), .A1(new_n6638_), .B0(new_n6642_), .Y(new_n6643_));
  INVX1    g05641(.A(\A[102] ), .Y(new_n6644_));
  INVX1    g05642(.A(\A[100] ), .Y(new_n6645_));
  OR2X1    g05643(.A(\A[101] ), .B(new_n6645_), .Y(new_n6646_));
  AOI21X1  g05644(.A0(\A[101] ), .A1(new_n6645_), .B0(new_n6644_), .Y(new_n6647_));
  XOR2X1   g05645(.A(\A[101] ), .B(\A[100] ), .Y(new_n6648_));
  AOI22X1  g05646(.A0(new_n6648_), .A1(new_n6644_), .B0(new_n6647_), .B1(new_n6646_), .Y(new_n6649_));
  AND2X1   g05647(.A(\A[101] ), .B(\A[100] ), .Y(new_n6650_));
  AOI21X1  g05648(.A0(new_n6648_), .A1(\A[102] ), .B0(new_n6650_), .Y(new_n6651_));
  AND2X1   g05649(.A(\A[98] ), .B(\A[97] ), .Y(new_n6652_));
  AOI21X1  g05650(.A0(new_n6641_), .A1(\A[99] ), .B0(new_n6652_), .Y(new_n6653_));
  XOR2X1   g05651(.A(new_n6649_), .B(new_n6643_), .Y(new_n6654_));
  INVX1    g05652(.A(\A[93] ), .Y(new_n6655_));
  INVX1    g05653(.A(\A[91] ), .Y(new_n6656_));
  OR2X1    g05654(.A(\A[92] ), .B(new_n6656_), .Y(new_n6657_));
  AOI21X1  g05655(.A0(\A[92] ), .A1(new_n6656_), .B0(new_n6655_), .Y(new_n6658_));
  XOR2X1   g05656(.A(\A[92] ), .B(\A[91] ), .Y(new_n6659_));
  AOI22X1  g05657(.A0(new_n6659_), .A1(new_n6655_), .B0(new_n6658_), .B1(new_n6657_), .Y(new_n6660_));
  INVX1    g05658(.A(\A[96] ), .Y(new_n6661_));
  INVX1    g05659(.A(\A[94] ), .Y(new_n6662_));
  OR2X1    g05660(.A(\A[95] ), .B(new_n6662_), .Y(new_n6663_));
  AOI21X1  g05661(.A0(\A[95] ), .A1(new_n6662_), .B0(new_n6661_), .Y(new_n6664_));
  XOR2X1   g05662(.A(\A[95] ), .B(\A[94] ), .Y(new_n6665_));
  AOI22X1  g05663(.A0(new_n6665_), .A1(new_n6661_), .B0(new_n6664_), .B1(new_n6663_), .Y(new_n6666_));
  AND2X1   g05664(.A(\A[95] ), .B(\A[94] ), .Y(new_n6667_));
  AOI21X1  g05665(.A0(new_n6665_), .A1(\A[96] ), .B0(new_n6667_), .Y(new_n6668_));
  AND2X1   g05666(.A(\A[92] ), .B(\A[91] ), .Y(new_n6669_));
  AOI21X1  g05667(.A0(new_n6659_), .A1(\A[93] ), .B0(new_n6669_), .Y(new_n6670_));
  XOR2X1   g05668(.A(new_n6666_), .B(new_n6660_), .Y(new_n6671_));
  XOR2X1   g05669(.A(new_n6671_), .B(new_n6654_), .Y(new_n6672_));
  INVX1    g05670(.A(new_n6672_), .Y(new_n6673_));
  INVX1    g05671(.A(\A[86] ), .Y(new_n6674_));
  AND2X1   g05672(.A(new_n6674_), .B(\A[85] ), .Y(new_n6675_));
  OAI21X1  g05673(.A0(new_n6674_), .A1(\A[85] ), .B0(\A[87] ), .Y(new_n6676_));
  INVX1    g05674(.A(\A[87] ), .Y(new_n6677_));
  XOR2X1   g05675(.A(\A[86] ), .B(\A[85] ), .Y(new_n6678_));
  NAND2X1  g05676(.A(new_n6678_), .B(new_n6677_), .Y(new_n6679_));
  OAI21X1  g05677(.A0(new_n6676_), .A1(new_n6675_), .B0(new_n6679_), .Y(new_n6680_));
  INVX1    g05678(.A(\A[90] ), .Y(new_n6681_));
  INVX1    g05679(.A(\A[88] ), .Y(new_n6682_));
  OR2X1    g05680(.A(\A[89] ), .B(new_n6682_), .Y(new_n6683_));
  AOI21X1  g05681(.A0(\A[89] ), .A1(new_n6682_), .B0(new_n6681_), .Y(new_n6684_));
  XOR2X1   g05682(.A(\A[89] ), .B(\A[88] ), .Y(new_n6685_));
  AOI22X1  g05683(.A0(new_n6685_), .A1(new_n6681_), .B0(new_n6684_), .B1(new_n6683_), .Y(new_n6686_));
  AND2X1   g05684(.A(\A[89] ), .B(\A[88] ), .Y(new_n6687_));
  AOI21X1  g05685(.A0(new_n6685_), .A1(\A[90] ), .B0(new_n6687_), .Y(new_n6688_));
  AND2X1   g05686(.A(\A[86] ), .B(\A[85] ), .Y(new_n6689_));
  AOI21X1  g05687(.A0(new_n6678_), .A1(\A[87] ), .B0(new_n6689_), .Y(new_n6690_));
  XOR2X1   g05688(.A(new_n6686_), .B(new_n6680_), .Y(new_n6691_));
  INVX1    g05689(.A(\A[81] ), .Y(new_n6692_));
  INVX1    g05690(.A(\A[79] ), .Y(new_n6693_));
  OR2X1    g05691(.A(\A[80] ), .B(new_n6693_), .Y(new_n6694_));
  AOI21X1  g05692(.A0(\A[80] ), .A1(new_n6693_), .B0(new_n6692_), .Y(new_n6695_));
  XOR2X1   g05693(.A(\A[80] ), .B(\A[79] ), .Y(new_n6696_));
  AOI22X1  g05694(.A0(new_n6696_), .A1(new_n6692_), .B0(new_n6695_), .B1(new_n6694_), .Y(new_n6697_));
  INVX1    g05695(.A(\A[84] ), .Y(new_n6698_));
  INVX1    g05696(.A(\A[82] ), .Y(new_n6699_));
  OR2X1    g05697(.A(\A[83] ), .B(new_n6699_), .Y(new_n6700_));
  AOI21X1  g05698(.A0(\A[83] ), .A1(new_n6699_), .B0(new_n6698_), .Y(new_n6701_));
  XOR2X1   g05699(.A(\A[83] ), .B(\A[82] ), .Y(new_n6702_));
  AOI22X1  g05700(.A0(new_n6702_), .A1(new_n6698_), .B0(new_n6701_), .B1(new_n6700_), .Y(new_n6703_));
  AND2X1   g05701(.A(\A[83] ), .B(\A[82] ), .Y(new_n6704_));
  AOI21X1  g05702(.A0(new_n6702_), .A1(\A[84] ), .B0(new_n6704_), .Y(new_n6705_));
  AND2X1   g05703(.A(\A[80] ), .B(\A[79] ), .Y(new_n6706_));
  AOI21X1  g05704(.A0(new_n6696_), .A1(\A[81] ), .B0(new_n6706_), .Y(new_n6707_));
  XOR2X1   g05705(.A(new_n6703_), .B(new_n6697_), .Y(new_n6708_));
  XOR2X1   g05706(.A(new_n6708_), .B(new_n6691_), .Y(new_n6709_));
  XOR2X1   g05707(.A(new_n6709_), .B(new_n6673_), .Y(new_n6710_));
  XOR2X1   g05708(.A(new_n6710_), .B(new_n6636_), .Y(new_n6711_));
  XOR2X1   g05709(.A(new_n6711_), .B(new_n6562_), .Y(new_n6712_));
  NOR2X1   g05710(.A(new_n6712_), .B(new_n6414_), .Y(new_n6713_));
  INVX1    g05711(.A(new_n6713_), .Y(new_n6714_));
  AND2X1   g05712(.A(new_n6410_), .B(new_n6407_), .Y(new_n6715_));
  AOI21X1  g05713(.A0(new_n6364_), .A1(new_n6256_), .B0(new_n6408_), .Y(new_n6716_));
  AOI22X1  g05714(.A0(new_n6716_), .A1(new_n6350_), .B0(new_n6369_), .B1(new_n6408_), .Y(new_n6717_));
  MX2X1    g05715(.A(new_n6717_), .B(new_n6370_), .S0(new_n6407_), .Y(new_n6718_));
  OAI21X1  g05716(.A0(new_n6717_), .A1(new_n6407_), .B0(new_n6376_), .Y(new_n6719_));
  OAI22X1  g05717(.A0(new_n6719_), .A1(new_n6715_), .B0(new_n6718_), .B1(new_n6376_), .Y(new_n6720_));
  AOI21X1  g05718(.A0(new_n6720_), .A1(new_n6013_), .B0(new_n6714_), .Y(new_n6721_));
  OR2X1    g05719(.A(new_n5909_), .B(new_n5906_), .Y(new_n6722_));
  OAI21X1  g05720(.A0(new_n5802_), .A1(new_n5751_), .B0(new_n5907_), .Y(new_n6723_));
  OAI22X1  g05721(.A0(new_n6723_), .A1(new_n5784_), .B0(new_n5806_), .B1(new_n5907_), .Y(new_n6724_));
  AOI21X1  g05722(.A0(new_n6724_), .A1(new_n5906_), .B0(new_n6010_), .Y(new_n6725_));
  MX2X1    g05723(.A(new_n5807_), .B(new_n6724_), .S0(new_n5906_), .Y(new_n6726_));
  AOI22X1  g05724(.A0(new_n6726_), .A1(new_n6010_), .B0(new_n6725_), .B1(new_n6722_), .Y(new_n6727_));
  AOI21X1  g05725(.A0(new_n6724_), .A1(new_n5906_), .B0(new_n5886_), .Y(new_n6728_));
  AOI22X1  g05726(.A0(new_n6728_), .A1(new_n6722_), .B0(new_n6726_), .B1(new_n5886_), .Y(new_n6729_));
  MX2X1    g05727(.A(new_n6729_), .B(new_n6727_), .S0(new_n6009_), .Y(new_n6730_));
  NOR2X1   g05728(.A(new_n6375_), .B(new_n6373_), .Y(new_n6731_));
  OAI21X1  g05729(.A0(new_n6717_), .A1(new_n6407_), .B0(new_n6731_), .Y(new_n6732_));
  OAI22X1  g05730(.A0(new_n6718_), .A1(new_n6731_), .B0(new_n6732_), .B1(new_n6715_), .Y(new_n6733_));
  MX2X1    g05731(.A(new_n6720_), .B(new_n6733_), .S0(new_n6730_), .Y(new_n6734_));
  AOI22X1  g05732(.A0(new_n6734_), .A1(new_n6714_), .B0(new_n6721_), .B1(new_n6413_), .Y(new_n6735_));
  INVX1    g05733(.A(\A[140] ), .Y(new_n6736_));
  AND2X1   g05734(.A(new_n6736_), .B(\A[139] ), .Y(new_n6737_));
  OAI21X1  g05735(.A0(new_n6736_), .A1(\A[139] ), .B0(\A[141] ), .Y(new_n6738_));
  NAND2X1  g05736(.A(new_n6510_), .B(new_n6506_), .Y(new_n6739_));
  OAI21X1  g05737(.A0(new_n6738_), .A1(new_n6737_), .B0(new_n6739_), .Y(new_n6740_));
  XOR2X1   g05738(.A(new_n6517_), .B(new_n6740_), .Y(new_n6741_));
  XOR2X1   g05739(.A(new_n6521_), .B(new_n6519_), .Y(new_n6742_));
  NOR2X1   g05740(.A(new_n6517_), .B(new_n6511_), .Y(new_n6743_));
  NOR2X1   g05741(.A(new_n6521_), .B(new_n6519_), .Y(new_n6744_));
  AOI21X1  g05742(.A0(new_n6743_), .A1(new_n6742_), .B0(new_n6744_), .Y(new_n6745_));
  XOR2X1   g05743(.A(new_n6743_), .B(new_n6742_), .Y(new_n6746_));
  OAI21X1  g05744(.A0(new_n6745_), .A1(new_n6741_), .B0(new_n6746_), .Y(new_n6747_));
  XOR2X1   g05745(.A(new_n6500_), .B(new_n6494_), .Y(new_n6748_));
  INVX1    g05746(.A(\A[145] ), .Y(new_n6749_));
  OR2X1    g05747(.A(\A[146] ), .B(new_n6749_), .Y(new_n6750_));
  AOI21X1  g05748(.A0(\A[146] ), .A1(new_n6749_), .B0(new_n6491_), .Y(new_n6751_));
  AOI22X1  g05749(.A0(new_n6492_), .A1(new_n6491_), .B0(new_n6751_), .B1(new_n6750_), .Y(new_n6752_));
  NOR4X1   g05750(.A(new_n6504_), .B(new_n6502_), .C(new_n6500_), .D(new_n6752_), .Y(new_n6753_));
  NOR4X1   g05751(.A(new_n6521_), .B(new_n6519_), .C(new_n6517_), .D(new_n6511_), .Y(new_n6754_));
  OR4X1    g05752(.A(new_n6754_), .B(new_n6741_), .C(new_n6753_), .D(new_n6748_), .Y(new_n6755_));
  XOR2X1   g05753(.A(new_n6504_), .B(new_n6502_), .Y(new_n6756_));
  NOR2X1   g05754(.A(new_n6500_), .B(new_n6752_), .Y(new_n6757_));
  NOR2X1   g05755(.A(new_n6504_), .B(new_n6502_), .Y(new_n6758_));
  AOI21X1  g05756(.A0(new_n6757_), .A1(new_n6756_), .B0(new_n6758_), .Y(new_n6759_));
  XOR2X1   g05757(.A(new_n6757_), .B(new_n6756_), .Y(new_n6760_));
  OAI21X1  g05758(.A0(new_n6759_), .A1(new_n6748_), .B0(new_n6760_), .Y(new_n6761_));
  XOR2X1   g05759(.A(new_n6761_), .B(new_n6755_), .Y(new_n6762_));
  AND2X1   g05760(.A(new_n6762_), .B(new_n6747_), .Y(new_n6763_));
  NOR2X1   g05761(.A(new_n6560_), .B(new_n6523_), .Y(new_n6764_));
  AND2X1   g05762(.A(new_n6499_), .B(\A[150] ), .Y(new_n6765_));
  OR2X1    g05763(.A(new_n6765_), .B(new_n6501_), .Y(new_n6766_));
  XOR2X1   g05764(.A(new_n6504_), .B(new_n6766_), .Y(new_n6767_));
  OR2X1    g05765(.A(new_n6500_), .B(new_n6752_), .Y(new_n6768_));
  OR2X1    g05766(.A(new_n6504_), .B(new_n6502_), .Y(new_n6769_));
  OAI21X1  g05767(.A0(new_n6768_), .A1(new_n6767_), .B0(new_n6769_), .Y(new_n6770_));
  XOR2X1   g05768(.A(new_n6768_), .B(new_n6756_), .Y(new_n6771_));
  NOR4X1   g05769(.A(new_n6741_), .B(new_n6771_), .C(new_n6770_), .D(new_n6748_), .Y(new_n6772_));
  XOR2X1   g05770(.A(new_n6500_), .B(new_n6752_), .Y(new_n6773_));
  AOI21X1  g05771(.A0(new_n6770_), .A1(new_n6773_), .B0(new_n6754_), .Y(new_n6774_));
  AOI22X1  g05772(.A0(new_n6774_), .A1(new_n6772_), .B0(new_n6761_), .B1(new_n6755_), .Y(new_n6775_));
  OAI21X1  g05773(.A0(new_n6775_), .A1(new_n6747_), .B0(new_n6764_), .Y(new_n6776_));
  AOI21X1  g05774(.A0(new_n6770_), .A1(new_n6773_), .B0(new_n6771_), .Y(new_n6777_));
  XOR2X1   g05775(.A(new_n6777_), .B(new_n6755_), .Y(new_n6778_));
  MX2X1    g05776(.A(new_n6775_), .B(new_n6778_), .S0(new_n6747_), .Y(new_n6779_));
  OAI22X1  g05777(.A0(new_n6779_), .A1(new_n6764_), .B0(new_n6776_), .B1(new_n6763_), .Y(new_n6780_));
  INVX1    g05778(.A(\A[128] ), .Y(new_n6781_));
  AND2X1   g05779(.A(new_n6781_), .B(\A[127] ), .Y(new_n6782_));
  OAI21X1  g05780(.A0(new_n6781_), .A1(\A[127] ), .B0(\A[129] ), .Y(new_n6783_));
  NAND2X1  g05781(.A(new_n6547_), .B(new_n6543_), .Y(new_n6784_));
  OAI21X1  g05782(.A0(new_n6783_), .A1(new_n6782_), .B0(new_n6784_), .Y(new_n6785_));
  XOR2X1   g05783(.A(new_n6554_), .B(new_n6785_), .Y(new_n6786_));
  XOR2X1   g05784(.A(new_n6558_), .B(new_n6556_), .Y(new_n6787_));
  NOR2X1   g05785(.A(new_n6554_), .B(new_n6548_), .Y(new_n6788_));
  NOR2X1   g05786(.A(new_n6558_), .B(new_n6556_), .Y(new_n6789_));
  AOI21X1  g05787(.A0(new_n6788_), .A1(new_n6787_), .B0(new_n6789_), .Y(new_n6790_));
  XOR2X1   g05788(.A(new_n6788_), .B(new_n6787_), .Y(new_n6791_));
  OAI21X1  g05789(.A0(new_n6790_), .A1(new_n6786_), .B0(new_n6791_), .Y(new_n6792_));
  XOR2X1   g05790(.A(new_n6537_), .B(new_n6531_), .Y(new_n6793_));
  INVX1    g05791(.A(\A[133] ), .Y(new_n6794_));
  OR2X1    g05792(.A(\A[134] ), .B(new_n6794_), .Y(new_n6795_));
  AOI21X1  g05793(.A0(\A[134] ), .A1(new_n6794_), .B0(new_n6528_), .Y(new_n6796_));
  AOI22X1  g05794(.A0(new_n6529_), .A1(new_n6528_), .B0(new_n6796_), .B1(new_n6795_), .Y(new_n6797_));
  NOR4X1   g05795(.A(new_n6541_), .B(new_n6539_), .C(new_n6537_), .D(new_n6797_), .Y(new_n6798_));
  NOR4X1   g05796(.A(new_n6558_), .B(new_n6556_), .C(new_n6554_), .D(new_n6548_), .Y(new_n6799_));
  OR4X1    g05797(.A(new_n6799_), .B(new_n6786_), .C(new_n6798_), .D(new_n6793_), .Y(new_n6800_));
  XOR2X1   g05798(.A(new_n6537_), .B(new_n6797_), .Y(new_n6801_));
  AND2X1   g05799(.A(new_n6536_), .B(\A[138] ), .Y(new_n6802_));
  OR2X1    g05800(.A(new_n6802_), .B(new_n6538_), .Y(new_n6803_));
  XOR2X1   g05801(.A(new_n6541_), .B(new_n6803_), .Y(new_n6804_));
  OR2X1    g05802(.A(new_n6537_), .B(new_n6797_), .Y(new_n6805_));
  OR2X1    g05803(.A(new_n6541_), .B(new_n6539_), .Y(new_n6806_));
  OAI21X1  g05804(.A0(new_n6805_), .A1(new_n6804_), .B0(new_n6806_), .Y(new_n6807_));
  NOR2X1   g05805(.A(new_n6537_), .B(new_n6797_), .Y(new_n6808_));
  XOR2X1   g05806(.A(new_n6808_), .B(new_n6804_), .Y(new_n6809_));
  AOI21X1  g05807(.A0(new_n6807_), .A1(new_n6801_), .B0(new_n6809_), .Y(new_n6810_));
  XOR2X1   g05808(.A(new_n6810_), .B(new_n6800_), .Y(new_n6811_));
  XOR2X1   g05809(.A(new_n6541_), .B(new_n6539_), .Y(new_n6812_));
  NOR2X1   g05810(.A(new_n6541_), .B(new_n6539_), .Y(new_n6813_));
  AOI21X1  g05811(.A0(new_n6808_), .A1(new_n6812_), .B0(new_n6813_), .Y(new_n6814_));
  XOR2X1   g05812(.A(new_n6808_), .B(new_n6812_), .Y(new_n6815_));
  OAI21X1  g05813(.A0(new_n6814_), .A1(new_n6793_), .B0(new_n6815_), .Y(new_n6816_));
  NOR4X1   g05814(.A(new_n6786_), .B(new_n6809_), .C(new_n6807_), .D(new_n6793_), .Y(new_n6817_));
  AOI21X1  g05815(.A0(new_n6807_), .A1(new_n6801_), .B0(new_n6799_), .Y(new_n6818_));
  AOI22X1  g05816(.A0(new_n6818_), .A1(new_n6817_), .B0(new_n6816_), .B1(new_n6800_), .Y(new_n6819_));
  MX2X1    g05817(.A(new_n6819_), .B(new_n6811_), .S0(new_n6792_), .Y(new_n6820_));
  OR2X1    g05818(.A(new_n6560_), .B(new_n6523_), .Y(new_n6821_));
  OAI21X1  g05819(.A0(new_n6775_), .A1(new_n6747_), .B0(new_n6821_), .Y(new_n6822_));
  OAI22X1  g05820(.A0(new_n6822_), .A1(new_n6763_), .B0(new_n6779_), .B1(new_n6821_), .Y(new_n6823_));
  MX2X1    g05821(.A(new_n6823_), .B(new_n6780_), .S0(new_n6820_), .Y(new_n6824_));
  INVX1    g05822(.A(\A[152] ), .Y(new_n6825_));
  AND2X1   g05823(.A(new_n6825_), .B(\A[151] ), .Y(new_n6826_));
  OAI21X1  g05824(.A0(new_n6825_), .A1(\A[151] ), .B0(\A[153] ), .Y(new_n6827_));
  NAND2X1  g05825(.A(new_n6473_), .B(new_n6469_), .Y(new_n6828_));
  OAI21X1  g05826(.A0(new_n6827_), .A1(new_n6826_), .B0(new_n6828_), .Y(new_n6829_));
  XOR2X1   g05827(.A(new_n6480_), .B(new_n6829_), .Y(new_n6830_));
  XOR2X1   g05828(.A(new_n6484_), .B(new_n6482_), .Y(new_n6831_));
  NOR2X1   g05829(.A(new_n6480_), .B(new_n6474_), .Y(new_n6832_));
  NOR2X1   g05830(.A(new_n6484_), .B(new_n6482_), .Y(new_n6833_));
  AOI21X1  g05831(.A0(new_n6832_), .A1(new_n6831_), .B0(new_n6833_), .Y(new_n6834_));
  XOR2X1   g05832(.A(new_n6832_), .B(new_n6831_), .Y(new_n6835_));
  OAI21X1  g05833(.A0(new_n6834_), .A1(new_n6830_), .B0(new_n6835_), .Y(new_n6836_));
  XOR2X1   g05834(.A(new_n6463_), .B(new_n6457_), .Y(new_n6837_));
  INVX1    g05835(.A(\A[157] ), .Y(new_n6838_));
  OR2X1    g05836(.A(\A[158] ), .B(new_n6838_), .Y(new_n6839_));
  AOI21X1  g05837(.A0(\A[158] ), .A1(new_n6838_), .B0(new_n6454_), .Y(new_n6840_));
  AOI22X1  g05838(.A0(new_n6455_), .A1(new_n6454_), .B0(new_n6840_), .B1(new_n6839_), .Y(new_n6841_));
  NOR4X1   g05839(.A(new_n6467_), .B(new_n6465_), .C(new_n6463_), .D(new_n6841_), .Y(new_n6842_));
  NOR4X1   g05840(.A(new_n6484_), .B(new_n6482_), .C(new_n6480_), .D(new_n6474_), .Y(new_n6843_));
  NOR4X1   g05841(.A(new_n6843_), .B(new_n6830_), .C(new_n6842_), .D(new_n6837_), .Y(new_n6844_));
  XOR2X1   g05842(.A(new_n6463_), .B(new_n6841_), .Y(new_n6845_));
  AND2X1   g05843(.A(new_n6462_), .B(\A[162] ), .Y(new_n6846_));
  OR2X1    g05844(.A(new_n6846_), .B(new_n6464_), .Y(new_n6847_));
  XOR2X1   g05845(.A(new_n6467_), .B(new_n6847_), .Y(new_n6848_));
  OR2X1    g05846(.A(new_n6463_), .B(new_n6841_), .Y(new_n6849_));
  OR2X1    g05847(.A(new_n6467_), .B(new_n6465_), .Y(new_n6850_));
  OAI21X1  g05848(.A0(new_n6849_), .A1(new_n6848_), .B0(new_n6850_), .Y(new_n6851_));
  NOR2X1   g05849(.A(new_n6463_), .B(new_n6841_), .Y(new_n6852_));
  XOR2X1   g05850(.A(new_n6852_), .B(new_n6848_), .Y(new_n6853_));
  AOI21X1  g05851(.A0(new_n6851_), .A1(new_n6845_), .B0(new_n6853_), .Y(new_n6854_));
  XOR2X1   g05852(.A(new_n6854_), .B(new_n6844_), .Y(new_n6855_));
  OR4X1    g05853(.A(new_n6830_), .B(new_n6842_), .C(new_n6853_), .D(new_n6837_), .Y(new_n6856_));
  XOR2X1   g05854(.A(new_n6467_), .B(new_n6465_), .Y(new_n6857_));
  NOR2X1   g05855(.A(new_n6467_), .B(new_n6465_), .Y(new_n6858_));
  AOI21X1  g05856(.A0(new_n6852_), .A1(new_n6857_), .B0(new_n6858_), .Y(new_n6859_));
  AND2X1   g05857(.A(new_n6479_), .B(\A[156] ), .Y(new_n6860_));
  OR2X1    g05858(.A(new_n6860_), .B(new_n6481_), .Y(new_n6861_));
  XOR2X1   g05859(.A(new_n6484_), .B(new_n6861_), .Y(new_n6862_));
  XOR2X1   g05860(.A(new_n6832_), .B(new_n6862_), .Y(new_n6863_));
  OAI22X1  g05861(.A0(new_n6863_), .A1(new_n6834_), .B0(new_n6859_), .B1(new_n6837_), .Y(new_n6864_));
  OAI22X1  g05862(.A0(new_n6864_), .A1(new_n6856_), .B0(new_n6854_), .B1(new_n6844_), .Y(new_n6865_));
  MX2X1    g05863(.A(new_n6865_), .B(new_n6855_), .S0(new_n6836_), .Y(new_n6866_));
  INVX1    g05864(.A(\A[164] ), .Y(new_n6867_));
  AND2X1   g05865(.A(new_n6867_), .B(\A[163] ), .Y(new_n6868_));
  OAI21X1  g05866(.A0(new_n6867_), .A1(\A[163] ), .B0(\A[165] ), .Y(new_n6869_));
  NAND2X1  g05867(.A(new_n6437_), .B(new_n6433_), .Y(new_n6870_));
  OAI21X1  g05868(.A0(new_n6869_), .A1(new_n6868_), .B0(new_n6870_), .Y(new_n6871_));
  XOR2X1   g05869(.A(new_n6444_), .B(new_n6871_), .Y(new_n6872_));
  XOR2X1   g05870(.A(new_n6448_), .B(new_n6446_), .Y(new_n6873_));
  NOR2X1   g05871(.A(new_n6444_), .B(new_n6438_), .Y(new_n6874_));
  NOR2X1   g05872(.A(new_n6448_), .B(new_n6446_), .Y(new_n6875_));
  AOI21X1  g05873(.A0(new_n6874_), .A1(new_n6873_), .B0(new_n6875_), .Y(new_n6876_));
  XOR2X1   g05874(.A(new_n6874_), .B(new_n6873_), .Y(new_n6877_));
  OAI21X1  g05875(.A0(new_n6876_), .A1(new_n6872_), .B0(new_n6877_), .Y(new_n6878_));
  XOR2X1   g05876(.A(new_n6427_), .B(new_n6421_), .Y(new_n6879_));
  INVX1    g05877(.A(\A[169] ), .Y(new_n6880_));
  OR2X1    g05878(.A(\A[170] ), .B(new_n6880_), .Y(new_n6881_));
  AOI21X1  g05879(.A0(\A[170] ), .A1(new_n6880_), .B0(new_n6418_), .Y(new_n6882_));
  AOI22X1  g05880(.A0(new_n6419_), .A1(new_n6418_), .B0(new_n6882_), .B1(new_n6881_), .Y(new_n6883_));
  NOR4X1   g05881(.A(new_n6431_), .B(new_n6429_), .C(new_n6427_), .D(new_n6883_), .Y(new_n6884_));
  NOR4X1   g05882(.A(new_n6448_), .B(new_n6446_), .C(new_n6444_), .D(new_n6438_), .Y(new_n6885_));
  OR4X1    g05883(.A(new_n6885_), .B(new_n6872_), .C(new_n6884_), .D(new_n6879_), .Y(new_n6886_));
  XOR2X1   g05884(.A(new_n6431_), .B(new_n6429_), .Y(new_n6887_));
  NOR2X1   g05885(.A(new_n6427_), .B(new_n6883_), .Y(new_n6888_));
  NOR2X1   g05886(.A(new_n6431_), .B(new_n6429_), .Y(new_n6889_));
  AOI21X1  g05887(.A0(new_n6888_), .A1(new_n6887_), .B0(new_n6889_), .Y(new_n6890_));
  XOR2X1   g05888(.A(new_n6888_), .B(new_n6887_), .Y(new_n6891_));
  OAI21X1  g05889(.A0(new_n6890_), .A1(new_n6879_), .B0(new_n6891_), .Y(new_n6892_));
  XOR2X1   g05890(.A(new_n6892_), .B(new_n6886_), .Y(new_n6893_));
  NAND2X1  g05891(.A(new_n6893_), .B(new_n6878_), .Y(new_n6894_));
  OR2X1    g05892(.A(new_n6486_), .B(new_n6450_), .Y(new_n6895_));
  XOR2X1   g05893(.A(new_n6444_), .B(new_n6438_), .Y(new_n6896_));
  AND2X1   g05894(.A(new_n6443_), .B(\A[168] ), .Y(new_n6897_));
  OR2X1    g05895(.A(new_n6897_), .B(new_n6445_), .Y(new_n6898_));
  XOR2X1   g05896(.A(new_n6448_), .B(new_n6898_), .Y(new_n6899_));
  OR2X1    g05897(.A(new_n6444_), .B(new_n6438_), .Y(new_n6900_));
  OR2X1    g05898(.A(new_n6448_), .B(new_n6446_), .Y(new_n6901_));
  OAI21X1  g05899(.A0(new_n6900_), .A1(new_n6899_), .B0(new_n6901_), .Y(new_n6902_));
  XOR2X1   g05900(.A(new_n6874_), .B(new_n6899_), .Y(new_n6903_));
  AOI21X1  g05901(.A0(new_n6902_), .A1(new_n6896_), .B0(new_n6903_), .Y(new_n6904_));
  NOR4X1   g05902(.A(new_n6885_), .B(new_n6872_), .C(new_n6884_), .D(new_n6879_), .Y(new_n6905_));
  XOR2X1   g05903(.A(new_n6427_), .B(new_n6883_), .Y(new_n6906_));
  AND2X1   g05904(.A(new_n6426_), .B(\A[174] ), .Y(new_n6907_));
  OR2X1    g05905(.A(new_n6907_), .B(new_n6428_), .Y(new_n6908_));
  XOR2X1   g05906(.A(new_n6431_), .B(new_n6908_), .Y(new_n6909_));
  OR2X1    g05907(.A(new_n6427_), .B(new_n6883_), .Y(new_n6910_));
  OR2X1    g05908(.A(new_n6431_), .B(new_n6429_), .Y(new_n6911_));
  OAI21X1  g05909(.A0(new_n6910_), .A1(new_n6909_), .B0(new_n6911_), .Y(new_n6912_));
  XOR2X1   g05910(.A(new_n6910_), .B(new_n6887_), .Y(new_n6913_));
  AOI21X1  g05911(.A0(new_n6912_), .A1(new_n6906_), .B0(new_n6913_), .Y(new_n6914_));
  OR4X1    g05912(.A(new_n6872_), .B(new_n6884_), .C(new_n6913_), .D(new_n6879_), .Y(new_n6915_));
  OAI22X1  g05913(.A0(new_n6903_), .A1(new_n6876_), .B0(new_n6890_), .B1(new_n6879_), .Y(new_n6916_));
  OAI22X1  g05914(.A0(new_n6916_), .A1(new_n6915_), .B0(new_n6914_), .B1(new_n6905_), .Y(new_n6917_));
  AOI21X1  g05915(.A0(new_n6917_), .A1(new_n6904_), .B0(new_n6895_), .Y(new_n6918_));
  MX2X1    g05916(.A(new_n6917_), .B(new_n6893_), .S0(new_n6878_), .Y(new_n6919_));
  AOI22X1  g05917(.A0(new_n6919_), .A1(new_n6895_), .B0(new_n6918_), .B1(new_n6894_), .Y(new_n6920_));
  OR2X1    g05918(.A(new_n6920_), .B(new_n6866_), .Y(new_n6921_));
  INVX1    g05919(.A(new_n6487_), .Y(new_n6922_));
  OR2X1    g05920(.A(new_n6561_), .B(new_n6922_), .Y(new_n6923_));
  AND2X1   g05921(.A(new_n6893_), .B(new_n6878_), .Y(new_n6924_));
  XOR2X1   g05922(.A(new_n6914_), .B(new_n6886_), .Y(new_n6925_));
  NOR4X1   g05923(.A(new_n6872_), .B(new_n6913_), .C(new_n6912_), .D(new_n6879_), .Y(new_n6926_));
  AOI21X1  g05924(.A0(new_n6912_), .A1(new_n6906_), .B0(new_n6885_), .Y(new_n6927_));
  AOI22X1  g05925(.A0(new_n6927_), .A1(new_n6926_), .B0(new_n6892_), .B1(new_n6886_), .Y(new_n6928_));
  MX2X1    g05926(.A(new_n6928_), .B(new_n6925_), .S0(new_n6878_), .Y(new_n6929_));
  OAI21X1  g05927(.A0(new_n6928_), .A1(new_n6878_), .B0(new_n6895_), .Y(new_n6930_));
  OAI22X1  g05928(.A0(new_n6930_), .A1(new_n6924_), .B0(new_n6929_), .B1(new_n6895_), .Y(new_n6931_));
  AOI21X1  g05929(.A0(new_n6931_), .A1(new_n6866_), .B0(new_n6923_), .Y(new_n6932_));
  OR4X1    g05930(.A(new_n6843_), .B(new_n6830_), .C(new_n6842_), .D(new_n6837_), .Y(new_n6933_));
  XOR2X1   g05931(.A(new_n6854_), .B(new_n6933_), .Y(new_n6934_));
  XOR2X1   g05932(.A(new_n6852_), .B(new_n6857_), .Y(new_n6935_));
  OAI21X1  g05933(.A0(new_n6859_), .A1(new_n6837_), .B0(new_n6935_), .Y(new_n6936_));
  NOR4X1   g05934(.A(new_n6830_), .B(new_n6853_), .C(new_n6851_), .D(new_n6837_), .Y(new_n6937_));
  AOI21X1  g05935(.A0(new_n6851_), .A1(new_n6845_), .B0(new_n6843_), .Y(new_n6938_));
  AOI22X1  g05936(.A0(new_n6938_), .A1(new_n6937_), .B0(new_n6936_), .B1(new_n6933_), .Y(new_n6939_));
  MX2X1    g05937(.A(new_n6939_), .B(new_n6934_), .S0(new_n6836_), .Y(new_n6940_));
  NOR2X1   g05938(.A(new_n6486_), .B(new_n6450_), .Y(new_n6941_));
  OAI21X1  g05939(.A0(new_n6928_), .A1(new_n6878_), .B0(new_n6941_), .Y(new_n6942_));
  OAI22X1  g05940(.A0(new_n6929_), .A1(new_n6941_), .B0(new_n6942_), .B1(new_n6924_), .Y(new_n6943_));
  MX2X1    g05941(.A(new_n6931_), .B(new_n6943_), .S0(new_n6940_), .Y(new_n6944_));
  AOI22X1  g05942(.A0(new_n6944_), .A1(new_n6923_), .B0(new_n6932_), .B1(new_n6921_), .Y(new_n6945_));
  OR2X1    g05943(.A(new_n6945_), .B(new_n6824_), .Y(new_n6946_));
  XOR2X1   g05944(.A(new_n6710_), .B(new_n6635_), .Y(new_n6947_));
  NOR2X1   g05945(.A(new_n6947_), .B(new_n6562_), .Y(new_n6948_));
  INVX1    g05946(.A(new_n6948_), .Y(new_n6949_));
  AND2X1   g05947(.A(new_n6943_), .B(new_n6940_), .Y(new_n6950_));
  AOI21X1  g05948(.A0(new_n6917_), .A1(new_n6904_), .B0(new_n6941_), .Y(new_n6951_));
  AOI22X1  g05949(.A0(new_n6951_), .A1(new_n6894_), .B0(new_n6919_), .B1(new_n6941_), .Y(new_n6952_));
  MX2X1    g05950(.A(new_n6952_), .B(new_n6920_), .S0(new_n6940_), .Y(new_n6953_));
  OAI21X1  g05951(.A0(new_n6952_), .A1(new_n6940_), .B0(new_n6923_), .Y(new_n6954_));
  OAI22X1  g05952(.A0(new_n6954_), .A1(new_n6950_), .B0(new_n6953_), .B1(new_n6923_), .Y(new_n6955_));
  AOI21X1  g05953(.A0(new_n6955_), .A1(new_n6824_), .B0(new_n6949_), .Y(new_n6956_));
  NAND2X1  g05954(.A(new_n6762_), .B(new_n6747_), .Y(new_n6957_));
  XOR2X1   g05955(.A(new_n6517_), .B(new_n6511_), .Y(new_n6958_));
  AND2X1   g05956(.A(new_n6516_), .B(\A[144] ), .Y(new_n6959_));
  OR2X1    g05957(.A(new_n6959_), .B(new_n6518_), .Y(new_n6960_));
  XOR2X1   g05958(.A(new_n6521_), .B(new_n6960_), .Y(new_n6961_));
  OR2X1    g05959(.A(new_n6517_), .B(new_n6511_), .Y(new_n6962_));
  OR2X1    g05960(.A(new_n6521_), .B(new_n6519_), .Y(new_n6963_));
  OAI21X1  g05961(.A0(new_n6962_), .A1(new_n6961_), .B0(new_n6963_), .Y(new_n6964_));
  XOR2X1   g05962(.A(new_n6743_), .B(new_n6961_), .Y(new_n6965_));
  AOI21X1  g05963(.A0(new_n6964_), .A1(new_n6958_), .B0(new_n6965_), .Y(new_n6966_));
  NOR4X1   g05964(.A(new_n6754_), .B(new_n6741_), .C(new_n6753_), .D(new_n6748_), .Y(new_n6967_));
  OR4X1    g05965(.A(new_n6741_), .B(new_n6753_), .C(new_n6771_), .D(new_n6748_), .Y(new_n6968_));
  OAI22X1  g05966(.A0(new_n6965_), .A1(new_n6745_), .B0(new_n6759_), .B1(new_n6748_), .Y(new_n6969_));
  OAI22X1  g05967(.A0(new_n6969_), .A1(new_n6968_), .B0(new_n6777_), .B1(new_n6967_), .Y(new_n6970_));
  AOI21X1  g05968(.A0(new_n6970_), .A1(new_n6966_), .B0(new_n6821_), .Y(new_n6971_));
  MX2X1    g05969(.A(new_n6970_), .B(new_n6762_), .S0(new_n6747_), .Y(new_n6972_));
  AOI22X1  g05970(.A0(new_n6972_), .A1(new_n6821_), .B0(new_n6971_), .B1(new_n6957_), .Y(new_n6973_));
  AOI21X1  g05971(.A0(new_n6970_), .A1(new_n6966_), .B0(new_n6764_), .Y(new_n6974_));
  AOI22X1  g05972(.A0(new_n6974_), .A1(new_n6957_), .B0(new_n6972_), .B1(new_n6764_), .Y(new_n6975_));
  MX2X1    g05973(.A(new_n6975_), .B(new_n6973_), .S0(new_n6820_), .Y(new_n6976_));
  NOR2X1   g05974(.A(new_n6561_), .B(new_n6922_), .Y(new_n6977_));
  OAI21X1  g05975(.A0(new_n6952_), .A1(new_n6940_), .B0(new_n6977_), .Y(new_n6978_));
  OAI22X1  g05976(.A0(new_n6953_), .A1(new_n6977_), .B0(new_n6978_), .B1(new_n6950_), .Y(new_n6979_));
  MX2X1    g05977(.A(new_n6955_), .B(new_n6979_), .S0(new_n6976_), .Y(new_n6980_));
  AOI22X1  g05978(.A0(new_n6980_), .A1(new_n6949_), .B0(new_n6956_), .B1(new_n6946_), .Y(new_n6981_));
  INVX1    g05979(.A(\A[104] ), .Y(new_n6982_));
  AND2X1   g05980(.A(new_n6982_), .B(\A[103] ), .Y(new_n6983_));
  OAI21X1  g05981(.A0(new_n6982_), .A1(\A[103] ), .B0(\A[105] ), .Y(new_n6984_));
  NAND2X1  g05982(.A(new_n6621_), .B(new_n6617_), .Y(new_n6985_));
  OAI21X1  g05983(.A0(new_n6984_), .A1(new_n6983_), .B0(new_n6985_), .Y(new_n6986_));
  XOR2X1   g05984(.A(new_n6628_), .B(new_n6986_), .Y(new_n6987_));
  XOR2X1   g05985(.A(new_n6632_), .B(new_n6630_), .Y(new_n6988_));
  NOR2X1   g05986(.A(new_n6628_), .B(new_n6622_), .Y(new_n6989_));
  NOR2X1   g05987(.A(new_n6632_), .B(new_n6630_), .Y(new_n6990_));
  AOI21X1  g05988(.A0(new_n6989_), .A1(new_n6988_), .B0(new_n6990_), .Y(new_n6991_));
  XOR2X1   g05989(.A(new_n6989_), .B(new_n6988_), .Y(new_n6992_));
  OAI21X1  g05990(.A0(new_n6991_), .A1(new_n6987_), .B0(new_n6992_), .Y(new_n6993_));
  XOR2X1   g05991(.A(new_n6611_), .B(new_n6605_), .Y(new_n6994_));
  INVX1    g05992(.A(\A[109] ), .Y(new_n6995_));
  OR2X1    g05993(.A(\A[110] ), .B(new_n6995_), .Y(new_n6996_));
  AOI21X1  g05994(.A0(\A[110] ), .A1(new_n6995_), .B0(new_n6602_), .Y(new_n6997_));
  AOI22X1  g05995(.A0(new_n6603_), .A1(new_n6602_), .B0(new_n6997_), .B1(new_n6996_), .Y(new_n6998_));
  NOR4X1   g05996(.A(new_n6615_), .B(new_n6613_), .C(new_n6611_), .D(new_n6998_), .Y(new_n6999_));
  NOR4X1   g05997(.A(new_n6632_), .B(new_n6630_), .C(new_n6628_), .D(new_n6622_), .Y(new_n7000_));
  NOR4X1   g05998(.A(new_n7000_), .B(new_n6987_), .C(new_n6999_), .D(new_n6994_), .Y(new_n7001_));
  XOR2X1   g05999(.A(new_n6611_), .B(new_n6998_), .Y(new_n7002_));
  AND2X1   g06000(.A(new_n6610_), .B(\A[114] ), .Y(new_n7003_));
  OR2X1    g06001(.A(new_n7003_), .B(new_n6612_), .Y(new_n7004_));
  XOR2X1   g06002(.A(new_n6615_), .B(new_n7004_), .Y(new_n7005_));
  OR2X1    g06003(.A(new_n6611_), .B(new_n6998_), .Y(new_n7006_));
  OR2X1    g06004(.A(new_n6615_), .B(new_n6613_), .Y(new_n7007_));
  OAI21X1  g06005(.A0(new_n7006_), .A1(new_n7005_), .B0(new_n7007_), .Y(new_n7008_));
  NOR2X1   g06006(.A(new_n6611_), .B(new_n6998_), .Y(new_n7009_));
  XOR2X1   g06007(.A(new_n7009_), .B(new_n7005_), .Y(new_n7010_));
  AOI21X1  g06008(.A0(new_n7008_), .A1(new_n7002_), .B0(new_n7010_), .Y(new_n7011_));
  XOR2X1   g06009(.A(new_n7011_), .B(new_n7001_), .Y(new_n7012_));
  OR4X1    g06010(.A(new_n6987_), .B(new_n6999_), .C(new_n7010_), .D(new_n6994_), .Y(new_n7013_));
  XOR2X1   g06011(.A(new_n6615_), .B(new_n6613_), .Y(new_n7014_));
  NOR2X1   g06012(.A(new_n6615_), .B(new_n6613_), .Y(new_n7015_));
  AOI21X1  g06013(.A0(new_n7009_), .A1(new_n7014_), .B0(new_n7015_), .Y(new_n7016_));
  AND2X1   g06014(.A(new_n6627_), .B(\A[108] ), .Y(new_n7017_));
  OR2X1    g06015(.A(new_n7017_), .B(new_n6629_), .Y(new_n7018_));
  XOR2X1   g06016(.A(new_n6632_), .B(new_n7018_), .Y(new_n7019_));
  XOR2X1   g06017(.A(new_n6989_), .B(new_n7019_), .Y(new_n7020_));
  OAI22X1  g06018(.A0(new_n7020_), .A1(new_n6991_), .B0(new_n7016_), .B1(new_n6994_), .Y(new_n7021_));
  OAI22X1  g06019(.A0(new_n7021_), .A1(new_n7013_), .B0(new_n7011_), .B1(new_n7001_), .Y(new_n7022_));
  MX2X1    g06020(.A(new_n7022_), .B(new_n7012_), .S0(new_n6993_), .Y(new_n7023_));
  INVX1    g06021(.A(\A[116] ), .Y(new_n7024_));
  AND2X1   g06022(.A(new_n7024_), .B(\A[115] ), .Y(new_n7025_));
  OAI21X1  g06023(.A0(new_n7024_), .A1(\A[115] ), .B0(\A[117] ), .Y(new_n7026_));
  NAND2X1  g06024(.A(new_n6585_), .B(new_n6581_), .Y(new_n7027_));
  OAI21X1  g06025(.A0(new_n7026_), .A1(new_n7025_), .B0(new_n7027_), .Y(new_n7028_));
  XOR2X1   g06026(.A(new_n6592_), .B(new_n7028_), .Y(new_n7029_));
  XOR2X1   g06027(.A(new_n6596_), .B(new_n6594_), .Y(new_n7030_));
  NOR2X1   g06028(.A(new_n6592_), .B(new_n6586_), .Y(new_n7031_));
  NOR2X1   g06029(.A(new_n6596_), .B(new_n6594_), .Y(new_n7032_));
  AOI21X1  g06030(.A0(new_n7031_), .A1(new_n7030_), .B0(new_n7032_), .Y(new_n7033_));
  XOR2X1   g06031(.A(new_n7031_), .B(new_n7030_), .Y(new_n7034_));
  OAI21X1  g06032(.A0(new_n7033_), .A1(new_n7029_), .B0(new_n7034_), .Y(new_n7035_));
  XOR2X1   g06033(.A(new_n6575_), .B(new_n6569_), .Y(new_n7036_));
  INVX1    g06034(.A(\A[121] ), .Y(new_n7037_));
  OR2X1    g06035(.A(\A[122] ), .B(new_n7037_), .Y(new_n7038_));
  AOI21X1  g06036(.A0(\A[122] ), .A1(new_n7037_), .B0(new_n6566_), .Y(new_n7039_));
  AOI22X1  g06037(.A0(new_n6567_), .A1(new_n6566_), .B0(new_n7039_), .B1(new_n7038_), .Y(new_n7040_));
  NOR4X1   g06038(.A(new_n6579_), .B(new_n6577_), .C(new_n6575_), .D(new_n7040_), .Y(new_n7041_));
  NOR4X1   g06039(.A(new_n6596_), .B(new_n6594_), .C(new_n6592_), .D(new_n6586_), .Y(new_n7042_));
  OR4X1    g06040(.A(new_n7042_), .B(new_n7029_), .C(new_n7041_), .D(new_n7036_), .Y(new_n7043_));
  XOR2X1   g06041(.A(new_n6579_), .B(new_n6577_), .Y(new_n7044_));
  NOR2X1   g06042(.A(new_n6575_), .B(new_n7040_), .Y(new_n7045_));
  NOR2X1   g06043(.A(new_n6579_), .B(new_n6577_), .Y(new_n7046_));
  AOI21X1  g06044(.A0(new_n7045_), .A1(new_n7044_), .B0(new_n7046_), .Y(new_n7047_));
  XOR2X1   g06045(.A(new_n7045_), .B(new_n7044_), .Y(new_n7048_));
  OAI21X1  g06046(.A0(new_n7047_), .A1(new_n7036_), .B0(new_n7048_), .Y(new_n7049_));
  XOR2X1   g06047(.A(new_n7049_), .B(new_n7043_), .Y(new_n7050_));
  NAND2X1  g06048(.A(new_n7050_), .B(new_n7035_), .Y(new_n7051_));
  OR2X1    g06049(.A(new_n6634_), .B(new_n6598_), .Y(new_n7052_));
  XOR2X1   g06050(.A(new_n6592_), .B(new_n6586_), .Y(new_n7053_));
  AND2X1   g06051(.A(new_n6591_), .B(\A[120] ), .Y(new_n7054_));
  OR2X1    g06052(.A(new_n7054_), .B(new_n6593_), .Y(new_n7055_));
  XOR2X1   g06053(.A(new_n6596_), .B(new_n7055_), .Y(new_n7056_));
  OR2X1    g06054(.A(new_n6592_), .B(new_n6586_), .Y(new_n7057_));
  OR2X1    g06055(.A(new_n6596_), .B(new_n6594_), .Y(new_n7058_));
  OAI21X1  g06056(.A0(new_n7057_), .A1(new_n7056_), .B0(new_n7058_), .Y(new_n7059_));
  XOR2X1   g06057(.A(new_n7031_), .B(new_n7056_), .Y(new_n7060_));
  AOI21X1  g06058(.A0(new_n7059_), .A1(new_n7053_), .B0(new_n7060_), .Y(new_n7061_));
  NOR4X1   g06059(.A(new_n7042_), .B(new_n7029_), .C(new_n7041_), .D(new_n7036_), .Y(new_n7062_));
  XOR2X1   g06060(.A(new_n6575_), .B(new_n7040_), .Y(new_n7063_));
  AND2X1   g06061(.A(new_n6574_), .B(\A[126] ), .Y(new_n7064_));
  OR2X1    g06062(.A(new_n7064_), .B(new_n6576_), .Y(new_n7065_));
  XOR2X1   g06063(.A(new_n6579_), .B(new_n7065_), .Y(new_n7066_));
  OR2X1    g06064(.A(new_n6575_), .B(new_n7040_), .Y(new_n7067_));
  OR2X1    g06065(.A(new_n6579_), .B(new_n6577_), .Y(new_n7068_));
  OAI21X1  g06066(.A0(new_n7067_), .A1(new_n7066_), .B0(new_n7068_), .Y(new_n7069_));
  XOR2X1   g06067(.A(new_n7067_), .B(new_n7044_), .Y(new_n7070_));
  AOI21X1  g06068(.A0(new_n7069_), .A1(new_n7063_), .B0(new_n7070_), .Y(new_n7071_));
  OR4X1    g06069(.A(new_n7029_), .B(new_n7041_), .C(new_n7070_), .D(new_n7036_), .Y(new_n7072_));
  OAI22X1  g06070(.A0(new_n7060_), .A1(new_n7033_), .B0(new_n7047_), .B1(new_n7036_), .Y(new_n7073_));
  OAI22X1  g06071(.A0(new_n7073_), .A1(new_n7072_), .B0(new_n7071_), .B1(new_n7062_), .Y(new_n7074_));
  AOI21X1  g06072(.A0(new_n7074_), .A1(new_n7061_), .B0(new_n7052_), .Y(new_n7075_));
  MX2X1    g06073(.A(new_n7074_), .B(new_n7050_), .S0(new_n7035_), .Y(new_n7076_));
  AOI22X1  g06074(.A0(new_n7076_), .A1(new_n7052_), .B0(new_n7075_), .B1(new_n7051_), .Y(new_n7077_));
  OR2X1    g06075(.A(new_n7077_), .B(new_n7023_), .Y(new_n7078_));
  OR2X1    g06076(.A(new_n6710_), .B(new_n6636_), .Y(new_n7079_));
  AND2X1   g06077(.A(new_n7050_), .B(new_n7035_), .Y(new_n7080_));
  XOR2X1   g06078(.A(new_n7071_), .B(new_n7043_), .Y(new_n7081_));
  NOR4X1   g06079(.A(new_n7029_), .B(new_n7070_), .C(new_n7069_), .D(new_n7036_), .Y(new_n7082_));
  AOI21X1  g06080(.A0(new_n7069_), .A1(new_n7063_), .B0(new_n7042_), .Y(new_n7083_));
  AOI22X1  g06081(.A0(new_n7083_), .A1(new_n7082_), .B0(new_n7049_), .B1(new_n7043_), .Y(new_n7084_));
  MX2X1    g06082(.A(new_n7084_), .B(new_n7081_), .S0(new_n7035_), .Y(new_n7085_));
  OAI21X1  g06083(.A0(new_n7084_), .A1(new_n7035_), .B0(new_n7052_), .Y(new_n7086_));
  OAI22X1  g06084(.A0(new_n7086_), .A1(new_n7080_), .B0(new_n7085_), .B1(new_n7052_), .Y(new_n7087_));
  AOI21X1  g06085(.A0(new_n7087_), .A1(new_n7023_), .B0(new_n7079_), .Y(new_n7088_));
  OR4X1    g06086(.A(new_n7000_), .B(new_n6987_), .C(new_n6999_), .D(new_n6994_), .Y(new_n7089_));
  XOR2X1   g06087(.A(new_n7011_), .B(new_n7089_), .Y(new_n7090_));
  XOR2X1   g06088(.A(new_n7009_), .B(new_n7014_), .Y(new_n7091_));
  OAI21X1  g06089(.A0(new_n7016_), .A1(new_n6994_), .B0(new_n7091_), .Y(new_n7092_));
  NOR4X1   g06090(.A(new_n6987_), .B(new_n7010_), .C(new_n7008_), .D(new_n6994_), .Y(new_n7093_));
  AOI21X1  g06091(.A0(new_n7008_), .A1(new_n7002_), .B0(new_n7000_), .Y(new_n7094_));
  AOI22X1  g06092(.A0(new_n7094_), .A1(new_n7093_), .B0(new_n7092_), .B1(new_n7089_), .Y(new_n7095_));
  MX2X1    g06093(.A(new_n7095_), .B(new_n7090_), .S0(new_n6993_), .Y(new_n7096_));
  NOR2X1   g06094(.A(new_n6634_), .B(new_n6598_), .Y(new_n7097_));
  OAI21X1  g06095(.A0(new_n7084_), .A1(new_n7035_), .B0(new_n7097_), .Y(new_n7098_));
  OAI22X1  g06096(.A0(new_n7085_), .A1(new_n7097_), .B0(new_n7098_), .B1(new_n7080_), .Y(new_n7099_));
  MX2X1    g06097(.A(new_n7087_), .B(new_n7099_), .S0(new_n7096_), .Y(new_n7100_));
  AOI22X1  g06098(.A0(new_n7100_), .A1(new_n7079_), .B0(new_n7088_), .B1(new_n7078_), .Y(new_n7101_));
  INVX1    g06099(.A(\A[92] ), .Y(new_n7102_));
  AND2X1   g06100(.A(new_n7102_), .B(\A[91] ), .Y(new_n7103_));
  OAI21X1  g06101(.A0(new_n7102_), .A1(\A[91] ), .B0(\A[93] ), .Y(new_n7104_));
  NAND2X1  g06102(.A(new_n6659_), .B(new_n6655_), .Y(new_n7105_));
  OAI21X1  g06103(.A0(new_n7104_), .A1(new_n7103_), .B0(new_n7105_), .Y(new_n7106_));
  XOR2X1   g06104(.A(new_n6666_), .B(new_n7106_), .Y(new_n7107_));
  XOR2X1   g06105(.A(new_n6670_), .B(new_n6668_), .Y(new_n7108_));
  NOR2X1   g06106(.A(new_n6666_), .B(new_n6660_), .Y(new_n7109_));
  NOR2X1   g06107(.A(new_n6670_), .B(new_n6668_), .Y(new_n7110_));
  AOI21X1  g06108(.A0(new_n7109_), .A1(new_n7108_), .B0(new_n7110_), .Y(new_n7111_));
  XOR2X1   g06109(.A(new_n7109_), .B(new_n7108_), .Y(new_n7112_));
  OAI21X1  g06110(.A0(new_n7111_), .A1(new_n7107_), .B0(new_n7112_), .Y(new_n7113_));
  XOR2X1   g06111(.A(new_n6649_), .B(new_n6643_), .Y(new_n7114_));
  INVX1    g06112(.A(\A[97] ), .Y(new_n7115_));
  OR2X1    g06113(.A(\A[98] ), .B(new_n7115_), .Y(new_n7116_));
  AOI21X1  g06114(.A0(\A[98] ), .A1(new_n7115_), .B0(new_n6640_), .Y(new_n7117_));
  AOI22X1  g06115(.A0(new_n6641_), .A1(new_n6640_), .B0(new_n7117_), .B1(new_n7116_), .Y(new_n7118_));
  NOR4X1   g06116(.A(new_n6653_), .B(new_n6651_), .C(new_n6649_), .D(new_n7118_), .Y(new_n7119_));
  NOR4X1   g06117(.A(new_n6670_), .B(new_n6668_), .C(new_n6666_), .D(new_n6660_), .Y(new_n7120_));
  OR4X1    g06118(.A(new_n7120_), .B(new_n7107_), .C(new_n7119_), .D(new_n7114_), .Y(new_n7121_));
  XOR2X1   g06119(.A(new_n6653_), .B(new_n6651_), .Y(new_n7122_));
  NOR2X1   g06120(.A(new_n6649_), .B(new_n7118_), .Y(new_n7123_));
  NOR2X1   g06121(.A(new_n6653_), .B(new_n6651_), .Y(new_n7124_));
  AOI21X1  g06122(.A0(new_n7123_), .A1(new_n7122_), .B0(new_n7124_), .Y(new_n7125_));
  XOR2X1   g06123(.A(new_n7123_), .B(new_n7122_), .Y(new_n7126_));
  OAI21X1  g06124(.A0(new_n7125_), .A1(new_n7114_), .B0(new_n7126_), .Y(new_n7127_));
  XOR2X1   g06125(.A(new_n7127_), .B(new_n7121_), .Y(new_n7128_));
  NAND2X1  g06126(.A(new_n7128_), .B(new_n7113_), .Y(new_n7129_));
  OR2X1    g06127(.A(new_n6709_), .B(new_n6672_), .Y(new_n7130_));
  XOR2X1   g06128(.A(new_n6666_), .B(new_n6660_), .Y(new_n7131_));
  AND2X1   g06129(.A(new_n6665_), .B(\A[96] ), .Y(new_n7132_));
  OR2X1    g06130(.A(new_n7132_), .B(new_n6667_), .Y(new_n7133_));
  XOR2X1   g06131(.A(new_n6670_), .B(new_n7133_), .Y(new_n7134_));
  OR2X1    g06132(.A(new_n6666_), .B(new_n6660_), .Y(new_n7135_));
  OR2X1    g06133(.A(new_n6670_), .B(new_n6668_), .Y(new_n7136_));
  OAI21X1  g06134(.A0(new_n7135_), .A1(new_n7134_), .B0(new_n7136_), .Y(new_n7137_));
  XOR2X1   g06135(.A(new_n7109_), .B(new_n7134_), .Y(new_n7138_));
  AOI21X1  g06136(.A0(new_n7137_), .A1(new_n7131_), .B0(new_n7138_), .Y(new_n7139_));
  NOR4X1   g06137(.A(new_n7120_), .B(new_n7107_), .C(new_n7119_), .D(new_n7114_), .Y(new_n7140_));
  XOR2X1   g06138(.A(new_n6649_), .B(new_n7118_), .Y(new_n7141_));
  AND2X1   g06139(.A(new_n6648_), .B(\A[102] ), .Y(new_n7142_));
  OR2X1    g06140(.A(new_n7142_), .B(new_n6650_), .Y(new_n7143_));
  XOR2X1   g06141(.A(new_n6653_), .B(new_n7143_), .Y(new_n7144_));
  OR2X1    g06142(.A(new_n6649_), .B(new_n7118_), .Y(new_n7145_));
  OR2X1    g06143(.A(new_n6653_), .B(new_n6651_), .Y(new_n7146_));
  OAI21X1  g06144(.A0(new_n7145_), .A1(new_n7144_), .B0(new_n7146_), .Y(new_n7147_));
  XOR2X1   g06145(.A(new_n7145_), .B(new_n7122_), .Y(new_n7148_));
  AOI21X1  g06146(.A0(new_n7147_), .A1(new_n7141_), .B0(new_n7148_), .Y(new_n7149_));
  OR4X1    g06147(.A(new_n7107_), .B(new_n7119_), .C(new_n7148_), .D(new_n7114_), .Y(new_n7150_));
  OAI22X1  g06148(.A0(new_n7138_), .A1(new_n7111_), .B0(new_n7125_), .B1(new_n7114_), .Y(new_n7151_));
  OAI22X1  g06149(.A0(new_n7151_), .A1(new_n7150_), .B0(new_n7149_), .B1(new_n7140_), .Y(new_n7152_));
  AOI21X1  g06150(.A0(new_n7152_), .A1(new_n7139_), .B0(new_n7130_), .Y(new_n7153_));
  MX2X1    g06151(.A(new_n7152_), .B(new_n7128_), .S0(new_n7113_), .Y(new_n7154_));
  AOI22X1  g06152(.A0(new_n7154_), .A1(new_n7130_), .B0(new_n7153_), .B1(new_n7129_), .Y(new_n7155_));
  INVX1    g06153(.A(\A[80] ), .Y(new_n7156_));
  AND2X1   g06154(.A(new_n7156_), .B(\A[79] ), .Y(new_n7157_));
  OAI21X1  g06155(.A0(new_n7156_), .A1(\A[79] ), .B0(\A[81] ), .Y(new_n7158_));
  NAND2X1  g06156(.A(new_n6696_), .B(new_n6692_), .Y(new_n7159_));
  OAI21X1  g06157(.A0(new_n7158_), .A1(new_n7157_), .B0(new_n7159_), .Y(new_n7160_));
  XOR2X1   g06158(.A(new_n6703_), .B(new_n7160_), .Y(new_n7161_));
  XOR2X1   g06159(.A(new_n6707_), .B(new_n6705_), .Y(new_n7162_));
  NOR2X1   g06160(.A(new_n6703_), .B(new_n6697_), .Y(new_n7163_));
  NOR2X1   g06161(.A(new_n6707_), .B(new_n6705_), .Y(new_n7164_));
  AOI21X1  g06162(.A0(new_n7163_), .A1(new_n7162_), .B0(new_n7164_), .Y(new_n7165_));
  XOR2X1   g06163(.A(new_n7163_), .B(new_n7162_), .Y(new_n7166_));
  OAI21X1  g06164(.A0(new_n7165_), .A1(new_n7161_), .B0(new_n7166_), .Y(new_n7167_));
  XOR2X1   g06165(.A(new_n6686_), .B(new_n6680_), .Y(new_n7168_));
  INVX1    g06166(.A(\A[85] ), .Y(new_n7169_));
  OR2X1    g06167(.A(\A[86] ), .B(new_n7169_), .Y(new_n7170_));
  AOI21X1  g06168(.A0(\A[86] ), .A1(new_n7169_), .B0(new_n6677_), .Y(new_n7171_));
  AOI22X1  g06169(.A0(new_n6678_), .A1(new_n6677_), .B0(new_n7171_), .B1(new_n7170_), .Y(new_n7172_));
  NOR4X1   g06170(.A(new_n6690_), .B(new_n6688_), .C(new_n6686_), .D(new_n7172_), .Y(new_n7173_));
  NOR4X1   g06171(.A(new_n6707_), .B(new_n6705_), .C(new_n6703_), .D(new_n6697_), .Y(new_n7174_));
  OR4X1    g06172(.A(new_n7174_), .B(new_n7161_), .C(new_n7173_), .D(new_n7168_), .Y(new_n7175_));
  XOR2X1   g06173(.A(new_n6686_), .B(new_n7172_), .Y(new_n7176_));
  AND2X1   g06174(.A(new_n6685_), .B(\A[90] ), .Y(new_n7177_));
  OR2X1    g06175(.A(new_n7177_), .B(new_n6687_), .Y(new_n7178_));
  XOR2X1   g06176(.A(new_n6690_), .B(new_n7178_), .Y(new_n7179_));
  OR2X1    g06177(.A(new_n6686_), .B(new_n7172_), .Y(new_n7180_));
  OR2X1    g06178(.A(new_n6690_), .B(new_n6688_), .Y(new_n7181_));
  OAI21X1  g06179(.A0(new_n7180_), .A1(new_n7179_), .B0(new_n7181_), .Y(new_n7182_));
  NOR2X1   g06180(.A(new_n6686_), .B(new_n7172_), .Y(new_n7183_));
  XOR2X1   g06181(.A(new_n7183_), .B(new_n7179_), .Y(new_n7184_));
  AOI21X1  g06182(.A0(new_n7182_), .A1(new_n7176_), .B0(new_n7184_), .Y(new_n7185_));
  XOR2X1   g06183(.A(new_n7185_), .B(new_n7175_), .Y(new_n7186_));
  XOR2X1   g06184(.A(new_n6690_), .B(new_n6688_), .Y(new_n7187_));
  NOR2X1   g06185(.A(new_n6690_), .B(new_n6688_), .Y(new_n7188_));
  AOI21X1  g06186(.A0(new_n7183_), .A1(new_n7187_), .B0(new_n7188_), .Y(new_n7189_));
  XOR2X1   g06187(.A(new_n7183_), .B(new_n7187_), .Y(new_n7190_));
  OAI21X1  g06188(.A0(new_n7189_), .A1(new_n7168_), .B0(new_n7190_), .Y(new_n7191_));
  NOR4X1   g06189(.A(new_n7161_), .B(new_n7184_), .C(new_n7182_), .D(new_n7168_), .Y(new_n7192_));
  AOI21X1  g06190(.A0(new_n7182_), .A1(new_n7176_), .B0(new_n7174_), .Y(new_n7193_));
  AOI22X1  g06191(.A0(new_n7193_), .A1(new_n7192_), .B0(new_n7191_), .B1(new_n7175_), .Y(new_n7194_));
  MX2X1    g06192(.A(new_n7194_), .B(new_n7186_), .S0(new_n7167_), .Y(new_n7195_));
  NOR2X1   g06193(.A(new_n6709_), .B(new_n6672_), .Y(new_n7196_));
  AOI21X1  g06194(.A0(new_n7152_), .A1(new_n7139_), .B0(new_n7196_), .Y(new_n7197_));
  AOI22X1  g06195(.A0(new_n7197_), .A1(new_n7129_), .B0(new_n7154_), .B1(new_n7196_), .Y(new_n7198_));
  MX2X1    g06196(.A(new_n7198_), .B(new_n7155_), .S0(new_n7195_), .Y(new_n7199_));
  NOR2X1   g06197(.A(new_n6710_), .B(new_n6636_), .Y(new_n7200_));
  AOI21X1  g06198(.A0(new_n7087_), .A1(new_n7023_), .B0(new_n7200_), .Y(new_n7201_));
  AOI22X1  g06199(.A0(new_n7201_), .A1(new_n7078_), .B0(new_n7100_), .B1(new_n7200_), .Y(new_n7202_));
  MX2X1    g06200(.A(new_n7202_), .B(new_n7101_), .S0(new_n7199_), .Y(new_n7203_));
  AOI21X1  g06201(.A0(new_n6955_), .A1(new_n6824_), .B0(new_n6948_), .Y(new_n7204_));
  AOI22X1  g06202(.A0(new_n7204_), .A1(new_n6946_), .B0(new_n6980_), .B1(new_n6948_), .Y(new_n7205_));
  MX2X1    g06203(.A(new_n7205_), .B(new_n6981_), .S0(new_n7203_), .Y(new_n7206_));
  AOI21X1  g06204(.A0(new_n6720_), .A1(new_n6013_), .B0(new_n6713_), .Y(new_n7207_));
  AOI22X1  g06205(.A0(new_n7207_), .A1(new_n6413_), .B0(new_n6734_), .B1(new_n6713_), .Y(new_n7208_));
  MX2X1    g06206(.A(new_n7208_), .B(new_n6735_), .S0(new_n7206_), .Y(new_n7209_));
  INVX1    g06207(.A(\A[333] ), .Y(new_n7210_));
  INVX1    g06208(.A(\A[332] ), .Y(new_n7211_));
  OR2X1    g06209(.A(new_n7211_), .B(\A[331] ), .Y(new_n7212_));
  AOI21X1  g06210(.A0(new_n7211_), .A1(\A[331] ), .B0(new_n7210_), .Y(new_n7213_));
  XOR2X1   g06211(.A(\A[332] ), .B(\A[331] ), .Y(new_n7214_));
  AOI22X1  g06212(.A0(new_n7214_), .A1(new_n7210_), .B0(new_n7213_), .B1(new_n7212_), .Y(new_n7215_));
  INVX1    g06213(.A(\A[336] ), .Y(new_n7216_));
  INVX1    g06214(.A(\A[335] ), .Y(new_n7217_));
  OR2X1    g06215(.A(new_n7217_), .B(\A[334] ), .Y(new_n7218_));
  AOI21X1  g06216(.A0(new_n7217_), .A1(\A[334] ), .B0(new_n7216_), .Y(new_n7219_));
  XOR2X1   g06217(.A(\A[335] ), .B(\A[334] ), .Y(new_n7220_));
  AOI22X1  g06218(.A0(new_n7220_), .A1(new_n7216_), .B0(new_n7219_), .B1(new_n7218_), .Y(new_n7221_));
  OR2X1    g06219(.A(new_n7221_), .B(new_n7215_), .Y(new_n7222_));
  AND2X1   g06220(.A(\A[335] ), .B(\A[334] ), .Y(new_n7223_));
  AND2X1   g06221(.A(new_n7220_), .B(\A[336] ), .Y(new_n7224_));
  OR2X1    g06222(.A(new_n7224_), .B(new_n7223_), .Y(new_n7225_));
  AND2X1   g06223(.A(\A[332] ), .B(\A[331] ), .Y(new_n7226_));
  AOI21X1  g06224(.A0(new_n7214_), .A1(\A[333] ), .B0(new_n7226_), .Y(new_n7227_));
  XOR2X1   g06225(.A(new_n7227_), .B(new_n7225_), .Y(new_n7228_));
  XOR2X1   g06226(.A(new_n7228_), .B(new_n7222_), .Y(new_n7229_));
  INVX1    g06227(.A(\A[331] ), .Y(new_n7230_));
  AND2X1   g06228(.A(\A[332] ), .B(new_n7230_), .Y(new_n7231_));
  OAI21X1  g06229(.A0(\A[332] ), .A1(new_n7230_), .B0(\A[333] ), .Y(new_n7232_));
  NAND2X1  g06230(.A(new_n7214_), .B(new_n7210_), .Y(new_n7233_));
  OAI21X1  g06231(.A0(new_n7232_), .A1(new_n7231_), .B0(new_n7233_), .Y(new_n7234_));
  XOR2X1   g06232(.A(new_n7221_), .B(new_n7234_), .Y(new_n7235_));
  NOR2X1   g06233(.A(new_n7221_), .B(new_n7215_), .Y(new_n7236_));
  AOI21X1  g06234(.A0(new_n7220_), .A1(\A[336] ), .B0(new_n7223_), .Y(new_n7237_));
  XOR2X1   g06235(.A(new_n7227_), .B(new_n7237_), .Y(new_n7238_));
  NOR2X1   g06236(.A(new_n7227_), .B(new_n7237_), .Y(new_n7239_));
  AOI21X1  g06237(.A0(new_n7238_), .A1(new_n7236_), .B0(new_n7239_), .Y(new_n7240_));
  OAI21X1  g06238(.A0(new_n7240_), .A1(new_n7235_), .B0(new_n7229_), .Y(new_n7241_));
  AND2X1   g06239(.A(\A[341] ), .B(\A[340] ), .Y(new_n7242_));
  XOR2X1   g06240(.A(\A[341] ), .B(\A[340] ), .Y(new_n7243_));
  AOI21X1  g06241(.A0(new_n7243_), .A1(\A[342] ), .B0(new_n7242_), .Y(new_n7244_));
  AND2X1   g06242(.A(\A[338] ), .B(\A[337] ), .Y(new_n7245_));
  XOR2X1   g06243(.A(\A[338] ), .B(\A[337] ), .Y(new_n7246_));
  AOI21X1  g06244(.A0(new_n7246_), .A1(\A[339] ), .B0(new_n7245_), .Y(new_n7247_));
  INVX1    g06245(.A(\A[339] ), .Y(new_n7248_));
  INVX1    g06246(.A(\A[338] ), .Y(new_n7249_));
  OR2X1    g06247(.A(new_n7249_), .B(\A[337] ), .Y(new_n7250_));
  AOI21X1  g06248(.A0(new_n7249_), .A1(\A[337] ), .B0(new_n7248_), .Y(new_n7251_));
  AOI22X1  g06249(.A0(new_n7251_), .A1(new_n7250_), .B0(new_n7246_), .B1(new_n7248_), .Y(new_n7252_));
  INVX1    g06250(.A(\A[342] ), .Y(new_n7253_));
  INVX1    g06251(.A(\A[341] ), .Y(new_n7254_));
  OR2X1    g06252(.A(new_n7254_), .B(\A[340] ), .Y(new_n7255_));
  AOI21X1  g06253(.A0(new_n7254_), .A1(\A[340] ), .B0(new_n7253_), .Y(new_n7256_));
  AOI22X1  g06254(.A0(new_n7256_), .A1(new_n7255_), .B0(new_n7243_), .B1(new_n7253_), .Y(new_n7257_));
  NOR4X1   g06255(.A(new_n7257_), .B(new_n7252_), .C(new_n7247_), .D(new_n7244_), .Y(new_n7258_));
  NOR4X1   g06256(.A(new_n7227_), .B(new_n7237_), .C(new_n7221_), .D(new_n7215_), .Y(new_n7259_));
  INVX1    g06257(.A(\A[337] ), .Y(new_n7260_));
  AND2X1   g06258(.A(\A[338] ), .B(new_n7260_), .Y(new_n7261_));
  OAI21X1  g06259(.A0(\A[338] ), .A1(new_n7260_), .B0(\A[339] ), .Y(new_n7262_));
  NAND2X1  g06260(.A(new_n7246_), .B(new_n7248_), .Y(new_n7263_));
  OAI21X1  g06261(.A0(new_n7262_), .A1(new_n7261_), .B0(new_n7263_), .Y(new_n7264_));
  XOR2X1   g06262(.A(new_n7257_), .B(new_n7264_), .Y(new_n7265_));
  OR4X1    g06263(.A(new_n7265_), .B(new_n7259_), .C(new_n7258_), .D(new_n7235_), .Y(new_n7266_));
  XOR2X1   g06264(.A(new_n7247_), .B(new_n7244_), .Y(new_n7267_));
  NOR2X1   g06265(.A(new_n7257_), .B(new_n7252_), .Y(new_n7268_));
  NOR2X1   g06266(.A(new_n7247_), .B(new_n7244_), .Y(new_n7269_));
  AOI21X1  g06267(.A0(new_n7268_), .A1(new_n7267_), .B0(new_n7269_), .Y(new_n7270_));
  XOR2X1   g06268(.A(new_n7268_), .B(new_n7267_), .Y(new_n7271_));
  OAI21X1  g06269(.A0(new_n7265_), .A1(new_n7270_), .B0(new_n7271_), .Y(new_n7272_));
  XOR2X1   g06270(.A(new_n7272_), .B(new_n7266_), .Y(new_n7273_));
  NAND2X1  g06271(.A(new_n7273_), .B(new_n7241_), .Y(new_n7274_));
  XOR2X1   g06272(.A(new_n7221_), .B(new_n7215_), .Y(new_n7275_));
  OAI21X1  g06273(.A0(new_n7265_), .A1(new_n7258_), .B0(new_n7275_), .Y(new_n7276_));
  OR4X1    g06274(.A(new_n7257_), .B(new_n7252_), .C(new_n7247_), .D(new_n7244_), .Y(new_n7277_));
  XOR2X1   g06275(.A(new_n7257_), .B(new_n7252_), .Y(new_n7278_));
  XOR2X1   g06276(.A(new_n7221_), .B(new_n7234_), .Y(new_n7279_));
  NAND3X1  g06277(.A(new_n7279_), .B(new_n7278_), .C(new_n7277_), .Y(new_n7280_));
  AND2X1   g06278(.A(new_n7280_), .B(new_n7276_), .Y(new_n7281_));
  INVX1    g06279(.A(\A[326] ), .Y(new_n7282_));
  AND2X1   g06280(.A(new_n7282_), .B(\A[325] ), .Y(new_n7283_));
  OAI21X1  g06281(.A0(new_n7282_), .A1(\A[325] ), .B0(\A[327] ), .Y(new_n7284_));
  INVX1    g06282(.A(\A[327] ), .Y(new_n7285_));
  XOR2X1   g06283(.A(\A[326] ), .B(\A[325] ), .Y(new_n7286_));
  NAND2X1  g06284(.A(new_n7286_), .B(new_n7285_), .Y(new_n7287_));
  OAI21X1  g06285(.A0(new_n7284_), .A1(new_n7283_), .B0(new_n7287_), .Y(new_n7288_));
  INVX1    g06286(.A(\A[330] ), .Y(new_n7289_));
  INVX1    g06287(.A(\A[328] ), .Y(new_n7290_));
  OR2X1    g06288(.A(\A[329] ), .B(new_n7290_), .Y(new_n7291_));
  AOI21X1  g06289(.A0(\A[329] ), .A1(new_n7290_), .B0(new_n7289_), .Y(new_n7292_));
  XOR2X1   g06290(.A(\A[329] ), .B(\A[328] ), .Y(new_n7293_));
  AOI22X1  g06291(.A0(new_n7293_), .A1(new_n7289_), .B0(new_n7292_), .B1(new_n7291_), .Y(new_n7294_));
  AND2X1   g06292(.A(\A[329] ), .B(\A[328] ), .Y(new_n7295_));
  AOI21X1  g06293(.A0(new_n7293_), .A1(\A[330] ), .B0(new_n7295_), .Y(new_n7296_));
  AND2X1   g06294(.A(\A[326] ), .B(\A[325] ), .Y(new_n7297_));
  AOI21X1  g06295(.A0(new_n7286_), .A1(\A[327] ), .B0(new_n7297_), .Y(new_n7298_));
  XOR2X1   g06296(.A(new_n7294_), .B(new_n7288_), .Y(new_n7299_));
  INVX1    g06297(.A(\A[321] ), .Y(new_n7300_));
  INVX1    g06298(.A(\A[319] ), .Y(new_n7301_));
  OR2X1    g06299(.A(\A[320] ), .B(new_n7301_), .Y(new_n7302_));
  AOI21X1  g06300(.A0(\A[320] ), .A1(new_n7301_), .B0(new_n7300_), .Y(new_n7303_));
  XOR2X1   g06301(.A(\A[320] ), .B(\A[319] ), .Y(new_n7304_));
  AOI22X1  g06302(.A0(new_n7304_), .A1(new_n7300_), .B0(new_n7303_), .B1(new_n7302_), .Y(new_n7305_));
  INVX1    g06303(.A(\A[324] ), .Y(new_n7306_));
  INVX1    g06304(.A(\A[322] ), .Y(new_n7307_));
  OR2X1    g06305(.A(\A[323] ), .B(new_n7307_), .Y(new_n7308_));
  AOI21X1  g06306(.A0(\A[323] ), .A1(new_n7307_), .B0(new_n7306_), .Y(new_n7309_));
  XOR2X1   g06307(.A(\A[323] ), .B(\A[322] ), .Y(new_n7310_));
  AOI22X1  g06308(.A0(new_n7310_), .A1(new_n7306_), .B0(new_n7309_), .B1(new_n7308_), .Y(new_n7311_));
  AND2X1   g06309(.A(\A[323] ), .B(\A[322] ), .Y(new_n7312_));
  AOI21X1  g06310(.A0(new_n7310_), .A1(\A[324] ), .B0(new_n7312_), .Y(new_n7313_));
  AND2X1   g06311(.A(\A[320] ), .B(\A[319] ), .Y(new_n7314_));
  AOI21X1  g06312(.A0(new_n7304_), .A1(\A[321] ), .B0(new_n7314_), .Y(new_n7315_));
  XOR2X1   g06313(.A(new_n7311_), .B(new_n7305_), .Y(new_n7316_));
  XOR2X1   g06314(.A(new_n7316_), .B(new_n7299_), .Y(new_n7317_));
  OR2X1    g06315(.A(new_n7317_), .B(new_n7281_), .Y(new_n7318_));
  XOR2X1   g06316(.A(new_n7228_), .B(new_n7236_), .Y(new_n7319_));
  XOR2X1   g06317(.A(new_n7221_), .B(new_n7215_), .Y(new_n7320_));
  OR2X1    g06318(.A(new_n7227_), .B(new_n7237_), .Y(new_n7321_));
  OAI21X1  g06319(.A0(new_n7228_), .A1(new_n7222_), .B0(new_n7321_), .Y(new_n7322_));
  AOI21X1  g06320(.A0(new_n7322_), .A1(new_n7320_), .B0(new_n7319_), .Y(new_n7323_));
  NOR4X1   g06321(.A(new_n7265_), .B(new_n7259_), .C(new_n7258_), .D(new_n7235_), .Y(new_n7324_));
  AND2X1   g06322(.A(new_n7243_), .B(\A[342] ), .Y(new_n7325_));
  OR2X1    g06323(.A(new_n7325_), .B(new_n7242_), .Y(new_n7326_));
  XOR2X1   g06324(.A(new_n7247_), .B(new_n7326_), .Y(new_n7327_));
  OR2X1    g06325(.A(new_n7257_), .B(new_n7252_), .Y(new_n7328_));
  OR2X1    g06326(.A(new_n7247_), .B(new_n7244_), .Y(new_n7329_));
  OAI21X1  g06327(.A0(new_n7328_), .A1(new_n7327_), .B0(new_n7329_), .Y(new_n7330_));
  XOR2X1   g06328(.A(new_n7268_), .B(new_n7327_), .Y(new_n7331_));
  AOI21X1  g06329(.A0(new_n7278_), .A1(new_n7330_), .B0(new_n7331_), .Y(new_n7332_));
  OR4X1    g06330(.A(new_n7265_), .B(new_n7259_), .C(new_n7331_), .D(new_n7235_), .Y(new_n7333_));
  AOI21X1  g06331(.A0(new_n7265_), .A1(new_n7331_), .B0(new_n7270_), .Y(new_n7334_));
  OAI22X1  g06332(.A0(new_n7334_), .A1(new_n7333_), .B0(new_n7332_), .B1(new_n7324_), .Y(new_n7335_));
  AOI21X1  g06333(.A0(new_n7335_), .A1(new_n7323_), .B0(new_n7318_), .Y(new_n7336_));
  MX2X1    g06334(.A(new_n7335_), .B(new_n7273_), .S0(new_n7241_), .Y(new_n7337_));
  AOI22X1  g06335(.A0(new_n7337_), .A1(new_n7318_), .B0(new_n7336_), .B1(new_n7274_), .Y(new_n7338_));
  INVX1    g06336(.A(\A[320] ), .Y(new_n7339_));
  AND2X1   g06337(.A(new_n7339_), .B(\A[319] ), .Y(new_n7340_));
  OAI21X1  g06338(.A0(new_n7339_), .A1(\A[319] ), .B0(\A[321] ), .Y(new_n7341_));
  NAND2X1  g06339(.A(new_n7304_), .B(new_n7300_), .Y(new_n7342_));
  OAI21X1  g06340(.A0(new_n7341_), .A1(new_n7340_), .B0(new_n7342_), .Y(new_n7343_));
  XOR2X1   g06341(.A(new_n7311_), .B(new_n7343_), .Y(new_n7344_));
  XOR2X1   g06342(.A(new_n7315_), .B(new_n7313_), .Y(new_n7345_));
  NOR2X1   g06343(.A(new_n7311_), .B(new_n7305_), .Y(new_n7346_));
  NOR2X1   g06344(.A(new_n7315_), .B(new_n7313_), .Y(new_n7347_));
  AOI21X1  g06345(.A0(new_n7346_), .A1(new_n7345_), .B0(new_n7347_), .Y(new_n7348_));
  XOR2X1   g06346(.A(new_n7346_), .B(new_n7345_), .Y(new_n7349_));
  OAI21X1  g06347(.A0(new_n7348_), .A1(new_n7344_), .B0(new_n7349_), .Y(new_n7350_));
  XOR2X1   g06348(.A(new_n7294_), .B(new_n7288_), .Y(new_n7351_));
  INVX1    g06349(.A(\A[325] ), .Y(new_n7352_));
  OR2X1    g06350(.A(\A[326] ), .B(new_n7352_), .Y(new_n7353_));
  AOI21X1  g06351(.A0(\A[326] ), .A1(new_n7352_), .B0(new_n7285_), .Y(new_n7354_));
  AOI22X1  g06352(.A0(new_n7286_), .A1(new_n7285_), .B0(new_n7354_), .B1(new_n7353_), .Y(new_n7355_));
  NOR4X1   g06353(.A(new_n7298_), .B(new_n7296_), .C(new_n7294_), .D(new_n7355_), .Y(new_n7356_));
  NOR4X1   g06354(.A(new_n7315_), .B(new_n7313_), .C(new_n7311_), .D(new_n7305_), .Y(new_n7357_));
  OR4X1    g06355(.A(new_n7357_), .B(new_n7344_), .C(new_n7356_), .D(new_n7351_), .Y(new_n7358_));
  XOR2X1   g06356(.A(new_n7294_), .B(new_n7355_), .Y(new_n7359_));
  AND2X1   g06357(.A(new_n7293_), .B(\A[330] ), .Y(new_n7360_));
  OR2X1    g06358(.A(new_n7360_), .B(new_n7295_), .Y(new_n7361_));
  XOR2X1   g06359(.A(new_n7298_), .B(new_n7361_), .Y(new_n7362_));
  OR2X1    g06360(.A(new_n7294_), .B(new_n7355_), .Y(new_n7363_));
  OR2X1    g06361(.A(new_n7298_), .B(new_n7296_), .Y(new_n7364_));
  OAI21X1  g06362(.A0(new_n7363_), .A1(new_n7362_), .B0(new_n7364_), .Y(new_n7365_));
  NOR2X1   g06363(.A(new_n7294_), .B(new_n7355_), .Y(new_n7366_));
  XOR2X1   g06364(.A(new_n7366_), .B(new_n7362_), .Y(new_n7367_));
  AOI21X1  g06365(.A0(new_n7365_), .A1(new_n7359_), .B0(new_n7367_), .Y(new_n7368_));
  XOR2X1   g06366(.A(new_n7368_), .B(new_n7358_), .Y(new_n7369_));
  XOR2X1   g06367(.A(new_n7298_), .B(new_n7296_), .Y(new_n7370_));
  NOR2X1   g06368(.A(new_n7298_), .B(new_n7296_), .Y(new_n7371_));
  AOI21X1  g06369(.A0(new_n7366_), .A1(new_n7370_), .B0(new_n7371_), .Y(new_n7372_));
  XOR2X1   g06370(.A(new_n7366_), .B(new_n7370_), .Y(new_n7373_));
  OAI21X1  g06371(.A0(new_n7372_), .A1(new_n7351_), .B0(new_n7373_), .Y(new_n7374_));
  NOR4X1   g06372(.A(new_n7344_), .B(new_n7367_), .C(new_n7365_), .D(new_n7351_), .Y(new_n7375_));
  AOI21X1  g06373(.A0(new_n7365_), .A1(new_n7359_), .B0(new_n7357_), .Y(new_n7376_));
  AOI22X1  g06374(.A0(new_n7376_), .A1(new_n7375_), .B0(new_n7374_), .B1(new_n7358_), .Y(new_n7377_));
  MX2X1    g06375(.A(new_n7377_), .B(new_n7369_), .S0(new_n7350_), .Y(new_n7378_));
  AOI21X1  g06376(.A0(new_n7280_), .A1(new_n7276_), .B0(new_n7317_), .Y(new_n7379_));
  AOI21X1  g06377(.A0(new_n7335_), .A1(new_n7323_), .B0(new_n7379_), .Y(new_n7380_));
  AOI22X1  g06378(.A0(new_n7380_), .A1(new_n7274_), .B0(new_n7337_), .B1(new_n7379_), .Y(new_n7381_));
  MX2X1    g06379(.A(new_n7381_), .B(new_n7338_), .S0(new_n7378_), .Y(new_n7382_));
  INVX1    g06380(.A(\A[345] ), .Y(new_n7383_));
  INVX1    g06381(.A(\A[344] ), .Y(new_n7384_));
  OR2X1    g06382(.A(new_n7384_), .B(\A[343] ), .Y(new_n7385_));
  AOI21X1  g06383(.A0(new_n7384_), .A1(\A[343] ), .B0(new_n7383_), .Y(new_n7386_));
  XOR2X1   g06384(.A(\A[344] ), .B(\A[343] ), .Y(new_n7387_));
  AOI22X1  g06385(.A0(new_n7387_), .A1(new_n7383_), .B0(new_n7386_), .B1(new_n7385_), .Y(new_n7388_));
  INVX1    g06386(.A(\A[348] ), .Y(new_n7389_));
  INVX1    g06387(.A(\A[347] ), .Y(new_n7390_));
  OR2X1    g06388(.A(new_n7390_), .B(\A[346] ), .Y(new_n7391_));
  AOI21X1  g06389(.A0(new_n7390_), .A1(\A[346] ), .B0(new_n7389_), .Y(new_n7392_));
  XOR2X1   g06390(.A(\A[347] ), .B(\A[346] ), .Y(new_n7393_));
  AOI22X1  g06391(.A0(new_n7393_), .A1(new_n7389_), .B0(new_n7392_), .B1(new_n7391_), .Y(new_n7394_));
  OR2X1    g06392(.A(new_n7394_), .B(new_n7388_), .Y(new_n7395_));
  AND2X1   g06393(.A(\A[347] ), .B(\A[346] ), .Y(new_n7396_));
  AND2X1   g06394(.A(new_n7393_), .B(\A[348] ), .Y(new_n7397_));
  OR2X1    g06395(.A(new_n7397_), .B(new_n7396_), .Y(new_n7398_));
  AND2X1   g06396(.A(\A[344] ), .B(\A[343] ), .Y(new_n7399_));
  AOI21X1  g06397(.A0(new_n7387_), .A1(\A[345] ), .B0(new_n7399_), .Y(new_n7400_));
  XOR2X1   g06398(.A(new_n7400_), .B(new_n7398_), .Y(new_n7401_));
  XOR2X1   g06399(.A(new_n7401_), .B(new_n7395_), .Y(new_n7402_));
  INVX1    g06400(.A(\A[343] ), .Y(new_n7403_));
  AND2X1   g06401(.A(\A[344] ), .B(new_n7403_), .Y(new_n7404_));
  OAI21X1  g06402(.A0(\A[344] ), .A1(new_n7403_), .B0(\A[345] ), .Y(new_n7405_));
  NAND2X1  g06403(.A(new_n7387_), .B(new_n7383_), .Y(new_n7406_));
  OAI21X1  g06404(.A0(new_n7405_), .A1(new_n7404_), .B0(new_n7406_), .Y(new_n7407_));
  XOR2X1   g06405(.A(new_n7394_), .B(new_n7407_), .Y(new_n7408_));
  NOR2X1   g06406(.A(new_n7394_), .B(new_n7388_), .Y(new_n7409_));
  AOI21X1  g06407(.A0(new_n7393_), .A1(\A[348] ), .B0(new_n7396_), .Y(new_n7410_));
  XOR2X1   g06408(.A(new_n7400_), .B(new_n7410_), .Y(new_n7411_));
  NOR2X1   g06409(.A(new_n7400_), .B(new_n7410_), .Y(new_n7412_));
  AOI21X1  g06410(.A0(new_n7411_), .A1(new_n7409_), .B0(new_n7412_), .Y(new_n7413_));
  OAI21X1  g06411(.A0(new_n7413_), .A1(new_n7408_), .B0(new_n7402_), .Y(new_n7414_));
  AND2X1   g06412(.A(\A[353] ), .B(\A[352] ), .Y(new_n7415_));
  XOR2X1   g06413(.A(\A[353] ), .B(\A[352] ), .Y(new_n7416_));
  AOI21X1  g06414(.A0(new_n7416_), .A1(\A[354] ), .B0(new_n7415_), .Y(new_n7417_));
  AND2X1   g06415(.A(\A[350] ), .B(\A[349] ), .Y(new_n7418_));
  XOR2X1   g06416(.A(\A[350] ), .B(\A[349] ), .Y(new_n7419_));
  AOI21X1  g06417(.A0(new_n7419_), .A1(\A[351] ), .B0(new_n7418_), .Y(new_n7420_));
  INVX1    g06418(.A(\A[351] ), .Y(new_n7421_));
  INVX1    g06419(.A(\A[350] ), .Y(new_n7422_));
  OR2X1    g06420(.A(new_n7422_), .B(\A[349] ), .Y(new_n7423_));
  AOI21X1  g06421(.A0(new_n7422_), .A1(\A[349] ), .B0(new_n7421_), .Y(new_n7424_));
  AOI22X1  g06422(.A0(new_n7424_), .A1(new_n7423_), .B0(new_n7419_), .B1(new_n7421_), .Y(new_n7425_));
  INVX1    g06423(.A(\A[354] ), .Y(new_n7426_));
  INVX1    g06424(.A(\A[353] ), .Y(new_n7427_));
  OR2X1    g06425(.A(new_n7427_), .B(\A[352] ), .Y(new_n7428_));
  AOI21X1  g06426(.A0(new_n7427_), .A1(\A[352] ), .B0(new_n7426_), .Y(new_n7429_));
  AOI22X1  g06427(.A0(new_n7429_), .A1(new_n7428_), .B0(new_n7416_), .B1(new_n7426_), .Y(new_n7430_));
  NOR4X1   g06428(.A(new_n7430_), .B(new_n7425_), .C(new_n7420_), .D(new_n7417_), .Y(new_n7431_));
  NOR4X1   g06429(.A(new_n7400_), .B(new_n7410_), .C(new_n7394_), .D(new_n7388_), .Y(new_n7432_));
  INVX1    g06430(.A(\A[349] ), .Y(new_n7433_));
  AND2X1   g06431(.A(\A[350] ), .B(new_n7433_), .Y(new_n7434_));
  OAI21X1  g06432(.A0(\A[350] ), .A1(new_n7433_), .B0(\A[351] ), .Y(new_n7435_));
  NAND2X1  g06433(.A(new_n7419_), .B(new_n7421_), .Y(new_n7436_));
  OAI21X1  g06434(.A0(new_n7435_), .A1(new_n7434_), .B0(new_n7436_), .Y(new_n7437_));
  XOR2X1   g06435(.A(new_n7430_), .B(new_n7437_), .Y(new_n7438_));
  OR4X1    g06436(.A(new_n7438_), .B(new_n7432_), .C(new_n7431_), .D(new_n7408_), .Y(new_n7439_));
  AND2X1   g06437(.A(new_n7416_), .B(\A[354] ), .Y(new_n7440_));
  OR2X1    g06438(.A(new_n7440_), .B(new_n7415_), .Y(new_n7441_));
  XOR2X1   g06439(.A(new_n7420_), .B(new_n7441_), .Y(new_n7442_));
  OR2X1    g06440(.A(new_n7430_), .B(new_n7425_), .Y(new_n7443_));
  OR2X1    g06441(.A(new_n7420_), .B(new_n7417_), .Y(new_n7444_));
  OAI21X1  g06442(.A0(new_n7443_), .A1(new_n7442_), .B0(new_n7444_), .Y(new_n7445_));
  NOR2X1   g06443(.A(new_n7430_), .B(new_n7425_), .Y(new_n7446_));
  XOR2X1   g06444(.A(new_n7446_), .B(new_n7442_), .Y(new_n7447_));
  XOR2X1   g06445(.A(new_n7430_), .B(new_n7425_), .Y(new_n7448_));
  AOI21X1  g06446(.A0(new_n7448_), .A1(new_n7445_), .B0(new_n7447_), .Y(new_n7449_));
  XOR2X1   g06447(.A(new_n7449_), .B(new_n7439_), .Y(new_n7450_));
  XOR2X1   g06448(.A(new_n7420_), .B(new_n7417_), .Y(new_n7451_));
  NOR2X1   g06449(.A(new_n7420_), .B(new_n7417_), .Y(new_n7452_));
  AOI21X1  g06450(.A0(new_n7446_), .A1(new_n7451_), .B0(new_n7452_), .Y(new_n7453_));
  XOR2X1   g06451(.A(new_n7446_), .B(new_n7451_), .Y(new_n7454_));
  OAI21X1  g06452(.A0(new_n7438_), .A1(new_n7453_), .B0(new_n7454_), .Y(new_n7455_));
  NOR4X1   g06453(.A(new_n7438_), .B(new_n7432_), .C(new_n7447_), .D(new_n7408_), .Y(new_n7456_));
  OAI21X1  g06454(.A0(new_n7448_), .A1(new_n7454_), .B0(new_n7445_), .Y(new_n7457_));
  AOI22X1  g06455(.A0(new_n7457_), .A1(new_n7456_), .B0(new_n7455_), .B1(new_n7439_), .Y(new_n7458_));
  MX2X1    g06456(.A(new_n7458_), .B(new_n7450_), .S0(new_n7414_), .Y(new_n7459_));
  INVX1    g06457(.A(\A[357] ), .Y(new_n7460_));
  INVX1    g06458(.A(\A[356] ), .Y(new_n7461_));
  OR2X1    g06459(.A(new_n7461_), .B(\A[355] ), .Y(new_n7462_));
  AOI21X1  g06460(.A0(new_n7461_), .A1(\A[355] ), .B0(new_n7460_), .Y(new_n7463_));
  XOR2X1   g06461(.A(\A[356] ), .B(\A[355] ), .Y(new_n7464_));
  AOI22X1  g06462(.A0(new_n7464_), .A1(new_n7460_), .B0(new_n7463_), .B1(new_n7462_), .Y(new_n7465_));
  INVX1    g06463(.A(\A[360] ), .Y(new_n7466_));
  INVX1    g06464(.A(\A[359] ), .Y(new_n7467_));
  OR2X1    g06465(.A(new_n7467_), .B(\A[358] ), .Y(new_n7468_));
  AOI21X1  g06466(.A0(new_n7467_), .A1(\A[358] ), .B0(new_n7466_), .Y(new_n7469_));
  XOR2X1   g06467(.A(\A[359] ), .B(\A[358] ), .Y(new_n7470_));
  AOI22X1  g06468(.A0(new_n7470_), .A1(new_n7466_), .B0(new_n7469_), .B1(new_n7468_), .Y(new_n7471_));
  OR2X1    g06469(.A(new_n7471_), .B(new_n7465_), .Y(new_n7472_));
  AND2X1   g06470(.A(\A[359] ), .B(\A[358] ), .Y(new_n7473_));
  AND2X1   g06471(.A(new_n7470_), .B(\A[360] ), .Y(new_n7474_));
  OR2X1    g06472(.A(new_n7474_), .B(new_n7473_), .Y(new_n7475_));
  AND2X1   g06473(.A(\A[356] ), .B(\A[355] ), .Y(new_n7476_));
  AOI21X1  g06474(.A0(new_n7464_), .A1(\A[357] ), .B0(new_n7476_), .Y(new_n7477_));
  XOR2X1   g06475(.A(new_n7477_), .B(new_n7475_), .Y(new_n7478_));
  XOR2X1   g06476(.A(new_n7478_), .B(new_n7472_), .Y(new_n7479_));
  INVX1    g06477(.A(\A[355] ), .Y(new_n7480_));
  AND2X1   g06478(.A(\A[356] ), .B(new_n7480_), .Y(new_n7481_));
  OAI21X1  g06479(.A0(\A[356] ), .A1(new_n7480_), .B0(\A[357] ), .Y(new_n7482_));
  NAND2X1  g06480(.A(new_n7464_), .B(new_n7460_), .Y(new_n7483_));
  OAI21X1  g06481(.A0(new_n7482_), .A1(new_n7481_), .B0(new_n7483_), .Y(new_n7484_));
  XOR2X1   g06482(.A(new_n7471_), .B(new_n7484_), .Y(new_n7485_));
  NOR2X1   g06483(.A(new_n7471_), .B(new_n7465_), .Y(new_n7486_));
  AOI21X1  g06484(.A0(new_n7470_), .A1(\A[360] ), .B0(new_n7473_), .Y(new_n7487_));
  XOR2X1   g06485(.A(new_n7477_), .B(new_n7487_), .Y(new_n7488_));
  NOR2X1   g06486(.A(new_n7477_), .B(new_n7487_), .Y(new_n7489_));
  AOI21X1  g06487(.A0(new_n7488_), .A1(new_n7486_), .B0(new_n7489_), .Y(new_n7490_));
  OAI21X1  g06488(.A0(new_n7490_), .A1(new_n7485_), .B0(new_n7479_), .Y(new_n7491_));
  AND2X1   g06489(.A(\A[365] ), .B(\A[364] ), .Y(new_n7492_));
  XOR2X1   g06490(.A(\A[365] ), .B(\A[364] ), .Y(new_n7493_));
  AOI21X1  g06491(.A0(new_n7493_), .A1(\A[366] ), .B0(new_n7492_), .Y(new_n7494_));
  AND2X1   g06492(.A(\A[362] ), .B(\A[361] ), .Y(new_n7495_));
  XOR2X1   g06493(.A(\A[362] ), .B(\A[361] ), .Y(new_n7496_));
  AOI21X1  g06494(.A0(new_n7496_), .A1(\A[363] ), .B0(new_n7495_), .Y(new_n7497_));
  INVX1    g06495(.A(\A[363] ), .Y(new_n7498_));
  INVX1    g06496(.A(\A[362] ), .Y(new_n7499_));
  OR2X1    g06497(.A(new_n7499_), .B(\A[361] ), .Y(new_n7500_));
  AOI21X1  g06498(.A0(new_n7499_), .A1(\A[361] ), .B0(new_n7498_), .Y(new_n7501_));
  AOI22X1  g06499(.A0(new_n7501_), .A1(new_n7500_), .B0(new_n7496_), .B1(new_n7498_), .Y(new_n7502_));
  INVX1    g06500(.A(\A[366] ), .Y(new_n7503_));
  INVX1    g06501(.A(\A[365] ), .Y(new_n7504_));
  OR2X1    g06502(.A(new_n7504_), .B(\A[364] ), .Y(new_n7505_));
  AOI21X1  g06503(.A0(new_n7504_), .A1(\A[364] ), .B0(new_n7503_), .Y(new_n7506_));
  AOI22X1  g06504(.A0(new_n7506_), .A1(new_n7505_), .B0(new_n7493_), .B1(new_n7503_), .Y(new_n7507_));
  NOR4X1   g06505(.A(new_n7507_), .B(new_n7502_), .C(new_n7497_), .D(new_n7494_), .Y(new_n7508_));
  NOR4X1   g06506(.A(new_n7477_), .B(new_n7487_), .C(new_n7471_), .D(new_n7465_), .Y(new_n7509_));
  INVX1    g06507(.A(\A[361] ), .Y(new_n7510_));
  AND2X1   g06508(.A(\A[362] ), .B(new_n7510_), .Y(new_n7511_));
  OAI21X1  g06509(.A0(\A[362] ), .A1(new_n7510_), .B0(\A[363] ), .Y(new_n7512_));
  NAND2X1  g06510(.A(new_n7496_), .B(new_n7498_), .Y(new_n7513_));
  OAI21X1  g06511(.A0(new_n7512_), .A1(new_n7511_), .B0(new_n7513_), .Y(new_n7514_));
  XOR2X1   g06512(.A(new_n7507_), .B(new_n7514_), .Y(new_n7515_));
  OR4X1    g06513(.A(new_n7515_), .B(new_n7509_), .C(new_n7508_), .D(new_n7485_), .Y(new_n7516_));
  XOR2X1   g06514(.A(new_n7497_), .B(new_n7494_), .Y(new_n7517_));
  NOR2X1   g06515(.A(new_n7507_), .B(new_n7502_), .Y(new_n7518_));
  NOR2X1   g06516(.A(new_n7497_), .B(new_n7494_), .Y(new_n7519_));
  AOI21X1  g06517(.A0(new_n7518_), .A1(new_n7517_), .B0(new_n7519_), .Y(new_n7520_));
  XOR2X1   g06518(.A(new_n7518_), .B(new_n7517_), .Y(new_n7521_));
  OAI21X1  g06519(.A0(new_n7515_), .A1(new_n7520_), .B0(new_n7521_), .Y(new_n7522_));
  XOR2X1   g06520(.A(new_n7522_), .B(new_n7516_), .Y(new_n7523_));
  AND2X1   g06521(.A(new_n7523_), .B(new_n7491_), .Y(new_n7524_));
  OR2X1    g06522(.A(new_n7515_), .B(new_n7508_), .Y(new_n7525_));
  XOR2X1   g06523(.A(new_n7471_), .B(new_n7465_), .Y(new_n7526_));
  XOR2X1   g06524(.A(new_n7526_), .B(new_n7525_), .Y(new_n7527_));
  OR2X1    g06525(.A(new_n7438_), .B(new_n7431_), .Y(new_n7528_));
  XOR2X1   g06526(.A(new_n7394_), .B(new_n7388_), .Y(new_n7529_));
  XOR2X1   g06527(.A(new_n7529_), .B(new_n7528_), .Y(new_n7530_));
  NOR2X1   g06528(.A(new_n7530_), .B(new_n7527_), .Y(new_n7531_));
  AND2X1   g06529(.A(new_n7493_), .B(\A[366] ), .Y(new_n7532_));
  OR2X1    g06530(.A(new_n7532_), .B(new_n7492_), .Y(new_n7533_));
  XOR2X1   g06531(.A(new_n7497_), .B(new_n7533_), .Y(new_n7534_));
  XOR2X1   g06532(.A(new_n7518_), .B(new_n7534_), .Y(new_n7535_));
  NOR4X1   g06533(.A(new_n7515_), .B(new_n7509_), .C(new_n7535_), .D(new_n7485_), .Y(new_n7536_));
  OR2X1    g06534(.A(new_n7507_), .B(new_n7502_), .Y(new_n7537_));
  OR2X1    g06535(.A(new_n7497_), .B(new_n7494_), .Y(new_n7538_));
  OAI21X1  g06536(.A0(new_n7537_), .A1(new_n7534_), .B0(new_n7538_), .Y(new_n7539_));
  XOR2X1   g06537(.A(new_n7507_), .B(new_n7502_), .Y(new_n7540_));
  OAI21X1  g06538(.A0(new_n7540_), .A1(new_n7521_), .B0(new_n7539_), .Y(new_n7541_));
  AOI22X1  g06539(.A0(new_n7541_), .A1(new_n7536_), .B0(new_n7522_), .B1(new_n7516_), .Y(new_n7542_));
  OAI21X1  g06540(.A0(new_n7542_), .A1(new_n7491_), .B0(new_n7531_), .Y(new_n7543_));
  AOI21X1  g06541(.A0(new_n7540_), .A1(new_n7539_), .B0(new_n7535_), .Y(new_n7544_));
  XOR2X1   g06542(.A(new_n7544_), .B(new_n7516_), .Y(new_n7545_));
  MX2X1    g06543(.A(new_n7542_), .B(new_n7545_), .S0(new_n7491_), .Y(new_n7546_));
  OAI22X1  g06544(.A0(new_n7546_), .A1(new_n7531_), .B0(new_n7543_), .B1(new_n7524_), .Y(new_n7547_));
  AND2X1   g06545(.A(new_n7547_), .B(new_n7459_), .Y(new_n7548_));
  XOR2X1   g06546(.A(new_n7471_), .B(new_n7484_), .Y(new_n7549_));
  XOR2X1   g06547(.A(new_n7549_), .B(new_n7525_), .Y(new_n7550_));
  XOR2X1   g06548(.A(new_n7530_), .B(new_n7550_), .Y(new_n7551_));
  INVX1    g06549(.A(new_n7317_), .Y(new_n7552_));
  XOR2X1   g06550(.A(new_n7552_), .B(new_n7281_), .Y(new_n7553_));
  NOR2X1   g06551(.A(new_n7553_), .B(new_n7551_), .Y(new_n7554_));
  NAND2X1  g06552(.A(new_n7523_), .B(new_n7491_), .Y(new_n7555_));
  NOR4X1   g06553(.A(new_n7515_), .B(new_n7509_), .C(new_n7508_), .D(new_n7485_), .Y(new_n7556_));
  OR4X1    g06554(.A(new_n7515_), .B(new_n7509_), .C(new_n7535_), .D(new_n7485_), .Y(new_n7557_));
  AOI21X1  g06555(.A0(new_n7515_), .A1(new_n7535_), .B0(new_n7520_), .Y(new_n7558_));
  OAI22X1  g06556(.A0(new_n7558_), .A1(new_n7557_), .B0(new_n7544_), .B1(new_n7556_), .Y(new_n7559_));
  MX2X1    g06557(.A(new_n7559_), .B(new_n7523_), .S0(new_n7491_), .Y(new_n7560_));
  XOR2X1   g06558(.A(new_n7478_), .B(new_n7486_), .Y(new_n7561_));
  XOR2X1   g06559(.A(new_n7471_), .B(new_n7465_), .Y(new_n7562_));
  OR2X1    g06560(.A(new_n7477_), .B(new_n7487_), .Y(new_n7563_));
  OAI21X1  g06561(.A0(new_n7478_), .A1(new_n7472_), .B0(new_n7563_), .Y(new_n7564_));
  AOI21X1  g06562(.A0(new_n7564_), .A1(new_n7562_), .B0(new_n7561_), .Y(new_n7565_));
  AOI21X1  g06563(.A0(new_n7559_), .A1(new_n7565_), .B0(new_n7531_), .Y(new_n7566_));
  AOI22X1  g06564(.A0(new_n7566_), .A1(new_n7555_), .B0(new_n7560_), .B1(new_n7531_), .Y(new_n7567_));
  OAI21X1  g06565(.A0(new_n7567_), .A1(new_n7459_), .B0(new_n7554_), .Y(new_n7568_));
  NOR4X1   g06566(.A(new_n7438_), .B(new_n7432_), .C(new_n7431_), .D(new_n7408_), .Y(new_n7569_));
  XOR2X1   g06567(.A(new_n7449_), .B(new_n7569_), .Y(new_n7570_));
  OR4X1    g06568(.A(new_n7438_), .B(new_n7432_), .C(new_n7447_), .D(new_n7408_), .Y(new_n7571_));
  AOI21X1  g06569(.A0(new_n7438_), .A1(new_n7447_), .B0(new_n7453_), .Y(new_n7572_));
  OAI22X1  g06570(.A0(new_n7572_), .A1(new_n7571_), .B0(new_n7449_), .B1(new_n7569_), .Y(new_n7573_));
  MX2X1    g06571(.A(new_n7573_), .B(new_n7570_), .S0(new_n7414_), .Y(new_n7574_));
  OR2X1    g06572(.A(new_n7530_), .B(new_n7527_), .Y(new_n7575_));
  AOI21X1  g06573(.A0(new_n7559_), .A1(new_n7565_), .B0(new_n7575_), .Y(new_n7576_));
  AOI22X1  g06574(.A0(new_n7560_), .A1(new_n7575_), .B0(new_n7576_), .B1(new_n7555_), .Y(new_n7577_));
  MX2X1    g06575(.A(new_n7577_), .B(new_n7567_), .S0(new_n7574_), .Y(new_n7578_));
  OAI22X1  g06576(.A0(new_n7578_), .A1(new_n7554_), .B0(new_n7568_), .B1(new_n7548_), .Y(new_n7579_));
  AND2X1   g06577(.A(new_n7579_), .B(new_n7382_), .Y(new_n7580_));
  XOR2X1   g06578(.A(new_n7553_), .B(new_n7551_), .Y(new_n7581_));
  INVX1    g06579(.A(new_n7581_), .Y(new_n7582_));
  INVX1    g06580(.A(\A[314] ), .Y(new_n7583_));
  AND2X1   g06581(.A(new_n7583_), .B(\A[313] ), .Y(new_n7584_));
  OAI21X1  g06582(.A0(new_n7583_), .A1(\A[313] ), .B0(\A[315] ), .Y(new_n7585_));
  INVX1    g06583(.A(\A[315] ), .Y(new_n7586_));
  XOR2X1   g06584(.A(\A[314] ), .B(\A[313] ), .Y(new_n7587_));
  NAND2X1  g06585(.A(new_n7587_), .B(new_n7586_), .Y(new_n7588_));
  OAI21X1  g06586(.A0(new_n7585_), .A1(new_n7584_), .B0(new_n7588_), .Y(new_n7589_));
  INVX1    g06587(.A(\A[318] ), .Y(new_n7590_));
  INVX1    g06588(.A(\A[316] ), .Y(new_n7591_));
  OR2X1    g06589(.A(\A[317] ), .B(new_n7591_), .Y(new_n7592_));
  AOI21X1  g06590(.A0(\A[317] ), .A1(new_n7591_), .B0(new_n7590_), .Y(new_n7593_));
  XOR2X1   g06591(.A(\A[317] ), .B(\A[316] ), .Y(new_n7594_));
  AOI22X1  g06592(.A0(new_n7594_), .A1(new_n7590_), .B0(new_n7593_), .B1(new_n7592_), .Y(new_n7595_));
  AND2X1   g06593(.A(\A[317] ), .B(\A[316] ), .Y(new_n7596_));
  AOI21X1  g06594(.A0(new_n7594_), .A1(\A[318] ), .B0(new_n7596_), .Y(new_n7597_));
  AND2X1   g06595(.A(\A[314] ), .B(\A[313] ), .Y(new_n7598_));
  AOI21X1  g06596(.A0(new_n7587_), .A1(\A[315] ), .B0(new_n7598_), .Y(new_n7599_));
  XOR2X1   g06597(.A(new_n7595_), .B(new_n7589_), .Y(new_n7600_));
  INVX1    g06598(.A(\A[309] ), .Y(new_n7601_));
  INVX1    g06599(.A(\A[307] ), .Y(new_n7602_));
  OR2X1    g06600(.A(\A[308] ), .B(new_n7602_), .Y(new_n7603_));
  AOI21X1  g06601(.A0(\A[308] ), .A1(new_n7602_), .B0(new_n7601_), .Y(new_n7604_));
  XOR2X1   g06602(.A(\A[308] ), .B(\A[307] ), .Y(new_n7605_));
  AOI22X1  g06603(.A0(new_n7605_), .A1(new_n7601_), .B0(new_n7604_), .B1(new_n7603_), .Y(new_n7606_));
  INVX1    g06604(.A(\A[312] ), .Y(new_n7607_));
  INVX1    g06605(.A(\A[310] ), .Y(new_n7608_));
  OR2X1    g06606(.A(\A[311] ), .B(new_n7608_), .Y(new_n7609_));
  AOI21X1  g06607(.A0(\A[311] ), .A1(new_n7608_), .B0(new_n7607_), .Y(new_n7610_));
  XOR2X1   g06608(.A(\A[311] ), .B(\A[310] ), .Y(new_n7611_));
  AOI22X1  g06609(.A0(new_n7611_), .A1(new_n7607_), .B0(new_n7610_), .B1(new_n7609_), .Y(new_n7612_));
  AND2X1   g06610(.A(\A[311] ), .B(\A[310] ), .Y(new_n7613_));
  AOI21X1  g06611(.A0(new_n7611_), .A1(\A[312] ), .B0(new_n7613_), .Y(new_n7614_));
  AND2X1   g06612(.A(\A[308] ), .B(\A[307] ), .Y(new_n7615_));
  AOI21X1  g06613(.A0(new_n7605_), .A1(\A[309] ), .B0(new_n7615_), .Y(new_n7616_));
  XOR2X1   g06614(.A(new_n7612_), .B(new_n7606_), .Y(new_n7617_));
  XOR2X1   g06615(.A(new_n7617_), .B(new_n7600_), .Y(new_n7618_));
  INVX1    g06616(.A(\A[302] ), .Y(new_n7619_));
  AND2X1   g06617(.A(new_n7619_), .B(\A[301] ), .Y(new_n7620_));
  OAI21X1  g06618(.A0(new_n7619_), .A1(\A[301] ), .B0(\A[303] ), .Y(new_n7621_));
  INVX1    g06619(.A(\A[303] ), .Y(new_n7622_));
  XOR2X1   g06620(.A(\A[302] ), .B(\A[301] ), .Y(new_n7623_));
  NAND2X1  g06621(.A(new_n7623_), .B(new_n7622_), .Y(new_n7624_));
  OAI21X1  g06622(.A0(new_n7621_), .A1(new_n7620_), .B0(new_n7624_), .Y(new_n7625_));
  INVX1    g06623(.A(\A[306] ), .Y(new_n7626_));
  INVX1    g06624(.A(\A[304] ), .Y(new_n7627_));
  OR2X1    g06625(.A(\A[305] ), .B(new_n7627_), .Y(new_n7628_));
  AOI21X1  g06626(.A0(\A[305] ), .A1(new_n7627_), .B0(new_n7626_), .Y(new_n7629_));
  XOR2X1   g06627(.A(\A[305] ), .B(\A[304] ), .Y(new_n7630_));
  AOI22X1  g06628(.A0(new_n7630_), .A1(new_n7626_), .B0(new_n7629_), .B1(new_n7628_), .Y(new_n7631_));
  AND2X1   g06629(.A(\A[305] ), .B(\A[304] ), .Y(new_n7632_));
  AOI21X1  g06630(.A0(new_n7630_), .A1(\A[306] ), .B0(new_n7632_), .Y(new_n7633_));
  AND2X1   g06631(.A(\A[302] ), .B(\A[301] ), .Y(new_n7634_));
  AOI21X1  g06632(.A0(new_n7623_), .A1(\A[303] ), .B0(new_n7634_), .Y(new_n7635_));
  XOR2X1   g06633(.A(new_n7631_), .B(new_n7625_), .Y(new_n7636_));
  INVX1    g06634(.A(\A[297] ), .Y(new_n7637_));
  INVX1    g06635(.A(\A[295] ), .Y(new_n7638_));
  OR2X1    g06636(.A(\A[296] ), .B(new_n7638_), .Y(new_n7639_));
  AOI21X1  g06637(.A0(\A[296] ), .A1(new_n7638_), .B0(new_n7637_), .Y(new_n7640_));
  XOR2X1   g06638(.A(\A[296] ), .B(\A[295] ), .Y(new_n7641_));
  AOI22X1  g06639(.A0(new_n7641_), .A1(new_n7637_), .B0(new_n7640_), .B1(new_n7639_), .Y(new_n7642_));
  INVX1    g06640(.A(\A[300] ), .Y(new_n7643_));
  INVX1    g06641(.A(\A[298] ), .Y(new_n7644_));
  OR2X1    g06642(.A(\A[299] ), .B(new_n7644_), .Y(new_n7645_));
  AOI21X1  g06643(.A0(\A[299] ), .A1(new_n7644_), .B0(new_n7643_), .Y(new_n7646_));
  XOR2X1   g06644(.A(\A[299] ), .B(\A[298] ), .Y(new_n7647_));
  AOI22X1  g06645(.A0(new_n7647_), .A1(new_n7643_), .B0(new_n7646_), .B1(new_n7645_), .Y(new_n7648_));
  AND2X1   g06646(.A(\A[299] ), .B(\A[298] ), .Y(new_n7649_));
  AOI21X1  g06647(.A0(new_n7647_), .A1(\A[300] ), .B0(new_n7649_), .Y(new_n7650_));
  AND2X1   g06648(.A(\A[296] ), .B(\A[295] ), .Y(new_n7651_));
  AOI21X1  g06649(.A0(new_n7641_), .A1(\A[297] ), .B0(new_n7651_), .Y(new_n7652_));
  XOR2X1   g06650(.A(new_n7648_), .B(new_n7642_), .Y(new_n7653_));
  XOR2X1   g06651(.A(new_n7653_), .B(new_n7636_), .Y(new_n7654_));
  XOR2X1   g06652(.A(new_n7654_), .B(new_n7618_), .Y(new_n7655_));
  INVX1    g06653(.A(\A[290] ), .Y(new_n7656_));
  AND2X1   g06654(.A(new_n7656_), .B(\A[289] ), .Y(new_n7657_));
  OAI21X1  g06655(.A0(new_n7656_), .A1(\A[289] ), .B0(\A[291] ), .Y(new_n7658_));
  INVX1    g06656(.A(\A[291] ), .Y(new_n7659_));
  XOR2X1   g06657(.A(\A[290] ), .B(\A[289] ), .Y(new_n7660_));
  NAND2X1  g06658(.A(new_n7660_), .B(new_n7659_), .Y(new_n7661_));
  OAI21X1  g06659(.A0(new_n7658_), .A1(new_n7657_), .B0(new_n7661_), .Y(new_n7662_));
  INVX1    g06660(.A(\A[294] ), .Y(new_n7663_));
  INVX1    g06661(.A(\A[292] ), .Y(new_n7664_));
  OR2X1    g06662(.A(\A[293] ), .B(new_n7664_), .Y(new_n7665_));
  AOI21X1  g06663(.A0(\A[293] ), .A1(new_n7664_), .B0(new_n7663_), .Y(new_n7666_));
  XOR2X1   g06664(.A(\A[293] ), .B(\A[292] ), .Y(new_n7667_));
  AOI22X1  g06665(.A0(new_n7667_), .A1(new_n7663_), .B0(new_n7666_), .B1(new_n7665_), .Y(new_n7668_));
  AND2X1   g06666(.A(\A[293] ), .B(\A[292] ), .Y(new_n7669_));
  AOI21X1  g06667(.A0(new_n7667_), .A1(\A[294] ), .B0(new_n7669_), .Y(new_n7670_));
  AND2X1   g06668(.A(\A[290] ), .B(\A[289] ), .Y(new_n7671_));
  AOI21X1  g06669(.A0(new_n7660_), .A1(\A[291] ), .B0(new_n7671_), .Y(new_n7672_));
  XOR2X1   g06670(.A(new_n7668_), .B(new_n7662_), .Y(new_n7673_));
  INVX1    g06671(.A(\A[285] ), .Y(new_n7674_));
  INVX1    g06672(.A(\A[283] ), .Y(new_n7675_));
  OR2X1    g06673(.A(\A[284] ), .B(new_n7675_), .Y(new_n7676_));
  AOI21X1  g06674(.A0(\A[284] ), .A1(new_n7675_), .B0(new_n7674_), .Y(new_n7677_));
  XOR2X1   g06675(.A(\A[284] ), .B(\A[283] ), .Y(new_n7678_));
  AOI22X1  g06676(.A0(new_n7678_), .A1(new_n7674_), .B0(new_n7677_), .B1(new_n7676_), .Y(new_n7679_));
  INVX1    g06677(.A(\A[288] ), .Y(new_n7680_));
  INVX1    g06678(.A(\A[286] ), .Y(new_n7681_));
  OR2X1    g06679(.A(\A[287] ), .B(new_n7681_), .Y(new_n7682_));
  AOI21X1  g06680(.A0(\A[287] ), .A1(new_n7681_), .B0(new_n7680_), .Y(new_n7683_));
  XOR2X1   g06681(.A(\A[287] ), .B(\A[286] ), .Y(new_n7684_));
  AOI22X1  g06682(.A0(new_n7684_), .A1(new_n7680_), .B0(new_n7683_), .B1(new_n7682_), .Y(new_n7685_));
  AND2X1   g06683(.A(\A[287] ), .B(\A[286] ), .Y(new_n7686_));
  AOI21X1  g06684(.A0(new_n7684_), .A1(\A[288] ), .B0(new_n7686_), .Y(new_n7687_));
  AND2X1   g06685(.A(\A[284] ), .B(\A[283] ), .Y(new_n7688_));
  AOI21X1  g06686(.A0(new_n7678_), .A1(\A[285] ), .B0(new_n7688_), .Y(new_n7689_));
  XOR2X1   g06687(.A(new_n7685_), .B(new_n7679_), .Y(new_n7690_));
  XOR2X1   g06688(.A(new_n7690_), .B(new_n7673_), .Y(new_n7691_));
  INVX1    g06689(.A(new_n7691_), .Y(new_n7692_));
  INVX1    g06690(.A(\A[278] ), .Y(new_n7693_));
  AND2X1   g06691(.A(new_n7693_), .B(\A[277] ), .Y(new_n7694_));
  OAI21X1  g06692(.A0(new_n7693_), .A1(\A[277] ), .B0(\A[279] ), .Y(new_n7695_));
  INVX1    g06693(.A(\A[279] ), .Y(new_n7696_));
  XOR2X1   g06694(.A(\A[278] ), .B(\A[277] ), .Y(new_n7697_));
  NAND2X1  g06695(.A(new_n7697_), .B(new_n7696_), .Y(new_n7698_));
  OAI21X1  g06696(.A0(new_n7695_), .A1(new_n7694_), .B0(new_n7698_), .Y(new_n7699_));
  INVX1    g06697(.A(\A[282] ), .Y(new_n7700_));
  INVX1    g06698(.A(\A[280] ), .Y(new_n7701_));
  OR2X1    g06699(.A(\A[281] ), .B(new_n7701_), .Y(new_n7702_));
  AOI21X1  g06700(.A0(\A[281] ), .A1(new_n7701_), .B0(new_n7700_), .Y(new_n7703_));
  XOR2X1   g06701(.A(\A[281] ), .B(\A[280] ), .Y(new_n7704_));
  AOI22X1  g06702(.A0(new_n7704_), .A1(new_n7700_), .B0(new_n7703_), .B1(new_n7702_), .Y(new_n7705_));
  AND2X1   g06703(.A(\A[281] ), .B(\A[280] ), .Y(new_n7706_));
  AOI21X1  g06704(.A0(new_n7704_), .A1(\A[282] ), .B0(new_n7706_), .Y(new_n7707_));
  AND2X1   g06705(.A(\A[278] ), .B(\A[277] ), .Y(new_n7708_));
  AOI21X1  g06706(.A0(new_n7697_), .A1(\A[279] ), .B0(new_n7708_), .Y(new_n7709_));
  XOR2X1   g06707(.A(new_n7705_), .B(new_n7699_), .Y(new_n7710_));
  INVX1    g06708(.A(\A[273] ), .Y(new_n7711_));
  INVX1    g06709(.A(\A[271] ), .Y(new_n7712_));
  OR2X1    g06710(.A(\A[272] ), .B(new_n7712_), .Y(new_n7713_));
  AOI21X1  g06711(.A0(\A[272] ), .A1(new_n7712_), .B0(new_n7711_), .Y(new_n7714_));
  XOR2X1   g06712(.A(\A[272] ), .B(\A[271] ), .Y(new_n7715_));
  AOI22X1  g06713(.A0(new_n7715_), .A1(new_n7711_), .B0(new_n7714_), .B1(new_n7713_), .Y(new_n7716_));
  INVX1    g06714(.A(\A[276] ), .Y(new_n7717_));
  INVX1    g06715(.A(\A[274] ), .Y(new_n7718_));
  OR2X1    g06716(.A(\A[275] ), .B(new_n7718_), .Y(new_n7719_));
  AOI21X1  g06717(.A0(\A[275] ), .A1(new_n7718_), .B0(new_n7717_), .Y(new_n7720_));
  XOR2X1   g06718(.A(\A[275] ), .B(\A[274] ), .Y(new_n7721_));
  AOI22X1  g06719(.A0(new_n7721_), .A1(new_n7717_), .B0(new_n7720_), .B1(new_n7719_), .Y(new_n7722_));
  AND2X1   g06720(.A(\A[275] ), .B(\A[274] ), .Y(new_n7723_));
  AOI21X1  g06721(.A0(new_n7721_), .A1(\A[276] ), .B0(new_n7723_), .Y(new_n7724_));
  AND2X1   g06722(.A(\A[272] ), .B(\A[271] ), .Y(new_n7725_));
  AOI21X1  g06723(.A0(new_n7715_), .A1(\A[273] ), .B0(new_n7725_), .Y(new_n7726_));
  XOR2X1   g06724(.A(new_n7722_), .B(new_n7716_), .Y(new_n7727_));
  XOR2X1   g06725(.A(new_n7727_), .B(new_n7710_), .Y(new_n7728_));
  XOR2X1   g06726(.A(new_n7728_), .B(new_n7692_), .Y(new_n7729_));
  XOR2X1   g06727(.A(new_n7729_), .B(new_n7655_), .Y(new_n7730_));
  NOR2X1   g06728(.A(new_n7730_), .B(new_n7582_), .Y(new_n7731_));
  OR2X1    g06729(.A(new_n7577_), .B(new_n7574_), .Y(new_n7732_));
  OAI21X1  g06730(.A0(new_n7542_), .A1(new_n7491_), .B0(new_n7575_), .Y(new_n7733_));
  OAI22X1  g06731(.A0(new_n7733_), .A1(new_n7524_), .B0(new_n7546_), .B1(new_n7575_), .Y(new_n7734_));
  MX2X1    g06732(.A(new_n7547_), .B(new_n7734_), .S0(new_n7574_), .Y(new_n7735_));
  AOI21X1  g06733(.A0(new_n7734_), .A1(new_n7574_), .B0(new_n7554_), .Y(new_n7736_));
  AOI22X1  g06734(.A0(new_n7736_), .A1(new_n7732_), .B0(new_n7735_), .B1(new_n7554_), .Y(new_n7737_));
  OAI21X1  g06735(.A0(new_n7737_), .A1(new_n7382_), .B0(new_n7731_), .Y(new_n7738_));
  OR2X1    g06736(.A(new_n7553_), .B(new_n7551_), .Y(new_n7739_));
  AOI21X1  g06737(.A0(new_n7734_), .A1(new_n7574_), .B0(new_n7739_), .Y(new_n7740_));
  AOI22X1  g06738(.A0(new_n7735_), .A1(new_n7739_), .B0(new_n7740_), .B1(new_n7732_), .Y(new_n7741_));
  MX2X1    g06739(.A(new_n7737_), .B(new_n7741_), .S0(new_n7382_), .Y(new_n7742_));
  OAI22X1  g06740(.A0(new_n7742_), .A1(new_n7731_), .B0(new_n7738_), .B1(new_n7580_), .Y(new_n7743_));
  INVX1    g06741(.A(\A[296] ), .Y(new_n7744_));
  AND2X1   g06742(.A(new_n7744_), .B(\A[295] ), .Y(new_n7745_));
  OAI21X1  g06743(.A0(new_n7744_), .A1(\A[295] ), .B0(\A[297] ), .Y(new_n7746_));
  NAND2X1  g06744(.A(new_n7641_), .B(new_n7637_), .Y(new_n7747_));
  OAI21X1  g06745(.A0(new_n7746_), .A1(new_n7745_), .B0(new_n7747_), .Y(new_n7748_));
  XOR2X1   g06746(.A(new_n7648_), .B(new_n7748_), .Y(new_n7749_));
  XOR2X1   g06747(.A(new_n7652_), .B(new_n7650_), .Y(new_n7750_));
  NOR2X1   g06748(.A(new_n7648_), .B(new_n7642_), .Y(new_n7751_));
  NOR2X1   g06749(.A(new_n7652_), .B(new_n7650_), .Y(new_n7752_));
  AOI21X1  g06750(.A0(new_n7751_), .A1(new_n7750_), .B0(new_n7752_), .Y(new_n7753_));
  XOR2X1   g06751(.A(new_n7751_), .B(new_n7750_), .Y(new_n7754_));
  OAI21X1  g06752(.A0(new_n7753_), .A1(new_n7749_), .B0(new_n7754_), .Y(new_n7755_));
  XOR2X1   g06753(.A(new_n7631_), .B(new_n7625_), .Y(new_n7756_));
  INVX1    g06754(.A(\A[301] ), .Y(new_n7757_));
  OR2X1    g06755(.A(\A[302] ), .B(new_n7757_), .Y(new_n7758_));
  AOI21X1  g06756(.A0(\A[302] ), .A1(new_n7757_), .B0(new_n7622_), .Y(new_n7759_));
  AOI22X1  g06757(.A0(new_n7623_), .A1(new_n7622_), .B0(new_n7759_), .B1(new_n7758_), .Y(new_n7760_));
  NOR4X1   g06758(.A(new_n7635_), .B(new_n7633_), .C(new_n7631_), .D(new_n7760_), .Y(new_n7761_));
  NOR4X1   g06759(.A(new_n7652_), .B(new_n7650_), .C(new_n7648_), .D(new_n7642_), .Y(new_n7762_));
  NOR4X1   g06760(.A(new_n7762_), .B(new_n7749_), .C(new_n7761_), .D(new_n7756_), .Y(new_n7763_));
  XOR2X1   g06761(.A(new_n7631_), .B(new_n7760_), .Y(new_n7764_));
  AND2X1   g06762(.A(new_n7630_), .B(\A[306] ), .Y(new_n7765_));
  OR2X1    g06763(.A(new_n7765_), .B(new_n7632_), .Y(new_n7766_));
  XOR2X1   g06764(.A(new_n7635_), .B(new_n7766_), .Y(new_n7767_));
  OR2X1    g06765(.A(new_n7631_), .B(new_n7760_), .Y(new_n7768_));
  OR2X1    g06766(.A(new_n7635_), .B(new_n7633_), .Y(new_n7769_));
  OAI21X1  g06767(.A0(new_n7768_), .A1(new_n7767_), .B0(new_n7769_), .Y(new_n7770_));
  NOR2X1   g06768(.A(new_n7631_), .B(new_n7760_), .Y(new_n7771_));
  XOR2X1   g06769(.A(new_n7771_), .B(new_n7767_), .Y(new_n7772_));
  AOI21X1  g06770(.A0(new_n7770_), .A1(new_n7764_), .B0(new_n7772_), .Y(new_n7773_));
  XOR2X1   g06771(.A(new_n7773_), .B(new_n7763_), .Y(new_n7774_));
  OR4X1    g06772(.A(new_n7749_), .B(new_n7761_), .C(new_n7772_), .D(new_n7756_), .Y(new_n7775_));
  XOR2X1   g06773(.A(new_n7635_), .B(new_n7633_), .Y(new_n7776_));
  NOR2X1   g06774(.A(new_n7635_), .B(new_n7633_), .Y(new_n7777_));
  AOI21X1  g06775(.A0(new_n7771_), .A1(new_n7776_), .B0(new_n7777_), .Y(new_n7778_));
  AND2X1   g06776(.A(new_n7647_), .B(\A[300] ), .Y(new_n7779_));
  OR2X1    g06777(.A(new_n7779_), .B(new_n7649_), .Y(new_n7780_));
  XOR2X1   g06778(.A(new_n7652_), .B(new_n7780_), .Y(new_n7781_));
  XOR2X1   g06779(.A(new_n7751_), .B(new_n7781_), .Y(new_n7782_));
  OAI22X1  g06780(.A0(new_n7782_), .A1(new_n7753_), .B0(new_n7778_), .B1(new_n7756_), .Y(new_n7783_));
  OAI22X1  g06781(.A0(new_n7783_), .A1(new_n7775_), .B0(new_n7773_), .B1(new_n7763_), .Y(new_n7784_));
  MX2X1    g06782(.A(new_n7784_), .B(new_n7774_), .S0(new_n7755_), .Y(new_n7785_));
  INVX1    g06783(.A(\A[308] ), .Y(new_n7786_));
  AND2X1   g06784(.A(new_n7786_), .B(\A[307] ), .Y(new_n7787_));
  OAI21X1  g06785(.A0(new_n7786_), .A1(\A[307] ), .B0(\A[309] ), .Y(new_n7788_));
  NAND2X1  g06786(.A(new_n7605_), .B(new_n7601_), .Y(new_n7789_));
  OAI21X1  g06787(.A0(new_n7788_), .A1(new_n7787_), .B0(new_n7789_), .Y(new_n7790_));
  XOR2X1   g06788(.A(new_n7612_), .B(new_n7790_), .Y(new_n7791_));
  XOR2X1   g06789(.A(new_n7616_), .B(new_n7614_), .Y(new_n7792_));
  NOR2X1   g06790(.A(new_n7612_), .B(new_n7606_), .Y(new_n7793_));
  NOR2X1   g06791(.A(new_n7616_), .B(new_n7614_), .Y(new_n7794_));
  AOI21X1  g06792(.A0(new_n7793_), .A1(new_n7792_), .B0(new_n7794_), .Y(new_n7795_));
  XOR2X1   g06793(.A(new_n7793_), .B(new_n7792_), .Y(new_n7796_));
  OAI21X1  g06794(.A0(new_n7795_), .A1(new_n7791_), .B0(new_n7796_), .Y(new_n7797_));
  XOR2X1   g06795(.A(new_n7595_), .B(new_n7589_), .Y(new_n7798_));
  INVX1    g06796(.A(\A[313] ), .Y(new_n7799_));
  OR2X1    g06797(.A(\A[314] ), .B(new_n7799_), .Y(new_n7800_));
  AOI21X1  g06798(.A0(\A[314] ), .A1(new_n7799_), .B0(new_n7586_), .Y(new_n7801_));
  AOI22X1  g06799(.A0(new_n7587_), .A1(new_n7586_), .B0(new_n7801_), .B1(new_n7800_), .Y(new_n7802_));
  NOR4X1   g06800(.A(new_n7599_), .B(new_n7597_), .C(new_n7595_), .D(new_n7802_), .Y(new_n7803_));
  NOR4X1   g06801(.A(new_n7616_), .B(new_n7614_), .C(new_n7612_), .D(new_n7606_), .Y(new_n7804_));
  OR4X1    g06802(.A(new_n7804_), .B(new_n7791_), .C(new_n7803_), .D(new_n7798_), .Y(new_n7805_));
  XOR2X1   g06803(.A(new_n7599_), .B(new_n7597_), .Y(new_n7806_));
  NOR2X1   g06804(.A(new_n7595_), .B(new_n7802_), .Y(new_n7807_));
  NOR2X1   g06805(.A(new_n7599_), .B(new_n7597_), .Y(new_n7808_));
  AOI21X1  g06806(.A0(new_n7807_), .A1(new_n7806_), .B0(new_n7808_), .Y(new_n7809_));
  XOR2X1   g06807(.A(new_n7807_), .B(new_n7806_), .Y(new_n7810_));
  OAI21X1  g06808(.A0(new_n7809_), .A1(new_n7798_), .B0(new_n7810_), .Y(new_n7811_));
  XOR2X1   g06809(.A(new_n7811_), .B(new_n7805_), .Y(new_n7812_));
  NAND2X1  g06810(.A(new_n7812_), .B(new_n7797_), .Y(new_n7813_));
  OR2X1    g06811(.A(new_n7654_), .B(new_n7618_), .Y(new_n7814_));
  XOR2X1   g06812(.A(new_n7612_), .B(new_n7606_), .Y(new_n7815_));
  AND2X1   g06813(.A(new_n7611_), .B(\A[312] ), .Y(new_n7816_));
  OR2X1    g06814(.A(new_n7816_), .B(new_n7613_), .Y(new_n7817_));
  XOR2X1   g06815(.A(new_n7616_), .B(new_n7817_), .Y(new_n7818_));
  OR2X1    g06816(.A(new_n7612_), .B(new_n7606_), .Y(new_n7819_));
  OR2X1    g06817(.A(new_n7616_), .B(new_n7614_), .Y(new_n7820_));
  OAI21X1  g06818(.A0(new_n7819_), .A1(new_n7818_), .B0(new_n7820_), .Y(new_n7821_));
  XOR2X1   g06819(.A(new_n7793_), .B(new_n7818_), .Y(new_n7822_));
  AOI21X1  g06820(.A0(new_n7821_), .A1(new_n7815_), .B0(new_n7822_), .Y(new_n7823_));
  NOR4X1   g06821(.A(new_n7804_), .B(new_n7791_), .C(new_n7803_), .D(new_n7798_), .Y(new_n7824_));
  XOR2X1   g06822(.A(new_n7595_), .B(new_n7802_), .Y(new_n7825_));
  AND2X1   g06823(.A(new_n7594_), .B(\A[318] ), .Y(new_n7826_));
  OR2X1    g06824(.A(new_n7826_), .B(new_n7596_), .Y(new_n7827_));
  XOR2X1   g06825(.A(new_n7599_), .B(new_n7827_), .Y(new_n7828_));
  OR2X1    g06826(.A(new_n7595_), .B(new_n7802_), .Y(new_n7829_));
  OR2X1    g06827(.A(new_n7599_), .B(new_n7597_), .Y(new_n7830_));
  OAI21X1  g06828(.A0(new_n7829_), .A1(new_n7828_), .B0(new_n7830_), .Y(new_n7831_));
  XOR2X1   g06829(.A(new_n7829_), .B(new_n7806_), .Y(new_n7832_));
  AOI21X1  g06830(.A0(new_n7831_), .A1(new_n7825_), .B0(new_n7832_), .Y(new_n7833_));
  OR4X1    g06831(.A(new_n7791_), .B(new_n7803_), .C(new_n7832_), .D(new_n7798_), .Y(new_n7834_));
  OAI22X1  g06832(.A0(new_n7822_), .A1(new_n7795_), .B0(new_n7809_), .B1(new_n7798_), .Y(new_n7835_));
  OAI22X1  g06833(.A0(new_n7835_), .A1(new_n7834_), .B0(new_n7833_), .B1(new_n7824_), .Y(new_n7836_));
  AOI21X1  g06834(.A0(new_n7836_), .A1(new_n7823_), .B0(new_n7814_), .Y(new_n7837_));
  MX2X1    g06835(.A(new_n7836_), .B(new_n7812_), .S0(new_n7797_), .Y(new_n7838_));
  AOI22X1  g06836(.A0(new_n7838_), .A1(new_n7814_), .B0(new_n7837_), .B1(new_n7813_), .Y(new_n7839_));
  OR2X1    g06837(.A(new_n7839_), .B(new_n7785_), .Y(new_n7840_));
  INVX1    g06838(.A(new_n7655_), .Y(new_n7841_));
  OR2X1    g06839(.A(new_n7729_), .B(new_n7841_), .Y(new_n7842_));
  AND2X1   g06840(.A(new_n7812_), .B(new_n7797_), .Y(new_n7843_));
  XOR2X1   g06841(.A(new_n7833_), .B(new_n7805_), .Y(new_n7844_));
  NOR4X1   g06842(.A(new_n7791_), .B(new_n7832_), .C(new_n7831_), .D(new_n7798_), .Y(new_n7845_));
  AOI21X1  g06843(.A0(new_n7831_), .A1(new_n7825_), .B0(new_n7804_), .Y(new_n7846_));
  AOI22X1  g06844(.A0(new_n7846_), .A1(new_n7845_), .B0(new_n7811_), .B1(new_n7805_), .Y(new_n7847_));
  MX2X1    g06845(.A(new_n7847_), .B(new_n7844_), .S0(new_n7797_), .Y(new_n7848_));
  OAI21X1  g06846(.A0(new_n7847_), .A1(new_n7797_), .B0(new_n7814_), .Y(new_n7849_));
  OAI22X1  g06847(.A0(new_n7849_), .A1(new_n7843_), .B0(new_n7848_), .B1(new_n7814_), .Y(new_n7850_));
  AOI21X1  g06848(.A0(new_n7850_), .A1(new_n7785_), .B0(new_n7842_), .Y(new_n7851_));
  OR4X1    g06849(.A(new_n7762_), .B(new_n7749_), .C(new_n7761_), .D(new_n7756_), .Y(new_n7852_));
  XOR2X1   g06850(.A(new_n7773_), .B(new_n7852_), .Y(new_n7853_));
  XOR2X1   g06851(.A(new_n7771_), .B(new_n7776_), .Y(new_n7854_));
  OAI21X1  g06852(.A0(new_n7778_), .A1(new_n7756_), .B0(new_n7854_), .Y(new_n7855_));
  NOR4X1   g06853(.A(new_n7749_), .B(new_n7772_), .C(new_n7770_), .D(new_n7756_), .Y(new_n7856_));
  AOI21X1  g06854(.A0(new_n7770_), .A1(new_n7764_), .B0(new_n7762_), .Y(new_n7857_));
  AOI22X1  g06855(.A0(new_n7857_), .A1(new_n7856_), .B0(new_n7855_), .B1(new_n7852_), .Y(new_n7858_));
  MX2X1    g06856(.A(new_n7858_), .B(new_n7853_), .S0(new_n7755_), .Y(new_n7859_));
  NOR2X1   g06857(.A(new_n7654_), .B(new_n7618_), .Y(new_n7860_));
  OAI21X1  g06858(.A0(new_n7847_), .A1(new_n7797_), .B0(new_n7860_), .Y(new_n7861_));
  OAI22X1  g06859(.A0(new_n7848_), .A1(new_n7860_), .B0(new_n7861_), .B1(new_n7843_), .Y(new_n7862_));
  MX2X1    g06860(.A(new_n7850_), .B(new_n7862_), .S0(new_n7859_), .Y(new_n7863_));
  AOI22X1  g06861(.A0(new_n7863_), .A1(new_n7842_), .B0(new_n7851_), .B1(new_n7840_), .Y(new_n7864_));
  INVX1    g06862(.A(\A[284] ), .Y(new_n7865_));
  AND2X1   g06863(.A(new_n7865_), .B(\A[283] ), .Y(new_n7866_));
  OAI21X1  g06864(.A0(new_n7865_), .A1(\A[283] ), .B0(\A[285] ), .Y(new_n7867_));
  NAND2X1  g06865(.A(new_n7678_), .B(new_n7674_), .Y(new_n7868_));
  OAI21X1  g06866(.A0(new_n7867_), .A1(new_n7866_), .B0(new_n7868_), .Y(new_n7869_));
  XOR2X1   g06867(.A(new_n7685_), .B(new_n7869_), .Y(new_n7870_));
  XOR2X1   g06868(.A(new_n7689_), .B(new_n7687_), .Y(new_n7871_));
  NOR2X1   g06869(.A(new_n7685_), .B(new_n7679_), .Y(new_n7872_));
  NOR2X1   g06870(.A(new_n7689_), .B(new_n7687_), .Y(new_n7873_));
  AOI21X1  g06871(.A0(new_n7872_), .A1(new_n7871_), .B0(new_n7873_), .Y(new_n7874_));
  XOR2X1   g06872(.A(new_n7872_), .B(new_n7871_), .Y(new_n7875_));
  OAI21X1  g06873(.A0(new_n7874_), .A1(new_n7870_), .B0(new_n7875_), .Y(new_n7876_));
  XOR2X1   g06874(.A(new_n7668_), .B(new_n7662_), .Y(new_n7877_));
  INVX1    g06875(.A(\A[289] ), .Y(new_n7878_));
  OR2X1    g06876(.A(\A[290] ), .B(new_n7878_), .Y(new_n7879_));
  AOI21X1  g06877(.A0(\A[290] ), .A1(new_n7878_), .B0(new_n7659_), .Y(new_n7880_));
  AOI22X1  g06878(.A0(new_n7660_), .A1(new_n7659_), .B0(new_n7880_), .B1(new_n7879_), .Y(new_n7881_));
  NOR4X1   g06879(.A(new_n7672_), .B(new_n7670_), .C(new_n7668_), .D(new_n7881_), .Y(new_n7882_));
  NOR4X1   g06880(.A(new_n7689_), .B(new_n7687_), .C(new_n7685_), .D(new_n7679_), .Y(new_n7883_));
  OR4X1    g06881(.A(new_n7883_), .B(new_n7870_), .C(new_n7882_), .D(new_n7877_), .Y(new_n7884_));
  XOR2X1   g06882(.A(new_n7672_), .B(new_n7670_), .Y(new_n7885_));
  NOR2X1   g06883(.A(new_n7668_), .B(new_n7881_), .Y(new_n7886_));
  NOR2X1   g06884(.A(new_n7672_), .B(new_n7670_), .Y(new_n7887_));
  AOI21X1  g06885(.A0(new_n7886_), .A1(new_n7885_), .B0(new_n7887_), .Y(new_n7888_));
  XOR2X1   g06886(.A(new_n7886_), .B(new_n7885_), .Y(new_n7889_));
  OAI21X1  g06887(.A0(new_n7888_), .A1(new_n7877_), .B0(new_n7889_), .Y(new_n7890_));
  XOR2X1   g06888(.A(new_n7890_), .B(new_n7884_), .Y(new_n7891_));
  NAND2X1  g06889(.A(new_n7891_), .B(new_n7876_), .Y(new_n7892_));
  OR2X1    g06890(.A(new_n7728_), .B(new_n7691_), .Y(new_n7893_));
  XOR2X1   g06891(.A(new_n7685_), .B(new_n7679_), .Y(new_n7894_));
  AND2X1   g06892(.A(new_n7684_), .B(\A[288] ), .Y(new_n7895_));
  OR2X1    g06893(.A(new_n7895_), .B(new_n7686_), .Y(new_n7896_));
  XOR2X1   g06894(.A(new_n7689_), .B(new_n7896_), .Y(new_n7897_));
  OR2X1    g06895(.A(new_n7685_), .B(new_n7679_), .Y(new_n7898_));
  OR2X1    g06896(.A(new_n7689_), .B(new_n7687_), .Y(new_n7899_));
  OAI21X1  g06897(.A0(new_n7898_), .A1(new_n7897_), .B0(new_n7899_), .Y(new_n7900_));
  XOR2X1   g06898(.A(new_n7872_), .B(new_n7897_), .Y(new_n7901_));
  AOI21X1  g06899(.A0(new_n7900_), .A1(new_n7894_), .B0(new_n7901_), .Y(new_n7902_));
  NOR4X1   g06900(.A(new_n7883_), .B(new_n7870_), .C(new_n7882_), .D(new_n7877_), .Y(new_n7903_));
  XOR2X1   g06901(.A(new_n7668_), .B(new_n7881_), .Y(new_n7904_));
  AND2X1   g06902(.A(new_n7667_), .B(\A[294] ), .Y(new_n7905_));
  OR2X1    g06903(.A(new_n7905_), .B(new_n7669_), .Y(new_n7906_));
  XOR2X1   g06904(.A(new_n7672_), .B(new_n7906_), .Y(new_n7907_));
  OR2X1    g06905(.A(new_n7668_), .B(new_n7881_), .Y(new_n7908_));
  OR2X1    g06906(.A(new_n7672_), .B(new_n7670_), .Y(new_n7909_));
  OAI21X1  g06907(.A0(new_n7908_), .A1(new_n7907_), .B0(new_n7909_), .Y(new_n7910_));
  XOR2X1   g06908(.A(new_n7908_), .B(new_n7885_), .Y(new_n7911_));
  AOI21X1  g06909(.A0(new_n7910_), .A1(new_n7904_), .B0(new_n7911_), .Y(new_n7912_));
  OR4X1    g06910(.A(new_n7870_), .B(new_n7882_), .C(new_n7911_), .D(new_n7877_), .Y(new_n7913_));
  OAI22X1  g06911(.A0(new_n7901_), .A1(new_n7874_), .B0(new_n7888_), .B1(new_n7877_), .Y(new_n7914_));
  OAI22X1  g06912(.A0(new_n7914_), .A1(new_n7913_), .B0(new_n7912_), .B1(new_n7903_), .Y(new_n7915_));
  AOI21X1  g06913(.A0(new_n7915_), .A1(new_n7902_), .B0(new_n7893_), .Y(new_n7916_));
  MX2X1    g06914(.A(new_n7915_), .B(new_n7891_), .S0(new_n7876_), .Y(new_n7917_));
  AOI22X1  g06915(.A0(new_n7917_), .A1(new_n7893_), .B0(new_n7916_), .B1(new_n7892_), .Y(new_n7918_));
  INVX1    g06916(.A(\A[272] ), .Y(new_n7919_));
  AND2X1   g06917(.A(new_n7919_), .B(\A[271] ), .Y(new_n7920_));
  OAI21X1  g06918(.A0(new_n7919_), .A1(\A[271] ), .B0(\A[273] ), .Y(new_n7921_));
  NAND2X1  g06919(.A(new_n7715_), .B(new_n7711_), .Y(new_n7922_));
  OAI21X1  g06920(.A0(new_n7921_), .A1(new_n7920_), .B0(new_n7922_), .Y(new_n7923_));
  XOR2X1   g06921(.A(new_n7722_), .B(new_n7923_), .Y(new_n7924_));
  XOR2X1   g06922(.A(new_n7726_), .B(new_n7724_), .Y(new_n7925_));
  NOR2X1   g06923(.A(new_n7722_), .B(new_n7716_), .Y(new_n7926_));
  NOR2X1   g06924(.A(new_n7726_), .B(new_n7724_), .Y(new_n7927_));
  AOI21X1  g06925(.A0(new_n7926_), .A1(new_n7925_), .B0(new_n7927_), .Y(new_n7928_));
  XOR2X1   g06926(.A(new_n7926_), .B(new_n7925_), .Y(new_n7929_));
  OAI21X1  g06927(.A0(new_n7928_), .A1(new_n7924_), .B0(new_n7929_), .Y(new_n7930_));
  XOR2X1   g06928(.A(new_n7705_), .B(new_n7699_), .Y(new_n7931_));
  INVX1    g06929(.A(\A[277] ), .Y(new_n7932_));
  OR2X1    g06930(.A(\A[278] ), .B(new_n7932_), .Y(new_n7933_));
  AOI21X1  g06931(.A0(\A[278] ), .A1(new_n7932_), .B0(new_n7696_), .Y(new_n7934_));
  AOI22X1  g06932(.A0(new_n7697_), .A1(new_n7696_), .B0(new_n7934_), .B1(new_n7933_), .Y(new_n7935_));
  NOR4X1   g06933(.A(new_n7709_), .B(new_n7707_), .C(new_n7705_), .D(new_n7935_), .Y(new_n7936_));
  NOR4X1   g06934(.A(new_n7726_), .B(new_n7724_), .C(new_n7722_), .D(new_n7716_), .Y(new_n7937_));
  OR4X1    g06935(.A(new_n7937_), .B(new_n7924_), .C(new_n7936_), .D(new_n7931_), .Y(new_n7938_));
  XOR2X1   g06936(.A(new_n7705_), .B(new_n7935_), .Y(new_n7939_));
  AND2X1   g06937(.A(new_n7704_), .B(\A[282] ), .Y(new_n7940_));
  OR2X1    g06938(.A(new_n7940_), .B(new_n7706_), .Y(new_n7941_));
  XOR2X1   g06939(.A(new_n7709_), .B(new_n7941_), .Y(new_n7942_));
  OR2X1    g06940(.A(new_n7705_), .B(new_n7935_), .Y(new_n7943_));
  OR2X1    g06941(.A(new_n7709_), .B(new_n7707_), .Y(new_n7944_));
  OAI21X1  g06942(.A0(new_n7943_), .A1(new_n7942_), .B0(new_n7944_), .Y(new_n7945_));
  NOR2X1   g06943(.A(new_n7705_), .B(new_n7935_), .Y(new_n7946_));
  XOR2X1   g06944(.A(new_n7946_), .B(new_n7942_), .Y(new_n7947_));
  AOI21X1  g06945(.A0(new_n7945_), .A1(new_n7939_), .B0(new_n7947_), .Y(new_n7948_));
  XOR2X1   g06946(.A(new_n7948_), .B(new_n7938_), .Y(new_n7949_));
  XOR2X1   g06947(.A(new_n7709_), .B(new_n7707_), .Y(new_n7950_));
  NOR2X1   g06948(.A(new_n7709_), .B(new_n7707_), .Y(new_n7951_));
  AOI21X1  g06949(.A0(new_n7946_), .A1(new_n7950_), .B0(new_n7951_), .Y(new_n7952_));
  XOR2X1   g06950(.A(new_n7946_), .B(new_n7950_), .Y(new_n7953_));
  OAI21X1  g06951(.A0(new_n7952_), .A1(new_n7931_), .B0(new_n7953_), .Y(new_n7954_));
  NOR4X1   g06952(.A(new_n7924_), .B(new_n7947_), .C(new_n7945_), .D(new_n7931_), .Y(new_n7955_));
  AOI21X1  g06953(.A0(new_n7945_), .A1(new_n7939_), .B0(new_n7937_), .Y(new_n7956_));
  AOI22X1  g06954(.A0(new_n7956_), .A1(new_n7955_), .B0(new_n7954_), .B1(new_n7938_), .Y(new_n7957_));
  MX2X1    g06955(.A(new_n7957_), .B(new_n7949_), .S0(new_n7930_), .Y(new_n7958_));
  NOR2X1   g06956(.A(new_n7728_), .B(new_n7691_), .Y(new_n7959_));
  AOI21X1  g06957(.A0(new_n7915_), .A1(new_n7902_), .B0(new_n7959_), .Y(new_n7960_));
  AOI22X1  g06958(.A0(new_n7960_), .A1(new_n7892_), .B0(new_n7917_), .B1(new_n7959_), .Y(new_n7961_));
  MX2X1    g06959(.A(new_n7961_), .B(new_n7918_), .S0(new_n7958_), .Y(new_n7962_));
  NOR2X1   g06960(.A(new_n7729_), .B(new_n7841_), .Y(new_n7963_));
  AOI21X1  g06961(.A0(new_n7850_), .A1(new_n7785_), .B0(new_n7963_), .Y(new_n7964_));
  AOI22X1  g06962(.A0(new_n7964_), .A1(new_n7840_), .B0(new_n7863_), .B1(new_n7963_), .Y(new_n7965_));
  MX2X1    g06963(.A(new_n7965_), .B(new_n7864_), .S0(new_n7962_), .Y(new_n7966_));
  OR2X1    g06964(.A(new_n7730_), .B(new_n7582_), .Y(new_n7967_));
  OAI21X1  g06965(.A0(new_n7737_), .A1(new_n7382_), .B0(new_n7967_), .Y(new_n7968_));
  OAI22X1  g06966(.A0(new_n7968_), .A1(new_n7580_), .B0(new_n7742_), .B1(new_n7967_), .Y(new_n7969_));
  MX2X1    g06967(.A(new_n7969_), .B(new_n7743_), .S0(new_n7966_), .Y(new_n7970_));
  INVX1    g06968(.A(\A[393] ), .Y(new_n7971_));
  INVX1    g06969(.A(\A[392] ), .Y(new_n7972_));
  OR2X1    g06970(.A(new_n7972_), .B(\A[391] ), .Y(new_n7973_));
  AOI21X1  g06971(.A0(new_n7972_), .A1(\A[391] ), .B0(new_n7971_), .Y(new_n7974_));
  XOR2X1   g06972(.A(\A[392] ), .B(\A[391] ), .Y(new_n7975_));
  AOI22X1  g06973(.A0(new_n7975_), .A1(new_n7971_), .B0(new_n7974_), .B1(new_n7973_), .Y(new_n7976_));
  INVX1    g06974(.A(\A[396] ), .Y(new_n7977_));
  INVX1    g06975(.A(\A[395] ), .Y(new_n7978_));
  OR2X1    g06976(.A(new_n7978_), .B(\A[394] ), .Y(new_n7979_));
  AOI21X1  g06977(.A0(new_n7978_), .A1(\A[394] ), .B0(new_n7977_), .Y(new_n7980_));
  XOR2X1   g06978(.A(\A[395] ), .B(\A[394] ), .Y(new_n7981_));
  AOI22X1  g06979(.A0(new_n7981_), .A1(new_n7977_), .B0(new_n7980_), .B1(new_n7979_), .Y(new_n7982_));
  OR2X1    g06980(.A(new_n7982_), .B(new_n7976_), .Y(new_n7983_));
  AND2X1   g06981(.A(\A[395] ), .B(\A[394] ), .Y(new_n7984_));
  AND2X1   g06982(.A(new_n7981_), .B(\A[396] ), .Y(new_n7985_));
  OR2X1    g06983(.A(new_n7985_), .B(new_n7984_), .Y(new_n7986_));
  AND2X1   g06984(.A(\A[392] ), .B(\A[391] ), .Y(new_n7987_));
  AOI21X1  g06985(.A0(new_n7975_), .A1(\A[393] ), .B0(new_n7987_), .Y(new_n7988_));
  XOR2X1   g06986(.A(new_n7988_), .B(new_n7986_), .Y(new_n7989_));
  XOR2X1   g06987(.A(new_n7989_), .B(new_n7983_), .Y(new_n7990_));
  INVX1    g06988(.A(\A[391] ), .Y(new_n7991_));
  AND2X1   g06989(.A(\A[392] ), .B(new_n7991_), .Y(new_n7992_));
  OAI21X1  g06990(.A0(\A[392] ), .A1(new_n7991_), .B0(\A[393] ), .Y(new_n7993_));
  NAND2X1  g06991(.A(new_n7975_), .B(new_n7971_), .Y(new_n7994_));
  OAI21X1  g06992(.A0(new_n7993_), .A1(new_n7992_), .B0(new_n7994_), .Y(new_n7995_));
  XOR2X1   g06993(.A(new_n7982_), .B(new_n7995_), .Y(new_n7996_));
  NOR2X1   g06994(.A(new_n7982_), .B(new_n7976_), .Y(new_n7997_));
  AOI21X1  g06995(.A0(new_n7981_), .A1(\A[396] ), .B0(new_n7984_), .Y(new_n7998_));
  XOR2X1   g06996(.A(new_n7988_), .B(new_n7998_), .Y(new_n7999_));
  NOR2X1   g06997(.A(new_n7988_), .B(new_n7998_), .Y(new_n8000_));
  AOI21X1  g06998(.A0(new_n7999_), .A1(new_n7997_), .B0(new_n8000_), .Y(new_n8001_));
  OAI21X1  g06999(.A0(new_n8001_), .A1(new_n7996_), .B0(new_n7990_), .Y(new_n8002_));
  AND2X1   g07000(.A(\A[401] ), .B(\A[400] ), .Y(new_n8003_));
  XOR2X1   g07001(.A(\A[401] ), .B(\A[400] ), .Y(new_n8004_));
  AOI21X1  g07002(.A0(new_n8004_), .A1(\A[402] ), .B0(new_n8003_), .Y(new_n8005_));
  AND2X1   g07003(.A(\A[398] ), .B(\A[397] ), .Y(new_n8006_));
  XOR2X1   g07004(.A(\A[398] ), .B(\A[397] ), .Y(new_n8007_));
  AOI21X1  g07005(.A0(new_n8007_), .A1(\A[399] ), .B0(new_n8006_), .Y(new_n8008_));
  INVX1    g07006(.A(\A[399] ), .Y(new_n8009_));
  INVX1    g07007(.A(\A[398] ), .Y(new_n8010_));
  OR2X1    g07008(.A(new_n8010_), .B(\A[397] ), .Y(new_n8011_));
  AOI21X1  g07009(.A0(new_n8010_), .A1(\A[397] ), .B0(new_n8009_), .Y(new_n8012_));
  AOI22X1  g07010(.A0(new_n8012_), .A1(new_n8011_), .B0(new_n8007_), .B1(new_n8009_), .Y(new_n8013_));
  INVX1    g07011(.A(\A[402] ), .Y(new_n8014_));
  INVX1    g07012(.A(\A[401] ), .Y(new_n8015_));
  OR2X1    g07013(.A(new_n8015_), .B(\A[400] ), .Y(new_n8016_));
  AOI21X1  g07014(.A0(new_n8015_), .A1(\A[400] ), .B0(new_n8014_), .Y(new_n8017_));
  AOI22X1  g07015(.A0(new_n8017_), .A1(new_n8016_), .B0(new_n8004_), .B1(new_n8014_), .Y(new_n8018_));
  NOR4X1   g07016(.A(new_n8018_), .B(new_n8013_), .C(new_n8008_), .D(new_n8005_), .Y(new_n8019_));
  NOR4X1   g07017(.A(new_n7988_), .B(new_n7998_), .C(new_n7982_), .D(new_n7976_), .Y(new_n8020_));
  INVX1    g07018(.A(\A[397] ), .Y(new_n8021_));
  AND2X1   g07019(.A(\A[398] ), .B(new_n8021_), .Y(new_n8022_));
  OAI21X1  g07020(.A0(\A[398] ), .A1(new_n8021_), .B0(\A[399] ), .Y(new_n8023_));
  NAND2X1  g07021(.A(new_n8007_), .B(new_n8009_), .Y(new_n8024_));
  OAI21X1  g07022(.A0(new_n8023_), .A1(new_n8022_), .B0(new_n8024_), .Y(new_n8025_));
  XOR2X1   g07023(.A(new_n8018_), .B(new_n8025_), .Y(new_n8026_));
  NOR4X1   g07024(.A(new_n8026_), .B(new_n8020_), .C(new_n8019_), .D(new_n7996_), .Y(new_n8027_));
  AND2X1   g07025(.A(new_n8004_), .B(\A[402] ), .Y(new_n8028_));
  OR2X1    g07026(.A(new_n8028_), .B(new_n8003_), .Y(new_n8029_));
  XOR2X1   g07027(.A(new_n8008_), .B(new_n8029_), .Y(new_n8030_));
  OR2X1    g07028(.A(new_n8018_), .B(new_n8013_), .Y(new_n8031_));
  OR2X1    g07029(.A(new_n8008_), .B(new_n8005_), .Y(new_n8032_));
  OAI21X1  g07030(.A0(new_n8031_), .A1(new_n8030_), .B0(new_n8032_), .Y(new_n8033_));
  NOR2X1   g07031(.A(new_n8018_), .B(new_n8013_), .Y(new_n8034_));
  XOR2X1   g07032(.A(new_n8034_), .B(new_n8030_), .Y(new_n8035_));
  XOR2X1   g07033(.A(new_n8018_), .B(new_n8013_), .Y(new_n8036_));
  AOI21X1  g07034(.A0(new_n8036_), .A1(new_n8033_), .B0(new_n8035_), .Y(new_n8037_));
  XOR2X1   g07035(.A(new_n8037_), .B(new_n8027_), .Y(new_n8038_));
  OR4X1    g07036(.A(new_n8026_), .B(new_n8020_), .C(new_n8035_), .D(new_n7996_), .Y(new_n8039_));
  XOR2X1   g07037(.A(new_n8008_), .B(new_n8005_), .Y(new_n8040_));
  NOR2X1   g07038(.A(new_n8008_), .B(new_n8005_), .Y(new_n8041_));
  AOI21X1  g07039(.A0(new_n8034_), .A1(new_n8040_), .B0(new_n8041_), .Y(new_n8042_));
  AOI21X1  g07040(.A0(new_n8026_), .A1(new_n8035_), .B0(new_n8042_), .Y(new_n8043_));
  OAI22X1  g07041(.A0(new_n8043_), .A1(new_n8039_), .B0(new_n8037_), .B1(new_n8027_), .Y(new_n8044_));
  MX2X1    g07042(.A(new_n8044_), .B(new_n8038_), .S0(new_n8002_), .Y(new_n8045_));
  INVX1    g07043(.A(\A[405] ), .Y(new_n8046_));
  INVX1    g07044(.A(\A[404] ), .Y(new_n8047_));
  OR2X1    g07045(.A(new_n8047_), .B(\A[403] ), .Y(new_n8048_));
  AOI21X1  g07046(.A0(new_n8047_), .A1(\A[403] ), .B0(new_n8046_), .Y(new_n8049_));
  XOR2X1   g07047(.A(\A[404] ), .B(\A[403] ), .Y(new_n8050_));
  AOI22X1  g07048(.A0(new_n8050_), .A1(new_n8046_), .B0(new_n8049_), .B1(new_n8048_), .Y(new_n8051_));
  INVX1    g07049(.A(\A[408] ), .Y(new_n8052_));
  INVX1    g07050(.A(\A[407] ), .Y(new_n8053_));
  OR2X1    g07051(.A(new_n8053_), .B(\A[406] ), .Y(new_n8054_));
  AOI21X1  g07052(.A0(new_n8053_), .A1(\A[406] ), .B0(new_n8052_), .Y(new_n8055_));
  XOR2X1   g07053(.A(\A[407] ), .B(\A[406] ), .Y(new_n8056_));
  AOI22X1  g07054(.A0(new_n8056_), .A1(new_n8052_), .B0(new_n8055_), .B1(new_n8054_), .Y(new_n8057_));
  OR2X1    g07055(.A(new_n8057_), .B(new_n8051_), .Y(new_n8058_));
  AND2X1   g07056(.A(\A[407] ), .B(\A[406] ), .Y(new_n8059_));
  AND2X1   g07057(.A(new_n8056_), .B(\A[408] ), .Y(new_n8060_));
  OR2X1    g07058(.A(new_n8060_), .B(new_n8059_), .Y(new_n8061_));
  AND2X1   g07059(.A(\A[404] ), .B(\A[403] ), .Y(new_n8062_));
  AOI21X1  g07060(.A0(new_n8050_), .A1(\A[405] ), .B0(new_n8062_), .Y(new_n8063_));
  XOR2X1   g07061(.A(new_n8063_), .B(new_n8061_), .Y(new_n8064_));
  XOR2X1   g07062(.A(new_n8064_), .B(new_n8058_), .Y(new_n8065_));
  INVX1    g07063(.A(\A[403] ), .Y(new_n8066_));
  AND2X1   g07064(.A(\A[404] ), .B(new_n8066_), .Y(new_n8067_));
  OAI21X1  g07065(.A0(\A[404] ), .A1(new_n8066_), .B0(\A[405] ), .Y(new_n8068_));
  NAND2X1  g07066(.A(new_n8050_), .B(new_n8046_), .Y(new_n8069_));
  OAI21X1  g07067(.A0(new_n8068_), .A1(new_n8067_), .B0(new_n8069_), .Y(new_n8070_));
  XOR2X1   g07068(.A(new_n8057_), .B(new_n8070_), .Y(new_n8071_));
  NOR2X1   g07069(.A(new_n8057_), .B(new_n8051_), .Y(new_n8072_));
  AOI21X1  g07070(.A0(new_n8056_), .A1(\A[408] ), .B0(new_n8059_), .Y(new_n8073_));
  XOR2X1   g07071(.A(new_n8063_), .B(new_n8073_), .Y(new_n8074_));
  NOR2X1   g07072(.A(new_n8063_), .B(new_n8073_), .Y(new_n8075_));
  AOI21X1  g07073(.A0(new_n8074_), .A1(new_n8072_), .B0(new_n8075_), .Y(new_n8076_));
  OAI21X1  g07074(.A0(new_n8076_), .A1(new_n8071_), .B0(new_n8065_), .Y(new_n8077_));
  AND2X1   g07075(.A(\A[413] ), .B(\A[412] ), .Y(new_n8078_));
  XOR2X1   g07076(.A(\A[413] ), .B(\A[412] ), .Y(new_n8079_));
  AOI21X1  g07077(.A0(new_n8079_), .A1(\A[414] ), .B0(new_n8078_), .Y(new_n8080_));
  AND2X1   g07078(.A(\A[410] ), .B(\A[409] ), .Y(new_n8081_));
  XOR2X1   g07079(.A(\A[410] ), .B(\A[409] ), .Y(new_n8082_));
  AOI21X1  g07080(.A0(new_n8082_), .A1(\A[411] ), .B0(new_n8081_), .Y(new_n8083_));
  INVX1    g07081(.A(\A[411] ), .Y(new_n8084_));
  INVX1    g07082(.A(\A[410] ), .Y(new_n8085_));
  OR2X1    g07083(.A(new_n8085_), .B(\A[409] ), .Y(new_n8086_));
  AOI21X1  g07084(.A0(new_n8085_), .A1(\A[409] ), .B0(new_n8084_), .Y(new_n8087_));
  AOI22X1  g07085(.A0(new_n8087_), .A1(new_n8086_), .B0(new_n8082_), .B1(new_n8084_), .Y(new_n8088_));
  INVX1    g07086(.A(\A[414] ), .Y(new_n8089_));
  INVX1    g07087(.A(\A[413] ), .Y(new_n8090_));
  OR2X1    g07088(.A(new_n8090_), .B(\A[412] ), .Y(new_n8091_));
  AOI21X1  g07089(.A0(new_n8090_), .A1(\A[412] ), .B0(new_n8089_), .Y(new_n8092_));
  AOI22X1  g07090(.A0(new_n8092_), .A1(new_n8091_), .B0(new_n8079_), .B1(new_n8089_), .Y(new_n8093_));
  NOR4X1   g07091(.A(new_n8093_), .B(new_n8088_), .C(new_n8083_), .D(new_n8080_), .Y(new_n8094_));
  NOR4X1   g07092(.A(new_n8063_), .B(new_n8073_), .C(new_n8057_), .D(new_n8051_), .Y(new_n8095_));
  INVX1    g07093(.A(\A[409] ), .Y(new_n8096_));
  AND2X1   g07094(.A(\A[410] ), .B(new_n8096_), .Y(new_n8097_));
  OAI21X1  g07095(.A0(\A[410] ), .A1(new_n8096_), .B0(\A[411] ), .Y(new_n8098_));
  NAND2X1  g07096(.A(new_n8082_), .B(new_n8084_), .Y(new_n8099_));
  OAI21X1  g07097(.A0(new_n8098_), .A1(new_n8097_), .B0(new_n8099_), .Y(new_n8100_));
  XOR2X1   g07098(.A(new_n8093_), .B(new_n8100_), .Y(new_n8101_));
  OR4X1    g07099(.A(new_n8101_), .B(new_n8095_), .C(new_n8094_), .D(new_n8071_), .Y(new_n8102_));
  XOR2X1   g07100(.A(new_n8083_), .B(new_n8080_), .Y(new_n8103_));
  NOR2X1   g07101(.A(new_n8093_), .B(new_n8088_), .Y(new_n8104_));
  NOR2X1   g07102(.A(new_n8083_), .B(new_n8080_), .Y(new_n8105_));
  AOI21X1  g07103(.A0(new_n8104_), .A1(new_n8103_), .B0(new_n8105_), .Y(new_n8106_));
  XOR2X1   g07104(.A(new_n8104_), .B(new_n8103_), .Y(new_n8107_));
  OAI21X1  g07105(.A0(new_n8101_), .A1(new_n8106_), .B0(new_n8107_), .Y(new_n8108_));
  XOR2X1   g07106(.A(new_n8108_), .B(new_n8102_), .Y(new_n8109_));
  NAND2X1  g07107(.A(new_n8109_), .B(new_n8077_), .Y(new_n8110_));
  OR2X1    g07108(.A(new_n8101_), .B(new_n8094_), .Y(new_n8111_));
  XOR2X1   g07109(.A(new_n8057_), .B(new_n8051_), .Y(new_n8112_));
  XOR2X1   g07110(.A(new_n8112_), .B(new_n8111_), .Y(new_n8113_));
  OR2X1    g07111(.A(new_n8026_), .B(new_n8019_), .Y(new_n8114_));
  XOR2X1   g07112(.A(new_n7982_), .B(new_n7976_), .Y(new_n8115_));
  XOR2X1   g07113(.A(new_n8115_), .B(new_n8114_), .Y(new_n8116_));
  OR2X1    g07114(.A(new_n8116_), .B(new_n8113_), .Y(new_n8117_));
  XOR2X1   g07115(.A(new_n8064_), .B(new_n8072_), .Y(new_n8118_));
  XOR2X1   g07116(.A(new_n8057_), .B(new_n8051_), .Y(new_n8119_));
  OR2X1    g07117(.A(new_n8063_), .B(new_n8073_), .Y(new_n8120_));
  OAI21X1  g07118(.A0(new_n8064_), .A1(new_n8058_), .B0(new_n8120_), .Y(new_n8121_));
  AOI21X1  g07119(.A0(new_n8121_), .A1(new_n8119_), .B0(new_n8118_), .Y(new_n8122_));
  NOR4X1   g07120(.A(new_n8101_), .B(new_n8095_), .C(new_n8094_), .D(new_n8071_), .Y(new_n8123_));
  AND2X1   g07121(.A(new_n8079_), .B(\A[414] ), .Y(new_n8124_));
  OR2X1    g07122(.A(new_n8124_), .B(new_n8078_), .Y(new_n8125_));
  XOR2X1   g07123(.A(new_n8083_), .B(new_n8125_), .Y(new_n8126_));
  OR2X1    g07124(.A(new_n8093_), .B(new_n8088_), .Y(new_n8127_));
  OR2X1    g07125(.A(new_n8083_), .B(new_n8080_), .Y(new_n8128_));
  OAI21X1  g07126(.A0(new_n8127_), .A1(new_n8126_), .B0(new_n8128_), .Y(new_n8129_));
  XOR2X1   g07127(.A(new_n8104_), .B(new_n8126_), .Y(new_n8130_));
  XOR2X1   g07128(.A(new_n8093_), .B(new_n8088_), .Y(new_n8131_));
  AOI21X1  g07129(.A0(new_n8131_), .A1(new_n8129_), .B0(new_n8130_), .Y(new_n8132_));
  OR4X1    g07130(.A(new_n8101_), .B(new_n8095_), .C(new_n8130_), .D(new_n8071_), .Y(new_n8133_));
  AOI21X1  g07131(.A0(new_n8101_), .A1(new_n8130_), .B0(new_n8106_), .Y(new_n8134_));
  OAI22X1  g07132(.A0(new_n8134_), .A1(new_n8133_), .B0(new_n8132_), .B1(new_n8123_), .Y(new_n8135_));
  AOI21X1  g07133(.A0(new_n8135_), .A1(new_n8122_), .B0(new_n8117_), .Y(new_n8136_));
  MX2X1    g07134(.A(new_n8135_), .B(new_n8109_), .S0(new_n8077_), .Y(new_n8137_));
  AOI22X1  g07135(.A0(new_n8137_), .A1(new_n8117_), .B0(new_n8136_), .B1(new_n8110_), .Y(new_n8138_));
  OR2X1    g07136(.A(new_n8138_), .B(new_n8045_), .Y(new_n8139_));
  XOR2X1   g07137(.A(new_n8057_), .B(new_n8070_), .Y(new_n8140_));
  XOR2X1   g07138(.A(new_n8140_), .B(new_n8111_), .Y(new_n8141_));
  XOR2X1   g07139(.A(new_n8116_), .B(new_n8141_), .Y(new_n8142_));
  INVX1    g07140(.A(\A[386] ), .Y(new_n8143_));
  AND2X1   g07141(.A(new_n8143_), .B(\A[385] ), .Y(new_n8144_));
  OAI21X1  g07142(.A0(new_n8143_), .A1(\A[385] ), .B0(\A[387] ), .Y(new_n8145_));
  INVX1    g07143(.A(\A[387] ), .Y(new_n8146_));
  XOR2X1   g07144(.A(\A[386] ), .B(\A[385] ), .Y(new_n8147_));
  NAND2X1  g07145(.A(new_n8147_), .B(new_n8146_), .Y(new_n8148_));
  OAI21X1  g07146(.A0(new_n8145_), .A1(new_n8144_), .B0(new_n8148_), .Y(new_n8149_));
  INVX1    g07147(.A(\A[390] ), .Y(new_n8150_));
  INVX1    g07148(.A(\A[388] ), .Y(new_n8151_));
  OR2X1    g07149(.A(\A[389] ), .B(new_n8151_), .Y(new_n8152_));
  AOI21X1  g07150(.A0(\A[389] ), .A1(new_n8151_), .B0(new_n8150_), .Y(new_n8153_));
  XOR2X1   g07151(.A(\A[389] ), .B(\A[388] ), .Y(new_n8154_));
  AOI22X1  g07152(.A0(new_n8154_), .A1(new_n8150_), .B0(new_n8153_), .B1(new_n8152_), .Y(new_n8155_));
  AND2X1   g07153(.A(\A[389] ), .B(\A[388] ), .Y(new_n8156_));
  AOI21X1  g07154(.A0(new_n8154_), .A1(\A[390] ), .B0(new_n8156_), .Y(new_n8157_));
  AND2X1   g07155(.A(\A[386] ), .B(\A[385] ), .Y(new_n8158_));
  AOI21X1  g07156(.A0(new_n8147_), .A1(\A[387] ), .B0(new_n8158_), .Y(new_n8159_));
  XOR2X1   g07157(.A(new_n8155_), .B(new_n8149_), .Y(new_n8160_));
  INVX1    g07158(.A(\A[381] ), .Y(new_n8161_));
  INVX1    g07159(.A(\A[379] ), .Y(new_n8162_));
  OR2X1    g07160(.A(\A[380] ), .B(new_n8162_), .Y(new_n8163_));
  AOI21X1  g07161(.A0(\A[380] ), .A1(new_n8162_), .B0(new_n8161_), .Y(new_n8164_));
  XOR2X1   g07162(.A(\A[380] ), .B(\A[379] ), .Y(new_n8165_));
  AOI22X1  g07163(.A0(new_n8165_), .A1(new_n8161_), .B0(new_n8164_), .B1(new_n8163_), .Y(new_n8166_));
  INVX1    g07164(.A(\A[384] ), .Y(new_n8167_));
  INVX1    g07165(.A(\A[382] ), .Y(new_n8168_));
  OR2X1    g07166(.A(\A[383] ), .B(new_n8168_), .Y(new_n8169_));
  AOI21X1  g07167(.A0(\A[383] ), .A1(new_n8168_), .B0(new_n8167_), .Y(new_n8170_));
  XOR2X1   g07168(.A(\A[383] ), .B(\A[382] ), .Y(new_n8171_));
  AOI22X1  g07169(.A0(new_n8171_), .A1(new_n8167_), .B0(new_n8170_), .B1(new_n8169_), .Y(new_n8172_));
  AND2X1   g07170(.A(\A[383] ), .B(\A[382] ), .Y(new_n8173_));
  AOI21X1  g07171(.A0(new_n8171_), .A1(\A[384] ), .B0(new_n8173_), .Y(new_n8174_));
  AND2X1   g07172(.A(\A[380] ), .B(\A[379] ), .Y(new_n8175_));
  AOI21X1  g07173(.A0(new_n8165_), .A1(\A[381] ), .B0(new_n8175_), .Y(new_n8176_));
  XOR2X1   g07174(.A(new_n8172_), .B(new_n8166_), .Y(new_n8177_));
  XOR2X1   g07175(.A(new_n8177_), .B(new_n8160_), .Y(new_n8178_));
  INVX1    g07176(.A(new_n8178_), .Y(new_n8179_));
  INVX1    g07177(.A(\A[374] ), .Y(new_n8180_));
  AND2X1   g07178(.A(new_n8180_), .B(\A[373] ), .Y(new_n8181_));
  OAI21X1  g07179(.A0(new_n8180_), .A1(\A[373] ), .B0(\A[375] ), .Y(new_n8182_));
  INVX1    g07180(.A(\A[375] ), .Y(new_n8183_));
  XOR2X1   g07181(.A(\A[374] ), .B(\A[373] ), .Y(new_n8184_));
  NAND2X1  g07182(.A(new_n8184_), .B(new_n8183_), .Y(new_n8185_));
  OAI21X1  g07183(.A0(new_n8182_), .A1(new_n8181_), .B0(new_n8185_), .Y(new_n8186_));
  INVX1    g07184(.A(\A[378] ), .Y(new_n8187_));
  INVX1    g07185(.A(\A[376] ), .Y(new_n8188_));
  OR2X1    g07186(.A(\A[377] ), .B(new_n8188_), .Y(new_n8189_));
  AOI21X1  g07187(.A0(\A[377] ), .A1(new_n8188_), .B0(new_n8187_), .Y(new_n8190_));
  XOR2X1   g07188(.A(\A[377] ), .B(\A[376] ), .Y(new_n8191_));
  AOI22X1  g07189(.A0(new_n8191_), .A1(new_n8187_), .B0(new_n8190_), .B1(new_n8189_), .Y(new_n8192_));
  AND2X1   g07190(.A(\A[377] ), .B(\A[376] ), .Y(new_n8193_));
  AOI21X1  g07191(.A0(new_n8191_), .A1(\A[378] ), .B0(new_n8193_), .Y(new_n8194_));
  AND2X1   g07192(.A(\A[374] ), .B(\A[373] ), .Y(new_n8195_));
  AOI21X1  g07193(.A0(new_n8184_), .A1(\A[375] ), .B0(new_n8195_), .Y(new_n8196_));
  XOR2X1   g07194(.A(new_n8192_), .B(new_n8186_), .Y(new_n8197_));
  INVX1    g07195(.A(\A[369] ), .Y(new_n8198_));
  INVX1    g07196(.A(\A[367] ), .Y(new_n8199_));
  OR2X1    g07197(.A(\A[368] ), .B(new_n8199_), .Y(new_n8200_));
  AOI21X1  g07198(.A0(\A[368] ), .A1(new_n8199_), .B0(new_n8198_), .Y(new_n8201_));
  XOR2X1   g07199(.A(\A[368] ), .B(\A[367] ), .Y(new_n8202_));
  AOI22X1  g07200(.A0(new_n8202_), .A1(new_n8198_), .B0(new_n8201_), .B1(new_n8200_), .Y(new_n8203_));
  INVX1    g07201(.A(\A[372] ), .Y(new_n8204_));
  INVX1    g07202(.A(\A[370] ), .Y(new_n8205_));
  OR2X1    g07203(.A(\A[371] ), .B(new_n8205_), .Y(new_n8206_));
  AOI21X1  g07204(.A0(\A[371] ), .A1(new_n8205_), .B0(new_n8204_), .Y(new_n8207_));
  XOR2X1   g07205(.A(\A[371] ), .B(\A[370] ), .Y(new_n8208_));
  AOI22X1  g07206(.A0(new_n8208_), .A1(new_n8204_), .B0(new_n8207_), .B1(new_n8206_), .Y(new_n8209_));
  AND2X1   g07207(.A(\A[371] ), .B(\A[370] ), .Y(new_n8210_));
  AOI21X1  g07208(.A0(new_n8208_), .A1(\A[372] ), .B0(new_n8210_), .Y(new_n8211_));
  AND2X1   g07209(.A(\A[368] ), .B(\A[367] ), .Y(new_n8212_));
  AOI21X1  g07210(.A0(new_n8202_), .A1(\A[369] ), .B0(new_n8212_), .Y(new_n8213_));
  XOR2X1   g07211(.A(new_n8209_), .B(new_n8203_), .Y(new_n8214_));
  XOR2X1   g07212(.A(new_n8214_), .B(new_n8197_), .Y(new_n8215_));
  XOR2X1   g07213(.A(new_n8215_), .B(new_n8179_), .Y(new_n8216_));
  OR2X1    g07214(.A(new_n8216_), .B(new_n8142_), .Y(new_n8217_));
  AND2X1   g07215(.A(new_n8109_), .B(new_n8077_), .Y(new_n8218_));
  XOR2X1   g07216(.A(new_n8132_), .B(new_n8102_), .Y(new_n8219_));
  NOR4X1   g07217(.A(new_n8101_), .B(new_n8095_), .C(new_n8130_), .D(new_n8071_), .Y(new_n8220_));
  OAI21X1  g07218(.A0(new_n8131_), .A1(new_n8107_), .B0(new_n8129_), .Y(new_n8221_));
  AOI22X1  g07219(.A0(new_n8221_), .A1(new_n8220_), .B0(new_n8108_), .B1(new_n8102_), .Y(new_n8222_));
  MX2X1    g07220(.A(new_n8222_), .B(new_n8219_), .S0(new_n8077_), .Y(new_n8223_));
  OAI21X1  g07221(.A0(new_n8222_), .A1(new_n8077_), .B0(new_n8117_), .Y(new_n8224_));
  OAI22X1  g07222(.A0(new_n8224_), .A1(new_n8218_), .B0(new_n8223_), .B1(new_n8117_), .Y(new_n8225_));
  AOI21X1  g07223(.A0(new_n8225_), .A1(new_n8045_), .B0(new_n8217_), .Y(new_n8226_));
  NOR2X1   g07224(.A(new_n8116_), .B(new_n8113_), .Y(new_n8227_));
  OAI21X1  g07225(.A0(new_n8222_), .A1(new_n8077_), .B0(new_n8227_), .Y(new_n8228_));
  OAI22X1  g07226(.A0(new_n8223_), .A1(new_n8227_), .B0(new_n8228_), .B1(new_n8218_), .Y(new_n8229_));
  MX2X1    g07227(.A(new_n8229_), .B(new_n8225_), .S0(new_n8045_), .Y(new_n8230_));
  AOI22X1  g07228(.A0(new_n8230_), .A1(new_n8217_), .B0(new_n8226_), .B1(new_n8139_), .Y(new_n8231_));
  INVX1    g07229(.A(\A[380] ), .Y(new_n8232_));
  AND2X1   g07230(.A(new_n8232_), .B(\A[379] ), .Y(new_n8233_));
  OAI21X1  g07231(.A0(new_n8232_), .A1(\A[379] ), .B0(\A[381] ), .Y(new_n8234_));
  NAND2X1  g07232(.A(new_n8165_), .B(new_n8161_), .Y(new_n8235_));
  OAI21X1  g07233(.A0(new_n8234_), .A1(new_n8233_), .B0(new_n8235_), .Y(new_n8236_));
  XOR2X1   g07234(.A(new_n8172_), .B(new_n8236_), .Y(new_n8237_));
  XOR2X1   g07235(.A(new_n8176_), .B(new_n8174_), .Y(new_n8238_));
  NOR2X1   g07236(.A(new_n8172_), .B(new_n8166_), .Y(new_n8239_));
  NOR2X1   g07237(.A(new_n8176_), .B(new_n8174_), .Y(new_n8240_));
  AOI21X1  g07238(.A0(new_n8239_), .A1(new_n8238_), .B0(new_n8240_), .Y(new_n8241_));
  XOR2X1   g07239(.A(new_n8239_), .B(new_n8238_), .Y(new_n8242_));
  OAI21X1  g07240(.A0(new_n8241_), .A1(new_n8237_), .B0(new_n8242_), .Y(new_n8243_));
  XOR2X1   g07241(.A(new_n8155_), .B(new_n8149_), .Y(new_n8244_));
  INVX1    g07242(.A(\A[385] ), .Y(new_n8245_));
  OR2X1    g07243(.A(\A[386] ), .B(new_n8245_), .Y(new_n8246_));
  AOI21X1  g07244(.A0(\A[386] ), .A1(new_n8245_), .B0(new_n8146_), .Y(new_n8247_));
  AOI22X1  g07245(.A0(new_n8147_), .A1(new_n8146_), .B0(new_n8247_), .B1(new_n8246_), .Y(new_n8248_));
  NOR4X1   g07246(.A(new_n8159_), .B(new_n8157_), .C(new_n8155_), .D(new_n8248_), .Y(new_n8249_));
  NOR4X1   g07247(.A(new_n8176_), .B(new_n8174_), .C(new_n8172_), .D(new_n8166_), .Y(new_n8250_));
  OR4X1    g07248(.A(new_n8250_), .B(new_n8237_), .C(new_n8249_), .D(new_n8244_), .Y(new_n8251_));
  XOR2X1   g07249(.A(new_n8159_), .B(new_n8157_), .Y(new_n8252_));
  NOR2X1   g07250(.A(new_n8155_), .B(new_n8248_), .Y(new_n8253_));
  NOR2X1   g07251(.A(new_n8159_), .B(new_n8157_), .Y(new_n8254_));
  AOI21X1  g07252(.A0(new_n8253_), .A1(new_n8252_), .B0(new_n8254_), .Y(new_n8255_));
  XOR2X1   g07253(.A(new_n8253_), .B(new_n8252_), .Y(new_n8256_));
  OAI21X1  g07254(.A0(new_n8255_), .A1(new_n8244_), .B0(new_n8256_), .Y(new_n8257_));
  XOR2X1   g07255(.A(new_n8257_), .B(new_n8251_), .Y(new_n8258_));
  NAND2X1  g07256(.A(new_n8258_), .B(new_n8243_), .Y(new_n8259_));
  OR2X1    g07257(.A(new_n8215_), .B(new_n8178_), .Y(new_n8260_));
  XOR2X1   g07258(.A(new_n8172_), .B(new_n8166_), .Y(new_n8261_));
  AND2X1   g07259(.A(new_n8171_), .B(\A[384] ), .Y(new_n8262_));
  OR2X1    g07260(.A(new_n8262_), .B(new_n8173_), .Y(new_n8263_));
  XOR2X1   g07261(.A(new_n8176_), .B(new_n8263_), .Y(new_n8264_));
  OR2X1    g07262(.A(new_n8172_), .B(new_n8166_), .Y(new_n8265_));
  OR2X1    g07263(.A(new_n8176_), .B(new_n8174_), .Y(new_n8266_));
  OAI21X1  g07264(.A0(new_n8265_), .A1(new_n8264_), .B0(new_n8266_), .Y(new_n8267_));
  XOR2X1   g07265(.A(new_n8239_), .B(new_n8264_), .Y(new_n8268_));
  AOI21X1  g07266(.A0(new_n8267_), .A1(new_n8261_), .B0(new_n8268_), .Y(new_n8269_));
  NOR4X1   g07267(.A(new_n8250_), .B(new_n8237_), .C(new_n8249_), .D(new_n8244_), .Y(new_n8270_));
  XOR2X1   g07268(.A(new_n8155_), .B(new_n8248_), .Y(new_n8271_));
  AND2X1   g07269(.A(new_n8154_), .B(\A[390] ), .Y(new_n8272_));
  OR2X1    g07270(.A(new_n8272_), .B(new_n8156_), .Y(new_n8273_));
  XOR2X1   g07271(.A(new_n8159_), .B(new_n8273_), .Y(new_n8274_));
  OR2X1    g07272(.A(new_n8155_), .B(new_n8248_), .Y(new_n8275_));
  OR2X1    g07273(.A(new_n8159_), .B(new_n8157_), .Y(new_n8276_));
  OAI21X1  g07274(.A0(new_n8275_), .A1(new_n8274_), .B0(new_n8276_), .Y(new_n8277_));
  XOR2X1   g07275(.A(new_n8275_), .B(new_n8252_), .Y(new_n8278_));
  AOI21X1  g07276(.A0(new_n8277_), .A1(new_n8271_), .B0(new_n8278_), .Y(new_n8279_));
  OR4X1    g07277(.A(new_n8237_), .B(new_n8249_), .C(new_n8278_), .D(new_n8244_), .Y(new_n8280_));
  OAI22X1  g07278(.A0(new_n8268_), .A1(new_n8241_), .B0(new_n8255_), .B1(new_n8244_), .Y(new_n8281_));
  OAI22X1  g07279(.A0(new_n8281_), .A1(new_n8280_), .B0(new_n8279_), .B1(new_n8270_), .Y(new_n8282_));
  AOI21X1  g07280(.A0(new_n8282_), .A1(new_n8269_), .B0(new_n8260_), .Y(new_n8283_));
  MX2X1    g07281(.A(new_n8282_), .B(new_n8258_), .S0(new_n8243_), .Y(new_n8284_));
  AOI22X1  g07282(.A0(new_n8284_), .A1(new_n8260_), .B0(new_n8283_), .B1(new_n8259_), .Y(new_n8285_));
  INVX1    g07283(.A(\A[368] ), .Y(new_n8286_));
  AND2X1   g07284(.A(new_n8286_), .B(\A[367] ), .Y(new_n8287_));
  OAI21X1  g07285(.A0(new_n8286_), .A1(\A[367] ), .B0(\A[369] ), .Y(new_n8288_));
  NAND2X1  g07286(.A(new_n8202_), .B(new_n8198_), .Y(new_n8289_));
  OAI21X1  g07287(.A0(new_n8288_), .A1(new_n8287_), .B0(new_n8289_), .Y(new_n8290_));
  XOR2X1   g07288(.A(new_n8209_), .B(new_n8290_), .Y(new_n8291_));
  XOR2X1   g07289(.A(new_n8213_), .B(new_n8211_), .Y(new_n8292_));
  NOR2X1   g07290(.A(new_n8209_), .B(new_n8203_), .Y(new_n8293_));
  NOR2X1   g07291(.A(new_n8213_), .B(new_n8211_), .Y(new_n8294_));
  AOI21X1  g07292(.A0(new_n8293_), .A1(new_n8292_), .B0(new_n8294_), .Y(new_n8295_));
  XOR2X1   g07293(.A(new_n8293_), .B(new_n8292_), .Y(new_n8296_));
  OAI21X1  g07294(.A0(new_n8295_), .A1(new_n8291_), .B0(new_n8296_), .Y(new_n8297_));
  XOR2X1   g07295(.A(new_n8192_), .B(new_n8186_), .Y(new_n8298_));
  INVX1    g07296(.A(\A[373] ), .Y(new_n8299_));
  OR2X1    g07297(.A(\A[374] ), .B(new_n8299_), .Y(new_n8300_));
  AOI21X1  g07298(.A0(\A[374] ), .A1(new_n8299_), .B0(new_n8183_), .Y(new_n8301_));
  AOI22X1  g07299(.A0(new_n8184_), .A1(new_n8183_), .B0(new_n8301_), .B1(new_n8300_), .Y(new_n8302_));
  NOR4X1   g07300(.A(new_n8196_), .B(new_n8194_), .C(new_n8192_), .D(new_n8302_), .Y(new_n8303_));
  NOR4X1   g07301(.A(new_n8213_), .B(new_n8211_), .C(new_n8209_), .D(new_n8203_), .Y(new_n8304_));
  OR4X1    g07302(.A(new_n8304_), .B(new_n8291_), .C(new_n8303_), .D(new_n8298_), .Y(new_n8305_));
  XOR2X1   g07303(.A(new_n8192_), .B(new_n8302_), .Y(new_n8306_));
  AND2X1   g07304(.A(new_n8191_), .B(\A[378] ), .Y(new_n8307_));
  OR2X1    g07305(.A(new_n8307_), .B(new_n8193_), .Y(new_n8308_));
  XOR2X1   g07306(.A(new_n8196_), .B(new_n8308_), .Y(new_n8309_));
  OR2X1    g07307(.A(new_n8192_), .B(new_n8302_), .Y(new_n8310_));
  OR2X1    g07308(.A(new_n8196_), .B(new_n8194_), .Y(new_n8311_));
  OAI21X1  g07309(.A0(new_n8310_), .A1(new_n8309_), .B0(new_n8311_), .Y(new_n8312_));
  NOR2X1   g07310(.A(new_n8192_), .B(new_n8302_), .Y(new_n8313_));
  XOR2X1   g07311(.A(new_n8313_), .B(new_n8309_), .Y(new_n8314_));
  AOI21X1  g07312(.A0(new_n8312_), .A1(new_n8306_), .B0(new_n8314_), .Y(new_n8315_));
  XOR2X1   g07313(.A(new_n8315_), .B(new_n8305_), .Y(new_n8316_));
  XOR2X1   g07314(.A(new_n8196_), .B(new_n8194_), .Y(new_n8317_));
  NOR2X1   g07315(.A(new_n8196_), .B(new_n8194_), .Y(new_n8318_));
  AOI21X1  g07316(.A0(new_n8313_), .A1(new_n8317_), .B0(new_n8318_), .Y(new_n8319_));
  XOR2X1   g07317(.A(new_n8313_), .B(new_n8317_), .Y(new_n8320_));
  OAI21X1  g07318(.A0(new_n8319_), .A1(new_n8298_), .B0(new_n8320_), .Y(new_n8321_));
  NOR4X1   g07319(.A(new_n8291_), .B(new_n8314_), .C(new_n8312_), .D(new_n8298_), .Y(new_n8322_));
  AOI21X1  g07320(.A0(new_n8312_), .A1(new_n8306_), .B0(new_n8304_), .Y(new_n8323_));
  AOI22X1  g07321(.A0(new_n8323_), .A1(new_n8322_), .B0(new_n8321_), .B1(new_n8305_), .Y(new_n8324_));
  MX2X1    g07322(.A(new_n8324_), .B(new_n8316_), .S0(new_n8297_), .Y(new_n8325_));
  NOR2X1   g07323(.A(new_n8215_), .B(new_n8178_), .Y(new_n8326_));
  AOI21X1  g07324(.A0(new_n8282_), .A1(new_n8269_), .B0(new_n8326_), .Y(new_n8327_));
  AOI22X1  g07325(.A0(new_n8327_), .A1(new_n8259_), .B0(new_n8284_), .B1(new_n8326_), .Y(new_n8328_));
  MX2X1    g07326(.A(new_n8328_), .B(new_n8285_), .S0(new_n8325_), .Y(new_n8329_));
  NOR2X1   g07327(.A(new_n8216_), .B(new_n8142_), .Y(new_n8330_));
  AOI21X1  g07328(.A0(new_n8225_), .A1(new_n8045_), .B0(new_n8330_), .Y(new_n8331_));
  AOI22X1  g07329(.A0(new_n8331_), .A1(new_n8139_), .B0(new_n8230_), .B1(new_n8330_), .Y(new_n8332_));
  MX2X1    g07330(.A(new_n8332_), .B(new_n8231_), .S0(new_n8329_), .Y(new_n8333_));
  INVX1    g07331(.A(\A[429] ), .Y(new_n8334_));
  INVX1    g07332(.A(\A[428] ), .Y(new_n8335_));
  OR2X1    g07333(.A(new_n8335_), .B(\A[427] ), .Y(new_n8336_));
  AOI21X1  g07334(.A0(new_n8335_), .A1(\A[427] ), .B0(new_n8334_), .Y(new_n8337_));
  XOR2X1   g07335(.A(\A[428] ), .B(\A[427] ), .Y(new_n8338_));
  AOI22X1  g07336(.A0(new_n8338_), .A1(new_n8334_), .B0(new_n8337_), .B1(new_n8336_), .Y(new_n8339_));
  INVX1    g07337(.A(\A[432] ), .Y(new_n8340_));
  INVX1    g07338(.A(\A[431] ), .Y(new_n8341_));
  OR2X1    g07339(.A(new_n8341_), .B(\A[430] ), .Y(new_n8342_));
  AOI21X1  g07340(.A0(new_n8341_), .A1(\A[430] ), .B0(new_n8340_), .Y(new_n8343_));
  XOR2X1   g07341(.A(\A[431] ), .B(\A[430] ), .Y(new_n8344_));
  AOI22X1  g07342(.A0(new_n8344_), .A1(new_n8340_), .B0(new_n8343_), .B1(new_n8342_), .Y(new_n8345_));
  OR2X1    g07343(.A(new_n8345_), .B(new_n8339_), .Y(new_n8346_));
  AND2X1   g07344(.A(\A[431] ), .B(\A[430] ), .Y(new_n8347_));
  AND2X1   g07345(.A(new_n8344_), .B(\A[432] ), .Y(new_n8348_));
  OR2X1    g07346(.A(new_n8348_), .B(new_n8347_), .Y(new_n8349_));
  AND2X1   g07347(.A(\A[428] ), .B(\A[427] ), .Y(new_n8350_));
  AOI21X1  g07348(.A0(new_n8338_), .A1(\A[429] ), .B0(new_n8350_), .Y(new_n8351_));
  XOR2X1   g07349(.A(new_n8351_), .B(new_n8349_), .Y(new_n8352_));
  XOR2X1   g07350(.A(new_n8352_), .B(new_n8346_), .Y(new_n8353_));
  INVX1    g07351(.A(\A[427] ), .Y(new_n8354_));
  AND2X1   g07352(.A(\A[428] ), .B(new_n8354_), .Y(new_n8355_));
  OAI21X1  g07353(.A0(\A[428] ), .A1(new_n8354_), .B0(\A[429] ), .Y(new_n8356_));
  NAND2X1  g07354(.A(new_n8338_), .B(new_n8334_), .Y(new_n8357_));
  OAI21X1  g07355(.A0(new_n8356_), .A1(new_n8355_), .B0(new_n8357_), .Y(new_n8358_));
  XOR2X1   g07356(.A(new_n8345_), .B(new_n8358_), .Y(new_n8359_));
  NOR2X1   g07357(.A(new_n8345_), .B(new_n8339_), .Y(new_n8360_));
  AOI21X1  g07358(.A0(new_n8344_), .A1(\A[432] ), .B0(new_n8347_), .Y(new_n8361_));
  XOR2X1   g07359(.A(new_n8351_), .B(new_n8361_), .Y(new_n8362_));
  NOR2X1   g07360(.A(new_n8351_), .B(new_n8361_), .Y(new_n8363_));
  AOI21X1  g07361(.A0(new_n8362_), .A1(new_n8360_), .B0(new_n8363_), .Y(new_n8364_));
  OAI21X1  g07362(.A0(new_n8364_), .A1(new_n8359_), .B0(new_n8353_), .Y(new_n8365_));
  AND2X1   g07363(.A(\A[437] ), .B(\A[436] ), .Y(new_n8366_));
  XOR2X1   g07364(.A(\A[437] ), .B(\A[436] ), .Y(new_n8367_));
  AOI21X1  g07365(.A0(new_n8367_), .A1(\A[438] ), .B0(new_n8366_), .Y(new_n8368_));
  AND2X1   g07366(.A(\A[434] ), .B(\A[433] ), .Y(new_n8369_));
  XOR2X1   g07367(.A(\A[434] ), .B(\A[433] ), .Y(new_n8370_));
  AOI21X1  g07368(.A0(new_n8370_), .A1(\A[435] ), .B0(new_n8369_), .Y(new_n8371_));
  INVX1    g07369(.A(\A[435] ), .Y(new_n8372_));
  INVX1    g07370(.A(\A[434] ), .Y(new_n8373_));
  OR2X1    g07371(.A(new_n8373_), .B(\A[433] ), .Y(new_n8374_));
  AOI21X1  g07372(.A0(new_n8373_), .A1(\A[433] ), .B0(new_n8372_), .Y(new_n8375_));
  AOI22X1  g07373(.A0(new_n8375_), .A1(new_n8374_), .B0(new_n8370_), .B1(new_n8372_), .Y(new_n8376_));
  INVX1    g07374(.A(\A[438] ), .Y(new_n8377_));
  INVX1    g07375(.A(\A[437] ), .Y(new_n8378_));
  OR2X1    g07376(.A(new_n8378_), .B(\A[436] ), .Y(new_n8379_));
  AOI21X1  g07377(.A0(new_n8378_), .A1(\A[436] ), .B0(new_n8377_), .Y(new_n8380_));
  AOI22X1  g07378(.A0(new_n8380_), .A1(new_n8379_), .B0(new_n8367_), .B1(new_n8377_), .Y(new_n8381_));
  NOR4X1   g07379(.A(new_n8381_), .B(new_n8376_), .C(new_n8371_), .D(new_n8368_), .Y(new_n8382_));
  NOR4X1   g07380(.A(new_n8351_), .B(new_n8361_), .C(new_n8345_), .D(new_n8339_), .Y(new_n8383_));
  INVX1    g07381(.A(\A[433] ), .Y(new_n8384_));
  AND2X1   g07382(.A(\A[434] ), .B(new_n8384_), .Y(new_n8385_));
  OAI21X1  g07383(.A0(\A[434] ), .A1(new_n8384_), .B0(\A[435] ), .Y(new_n8386_));
  NAND2X1  g07384(.A(new_n8370_), .B(new_n8372_), .Y(new_n8387_));
  OAI21X1  g07385(.A0(new_n8386_), .A1(new_n8385_), .B0(new_n8387_), .Y(new_n8388_));
  XOR2X1   g07386(.A(new_n8381_), .B(new_n8388_), .Y(new_n8389_));
  OR4X1    g07387(.A(new_n8389_), .B(new_n8383_), .C(new_n8382_), .D(new_n8359_), .Y(new_n8390_));
  XOR2X1   g07388(.A(new_n8371_), .B(new_n8368_), .Y(new_n8391_));
  NOR2X1   g07389(.A(new_n8381_), .B(new_n8376_), .Y(new_n8392_));
  NOR2X1   g07390(.A(new_n8371_), .B(new_n8368_), .Y(new_n8393_));
  AOI21X1  g07391(.A0(new_n8392_), .A1(new_n8391_), .B0(new_n8393_), .Y(new_n8394_));
  XOR2X1   g07392(.A(new_n8392_), .B(new_n8391_), .Y(new_n8395_));
  OAI21X1  g07393(.A0(new_n8389_), .A1(new_n8394_), .B0(new_n8395_), .Y(new_n8396_));
  XOR2X1   g07394(.A(new_n8396_), .B(new_n8390_), .Y(new_n8397_));
  NAND2X1  g07395(.A(new_n8397_), .B(new_n8365_), .Y(new_n8398_));
  XOR2X1   g07396(.A(new_n8345_), .B(new_n8339_), .Y(new_n8399_));
  OAI21X1  g07397(.A0(new_n8389_), .A1(new_n8382_), .B0(new_n8399_), .Y(new_n8400_));
  OR4X1    g07398(.A(new_n8381_), .B(new_n8376_), .C(new_n8371_), .D(new_n8368_), .Y(new_n8401_));
  XOR2X1   g07399(.A(new_n8381_), .B(new_n8376_), .Y(new_n8402_));
  XOR2X1   g07400(.A(new_n8345_), .B(new_n8358_), .Y(new_n8403_));
  NAND3X1  g07401(.A(new_n8403_), .B(new_n8402_), .C(new_n8401_), .Y(new_n8404_));
  AND2X1   g07402(.A(new_n8404_), .B(new_n8400_), .Y(new_n8405_));
  INVX1    g07403(.A(\A[422] ), .Y(new_n8406_));
  AND2X1   g07404(.A(new_n8406_), .B(\A[421] ), .Y(new_n8407_));
  OAI21X1  g07405(.A0(new_n8406_), .A1(\A[421] ), .B0(\A[423] ), .Y(new_n8408_));
  INVX1    g07406(.A(\A[423] ), .Y(new_n8409_));
  XOR2X1   g07407(.A(\A[422] ), .B(\A[421] ), .Y(new_n8410_));
  NAND2X1  g07408(.A(new_n8410_), .B(new_n8409_), .Y(new_n8411_));
  OAI21X1  g07409(.A0(new_n8408_), .A1(new_n8407_), .B0(new_n8411_), .Y(new_n8412_));
  INVX1    g07410(.A(\A[426] ), .Y(new_n8413_));
  INVX1    g07411(.A(\A[424] ), .Y(new_n8414_));
  OR2X1    g07412(.A(\A[425] ), .B(new_n8414_), .Y(new_n8415_));
  AOI21X1  g07413(.A0(\A[425] ), .A1(new_n8414_), .B0(new_n8413_), .Y(new_n8416_));
  XOR2X1   g07414(.A(\A[425] ), .B(\A[424] ), .Y(new_n8417_));
  AOI22X1  g07415(.A0(new_n8417_), .A1(new_n8413_), .B0(new_n8416_), .B1(new_n8415_), .Y(new_n8418_));
  AND2X1   g07416(.A(\A[425] ), .B(\A[424] ), .Y(new_n8419_));
  AOI21X1  g07417(.A0(new_n8417_), .A1(\A[426] ), .B0(new_n8419_), .Y(new_n8420_));
  AND2X1   g07418(.A(\A[422] ), .B(\A[421] ), .Y(new_n8421_));
  AOI21X1  g07419(.A0(new_n8410_), .A1(\A[423] ), .B0(new_n8421_), .Y(new_n8422_));
  XOR2X1   g07420(.A(new_n8418_), .B(new_n8412_), .Y(new_n8423_));
  INVX1    g07421(.A(\A[417] ), .Y(new_n8424_));
  INVX1    g07422(.A(\A[415] ), .Y(new_n8425_));
  OR2X1    g07423(.A(\A[416] ), .B(new_n8425_), .Y(new_n8426_));
  AOI21X1  g07424(.A0(\A[416] ), .A1(new_n8425_), .B0(new_n8424_), .Y(new_n8427_));
  XOR2X1   g07425(.A(\A[416] ), .B(\A[415] ), .Y(new_n8428_));
  AOI22X1  g07426(.A0(new_n8428_), .A1(new_n8424_), .B0(new_n8427_), .B1(new_n8426_), .Y(new_n8429_));
  INVX1    g07427(.A(\A[420] ), .Y(new_n8430_));
  INVX1    g07428(.A(\A[418] ), .Y(new_n8431_));
  OR2X1    g07429(.A(\A[419] ), .B(new_n8431_), .Y(new_n8432_));
  AOI21X1  g07430(.A0(\A[419] ), .A1(new_n8431_), .B0(new_n8430_), .Y(new_n8433_));
  XOR2X1   g07431(.A(\A[419] ), .B(\A[418] ), .Y(new_n8434_));
  AOI22X1  g07432(.A0(new_n8434_), .A1(new_n8430_), .B0(new_n8433_), .B1(new_n8432_), .Y(new_n8435_));
  AND2X1   g07433(.A(\A[419] ), .B(\A[418] ), .Y(new_n8436_));
  AOI21X1  g07434(.A0(new_n8434_), .A1(\A[420] ), .B0(new_n8436_), .Y(new_n8437_));
  AND2X1   g07435(.A(\A[416] ), .B(\A[415] ), .Y(new_n8438_));
  AOI21X1  g07436(.A0(new_n8428_), .A1(\A[417] ), .B0(new_n8438_), .Y(new_n8439_));
  XOR2X1   g07437(.A(new_n8435_), .B(new_n8429_), .Y(new_n8440_));
  XOR2X1   g07438(.A(new_n8440_), .B(new_n8423_), .Y(new_n8441_));
  OR2X1    g07439(.A(new_n8441_), .B(new_n8405_), .Y(new_n8442_));
  XOR2X1   g07440(.A(new_n8352_), .B(new_n8360_), .Y(new_n8443_));
  XOR2X1   g07441(.A(new_n8345_), .B(new_n8339_), .Y(new_n8444_));
  OR2X1    g07442(.A(new_n8351_), .B(new_n8361_), .Y(new_n8445_));
  OAI21X1  g07443(.A0(new_n8352_), .A1(new_n8346_), .B0(new_n8445_), .Y(new_n8446_));
  AOI21X1  g07444(.A0(new_n8446_), .A1(new_n8444_), .B0(new_n8443_), .Y(new_n8447_));
  NOR4X1   g07445(.A(new_n8389_), .B(new_n8383_), .C(new_n8382_), .D(new_n8359_), .Y(new_n8448_));
  AND2X1   g07446(.A(new_n8367_), .B(\A[438] ), .Y(new_n8449_));
  OR2X1    g07447(.A(new_n8449_), .B(new_n8366_), .Y(new_n8450_));
  XOR2X1   g07448(.A(new_n8371_), .B(new_n8450_), .Y(new_n8451_));
  OR2X1    g07449(.A(new_n8381_), .B(new_n8376_), .Y(new_n8452_));
  OR2X1    g07450(.A(new_n8371_), .B(new_n8368_), .Y(new_n8453_));
  OAI21X1  g07451(.A0(new_n8452_), .A1(new_n8451_), .B0(new_n8453_), .Y(new_n8454_));
  XOR2X1   g07452(.A(new_n8392_), .B(new_n8451_), .Y(new_n8455_));
  AOI21X1  g07453(.A0(new_n8402_), .A1(new_n8454_), .B0(new_n8455_), .Y(new_n8456_));
  OR4X1    g07454(.A(new_n8389_), .B(new_n8383_), .C(new_n8455_), .D(new_n8359_), .Y(new_n8457_));
  AOI21X1  g07455(.A0(new_n8389_), .A1(new_n8455_), .B0(new_n8394_), .Y(new_n8458_));
  OAI22X1  g07456(.A0(new_n8458_), .A1(new_n8457_), .B0(new_n8456_), .B1(new_n8448_), .Y(new_n8459_));
  AOI21X1  g07457(.A0(new_n8459_), .A1(new_n8447_), .B0(new_n8442_), .Y(new_n8460_));
  MX2X1    g07458(.A(new_n8459_), .B(new_n8397_), .S0(new_n8365_), .Y(new_n8461_));
  AOI22X1  g07459(.A0(new_n8461_), .A1(new_n8442_), .B0(new_n8460_), .B1(new_n8398_), .Y(new_n8462_));
  INVX1    g07460(.A(\A[416] ), .Y(new_n8463_));
  AND2X1   g07461(.A(new_n8463_), .B(\A[415] ), .Y(new_n8464_));
  OAI21X1  g07462(.A0(new_n8463_), .A1(\A[415] ), .B0(\A[417] ), .Y(new_n8465_));
  NAND2X1  g07463(.A(new_n8428_), .B(new_n8424_), .Y(new_n8466_));
  OAI21X1  g07464(.A0(new_n8465_), .A1(new_n8464_), .B0(new_n8466_), .Y(new_n8467_));
  XOR2X1   g07465(.A(new_n8435_), .B(new_n8467_), .Y(new_n8468_));
  XOR2X1   g07466(.A(new_n8439_), .B(new_n8437_), .Y(new_n8469_));
  NOR2X1   g07467(.A(new_n8435_), .B(new_n8429_), .Y(new_n8470_));
  NOR2X1   g07468(.A(new_n8439_), .B(new_n8437_), .Y(new_n8471_));
  AOI21X1  g07469(.A0(new_n8470_), .A1(new_n8469_), .B0(new_n8471_), .Y(new_n8472_));
  XOR2X1   g07470(.A(new_n8470_), .B(new_n8469_), .Y(new_n8473_));
  OAI21X1  g07471(.A0(new_n8472_), .A1(new_n8468_), .B0(new_n8473_), .Y(new_n8474_));
  XOR2X1   g07472(.A(new_n8418_), .B(new_n8412_), .Y(new_n8475_));
  INVX1    g07473(.A(\A[421] ), .Y(new_n8476_));
  OR2X1    g07474(.A(\A[422] ), .B(new_n8476_), .Y(new_n8477_));
  AOI21X1  g07475(.A0(\A[422] ), .A1(new_n8476_), .B0(new_n8409_), .Y(new_n8478_));
  AOI22X1  g07476(.A0(new_n8410_), .A1(new_n8409_), .B0(new_n8478_), .B1(new_n8477_), .Y(new_n8479_));
  NOR4X1   g07477(.A(new_n8422_), .B(new_n8420_), .C(new_n8418_), .D(new_n8479_), .Y(new_n8480_));
  NOR4X1   g07478(.A(new_n8439_), .B(new_n8437_), .C(new_n8435_), .D(new_n8429_), .Y(new_n8481_));
  OR4X1    g07479(.A(new_n8481_), .B(new_n8468_), .C(new_n8480_), .D(new_n8475_), .Y(new_n8482_));
  XOR2X1   g07480(.A(new_n8418_), .B(new_n8479_), .Y(new_n8483_));
  AND2X1   g07481(.A(new_n8417_), .B(\A[426] ), .Y(new_n8484_));
  OR2X1    g07482(.A(new_n8484_), .B(new_n8419_), .Y(new_n8485_));
  XOR2X1   g07483(.A(new_n8422_), .B(new_n8485_), .Y(new_n8486_));
  OR2X1    g07484(.A(new_n8418_), .B(new_n8479_), .Y(new_n8487_));
  OR2X1    g07485(.A(new_n8422_), .B(new_n8420_), .Y(new_n8488_));
  OAI21X1  g07486(.A0(new_n8487_), .A1(new_n8486_), .B0(new_n8488_), .Y(new_n8489_));
  NOR2X1   g07487(.A(new_n8418_), .B(new_n8479_), .Y(new_n8490_));
  XOR2X1   g07488(.A(new_n8490_), .B(new_n8486_), .Y(new_n8491_));
  AOI21X1  g07489(.A0(new_n8489_), .A1(new_n8483_), .B0(new_n8491_), .Y(new_n8492_));
  XOR2X1   g07490(.A(new_n8492_), .B(new_n8482_), .Y(new_n8493_));
  XOR2X1   g07491(.A(new_n8422_), .B(new_n8420_), .Y(new_n8494_));
  NOR2X1   g07492(.A(new_n8422_), .B(new_n8420_), .Y(new_n8495_));
  AOI21X1  g07493(.A0(new_n8490_), .A1(new_n8494_), .B0(new_n8495_), .Y(new_n8496_));
  XOR2X1   g07494(.A(new_n8490_), .B(new_n8494_), .Y(new_n8497_));
  OAI21X1  g07495(.A0(new_n8496_), .A1(new_n8475_), .B0(new_n8497_), .Y(new_n8498_));
  NOR4X1   g07496(.A(new_n8468_), .B(new_n8491_), .C(new_n8489_), .D(new_n8475_), .Y(new_n8499_));
  AOI21X1  g07497(.A0(new_n8489_), .A1(new_n8483_), .B0(new_n8481_), .Y(new_n8500_));
  AOI22X1  g07498(.A0(new_n8500_), .A1(new_n8499_), .B0(new_n8498_), .B1(new_n8482_), .Y(new_n8501_));
  MX2X1    g07499(.A(new_n8501_), .B(new_n8493_), .S0(new_n8474_), .Y(new_n8502_));
  AOI21X1  g07500(.A0(new_n8404_), .A1(new_n8400_), .B0(new_n8441_), .Y(new_n8503_));
  AOI21X1  g07501(.A0(new_n8459_), .A1(new_n8447_), .B0(new_n8503_), .Y(new_n8504_));
  AOI22X1  g07502(.A0(new_n8504_), .A1(new_n8398_), .B0(new_n8461_), .B1(new_n8503_), .Y(new_n8505_));
  MX2X1    g07503(.A(new_n8505_), .B(new_n8462_), .S0(new_n8502_), .Y(new_n8506_));
  INVX1    g07504(.A(\A[441] ), .Y(new_n8507_));
  INVX1    g07505(.A(\A[440] ), .Y(new_n8508_));
  OR2X1    g07506(.A(new_n8508_), .B(\A[439] ), .Y(new_n8509_));
  AOI21X1  g07507(.A0(new_n8508_), .A1(\A[439] ), .B0(new_n8507_), .Y(new_n8510_));
  XOR2X1   g07508(.A(\A[440] ), .B(\A[439] ), .Y(new_n8511_));
  AOI22X1  g07509(.A0(new_n8511_), .A1(new_n8507_), .B0(new_n8510_), .B1(new_n8509_), .Y(new_n8512_));
  INVX1    g07510(.A(\A[444] ), .Y(new_n8513_));
  INVX1    g07511(.A(\A[443] ), .Y(new_n8514_));
  OR2X1    g07512(.A(new_n8514_), .B(\A[442] ), .Y(new_n8515_));
  AOI21X1  g07513(.A0(new_n8514_), .A1(\A[442] ), .B0(new_n8513_), .Y(new_n8516_));
  XOR2X1   g07514(.A(\A[443] ), .B(\A[442] ), .Y(new_n8517_));
  AOI22X1  g07515(.A0(new_n8517_), .A1(new_n8513_), .B0(new_n8516_), .B1(new_n8515_), .Y(new_n8518_));
  OR2X1    g07516(.A(new_n8518_), .B(new_n8512_), .Y(new_n8519_));
  AND2X1   g07517(.A(\A[443] ), .B(\A[442] ), .Y(new_n8520_));
  AND2X1   g07518(.A(new_n8517_), .B(\A[444] ), .Y(new_n8521_));
  OR2X1    g07519(.A(new_n8521_), .B(new_n8520_), .Y(new_n8522_));
  AND2X1   g07520(.A(\A[440] ), .B(\A[439] ), .Y(new_n8523_));
  AOI21X1  g07521(.A0(new_n8511_), .A1(\A[441] ), .B0(new_n8523_), .Y(new_n8524_));
  XOR2X1   g07522(.A(new_n8524_), .B(new_n8522_), .Y(new_n8525_));
  XOR2X1   g07523(.A(new_n8525_), .B(new_n8519_), .Y(new_n8526_));
  INVX1    g07524(.A(\A[439] ), .Y(new_n8527_));
  AND2X1   g07525(.A(\A[440] ), .B(new_n8527_), .Y(new_n8528_));
  OAI21X1  g07526(.A0(\A[440] ), .A1(new_n8527_), .B0(\A[441] ), .Y(new_n8529_));
  NAND2X1  g07527(.A(new_n8511_), .B(new_n8507_), .Y(new_n8530_));
  OAI21X1  g07528(.A0(new_n8529_), .A1(new_n8528_), .B0(new_n8530_), .Y(new_n8531_));
  XOR2X1   g07529(.A(new_n8518_), .B(new_n8531_), .Y(new_n8532_));
  NOR2X1   g07530(.A(new_n8518_), .B(new_n8512_), .Y(new_n8533_));
  AOI21X1  g07531(.A0(new_n8517_), .A1(\A[444] ), .B0(new_n8520_), .Y(new_n8534_));
  XOR2X1   g07532(.A(new_n8524_), .B(new_n8534_), .Y(new_n8535_));
  NOR2X1   g07533(.A(new_n8524_), .B(new_n8534_), .Y(new_n8536_));
  AOI21X1  g07534(.A0(new_n8535_), .A1(new_n8533_), .B0(new_n8536_), .Y(new_n8537_));
  OAI21X1  g07535(.A0(new_n8537_), .A1(new_n8532_), .B0(new_n8526_), .Y(new_n8538_));
  AND2X1   g07536(.A(\A[449] ), .B(\A[448] ), .Y(new_n8539_));
  XOR2X1   g07537(.A(\A[449] ), .B(\A[448] ), .Y(new_n8540_));
  AOI21X1  g07538(.A0(new_n8540_), .A1(\A[450] ), .B0(new_n8539_), .Y(new_n8541_));
  AND2X1   g07539(.A(\A[446] ), .B(\A[445] ), .Y(new_n8542_));
  XOR2X1   g07540(.A(\A[446] ), .B(\A[445] ), .Y(new_n8543_));
  AOI21X1  g07541(.A0(new_n8543_), .A1(\A[447] ), .B0(new_n8542_), .Y(new_n8544_));
  INVX1    g07542(.A(\A[447] ), .Y(new_n8545_));
  INVX1    g07543(.A(\A[446] ), .Y(new_n8546_));
  OR2X1    g07544(.A(new_n8546_), .B(\A[445] ), .Y(new_n8547_));
  AOI21X1  g07545(.A0(new_n8546_), .A1(\A[445] ), .B0(new_n8545_), .Y(new_n8548_));
  AOI22X1  g07546(.A0(new_n8548_), .A1(new_n8547_), .B0(new_n8543_), .B1(new_n8545_), .Y(new_n8549_));
  INVX1    g07547(.A(\A[450] ), .Y(new_n8550_));
  INVX1    g07548(.A(\A[449] ), .Y(new_n8551_));
  OR2X1    g07549(.A(new_n8551_), .B(\A[448] ), .Y(new_n8552_));
  AOI21X1  g07550(.A0(new_n8551_), .A1(\A[448] ), .B0(new_n8550_), .Y(new_n8553_));
  AOI22X1  g07551(.A0(new_n8553_), .A1(new_n8552_), .B0(new_n8540_), .B1(new_n8550_), .Y(new_n8554_));
  NOR4X1   g07552(.A(new_n8554_), .B(new_n8549_), .C(new_n8544_), .D(new_n8541_), .Y(new_n8555_));
  NOR4X1   g07553(.A(new_n8524_), .B(new_n8534_), .C(new_n8518_), .D(new_n8512_), .Y(new_n8556_));
  INVX1    g07554(.A(\A[445] ), .Y(new_n8557_));
  AND2X1   g07555(.A(\A[446] ), .B(new_n8557_), .Y(new_n8558_));
  OAI21X1  g07556(.A0(\A[446] ), .A1(new_n8557_), .B0(\A[447] ), .Y(new_n8559_));
  NAND2X1  g07557(.A(new_n8543_), .B(new_n8545_), .Y(new_n8560_));
  OAI21X1  g07558(.A0(new_n8559_), .A1(new_n8558_), .B0(new_n8560_), .Y(new_n8561_));
  XOR2X1   g07559(.A(new_n8554_), .B(new_n8561_), .Y(new_n8562_));
  OR4X1    g07560(.A(new_n8562_), .B(new_n8556_), .C(new_n8555_), .D(new_n8532_), .Y(new_n8563_));
  AND2X1   g07561(.A(new_n8540_), .B(\A[450] ), .Y(new_n8564_));
  OR2X1    g07562(.A(new_n8564_), .B(new_n8539_), .Y(new_n8565_));
  XOR2X1   g07563(.A(new_n8544_), .B(new_n8565_), .Y(new_n8566_));
  OR2X1    g07564(.A(new_n8554_), .B(new_n8549_), .Y(new_n8567_));
  OR2X1    g07565(.A(new_n8544_), .B(new_n8541_), .Y(new_n8568_));
  OAI21X1  g07566(.A0(new_n8567_), .A1(new_n8566_), .B0(new_n8568_), .Y(new_n8569_));
  NOR2X1   g07567(.A(new_n8554_), .B(new_n8549_), .Y(new_n8570_));
  XOR2X1   g07568(.A(new_n8570_), .B(new_n8566_), .Y(new_n8571_));
  XOR2X1   g07569(.A(new_n8554_), .B(new_n8549_), .Y(new_n8572_));
  AOI21X1  g07570(.A0(new_n8572_), .A1(new_n8569_), .B0(new_n8571_), .Y(new_n8573_));
  XOR2X1   g07571(.A(new_n8573_), .B(new_n8563_), .Y(new_n8574_));
  XOR2X1   g07572(.A(new_n8544_), .B(new_n8541_), .Y(new_n8575_));
  NOR2X1   g07573(.A(new_n8544_), .B(new_n8541_), .Y(new_n8576_));
  AOI21X1  g07574(.A0(new_n8570_), .A1(new_n8575_), .B0(new_n8576_), .Y(new_n8577_));
  XOR2X1   g07575(.A(new_n8570_), .B(new_n8575_), .Y(new_n8578_));
  OAI21X1  g07576(.A0(new_n8562_), .A1(new_n8577_), .B0(new_n8578_), .Y(new_n8579_));
  NOR4X1   g07577(.A(new_n8562_), .B(new_n8556_), .C(new_n8571_), .D(new_n8532_), .Y(new_n8580_));
  OAI21X1  g07578(.A0(new_n8572_), .A1(new_n8578_), .B0(new_n8569_), .Y(new_n8581_));
  AOI22X1  g07579(.A0(new_n8581_), .A1(new_n8580_), .B0(new_n8579_), .B1(new_n8563_), .Y(new_n8582_));
  MX2X1    g07580(.A(new_n8582_), .B(new_n8574_), .S0(new_n8538_), .Y(new_n8583_));
  INVX1    g07581(.A(\A[453] ), .Y(new_n8584_));
  INVX1    g07582(.A(\A[452] ), .Y(new_n8585_));
  OR2X1    g07583(.A(new_n8585_), .B(\A[451] ), .Y(new_n8586_));
  AOI21X1  g07584(.A0(new_n8585_), .A1(\A[451] ), .B0(new_n8584_), .Y(new_n8587_));
  XOR2X1   g07585(.A(\A[452] ), .B(\A[451] ), .Y(new_n8588_));
  AOI22X1  g07586(.A0(new_n8588_), .A1(new_n8584_), .B0(new_n8587_), .B1(new_n8586_), .Y(new_n8589_));
  INVX1    g07587(.A(\A[456] ), .Y(new_n8590_));
  INVX1    g07588(.A(\A[455] ), .Y(new_n8591_));
  OR2X1    g07589(.A(new_n8591_), .B(\A[454] ), .Y(new_n8592_));
  AOI21X1  g07590(.A0(new_n8591_), .A1(\A[454] ), .B0(new_n8590_), .Y(new_n8593_));
  XOR2X1   g07591(.A(\A[455] ), .B(\A[454] ), .Y(new_n8594_));
  AOI22X1  g07592(.A0(new_n8594_), .A1(new_n8590_), .B0(new_n8593_), .B1(new_n8592_), .Y(new_n8595_));
  OR2X1    g07593(.A(new_n8595_), .B(new_n8589_), .Y(new_n8596_));
  AND2X1   g07594(.A(\A[455] ), .B(\A[454] ), .Y(new_n8597_));
  AND2X1   g07595(.A(new_n8594_), .B(\A[456] ), .Y(new_n8598_));
  OR2X1    g07596(.A(new_n8598_), .B(new_n8597_), .Y(new_n8599_));
  AND2X1   g07597(.A(\A[452] ), .B(\A[451] ), .Y(new_n8600_));
  AOI21X1  g07598(.A0(new_n8588_), .A1(\A[453] ), .B0(new_n8600_), .Y(new_n8601_));
  XOR2X1   g07599(.A(new_n8601_), .B(new_n8599_), .Y(new_n8602_));
  XOR2X1   g07600(.A(new_n8602_), .B(new_n8596_), .Y(new_n8603_));
  INVX1    g07601(.A(\A[451] ), .Y(new_n8604_));
  AND2X1   g07602(.A(\A[452] ), .B(new_n8604_), .Y(new_n8605_));
  OAI21X1  g07603(.A0(\A[452] ), .A1(new_n8604_), .B0(\A[453] ), .Y(new_n8606_));
  NAND2X1  g07604(.A(new_n8588_), .B(new_n8584_), .Y(new_n8607_));
  OAI21X1  g07605(.A0(new_n8606_), .A1(new_n8605_), .B0(new_n8607_), .Y(new_n8608_));
  XOR2X1   g07606(.A(new_n8595_), .B(new_n8608_), .Y(new_n8609_));
  NOR2X1   g07607(.A(new_n8595_), .B(new_n8589_), .Y(new_n8610_));
  AOI21X1  g07608(.A0(new_n8594_), .A1(\A[456] ), .B0(new_n8597_), .Y(new_n8611_));
  XOR2X1   g07609(.A(new_n8601_), .B(new_n8611_), .Y(new_n8612_));
  NOR2X1   g07610(.A(new_n8601_), .B(new_n8611_), .Y(new_n8613_));
  AOI21X1  g07611(.A0(new_n8612_), .A1(new_n8610_), .B0(new_n8613_), .Y(new_n8614_));
  OAI21X1  g07612(.A0(new_n8614_), .A1(new_n8609_), .B0(new_n8603_), .Y(new_n8615_));
  AND2X1   g07613(.A(\A[461] ), .B(\A[460] ), .Y(new_n8616_));
  XOR2X1   g07614(.A(\A[461] ), .B(\A[460] ), .Y(new_n8617_));
  AOI21X1  g07615(.A0(new_n8617_), .A1(\A[462] ), .B0(new_n8616_), .Y(new_n8618_));
  AND2X1   g07616(.A(\A[458] ), .B(\A[457] ), .Y(new_n8619_));
  XOR2X1   g07617(.A(\A[458] ), .B(\A[457] ), .Y(new_n8620_));
  AOI21X1  g07618(.A0(new_n8620_), .A1(\A[459] ), .B0(new_n8619_), .Y(new_n8621_));
  INVX1    g07619(.A(\A[459] ), .Y(new_n8622_));
  INVX1    g07620(.A(\A[458] ), .Y(new_n8623_));
  OR2X1    g07621(.A(new_n8623_), .B(\A[457] ), .Y(new_n8624_));
  AOI21X1  g07622(.A0(new_n8623_), .A1(\A[457] ), .B0(new_n8622_), .Y(new_n8625_));
  AOI22X1  g07623(.A0(new_n8625_), .A1(new_n8624_), .B0(new_n8620_), .B1(new_n8622_), .Y(new_n8626_));
  INVX1    g07624(.A(\A[462] ), .Y(new_n8627_));
  INVX1    g07625(.A(\A[461] ), .Y(new_n8628_));
  OR2X1    g07626(.A(new_n8628_), .B(\A[460] ), .Y(new_n8629_));
  AOI21X1  g07627(.A0(new_n8628_), .A1(\A[460] ), .B0(new_n8627_), .Y(new_n8630_));
  AOI22X1  g07628(.A0(new_n8630_), .A1(new_n8629_), .B0(new_n8617_), .B1(new_n8627_), .Y(new_n8631_));
  NOR4X1   g07629(.A(new_n8631_), .B(new_n8626_), .C(new_n8621_), .D(new_n8618_), .Y(new_n8632_));
  NOR4X1   g07630(.A(new_n8601_), .B(new_n8611_), .C(new_n8595_), .D(new_n8589_), .Y(new_n8633_));
  INVX1    g07631(.A(\A[457] ), .Y(new_n8634_));
  AND2X1   g07632(.A(\A[458] ), .B(new_n8634_), .Y(new_n8635_));
  OAI21X1  g07633(.A0(\A[458] ), .A1(new_n8634_), .B0(\A[459] ), .Y(new_n8636_));
  NAND2X1  g07634(.A(new_n8620_), .B(new_n8622_), .Y(new_n8637_));
  OAI21X1  g07635(.A0(new_n8636_), .A1(new_n8635_), .B0(new_n8637_), .Y(new_n8638_));
  XOR2X1   g07636(.A(new_n8631_), .B(new_n8638_), .Y(new_n8639_));
  OR4X1    g07637(.A(new_n8639_), .B(new_n8633_), .C(new_n8632_), .D(new_n8609_), .Y(new_n8640_));
  XOR2X1   g07638(.A(new_n8621_), .B(new_n8618_), .Y(new_n8641_));
  NOR2X1   g07639(.A(new_n8631_), .B(new_n8626_), .Y(new_n8642_));
  NOR2X1   g07640(.A(new_n8621_), .B(new_n8618_), .Y(new_n8643_));
  AOI21X1  g07641(.A0(new_n8642_), .A1(new_n8641_), .B0(new_n8643_), .Y(new_n8644_));
  XOR2X1   g07642(.A(new_n8642_), .B(new_n8641_), .Y(new_n8645_));
  OAI21X1  g07643(.A0(new_n8639_), .A1(new_n8644_), .B0(new_n8645_), .Y(new_n8646_));
  XOR2X1   g07644(.A(new_n8646_), .B(new_n8640_), .Y(new_n8647_));
  AND2X1   g07645(.A(new_n8647_), .B(new_n8615_), .Y(new_n8648_));
  OR2X1    g07646(.A(new_n8639_), .B(new_n8632_), .Y(new_n8649_));
  XOR2X1   g07647(.A(new_n8595_), .B(new_n8589_), .Y(new_n8650_));
  XOR2X1   g07648(.A(new_n8650_), .B(new_n8649_), .Y(new_n8651_));
  OR2X1    g07649(.A(new_n8562_), .B(new_n8555_), .Y(new_n8652_));
  XOR2X1   g07650(.A(new_n8518_), .B(new_n8512_), .Y(new_n8653_));
  XOR2X1   g07651(.A(new_n8653_), .B(new_n8652_), .Y(new_n8654_));
  NOR2X1   g07652(.A(new_n8654_), .B(new_n8651_), .Y(new_n8655_));
  AND2X1   g07653(.A(new_n8617_), .B(\A[462] ), .Y(new_n8656_));
  OR2X1    g07654(.A(new_n8656_), .B(new_n8616_), .Y(new_n8657_));
  XOR2X1   g07655(.A(new_n8621_), .B(new_n8657_), .Y(new_n8658_));
  XOR2X1   g07656(.A(new_n8642_), .B(new_n8658_), .Y(new_n8659_));
  NOR4X1   g07657(.A(new_n8639_), .B(new_n8633_), .C(new_n8659_), .D(new_n8609_), .Y(new_n8660_));
  OR2X1    g07658(.A(new_n8631_), .B(new_n8626_), .Y(new_n8661_));
  OR2X1    g07659(.A(new_n8621_), .B(new_n8618_), .Y(new_n8662_));
  OAI21X1  g07660(.A0(new_n8661_), .A1(new_n8658_), .B0(new_n8662_), .Y(new_n8663_));
  XOR2X1   g07661(.A(new_n8631_), .B(new_n8626_), .Y(new_n8664_));
  OAI21X1  g07662(.A0(new_n8664_), .A1(new_n8645_), .B0(new_n8663_), .Y(new_n8665_));
  AOI22X1  g07663(.A0(new_n8665_), .A1(new_n8660_), .B0(new_n8646_), .B1(new_n8640_), .Y(new_n8666_));
  OAI21X1  g07664(.A0(new_n8666_), .A1(new_n8615_), .B0(new_n8655_), .Y(new_n8667_));
  AOI21X1  g07665(.A0(new_n8664_), .A1(new_n8663_), .B0(new_n8659_), .Y(new_n8668_));
  XOR2X1   g07666(.A(new_n8668_), .B(new_n8640_), .Y(new_n8669_));
  MX2X1    g07667(.A(new_n8666_), .B(new_n8669_), .S0(new_n8615_), .Y(new_n8670_));
  OAI22X1  g07668(.A0(new_n8670_), .A1(new_n8655_), .B0(new_n8667_), .B1(new_n8648_), .Y(new_n8671_));
  AND2X1   g07669(.A(new_n8671_), .B(new_n8583_), .Y(new_n8672_));
  XOR2X1   g07670(.A(new_n8595_), .B(new_n8608_), .Y(new_n8673_));
  XOR2X1   g07671(.A(new_n8673_), .B(new_n8649_), .Y(new_n8674_));
  XOR2X1   g07672(.A(new_n8654_), .B(new_n8674_), .Y(new_n8675_));
  INVX1    g07673(.A(new_n8441_), .Y(new_n8676_));
  XOR2X1   g07674(.A(new_n8676_), .B(new_n8405_), .Y(new_n8677_));
  NOR2X1   g07675(.A(new_n8677_), .B(new_n8675_), .Y(new_n8678_));
  NAND2X1  g07676(.A(new_n8647_), .B(new_n8615_), .Y(new_n8679_));
  NOR4X1   g07677(.A(new_n8639_), .B(new_n8633_), .C(new_n8632_), .D(new_n8609_), .Y(new_n8680_));
  OR4X1    g07678(.A(new_n8639_), .B(new_n8633_), .C(new_n8659_), .D(new_n8609_), .Y(new_n8681_));
  AOI21X1  g07679(.A0(new_n8639_), .A1(new_n8659_), .B0(new_n8644_), .Y(new_n8682_));
  OAI22X1  g07680(.A0(new_n8682_), .A1(new_n8681_), .B0(new_n8668_), .B1(new_n8680_), .Y(new_n8683_));
  MX2X1    g07681(.A(new_n8683_), .B(new_n8647_), .S0(new_n8615_), .Y(new_n8684_));
  XOR2X1   g07682(.A(new_n8602_), .B(new_n8610_), .Y(new_n8685_));
  XOR2X1   g07683(.A(new_n8595_), .B(new_n8589_), .Y(new_n8686_));
  OR2X1    g07684(.A(new_n8601_), .B(new_n8611_), .Y(new_n8687_));
  OAI21X1  g07685(.A0(new_n8602_), .A1(new_n8596_), .B0(new_n8687_), .Y(new_n8688_));
  AOI21X1  g07686(.A0(new_n8688_), .A1(new_n8686_), .B0(new_n8685_), .Y(new_n8689_));
  AOI21X1  g07687(.A0(new_n8683_), .A1(new_n8689_), .B0(new_n8655_), .Y(new_n8690_));
  AOI22X1  g07688(.A0(new_n8690_), .A1(new_n8679_), .B0(new_n8684_), .B1(new_n8655_), .Y(new_n8691_));
  OAI21X1  g07689(.A0(new_n8691_), .A1(new_n8583_), .B0(new_n8678_), .Y(new_n8692_));
  NOR4X1   g07690(.A(new_n8562_), .B(new_n8556_), .C(new_n8555_), .D(new_n8532_), .Y(new_n8693_));
  XOR2X1   g07691(.A(new_n8573_), .B(new_n8693_), .Y(new_n8694_));
  OR4X1    g07692(.A(new_n8562_), .B(new_n8556_), .C(new_n8571_), .D(new_n8532_), .Y(new_n8695_));
  AOI21X1  g07693(.A0(new_n8562_), .A1(new_n8571_), .B0(new_n8577_), .Y(new_n8696_));
  OAI22X1  g07694(.A0(new_n8696_), .A1(new_n8695_), .B0(new_n8573_), .B1(new_n8693_), .Y(new_n8697_));
  MX2X1    g07695(.A(new_n8697_), .B(new_n8694_), .S0(new_n8538_), .Y(new_n8698_));
  OR2X1    g07696(.A(new_n8654_), .B(new_n8651_), .Y(new_n8699_));
  AOI21X1  g07697(.A0(new_n8683_), .A1(new_n8689_), .B0(new_n8699_), .Y(new_n8700_));
  AOI22X1  g07698(.A0(new_n8684_), .A1(new_n8699_), .B0(new_n8700_), .B1(new_n8679_), .Y(new_n8701_));
  MX2X1    g07699(.A(new_n8701_), .B(new_n8691_), .S0(new_n8698_), .Y(new_n8702_));
  OAI22X1  g07700(.A0(new_n8702_), .A1(new_n8678_), .B0(new_n8692_), .B1(new_n8672_), .Y(new_n8703_));
  AND2X1   g07701(.A(new_n8703_), .B(new_n8506_), .Y(new_n8704_));
  XOR2X1   g07702(.A(new_n8677_), .B(new_n8675_), .Y(new_n8705_));
  INVX1    g07703(.A(new_n8705_), .Y(new_n8706_));
  XOR2X1   g07704(.A(new_n8215_), .B(new_n8178_), .Y(new_n8707_));
  XOR2X1   g07705(.A(new_n8707_), .B(new_n8142_), .Y(new_n8708_));
  NOR2X1   g07706(.A(new_n8708_), .B(new_n8706_), .Y(new_n8709_));
  OR2X1    g07707(.A(new_n8701_), .B(new_n8698_), .Y(new_n8710_));
  OAI21X1  g07708(.A0(new_n8666_), .A1(new_n8615_), .B0(new_n8699_), .Y(new_n8711_));
  OAI22X1  g07709(.A0(new_n8711_), .A1(new_n8648_), .B0(new_n8670_), .B1(new_n8699_), .Y(new_n8712_));
  MX2X1    g07710(.A(new_n8671_), .B(new_n8712_), .S0(new_n8698_), .Y(new_n8713_));
  AOI21X1  g07711(.A0(new_n8712_), .A1(new_n8698_), .B0(new_n8678_), .Y(new_n8714_));
  AOI22X1  g07712(.A0(new_n8714_), .A1(new_n8710_), .B0(new_n8713_), .B1(new_n8678_), .Y(new_n8715_));
  OAI21X1  g07713(.A0(new_n8715_), .A1(new_n8506_), .B0(new_n8709_), .Y(new_n8716_));
  OR2X1    g07714(.A(new_n8677_), .B(new_n8675_), .Y(new_n8717_));
  AOI21X1  g07715(.A0(new_n8712_), .A1(new_n8698_), .B0(new_n8717_), .Y(new_n8718_));
  AOI22X1  g07716(.A0(new_n8713_), .A1(new_n8717_), .B0(new_n8718_), .B1(new_n8710_), .Y(new_n8719_));
  MX2X1    g07717(.A(new_n8715_), .B(new_n8719_), .S0(new_n8506_), .Y(new_n8720_));
  OAI22X1  g07718(.A0(new_n8720_), .A1(new_n8709_), .B0(new_n8716_), .B1(new_n8704_), .Y(new_n8721_));
  AND2X1   g07719(.A(new_n8721_), .B(new_n8333_), .Y(new_n8722_));
  OR4X1    g07720(.A(new_n8026_), .B(new_n8020_), .C(new_n8019_), .D(new_n7996_), .Y(new_n8723_));
  XOR2X1   g07721(.A(new_n8037_), .B(new_n8723_), .Y(new_n8724_));
  XOR2X1   g07722(.A(new_n8034_), .B(new_n8040_), .Y(new_n8725_));
  OAI21X1  g07723(.A0(new_n8026_), .A1(new_n8042_), .B0(new_n8725_), .Y(new_n8726_));
  NOR4X1   g07724(.A(new_n8026_), .B(new_n8020_), .C(new_n8035_), .D(new_n7996_), .Y(new_n8727_));
  OAI21X1  g07725(.A0(new_n8036_), .A1(new_n8725_), .B0(new_n8033_), .Y(new_n8728_));
  AOI22X1  g07726(.A0(new_n8728_), .A1(new_n8727_), .B0(new_n8726_), .B1(new_n8723_), .Y(new_n8729_));
  MX2X1    g07727(.A(new_n8729_), .B(new_n8724_), .S0(new_n8002_), .Y(new_n8730_));
  AND2X1   g07728(.A(new_n8229_), .B(new_n8730_), .Y(new_n8731_));
  AOI21X1  g07729(.A0(new_n8135_), .A1(new_n8122_), .B0(new_n8227_), .Y(new_n8732_));
  AOI22X1  g07730(.A0(new_n8732_), .A1(new_n8110_), .B0(new_n8137_), .B1(new_n8227_), .Y(new_n8733_));
  OAI21X1  g07731(.A0(new_n8733_), .A1(new_n8730_), .B0(new_n8330_), .Y(new_n8734_));
  MX2X1    g07732(.A(new_n8138_), .B(new_n8733_), .S0(new_n8045_), .Y(new_n8735_));
  OAI22X1  g07733(.A0(new_n8735_), .A1(new_n8330_), .B0(new_n8734_), .B1(new_n8731_), .Y(new_n8736_));
  OAI21X1  g07734(.A0(new_n8733_), .A1(new_n8730_), .B0(new_n8217_), .Y(new_n8737_));
  OAI22X1  g07735(.A0(new_n8737_), .A1(new_n8731_), .B0(new_n8735_), .B1(new_n8217_), .Y(new_n8738_));
  MX2X1    g07736(.A(new_n8738_), .B(new_n8736_), .S0(new_n8329_), .Y(new_n8739_));
  OR2X1    g07737(.A(new_n8708_), .B(new_n8706_), .Y(new_n8740_));
  OAI21X1  g07738(.A0(new_n8715_), .A1(new_n8506_), .B0(new_n8740_), .Y(new_n8741_));
  OAI22X1  g07739(.A0(new_n8741_), .A1(new_n8704_), .B0(new_n8720_), .B1(new_n8740_), .Y(new_n8742_));
  AND2X1   g07740(.A(new_n8742_), .B(new_n8739_), .Y(new_n8743_));
  XOR2X1   g07741(.A(new_n8708_), .B(new_n8705_), .Y(new_n8744_));
  XOR2X1   g07742(.A(new_n7730_), .B(new_n7581_), .Y(new_n8745_));
  OR4X1    g07743(.A(new_n8745_), .B(new_n8744_), .C(new_n8743_), .D(new_n8722_), .Y(new_n8746_));
  NOR2X1   g07744(.A(new_n8745_), .B(new_n8744_), .Y(new_n8747_));
  AND2X1   g07745(.A(new_n8397_), .B(new_n8365_), .Y(new_n8748_));
  NOR4X1   g07746(.A(new_n8389_), .B(new_n8383_), .C(new_n8455_), .D(new_n8359_), .Y(new_n8749_));
  OAI21X1  g07747(.A0(new_n8402_), .A1(new_n8395_), .B0(new_n8454_), .Y(new_n8750_));
  AOI22X1  g07748(.A0(new_n8750_), .A1(new_n8749_), .B0(new_n8396_), .B1(new_n8390_), .Y(new_n8751_));
  OAI21X1  g07749(.A0(new_n8751_), .A1(new_n8365_), .B0(new_n8503_), .Y(new_n8752_));
  XOR2X1   g07750(.A(new_n8456_), .B(new_n8390_), .Y(new_n8753_));
  MX2X1    g07751(.A(new_n8751_), .B(new_n8753_), .S0(new_n8365_), .Y(new_n8754_));
  OAI22X1  g07752(.A0(new_n8754_), .A1(new_n8503_), .B0(new_n8752_), .B1(new_n8748_), .Y(new_n8755_));
  OAI21X1  g07753(.A0(new_n8751_), .A1(new_n8365_), .B0(new_n8442_), .Y(new_n8756_));
  OAI22X1  g07754(.A0(new_n8756_), .A1(new_n8748_), .B0(new_n8754_), .B1(new_n8442_), .Y(new_n8757_));
  MX2X1    g07755(.A(new_n8757_), .B(new_n8755_), .S0(new_n8502_), .Y(new_n8758_));
  OR2X1    g07756(.A(new_n8719_), .B(new_n8758_), .Y(new_n8759_));
  OAI21X1  g07757(.A0(new_n8691_), .A1(new_n8583_), .B0(new_n8717_), .Y(new_n8760_));
  OAI22X1  g07758(.A0(new_n8760_), .A1(new_n8672_), .B0(new_n8702_), .B1(new_n8717_), .Y(new_n8761_));
  AOI21X1  g07759(.A0(new_n8761_), .A1(new_n8758_), .B0(new_n8740_), .Y(new_n8762_));
  MX2X1    g07760(.A(new_n8761_), .B(new_n8703_), .S0(new_n8506_), .Y(new_n8763_));
  AOI22X1  g07761(.A0(new_n8763_), .A1(new_n8740_), .B0(new_n8762_), .B1(new_n8759_), .Y(new_n8764_));
  AOI21X1  g07762(.A0(new_n8761_), .A1(new_n8758_), .B0(new_n8709_), .Y(new_n8765_));
  AOI22X1  g07763(.A0(new_n8765_), .A1(new_n8759_), .B0(new_n8763_), .B1(new_n8709_), .Y(new_n8766_));
  MX2X1    g07764(.A(new_n8766_), .B(new_n8764_), .S0(new_n8333_), .Y(new_n8767_));
  OR2X1    g07765(.A(new_n8767_), .B(new_n8747_), .Y(new_n8768_));
  AOI21X1  g07766(.A0(new_n8768_), .A1(new_n8746_), .B0(new_n7970_), .Y(new_n8769_));
  INVX1    g07767(.A(new_n8747_), .Y(new_n8770_));
  OAI21X1  g07768(.A0(new_n8766_), .A1(new_n8333_), .B0(new_n8770_), .Y(new_n8771_));
  OAI22X1  g07769(.A0(new_n8771_), .A1(new_n8722_), .B0(new_n8767_), .B1(new_n8770_), .Y(new_n8772_));
  AND2X1   g07770(.A(new_n8772_), .B(new_n7970_), .Y(new_n8773_));
  INVX1    g07771(.A(new_n8744_), .Y(new_n8774_));
  XOR2X1   g07772(.A(new_n8745_), .B(new_n8774_), .Y(new_n8775_));
  XOR2X1   g07773(.A(new_n6947_), .B(new_n6562_), .Y(new_n8776_));
  XOR2X1   g07774(.A(new_n8776_), .B(new_n6414_), .Y(new_n8777_));
  NOR2X1   g07775(.A(new_n8777_), .B(new_n8775_), .Y(new_n8778_));
  INVX1    g07776(.A(new_n8778_), .Y(new_n8779_));
  NOR3X1   g07777(.A(new_n8779_), .B(new_n8773_), .C(new_n8769_), .Y(new_n8780_));
  AND2X1   g07778(.A(new_n7273_), .B(new_n7241_), .Y(new_n8781_));
  NOR4X1   g07779(.A(new_n7265_), .B(new_n7259_), .C(new_n7331_), .D(new_n7235_), .Y(new_n8782_));
  OAI21X1  g07780(.A0(new_n7278_), .A1(new_n7271_), .B0(new_n7330_), .Y(new_n8783_));
  AOI22X1  g07781(.A0(new_n8783_), .A1(new_n8782_), .B0(new_n7272_), .B1(new_n7266_), .Y(new_n8784_));
  OAI21X1  g07782(.A0(new_n8784_), .A1(new_n7241_), .B0(new_n7379_), .Y(new_n8785_));
  XOR2X1   g07783(.A(new_n7332_), .B(new_n7266_), .Y(new_n8786_));
  MX2X1    g07784(.A(new_n8784_), .B(new_n8786_), .S0(new_n7241_), .Y(new_n8787_));
  OAI22X1  g07785(.A0(new_n8787_), .A1(new_n7379_), .B0(new_n8785_), .B1(new_n8781_), .Y(new_n8788_));
  OAI21X1  g07786(.A0(new_n8784_), .A1(new_n7241_), .B0(new_n7318_), .Y(new_n8789_));
  OAI22X1  g07787(.A0(new_n8789_), .A1(new_n8781_), .B0(new_n8787_), .B1(new_n7318_), .Y(new_n8790_));
  MX2X1    g07788(.A(new_n8790_), .B(new_n8788_), .S0(new_n7378_), .Y(new_n8791_));
  OR2X1    g07789(.A(new_n7741_), .B(new_n8791_), .Y(new_n8792_));
  OAI21X1  g07790(.A0(new_n7567_), .A1(new_n7459_), .B0(new_n7739_), .Y(new_n8793_));
  OAI22X1  g07791(.A0(new_n8793_), .A1(new_n7548_), .B0(new_n7578_), .B1(new_n7739_), .Y(new_n8794_));
  AOI21X1  g07792(.A0(new_n8794_), .A1(new_n8791_), .B0(new_n7967_), .Y(new_n8795_));
  MX2X1    g07793(.A(new_n8794_), .B(new_n7579_), .S0(new_n7382_), .Y(new_n8796_));
  AOI22X1  g07794(.A0(new_n8796_), .A1(new_n7967_), .B0(new_n8795_), .B1(new_n8792_), .Y(new_n8797_));
  AOI21X1  g07795(.A0(new_n8794_), .A1(new_n8791_), .B0(new_n7731_), .Y(new_n8798_));
  AOI22X1  g07796(.A0(new_n8798_), .A1(new_n8792_), .B0(new_n8796_), .B1(new_n7731_), .Y(new_n8799_));
  MX2X1    g07797(.A(new_n8799_), .B(new_n8797_), .S0(new_n7966_), .Y(new_n8800_));
  NOR3X1   g07798(.A(new_n8770_), .B(new_n8743_), .C(new_n8722_), .Y(new_n8801_));
  MX2X1    g07799(.A(new_n8742_), .B(new_n8721_), .S0(new_n8333_), .Y(new_n8802_));
  AND2X1   g07800(.A(new_n8802_), .B(new_n8770_), .Y(new_n8803_));
  OAI21X1  g07801(.A0(new_n8803_), .A1(new_n8801_), .B0(new_n8800_), .Y(new_n8804_));
  OR2X1    g07802(.A(new_n8764_), .B(new_n8739_), .Y(new_n8805_));
  AOI21X1  g07803(.A0(new_n8742_), .A1(new_n8739_), .B0(new_n8747_), .Y(new_n8806_));
  AOI22X1  g07804(.A0(new_n8806_), .A1(new_n8805_), .B0(new_n8802_), .B1(new_n8747_), .Y(new_n8807_));
  OR2X1    g07805(.A(new_n8807_), .B(new_n8800_), .Y(new_n8808_));
  AOI21X1  g07806(.A0(new_n8808_), .A1(new_n8804_), .B0(new_n8778_), .Y(new_n8809_));
  OAI21X1  g07807(.A0(new_n8809_), .A1(new_n8780_), .B0(new_n7209_), .Y(new_n8810_));
  AND2X1   g07808(.A(new_n6733_), .B(new_n6730_), .Y(new_n8811_));
  AOI21X1  g07809(.A0(new_n6390_), .A1(new_n6181_), .B0(new_n6731_), .Y(new_n8812_));
  AOI22X1  g07810(.A0(new_n8812_), .A1(new_n6371_), .B0(new_n6411_), .B1(new_n6731_), .Y(new_n8813_));
  OAI21X1  g07811(.A0(new_n8813_), .A1(new_n6730_), .B0(new_n6713_), .Y(new_n8814_));
  MX2X1    g07812(.A(new_n8813_), .B(new_n6412_), .S0(new_n6730_), .Y(new_n8815_));
  OAI22X1  g07813(.A0(new_n8815_), .A1(new_n6713_), .B0(new_n8814_), .B1(new_n8811_), .Y(new_n8816_));
  OAI21X1  g07814(.A0(new_n8813_), .A1(new_n6730_), .B0(new_n6714_), .Y(new_n8817_));
  OAI22X1  g07815(.A0(new_n8817_), .A1(new_n8811_), .B0(new_n8815_), .B1(new_n6714_), .Y(new_n8818_));
  MX2X1    g07816(.A(new_n8818_), .B(new_n8816_), .S0(new_n7206_), .Y(new_n8819_));
  AOI21X1  g07817(.A0(new_n8772_), .A1(new_n7970_), .B0(new_n8778_), .Y(new_n8820_));
  AND2X1   g07818(.A(new_n8820_), .B(new_n8804_), .Y(new_n8821_));
  AOI21X1  g07819(.A0(new_n8808_), .A1(new_n8804_), .B0(new_n8779_), .Y(new_n8822_));
  OAI21X1  g07820(.A0(new_n8822_), .A1(new_n8821_), .B0(new_n8819_), .Y(new_n8823_));
  XOR2X1   g07821(.A(new_n8777_), .B(new_n8775_), .Y(new_n8824_));
  INVX1    g07822(.A(new_n8824_), .Y(new_n8825_));
  AOI21X1  g07823(.A0(new_n4926_), .A1(new_n4924_), .B0(new_n5236_), .Y(new_n8826_));
  AND2X1   g07824(.A(new_n5236_), .B(new_n4924_), .Y(new_n8827_));
  AOI21X1  g07825(.A0(new_n8827_), .A1(new_n4926_), .B0(new_n8826_), .Y(new_n8828_));
  NOR2X1   g07826(.A(new_n8828_), .B(new_n8825_), .Y(new_n8829_));
  NAND3X1  g07827(.A(new_n8829_), .B(new_n8823_), .C(new_n8810_), .Y(new_n8830_));
  NAND3X1  g07828(.A(new_n8778_), .B(new_n8808_), .C(new_n8804_), .Y(new_n8831_));
  OAI21X1  g07829(.A0(new_n8773_), .A1(new_n8769_), .B0(new_n8779_), .Y(new_n8832_));
  AOI21X1  g07830(.A0(new_n8832_), .A1(new_n8831_), .B0(new_n8819_), .Y(new_n8833_));
  OAI21X1  g07831(.A0(new_n8807_), .A1(new_n8800_), .B0(new_n8779_), .Y(new_n8834_));
  OR2X1    g07832(.A(new_n8834_), .B(new_n8769_), .Y(new_n8835_));
  OAI21X1  g07833(.A0(new_n8773_), .A1(new_n8769_), .B0(new_n8778_), .Y(new_n8836_));
  AOI21X1  g07834(.A0(new_n8836_), .A1(new_n8835_), .B0(new_n7209_), .Y(new_n8837_));
  INVX1    g07835(.A(new_n8829_), .Y(new_n8838_));
  OAI21X1  g07836(.A0(new_n8837_), .A1(new_n8833_), .B0(new_n8838_), .Y(new_n8839_));
  AOI21X1  g07837(.A0(new_n8839_), .A1(new_n8830_), .B0(new_n5642_), .Y(new_n8840_));
  AND2X1   g07838(.A(new_n5641_), .B(new_n5630_), .Y(new_n8841_));
  NAND3X1  g07839(.A(new_n8838_), .B(new_n8823_), .C(new_n8810_), .Y(new_n8842_));
  OAI21X1  g07840(.A0(new_n8837_), .A1(new_n8833_), .B0(new_n8829_), .Y(new_n8843_));
  AOI21X1  g07841(.A0(new_n8843_), .A1(new_n8842_), .B0(new_n8841_), .Y(new_n8844_));
  XOR2X1   g07842(.A(new_n3042_), .B(new_n3041_), .Y(new_n8845_));
  XOR2X1   g07843(.A(new_n8828_), .B(new_n8824_), .Y(new_n8846_));
  NOR2X1   g07844(.A(new_n8846_), .B(new_n8845_), .Y(new_n8847_));
  NOR3X1   g07845(.A(new_n8847_), .B(new_n8844_), .C(new_n8840_), .Y(new_n8848_));
  OAI21X1  g07846(.A0(new_n8844_), .A1(new_n8840_), .B0(new_n8847_), .Y(new_n8849_));
  OAI21X1  g07847(.A0(new_n8848_), .A1(new_n3849_), .B0(new_n8849_), .Y(new_n8850_));
  NOR3X1   g07848(.A(new_n8829_), .B(new_n8837_), .C(new_n8833_), .Y(new_n8851_));
  OAI21X1  g07849(.A0(new_n8851_), .A1(new_n8841_), .B0(new_n8843_), .Y(new_n8852_));
  AOI21X1  g07850(.A0(new_n5638_), .A1(new_n5243_), .B0(new_n5629_), .Y(new_n8853_));
  OR2X1    g07851(.A(new_n8853_), .B(new_n5640_), .Y(new_n8854_));
  OR2X1    g07852(.A(new_n4917_), .B(new_n4920_), .Y(new_n8855_));
  OAI21X1  g07853(.A0(new_n4921_), .A1(new_n4878_), .B0(new_n4186_), .Y(new_n8856_));
  AND2X1   g07854(.A(new_n8856_), .B(new_n8855_), .Y(new_n8857_));
  AND2X1   g07855(.A(new_n4913_), .B(new_n4865_), .Y(new_n8858_));
  AOI21X1  g07856(.A0(new_n4915_), .A1(new_n4909_), .B0(new_n4483_), .Y(new_n8859_));
  OR2X1    g07857(.A(new_n8859_), .B(new_n8858_), .Y(new_n8860_));
  OR2X1    g07858(.A(new_n4884_), .B(new_n4423_), .Y(new_n8861_));
  OAI21X1  g07859(.A0(new_n4886_), .A1(new_n4880_), .B0(new_n4479_), .Y(new_n8862_));
  AND2X1   g07860(.A(new_n8862_), .B(new_n8861_), .Y(new_n8863_));
  OR2X1    g07861(.A(new_n4474_), .B(new_n4476_), .Y(new_n8864_));
  INVX1    g07862(.A(new_n4445_), .Y(new_n8865_));
  OAI21X1  g07863(.A0(new_n4477_), .A1(new_n4463_), .B0(new_n8865_), .Y(new_n8866_));
  NOR2X1   g07864(.A(new_n4465_), .B(new_n4459_), .Y(new_n8867_));
  AOI21X1  g07865(.A0(new_n4465_), .A1(new_n4459_), .B0(new_n4447_), .Y(new_n8868_));
  NOR2X1   g07866(.A(new_n4453_), .B(new_n4451_), .Y(new_n8869_));
  AOI21X1  g07867(.A0(new_n4471_), .A1(new_n4454_), .B0(new_n8869_), .Y(new_n8870_));
  OAI21X1  g07868(.A0(new_n8868_), .A1(new_n8867_), .B0(new_n8870_), .Y(new_n8871_));
  OR2X1    g07869(.A(new_n4465_), .B(new_n4459_), .Y(new_n8872_));
  OAI21X1  g07870(.A0(new_n4461_), .A1(new_n4472_), .B0(new_n4448_), .Y(new_n8873_));
  INVX1    g07871(.A(new_n8869_), .Y(new_n8874_));
  OAI21X1  g07872(.A0(new_n4458_), .A1(new_n4455_), .B0(new_n8874_), .Y(new_n8875_));
  NAND3X1  g07873(.A(new_n8875_), .B(new_n8873_), .C(new_n8872_), .Y(new_n8876_));
  INVX1    g07874(.A(new_n4439_), .Y(new_n8877_));
  AOI21X1  g07875(.A0(new_n4444_), .A1(new_n8877_), .B0(new_n4443_), .Y(new_n8878_));
  NAND3X1  g07876(.A(new_n8878_), .B(new_n8876_), .C(new_n8871_), .Y(new_n8879_));
  AOI21X1  g07877(.A0(new_n8873_), .A1(new_n8872_), .B0(new_n8875_), .Y(new_n8880_));
  NOR3X1   g07878(.A(new_n8870_), .B(new_n8868_), .C(new_n8867_), .Y(new_n8881_));
  AND2X1   g07879(.A(new_n4444_), .B(new_n8877_), .Y(new_n8882_));
  OR2X1    g07880(.A(new_n8882_), .B(new_n4443_), .Y(new_n8883_));
  OAI21X1  g07881(.A0(new_n8881_), .A1(new_n8880_), .B0(new_n8883_), .Y(new_n8884_));
  AOI22X1  g07882(.A0(new_n8884_), .A1(new_n8879_), .B0(new_n8866_), .B1(new_n8864_), .Y(new_n8885_));
  XOR2X1   g07883(.A(new_n4465_), .B(new_n4459_), .Y(new_n8886_));
  OAI22X1  g07884(.A0(new_n4467_), .A1(new_n4466_), .B0(new_n8886_), .B1(new_n4447_), .Y(new_n8887_));
  AND2X1   g07885(.A(new_n8887_), .B(new_n4464_), .Y(new_n8888_));
  OR2X1    g07886(.A(new_n8886_), .B(new_n4447_), .Y(new_n8889_));
  AOI21X1  g07887(.A0(new_n4473_), .A1(new_n4469_), .B0(new_n4464_), .Y(new_n8890_));
  AOI21X1  g07888(.A0(new_n8890_), .A1(new_n8889_), .B0(new_n4445_), .Y(new_n8891_));
  NOR3X1   g07889(.A(new_n8883_), .B(new_n8881_), .C(new_n8880_), .Y(new_n8892_));
  AOI21X1  g07890(.A0(new_n8876_), .A1(new_n8871_), .B0(new_n8878_), .Y(new_n8893_));
  NOR4X1   g07891(.A(new_n8893_), .B(new_n8892_), .C(new_n8891_), .D(new_n8888_), .Y(new_n8894_));
  OR2X1    g07892(.A(new_n8894_), .B(new_n8885_), .Y(new_n8895_));
  AND2X1   g07893(.A(new_n4361_), .B(new_n4433_), .Y(new_n8896_));
  AOI21X1  g07894(.A0(new_n4881_), .A1(new_n4334_), .B0(new_n4879_), .Y(new_n8897_));
  NOR2X1   g07895(.A(new_n8897_), .B(new_n8896_), .Y(new_n8898_));
  OR4X1    g07896(.A(new_n4242_), .B(new_n4236_), .C(new_n4251_), .D(new_n4218_), .Y(new_n8899_));
  AOI21X1  g07897(.A0(new_n4242_), .A1(new_n4251_), .B0(new_n4262_), .Y(new_n8900_));
  OR2X1    g07898(.A(new_n8900_), .B(new_n8899_), .Y(new_n8901_));
  NOR4X1   g07899(.A(new_n4242_), .B(new_n4236_), .C(new_n4235_), .D(new_n4218_), .Y(new_n8902_));
  OAI21X1  g07900(.A0(new_n4253_), .A1(new_n8902_), .B0(new_n4212_), .Y(new_n8903_));
  OAI21X1  g07901(.A0(new_n4242_), .A1(new_n4251_), .B0(new_n4249_), .Y(new_n8904_));
  AOI21X1  g07902(.A0(new_n4207_), .A1(new_n4255_), .B0(new_n4258_), .Y(new_n8905_));
  XOR2X1   g07903(.A(new_n8905_), .B(new_n8904_), .Y(new_n8906_));
  AOI21X1  g07904(.A0(new_n8903_), .A1(new_n8901_), .B0(new_n8906_), .Y(new_n8907_));
  AOI21X1  g07905(.A0(new_n4264_), .A1(new_n4243_), .B0(new_n4259_), .Y(new_n8908_));
  NOR2X1   g07906(.A(new_n8905_), .B(new_n8904_), .Y(new_n8909_));
  AOI21X1  g07907(.A0(new_n4252_), .A1(new_n4263_), .B0(new_n4262_), .Y(new_n8910_));
  OAI21X1  g07908(.A0(new_n4218_), .A1(new_n4206_), .B0(new_n4211_), .Y(new_n8911_));
  OAI22X1  g07909(.A0(new_n8911_), .A1(new_n8910_), .B0(new_n8900_), .B1(new_n8899_), .Y(new_n8912_));
  NOR3X1   g07910(.A(new_n8912_), .B(new_n8909_), .C(new_n8908_), .Y(new_n8913_));
  OR2X1    g07911(.A(new_n8913_), .B(new_n8907_), .Y(new_n8914_));
  OR2X1    g07912(.A(new_n4358_), .B(new_n4357_), .Y(new_n8915_));
  OAI21X1  g07913(.A0(new_n4356_), .A1(new_n4347_), .B0(new_n4346_), .Y(new_n8916_));
  OAI21X1  g07914(.A0(new_n4325_), .A1(new_n4354_), .B0(new_n4353_), .Y(new_n8917_));
  AOI21X1  g07915(.A0(new_n4343_), .A1(new_n4289_), .B0(new_n4300_), .Y(new_n8918_));
  XOR2X1   g07916(.A(new_n8918_), .B(new_n8917_), .Y(new_n8919_));
  AOI21X1  g07917(.A0(new_n8916_), .A1(new_n8915_), .B0(new_n8919_), .Y(new_n8920_));
  AOI21X1  g07918(.A0(new_n4332_), .A1(new_n4326_), .B0(new_n4301_), .Y(new_n8921_));
  NOR2X1   g07919(.A(new_n8918_), .B(new_n8917_), .Y(new_n8922_));
  AOI21X1  g07920(.A0(new_n4355_), .A1(new_n4331_), .B0(new_n4330_), .Y(new_n8923_));
  OAI21X1  g07921(.A0(new_n4295_), .A1(new_n4342_), .B0(new_n4345_), .Y(new_n8924_));
  OAI22X1  g07922(.A0(new_n8924_), .A1(new_n8923_), .B0(new_n4358_), .B1(new_n4357_), .Y(new_n8925_));
  NOR3X1   g07923(.A(new_n8925_), .B(new_n8922_), .C(new_n8921_), .Y(new_n8926_));
  NOR2X1   g07924(.A(new_n8926_), .B(new_n8920_), .Y(new_n8927_));
  XOR2X1   g07925(.A(new_n8927_), .B(new_n8914_), .Y(new_n8928_));
  XOR2X1   g07926(.A(new_n8928_), .B(new_n8898_), .Y(new_n8929_));
  XOR2X1   g07927(.A(new_n8929_), .B(new_n8895_), .Y(new_n8930_));
  XOR2X1   g07928(.A(new_n8930_), .B(new_n8863_), .Y(new_n8931_));
  OR2X1    g07929(.A(new_n4852_), .B(new_n4873_), .Y(new_n8932_));
  OAI21X1  g07930(.A0(new_n4910_), .A1(new_n4822_), .B0(new_n4908_), .Y(new_n8933_));
  AND2X1   g07931(.A(new_n8933_), .B(new_n8932_), .Y(new_n8934_));
  OR2X1    g07932(.A(new_n4904_), .B(new_n4592_), .Y(new_n8935_));
  NOR4X1   g07933(.A(new_n4631_), .B(new_n4618_), .C(new_n4630_), .D(new_n4625_), .Y(new_n8936_));
  XOR2X1   g07934(.A(new_n4642_), .B(new_n8936_), .Y(new_n8937_));
  OR4X1    g07935(.A(new_n4618_), .B(new_n4630_), .C(new_n4641_), .D(new_n4625_), .Y(new_n8938_));
  AND2X1   g07936(.A(new_n4584_), .B(\A[36] ), .Y(new_n8939_));
  OR2X1    g07937(.A(new_n8939_), .B(new_n4586_), .Y(new_n8940_));
  XOR2X1   g07938(.A(new_n4589_), .B(new_n8940_), .Y(new_n8941_));
  XOR2X1   g07939(.A(new_n4620_), .B(new_n8941_), .Y(new_n8942_));
  OAI22X1  g07940(.A0(new_n8942_), .A1(new_n4622_), .B0(new_n4646_), .B1(new_n4625_), .Y(new_n8943_));
  OAI22X1  g07941(.A0(new_n8943_), .A1(new_n8938_), .B0(new_n4642_), .B1(new_n8936_), .Y(new_n8944_));
  MX2X1    g07942(.A(new_n8944_), .B(new_n8937_), .S0(new_n4624_), .Y(new_n8945_));
  OAI21X1  g07943(.A0(new_n4906_), .A1(new_n4898_), .B0(new_n8945_), .Y(new_n8946_));
  AND2X1   g07944(.A(new_n8946_), .B(new_n8935_), .Y(new_n8947_));
  OR2X1    g07945(.A(new_n8943_), .B(new_n8938_), .Y(new_n8948_));
  XOR2X1   g07946(.A(new_n4585_), .B(new_n4579_), .Y(new_n8949_));
  OR2X1    g07947(.A(new_n4585_), .B(new_n4579_), .Y(new_n8950_));
  OR2X1    g07948(.A(new_n4589_), .B(new_n4587_), .Y(new_n8951_));
  OAI21X1  g07949(.A0(new_n8950_), .A1(new_n8941_), .B0(new_n8951_), .Y(new_n8952_));
  AOI21X1  g07950(.A0(new_n8952_), .A1(new_n8949_), .B0(new_n8942_), .Y(new_n8953_));
  OAI21X1  g07951(.A0(new_n4642_), .A1(new_n8936_), .B0(new_n8953_), .Y(new_n8954_));
  OAI21X1  g07952(.A0(new_n4641_), .A1(new_n4625_), .B0(new_n4639_), .Y(new_n8955_));
  AOI21X1  g07953(.A0(new_n4623_), .A1(new_n8949_), .B0(new_n4622_), .Y(new_n8956_));
  XOR2X1   g07954(.A(new_n8956_), .B(new_n8955_), .Y(new_n8957_));
  AOI21X1  g07955(.A0(new_n8954_), .A1(new_n8948_), .B0(new_n8957_), .Y(new_n8958_));
  AOI21X1  g07956(.A0(new_n4648_), .A1(new_n4632_), .B0(new_n4624_), .Y(new_n8959_));
  NOR2X1   g07957(.A(new_n8956_), .B(new_n8955_), .Y(new_n8960_));
  AOI21X1  g07958(.A0(new_n4647_), .A1(new_n4633_), .B0(new_n4646_), .Y(new_n8961_));
  OAI21X1  g07959(.A0(new_n8942_), .A1(new_n4618_), .B0(new_n8952_), .Y(new_n8962_));
  OAI22X1  g07960(.A0(new_n8962_), .A1(new_n8961_), .B0(new_n8943_), .B1(new_n8938_), .Y(new_n8963_));
  NOR3X1   g07961(.A(new_n8963_), .B(new_n8960_), .C(new_n8959_), .Y(new_n8964_));
  NOR2X1   g07962(.A(new_n8964_), .B(new_n8958_), .Y(new_n8965_));
  OR2X1    g07963(.A(new_n4608_), .B(new_n4607_), .Y(new_n8966_));
  OAI21X1  g07964(.A0(new_n4606_), .A1(new_n4598_), .B0(new_n4597_), .Y(new_n8967_));
  OAI21X1  g07965(.A0(new_n4539_), .A1(new_n4605_), .B0(new_n4604_), .Y(new_n8968_));
  AOI21X1  g07966(.A0(new_n4594_), .A1(new_n4503_), .B0(new_n4514_), .Y(new_n8969_));
  XOR2X1   g07967(.A(new_n8969_), .B(new_n8968_), .Y(new_n8970_));
  AOI21X1  g07968(.A0(new_n8967_), .A1(new_n8966_), .B0(new_n8970_), .Y(new_n8971_));
  AOI21X1  g07969(.A0(new_n4546_), .A1(new_n4540_), .B0(new_n4515_), .Y(new_n8972_));
  NOR2X1   g07970(.A(new_n8969_), .B(new_n8968_), .Y(new_n8973_));
  AOI21X1  g07971(.A0(new_n4552_), .A1(new_n4545_), .B0(new_n4544_), .Y(new_n8974_));
  OAI21X1  g07972(.A0(new_n4509_), .A1(new_n4593_), .B0(new_n4596_), .Y(new_n8975_));
  OAI22X1  g07973(.A0(new_n8975_), .A1(new_n8974_), .B0(new_n4608_), .B1(new_n4607_), .Y(new_n8976_));
  NOR3X1   g07974(.A(new_n8976_), .B(new_n8973_), .C(new_n8972_), .Y(new_n8977_));
  NOR2X1   g07975(.A(new_n8977_), .B(new_n8971_), .Y(new_n8978_));
  XOR2X1   g07976(.A(new_n8978_), .B(new_n8965_), .Y(new_n8979_));
  XOR2X1   g07977(.A(new_n8979_), .B(new_n8947_), .Y(new_n8980_));
  OR2X1    g07978(.A(new_n4820_), .B(new_n4849_), .Y(new_n8981_));
  OAI21X1  g07979(.A0(new_n4867_), .A1(new_n4798_), .B0(new_n4848_), .Y(new_n8982_));
  AND2X1   g07980(.A(new_n8982_), .B(new_n8981_), .Y(new_n8983_));
  OR2X1    g07981(.A(new_n4846_), .B(new_n4845_), .Y(new_n8984_));
  XOR2X1   g07982(.A(new_n4675_), .B(new_n4683_), .Y(new_n8985_));
  XOR2X1   g07983(.A(new_n4668_), .B(new_n4662_), .Y(new_n8986_));
  OR2X1    g07984(.A(new_n4674_), .B(new_n4684_), .Y(new_n8987_));
  OAI21X1  g07985(.A0(new_n4675_), .A1(new_n4669_), .B0(new_n8987_), .Y(new_n8988_));
  AOI21X1  g07986(.A0(new_n8988_), .A1(new_n8986_), .B0(new_n8985_), .Y(new_n8989_));
  OAI21X1  g07987(.A0(new_n4723_), .A1(new_n4843_), .B0(new_n8989_), .Y(new_n8990_));
  OAI21X1  g07988(.A0(new_n4712_), .A1(new_n4721_), .B0(new_n4719_), .Y(new_n8991_));
  AOI21X1  g07989(.A0(new_n8986_), .A1(new_n4676_), .B0(new_n4687_), .Y(new_n8992_));
  XOR2X1   g07990(.A(new_n8992_), .B(new_n8991_), .Y(new_n8993_));
  AOI21X1  g07991(.A0(new_n8990_), .A1(new_n8984_), .B0(new_n8993_), .Y(new_n8994_));
  AND2X1   g07992(.A(new_n4731_), .B(new_n4730_), .Y(new_n8995_));
  AOI21X1  g07993(.A0(new_n4729_), .A1(new_n4713_), .B0(new_n4688_), .Y(new_n8996_));
  AND2X1   g07994(.A(new_n8992_), .B(new_n8991_), .Y(new_n8997_));
  NOR2X1   g07995(.A(new_n8992_), .B(new_n8991_), .Y(new_n8998_));
  NOR4X1   g07996(.A(new_n8998_), .B(new_n8997_), .C(new_n8996_), .D(new_n8995_), .Y(new_n8999_));
  OR2X1    g07997(.A(new_n8999_), .B(new_n8994_), .Y(new_n9000_));
  OR2X1    g07998(.A(new_n4832_), .B(new_n4831_), .Y(new_n9001_));
  OAI21X1  g07999(.A0(new_n4818_), .A1(new_n4830_), .B0(new_n4839_), .Y(new_n9002_));
  OAI21X1  g08000(.A0(new_n4789_), .A1(new_n4809_), .B0(new_n4813_), .Y(new_n9003_));
  AOI21X1  g08001(.A0(new_n4836_), .A1(new_n4753_), .B0(new_n4764_), .Y(new_n9004_));
  XOR2X1   g08002(.A(new_n9004_), .B(new_n9003_), .Y(new_n9005_));
  AOI21X1  g08003(.A0(new_n9002_), .A1(new_n9001_), .B0(new_n9005_), .Y(new_n9006_));
  AOI21X1  g08004(.A0(new_n4796_), .A1(new_n4790_), .B0(new_n4765_), .Y(new_n9007_));
  NOR2X1   g08005(.A(new_n9004_), .B(new_n9003_), .Y(new_n9008_));
  AOI21X1  g08006(.A0(new_n4814_), .A1(new_n4795_), .B0(new_n4794_), .Y(new_n9009_));
  OAI21X1  g08007(.A0(new_n4759_), .A1(new_n4835_), .B0(new_n4838_), .Y(new_n9010_));
  OAI22X1  g08008(.A0(new_n9010_), .A1(new_n9009_), .B0(new_n4832_), .B1(new_n4831_), .Y(new_n9011_));
  NOR3X1   g08009(.A(new_n9011_), .B(new_n9008_), .C(new_n9007_), .Y(new_n9012_));
  NOR2X1   g08010(.A(new_n9012_), .B(new_n9006_), .Y(new_n9013_));
  XOR2X1   g08011(.A(new_n9013_), .B(new_n9000_), .Y(new_n9014_));
  XOR2X1   g08012(.A(new_n9014_), .B(new_n8983_), .Y(new_n9015_));
  XOR2X1   g08013(.A(new_n9015_), .B(new_n8980_), .Y(new_n9016_));
  XOR2X1   g08014(.A(new_n9016_), .B(new_n8934_), .Y(new_n9017_));
  XOR2X1   g08015(.A(new_n9017_), .B(new_n8931_), .Y(new_n9018_));
  NAND2X1  g08016(.A(new_n9018_), .B(new_n8860_), .Y(new_n9019_));
  OAI21X1  g08017(.A0(new_n4008_), .A1(new_n4002_), .B0(new_n4181_), .Y(new_n9020_));
  OAI21X1  g08018(.A0(new_n4183_), .A1(new_n4179_), .B0(new_n9020_), .Y(new_n9021_));
  AOI21X1  g08019(.A0(new_n4129_), .A1(new_n4113_), .B0(new_n4137_), .Y(new_n9022_));
  AOI21X1  g08020(.A0(new_n4176_), .A1(new_n4171_), .B0(new_n9022_), .Y(new_n9023_));
  AOI21X1  g08021(.A0(new_n4158_), .A1(new_n4152_), .B0(new_n4147_), .Y(new_n9024_));
  OR2X1    g08022(.A(new_n9024_), .B(new_n4169_), .Y(new_n9025_));
  XOR2X1   g08023(.A(new_n4062_), .B(new_n4149_), .Y(new_n9026_));
  AOI21X1  g08024(.A0(new_n4157_), .A1(new_n9026_), .B0(new_n4156_), .Y(new_n9027_));
  XOR2X1   g08025(.A(new_n4080_), .B(new_n4074_), .Y(new_n9028_));
  AOI21X1  g08026(.A0(new_n4146_), .A1(new_n9028_), .B0(new_n4145_), .Y(new_n9029_));
  XOR2X1   g08027(.A(new_n9029_), .B(new_n9027_), .Y(new_n9030_));
  AND2X1   g08028(.A(new_n4154_), .B(new_n4153_), .Y(new_n9031_));
  OAI22X1  g08029(.A0(new_n4162_), .A1(new_n4148_), .B0(new_n4155_), .B1(new_n9031_), .Y(new_n9032_));
  AND2X1   g08030(.A(new_n9029_), .B(new_n9032_), .Y(new_n9033_));
  NOR2X1   g08031(.A(new_n9029_), .B(new_n9032_), .Y(new_n9034_));
  NOR4X1   g08032(.A(new_n9034_), .B(new_n9033_), .C(new_n9024_), .D(new_n4169_), .Y(new_n9035_));
  AOI21X1  g08033(.A0(new_n9030_), .A1(new_n9025_), .B0(new_n9035_), .Y(new_n9036_));
  AOI21X1  g08034(.A0(new_n4111_), .A1(new_n4105_), .B0(new_n4099_), .Y(new_n9037_));
  OR2X1    g08035(.A(new_n9037_), .B(new_n4128_), .Y(new_n9038_));
  XOR2X1   g08036(.A(new_n4024_), .B(new_n4018_), .Y(new_n9039_));
  AOI21X1  g08037(.A0(new_n4110_), .A1(new_n9039_), .B0(new_n4109_), .Y(new_n9040_));
  AOI21X1  g08038(.A0(new_n4098_), .A1(new_n4114_), .B0(new_n4097_), .Y(new_n9041_));
  XOR2X1   g08039(.A(new_n9041_), .B(new_n9040_), .Y(new_n9042_));
  AND2X1   g08040(.A(new_n4107_), .B(new_n4106_), .Y(new_n9043_));
  OAI22X1  g08041(.A0(new_n4125_), .A1(new_n4102_), .B0(new_n4108_), .B1(new_n9043_), .Y(new_n9044_));
  AND2X1   g08042(.A(new_n9041_), .B(new_n9044_), .Y(new_n9045_));
  NOR2X1   g08043(.A(new_n9041_), .B(new_n9044_), .Y(new_n9046_));
  NOR4X1   g08044(.A(new_n9046_), .B(new_n9045_), .C(new_n9037_), .D(new_n4128_), .Y(new_n9047_));
  AOI21X1  g08045(.A0(new_n9042_), .A1(new_n9038_), .B0(new_n9047_), .Y(new_n9048_));
  XOR2X1   g08046(.A(new_n9048_), .B(new_n9036_), .Y(new_n9049_));
  XOR2X1   g08047(.A(new_n9049_), .B(new_n9023_), .Y(new_n9050_));
  AOI21X1  g08048(.A0(new_n3989_), .A1(new_n3981_), .B0(new_n4000_), .Y(new_n9051_));
  AOI21X1  g08049(.A0(new_n4006_), .A1(new_n3919_), .B0(new_n9051_), .Y(new_n9052_));
  OAI21X1  g08050(.A0(new_n3913_), .A1(new_n3909_), .B0(new_n4003_), .Y(new_n9053_));
  AND2X1   g08051(.A(new_n3900_), .B(new_n3899_), .Y(new_n9054_));
  OAI22X1  g08052(.A0(new_n3906_), .A1(new_n3911_), .B0(new_n3901_), .B1(new_n9054_), .Y(new_n9055_));
  XOR2X1   g08053(.A(new_n3869_), .B(new_n3872_), .Y(new_n9056_));
  OR2X1    g08054(.A(new_n3869_), .B(new_n3872_), .Y(new_n9057_));
  AOI22X1  g08055(.A0(new_n3874_), .A1(new_n9057_), .B0(new_n3871_), .B1(new_n9056_), .Y(new_n9058_));
  XOR2X1   g08056(.A(new_n9058_), .B(new_n9055_), .Y(new_n9059_));
  AOI21X1  g08057(.A0(new_n9053_), .A1(new_n3917_), .B0(new_n9059_), .Y(new_n9060_));
  NOR4X1   g08058(.A(new_n3916_), .B(new_n3915_), .C(new_n3914_), .D(new_n3911_), .Y(new_n9061_));
  AND2X1   g08059(.A(new_n9058_), .B(new_n9055_), .Y(new_n9062_));
  NOR2X1   g08060(.A(new_n9058_), .B(new_n9055_), .Y(new_n9063_));
  NOR3X1   g08061(.A(new_n9063_), .B(new_n9062_), .C(new_n9061_), .Y(new_n9064_));
  AND2X1   g08062(.A(new_n9064_), .B(new_n9053_), .Y(new_n9065_));
  NOR2X1   g08063(.A(new_n9065_), .B(new_n9060_), .Y(new_n9066_));
  AND2X1   g08064(.A(new_n3979_), .B(new_n3973_), .Y(new_n9067_));
  OR4X1    g08065(.A(new_n3972_), .B(new_n3969_), .C(new_n3983_), .D(new_n3950_), .Y(new_n9068_));
  AOI21X1  g08066(.A0(new_n3972_), .A1(new_n3983_), .B0(new_n3977_), .Y(new_n9069_));
  OAI22X1  g08067(.A0(new_n9069_), .A1(new_n9068_), .B0(new_n9067_), .B1(new_n3947_), .Y(new_n9070_));
  AOI21X1  g08068(.A0(new_n3986_), .A1(new_n3978_), .B0(new_n3977_), .Y(new_n9071_));
  OR2X1    g08069(.A(new_n3950_), .B(new_n3940_), .Y(new_n9072_));
  AND2X1   g08070(.A(new_n9072_), .B(new_n3945_), .Y(new_n9073_));
  XOR2X1   g08071(.A(new_n9073_), .B(new_n9071_), .Y(new_n9074_));
  AND2X1   g08072(.A(new_n9074_), .B(new_n9070_), .Y(new_n9075_));
  NOR2X1   g08073(.A(new_n9067_), .B(new_n3947_), .Y(new_n9076_));
  OAI21X1  g08074(.A0(new_n3950_), .A1(new_n3940_), .B0(new_n3945_), .Y(new_n9077_));
  AND2X1   g08075(.A(new_n9077_), .B(new_n9071_), .Y(new_n9078_));
  OAI22X1  g08076(.A0(new_n9077_), .A1(new_n9071_), .B0(new_n9069_), .B1(new_n9068_), .Y(new_n9079_));
  NOR3X1   g08077(.A(new_n9079_), .B(new_n9078_), .C(new_n9076_), .Y(new_n9080_));
  NOR2X1   g08078(.A(new_n9080_), .B(new_n9075_), .Y(new_n9081_));
  XOR2X1   g08079(.A(new_n9081_), .B(new_n9066_), .Y(new_n9082_));
  XOR2X1   g08080(.A(new_n9082_), .B(new_n9052_), .Y(new_n9083_));
  XOR2X1   g08081(.A(new_n9083_), .B(new_n9050_), .Y(new_n9084_));
  XOR2X1   g08082(.A(new_n9084_), .B(new_n9021_), .Y(new_n9085_));
  OR2X1    g08083(.A(new_n4876_), .B(new_n4889_), .Y(new_n9086_));
  OAI21X1  g08084(.A0(new_n4890_), .A1(new_n4854_), .B0(new_n4888_), .Y(new_n9087_));
  AND2X1   g08085(.A(new_n9087_), .B(new_n9086_), .Y(new_n9088_));
  AND2X1   g08086(.A(new_n4436_), .B(new_n4480_), .Y(new_n9089_));
  AOI21X1  g08087(.A0(new_n4473_), .A1(new_n4469_), .B0(new_n4476_), .Y(new_n9090_));
  AOI22X1  g08088(.A0(new_n8887_), .A1(new_n4476_), .B0(new_n9090_), .B1(new_n8889_), .Y(new_n9091_));
  AOI22X1  g08089(.A0(new_n8890_), .A1(new_n8889_), .B0(new_n8887_), .B1(new_n4464_), .Y(new_n9092_));
  MX2X1    g08090(.A(new_n9092_), .B(new_n9091_), .S0(new_n4445_), .Y(new_n9093_));
  AOI21X1  g08091(.A0(new_n4481_), .A1(new_n4363_), .B0(new_n9093_), .Y(new_n9094_));
  OR2X1    g08092(.A(new_n9094_), .B(new_n9089_), .Y(new_n9095_));
  XOR2X1   g08093(.A(new_n8930_), .B(new_n9095_), .Y(new_n9096_));
  XOR2X1   g08094(.A(new_n9017_), .B(new_n9096_), .Y(new_n9097_));
  AOI21X1  g08095(.A0(new_n9097_), .A1(new_n9088_), .B0(new_n9085_), .Y(new_n9098_));
  XOR2X1   g08096(.A(new_n9097_), .B(new_n8860_), .Y(new_n9099_));
  AOI22X1  g08097(.A0(new_n9099_), .A1(new_n9085_), .B0(new_n9098_), .B1(new_n9019_), .Y(new_n9100_));
  OR2X1    g08098(.A(new_n9100_), .B(new_n8857_), .Y(new_n9101_));
  NOR3X1   g08099(.A(new_n5625_), .B(new_n5621_), .C(new_n5617_), .Y(new_n9102_));
  OAI21X1  g08100(.A0(new_n9102_), .A1(new_n5636_), .B0(new_n5627_), .Y(new_n9103_));
  AOI21X1  g08101(.A0(new_n5633_), .A1(new_n5431_), .B0(new_n5433_), .Y(new_n9104_));
  AOI21X1  g08102(.A0(new_n5385_), .A1(new_n5369_), .B0(new_n5392_), .Y(new_n9105_));
  AOI21X1  g08103(.A0(new_n5428_), .A1(new_n5423_), .B0(new_n9105_), .Y(new_n9106_));
  AOI21X1  g08104(.A0(new_n5413_), .A1(new_n5407_), .B0(new_n5402_), .Y(new_n9107_));
  OR2X1    g08105(.A(new_n9107_), .B(new_n5421_), .Y(new_n9108_));
  XOR2X1   g08106(.A(new_n5209_), .B(new_n5404_), .Y(new_n9109_));
  AOI21X1  g08107(.A0(new_n5412_), .A1(new_n9109_), .B0(new_n5411_), .Y(new_n9110_));
  XOR2X1   g08108(.A(new_n5227_), .B(new_n5221_), .Y(new_n9111_));
  AOI21X1  g08109(.A0(new_n5401_), .A1(new_n9111_), .B0(new_n5400_), .Y(new_n9112_));
  XOR2X1   g08110(.A(new_n9112_), .B(new_n9110_), .Y(new_n9113_));
  AND2X1   g08111(.A(new_n5409_), .B(new_n5408_), .Y(new_n9114_));
  OAI22X1  g08112(.A0(new_n5417_), .A1(new_n5403_), .B0(new_n5410_), .B1(new_n9114_), .Y(new_n9115_));
  AND2X1   g08113(.A(new_n9112_), .B(new_n9115_), .Y(new_n9116_));
  NOR2X1   g08114(.A(new_n9112_), .B(new_n9115_), .Y(new_n9117_));
  NOR4X1   g08115(.A(new_n9117_), .B(new_n9116_), .C(new_n9107_), .D(new_n5421_), .Y(new_n9118_));
  AOI21X1  g08116(.A0(new_n9113_), .A1(new_n9108_), .B0(new_n9118_), .Y(new_n9119_));
  AOI21X1  g08117(.A0(new_n5367_), .A1(new_n5361_), .B0(new_n5355_), .Y(new_n9120_));
  OR2X1    g08118(.A(new_n9120_), .B(new_n5384_), .Y(new_n9121_));
  XOR2X1   g08119(.A(new_n5170_), .B(new_n5164_), .Y(new_n9122_));
  AOI21X1  g08120(.A0(new_n5366_), .A1(new_n9122_), .B0(new_n5365_), .Y(new_n9123_));
  AOI21X1  g08121(.A0(new_n5354_), .A1(new_n5370_), .B0(new_n5353_), .Y(new_n9124_));
  XOR2X1   g08122(.A(new_n9124_), .B(new_n9123_), .Y(new_n9125_));
  AND2X1   g08123(.A(new_n5363_), .B(new_n5362_), .Y(new_n9126_));
  OAI22X1  g08124(.A0(new_n5381_), .A1(new_n5358_), .B0(new_n5364_), .B1(new_n9126_), .Y(new_n9127_));
  AND2X1   g08125(.A(new_n9124_), .B(new_n9127_), .Y(new_n9128_));
  NOR2X1   g08126(.A(new_n9124_), .B(new_n9127_), .Y(new_n9129_));
  NOR4X1   g08127(.A(new_n9129_), .B(new_n9128_), .C(new_n9120_), .D(new_n5384_), .Y(new_n9130_));
  AOI21X1  g08128(.A0(new_n9125_), .A1(new_n9121_), .B0(new_n9130_), .Y(new_n9131_));
  XOR2X1   g08129(.A(new_n9131_), .B(new_n9119_), .Y(new_n9132_));
  XOR2X1   g08130(.A(new_n9132_), .B(new_n9106_), .Y(new_n9133_));
  AOI21X1  g08131(.A0(new_n5341_), .A1(new_n5331_), .B0(new_n5333_), .Y(new_n9134_));
  AOI21X1  g08132(.A0(new_n5270_), .A1(new_n5264_), .B0(new_n5258_), .Y(new_n9135_));
  OR2X1    g08133(.A(new_n9135_), .B(new_n5279_), .Y(new_n9136_));
  XOR2X1   g08134(.A(new_n5132_), .B(new_n5261_), .Y(new_n9137_));
  AOI21X1  g08135(.A0(new_n5269_), .A1(new_n9137_), .B0(new_n5268_), .Y(new_n9138_));
  XOR2X1   g08136(.A(new_n5150_), .B(new_n5144_), .Y(new_n9139_));
  AOI21X1  g08137(.A0(new_n5257_), .A1(new_n9139_), .B0(new_n5256_), .Y(new_n9140_));
  XOR2X1   g08138(.A(new_n9140_), .B(new_n9138_), .Y(new_n9141_));
  AND2X1   g08139(.A(new_n5266_), .B(new_n5265_), .Y(new_n9142_));
  OAI22X1  g08140(.A0(new_n5275_), .A1(new_n5260_), .B0(new_n5267_), .B1(new_n9142_), .Y(new_n9143_));
  AND2X1   g08141(.A(new_n9140_), .B(new_n9143_), .Y(new_n9144_));
  NOR2X1   g08142(.A(new_n9140_), .B(new_n9143_), .Y(new_n9145_));
  NOR4X1   g08143(.A(new_n9145_), .B(new_n9144_), .C(new_n9135_), .D(new_n5279_), .Y(new_n9146_));
  AOI21X1  g08144(.A0(new_n9141_), .A1(new_n9136_), .B0(new_n9146_), .Y(new_n9147_));
  AOI21X1  g08145(.A0(new_n5302_), .A1(new_n5296_), .B0(new_n5290_), .Y(new_n9148_));
  OR2X1    g08146(.A(new_n9148_), .B(new_n5326_), .Y(new_n9149_));
  XOR2X1   g08147(.A(new_n5094_), .B(new_n5088_), .Y(new_n9150_));
  AOI21X1  g08148(.A0(new_n5301_), .A1(new_n9150_), .B0(new_n5300_), .Y(new_n9151_));
  AOI21X1  g08149(.A0(new_n5289_), .A1(new_n5320_), .B0(new_n5288_), .Y(new_n9152_));
  XOR2X1   g08150(.A(new_n9152_), .B(new_n9151_), .Y(new_n9153_));
  AND2X1   g08151(.A(new_n5298_), .B(new_n5297_), .Y(new_n9154_));
  OAI22X1  g08152(.A0(new_n5307_), .A1(new_n5293_), .B0(new_n5299_), .B1(new_n9154_), .Y(new_n9155_));
  AND2X1   g08153(.A(new_n9152_), .B(new_n9155_), .Y(new_n9156_));
  NOR2X1   g08154(.A(new_n9152_), .B(new_n9155_), .Y(new_n9157_));
  NOR4X1   g08155(.A(new_n9157_), .B(new_n9156_), .C(new_n9148_), .D(new_n5326_), .Y(new_n9158_));
  AOI21X1  g08156(.A0(new_n9153_), .A1(new_n9149_), .B0(new_n9158_), .Y(new_n9159_));
  XOR2X1   g08157(.A(new_n9159_), .B(new_n9147_), .Y(new_n9160_));
  XOR2X1   g08158(.A(new_n9160_), .B(new_n9134_), .Y(new_n9161_));
  XOR2X1   g08159(.A(new_n9161_), .B(new_n9133_), .Y(new_n9162_));
  XOR2X1   g08160(.A(new_n9162_), .B(new_n9104_), .Y(new_n9163_));
  AOI21X1  g08161(.A0(new_n5605_), .A1(new_n5601_), .B0(new_n5615_), .Y(new_n9164_));
  AOI21X1  g08162(.A0(new_n5619_), .A1(new_n5520_), .B0(new_n9164_), .Y(new_n9165_));
  AOI21X1  g08163(.A0(new_n5474_), .A1(new_n5458_), .B0(new_n5481_), .Y(new_n9166_));
  AOI21X1  g08164(.A0(new_n5517_), .A1(new_n5512_), .B0(new_n9166_), .Y(new_n9167_));
  AOI21X1  g08165(.A0(new_n5502_), .A1(new_n5496_), .B0(new_n5491_), .Y(new_n9168_));
  OR2X1    g08166(.A(new_n9168_), .B(new_n5510_), .Y(new_n9169_));
  XOR2X1   g08167(.A(new_n5055_), .B(new_n5493_), .Y(new_n9170_));
  AOI21X1  g08168(.A0(new_n5501_), .A1(new_n9170_), .B0(new_n5500_), .Y(new_n9171_));
  XOR2X1   g08169(.A(new_n5073_), .B(new_n5067_), .Y(new_n9172_));
  AOI21X1  g08170(.A0(new_n5490_), .A1(new_n9172_), .B0(new_n5489_), .Y(new_n9173_));
  XOR2X1   g08171(.A(new_n9173_), .B(new_n9171_), .Y(new_n9174_));
  AND2X1   g08172(.A(new_n5498_), .B(new_n5497_), .Y(new_n9175_));
  OAI22X1  g08173(.A0(new_n5506_), .A1(new_n5492_), .B0(new_n5499_), .B1(new_n9175_), .Y(new_n9176_));
  AND2X1   g08174(.A(new_n9173_), .B(new_n9176_), .Y(new_n9177_));
  NOR2X1   g08175(.A(new_n9173_), .B(new_n9176_), .Y(new_n9178_));
  NOR4X1   g08176(.A(new_n9178_), .B(new_n9177_), .C(new_n9168_), .D(new_n5510_), .Y(new_n9179_));
  AOI21X1  g08177(.A0(new_n9174_), .A1(new_n9169_), .B0(new_n9179_), .Y(new_n9180_));
  AOI21X1  g08178(.A0(new_n5456_), .A1(new_n5450_), .B0(new_n5444_), .Y(new_n9181_));
  OR2X1    g08179(.A(new_n9181_), .B(new_n5473_), .Y(new_n9182_));
  XOR2X1   g08180(.A(new_n5016_), .B(new_n5010_), .Y(new_n9183_));
  AOI21X1  g08181(.A0(new_n5455_), .A1(new_n9183_), .B0(new_n5454_), .Y(new_n9184_));
  AOI21X1  g08182(.A0(new_n5443_), .A1(new_n5459_), .B0(new_n5442_), .Y(new_n9185_));
  XOR2X1   g08183(.A(new_n9185_), .B(new_n9184_), .Y(new_n9186_));
  AND2X1   g08184(.A(new_n5452_), .B(new_n5451_), .Y(new_n9187_));
  OAI22X1  g08185(.A0(new_n5470_), .A1(new_n5447_), .B0(new_n5453_), .B1(new_n9187_), .Y(new_n9188_));
  AND2X1   g08186(.A(new_n9185_), .B(new_n9188_), .Y(new_n9189_));
  NOR2X1   g08187(.A(new_n9185_), .B(new_n9188_), .Y(new_n9190_));
  NOR4X1   g08188(.A(new_n9190_), .B(new_n9189_), .C(new_n9181_), .D(new_n5473_), .Y(new_n9191_));
  AOI21X1  g08189(.A0(new_n9186_), .A1(new_n9182_), .B0(new_n9191_), .Y(new_n9192_));
  XOR2X1   g08190(.A(new_n9192_), .B(new_n9180_), .Y(new_n9193_));
  XOR2X1   g08191(.A(new_n9193_), .B(new_n9167_), .Y(new_n9194_));
  AOI21X1  g08192(.A0(new_n5612_), .A1(new_n5602_), .B0(new_n5604_), .Y(new_n9195_));
  AOI21X1  g08193(.A0(new_n5541_), .A1(new_n5535_), .B0(new_n5529_), .Y(new_n9196_));
  OR2X1    g08194(.A(new_n9196_), .B(new_n5550_), .Y(new_n9197_));
  XOR2X1   g08195(.A(new_n4978_), .B(new_n5532_), .Y(new_n9198_));
  AOI21X1  g08196(.A0(new_n5540_), .A1(new_n9198_), .B0(new_n5539_), .Y(new_n9199_));
  XOR2X1   g08197(.A(new_n4996_), .B(new_n4990_), .Y(new_n9200_));
  AOI21X1  g08198(.A0(new_n5528_), .A1(new_n9200_), .B0(new_n5527_), .Y(new_n9201_));
  XOR2X1   g08199(.A(new_n9201_), .B(new_n9199_), .Y(new_n9202_));
  AND2X1   g08200(.A(new_n5537_), .B(new_n5536_), .Y(new_n9203_));
  OAI22X1  g08201(.A0(new_n5546_), .A1(new_n5531_), .B0(new_n5538_), .B1(new_n9203_), .Y(new_n9204_));
  AND2X1   g08202(.A(new_n9201_), .B(new_n9204_), .Y(new_n9205_));
  NOR2X1   g08203(.A(new_n9201_), .B(new_n9204_), .Y(new_n9206_));
  NOR4X1   g08204(.A(new_n9206_), .B(new_n9205_), .C(new_n9196_), .D(new_n5550_), .Y(new_n9207_));
  AOI21X1  g08205(.A0(new_n9202_), .A1(new_n9197_), .B0(new_n9207_), .Y(new_n9208_));
  AOI21X1  g08206(.A0(new_n5573_), .A1(new_n5567_), .B0(new_n5561_), .Y(new_n9209_));
  OR2X1    g08207(.A(new_n9209_), .B(new_n5597_), .Y(new_n9210_));
  XOR2X1   g08208(.A(new_n4940_), .B(new_n4934_), .Y(new_n9211_));
  AOI21X1  g08209(.A0(new_n5572_), .A1(new_n9211_), .B0(new_n5571_), .Y(new_n9212_));
  AOI21X1  g08210(.A0(new_n5560_), .A1(new_n5591_), .B0(new_n5559_), .Y(new_n9213_));
  XOR2X1   g08211(.A(new_n9213_), .B(new_n9212_), .Y(new_n9214_));
  AND2X1   g08212(.A(new_n5569_), .B(new_n5568_), .Y(new_n9215_));
  OAI22X1  g08213(.A0(new_n5578_), .A1(new_n5564_), .B0(new_n5570_), .B1(new_n9215_), .Y(new_n9216_));
  AND2X1   g08214(.A(new_n9213_), .B(new_n9216_), .Y(new_n9217_));
  NOR2X1   g08215(.A(new_n9213_), .B(new_n9216_), .Y(new_n9218_));
  NOR4X1   g08216(.A(new_n9218_), .B(new_n9217_), .C(new_n9209_), .D(new_n5597_), .Y(new_n9219_));
  AOI21X1  g08217(.A0(new_n9214_), .A1(new_n9210_), .B0(new_n9219_), .Y(new_n9220_));
  XOR2X1   g08218(.A(new_n9220_), .B(new_n9208_), .Y(new_n9221_));
  XOR2X1   g08219(.A(new_n9221_), .B(new_n9195_), .Y(new_n9222_));
  XOR2X1   g08220(.A(new_n9222_), .B(new_n9194_), .Y(new_n9223_));
  XOR2X1   g08221(.A(new_n9223_), .B(new_n9165_), .Y(new_n9224_));
  XOR2X1   g08222(.A(new_n9224_), .B(new_n9163_), .Y(new_n9225_));
  XOR2X1   g08223(.A(new_n9225_), .B(new_n9103_), .Y(new_n9226_));
  AOI21X1  g08224(.A0(new_n9100_), .A1(new_n8857_), .B0(new_n9226_), .Y(new_n9227_));
  AND2X1   g08225(.A(new_n5241_), .B(new_n4897_), .Y(new_n9228_));
  AOI21X1  g08226(.A0(new_n5245_), .A1(new_n5244_), .B0(new_n5239_), .Y(new_n9229_));
  OR2X1    g08227(.A(new_n9229_), .B(new_n9228_), .Y(new_n9230_));
  XOR2X1   g08228(.A(new_n9100_), .B(new_n9230_), .Y(new_n9231_));
  AOI22X1  g08229(.A0(new_n9231_), .A1(new_n9226_), .B0(new_n9227_), .B1(new_n9101_), .Y(new_n9232_));
  XOR2X1   g08230(.A(new_n9232_), .B(new_n8854_), .Y(new_n9233_));
  AOI21X1  g08231(.A0(new_n8820_), .A1(new_n8804_), .B0(new_n7209_), .Y(new_n9234_));
  OR2X1    g08232(.A(new_n9234_), .B(new_n8822_), .Y(new_n9235_));
  OR2X1    g08233(.A(new_n8815_), .B(new_n6714_), .Y(new_n9236_));
  AND2X1   g08234(.A(new_n6979_), .B(new_n6976_), .Y(new_n9237_));
  AOI21X1  g08235(.A0(new_n6931_), .A1(new_n6866_), .B0(new_n6977_), .Y(new_n9238_));
  AOI22X1  g08236(.A0(new_n9238_), .A1(new_n6921_), .B0(new_n6944_), .B1(new_n6977_), .Y(new_n9239_));
  OAI21X1  g08237(.A0(new_n9239_), .A1(new_n6976_), .B0(new_n6948_), .Y(new_n9240_));
  MX2X1    g08238(.A(new_n9239_), .B(new_n6945_), .S0(new_n6976_), .Y(new_n9241_));
  OAI22X1  g08239(.A0(new_n9241_), .A1(new_n6948_), .B0(new_n9240_), .B1(new_n9237_), .Y(new_n9242_));
  OAI21X1  g08240(.A0(new_n9239_), .A1(new_n6976_), .B0(new_n6949_), .Y(new_n9243_));
  OAI22X1  g08241(.A0(new_n9243_), .A1(new_n9237_), .B0(new_n9241_), .B1(new_n6949_), .Y(new_n9244_));
  MX2X1    g08242(.A(new_n9244_), .B(new_n9242_), .S0(new_n7203_), .Y(new_n9245_));
  OAI21X1  g08243(.A0(new_n8817_), .A1(new_n8811_), .B0(new_n9245_), .Y(new_n9246_));
  AND2X1   g08244(.A(new_n9246_), .B(new_n9236_), .Y(new_n9247_));
  OR2X1    g08245(.A(new_n9241_), .B(new_n6949_), .Y(new_n9248_));
  AND2X1   g08246(.A(new_n7099_), .B(new_n7096_), .Y(new_n9249_));
  AOI21X1  g08247(.A0(new_n7074_), .A1(new_n7061_), .B0(new_n7097_), .Y(new_n9250_));
  AOI22X1  g08248(.A0(new_n9250_), .A1(new_n7051_), .B0(new_n7076_), .B1(new_n7097_), .Y(new_n9251_));
  OAI21X1  g08249(.A0(new_n9251_), .A1(new_n7096_), .B0(new_n7200_), .Y(new_n9252_));
  MX2X1    g08250(.A(new_n9251_), .B(new_n7077_), .S0(new_n7096_), .Y(new_n9253_));
  OAI22X1  g08251(.A0(new_n9253_), .A1(new_n7200_), .B0(new_n9252_), .B1(new_n9249_), .Y(new_n9254_));
  OAI21X1  g08252(.A0(new_n9251_), .A1(new_n7096_), .B0(new_n7079_), .Y(new_n9255_));
  OAI22X1  g08253(.A0(new_n9255_), .A1(new_n9249_), .B0(new_n9253_), .B1(new_n7079_), .Y(new_n9256_));
  MX2X1    g08254(.A(new_n9256_), .B(new_n9254_), .S0(new_n7199_), .Y(new_n9257_));
  OAI21X1  g08255(.A0(new_n9243_), .A1(new_n9237_), .B0(new_n9257_), .Y(new_n9258_));
  AND2X1   g08256(.A(new_n9258_), .B(new_n9248_), .Y(new_n9259_));
  AND2X1   g08257(.A(new_n7100_), .B(new_n7200_), .Y(new_n9260_));
  AOI21X1  g08258(.A0(new_n7201_), .A1(new_n7078_), .B0(new_n7199_), .Y(new_n9261_));
  OR2X1    g08259(.A(new_n9261_), .B(new_n9260_), .Y(new_n9262_));
  XOR2X1   g08260(.A(new_n7149_), .B(new_n7121_), .Y(new_n9263_));
  NOR4X1   g08261(.A(new_n7107_), .B(new_n7148_), .C(new_n7147_), .D(new_n7114_), .Y(new_n9264_));
  AOI21X1  g08262(.A0(new_n7147_), .A1(new_n7141_), .B0(new_n7120_), .Y(new_n9265_));
  AOI22X1  g08263(.A0(new_n9265_), .A1(new_n9264_), .B0(new_n7127_), .B1(new_n7121_), .Y(new_n9266_));
  MX2X1    g08264(.A(new_n9266_), .B(new_n9263_), .S0(new_n7113_), .Y(new_n9267_));
  OR2X1    g08265(.A(new_n9267_), .B(new_n7130_), .Y(new_n9268_));
  AND2X1   g08266(.A(new_n7128_), .B(new_n7113_), .Y(new_n9269_));
  NOR4X1   g08267(.A(new_n7174_), .B(new_n7161_), .C(new_n7173_), .D(new_n7168_), .Y(new_n9270_));
  XOR2X1   g08268(.A(new_n7185_), .B(new_n9270_), .Y(new_n9271_));
  OR4X1    g08269(.A(new_n7161_), .B(new_n7173_), .C(new_n7184_), .D(new_n7168_), .Y(new_n9272_));
  AND2X1   g08270(.A(new_n6702_), .B(\A[84] ), .Y(new_n9273_));
  OR2X1    g08271(.A(new_n9273_), .B(new_n6704_), .Y(new_n9274_));
  XOR2X1   g08272(.A(new_n6707_), .B(new_n9274_), .Y(new_n9275_));
  XOR2X1   g08273(.A(new_n7163_), .B(new_n9275_), .Y(new_n9276_));
  OAI22X1  g08274(.A0(new_n9276_), .A1(new_n7165_), .B0(new_n7189_), .B1(new_n7168_), .Y(new_n9277_));
  OAI22X1  g08275(.A0(new_n9277_), .A1(new_n9272_), .B0(new_n7185_), .B1(new_n9270_), .Y(new_n9278_));
  MX2X1    g08276(.A(new_n9278_), .B(new_n9271_), .S0(new_n7167_), .Y(new_n9279_));
  OAI21X1  g08277(.A0(new_n9266_), .A1(new_n7113_), .B0(new_n7130_), .Y(new_n9280_));
  OAI21X1  g08278(.A0(new_n9280_), .A1(new_n9269_), .B0(new_n9279_), .Y(new_n9281_));
  AND2X1   g08279(.A(new_n9281_), .B(new_n9268_), .Y(new_n9282_));
  OR2X1    g08280(.A(new_n9277_), .B(new_n9272_), .Y(new_n9283_));
  XOR2X1   g08281(.A(new_n6703_), .B(new_n6697_), .Y(new_n9284_));
  OR2X1    g08282(.A(new_n6703_), .B(new_n6697_), .Y(new_n9285_));
  OR2X1    g08283(.A(new_n6707_), .B(new_n6705_), .Y(new_n9286_));
  OAI21X1  g08284(.A0(new_n9285_), .A1(new_n9275_), .B0(new_n9286_), .Y(new_n9287_));
  AOI21X1  g08285(.A0(new_n9287_), .A1(new_n9284_), .B0(new_n9276_), .Y(new_n9288_));
  OAI21X1  g08286(.A0(new_n7185_), .A1(new_n9270_), .B0(new_n9288_), .Y(new_n9289_));
  OAI21X1  g08287(.A0(new_n7184_), .A1(new_n7168_), .B0(new_n7182_), .Y(new_n9290_));
  AOI21X1  g08288(.A0(new_n7166_), .A1(new_n9284_), .B0(new_n7165_), .Y(new_n9291_));
  XOR2X1   g08289(.A(new_n9291_), .B(new_n9290_), .Y(new_n9292_));
  AOI21X1  g08290(.A0(new_n9289_), .A1(new_n9283_), .B0(new_n9292_), .Y(new_n9293_));
  AND2X1   g08291(.A(new_n7193_), .B(new_n7192_), .Y(new_n9294_));
  AOI21X1  g08292(.A0(new_n7191_), .A1(new_n7175_), .B0(new_n7167_), .Y(new_n9295_));
  AND2X1   g08293(.A(new_n9291_), .B(new_n9290_), .Y(new_n9296_));
  NOR2X1   g08294(.A(new_n9291_), .B(new_n9290_), .Y(new_n9297_));
  NOR4X1   g08295(.A(new_n9297_), .B(new_n9296_), .C(new_n9295_), .D(new_n9294_), .Y(new_n9298_));
  NOR2X1   g08296(.A(new_n9298_), .B(new_n9293_), .Y(new_n9299_));
  OR2X1    g08297(.A(new_n7151_), .B(new_n7150_), .Y(new_n9300_));
  OAI21X1  g08298(.A0(new_n7149_), .A1(new_n7140_), .B0(new_n7139_), .Y(new_n9301_));
  OAI21X1  g08299(.A0(new_n7148_), .A1(new_n7114_), .B0(new_n7147_), .Y(new_n9302_));
  AOI21X1  g08300(.A0(new_n7112_), .A1(new_n7131_), .B0(new_n7111_), .Y(new_n9303_));
  XOR2X1   g08301(.A(new_n9303_), .B(new_n9302_), .Y(new_n9304_));
  AOI21X1  g08302(.A0(new_n9301_), .A1(new_n9300_), .B0(new_n9304_), .Y(new_n9305_));
  AOI21X1  g08303(.A0(new_n7127_), .A1(new_n7121_), .B0(new_n7113_), .Y(new_n9306_));
  NOR2X1   g08304(.A(new_n9303_), .B(new_n9302_), .Y(new_n9307_));
  AOI21X1  g08305(.A0(new_n7126_), .A1(new_n7141_), .B0(new_n7125_), .Y(new_n9308_));
  OAI21X1  g08306(.A0(new_n7138_), .A1(new_n7107_), .B0(new_n7137_), .Y(new_n9309_));
  OAI22X1  g08307(.A0(new_n9309_), .A1(new_n9308_), .B0(new_n7151_), .B1(new_n7150_), .Y(new_n9310_));
  NOR3X1   g08308(.A(new_n9310_), .B(new_n9307_), .C(new_n9306_), .Y(new_n9311_));
  NOR2X1   g08309(.A(new_n9311_), .B(new_n9305_), .Y(new_n9312_));
  XOR2X1   g08310(.A(new_n9312_), .B(new_n9299_), .Y(new_n9313_));
  XOR2X1   g08311(.A(new_n9313_), .B(new_n9282_), .Y(new_n9314_));
  OR2X1    g08312(.A(new_n7085_), .B(new_n7052_), .Y(new_n9315_));
  OAI21X1  g08313(.A0(new_n7086_), .A1(new_n7080_), .B0(new_n7023_), .Y(new_n9316_));
  AND2X1   g08314(.A(new_n9316_), .B(new_n9315_), .Y(new_n9317_));
  OR2X1    g08315(.A(new_n7021_), .B(new_n7013_), .Y(new_n9318_));
  XOR2X1   g08316(.A(new_n6628_), .B(new_n6622_), .Y(new_n9319_));
  OR2X1    g08317(.A(new_n6628_), .B(new_n6622_), .Y(new_n9320_));
  OR2X1    g08318(.A(new_n6632_), .B(new_n6630_), .Y(new_n9321_));
  OAI21X1  g08319(.A0(new_n9320_), .A1(new_n7019_), .B0(new_n9321_), .Y(new_n9322_));
  AOI21X1  g08320(.A0(new_n9322_), .A1(new_n9319_), .B0(new_n7020_), .Y(new_n9323_));
  OAI21X1  g08321(.A0(new_n7011_), .A1(new_n7001_), .B0(new_n9323_), .Y(new_n9324_));
  OAI21X1  g08322(.A0(new_n7010_), .A1(new_n6994_), .B0(new_n7008_), .Y(new_n9325_));
  AOI21X1  g08323(.A0(new_n6992_), .A1(new_n9319_), .B0(new_n6991_), .Y(new_n9326_));
  XOR2X1   g08324(.A(new_n9326_), .B(new_n9325_), .Y(new_n9327_));
  AOI21X1  g08325(.A0(new_n9324_), .A1(new_n9318_), .B0(new_n9327_), .Y(new_n9328_));
  AND2X1   g08326(.A(new_n7094_), .B(new_n7093_), .Y(new_n9329_));
  AOI21X1  g08327(.A0(new_n7092_), .A1(new_n7089_), .B0(new_n6993_), .Y(new_n9330_));
  AND2X1   g08328(.A(new_n9326_), .B(new_n9325_), .Y(new_n9331_));
  NOR2X1   g08329(.A(new_n9326_), .B(new_n9325_), .Y(new_n9332_));
  NOR4X1   g08330(.A(new_n9332_), .B(new_n9331_), .C(new_n9330_), .D(new_n9329_), .Y(new_n9333_));
  OR2X1    g08331(.A(new_n9333_), .B(new_n9328_), .Y(new_n9334_));
  OR2X1    g08332(.A(new_n7073_), .B(new_n7072_), .Y(new_n9335_));
  OAI21X1  g08333(.A0(new_n7071_), .A1(new_n7062_), .B0(new_n7061_), .Y(new_n9336_));
  OAI21X1  g08334(.A0(new_n7070_), .A1(new_n7036_), .B0(new_n7069_), .Y(new_n9337_));
  AOI21X1  g08335(.A0(new_n7034_), .A1(new_n7053_), .B0(new_n7033_), .Y(new_n9338_));
  XOR2X1   g08336(.A(new_n9338_), .B(new_n9337_), .Y(new_n9339_));
  AOI21X1  g08337(.A0(new_n9336_), .A1(new_n9335_), .B0(new_n9339_), .Y(new_n9340_));
  AOI21X1  g08338(.A0(new_n7049_), .A1(new_n7043_), .B0(new_n7035_), .Y(new_n9341_));
  NOR2X1   g08339(.A(new_n9338_), .B(new_n9337_), .Y(new_n9342_));
  AOI21X1  g08340(.A0(new_n7048_), .A1(new_n7063_), .B0(new_n7047_), .Y(new_n9343_));
  OAI21X1  g08341(.A0(new_n7060_), .A1(new_n7029_), .B0(new_n7059_), .Y(new_n9344_));
  OAI22X1  g08342(.A0(new_n9344_), .A1(new_n9343_), .B0(new_n7073_), .B1(new_n7072_), .Y(new_n9345_));
  NOR3X1   g08343(.A(new_n9345_), .B(new_n9342_), .C(new_n9341_), .Y(new_n9346_));
  NOR2X1   g08344(.A(new_n9346_), .B(new_n9340_), .Y(new_n9347_));
  XOR2X1   g08345(.A(new_n9347_), .B(new_n9334_), .Y(new_n9348_));
  XOR2X1   g08346(.A(new_n9348_), .B(new_n9317_), .Y(new_n9349_));
  XOR2X1   g08347(.A(new_n9349_), .B(new_n9314_), .Y(new_n9350_));
  XOR2X1   g08348(.A(new_n9350_), .B(new_n9262_), .Y(new_n9351_));
  AND2X1   g08349(.A(new_n6944_), .B(new_n6977_), .Y(new_n9352_));
  AOI21X1  g08350(.A0(new_n9238_), .A1(new_n6921_), .B0(new_n6976_), .Y(new_n9353_));
  OR2X1    g08351(.A(new_n9353_), .B(new_n9352_), .Y(new_n9354_));
  OR2X1    g08352(.A(new_n6779_), .B(new_n6821_), .Y(new_n9355_));
  NOR4X1   g08353(.A(new_n6799_), .B(new_n6786_), .C(new_n6798_), .D(new_n6793_), .Y(new_n9356_));
  XOR2X1   g08354(.A(new_n6810_), .B(new_n9356_), .Y(new_n9357_));
  OR4X1    g08355(.A(new_n6786_), .B(new_n6798_), .C(new_n6809_), .D(new_n6793_), .Y(new_n9358_));
  AND2X1   g08356(.A(new_n6553_), .B(\A[132] ), .Y(new_n9359_));
  OR2X1    g08357(.A(new_n9359_), .B(new_n6555_), .Y(new_n9360_));
  XOR2X1   g08358(.A(new_n6558_), .B(new_n9360_), .Y(new_n9361_));
  XOR2X1   g08359(.A(new_n6788_), .B(new_n9361_), .Y(new_n9362_));
  OAI22X1  g08360(.A0(new_n9362_), .A1(new_n6790_), .B0(new_n6814_), .B1(new_n6793_), .Y(new_n9363_));
  OAI22X1  g08361(.A0(new_n9363_), .A1(new_n9358_), .B0(new_n6810_), .B1(new_n9356_), .Y(new_n9364_));
  MX2X1    g08362(.A(new_n9364_), .B(new_n9357_), .S0(new_n6792_), .Y(new_n9365_));
  OAI21X1  g08363(.A0(new_n6822_), .A1(new_n6763_), .B0(new_n9365_), .Y(new_n9366_));
  AND2X1   g08364(.A(new_n9366_), .B(new_n9355_), .Y(new_n9367_));
  OR2X1    g08365(.A(new_n9363_), .B(new_n9358_), .Y(new_n9368_));
  XOR2X1   g08366(.A(new_n6554_), .B(new_n6548_), .Y(new_n9369_));
  OR2X1    g08367(.A(new_n6554_), .B(new_n6548_), .Y(new_n9370_));
  OR2X1    g08368(.A(new_n6558_), .B(new_n6556_), .Y(new_n9371_));
  OAI21X1  g08369(.A0(new_n9370_), .A1(new_n9361_), .B0(new_n9371_), .Y(new_n9372_));
  AOI21X1  g08370(.A0(new_n9372_), .A1(new_n9369_), .B0(new_n9362_), .Y(new_n9373_));
  OAI21X1  g08371(.A0(new_n6810_), .A1(new_n9356_), .B0(new_n9373_), .Y(new_n9374_));
  OAI21X1  g08372(.A0(new_n6809_), .A1(new_n6793_), .B0(new_n6807_), .Y(new_n9375_));
  AOI21X1  g08373(.A0(new_n6791_), .A1(new_n9369_), .B0(new_n6790_), .Y(new_n9376_));
  XOR2X1   g08374(.A(new_n9376_), .B(new_n9375_), .Y(new_n9377_));
  AOI21X1  g08375(.A0(new_n9374_), .A1(new_n9368_), .B0(new_n9377_), .Y(new_n9378_));
  AND2X1   g08376(.A(new_n6818_), .B(new_n6817_), .Y(new_n9379_));
  AOI21X1  g08377(.A0(new_n6816_), .A1(new_n6800_), .B0(new_n6792_), .Y(new_n9380_));
  AND2X1   g08378(.A(new_n9376_), .B(new_n9375_), .Y(new_n9381_));
  NOR2X1   g08379(.A(new_n9376_), .B(new_n9375_), .Y(new_n9382_));
  NOR4X1   g08380(.A(new_n9382_), .B(new_n9381_), .C(new_n9380_), .D(new_n9379_), .Y(new_n9383_));
  NOR2X1   g08381(.A(new_n9383_), .B(new_n9378_), .Y(new_n9384_));
  OR2X1    g08382(.A(new_n6969_), .B(new_n6968_), .Y(new_n9385_));
  OAI21X1  g08383(.A0(new_n6777_), .A1(new_n6967_), .B0(new_n6966_), .Y(new_n9386_));
  OAI21X1  g08384(.A0(new_n6771_), .A1(new_n6748_), .B0(new_n6770_), .Y(new_n9387_));
  AOI21X1  g08385(.A0(new_n6746_), .A1(new_n6958_), .B0(new_n6745_), .Y(new_n9388_));
  XOR2X1   g08386(.A(new_n9388_), .B(new_n9387_), .Y(new_n9389_));
  AOI21X1  g08387(.A0(new_n9386_), .A1(new_n9385_), .B0(new_n9389_), .Y(new_n9390_));
  AOI21X1  g08388(.A0(new_n6761_), .A1(new_n6755_), .B0(new_n6747_), .Y(new_n9391_));
  NOR2X1   g08389(.A(new_n9388_), .B(new_n9387_), .Y(new_n9392_));
  AOI21X1  g08390(.A0(new_n6760_), .A1(new_n6773_), .B0(new_n6759_), .Y(new_n9393_));
  OAI21X1  g08391(.A0(new_n6965_), .A1(new_n6741_), .B0(new_n6964_), .Y(new_n9394_));
  OAI22X1  g08392(.A0(new_n9394_), .A1(new_n9393_), .B0(new_n6969_), .B1(new_n6968_), .Y(new_n9395_));
  NOR3X1   g08393(.A(new_n9395_), .B(new_n9392_), .C(new_n9391_), .Y(new_n9396_));
  NOR2X1   g08394(.A(new_n9396_), .B(new_n9390_), .Y(new_n9397_));
  XOR2X1   g08395(.A(new_n9397_), .B(new_n9384_), .Y(new_n9398_));
  XOR2X1   g08396(.A(new_n9398_), .B(new_n9367_), .Y(new_n9399_));
  OR2X1    g08397(.A(new_n6929_), .B(new_n6895_), .Y(new_n9400_));
  OAI21X1  g08398(.A0(new_n6930_), .A1(new_n6924_), .B0(new_n6866_), .Y(new_n9401_));
  AND2X1   g08399(.A(new_n9401_), .B(new_n9400_), .Y(new_n9402_));
  OR2X1    g08400(.A(new_n6864_), .B(new_n6856_), .Y(new_n9403_));
  XOR2X1   g08401(.A(new_n6480_), .B(new_n6474_), .Y(new_n9404_));
  OR2X1    g08402(.A(new_n6480_), .B(new_n6474_), .Y(new_n9405_));
  OR2X1    g08403(.A(new_n6484_), .B(new_n6482_), .Y(new_n9406_));
  OAI21X1  g08404(.A0(new_n9405_), .A1(new_n6862_), .B0(new_n9406_), .Y(new_n9407_));
  AOI21X1  g08405(.A0(new_n9407_), .A1(new_n9404_), .B0(new_n6863_), .Y(new_n9408_));
  OAI21X1  g08406(.A0(new_n6854_), .A1(new_n6844_), .B0(new_n9408_), .Y(new_n9409_));
  OAI21X1  g08407(.A0(new_n6853_), .A1(new_n6837_), .B0(new_n6851_), .Y(new_n9410_));
  AOI21X1  g08408(.A0(new_n6835_), .A1(new_n9404_), .B0(new_n6834_), .Y(new_n9411_));
  XOR2X1   g08409(.A(new_n9411_), .B(new_n9410_), .Y(new_n9412_));
  AOI21X1  g08410(.A0(new_n9409_), .A1(new_n9403_), .B0(new_n9412_), .Y(new_n9413_));
  AND2X1   g08411(.A(new_n6938_), .B(new_n6937_), .Y(new_n9414_));
  AOI21X1  g08412(.A0(new_n6936_), .A1(new_n6933_), .B0(new_n6836_), .Y(new_n9415_));
  AND2X1   g08413(.A(new_n9411_), .B(new_n9410_), .Y(new_n9416_));
  NOR2X1   g08414(.A(new_n9411_), .B(new_n9410_), .Y(new_n9417_));
  NOR4X1   g08415(.A(new_n9417_), .B(new_n9416_), .C(new_n9415_), .D(new_n9414_), .Y(new_n9418_));
  OR2X1    g08416(.A(new_n9418_), .B(new_n9413_), .Y(new_n9419_));
  OR2X1    g08417(.A(new_n6916_), .B(new_n6915_), .Y(new_n9420_));
  OAI21X1  g08418(.A0(new_n6914_), .A1(new_n6905_), .B0(new_n6904_), .Y(new_n9421_));
  OAI21X1  g08419(.A0(new_n6913_), .A1(new_n6879_), .B0(new_n6912_), .Y(new_n9422_));
  AOI21X1  g08420(.A0(new_n6877_), .A1(new_n6896_), .B0(new_n6876_), .Y(new_n9423_));
  XOR2X1   g08421(.A(new_n9423_), .B(new_n9422_), .Y(new_n9424_));
  AOI21X1  g08422(.A0(new_n9421_), .A1(new_n9420_), .B0(new_n9424_), .Y(new_n9425_));
  AOI21X1  g08423(.A0(new_n6892_), .A1(new_n6886_), .B0(new_n6878_), .Y(new_n9426_));
  NOR2X1   g08424(.A(new_n9423_), .B(new_n9422_), .Y(new_n9427_));
  AOI21X1  g08425(.A0(new_n6891_), .A1(new_n6906_), .B0(new_n6890_), .Y(new_n9428_));
  OAI21X1  g08426(.A0(new_n6903_), .A1(new_n6872_), .B0(new_n6902_), .Y(new_n9429_));
  OAI22X1  g08427(.A0(new_n9429_), .A1(new_n9428_), .B0(new_n6916_), .B1(new_n6915_), .Y(new_n9430_));
  NOR3X1   g08428(.A(new_n9430_), .B(new_n9427_), .C(new_n9426_), .Y(new_n9431_));
  NOR2X1   g08429(.A(new_n9431_), .B(new_n9425_), .Y(new_n9432_));
  XOR2X1   g08430(.A(new_n9432_), .B(new_n9419_), .Y(new_n9433_));
  XOR2X1   g08431(.A(new_n9433_), .B(new_n9402_), .Y(new_n9434_));
  XOR2X1   g08432(.A(new_n9434_), .B(new_n9399_), .Y(new_n9435_));
  XOR2X1   g08433(.A(new_n9435_), .B(new_n9354_), .Y(new_n9436_));
  XOR2X1   g08434(.A(new_n9436_), .B(new_n9351_), .Y(new_n9437_));
  XOR2X1   g08435(.A(new_n9437_), .B(new_n9259_), .Y(new_n9438_));
  AND2X1   g08436(.A(new_n6411_), .B(new_n6731_), .Y(new_n9439_));
  AOI21X1  g08437(.A0(new_n8812_), .A1(new_n6371_), .B0(new_n6730_), .Y(new_n9440_));
  OR2X1    g08438(.A(new_n9440_), .B(new_n9439_), .Y(new_n9441_));
  AND2X1   g08439(.A(new_n6726_), .B(new_n5886_), .Y(new_n9442_));
  AOI21X1  g08440(.A0(new_n6728_), .A1(new_n6722_), .B0(new_n6009_), .Y(new_n9443_));
  OR2X1    g08441(.A(new_n9443_), .B(new_n9442_), .Y(new_n9444_));
  XOR2X1   g08442(.A(new_n5959_), .B(new_n5931_), .Y(new_n9445_));
  NOR4X1   g08443(.A(new_n5917_), .B(new_n5958_), .C(new_n5957_), .D(new_n5924_), .Y(new_n9446_));
  AOI21X1  g08444(.A0(new_n5957_), .A1(new_n5951_), .B0(new_n5930_), .Y(new_n9447_));
  AOI22X1  g08445(.A0(new_n9447_), .A1(new_n9446_), .B0(new_n5937_), .B1(new_n5931_), .Y(new_n9448_));
  MX2X1    g08446(.A(new_n9448_), .B(new_n9445_), .S0(new_n5923_), .Y(new_n9449_));
  OR2X1    g08447(.A(new_n9449_), .B(new_n5940_), .Y(new_n9450_));
  AND2X1   g08448(.A(new_n5938_), .B(new_n5923_), .Y(new_n9451_));
  NOR4X1   g08449(.A(new_n5984_), .B(new_n5971_), .C(new_n5983_), .D(new_n5978_), .Y(new_n9452_));
  XOR2X1   g08450(.A(new_n5995_), .B(new_n9452_), .Y(new_n9453_));
  OR4X1    g08451(.A(new_n5971_), .B(new_n5983_), .C(new_n5994_), .D(new_n5978_), .Y(new_n9454_));
  AND2X1   g08452(.A(new_n5877_), .B(\A[180] ), .Y(new_n9455_));
  OR2X1    g08453(.A(new_n9455_), .B(new_n5879_), .Y(new_n9456_));
  XOR2X1   g08454(.A(new_n5882_), .B(new_n9456_), .Y(new_n9457_));
  XOR2X1   g08455(.A(new_n5973_), .B(new_n9457_), .Y(new_n9458_));
  OAI22X1  g08456(.A0(new_n9458_), .A1(new_n5975_), .B0(new_n5999_), .B1(new_n5978_), .Y(new_n9459_));
  OAI22X1  g08457(.A0(new_n9459_), .A1(new_n9454_), .B0(new_n5995_), .B1(new_n9452_), .Y(new_n9460_));
  MX2X1    g08458(.A(new_n9460_), .B(new_n9453_), .S0(new_n5977_), .Y(new_n9461_));
  OAI21X1  g08459(.A0(new_n9448_), .A1(new_n5923_), .B0(new_n5940_), .Y(new_n9462_));
  OAI21X1  g08460(.A0(new_n9462_), .A1(new_n9451_), .B0(new_n9461_), .Y(new_n9463_));
  AND2X1   g08461(.A(new_n9463_), .B(new_n9450_), .Y(new_n9464_));
  OR2X1    g08462(.A(new_n9459_), .B(new_n9454_), .Y(new_n9465_));
  XOR2X1   g08463(.A(new_n5878_), .B(new_n5872_), .Y(new_n9466_));
  OR2X1    g08464(.A(new_n5878_), .B(new_n5872_), .Y(new_n9467_));
  OR2X1    g08465(.A(new_n5882_), .B(new_n5880_), .Y(new_n9468_));
  OAI21X1  g08466(.A0(new_n9467_), .A1(new_n9457_), .B0(new_n9468_), .Y(new_n9469_));
  AOI21X1  g08467(.A0(new_n9469_), .A1(new_n9466_), .B0(new_n9458_), .Y(new_n9470_));
  OAI21X1  g08468(.A0(new_n5995_), .A1(new_n9452_), .B0(new_n9470_), .Y(new_n9471_));
  OAI21X1  g08469(.A0(new_n5994_), .A1(new_n5978_), .B0(new_n5992_), .Y(new_n9472_));
  AOI21X1  g08470(.A0(new_n5976_), .A1(new_n9466_), .B0(new_n5975_), .Y(new_n9473_));
  XOR2X1   g08471(.A(new_n9473_), .B(new_n9472_), .Y(new_n9474_));
  AOI21X1  g08472(.A0(new_n9471_), .A1(new_n9465_), .B0(new_n9474_), .Y(new_n9475_));
  AND2X1   g08473(.A(new_n6003_), .B(new_n6002_), .Y(new_n9476_));
  AOI21X1  g08474(.A0(new_n6001_), .A1(new_n5985_), .B0(new_n5977_), .Y(new_n9477_));
  AND2X1   g08475(.A(new_n9473_), .B(new_n9472_), .Y(new_n9478_));
  NOR2X1   g08476(.A(new_n9473_), .B(new_n9472_), .Y(new_n9479_));
  NOR4X1   g08477(.A(new_n9479_), .B(new_n9478_), .C(new_n9477_), .D(new_n9476_), .Y(new_n9480_));
  NOR2X1   g08478(.A(new_n9480_), .B(new_n9475_), .Y(new_n9481_));
  OR2X1    g08479(.A(new_n5961_), .B(new_n5960_), .Y(new_n9482_));
  OAI21X1  g08480(.A0(new_n5959_), .A1(new_n5950_), .B0(new_n5949_), .Y(new_n9483_));
  OAI21X1  g08481(.A0(new_n5958_), .A1(new_n5924_), .B0(new_n5957_), .Y(new_n9484_));
  AOI21X1  g08482(.A0(new_n5922_), .A1(new_n5941_), .B0(new_n5921_), .Y(new_n9485_));
  XOR2X1   g08483(.A(new_n9485_), .B(new_n9484_), .Y(new_n9486_));
  AOI21X1  g08484(.A0(new_n9483_), .A1(new_n9482_), .B0(new_n9486_), .Y(new_n9487_));
  AOI21X1  g08485(.A0(new_n5937_), .A1(new_n5931_), .B0(new_n5923_), .Y(new_n9488_));
  NOR2X1   g08486(.A(new_n9485_), .B(new_n9484_), .Y(new_n9489_));
  AOI21X1  g08487(.A0(new_n5936_), .A1(new_n5951_), .B0(new_n5935_), .Y(new_n9490_));
  OAI21X1  g08488(.A0(new_n5948_), .A1(new_n5917_), .B0(new_n5947_), .Y(new_n9491_));
  OAI22X1  g08489(.A0(new_n9491_), .A1(new_n9490_), .B0(new_n5961_), .B1(new_n5960_), .Y(new_n9492_));
  NOR3X1   g08490(.A(new_n9492_), .B(new_n9489_), .C(new_n9488_), .Y(new_n9493_));
  NOR2X1   g08491(.A(new_n9493_), .B(new_n9487_), .Y(new_n9494_));
  XOR2X1   g08492(.A(new_n9494_), .B(new_n9481_), .Y(new_n9495_));
  XOR2X1   g08493(.A(new_n9495_), .B(new_n9464_), .Y(new_n9496_));
  OR2X1    g08494(.A(new_n5806_), .B(new_n5907_), .Y(new_n9497_));
  OAI21X1  g08495(.A0(new_n6723_), .A1(new_n5784_), .B0(new_n5906_), .Y(new_n9498_));
  AND2X1   g08496(.A(new_n9498_), .B(new_n9497_), .Y(new_n9499_));
  OR2X1    g08497(.A(new_n5904_), .B(new_n5903_), .Y(new_n9500_));
  XOR2X1   g08498(.A(new_n5661_), .B(new_n5669_), .Y(new_n9501_));
  XOR2X1   g08499(.A(new_n5654_), .B(new_n5648_), .Y(new_n9502_));
  OR2X1    g08500(.A(new_n5660_), .B(new_n5670_), .Y(new_n9503_));
  OAI21X1  g08501(.A0(new_n5661_), .A1(new_n5655_), .B0(new_n9503_), .Y(new_n9504_));
  AOI21X1  g08502(.A0(new_n9504_), .A1(new_n9502_), .B0(new_n9501_), .Y(new_n9505_));
  OAI21X1  g08503(.A0(new_n5709_), .A1(new_n5901_), .B0(new_n9505_), .Y(new_n9506_));
  OAI21X1  g08504(.A0(new_n5698_), .A1(new_n5707_), .B0(new_n5705_), .Y(new_n9507_));
  AOI21X1  g08505(.A0(new_n9502_), .A1(new_n5662_), .B0(new_n5673_), .Y(new_n9508_));
  XOR2X1   g08506(.A(new_n9508_), .B(new_n9507_), .Y(new_n9509_));
  AOI21X1  g08507(.A0(new_n9506_), .A1(new_n9500_), .B0(new_n9509_), .Y(new_n9510_));
  AND2X1   g08508(.A(new_n5717_), .B(new_n5716_), .Y(new_n9511_));
  AOI21X1  g08509(.A0(new_n5715_), .A1(new_n5699_), .B0(new_n5674_), .Y(new_n9512_));
  AND2X1   g08510(.A(new_n9508_), .B(new_n9507_), .Y(new_n9513_));
  NOR2X1   g08511(.A(new_n9508_), .B(new_n9507_), .Y(new_n9514_));
  NOR4X1   g08512(.A(new_n9514_), .B(new_n9513_), .C(new_n9512_), .D(new_n9511_), .Y(new_n9515_));
  OR2X1    g08513(.A(new_n9515_), .B(new_n9510_), .Y(new_n9516_));
  OR2X1    g08514(.A(new_n5890_), .B(new_n5889_), .Y(new_n9517_));
  OAI21X1  g08515(.A0(new_n5804_), .A1(new_n5888_), .B0(new_n5897_), .Y(new_n9518_));
  OAI21X1  g08516(.A0(new_n5775_), .A1(new_n5795_), .B0(new_n5799_), .Y(new_n9519_));
  AOI21X1  g08517(.A0(new_n5894_), .A1(new_n5739_), .B0(new_n5750_), .Y(new_n9520_));
  XOR2X1   g08518(.A(new_n9520_), .B(new_n9519_), .Y(new_n9521_));
  AOI21X1  g08519(.A0(new_n9518_), .A1(new_n9517_), .B0(new_n9521_), .Y(new_n9522_));
  AOI21X1  g08520(.A0(new_n5782_), .A1(new_n5776_), .B0(new_n5751_), .Y(new_n9523_));
  NOR2X1   g08521(.A(new_n9520_), .B(new_n9519_), .Y(new_n9524_));
  AOI21X1  g08522(.A0(new_n5800_), .A1(new_n5781_), .B0(new_n5780_), .Y(new_n9525_));
  OAI21X1  g08523(.A0(new_n5745_), .A1(new_n5893_), .B0(new_n5896_), .Y(new_n9526_));
  OAI22X1  g08524(.A0(new_n9526_), .A1(new_n9525_), .B0(new_n5890_), .B1(new_n5889_), .Y(new_n9527_));
  NOR3X1   g08525(.A(new_n9527_), .B(new_n9524_), .C(new_n9523_), .Y(new_n9528_));
  NOR2X1   g08526(.A(new_n9528_), .B(new_n9522_), .Y(new_n9529_));
  XOR2X1   g08527(.A(new_n9529_), .B(new_n9516_), .Y(new_n9530_));
  XOR2X1   g08528(.A(new_n9530_), .B(new_n9499_), .Y(new_n9531_));
  XOR2X1   g08529(.A(new_n9531_), .B(new_n9496_), .Y(new_n9532_));
  XOR2X1   g08530(.A(new_n9532_), .B(new_n9444_), .Y(new_n9533_));
  OR2X1    g08531(.A(new_n6388_), .B(new_n6356_), .Y(new_n9534_));
  OAI21X1  g08532(.A0(new_n6389_), .A1(new_n6385_), .B0(new_n6181_), .Y(new_n9535_));
  AND2X1   g08533(.A(new_n9535_), .B(new_n9534_), .Y(new_n9536_));
  OR2X1    g08534(.A(new_n6135_), .B(new_n6178_), .Y(new_n9537_));
  NOR4X1   g08535(.A(new_n6155_), .B(new_n6142_), .C(new_n6154_), .D(new_n6149_), .Y(new_n9538_));
  XOR2X1   g08536(.A(new_n6166_), .B(new_n9538_), .Y(new_n9539_));
  OR4X1    g08537(.A(new_n6142_), .B(new_n6154_), .C(new_n6165_), .D(new_n6149_), .Y(new_n9540_));
  AND2X1   g08538(.A(new_n6113_), .B(\A[228] ), .Y(new_n9541_));
  OR2X1    g08539(.A(new_n9541_), .B(new_n6115_), .Y(new_n9542_));
  XOR2X1   g08540(.A(new_n6118_), .B(new_n9542_), .Y(new_n9543_));
  XOR2X1   g08541(.A(new_n6144_), .B(new_n9543_), .Y(new_n9544_));
  OAI22X1  g08542(.A0(new_n9544_), .A1(new_n6146_), .B0(new_n6170_), .B1(new_n6149_), .Y(new_n9545_));
  OAI22X1  g08543(.A0(new_n9545_), .A1(new_n9540_), .B0(new_n6166_), .B1(new_n9538_), .Y(new_n9546_));
  MX2X1    g08544(.A(new_n9546_), .B(new_n9539_), .S0(new_n6148_), .Y(new_n9547_));
  OAI21X1  g08545(.A0(new_n6179_), .A1(new_n6078_), .B0(new_n9547_), .Y(new_n9548_));
  AND2X1   g08546(.A(new_n9548_), .B(new_n9537_), .Y(new_n9549_));
  OR2X1    g08547(.A(new_n9545_), .B(new_n9540_), .Y(new_n9550_));
  XOR2X1   g08548(.A(new_n6114_), .B(new_n6108_), .Y(new_n9551_));
  OR2X1    g08549(.A(new_n6114_), .B(new_n6108_), .Y(new_n9552_));
  OR2X1    g08550(.A(new_n6118_), .B(new_n6116_), .Y(new_n9553_));
  OAI21X1  g08551(.A0(new_n9552_), .A1(new_n9543_), .B0(new_n9553_), .Y(new_n9554_));
  AOI21X1  g08552(.A0(new_n9554_), .A1(new_n9551_), .B0(new_n9544_), .Y(new_n9555_));
  OAI21X1  g08553(.A0(new_n6166_), .A1(new_n9538_), .B0(new_n9555_), .Y(new_n9556_));
  OAI21X1  g08554(.A0(new_n6165_), .A1(new_n6149_), .B0(new_n6163_), .Y(new_n9557_));
  AOI21X1  g08555(.A0(new_n6147_), .A1(new_n9551_), .B0(new_n6146_), .Y(new_n9558_));
  XOR2X1   g08556(.A(new_n9558_), .B(new_n9557_), .Y(new_n9559_));
  AOI21X1  g08557(.A0(new_n9556_), .A1(new_n9550_), .B0(new_n9559_), .Y(new_n9560_));
  AOI21X1  g08558(.A0(new_n6172_), .A1(new_n6156_), .B0(new_n6148_), .Y(new_n9561_));
  NOR2X1   g08559(.A(new_n9558_), .B(new_n9557_), .Y(new_n9562_));
  AOI21X1  g08560(.A0(new_n6171_), .A1(new_n6157_), .B0(new_n6170_), .Y(new_n9563_));
  OAI21X1  g08561(.A0(new_n9544_), .A1(new_n6142_), .B0(new_n9554_), .Y(new_n9564_));
  OAI22X1  g08562(.A0(new_n9564_), .A1(new_n9563_), .B0(new_n9545_), .B1(new_n9540_), .Y(new_n9565_));
  NOR3X1   g08563(.A(new_n9565_), .B(new_n9562_), .C(new_n9561_), .Y(new_n9566_));
  NOR2X1   g08564(.A(new_n9566_), .B(new_n9560_), .Y(new_n9567_));
  OR2X1    g08565(.A(new_n6400_), .B(new_n6399_), .Y(new_n9568_));
  OAI21X1  g08566(.A0(new_n6133_), .A1(new_n6398_), .B0(new_n6397_), .Y(new_n9569_));
  OAI21X1  g08567(.A0(new_n6069_), .A1(new_n6125_), .B0(new_n6129_), .Y(new_n9570_));
  AOI21X1  g08568(.A0(new_n6394_), .A1(new_n6033_), .B0(new_n6044_), .Y(new_n9571_));
  XOR2X1   g08569(.A(new_n9571_), .B(new_n9570_), .Y(new_n9572_));
  AOI21X1  g08570(.A0(new_n9569_), .A1(new_n9568_), .B0(new_n9572_), .Y(new_n9573_));
  AOI21X1  g08571(.A0(new_n6076_), .A1(new_n6070_), .B0(new_n6045_), .Y(new_n9574_));
  NOR2X1   g08572(.A(new_n9571_), .B(new_n9570_), .Y(new_n9575_));
  AOI21X1  g08573(.A0(new_n6082_), .A1(new_n6075_), .B0(new_n6074_), .Y(new_n9576_));
  OAI21X1  g08574(.A0(new_n6039_), .A1(new_n6393_), .B0(new_n6396_), .Y(new_n9577_));
  OAI22X1  g08575(.A0(new_n9577_), .A1(new_n9576_), .B0(new_n6400_), .B1(new_n6399_), .Y(new_n9578_));
  NOR3X1   g08576(.A(new_n9578_), .B(new_n9575_), .C(new_n9574_), .Y(new_n9579_));
  NOR2X1   g08577(.A(new_n9579_), .B(new_n9573_), .Y(new_n9580_));
  XOR2X1   g08578(.A(new_n9580_), .B(new_n9567_), .Y(new_n9581_));
  XOR2X1   g08579(.A(new_n9581_), .B(new_n9549_), .Y(new_n9582_));
  OR2X1    g08580(.A(new_n6362_), .B(new_n6328_), .Y(new_n9583_));
  OAI21X1  g08581(.A0(new_n6363_), .A1(new_n6357_), .B0(new_n6256_), .Y(new_n9584_));
  AND2X1   g08582(.A(new_n9584_), .B(new_n9583_), .Y(new_n9585_));
  OR2X1    g08583(.A(new_n6254_), .B(new_n6250_), .Y(new_n9586_));
  XOR2X1   g08584(.A(new_n6200_), .B(new_n6208_), .Y(new_n9587_));
  XOR2X1   g08585(.A(new_n6193_), .B(new_n6187_), .Y(new_n9588_));
  OR2X1    g08586(.A(new_n6199_), .B(new_n6209_), .Y(new_n9589_));
  OAI21X1  g08587(.A0(new_n6200_), .A1(new_n6194_), .B0(new_n9589_), .Y(new_n9590_));
  AOI21X1  g08588(.A0(new_n9590_), .A1(new_n9588_), .B0(new_n9587_), .Y(new_n9591_));
  OAI21X1  g08589(.A0(new_n6248_), .A1(new_n6238_), .B0(new_n9591_), .Y(new_n9592_));
  OAI21X1  g08590(.A0(new_n6237_), .A1(new_n6246_), .B0(new_n6244_), .Y(new_n9593_));
  AOI21X1  g08591(.A0(new_n9588_), .A1(new_n6201_), .B0(new_n6212_), .Y(new_n9594_));
  XOR2X1   g08592(.A(new_n9594_), .B(new_n9593_), .Y(new_n9595_));
  AOI21X1  g08593(.A0(new_n9592_), .A1(new_n9586_), .B0(new_n9595_), .Y(new_n9596_));
  AND2X1   g08594(.A(new_n6382_), .B(new_n6381_), .Y(new_n9597_));
  AOI21X1  g08595(.A0(new_n6380_), .A1(new_n6377_), .B0(new_n6213_), .Y(new_n9598_));
  AND2X1   g08596(.A(new_n9594_), .B(new_n9593_), .Y(new_n9599_));
  NOR2X1   g08597(.A(new_n9594_), .B(new_n9593_), .Y(new_n9600_));
  NOR4X1   g08598(.A(new_n9600_), .B(new_n9599_), .C(new_n9598_), .D(new_n9597_), .Y(new_n9601_));
  OR2X1    g08599(.A(new_n9601_), .B(new_n9596_), .Y(new_n9602_));
  OR2X1    g08600(.A(new_n6345_), .B(new_n6344_), .Y(new_n9603_));
  OAI21X1  g08601(.A0(new_n6343_), .A1(new_n6334_), .B0(new_n6333_), .Y(new_n9604_));
  OAI21X1  g08602(.A0(new_n6312_), .A1(new_n6341_), .B0(new_n6340_), .Y(new_n9605_));
  AOI21X1  g08603(.A0(new_n6330_), .A1(new_n6276_), .B0(new_n6287_), .Y(new_n9606_));
  XOR2X1   g08604(.A(new_n9606_), .B(new_n9605_), .Y(new_n9607_));
  AOI21X1  g08605(.A0(new_n9604_), .A1(new_n9603_), .B0(new_n9607_), .Y(new_n9608_));
  AOI21X1  g08606(.A0(new_n6319_), .A1(new_n6313_), .B0(new_n6288_), .Y(new_n9609_));
  NOR2X1   g08607(.A(new_n9606_), .B(new_n9605_), .Y(new_n9610_));
  AOI21X1  g08608(.A0(new_n6342_), .A1(new_n6318_), .B0(new_n6317_), .Y(new_n9611_));
  OAI21X1  g08609(.A0(new_n6282_), .A1(new_n6329_), .B0(new_n6332_), .Y(new_n9612_));
  OAI22X1  g08610(.A0(new_n9612_), .A1(new_n9611_), .B0(new_n6345_), .B1(new_n6344_), .Y(new_n9613_));
  NOR3X1   g08611(.A(new_n9613_), .B(new_n9610_), .C(new_n9609_), .Y(new_n9614_));
  NOR2X1   g08612(.A(new_n9614_), .B(new_n9608_), .Y(new_n9615_));
  XOR2X1   g08613(.A(new_n9615_), .B(new_n9602_), .Y(new_n9616_));
  XOR2X1   g08614(.A(new_n9616_), .B(new_n9585_), .Y(new_n9617_));
  XOR2X1   g08615(.A(new_n9617_), .B(new_n9582_), .Y(new_n9618_));
  XOR2X1   g08616(.A(new_n9618_), .B(new_n9536_), .Y(new_n9619_));
  XOR2X1   g08617(.A(new_n9619_), .B(new_n9533_), .Y(new_n9620_));
  XOR2X1   g08618(.A(new_n9620_), .B(new_n9441_), .Y(new_n9621_));
  XOR2X1   g08619(.A(new_n9621_), .B(new_n9438_), .Y(new_n9622_));
  XOR2X1   g08620(.A(new_n9622_), .B(new_n9247_), .Y(new_n9623_));
  OR2X1    g08621(.A(new_n8767_), .B(new_n8770_), .Y(new_n9624_));
  OAI21X1  g08622(.A0(new_n8771_), .A1(new_n8722_), .B0(new_n7970_), .Y(new_n9625_));
  AND2X1   g08623(.A(new_n9625_), .B(new_n9624_), .Y(new_n9626_));
  OR2X1    g08624(.A(new_n7742_), .B(new_n7967_), .Y(new_n9627_));
  AND2X1   g08625(.A(new_n7862_), .B(new_n7859_), .Y(new_n9628_));
  AOI21X1  g08626(.A0(new_n7836_), .A1(new_n7823_), .B0(new_n7860_), .Y(new_n9629_));
  AOI22X1  g08627(.A0(new_n9629_), .A1(new_n7813_), .B0(new_n7838_), .B1(new_n7860_), .Y(new_n9630_));
  OAI21X1  g08628(.A0(new_n9630_), .A1(new_n7859_), .B0(new_n7963_), .Y(new_n9631_));
  MX2X1    g08629(.A(new_n9630_), .B(new_n7839_), .S0(new_n7859_), .Y(new_n9632_));
  OAI22X1  g08630(.A0(new_n9632_), .A1(new_n7963_), .B0(new_n9631_), .B1(new_n9628_), .Y(new_n9633_));
  OAI21X1  g08631(.A0(new_n9630_), .A1(new_n7859_), .B0(new_n7842_), .Y(new_n9634_));
  OAI22X1  g08632(.A0(new_n9634_), .A1(new_n9628_), .B0(new_n9632_), .B1(new_n7842_), .Y(new_n9635_));
  MX2X1    g08633(.A(new_n9635_), .B(new_n9633_), .S0(new_n7962_), .Y(new_n9636_));
  OAI21X1  g08634(.A0(new_n7968_), .A1(new_n7580_), .B0(new_n9636_), .Y(new_n9637_));
  AND2X1   g08635(.A(new_n9637_), .B(new_n9627_), .Y(new_n9638_));
  AND2X1   g08636(.A(new_n7863_), .B(new_n7963_), .Y(new_n9639_));
  AOI21X1  g08637(.A0(new_n7964_), .A1(new_n7840_), .B0(new_n7962_), .Y(new_n9640_));
  OR2X1    g08638(.A(new_n9640_), .B(new_n9639_), .Y(new_n9641_));
  XOR2X1   g08639(.A(new_n7912_), .B(new_n7884_), .Y(new_n9642_));
  NOR4X1   g08640(.A(new_n7870_), .B(new_n7911_), .C(new_n7910_), .D(new_n7877_), .Y(new_n9643_));
  AOI21X1  g08641(.A0(new_n7910_), .A1(new_n7904_), .B0(new_n7883_), .Y(new_n9644_));
  AOI22X1  g08642(.A0(new_n9644_), .A1(new_n9643_), .B0(new_n7890_), .B1(new_n7884_), .Y(new_n9645_));
  MX2X1    g08643(.A(new_n9645_), .B(new_n9642_), .S0(new_n7876_), .Y(new_n9646_));
  OR2X1    g08644(.A(new_n9646_), .B(new_n7893_), .Y(new_n9647_));
  AND2X1   g08645(.A(new_n7891_), .B(new_n7876_), .Y(new_n9648_));
  NOR4X1   g08646(.A(new_n7937_), .B(new_n7924_), .C(new_n7936_), .D(new_n7931_), .Y(new_n9649_));
  XOR2X1   g08647(.A(new_n7948_), .B(new_n9649_), .Y(new_n9650_));
  OR4X1    g08648(.A(new_n7924_), .B(new_n7936_), .C(new_n7947_), .D(new_n7931_), .Y(new_n9651_));
  AND2X1   g08649(.A(new_n7721_), .B(\A[276] ), .Y(new_n9652_));
  OR2X1    g08650(.A(new_n9652_), .B(new_n7723_), .Y(new_n9653_));
  XOR2X1   g08651(.A(new_n7726_), .B(new_n9653_), .Y(new_n9654_));
  XOR2X1   g08652(.A(new_n7926_), .B(new_n9654_), .Y(new_n9655_));
  OAI22X1  g08653(.A0(new_n9655_), .A1(new_n7928_), .B0(new_n7952_), .B1(new_n7931_), .Y(new_n9656_));
  OAI22X1  g08654(.A0(new_n9656_), .A1(new_n9651_), .B0(new_n7948_), .B1(new_n9649_), .Y(new_n9657_));
  MX2X1    g08655(.A(new_n9657_), .B(new_n9650_), .S0(new_n7930_), .Y(new_n9658_));
  OAI21X1  g08656(.A0(new_n9645_), .A1(new_n7876_), .B0(new_n7893_), .Y(new_n9659_));
  OAI21X1  g08657(.A0(new_n9659_), .A1(new_n9648_), .B0(new_n9658_), .Y(new_n9660_));
  AND2X1   g08658(.A(new_n9660_), .B(new_n9647_), .Y(new_n9661_));
  OR2X1    g08659(.A(new_n9656_), .B(new_n9651_), .Y(new_n9662_));
  XOR2X1   g08660(.A(new_n7722_), .B(new_n7716_), .Y(new_n9663_));
  OR2X1    g08661(.A(new_n7722_), .B(new_n7716_), .Y(new_n9664_));
  OR2X1    g08662(.A(new_n7726_), .B(new_n7724_), .Y(new_n9665_));
  OAI21X1  g08663(.A0(new_n9664_), .A1(new_n9654_), .B0(new_n9665_), .Y(new_n9666_));
  AOI21X1  g08664(.A0(new_n9666_), .A1(new_n9663_), .B0(new_n9655_), .Y(new_n9667_));
  OAI21X1  g08665(.A0(new_n7948_), .A1(new_n9649_), .B0(new_n9667_), .Y(new_n9668_));
  OAI21X1  g08666(.A0(new_n7947_), .A1(new_n7931_), .B0(new_n7945_), .Y(new_n9669_));
  AOI21X1  g08667(.A0(new_n7929_), .A1(new_n9663_), .B0(new_n7928_), .Y(new_n9670_));
  XOR2X1   g08668(.A(new_n9670_), .B(new_n9669_), .Y(new_n9671_));
  AOI21X1  g08669(.A0(new_n9668_), .A1(new_n9662_), .B0(new_n9671_), .Y(new_n9672_));
  AND2X1   g08670(.A(new_n7956_), .B(new_n7955_), .Y(new_n9673_));
  AOI21X1  g08671(.A0(new_n7954_), .A1(new_n7938_), .B0(new_n7930_), .Y(new_n9674_));
  AND2X1   g08672(.A(new_n9670_), .B(new_n9669_), .Y(new_n9675_));
  NOR2X1   g08673(.A(new_n9670_), .B(new_n9669_), .Y(new_n9676_));
  NOR4X1   g08674(.A(new_n9676_), .B(new_n9675_), .C(new_n9674_), .D(new_n9673_), .Y(new_n9677_));
  NOR2X1   g08675(.A(new_n9677_), .B(new_n9672_), .Y(new_n9678_));
  OR2X1    g08676(.A(new_n7914_), .B(new_n7913_), .Y(new_n9679_));
  OAI21X1  g08677(.A0(new_n7912_), .A1(new_n7903_), .B0(new_n7902_), .Y(new_n9680_));
  OAI21X1  g08678(.A0(new_n7911_), .A1(new_n7877_), .B0(new_n7910_), .Y(new_n9681_));
  AOI21X1  g08679(.A0(new_n7875_), .A1(new_n7894_), .B0(new_n7874_), .Y(new_n9682_));
  XOR2X1   g08680(.A(new_n9682_), .B(new_n9681_), .Y(new_n9683_));
  AOI21X1  g08681(.A0(new_n9680_), .A1(new_n9679_), .B0(new_n9683_), .Y(new_n9684_));
  AOI21X1  g08682(.A0(new_n7890_), .A1(new_n7884_), .B0(new_n7876_), .Y(new_n9685_));
  NOR2X1   g08683(.A(new_n9682_), .B(new_n9681_), .Y(new_n9686_));
  AOI21X1  g08684(.A0(new_n7889_), .A1(new_n7904_), .B0(new_n7888_), .Y(new_n9687_));
  OAI21X1  g08685(.A0(new_n7901_), .A1(new_n7870_), .B0(new_n7900_), .Y(new_n9688_));
  OAI22X1  g08686(.A0(new_n9688_), .A1(new_n9687_), .B0(new_n7914_), .B1(new_n7913_), .Y(new_n9689_));
  NOR3X1   g08687(.A(new_n9689_), .B(new_n9686_), .C(new_n9685_), .Y(new_n9690_));
  NOR2X1   g08688(.A(new_n9690_), .B(new_n9684_), .Y(new_n9691_));
  XOR2X1   g08689(.A(new_n9691_), .B(new_n9678_), .Y(new_n9692_));
  XOR2X1   g08690(.A(new_n9692_), .B(new_n9661_), .Y(new_n9693_));
  OR2X1    g08691(.A(new_n7848_), .B(new_n7814_), .Y(new_n9694_));
  OAI21X1  g08692(.A0(new_n7849_), .A1(new_n7843_), .B0(new_n7785_), .Y(new_n9695_));
  AND2X1   g08693(.A(new_n9695_), .B(new_n9694_), .Y(new_n9696_));
  OR2X1    g08694(.A(new_n7783_), .B(new_n7775_), .Y(new_n9697_));
  XOR2X1   g08695(.A(new_n7648_), .B(new_n7642_), .Y(new_n9698_));
  OR2X1    g08696(.A(new_n7648_), .B(new_n7642_), .Y(new_n9699_));
  OR2X1    g08697(.A(new_n7652_), .B(new_n7650_), .Y(new_n9700_));
  OAI21X1  g08698(.A0(new_n9699_), .A1(new_n7781_), .B0(new_n9700_), .Y(new_n9701_));
  AOI21X1  g08699(.A0(new_n9701_), .A1(new_n9698_), .B0(new_n7782_), .Y(new_n9702_));
  OAI21X1  g08700(.A0(new_n7773_), .A1(new_n7763_), .B0(new_n9702_), .Y(new_n9703_));
  OAI21X1  g08701(.A0(new_n7772_), .A1(new_n7756_), .B0(new_n7770_), .Y(new_n9704_));
  AOI21X1  g08702(.A0(new_n7754_), .A1(new_n9698_), .B0(new_n7753_), .Y(new_n9705_));
  XOR2X1   g08703(.A(new_n9705_), .B(new_n9704_), .Y(new_n9706_));
  AOI21X1  g08704(.A0(new_n9703_), .A1(new_n9697_), .B0(new_n9706_), .Y(new_n9707_));
  AND2X1   g08705(.A(new_n7857_), .B(new_n7856_), .Y(new_n9708_));
  AOI21X1  g08706(.A0(new_n7855_), .A1(new_n7852_), .B0(new_n7755_), .Y(new_n9709_));
  AND2X1   g08707(.A(new_n9705_), .B(new_n9704_), .Y(new_n9710_));
  NOR2X1   g08708(.A(new_n9705_), .B(new_n9704_), .Y(new_n9711_));
  NOR4X1   g08709(.A(new_n9711_), .B(new_n9710_), .C(new_n9709_), .D(new_n9708_), .Y(new_n9712_));
  OR2X1    g08710(.A(new_n9712_), .B(new_n9707_), .Y(new_n9713_));
  OR2X1    g08711(.A(new_n7835_), .B(new_n7834_), .Y(new_n9714_));
  OAI21X1  g08712(.A0(new_n7833_), .A1(new_n7824_), .B0(new_n7823_), .Y(new_n9715_));
  OAI21X1  g08713(.A0(new_n7832_), .A1(new_n7798_), .B0(new_n7831_), .Y(new_n9716_));
  AOI21X1  g08714(.A0(new_n7796_), .A1(new_n7815_), .B0(new_n7795_), .Y(new_n9717_));
  XOR2X1   g08715(.A(new_n9717_), .B(new_n9716_), .Y(new_n9718_));
  AOI21X1  g08716(.A0(new_n9715_), .A1(new_n9714_), .B0(new_n9718_), .Y(new_n9719_));
  AOI21X1  g08717(.A0(new_n7811_), .A1(new_n7805_), .B0(new_n7797_), .Y(new_n9720_));
  NOR2X1   g08718(.A(new_n9717_), .B(new_n9716_), .Y(new_n9721_));
  AOI21X1  g08719(.A0(new_n7810_), .A1(new_n7825_), .B0(new_n7809_), .Y(new_n9722_));
  OAI21X1  g08720(.A0(new_n7822_), .A1(new_n7791_), .B0(new_n7821_), .Y(new_n9723_));
  OAI22X1  g08721(.A0(new_n9723_), .A1(new_n9722_), .B0(new_n7835_), .B1(new_n7834_), .Y(new_n9724_));
  NOR3X1   g08722(.A(new_n9724_), .B(new_n9721_), .C(new_n9720_), .Y(new_n9725_));
  NOR2X1   g08723(.A(new_n9725_), .B(new_n9719_), .Y(new_n9726_));
  XOR2X1   g08724(.A(new_n9726_), .B(new_n9713_), .Y(new_n9727_));
  XOR2X1   g08725(.A(new_n9727_), .B(new_n9696_), .Y(new_n9728_));
  XOR2X1   g08726(.A(new_n9728_), .B(new_n9693_), .Y(new_n9729_));
  XOR2X1   g08727(.A(new_n9729_), .B(new_n9641_), .Y(new_n9730_));
  AND2X1   g08728(.A(new_n7735_), .B(new_n7554_), .Y(new_n9731_));
  AOI21X1  g08729(.A0(new_n7736_), .A1(new_n7732_), .B0(new_n7382_), .Y(new_n9732_));
  OR2X1    g08730(.A(new_n9732_), .B(new_n9731_), .Y(new_n9733_));
  OR2X1    g08731(.A(new_n8787_), .B(new_n7318_), .Y(new_n9734_));
  NOR4X1   g08732(.A(new_n7357_), .B(new_n7344_), .C(new_n7356_), .D(new_n7351_), .Y(new_n9735_));
  XOR2X1   g08733(.A(new_n7368_), .B(new_n9735_), .Y(new_n9736_));
  OR4X1    g08734(.A(new_n7344_), .B(new_n7356_), .C(new_n7367_), .D(new_n7351_), .Y(new_n9737_));
  AND2X1   g08735(.A(new_n7310_), .B(\A[324] ), .Y(new_n9738_));
  OR2X1    g08736(.A(new_n9738_), .B(new_n7312_), .Y(new_n9739_));
  XOR2X1   g08737(.A(new_n7315_), .B(new_n9739_), .Y(new_n9740_));
  XOR2X1   g08738(.A(new_n7346_), .B(new_n9740_), .Y(new_n9741_));
  OAI22X1  g08739(.A0(new_n9741_), .A1(new_n7348_), .B0(new_n7372_), .B1(new_n7351_), .Y(new_n9742_));
  OAI22X1  g08740(.A0(new_n9742_), .A1(new_n9737_), .B0(new_n7368_), .B1(new_n9735_), .Y(new_n9743_));
  MX2X1    g08741(.A(new_n9743_), .B(new_n9736_), .S0(new_n7350_), .Y(new_n9744_));
  OAI21X1  g08742(.A0(new_n8789_), .A1(new_n8781_), .B0(new_n9744_), .Y(new_n9745_));
  AND2X1   g08743(.A(new_n9745_), .B(new_n9734_), .Y(new_n9746_));
  OR2X1    g08744(.A(new_n9742_), .B(new_n9737_), .Y(new_n9747_));
  XOR2X1   g08745(.A(new_n7311_), .B(new_n7305_), .Y(new_n9748_));
  OR2X1    g08746(.A(new_n7311_), .B(new_n7305_), .Y(new_n9749_));
  OR2X1    g08747(.A(new_n7315_), .B(new_n7313_), .Y(new_n9750_));
  OAI21X1  g08748(.A0(new_n9749_), .A1(new_n9740_), .B0(new_n9750_), .Y(new_n9751_));
  AOI21X1  g08749(.A0(new_n9751_), .A1(new_n9748_), .B0(new_n9741_), .Y(new_n9752_));
  OAI21X1  g08750(.A0(new_n7368_), .A1(new_n9735_), .B0(new_n9752_), .Y(new_n9753_));
  OAI21X1  g08751(.A0(new_n7367_), .A1(new_n7351_), .B0(new_n7365_), .Y(new_n9754_));
  AOI21X1  g08752(.A0(new_n7349_), .A1(new_n9748_), .B0(new_n7348_), .Y(new_n9755_));
  XOR2X1   g08753(.A(new_n9755_), .B(new_n9754_), .Y(new_n9756_));
  AOI21X1  g08754(.A0(new_n9753_), .A1(new_n9747_), .B0(new_n9756_), .Y(new_n9757_));
  AOI21X1  g08755(.A0(new_n7374_), .A1(new_n7358_), .B0(new_n7350_), .Y(new_n9758_));
  NOR2X1   g08756(.A(new_n9755_), .B(new_n9754_), .Y(new_n9759_));
  AOI21X1  g08757(.A0(new_n7373_), .A1(new_n7359_), .B0(new_n7372_), .Y(new_n9760_));
  OAI21X1  g08758(.A0(new_n9741_), .A1(new_n7344_), .B0(new_n9751_), .Y(new_n9761_));
  OAI22X1  g08759(.A0(new_n9761_), .A1(new_n9760_), .B0(new_n9742_), .B1(new_n9737_), .Y(new_n9762_));
  NOR3X1   g08760(.A(new_n9762_), .B(new_n9759_), .C(new_n9758_), .Y(new_n9763_));
  NOR2X1   g08761(.A(new_n9763_), .B(new_n9757_), .Y(new_n9764_));
  OR2X1    g08762(.A(new_n7334_), .B(new_n7333_), .Y(new_n9765_));
  OAI21X1  g08763(.A0(new_n7332_), .A1(new_n7324_), .B0(new_n7323_), .Y(new_n9766_));
  OAI21X1  g08764(.A0(new_n7265_), .A1(new_n7331_), .B0(new_n7330_), .Y(new_n9767_));
  AOI21X1  g08765(.A0(new_n7320_), .A1(new_n7229_), .B0(new_n7240_), .Y(new_n9768_));
  XOR2X1   g08766(.A(new_n9768_), .B(new_n9767_), .Y(new_n9769_));
  AOI21X1  g08767(.A0(new_n9766_), .A1(new_n9765_), .B0(new_n9769_), .Y(new_n9770_));
  AOI21X1  g08768(.A0(new_n7272_), .A1(new_n7266_), .B0(new_n7241_), .Y(new_n9771_));
  NOR2X1   g08769(.A(new_n9768_), .B(new_n9767_), .Y(new_n9772_));
  AOI21X1  g08770(.A0(new_n7278_), .A1(new_n7271_), .B0(new_n7270_), .Y(new_n9773_));
  OAI21X1  g08771(.A0(new_n7235_), .A1(new_n7319_), .B0(new_n7322_), .Y(new_n9774_));
  OAI22X1  g08772(.A0(new_n9774_), .A1(new_n9773_), .B0(new_n7334_), .B1(new_n7333_), .Y(new_n9775_));
  NOR3X1   g08773(.A(new_n9775_), .B(new_n9772_), .C(new_n9771_), .Y(new_n9776_));
  NOR2X1   g08774(.A(new_n9776_), .B(new_n9770_), .Y(new_n9777_));
  XOR2X1   g08775(.A(new_n9777_), .B(new_n9764_), .Y(new_n9778_));
  XOR2X1   g08776(.A(new_n9778_), .B(new_n9746_), .Y(new_n9779_));
  OR2X1    g08777(.A(new_n7546_), .B(new_n7575_), .Y(new_n9780_));
  OAI21X1  g08778(.A0(new_n7733_), .A1(new_n7524_), .B0(new_n7574_), .Y(new_n9781_));
  AND2X1   g08779(.A(new_n9781_), .B(new_n9780_), .Y(new_n9782_));
  OR2X1    g08780(.A(new_n7572_), .B(new_n7571_), .Y(new_n9783_));
  XOR2X1   g08781(.A(new_n7401_), .B(new_n7409_), .Y(new_n9784_));
  XOR2X1   g08782(.A(new_n7394_), .B(new_n7388_), .Y(new_n9785_));
  OR2X1    g08783(.A(new_n7400_), .B(new_n7410_), .Y(new_n9786_));
  OAI21X1  g08784(.A0(new_n7401_), .A1(new_n7395_), .B0(new_n9786_), .Y(new_n9787_));
  AOI21X1  g08785(.A0(new_n9787_), .A1(new_n9785_), .B0(new_n9784_), .Y(new_n9788_));
  OAI21X1  g08786(.A0(new_n7449_), .A1(new_n7569_), .B0(new_n9788_), .Y(new_n9789_));
  OAI21X1  g08787(.A0(new_n7438_), .A1(new_n7447_), .B0(new_n7445_), .Y(new_n9790_));
  AOI21X1  g08788(.A0(new_n9785_), .A1(new_n7402_), .B0(new_n7413_), .Y(new_n9791_));
  XOR2X1   g08789(.A(new_n9791_), .B(new_n9790_), .Y(new_n9792_));
  AOI21X1  g08790(.A0(new_n9789_), .A1(new_n9783_), .B0(new_n9792_), .Y(new_n9793_));
  AND2X1   g08791(.A(new_n7457_), .B(new_n7456_), .Y(new_n9794_));
  AOI21X1  g08792(.A0(new_n7455_), .A1(new_n7439_), .B0(new_n7414_), .Y(new_n9795_));
  AND2X1   g08793(.A(new_n9791_), .B(new_n9790_), .Y(new_n9796_));
  NOR2X1   g08794(.A(new_n9791_), .B(new_n9790_), .Y(new_n9797_));
  NOR4X1   g08795(.A(new_n9797_), .B(new_n9796_), .C(new_n9795_), .D(new_n9794_), .Y(new_n9798_));
  OR2X1    g08796(.A(new_n9798_), .B(new_n9793_), .Y(new_n9799_));
  OR2X1    g08797(.A(new_n7558_), .B(new_n7557_), .Y(new_n9800_));
  OAI21X1  g08798(.A0(new_n7544_), .A1(new_n7556_), .B0(new_n7565_), .Y(new_n9801_));
  OAI21X1  g08799(.A0(new_n7515_), .A1(new_n7535_), .B0(new_n7539_), .Y(new_n9802_));
  AOI21X1  g08800(.A0(new_n7562_), .A1(new_n7479_), .B0(new_n7490_), .Y(new_n9803_));
  XOR2X1   g08801(.A(new_n9803_), .B(new_n9802_), .Y(new_n9804_));
  AOI21X1  g08802(.A0(new_n9801_), .A1(new_n9800_), .B0(new_n9804_), .Y(new_n9805_));
  AOI21X1  g08803(.A0(new_n7522_), .A1(new_n7516_), .B0(new_n7491_), .Y(new_n9806_));
  NOR2X1   g08804(.A(new_n9803_), .B(new_n9802_), .Y(new_n9807_));
  AOI21X1  g08805(.A0(new_n7540_), .A1(new_n7521_), .B0(new_n7520_), .Y(new_n9808_));
  OAI21X1  g08806(.A0(new_n7485_), .A1(new_n7561_), .B0(new_n7564_), .Y(new_n9809_));
  OAI22X1  g08807(.A0(new_n9809_), .A1(new_n9808_), .B0(new_n7558_), .B1(new_n7557_), .Y(new_n9810_));
  NOR3X1   g08808(.A(new_n9810_), .B(new_n9807_), .C(new_n9806_), .Y(new_n9811_));
  NOR2X1   g08809(.A(new_n9811_), .B(new_n9805_), .Y(new_n9812_));
  XOR2X1   g08810(.A(new_n9812_), .B(new_n9799_), .Y(new_n9813_));
  XOR2X1   g08811(.A(new_n9813_), .B(new_n9782_), .Y(new_n9814_));
  XOR2X1   g08812(.A(new_n9814_), .B(new_n9779_), .Y(new_n9815_));
  XOR2X1   g08813(.A(new_n9815_), .B(new_n9733_), .Y(new_n9816_));
  XOR2X1   g08814(.A(new_n9816_), .B(new_n9730_), .Y(new_n9817_));
  XOR2X1   g08815(.A(new_n9817_), .B(new_n9638_), .Y(new_n9818_));
  AND2X1   g08816(.A(new_n8763_), .B(new_n8709_), .Y(new_n9819_));
  AOI21X1  g08817(.A0(new_n8765_), .A1(new_n8759_), .B0(new_n8333_), .Y(new_n9820_));
  OR2X1    g08818(.A(new_n9820_), .B(new_n9819_), .Y(new_n9821_));
  AND2X1   g08819(.A(new_n8230_), .B(new_n8330_), .Y(new_n9822_));
  AOI21X1  g08820(.A0(new_n8331_), .A1(new_n8139_), .B0(new_n8329_), .Y(new_n9823_));
  OR2X1    g08821(.A(new_n9823_), .B(new_n9822_), .Y(new_n9824_));
  XOR2X1   g08822(.A(new_n8279_), .B(new_n8251_), .Y(new_n9825_));
  NOR4X1   g08823(.A(new_n8237_), .B(new_n8278_), .C(new_n8277_), .D(new_n8244_), .Y(new_n9826_));
  AOI21X1  g08824(.A0(new_n8277_), .A1(new_n8271_), .B0(new_n8250_), .Y(new_n9827_));
  AOI22X1  g08825(.A0(new_n9827_), .A1(new_n9826_), .B0(new_n8257_), .B1(new_n8251_), .Y(new_n9828_));
  MX2X1    g08826(.A(new_n9828_), .B(new_n9825_), .S0(new_n8243_), .Y(new_n9829_));
  OR2X1    g08827(.A(new_n9829_), .B(new_n8260_), .Y(new_n9830_));
  AND2X1   g08828(.A(new_n8258_), .B(new_n8243_), .Y(new_n9831_));
  NOR4X1   g08829(.A(new_n8304_), .B(new_n8291_), .C(new_n8303_), .D(new_n8298_), .Y(new_n9832_));
  XOR2X1   g08830(.A(new_n8315_), .B(new_n9832_), .Y(new_n9833_));
  OR4X1    g08831(.A(new_n8291_), .B(new_n8303_), .C(new_n8314_), .D(new_n8298_), .Y(new_n9834_));
  AND2X1   g08832(.A(new_n8208_), .B(\A[372] ), .Y(new_n9835_));
  OR2X1    g08833(.A(new_n9835_), .B(new_n8210_), .Y(new_n9836_));
  XOR2X1   g08834(.A(new_n8213_), .B(new_n9836_), .Y(new_n9837_));
  XOR2X1   g08835(.A(new_n8293_), .B(new_n9837_), .Y(new_n9838_));
  OAI22X1  g08836(.A0(new_n9838_), .A1(new_n8295_), .B0(new_n8319_), .B1(new_n8298_), .Y(new_n9839_));
  OAI22X1  g08837(.A0(new_n9839_), .A1(new_n9834_), .B0(new_n8315_), .B1(new_n9832_), .Y(new_n9840_));
  MX2X1    g08838(.A(new_n9840_), .B(new_n9833_), .S0(new_n8297_), .Y(new_n9841_));
  OAI21X1  g08839(.A0(new_n9828_), .A1(new_n8243_), .B0(new_n8260_), .Y(new_n9842_));
  OAI21X1  g08840(.A0(new_n9842_), .A1(new_n9831_), .B0(new_n9841_), .Y(new_n9843_));
  AND2X1   g08841(.A(new_n9843_), .B(new_n9830_), .Y(new_n9844_));
  OR2X1    g08842(.A(new_n9839_), .B(new_n9834_), .Y(new_n9845_));
  XOR2X1   g08843(.A(new_n8209_), .B(new_n8203_), .Y(new_n9846_));
  OR2X1    g08844(.A(new_n8209_), .B(new_n8203_), .Y(new_n9847_));
  OR2X1    g08845(.A(new_n8213_), .B(new_n8211_), .Y(new_n9848_));
  OAI21X1  g08846(.A0(new_n9847_), .A1(new_n9837_), .B0(new_n9848_), .Y(new_n9849_));
  AOI21X1  g08847(.A0(new_n9849_), .A1(new_n9846_), .B0(new_n9838_), .Y(new_n9850_));
  OAI21X1  g08848(.A0(new_n8315_), .A1(new_n9832_), .B0(new_n9850_), .Y(new_n9851_));
  OAI21X1  g08849(.A0(new_n8314_), .A1(new_n8298_), .B0(new_n8312_), .Y(new_n9852_));
  AOI21X1  g08850(.A0(new_n8296_), .A1(new_n9846_), .B0(new_n8295_), .Y(new_n9853_));
  XOR2X1   g08851(.A(new_n9853_), .B(new_n9852_), .Y(new_n9854_));
  AOI21X1  g08852(.A0(new_n9851_), .A1(new_n9845_), .B0(new_n9854_), .Y(new_n9855_));
  AND2X1   g08853(.A(new_n8323_), .B(new_n8322_), .Y(new_n9856_));
  AOI21X1  g08854(.A0(new_n8321_), .A1(new_n8305_), .B0(new_n8297_), .Y(new_n9857_));
  AND2X1   g08855(.A(new_n9853_), .B(new_n9852_), .Y(new_n9858_));
  NOR2X1   g08856(.A(new_n9853_), .B(new_n9852_), .Y(new_n9859_));
  NOR4X1   g08857(.A(new_n9859_), .B(new_n9858_), .C(new_n9857_), .D(new_n9856_), .Y(new_n9860_));
  NOR2X1   g08858(.A(new_n9860_), .B(new_n9855_), .Y(new_n9861_));
  OR2X1    g08859(.A(new_n8281_), .B(new_n8280_), .Y(new_n9862_));
  OAI21X1  g08860(.A0(new_n8279_), .A1(new_n8270_), .B0(new_n8269_), .Y(new_n9863_));
  OAI21X1  g08861(.A0(new_n8278_), .A1(new_n8244_), .B0(new_n8277_), .Y(new_n9864_));
  AOI21X1  g08862(.A0(new_n8242_), .A1(new_n8261_), .B0(new_n8241_), .Y(new_n9865_));
  XOR2X1   g08863(.A(new_n9865_), .B(new_n9864_), .Y(new_n9866_));
  AOI21X1  g08864(.A0(new_n9863_), .A1(new_n9862_), .B0(new_n9866_), .Y(new_n9867_));
  AOI21X1  g08865(.A0(new_n8257_), .A1(new_n8251_), .B0(new_n8243_), .Y(new_n9868_));
  NOR2X1   g08866(.A(new_n9865_), .B(new_n9864_), .Y(new_n9869_));
  AOI21X1  g08867(.A0(new_n8256_), .A1(new_n8271_), .B0(new_n8255_), .Y(new_n9870_));
  OAI21X1  g08868(.A0(new_n8268_), .A1(new_n8237_), .B0(new_n8267_), .Y(new_n9871_));
  OAI22X1  g08869(.A0(new_n9871_), .A1(new_n9870_), .B0(new_n8281_), .B1(new_n8280_), .Y(new_n9872_));
  NOR3X1   g08870(.A(new_n9872_), .B(new_n9869_), .C(new_n9868_), .Y(new_n9873_));
  NOR2X1   g08871(.A(new_n9873_), .B(new_n9867_), .Y(new_n9874_));
  XOR2X1   g08872(.A(new_n9874_), .B(new_n9861_), .Y(new_n9875_));
  XOR2X1   g08873(.A(new_n9875_), .B(new_n9844_), .Y(new_n9876_));
  OR2X1    g08874(.A(new_n8223_), .B(new_n8117_), .Y(new_n9877_));
  OAI21X1  g08875(.A0(new_n8224_), .A1(new_n8218_), .B0(new_n8045_), .Y(new_n9878_));
  AND2X1   g08876(.A(new_n9878_), .B(new_n9877_), .Y(new_n9879_));
  OR2X1    g08877(.A(new_n8043_), .B(new_n8039_), .Y(new_n9880_));
  XOR2X1   g08878(.A(new_n7989_), .B(new_n7997_), .Y(new_n9881_));
  XOR2X1   g08879(.A(new_n7982_), .B(new_n7976_), .Y(new_n9882_));
  OR2X1    g08880(.A(new_n7988_), .B(new_n7998_), .Y(new_n9883_));
  OAI21X1  g08881(.A0(new_n7989_), .A1(new_n7983_), .B0(new_n9883_), .Y(new_n9884_));
  AOI21X1  g08882(.A0(new_n9884_), .A1(new_n9882_), .B0(new_n9881_), .Y(new_n9885_));
  OAI21X1  g08883(.A0(new_n8037_), .A1(new_n8027_), .B0(new_n9885_), .Y(new_n9886_));
  OAI21X1  g08884(.A0(new_n8026_), .A1(new_n8035_), .B0(new_n8033_), .Y(new_n9887_));
  AOI21X1  g08885(.A0(new_n9882_), .A1(new_n7990_), .B0(new_n8001_), .Y(new_n9888_));
  XOR2X1   g08886(.A(new_n9888_), .B(new_n9887_), .Y(new_n9889_));
  AOI21X1  g08887(.A0(new_n9886_), .A1(new_n9880_), .B0(new_n9889_), .Y(new_n9890_));
  AND2X1   g08888(.A(new_n8728_), .B(new_n8727_), .Y(new_n9891_));
  AOI21X1  g08889(.A0(new_n8726_), .A1(new_n8723_), .B0(new_n8002_), .Y(new_n9892_));
  AND2X1   g08890(.A(new_n9888_), .B(new_n9887_), .Y(new_n9893_));
  NOR2X1   g08891(.A(new_n9888_), .B(new_n9887_), .Y(new_n9894_));
  NOR4X1   g08892(.A(new_n9894_), .B(new_n9893_), .C(new_n9892_), .D(new_n9891_), .Y(new_n9895_));
  OR2X1    g08893(.A(new_n9895_), .B(new_n9890_), .Y(new_n9896_));
  OR2X1    g08894(.A(new_n8134_), .B(new_n8133_), .Y(new_n9897_));
  OAI21X1  g08895(.A0(new_n8132_), .A1(new_n8123_), .B0(new_n8122_), .Y(new_n9898_));
  OAI21X1  g08896(.A0(new_n8101_), .A1(new_n8130_), .B0(new_n8129_), .Y(new_n9899_));
  AOI21X1  g08897(.A0(new_n8119_), .A1(new_n8065_), .B0(new_n8076_), .Y(new_n9900_));
  XOR2X1   g08898(.A(new_n9900_), .B(new_n9899_), .Y(new_n9901_));
  AOI21X1  g08899(.A0(new_n9898_), .A1(new_n9897_), .B0(new_n9901_), .Y(new_n9902_));
  AOI21X1  g08900(.A0(new_n8108_), .A1(new_n8102_), .B0(new_n8077_), .Y(new_n9903_));
  NOR2X1   g08901(.A(new_n9900_), .B(new_n9899_), .Y(new_n9904_));
  AOI21X1  g08902(.A0(new_n8131_), .A1(new_n8107_), .B0(new_n8106_), .Y(new_n9905_));
  OAI21X1  g08903(.A0(new_n8071_), .A1(new_n8118_), .B0(new_n8121_), .Y(new_n9906_));
  OAI22X1  g08904(.A0(new_n9906_), .A1(new_n9905_), .B0(new_n8134_), .B1(new_n8133_), .Y(new_n9907_));
  NOR3X1   g08905(.A(new_n9907_), .B(new_n9904_), .C(new_n9903_), .Y(new_n9908_));
  NOR2X1   g08906(.A(new_n9908_), .B(new_n9902_), .Y(new_n9909_));
  XOR2X1   g08907(.A(new_n9909_), .B(new_n9896_), .Y(new_n9910_));
  XOR2X1   g08908(.A(new_n9910_), .B(new_n9879_), .Y(new_n9911_));
  XOR2X1   g08909(.A(new_n9911_), .B(new_n9876_), .Y(new_n9912_));
  XOR2X1   g08910(.A(new_n9912_), .B(new_n9824_), .Y(new_n9913_));
  OR2X1    g08911(.A(new_n8702_), .B(new_n8717_), .Y(new_n9914_));
  OAI21X1  g08912(.A0(new_n8760_), .A1(new_n8672_), .B0(new_n8758_), .Y(new_n9915_));
  AND2X1   g08913(.A(new_n9915_), .B(new_n9914_), .Y(new_n9916_));
  OR2X1    g08914(.A(new_n8754_), .B(new_n8442_), .Y(new_n9917_));
  NOR4X1   g08915(.A(new_n8481_), .B(new_n8468_), .C(new_n8480_), .D(new_n8475_), .Y(new_n9918_));
  XOR2X1   g08916(.A(new_n8492_), .B(new_n9918_), .Y(new_n9919_));
  OR4X1    g08917(.A(new_n8468_), .B(new_n8480_), .C(new_n8491_), .D(new_n8475_), .Y(new_n9920_));
  AND2X1   g08918(.A(new_n8434_), .B(\A[420] ), .Y(new_n9921_));
  OR2X1    g08919(.A(new_n9921_), .B(new_n8436_), .Y(new_n9922_));
  XOR2X1   g08920(.A(new_n8439_), .B(new_n9922_), .Y(new_n9923_));
  XOR2X1   g08921(.A(new_n8470_), .B(new_n9923_), .Y(new_n9924_));
  OAI22X1  g08922(.A0(new_n9924_), .A1(new_n8472_), .B0(new_n8496_), .B1(new_n8475_), .Y(new_n9925_));
  OAI22X1  g08923(.A0(new_n9925_), .A1(new_n9920_), .B0(new_n8492_), .B1(new_n9918_), .Y(new_n9926_));
  MX2X1    g08924(.A(new_n9926_), .B(new_n9919_), .S0(new_n8474_), .Y(new_n9927_));
  OAI21X1  g08925(.A0(new_n8756_), .A1(new_n8748_), .B0(new_n9927_), .Y(new_n9928_));
  AND2X1   g08926(.A(new_n9928_), .B(new_n9917_), .Y(new_n9929_));
  OR2X1    g08927(.A(new_n9925_), .B(new_n9920_), .Y(new_n9930_));
  XOR2X1   g08928(.A(new_n8435_), .B(new_n8429_), .Y(new_n9931_));
  OR2X1    g08929(.A(new_n8435_), .B(new_n8429_), .Y(new_n9932_));
  OR2X1    g08930(.A(new_n8439_), .B(new_n8437_), .Y(new_n9933_));
  OAI21X1  g08931(.A0(new_n9932_), .A1(new_n9923_), .B0(new_n9933_), .Y(new_n9934_));
  AOI21X1  g08932(.A0(new_n9934_), .A1(new_n9931_), .B0(new_n9924_), .Y(new_n9935_));
  OAI21X1  g08933(.A0(new_n8492_), .A1(new_n9918_), .B0(new_n9935_), .Y(new_n9936_));
  OAI21X1  g08934(.A0(new_n8491_), .A1(new_n8475_), .B0(new_n8489_), .Y(new_n9937_));
  AOI21X1  g08935(.A0(new_n8473_), .A1(new_n9931_), .B0(new_n8472_), .Y(new_n9938_));
  XOR2X1   g08936(.A(new_n9938_), .B(new_n9937_), .Y(new_n9939_));
  AOI21X1  g08937(.A0(new_n9936_), .A1(new_n9930_), .B0(new_n9939_), .Y(new_n9940_));
  AOI21X1  g08938(.A0(new_n8498_), .A1(new_n8482_), .B0(new_n8474_), .Y(new_n9941_));
  NOR2X1   g08939(.A(new_n9938_), .B(new_n9937_), .Y(new_n9942_));
  AOI21X1  g08940(.A0(new_n8497_), .A1(new_n8483_), .B0(new_n8496_), .Y(new_n9943_));
  OAI21X1  g08941(.A0(new_n9924_), .A1(new_n8468_), .B0(new_n9934_), .Y(new_n9944_));
  OAI22X1  g08942(.A0(new_n9944_), .A1(new_n9943_), .B0(new_n9925_), .B1(new_n9920_), .Y(new_n9945_));
  NOR3X1   g08943(.A(new_n9945_), .B(new_n9942_), .C(new_n9941_), .Y(new_n9946_));
  NOR2X1   g08944(.A(new_n9946_), .B(new_n9940_), .Y(new_n9947_));
  OR2X1    g08945(.A(new_n8458_), .B(new_n8457_), .Y(new_n9948_));
  OAI21X1  g08946(.A0(new_n8456_), .A1(new_n8448_), .B0(new_n8447_), .Y(new_n9949_));
  OAI21X1  g08947(.A0(new_n8389_), .A1(new_n8455_), .B0(new_n8454_), .Y(new_n9950_));
  AOI21X1  g08948(.A0(new_n8444_), .A1(new_n8353_), .B0(new_n8364_), .Y(new_n9951_));
  XOR2X1   g08949(.A(new_n9951_), .B(new_n9950_), .Y(new_n9952_));
  AOI21X1  g08950(.A0(new_n9949_), .A1(new_n9948_), .B0(new_n9952_), .Y(new_n9953_));
  AOI21X1  g08951(.A0(new_n8396_), .A1(new_n8390_), .B0(new_n8365_), .Y(new_n9954_));
  NOR2X1   g08952(.A(new_n9951_), .B(new_n9950_), .Y(new_n9955_));
  AOI21X1  g08953(.A0(new_n8402_), .A1(new_n8395_), .B0(new_n8394_), .Y(new_n9956_));
  OAI21X1  g08954(.A0(new_n8359_), .A1(new_n8443_), .B0(new_n8446_), .Y(new_n9957_));
  OAI22X1  g08955(.A0(new_n9957_), .A1(new_n9956_), .B0(new_n8458_), .B1(new_n8457_), .Y(new_n9958_));
  NOR3X1   g08956(.A(new_n9958_), .B(new_n9955_), .C(new_n9954_), .Y(new_n9959_));
  NOR2X1   g08957(.A(new_n9959_), .B(new_n9953_), .Y(new_n9960_));
  XOR2X1   g08958(.A(new_n9960_), .B(new_n9947_), .Y(new_n9961_));
  XOR2X1   g08959(.A(new_n9961_), .B(new_n9929_), .Y(new_n9962_));
  OR2X1    g08960(.A(new_n8670_), .B(new_n8699_), .Y(new_n9963_));
  OAI21X1  g08961(.A0(new_n8711_), .A1(new_n8648_), .B0(new_n8698_), .Y(new_n9964_));
  AND2X1   g08962(.A(new_n9964_), .B(new_n9963_), .Y(new_n9965_));
  OR2X1    g08963(.A(new_n8696_), .B(new_n8695_), .Y(new_n9966_));
  XOR2X1   g08964(.A(new_n8525_), .B(new_n8533_), .Y(new_n9967_));
  XOR2X1   g08965(.A(new_n8518_), .B(new_n8512_), .Y(new_n9968_));
  OR2X1    g08966(.A(new_n8524_), .B(new_n8534_), .Y(new_n9969_));
  OAI21X1  g08967(.A0(new_n8525_), .A1(new_n8519_), .B0(new_n9969_), .Y(new_n9970_));
  AOI21X1  g08968(.A0(new_n9970_), .A1(new_n9968_), .B0(new_n9967_), .Y(new_n9971_));
  OAI21X1  g08969(.A0(new_n8573_), .A1(new_n8693_), .B0(new_n9971_), .Y(new_n9972_));
  OAI21X1  g08970(.A0(new_n8562_), .A1(new_n8571_), .B0(new_n8569_), .Y(new_n9973_));
  AOI21X1  g08971(.A0(new_n9968_), .A1(new_n8526_), .B0(new_n8537_), .Y(new_n9974_));
  XOR2X1   g08972(.A(new_n9974_), .B(new_n9973_), .Y(new_n9975_));
  AOI21X1  g08973(.A0(new_n9972_), .A1(new_n9966_), .B0(new_n9975_), .Y(new_n9976_));
  AND2X1   g08974(.A(new_n8581_), .B(new_n8580_), .Y(new_n9977_));
  AOI21X1  g08975(.A0(new_n8579_), .A1(new_n8563_), .B0(new_n8538_), .Y(new_n9978_));
  AND2X1   g08976(.A(new_n9974_), .B(new_n9973_), .Y(new_n9979_));
  NOR2X1   g08977(.A(new_n9974_), .B(new_n9973_), .Y(new_n9980_));
  NOR4X1   g08978(.A(new_n9980_), .B(new_n9979_), .C(new_n9978_), .D(new_n9977_), .Y(new_n9981_));
  OR2X1    g08979(.A(new_n9981_), .B(new_n9976_), .Y(new_n9982_));
  OR2X1    g08980(.A(new_n8682_), .B(new_n8681_), .Y(new_n9983_));
  OAI21X1  g08981(.A0(new_n8668_), .A1(new_n8680_), .B0(new_n8689_), .Y(new_n9984_));
  OAI21X1  g08982(.A0(new_n8639_), .A1(new_n8659_), .B0(new_n8663_), .Y(new_n9985_));
  AOI21X1  g08983(.A0(new_n8686_), .A1(new_n8603_), .B0(new_n8614_), .Y(new_n9986_));
  XOR2X1   g08984(.A(new_n9986_), .B(new_n9985_), .Y(new_n9987_));
  AOI21X1  g08985(.A0(new_n9984_), .A1(new_n9983_), .B0(new_n9987_), .Y(new_n9988_));
  AOI21X1  g08986(.A0(new_n8646_), .A1(new_n8640_), .B0(new_n8615_), .Y(new_n9989_));
  NOR2X1   g08987(.A(new_n9986_), .B(new_n9985_), .Y(new_n9990_));
  AOI21X1  g08988(.A0(new_n8664_), .A1(new_n8645_), .B0(new_n8644_), .Y(new_n9991_));
  OAI21X1  g08989(.A0(new_n8609_), .A1(new_n8685_), .B0(new_n8688_), .Y(new_n9992_));
  OAI22X1  g08990(.A0(new_n9992_), .A1(new_n9991_), .B0(new_n8682_), .B1(new_n8681_), .Y(new_n9993_));
  NOR3X1   g08991(.A(new_n9993_), .B(new_n9990_), .C(new_n9989_), .Y(new_n9994_));
  NOR2X1   g08992(.A(new_n9994_), .B(new_n9988_), .Y(new_n9995_));
  XOR2X1   g08993(.A(new_n9995_), .B(new_n9982_), .Y(new_n9996_));
  XOR2X1   g08994(.A(new_n9996_), .B(new_n9965_), .Y(new_n9997_));
  XOR2X1   g08995(.A(new_n9997_), .B(new_n9962_), .Y(new_n9998_));
  XOR2X1   g08996(.A(new_n9998_), .B(new_n9916_), .Y(new_n9999_));
  XOR2X1   g08997(.A(new_n9999_), .B(new_n9913_), .Y(new_n10000_));
  XOR2X1   g08998(.A(new_n10000_), .B(new_n9821_), .Y(new_n10001_));
  XOR2X1   g08999(.A(new_n10001_), .B(new_n9818_), .Y(new_n10002_));
  XOR2X1   g09000(.A(new_n10002_), .B(new_n9626_), .Y(new_n10003_));
  XOR2X1   g09001(.A(new_n10003_), .B(new_n9623_), .Y(new_n10004_));
  XOR2X1   g09002(.A(new_n10004_), .B(new_n9235_), .Y(new_n10005_));
  XOR2X1   g09003(.A(new_n10005_), .B(new_n9233_), .Y(new_n10006_));
  XOR2X1   g09004(.A(new_n10006_), .B(new_n8852_), .Y(new_n10007_));
  NOR3X1   g09005(.A(new_n3844_), .B(new_n2423_), .C(new_n2411_), .Y(new_n10008_));
  OR2X1    g09006(.A(new_n10008_), .B(new_n3842_), .Y(new_n10009_));
  AND2X1   g09007(.A(new_n10009_), .B(new_n3846_), .Y(new_n10010_));
  OR2X1    g09008(.A(new_n3829_), .B(new_n3823_), .Y(new_n10011_));
  NOR3X1   g09009(.A(new_n3733_), .B(new_n3740_), .C(new_n3737_), .Y(new_n10012_));
  AOI21X1  g09010(.A0(new_n3731_), .A1(new_n3727_), .B0(new_n3741_), .Y(new_n10013_));
  OAI21X1  g09011(.A0(new_n10013_), .A1(new_n10012_), .B0(new_n10011_), .Y(new_n10014_));
  OAI21X1  g09012(.A0(new_n10011_), .A1(new_n3743_), .B0(new_n10014_), .Y(new_n10015_));
  NOR3X1   g09013(.A(new_n3637_), .B(new_n3644_), .C(new_n3641_), .Y(new_n10016_));
  AOI21X1  g09014(.A0(new_n3636_), .A1(new_n3632_), .B0(new_n3645_), .Y(new_n10017_));
  OAI21X1  g09015(.A0(new_n10017_), .A1(new_n10016_), .B0(new_n10015_), .Y(new_n10018_));
  OAI21X1  g09016(.A0(new_n10015_), .A1(new_n3647_), .B0(new_n10018_), .Y(new_n10019_));
  AOI21X1  g09017(.A0(new_n3438_), .A1(new_n3430_), .B0(new_n3448_), .Y(new_n10020_));
  AOI21X1  g09018(.A0(new_n3839_), .A1(new_n10019_), .B0(new_n10020_), .Y(new_n10021_));
  AOI21X1  g09019(.A0(new_n3835_), .A1(new_n10015_), .B0(new_n10017_), .Y(new_n10022_));
  OAI21X1  g09020(.A0(new_n10012_), .A1(new_n3830_), .B0(new_n3832_), .Y(new_n10023_));
  AOI21X1  g09021(.A0(new_n3778_), .A1(new_n3765_), .B0(new_n3786_), .Y(new_n10024_));
  AOI21X1  g09022(.A0(new_n3827_), .A1(new_n3822_), .B0(new_n10024_), .Y(new_n10025_));
  OR2X1    g09023(.A(new_n3820_), .B(new_n3819_), .Y(new_n10026_));
  OAI21X1  g09024(.A0(new_n3818_), .A1(new_n3814_), .B0(new_n3824_), .Y(new_n10027_));
  AND2X1   g09025(.A(new_n3808_), .B(new_n3807_), .Y(new_n10028_));
  OAI22X1  g09026(.A0(new_n3816_), .A1(new_n3800_), .B0(new_n3809_), .B1(new_n10028_), .Y(new_n10029_));
  OR2X1    g09027(.A(new_n3791_), .B(new_n3788_), .Y(new_n10030_));
  AOI22X1  g09028(.A0(new_n3794_), .A1(new_n10030_), .B0(new_n3792_), .B1(new_n3793_), .Y(new_n10031_));
  XOR2X1   g09029(.A(new_n10031_), .B(new_n10029_), .Y(new_n10032_));
  AOI21X1  g09030(.A0(new_n10027_), .A1(new_n10026_), .B0(new_n10032_), .Y(new_n10033_));
  NOR3X1   g09031(.A(new_n3819_), .B(new_n3817_), .C(new_n3805_), .Y(new_n10034_));
  AND2X1   g09032(.A(new_n10031_), .B(new_n10029_), .Y(new_n10035_));
  NOR2X1   g09033(.A(new_n10031_), .B(new_n10029_), .Y(new_n10036_));
  NOR3X1   g09034(.A(new_n10036_), .B(new_n10035_), .C(new_n10034_), .Y(new_n10037_));
  AND2X1   g09035(.A(new_n10037_), .B(new_n10027_), .Y(new_n10038_));
  NOR2X1   g09036(.A(new_n10038_), .B(new_n10033_), .Y(new_n10039_));
  AOI21X1  g09037(.A0(new_n3763_), .A1(new_n3757_), .B0(new_n3752_), .Y(new_n10040_));
  OR2X1    g09038(.A(new_n10040_), .B(new_n3777_), .Y(new_n10041_));
  XOR2X1   g09039(.A(new_n2474_), .B(new_n3754_), .Y(new_n10042_));
  AOI21X1  g09040(.A0(new_n3762_), .A1(new_n10042_), .B0(new_n3761_), .Y(new_n10043_));
  AOI21X1  g09041(.A0(new_n3751_), .A1(new_n3766_), .B0(new_n3750_), .Y(new_n10044_));
  XOR2X1   g09042(.A(new_n10044_), .B(new_n10043_), .Y(new_n10045_));
  AND2X1   g09043(.A(new_n3759_), .B(new_n3758_), .Y(new_n10046_));
  OAI22X1  g09044(.A0(new_n3774_), .A1(new_n3753_), .B0(new_n3760_), .B1(new_n10046_), .Y(new_n10047_));
  AND2X1   g09045(.A(new_n10044_), .B(new_n10047_), .Y(new_n10048_));
  NOR2X1   g09046(.A(new_n10044_), .B(new_n10047_), .Y(new_n10049_));
  NOR4X1   g09047(.A(new_n10049_), .B(new_n10048_), .C(new_n10040_), .D(new_n3777_), .Y(new_n10050_));
  AOI21X1  g09048(.A0(new_n10045_), .A1(new_n10041_), .B0(new_n10050_), .Y(new_n10051_));
  XOR2X1   g09049(.A(new_n10051_), .B(new_n10039_), .Y(new_n10052_));
  XOR2X1   g09050(.A(new_n10052_), .B(new_n10025_), .Y(new_n10053_));
  OAI21X1  g09051(.A0(new_n3729_), .A1(new_n3679_), .B0(new_n3739_), .Y(new_n10054_));
  AOI21X1  g09052(.A0(new_n3668_), .A1(new_n3662_), .B0(new_n3656_), .Y(new_n10055_));
  OR2X1    g09053(.A(new_n10055_), .B(new_n3677_), .Y(new_n10056_));
  XOR2X1   g09054(.A(new_n2551_), .B(new_n3659_), .Y(new_n10057_));
  AOI21X1  g09055(.A0(new_n3667_), .A1(new_n10057_), .B0(new_n3666_), .Y(new_n10058_));
  XOR2X1   g09056(.A(new_n2569_), .B(new_n2563_), .Y(new_n10059_));
  AOI21X1  g09057(.A0(new_n3655_), .A1(new_n10059_), .B0(new_n3654_), .Y(new_n10060_));
  XOR2X1   g09058(.A(new_n10060_), .B(new_n10058_), .Y(new_n10061_));
  AND2X1   g09059(.A(new_n3664_), .B(new_n3663_), .Y(new_n10062_));
  OAI22X1  g09060(.A0(new_n3673_), .A1(new_n3658_), .B0(new_n3665_), .B1(new_n10062_), .Y(new_n10063_));
  AND2X1   g09061(.A(new_n10060_), .B(new_n10063_), .Y(new_n10064_));
  NOR2X1   g09062(.A(new_n10060_), .B(new_n10063_), .Y(new_n10065_));
  NOR4X1   g09063(.A(new_n10065_), .B(new_n10064_), .C(new_n10055_), .D(new_n3677_), .Y(new_n10066_));
  AOI21X1  g09064(.A0(new_n10061_), .A1(new_n10056_), .B0(new_n10066_), .Y(new_n10067_));
  AOI21X1  g09065(.A0(new_n3700_), .A1(new_n3694_), .B0(new_n3688_), .Y(new_n10068_));
  OR2X1    g09066(.A(new_n10068_), .B(new_n3723_), .Y(new_n10069_));
  XOR2X1   g09067(.A(new_n2512_), .B(new_n2506_), .Y(new_n10070_));
  AOI21X1  g09068(.A0(new_n3699_), .A1(new_n10070_), .B0(new_n3698_), .Y(new_n10071_));
  AOI21X1  g09069(.A0(new_n3687_), .A1(new_n3717_), .B0(new_n3686_), .Y(new_n10072_));
  XOR2X1   g09070(.A(new_n10072_), .B(new_n10071_), .Y(new_n10073_));
  AND2X1   g09071(.A(new_n3696_), .B(new_n3695_), .Y(new_n10074_));
  OAI22X1  g09072(.A0(new_n3705_), .A1(new_n3691_), .B0(new_n3697_), .B1(new_n10074_), .Y(new_n10075_));
  AND2X1   g09073(.A(new_n10072_), .B(new_n10075_), .Y(new_n10076_));
  NOR2X1   g09074(.A(new_n10072_), .B(new_n10075_), .Y(new_n10077_));
  NOR4X1   g09075(.A(new_n10077_), .B(new_n10076_), .C(new_n10068_), .D(new_n3723_), .Y(new_n10078_));
  AOI21X1  g09076(.A0(new_n10073_), .A1(new_n10069_), .B0(new_n10078_), .Y(new_n10079_));
  XOR2X1   g09077(.A(new_n10079_), .B(new_n10067_), .Y(new_n10080_));
  XOR2X1   g09078(.A(new_n10080_), .B(new_n10054_), .Y(new_n10081_));
  XOR2X1   g09079(.A(new_n10081_), .B(new_n10053_), .Y(new_n10082_));
  XOR2X1   g09080(.A(new_n10082_), .B(new_n10023_), .Y(new_n10083_));
  OAI21X1  g09081(.A0(new_n3634_), .A1(new_n3535_), .B0(new_n3643_), .Y(new_n10084_));
  AOI21X1  g09082(.A0(new_n3489_), .A1(new_n3473_), .B0(new_n3496_), .Y(new_n10085_));
  AOI21X1  g09083(.A0(new_n3532_), .A1(new_n3527_), .B0(new_n10085_), .Y(new_n10086_));
  AOI21X1  g09084(.A0(new_n3517_), .A1(new_n3511_), .B0(new_n3506_), .Y(new_n10087_));
  OR2X1    g09085(.A(new_n10087_), .B(new_n3525_), .Y(new_n10088_));
  XOR2X1   g09086(.A(new_n2705_), .B(new_n3508_), .Y(new_n10089_));
  AOI21X1  g09087(.A0(new_n3516_), .A1(new_n10089_), .B0(new_n3515_), .Y(new_n10090_));
  XOR2X1   g09088(.A(new_n2723_), .B(new_n2717_), .Y(new_n10091_));
  AOI21X1  g09089(.A0(new_n3505_), .A1(new_n10091_), .B0(new_n3504_), .Y(new_n10092_));
  XOR2X1   g09090(.A(new_n10092_), .B(new_n10090_), .Y(new_n10093_));
  AND2X1   g09091(.A(new_n3513_), .B(new_n3512_), .Y(new_n10094_));
  OAI22X1  g09092(.A0(new_n3521_), .A1(new_n3507_), .B0(new_n3514_), .B1(new_n10094_), .Y(new_n10095_));
  AND2X1   g09093(.A(new_n10092_), .B(new_n10095_), .Y(new_n10096_));
  NOR2X1   g09094(.A(new_n10092_), .B(new_n10095_), .Y(new_n10097_));
  NOR4X1   g09095(.A(new_n10097_), .B(new_n10096_), .C(new_n10087_), .D(new_n3525_), .Y(new_n10098_));
  AOI21X1  g09096(.A0(new_n10093_), .A1(new_n10088_), .B0(new_n10098_), .Y(new_n10099_));
  AOI21X1  g09097(.A0(new_n3471_), .A1(new_n3465_), .B0(new_n3459_), .Y(new_n10100_));
  OR2X1    g09098(.A(new_n10100_), .B(new_n3488_), .Y(new_n10101_));
  XOR2X1   g09099(.A(new_n2666_), .B(new_n2660_), .Y(new_n10102_));
  AOI21X1  g09100(.A0(new_n3470_), .A1(new_n10102_), .B0(new_n3469_), .Y(new_n10103_));
  AOI21X1  g09101(.A0(new_n3458_), .A1(new_n3474_), .B0(new_n3457_), .Y(new_n10104_));
  XOR2X1   g09102(.A(new_n10104_), .B(new_n10103_), .Y(new_n10105_));
  AND2X1   g09103(.A(new_n3467_), .B(new_n3466_), .Y(new_n10106_));
  OAI22X1  g09104(.A0(new_n3485_), .A1(new_n3462_), .B0(new_n3468_), .B1(new_n10106_), .Y(new_n10107_));
  AND2X1   g09105(.A(new_n10104_), .B(new_n10107_), .Y(new_n10108_));
  NOR2X1   g09106(.A(new_n10104_), .B(new_n10107_), .Y(new_n10109_));
  NOR4X1   g09107(.A(new_n10109_), .B(new_n10108_), .C(new_n10100_), .D(new_n3488_), .Y(new_n10110_));
  AOI21X1  g09108(.A0(new_n10105_), .A1(new_n10101_), .B0(new_n10110_), .Y(new_n10111_));
  XOR2X1   g09109(.A(new_n10111_), .B(new_n10099_), .Y(new_n10112_));
  XOR2X1   g09110(.A(new_n10112_), .B(new_n10086_), .Y(new_n10113_));
  OAI21X1  g09111(.A0(new_n3628_), .A1(new_n3617_), .B0(new_n3619_), .Y(new_n10114_));
  AOI21X1  g09112(.A0(new_n3555_), .A1(new_n3549_), .B0(new_n3544_), .Y(new_n10115_));
  OR2X1    g09113(.A(new_n10115_), .B(new_n3563_), .Y(new_n10116_));
  XOR2X1   g09114(.A(new_n2628_), .B(new_n3546_), .Y(new_n10117_));
  AOI21X1  g09115(.A0(new_n3554_), .A1(new_n10117_), .B0(new_n3553_), .Y(new_n10118_));
  XOR2X1   g09116(.A(new_n2646_), .B(new_n2640_), .Y(new_n10119_));
  AOI21X1  g09117(.A0(new_n3543_), .A1(new_n10119_), .B0(new_n3542_), .Y(new_n10120_));
  XOR2X1   g09118(.A(new_n10120_), .B(new_n10118_), .Y(new_n10121_));
  AND2X1   g09119(.A(new_n3551_), .B(new_n3550_), .Y(new_n10122_));
  OAI22X1  g09120(.A0(new_n3559_), .A1(new_n3545_), .B0(new_n3552_), .B1(new_n10122_), .Y(new_n10123_));
  AND2X1   g09121(.A(new_n10120_), .B(new_n10123_), .Y(new_n10124_));
  NOR2X1   g09122(.A(new_n10120_), .B(new_n10123_), .Y(new_n10125_));
  NOR4X1   g09123(.A(new_n10125_), .B(new_n10124_), .C(new_n10115_), .D(new_n3563_), .Y(new_n10126_));
  AOI21X1  g09124(.A0(new_n10121_), .A1(new_n10116_), .B0(new_n10126_), .Y(new_n10127_));
  AOI21X1  g09125(.A0(new_n3586_), .A1(new_n3580_), .B0(new_n3574_), .Y(new_n10128_));
  OR2X1    g09126(.A(new_n10128_), .B(new_n3603_), .Y(new_n10129_));
  XOR2X1   g09127(.A(new_n2590_), .B(new_n2584_), .Y(new_n10130_));
  AOI21X1  g09128(.A0(new_n3585_), .A1(new_n10130_), .B0(new_n3584_), .Y(new_n10131_));
  AOI21X1  g09129(.A0(new_n3573_), .A1(new_n3589_), .B0(new_n3572_), .Y(new_n10132_));
  XOR2X1   g09130(.A(new_n10132_), .B(new_n10131_), .Y(new_n10133_));
  AND2X1   g09131(.A(new_n3582_), .B(new_n3581_), .Y(new_n10134_));
  OAI22X1  g09132(.A0(new_n3600_), .A1(new_n3577_), .B0(new_n3583_), .B1(new_n10134_), .Y(new_n10135_));
  AND2X1   g09133(.A(new_n10132_), .B(new_n10135_), .Y(new_n10136_));
  NOR2X1   g09134(.A(new_n10132_), .B(new_n10135_), .Y(new_n10137_));
  NOR4X1   g09135(.A(new_n10137_), .B(new_n10136_), .C(new_n10128_), .D(new_n3603_), .Y(new_n10138_));
  AOI21X1  g09136(.A0(new_n10133_), .A1(new_n10129_), .B0(new_n10138_), .Y(new_n10139_));
  XOR2X1   g09137(.A(new_n10139_), .B(new_n10127_), .Y(new_n10140_));
  XOR2X1   g09138(.A(new_n10140_), .B(new_n10114_), .Y(new_n10141_));
  XOR2X1   g09139(.A(new_n10141_), .B(new_n10113_), .Y(new_n10142_));
  XOR2X1   g09140(.A(new_n10142_), .B(new_n10084_), .Y(new_n10143_));
  XOR2X1   g09141(.A(new_n10143_), .B(new_n10083_), .Y(new_n10144_));
  XOR2X1   g09142(.A(new_n10144_), .B(new_n10022_), .Y(new_n10145_));
  OAI21X1  g09143(.A0(new_n3436_), .A1(new_n3232_), .B0(new_n3446_), .Y(new_n10146_));
  AOI21X1  g09144(.A0(new_n3229_), .A1(new_n3431_), .B0(new_n3433_), .Y(new_n10147_));
  AOI21X1  g09145(.A0(new_n3182_), .A1(new_n3166_), .B0(new_n3189_), .Y(new_n10148_));
  AOI21X1  g09146(.A0(new_n3225_), .A1(new_n3220_), .B0(new_n10148_), .Y(new_n10149_));
  AOI21X1  g09147(.A0(new_n3210_), .A1(new_n3204_), .B0(new_n3199_), .Y(new_n10150_));
  OR2X1    g09148(.A(new_n10150_), .B(new_n3218_), .Y(new_n10151_));
  XOR2X1   g09149(.A(new_n3013_), .B(new_n3201_), .Y(new_n10152_));
  AOI21X1  g09150(.A0(new_n3209_), .A1(new_n10152_), .B0(new_n3208_), .Y(new_n10153_));
  XOR2X1   g09151(.A(new_n3031_), .B(new_n3025_), .Y(new_n10154_));
  AOI21X1  g09152(.A0(new_n3198_), .A1(new_n10154_), .B0(new_n3197_), .Y(new_n10155_));
  XOR2X1   g09153(.A(new_n10155_), .B(new_n10153_), .Y(new_n10156_));
  AND2X1   g09154(.A(new_n3206_), .B(new_n3205_), .Y(new_n10157_));
  OAI22X1  g09155(.A0(new_n3214_), .A1(new_n3200_), .B0(new_n3207_), .B1(new_n10157_), .Y(new_n10158_));
  AND2X1   g09156(.A(new_n10155_), .B(new_n10158_), .Y(new_n10159_));
  NOR2X1   g09157(.A(new_n10155_), .B(new_n10158_), .Y(new_n10160_));
  NOR4X1   g09158(.A(new_n10160_), .B(new_n10159_), .C(new_n10150_), .D(new_n3218_), .Y(new_n10161_));
  AOI21X1  g09159(.A0(new_n10156_), .A1(new_n10151_), .B0(new_n10161_), .Y(new_n10162_));
  AOI21X1  g09160(.A0(new_n3164_), .A1(new_n3158_), .B0(new_n3152_), .Y(new_n10163_));
  OR2X1    g09161(.A(new_n10163_), .B(new_n3181_), .Y(new_n10164_));
  XOR2X1   g09162(.A(new_n2974_), .B(new_n2968_), .Y(new_n10165_));
  AOI21X1  g09163(.A0(new_n3163_), .A1(new_n10165_), .B0(new_n3162_), .Y(new_n10166_));
  AOI21X1  g09164(.A0(new_n3151_), .A1(new_n3167_), .B0(new_n3150_), .Y(new_n10167_));
  XOR2X1   g09165(.A(new_n10167_), .B(new_n10166_), .Y(new_n10168_));
  AND2X1   g09166(.A(new_n3160_), .B(new_n3159_), .Y(new_n10169_));
  OAI22X1  g09167(.A0(new_n3178_), .A1(new_n3155_), .B0(new_n3161_), .B1(new_n10169_), .Y(new_n10170_));
  AND2X1   g09168(.A(new_n10167_), .B(new_n10170_), .Y(new_n10171_));
  NOR2X1   g09169(.A(new_n10167_), .B(new_n10170_), .Y(new_n10172_));
  NOR4X1   g09170(.A(new_n10172_), .B(new_n10171_), .C(new_n10163_), .D(new_n3181_), .Y(new_n10173_));
  AOI21X1  g09171(.A0(new_n10168_), .A1(new_n10164_), .B0(new_n10173_), .Y(new_n10174_));
  XOR2X1   g09172(.A(new_n10174_), .B(new_n10162_), .Y(new_n10175_));
  XOR2X1   g09173(.A(new_n10175_), .B(new_n10149_), .Y(new_n10176_));
  AOI21X1  g09174(.A0(new_n3138_), .A1(new_n3128_), .B0(new_n3130_), .Y(new_n10177_));
  AOI21X1  g09175(.A0(new_n3067_), .A1(new_n3061_), .B0(new_n3055_), .Y(new_n10178_));
  OR2X1    g09176(.A(new_n10178_), .B(new_n3076_), .Y(new_n10179_));
  XOR2X1   g09177(.A(new_n2936_), .B(new_n3058_), .Y(new_n10180_));
  AOI21X1  g09178(.A0(new_n3066_), .A1(new_n10180_), .B0(new_n3065_), .Y(new_n10181_));
  XOR2X1   g09179(.A(new_n2954_), .B(new_n2948_), .Y(new_n10182_));
  AOI21X1  g09180(.A0(new_n3054_), .A1(new_n10182_), .B0(new_n3053_), .Y(new_n10183_));
  XOR2X1   g09181(.A(new_n10183_), .B(new_n10181_), .Y(new_n10184_));
  AND2X1   g09182(.A(new_n3063_), .B(new_n3062_), .Y(new_n10185_));
  OAI22X1  g09183(.A0(new_n3072_), .A1(new_n3057_), .B0(new_n3064_), .B1(new_n10185_), .Y(new_n10186_));
  AND2X1   g09184(.A(new_n10183_), .B(new_n10186_), .Y(new_n10187_));
  NOR2X1   g09185(.A(new_n10183_), .B(new_n10186_), .Y(new_n10188_));
  NOR4X1   g09186(.A(new_n10188_), .B(new_n10187_), .C(new_n10178_), .D(new_n3076_), .Y(new_n10189_));
  AOI21X1  g09187(.A0(new_n10184_), .A1(new_n10179_), .B0(new_n10189_), .Y(new_n10190_));
  AOI21X1  g09188(.A0(new_n3099_), .A1(new_n3093_), .B0(new_n3087_), .Y(new_n10191_));
  OR2X1    g09189(.A(new_n10191_), .B(new_n3123_), .Y(new_n10192_));
  XOR2X1   g09190(.A(new_n2898_), .B(new_n2892_), .Y(new_n10193_));
  AOI21X1  g09191(.A0(new_n3098_), .A1(new_n10193_), .B0(new_n3097_), .Y(new_n10194_));
  AOI21X1  g09192(.A0(new_n3086_), .A1(new_n3117_), .B0(new_n3085_), .Y(new_n10195_));
  XOR2X1   g09193(.A(new_n10195_), .B(new_n10194_), .Y(new_n10196_));
  AND2X1   g09194(.A(new_n3095_), .B(new_n3094_), .Y(new_n10197_));
  OAI22X1  g09195(.A0(new_n3104_), .A1(new_n3090_), .B0(new_n3096_), .B1(new_n10197_), .Y(new_n10198_));
  AND2X1   g09196(.A(new_n10195_), .B(new_n10198_), .Y(new_n10199_));
  NOR2X1   g09197(.A(new_n10195_), .B(new_n10198_), .Y(new_n10200_));
  NOR4X1   g09198(.A(new_n10200_), .B(new_n10199_), .C(new_n10191_), .D(new_n3123_), .Y(new_n10201_));
  AOI21X1  g09199(.A0(new_n10196_), .A1(new_n10192_), .B0(new_n10201_), .Y(new_n10202_));
  XOR2X1   g09200(.A(new_n10202_), .B(new_n10190_), .Y(new_n10203_));
  XOR2X1   g09201(.A(new_n10203_), .B(new_n10177_), .Y(new_n10204_));
  XOR2X1   g09202(.A(new_n10204_), .B(new_n10176_), .Y(new_n10205_));
  XOR2X1   g09203(.A(new_n10205_), .B(new_n10147_), .Y(new_n10206_));
  AOI21X1  g09204(.A0(new_n3416_), .A1(new_n3318_), .B0(new_n3427_), .Y(new_n10207_));
  AOI21X1  g09205(.A0(new_n3271_), .A1(new_n3255_), .B0(new_n3279_), .Y(new_n10208_));
  AOI21X1  g09206(.A0(new_n3315_), .A1(new_n3310_), .B0(new_n10208_), .Y(new_n10209_));
  AOI21X1  g09207(.A0(new_n3300_), .A1(new_n3294_), .B0(new_n3289_), .Y(new_n10210_));
  OR2X1    g09208(.A(new_n10210_), .B(new_n3308_), .Y(new_n10211_));
  XOR2X1   g09209(.A(new_n2859_), .B(new_n3291_), .Y(new_n10212_));
  AOI21X1  g09210(.A0(new_n3299_), .A1(new_n10212_), .B0(new_n3298_), .Y(new_n10213_));
  XOR2X1   g09211(.A(new_n2877_), .B(new_n2871_), .Y(new_n10214_));
  AOI21X1  g09212(.A0(new_n3288_), .A1(new_n10214_), .B0(new_n3287_), .Y(new_n10215_));
  XOR2X1   g09213(.A(new_n10215_), .B(new_n10213_), .Y(new_n10216_));
  AND2X1   g09214(.A(new_n3296_), .B(new_n3295_), .Y(new_n10217_));
  OAI22X1  g09215(.A0(new_n3304_), .A1(new_n3290_), .B0(new_n3297_), .B1(new_n10217_), .Y(new_n10218_));
  AND2X1   g09216(.A(new_n10215_), .B(new_n10218_), .Y(new_n10219_));
  NOR2X1   g09217(.A(new_n10215_), .B(new_n10218_), .Y(new_n10220_));
  NOR4X1   g09218(.A(new_n10220_), .B(new_n10219_), .C(new_n10210_), .D(new_n3308_), .Y(new_n10221_));
  AOI21X1  g09219(.A0(new_n10216_), .A1(new_n10211_), .B0(new_n10221_), .Y(new_n10222_));
  AOI21X1  g09220(.A0(new_n3253_), .A1(new_n3247_), .B0(new_n3241_), .Y(new_n10223_));
  OR2X1    g09221(.A(new_n10223_), .B(new_n3270_), .Y(new_n10224_));
  XOR2X1   g09222(.A(new_n2821_), .B(new_n2815_), .Y(new_n10225_));
  AOI21X1  g09223(.A0(new_n3252_), .A1(new_n10225_), .B0(new_n3251_), .Y(new_n10226_));
  AOI21X1  g09224(.A0(new_n3240_), .A1(new_n3256_), .B0(new_n3239_), .Y(new_n10227_));
  XOR2X1   g09225(.A(new_n10227_), .B(new_n10226_), .Y(new_n10228_));
  AND2X1   g09226(.A(new_n3249_), .B(new_n3248_), .Y(new_n10229_));
  OAI22X1  g09227(.A0(new_n3267_), .A1(new_n3244_), .B0(new_n3250_), .B1(new_n10229_), .Y(new_n10230_));
  AND2X1   g09228(.A(new_n10227_), .B(new_n10230_), .Y(new_n10231_));
  NOR2X1   g09229(.A(new_n10227_), .B(new_n10230_), .Y(new_n10232_));
  NOR4X1   g09230(.A(new_n10232_), .B(new_n10231_), .C(new_n10223_), .D(new_n3270_), .Y(new_n10233_));
  AOI21X1  g09231(.A0(new_n10228_), .A1(new_n10224_), .B0(new_n10233_), .Y(new_n10234_));
  XOR2X1   g09232(.A(new_n10234_), .B(new_n10222_), .Y(new_n10235_));
  XOR2X1   g09233(.A(new_n10235_), .B(new_n10209_), .Y(new_n10236_));
  OAI21X1  g09234(.A0(new_n3401_), .A1(new_n3350_), .B0(new_n3410_), .Y(new_n10237_));
  AOI21X1  g09235(.A0(new_n3339_), .A1(new_n3333_), .B0(new_n3327_), .Y(new_n10238_));
  OR2X1    g09236(.A(new_n10238_), .B(new_n3348_), .Y(new_n10239_));
  XOR2X1   g09237(.A(new_n2783_), .B(new_n3330_), .Y(new_n10240_));
  AOI21X1  g09238(.A0(new_n3338_), .A1(new_n10240_), .B0(new_n3337_), .Y(new_n10241_));
  XOR2X1   g09239(.A(new_n2801_), .B(new_n2795_), .Y(new_n10242_));
  AOI21X1  g09240(.A0(new_n3326_), .A1(new_n10242_), .B0(new_n3325_), .Y(new_n10243_));
  XOR2X1   g09241(.A(new_n10243_), .B(new_n10241_), .Y(new_n10244_));
  AND2X1   g09242(.A(new_n3335_), .B(new_n3334_), .Y(new_n10245_));
  OAI22X1  g09243(.A0(new_n3344_), .A1(new_n3329_), .B0(new_n3336_), .B1(new_n10245_), .Y(new_n10246_));
  AND2X1   g09244(.A(new_n10243_), .B(new_n10246_), .Y(new_n10247_));
  NOR2X1   g09245(.A(new_n10243_), .B(new_n10246_), .Y(new_n10248_));
  NOR4X1   g09246(.A(new_n10248_), .B(new_n10247_), .C(new_n10238_), .D(new_n3348_), .Y(new_n10249_));
  AOI21X1  g09247(.A0(new_n10244_), .A1(new_n10239_), .B0(new_n10249_), .Y(new_n10250_));
  AOI21X1  g09248(.A0(new_n3371_), .A1(new_n3365_), .B0(new_n3359_), .Y(new_n10251_));
  OR2X1    g09249(.A(new_n10251_), .B(new_n3395_), .Y(new_n10252_));
  XOR2X1   g09250(.A(new_n2745_), .B(new_n2739_), .Y(new_n10253_));
  AOI21X1  g09251(.A0(new_n3370_), .A1(new_n10253_), .B0(new_n3369_), .Y(new_n10254_));
  AOI21X1  g09252(.A0(new_n3358_), .A1(new_n3389_), .B0(new_n3357_), .Y(new_n10255_));
  XOR2X1   g09253(.A(new_n10255_), .B(new_n10254_), .Y(new_n10256_));
  AND2X1   g09254(.A(new_n3367_), .B(new_n3366_), .Y(new_n10257_));
  OAI22X1  g09255(.A0(new_n3376_), .A1(new_n3362_), .B0(new_n3368_), .B1(new_n10257_), .Y(new_n10258_));
  AND2X1   g09256(.A(new_n10255_), .B(new_n10258_), .Y(new_n10259_));
  NOR2X1   g09257(.A(new_n10255_), .B(new_n10258_), .Y(new_n10260_));
  NOR4X1   g09258(.A(new_n10260_), .B(new_n10259_), .C(new_n10251_), .D(new_n3395_), .Y(new_n10261_));
  AOI21X1  g09259(.A0(new_n10256_), .A1(new_n10252_), .B0(new_n10261_), .Y(new_n10262_));
  XOR2X1   g09260(.A(new_n10262_), .B(new_n10250_), .Y(new_n10263_));
  XOR2X1   g09261(.A(new_n10263_), .B(new_n10237_), .Y(new_n10264_));
  XOR2X1   g09262(.A(new_n10264_), .B(new_n10236_), .Y(new_n10265_));
  XOR2X1   g09263(.A(new_n10265_), .B(new_n10207_), .Y(new_n10266_));
  XOR2X1   g09264(.A(new_n10266_), .B(new_n10206_), .Y(new_n10267_));
  XOR2X1   g09265(.A(new_n10267_), .B(new_n10146_), .Y(new_n10268_));
  XOR2X1   g09266(.A(new_n10268_), .B(new_n10145_), .Y(new_n10269_));
  XOR2X1   g09267(.A(new_n10269_), .B(new_n10021_), .Y(new_n10270_));
  AOI21X1  g09268(.A0(new_n2396_), .A1(new_n2388_), .B0(new_n2409_), .Y(new_n10271_));
  AOI21X1  g09269(.A0(new_n2421_), .A1(new_n1695_), .B0(new_n10271_), .Y(new_n10272_));
  AOI21X1  g09270(.A0(new_n2417_), .A1(new_n1691_), .B0(new_n1693_), .Y(new_n10273_));
  OAI21X1  g09271(.A0(new_n1688_), .A1(new_n2412_), .B0(new_n2414_), .Y(new_n10274_));
  AOI21X1  g09272(.A0(new_n1641_), .A1(new_n1625_), .B0(new_n1648_), .Y(new_n10275_));
  AOI21X1  g09273(.A0(new_n1684_), .A1(new_n1679_), .B0(new_n10275_), .Y(new_n10276_));
  AOI21X1  g09274(.A0(new_n1669_), .A1(new_n1663_), .B0(new_n1658_), .Y(new_n10277_));
  OR2X1    g09275(.A(new_n10277_), .B(new_n1677_), .Y(new_n10278_));
  XOR2X1   g09276(.A(new_n1468_), .B(new_n1660_), .Y(new_n10279_));
  AOI21X1  g09277(.A0(new_n1668_), .A1(new_n10279_), .B0(new_n1667_), .Y(new_n10280_));
  XOR2X1   g09278(.A(new_n1486_), .B(new_n1480_), .Y(new_n10281_));
  AOI21X1  g09279(.A0(new_n1657_), .A1(new_n10281_), .B0(new_n1656_), .Y(new_n10282_));
  XOR2X1   g09280(.A(new_n10282_), .B(new_n10280_), .Y(new_n10283_));
  AND2X1   g09281(.A(new_n1665_), .B(new_n1664_), .Y(new_n10284_));
  OAI22X1  g09282(.A0(new_n1673_), .A1(new_n1659_), .B0(new_n1666_), .B1(new_n10284_), .Y(new_n10285_));
  AND2X1   g09283(.A(new_n10282_), .B(new_n10285_), .Y(new_n10286_));
  NOR2X1   g09284(.A(new_n10282_), .B(new_n10285_), .Y(new_n10287_));
  NOR4X1   g09285(.A(new_n10287_), .B(new_n10286_), .C(new_n10277_), .D(new_n1677_), .Y(new_n10288_));
  AOI21X1  g09286(.A0(new_n10283_), .A1(new_n10278_), .B0(new_n10288_), .Y(new_n10289_));
  AOI21X1  g09287(.A0(new_n1623_), .A1(new_n1617_), .B0(new_n1611_), .Y(new_n10290_));
  OR2X1    g09288(.A(new_n10290_), .B(new_n1640_), .Y(new_n10291_));
  XOR2X1   g09289(.A(new_n1429_), .B(new_n1423_), .Y(new_n10292_));
  AOI21X1  g09290(.A0(new_n1622_), .A1(new_n10292_), .B0(new_n1621_), .Y(new_n10293_));
  AOI21X1  g09291(.A0(new_n1610_), .A1(new_n1626_), .B0(new_n1609_), .Y(new_n10294_));
  XOR2X1   g09292(.A(new_n10294_), .B(new_n10293_), .Y(new_n10295_));
  AND2X1   g09293(.A(new_n1619_), .B(new_n1618_), .Y(new_n10296_));
  OAI22X1  g09294(.A0(new_n1637_), .A1(new_n1614_), .B0(new_n1620_), .B1(new_n10296_), .Y(new_n10297_));
  AND2X1   g09295(.A(new_n10294_), .B(new_n10297_), .Y(new_n10298_));
  NOR2X1   g09296(.A(new_n10294_), .B(new_n10297_), .Y(new_n10299_));
  NOR4X1   g09297(.A(new_n10299_), .B(new_n10298_), .C(new_n10290_), .D(new_n1640_), .Y(new_n10300_));
  AOI21X1  g09298(.A0(new_n10295_), .A1(new_n10291_), .B0(new_n10300_), .Y(new_n10301_));
  XOR2X1   g09299(.A(new_n10301_), .B(new_n10289_), .Y(new_n10302_));
  XOR2X1   g09300(.A(new_n10302_), .B(new_n10276_), .Y(new_n10303_));
  OAI21X1  g09301(.A0(new_n1588_), .A1(new_n1537_), .B0(new_n1598_), .Y(new_n10304_));
  AOI21X1  g09302(.A0(new_n1526_), .A1(new_n1520_), .B0(new_n1514_), .Y(new_n10305_));
  OR2X1    g09303(.A(new_n10305_), .B(new_n1535_), .Y(new_n10306_));
  XOR2X1   g09304(.A(new_n1391_), .B(new_n1517_), .Y(new_n10307_));
  AOI21X1  g09305(.A0(new_n1525_), .A1(new_n10307_), .B0(new_n1524_), .Y(new_n10308_));
  XOR2X1   g09306(.A(new_n1409_), .B(new_n1403_), .Y(new_n10309_));
  AOI21X1  g09307(.A0(new_n1513_), .A1(new_n10309_), .B0(new_n1512_), .Y(new_n10310_));
  XOR2X1   g09308(.A(new_n10310_), .B(new_n10308_), .Y(new_n10311_));
  AND2X1   g09309(.A(new_n1522_), .B(new_n1521_), .Y(new_n10312_));
  OAI22X1  g09310(.A0(new_n1531_), .A1(new_n1516_), .B0(new_n1523_), .B1(new_n10312_), .Y(new_n10313_));
  AND2X1   g09311(.A(new_n10310_), .B(new_n10313_), .Y(new_n10314_));
  NOR2X1   g09312(.A(new_n10310_), .B(new_n10313_), .Y(new_n10315_));
  NOR4X1   g09313(.A(new_n10315_), .B(new_n10314_), .C(new_n10305_), .D(new_n1535_), .Y(new_n10316_));
  AOI21X1  g09314(.A0(new_n10311_), .A1(new_n10306_), .B0(new_n10316_), .Y(new_n10317_));
  AOI21X1  g09315(.A0(new_n1558_), .A1(new_n1552_), .B0(new_n1546_), .Y(new_n10318_));
  OR2X1    g09316(.A(new_n10318_), .B(new_n1582_), .Y(new_n10319_));
  XOR2X1   g09317(.A(new_n1353_), .B(new_n1347_), .Y(new_n10320_));
  AOI21X1  g09318(.A0(new_n1557_), .A1(new_n10320_), .B0(new_n1556_), .Y(new_n10321_));
  AOI21X1  g09319(.A0(new_n1545_), .A1(new_n1576_), .B0(new_n1544_), .Y(new_n10322_));
  XOR2X1   g09320(.A(new_n10322_), .B(new_n10321_), .Y(new_n10323_));
  AND2X1   g09321(.A(new_n1554_), .B(new_n1553_), .Y(new_n10324_));
  OAI22X1  g09322(.A0(new_n1563_), .A1(new_n1549_), .B0(new_n1555_), .B1(new_n10324_), .Y(new_n10325_));
  AND2X1   g09323(.A(new_n10322_), .B(new_n10325_), .Y(new_n10326_));
  NOR2X1   g09324(.A(new_n10322_), .B(new_n10325_), .Y(new_n10327_));
  NOR4X1   g09325(.A(new_n10327_), .B(new_n10326_), .C(new_n10318_), .D(new_n1582_), .Y(new_n10328_));
  AOI21X1  g09326(.A0(new_n10323_), .A1(new_n10319_), .B0(new_n10328_), .Y(new_n10329_));
  XOR2X1   g09327(.A(new_n10329_), .B(new_n10317_), .Y(new_n10330_));
  XOR2X1   g09328(.A(new_n10330_), .B(new_n10304_), .Y(new_n10331_));
  XOR2X1   g09329(.A(new_n10331_), .B(new_n10303_), .Y(new_n10332_));
  XOR2X1   g09330(.A(new_n10332_), .B(new_n10274_), .Y(new_n10333_));
  OAI21X1  g09331(.A0(new_n1337_), .A1(new_n1158_), .B0(new_n1501_), .Y(new_n10334_));
  MX2X1    g09332(.A(new_n1151_), .B(new_n1141_), .S0(new_n1128_), .Y(new_n10335_));
  AOI21X1  g09333(.A0(new_n1154_), .A1(new_n1153_), .B0(new_n1117_), .Y(new_n10336_));
  AOI21X1  g09334(.A0(new_n1155_), .A1(new_n10335_), .B0(new_n10336_), .Y(new_n10337_));
  AOI21X1  g09335(.A0(new_n1140_), .A1(new_n1134_), .B0(new_n1128_), .Y(new_n10338_));
  OR2X1    g09336(.A(new_n10338_), .B(new_n1150_), .Y(new_n10339_));
  XOR2X1   g09337(.A(new_n1089_), .B(new_n1131_), .Y(new_n10340_));
  AOI21X1  g09338(.A0(new_n1139_), .A1(new_n10340_), .B0(new_n1138_), .Y(new_n10341_));
  XOR2X1   g09339(.A(new_n1107_), .B(new_n1101_), .Y(new_n10342_));
  AOI21X1  g09340(.A0(new_n1127_), .A1(new_n10342_), .B0(new_n1126_), .Y(new_n10343_));
  XOR2X1   g09341(.A(new_n10343_), .B(new_n10341_), .Y(new_n10344_));
  AND2X1   g09342(.A(new_n1136_), .B(new_n1135_), .Y(new_n10345_));
  OAI22X1  g09343(.A0(new_n1145_), .A1(new_n1130_), .B0(new_n1137_), .B1(new_n10345_), .Y(new_n10346_));
  AND2X1   g09344(.A(new_n10343_), .B(new_n10346_), .Y(new_n10347_));
  NOR2X1   g09345(.A(new_n10343_), .B(new_n10346_), .Y(new_n10348_));
  NOR4X1   g09346(.A(new_n10348_), .B(new_n10347_), .C(new_n10338_), .D(new_n1150_), .Y(new_n10349_));
  AOI21X1  g09347(.A0(new_n10344_), .A1(new_n10339_), .B0(new_n10349_), .Y(new_n10350_));
  AND2X1   g09348(.A(new_n1060_), .B(new_n1051_), .Y(new_n10351_));
  OR4X1    g09349(.A(new_n1059_), .B(new_n1068_), .C(new_n1067_), .D(new_n1065_), .Y(new_n10352_));
  OAI21X1  g09350(.A0(new_n1059_), .A1(new_n1055_), .B0(new_n1048_), .Y(new_n10353_));
  OAI22X1  g09351(.A0(new_n10353_), .A1(new_n10352_), .B0(new_n10351_), .B1(new_n1030_), .Y(new_n10354_));
  AOI21X1  g09352(.A0(new_n1050_), .A1(new_n1056_), .B0(new_n1055_), .Y(new_n10355_));
  OR2X1    g09353(.A(new_n1065_), .B(new_n1023_), .Y(new_n10356_));
  AND2X1   g09354(.A(new_n10356_), .B(new_n1028_), .Y(new_n10357_));
  XOR2X1   g09355(.A(new_n10357_), .B(new_n10355_), .Y(new_n10358_));
  AND2X1   g09356(.A(new_n10358_), .B(new_n10354_), .Y(new_n10359_));
  NOR2X1   g09357(.A(new_n10351_), .B(new_n1030_), .Y(new_n10360_));
  OAI21X1  g09358(.A0(new_n1065_), .A1(new_n1023_), .B0(new_n1028_), .Y(new_n10361_));
  AND2X1   g09359(.A(new_n10361_), .B(new_n10355_), .Y(new_n10362_));
  OAI22X1  g09360(.A0(new_n10361_), .A1(new_n10355_), .B0(new_n10353_), .B1(new_n10352_), .Y(new_n10363_));
  NOR3X1   g09361(.A(new_n10363_), .B(new_n10362_), .C(new_n10360_), .Y(new_n10364_));
  NOR2X1   g09362(.A(new_n10364_), .B(new_n10359_), .Y(new_n10365_));
  XOR2X1   g09363(.A(new_n10365_), .B(new_n10350_), .Y(new_n10366_));
  XOR2X1   g09364(.A(new_n10366_), .B(new_n10337_), .Y(new_n10367_));
  AOI21X1  g09365(.A0(new_n1315_), .A1(new_n1227_), .B0(new_n1330_), .Y(new_n10368_));
  OAI21X1  g09366(.A0(new_n1221_), .A1(new_n1217_), .B0(new_n1311_), .Y(new_n10369_));
  AND2X1   g09367(.A(new_n1208_), .B(new_n1207_), .Y(new_n10370_));
  OAI22X1  g09368(.A0(new_n1214_), .A1(new_n1219_), .B0(new_n1209_), .B1(new_n10370_), .Y(new_n10371_));
  OR2X1    g09369(.A(new_n1178_), .B(new_n1172_), .Y(new_n10372_));
  AOI22X1  g09370(.A0(new_n1182_), .A1(new_n10372_), .B0(new_n1180_), .B1(new_n1179_), .Y(new_n10373_));
  XOR2X1   g09371(.A(new_n10373_), .B(new_n10371_), .Y(new_n10374_));
  AOI21X1  g09372(.A0(new_n10369_), .A1(new_n1225_), .B0(new_n10374_), .Y(new_n10375_));
  NOR4X1   g09373(.A(new_n1224_), .B(new_n1223_), .C(new_n1222_), .D(new_n1219_), .Y(new_n10376_));
  AND2X1   g09374(.A(new_n10373_), .B(new_n10371_), .Y(new_n10377_));
  NOR2X1   g09375(.A(new_n10373_), .B(new_n10371_), .Y(new_n10378_));
  NOR3X1   g09376(.A(new_n10378_), .B(new_n10377_), .C(new_n10376_), .Y(new_n10379_));
  AND2X1   g09377(.A(new_n10379_), .B(new_n10369_), .Y(new_n10380_));
  OR2X1    g09378(.A(new_n10380_), .B(new_n10375_), .Y(new_n10381_));
  AND2X1   g09379(.A(new_n1285_), .B(new_n1276_), .Y(new_n10382_));
  OR4X1    g09380(.A(new_n1284_), .B(new_n1293_), .C(new_n1292_), .D(new_n1290_), .Y(new_n10383_));
  OAI21X1  g09381(.A0(new_n1284_), .A1(new_n1280_), .B0(new_n1273_), .Y(new_n10384_));
  OAI22X1  g09382(.A0(new_n10384_), .A1(new_n10383_), .B0(new_n10382_), .B1(new_n1255_), .Y(new_n10385_));
  AOI21X1  g09383(.A0(new_n1275_), .A1(new_n1281_), .B0(new_n1280_), .Y(new_n10386_));
  OR2X1    g09384(.A(new_n1290_), .B(new_n1248_), .Y(new_n10387_));
  AND2X1   g09385(.A(new_n10387_), .B(new_n1253_), .Y(new_n10388_));
  XOR2X1   g09386(.A(new_n10388_), .B(new_n10386_), .Y(new_n10389_));
  AND2X1   g09387(.A(new_n10389_), .B(new_n10385_), .Y(new_n10390_));
  NOR2X1   g09388(.A(new_n10382_), .B(new_n1255_), .Y(new_n10391_));
  OAI21X1  g09389(.A0(new_n1290_), .A1(new_n1248_), .B0(new_n1253_), .Y(new_n10392_));
  AND2X1   g09390(.A(new_n10392_), .B(new_n10386_), .Y(new_n10393_));
  OAI22X1  g09391(.A0(new_n10392_), .A1(new_n10386_), .B0(new_n10384_), .B1(new_n10383_), .Y(new_n10394_));
  NOR3X1   g09392(.A(new_n10394_), .B(new_n10393_), .C(new_n10391_), .Y(new_n10395_));
  NOR2X1   g09393(.A(new_n10395_), .B(new_n10390_), .Y(new_n10396_));
  XOR2X1   g09394(.A(new_n10396_), .B(new_n10381_), .Y(new_n10397_));
  XOR2X1   g09395(.A(new_n10397_), .B(new_n10368_), .Y(new_n10398_));
  XOR2X1   g09396(.A(new_n10398_), .B(new_n10367_), .Y(new_n10399_));
  XOR2X1   g09397(.A(new_n10399_), .B(new_n10334_), .Y(new_n10400_));
  XOR2X1   g09398(.A(new_n10400_), .B(new_n10333_), .Y(new_n10401_));
  XOR2X1   g09399(.A(new_n10401_), .B(new_n10273_), .Y(new_n10402_));
  OAI21X1  g09400(.A0(new_n2394_), .A1(new_n2038_), .B0(new_n2407_), .Y(new_n10403_));
  OAI21X1  g09401(.A0(new_n2390_), .A1(new_n2034_), .B0(new_n2036_), .Y(new_n10404_));
  AOI21X1  g09402(.A0(new_n1984_), .A1(new_n1968_), .B0(new_n1992_), .Y(new_n10405_));
  AOI21X1  g09403(.A0(new_n2031_), .A1(new_n2026_), .B0(new_n10405_), .Y(new_n10406_));
  AOI21X1  g09404(.A0(new_n2013_), .A1(new_n2007_), .B0(new_n2002_), .Y(new_n10407_));
  OR2X1    g09405(.A(new_n10407_), .B(new_n2024_), .Y(new_n10408_));
  XOR2X1   g09406(.A(new_n1908_), .B(new_n2004_), .Y(new_n10409_));
  AOI21X1  g09407(.A0(new_n2012_), .A1(new_n10409_), .B0(new_n2011_), .Y(new_n10410_));
  XOR2X1   g09408(.A(new_n1926_), .B(new_n1920_), .Y(new_n10411_));
  AOI21X1  g09409(.A0(new_n2001_), .A1(new_n10411_), .B0(new_n2000_), .Y(new_n10412_));
  XOR2X1   g09410(.A(new_n10412_), .B(new_n10410_), .Y(new_n10413_));
  AND2X1   g09411(.A(new_n2009_), .B(new_n2008_), .Y(new_n10414_));
  OAI22X1  g09412(.A0(new_n2017_), .A1(new_n2003_), .B0(new_n2010_), .B1(new_n10414_), .Y(new_n10415_));
  AND2X1   g09413(.A(new_n10412_), .B(new_n10415_), .Y(new_n10416_));
  NOR2X1   g09414(.A(new_n10412_), .B(new_n10415_), .Y(new_n10417_));
  NOR4X1   g09415(.A(new_n10417_), .B(new_n10416_), .C(new_n10407_), .D(new_n2024_), .Y(new_n10418_));
  AOI21X1  g09416(.A0(new_n10413_), .A1(new_n10408_), .B0(new_n10418_), .Y(new_n10419_));
  AOI21X1  g09417(.A0(new_n1966_), .A1(new_n1960_), .B0(new_n1954_), .Y(new_n10420_));
  OR2X1    g09418(.A(new_n10420_), .B(new_n1983_), .Y(new_n10421_));
  XOR2X1   g09419(.A(new_n1870_), .B(new_n1864_), .Y(new_n10422_));
  AOI21X1  g09420(.A0(new_n1965_), .A1(new_n10422_), .B0(new_n1964_), .Y(new_n10423_));
  AOI21X1  g09421(.A0(new_n1953_), .A1(new_n1969_), .B0(new_n1952_), .Y(new_n10424_));
  XOR2X1   g09422(.A(new_n10424_), .B(new_n10423_), .Y(new_n10425_));
  AND2X1   g09423(.A(new_n1962_), .B(new_n1961_), .Y(new_n10426_));
  OAI22X1  g09424(.A0(new_n1980_), .A1(new_n1957_), .B0(new_n1963_), .B1(new_n10426_), .Y(new_n10427_));
  AND2X1   g09425(.A(new_n10424_), .B(new_n10427_), .Y(new_n10428_));
  NOR2X1   g09426(.A(new_n10424_), .B(new_n10427_), .Y(new_n10429_));
  NOR4X1   g09427(.A(new_n10429_), .B(new_n10428_), .C(new_n10420_), .D(new_n1983_), .Y(new_n10430_));
  AOI21X1  g09428(.A0(new_n10425_), .A1(new_n10421_), .B0(new_n10430_), .Y(new_n10431_));
  XOR2X1   g09429(.A(new_n10431_), .B(new_n10419_), .Y(new_n10432_));
  XOR2X1   g09430(.A(new_n10432_), .B(new_n10406_), .Y(new_n10433_));
  AOI21X1  g09431(.A0(new_n1940_), .A1(new_n1850_), .B0(new_n1854_), .Y(new_n10434_));
  OAI21X1  g09432(.A0(new_n1760_), .A1(new_n1756_), .B0(new_n1722_), .Y(new_n10435_));
  AND2X1   g09433(.A(new_n1746_), .B(new_n1745_), .Y(new_n10436_));
  OAI22X1  g09434(.A0(new_n1752_), .A1(new_n1758_), .B0(new_n1747_), .B1(new_n10436_), .Y(new_n10437_));
  OR2X1    g09435(.A(new_n1715_), .B(new_n1709_), .Y(new_n10438_));
  AOI22X1  g09436(.A0(new_n1719_), .A1(new_n10438_), .B0(new_n1717_), .B1(new_n1716_), .Y(new_n10439_));
  XOR2X1   g09437(.A(new_n10439_), .B(new_n10437_), .Y(new_n10440_));
  AOI21X1  g09438(.A0(new_n10435_), .A1(new_n1764_), .B0(new_n10440_), .Y(new_n10441_));
  NOR4X1   g09439(.A(new_n1763_), .B(new_n1762_), .C(new_n1761_), .D(new_n1758_), .Y(new_n10442_));
  AND2X1   g09440(.A(new_n10439_), .B(new_n10437_), .Y(new_n10443_));
  NOR2X1   g09441(.A(new_n10439_), .B(new_n10437_), .Y(new_n10444_));
  NOR3X1   g09442(.A(new_n10444_), .B(new_n10443_), .C(new_n10442_), .Y(new_n10445_));
  AND2X1   g09443(.A(new_n10445_), .B(new_n10435_), .Y(new_n10446_));
  OR2X1    g09444(.A(new_n10446_), .B(new_n10441_), .Y(new_n10447_));
  AND2X1   g09445(.A(new_n1824_), .B(new_n1815_), .Y(new_n10448_));
  OR4X1    g09446(.A(new_n1823_), .B(new_n1832_), .C(new_n1831_), .D(new_n1829_), .Y(new_n10449_));
  OAI21X1  g09447(.A0(new_n1823_), .A1(new_n1819_), .B0(new_n1812_), .Y(new_n10450_));
  OAI22X1  g09448(.A0(new_n10450_), .A1(new_n10449_), .B0(new_n10448_), .B1(new_n1794_), .Y(new_n10451_));
  AOI21X1  g09449(.A0(new_n1814_), .A1(new_n1820_), .B0(new_n1819_), .Y(new_n10452_));
  OR2X1    g09450(.A(new_n1829_), .B(new_n1787_), .Y(new_n10453_));
  AND2X1   g09451(.A(new_n10453_), .B(new_n1792_), .Y(new_n10454_));
  XOR2X1   g09452(.A(new_n10454_), .B(new_n10452_), .Y(new_n10455_));
  AND2X1   g09453(.A(new_n10455_), .B(new_n10451_), .Y(new_n10456_));
  NOR2X1   g09454(.A(new_n10448_), .B(new_n1794_), .Y(new_n10457_));
  OAI21X1  g09455(.A0(new_n1829_), .A1(new_n1787_), .B0(new_n1792_), .Y(new_n10458_));
  AND2X1   g09456(.A(new_n10458_), .B(new_n10452_), .Y(new_n10459_));
  OAI22X1  g09457(.A0(new_n10458_), .A1(new_n10452_), .B0(new_n10450_), .B1(new_n10449_), .Y(new_n10460_));
  NOR3X1   g09458(.A(new_n10460_), .B(new_n10459_), .C(new_n10457_), .Y(new_n10461_));
  NOR2X1   g09459(.A(new_n10461_), .B(new_n10456_), .Y(new_n10462_));
  XOR2X1   g09460(.A(new_n10462_), .B(new_n10447_), .Y(new_n10463_));
  XOR2X1   g09461(.A(new_n10463_), .B(new_n10434_), .Y(new_n10464_));
  XOR2X1   g09462(.A(new_n10464_), .B(new_n10433_), .Y(new_n10465_));
  XOR2X1   g09463(.A(new_n10465_), .B(new_n10404_), .Y(new_n10466_));
  AOI21X1  g09464(.A0(new_n2373_), .A1(new_n2194_), .B0(new_n2385_), .Y(new_n10467_));
  MX2X1    g09465(.A(new_n2187_), .B(new_n2177_), .S0(new_n2164_), .Y(new_n10468_));
  AOI21X1  g09466(.A0(new_n2190_), .A1(new_n2189_), .B0(new_n2153_), .Y(new_n10469_));
  AOI21X1  g09467(.A0(new_n2191_), .A1(new_n10468_), .B0(new_n10469_), .Y(new_n10470_));
  AOI21X1  g09468(.A0(new_n2176_), .A1(new_n2170_), .B0(new_n2164_), .Y(new_n10471_));
  OR2X1    g09469(.A(new_n10471_), .B(new_n2186_), .Y(new_n10472_));
  XOR2X1   g09470(.A(new_n2125_), .B(new_n2167_), .Y(new_n10473_));
  AOI21X1  g09471(.A0(new_n2175_), .A1(new_n10473_), .B0(new_n2174_), .Y(new_n10474_));
  XOR2X1   g09472(.A(new_n2143_), .B(new_n2137_), .Y(new_n10475_));
  AOI21X1  g09473(.A0(new_n2163_), .A1(new_n10475_), .B0(new_n2162_), .Y(new_n10476_));
  XOR2X1   g09474(.A(new_n10476_), .B(new_n10474_), .Y(new_n10477_));
  AND2X1   g09475(.A(new_n2172_), .B(new_n2171_), .Y(new_n10478_));
  OAI22X1  g09476(.A0(new_n2181_), .A1(new_n2166_), .B0(new_n2173_), .B1(new_n10478_), .Y(new_n10479_));
  AND2X1   g09477(.A(new_n10476_), .B(new_n10479_), .Y(new_n10480_));
  NOR2X1   g09478(.A(new_n10476_), .B(new_n10479_), .Y(new_n10481_));
  NOR4X1   g09479(.A(new_n10481_), .B(new_n10480_), .C(new_n10471_), .D(new_n2186_), .Y(new_n10482_));
  AOI21X1  g09480(.A0(new_n10477_), .A1(new_n10472_), .B0(new_n10482_), .Y(new_n10483_));
  AND2X1   g09481(.A(new_n2096_), .B(new_n2087_), .Y(new_n10484_));
  OR4X1    g09482(.A(new_n2095_), .B(new_n2104_), .C(new_n2103_), .D(new_n2101_), .Y(new_n10485_));
  OAI21X1  g09483(.A0(new_n2095_), .A1(new_n2091_), .B0(new_n2084_), .Y(new_n10486_));
  OAI22X1  g09484(.A0(new_n10486_), .A1(new_n10485_), .B0(new_n10484_), .B1(new_n2066_), .Y(new_n10487_));
  AOI21X1  g09485(.A0(new_n2086_), .A1(new_n2092_), .B0(new_n2091_), .Y(new_n10488_));
  OR2X1    g09486(.A(new_n2101_), .B(new_n2059_), .Y(new_n10489_));
  AND2X1   g09487(.A(new_n10489_), .B(new_n2064_), .Y(new_n10490_));
  XOR2X1   g09488(.A(new_n10490_), .B(new_n10488_), .Y(new_n10491_));
  AND2X1   g09489(.A(new_n10491_), .B(new_n10487_), .Y(new_n10492_));
  NOR2X1   g09490(.A(new_n10484_), .B(new_n2066_), .Y(new_n10493_));
  OAI21X1  g09491(.A0(new_n2101_), .A1(new_n2059_), .B0(new_n2064_), .Y(new_n10494_));
  AND2X1   g09492(.A(new_n10494_), .B(new_n10488_), .Y(new_n10495_));
  OAI22X1  g09493(.A0(new_n10494_), .A1(new_n10488_), .B0(new_n10486_), .B1(new_n10485_), .Y(new_n10496_));
  NOR3X1   g09494(.A(new_n10496_), .B(new_n10495_), .C(new_n10493_), .Y(new_n10497_));
  NOR2X1   g09495(.A(new_n10497_), .B(new_n10492_), .Y(new_n10498_));
  XOR2X1   g09496(.A(new_n10498_), .B(new_n10483_), .Y(new_n10499_));
  XOR2X1   g09497(.A(new_n10499_), .B(new_n10470_), .Y(new_n10500_));
  AOI21X1  g09498(.A0(new_n2365_), .A1(new_n2349_), .B0(new_n2353_), .Y(new_n10501_));
  OAI21X1  g09499(.A0(new_n2259_), .A1(new_n2255_), .B0(new_n2221_), .Y(new_n10502_));
  AND2X1   g09500(.A(new_n2245_), .B(new_n2244_), .Y(new_n10503_));
  OAI22X1  g09501(.A0(new_n2251_), .A1(new_n2257_), .B0(new_n2246_), .B1(new_n10503_), .Y(new_n10504_));
  OR2X1    g09502(.A(new_n2214_), .B(new_n2208_), .Y(new_n10505_));
  AOI22X1  g09503(.A0(new_n2218_), .A1(new_n10505_), .B0(new_n2216_), .B1(new_n2215_), .Y(new_n10506_));
  XOR2X1   g09504(.A(new_n10506_), .B(new_n10504_), .Y(new_n10507_));
  AOI21X1  g09505(.A0(new_n10502_), .A1(new_n2263_), .B0(new_n10507_), .Y(new_n10508_));
  NOR4X1   g09506(.A(new_n2262_), .B(new_n2261_), .C(new_n2260_), .D(new_n2257_), .Y(new_n10509_));
  AND2X1   g09507(.A(new_n10506_), .B(new_n10504_), .Y(new_n10510_));
  NOR2X1   g09508(.A(new_n10506_), .B(new_n10504_), .Y(new_n10511_));
  NOR3X1   g09509(.A(new_n10511_), .B(new_n10510_), .C(new_n10509_), .Y(new_n10512_));
  AND2X1   g09510(.A(new_n10512_), .B(new_n10502_), .Y(new_n10513_));
  OR2X1    g09511(.A(new_n10513_), .B(new_n10508_), .Y(new_n10514_));
  AND2X1   g09512(.A(new_n2323_), .B(new_n2314_), .Y(new_n10515_));
  OR4X1    g09513(.A(new_n2322_), .B(new_n2331_), .C(new_n2330_), .D(new_n2328_), .Y(new_n10516_));
  OAI21X1  g09514(.A0(new_n2322_), .A1(new_n2318_), .B0(new_n2311_), .Y(new_n10517_));
  OAI22X1  g09515(.A0(new_n10517_), .A1(new_n10516_), .B0(new_n10515_), .B1(new_n2293_), .Y(new_n10518_));
  AOI21X1  g09516(.A0(new_n2313_), .A1(new_n2319_), .B0(new_n2318_), .Y(new_n10519_));
  OR2X1    g09517(.A(new_n2328_), .B(new_n2286_), .Y(new_n10520_));
  AND2X1   g09518(.A(new_n10520_), .B(new_n2291_), .Y(new_n10521_));
  XOR2X1   g09519(.A(new_n10521_), .B(new_n10519_), .Y(new_n10522_));
  AND2X1   g09520(.A(new_n10522_), .B(new_n10518_), .Y(new_n10523_));
  NOR2X1   g09521(.A(new_n10515_), .B(new_n2293_), .Y(new_n10524_));
  OAI21X1  g09522(.A0(new_n2328_), .A1(new_n2286_), .B0(new_n2291_), .Y(new_n10525_));
  AND2X1   g09523(.A(new_n10525_), .B(new_n10519_), .Y(new_n10526_));
  OAI22X1  g09524(.A0(new_n10525_), .A1(new_n10519_), .B0(new_n10517_), .B1(new_n10516_), .Y(new_n10527_));
  NOR3X1   g09525(.A(new_n10527_), .B(new_n10526_), .C(new_n10524_), .Y(new_n10528_));
  NOR2X1   g09526(.A(new_n10528_), .B(new_n10523_), .Y(new_n10529_));
  XOR2X1   g09527(.A(new_n10529_), .B(new_n10514_), .Y(new_n10530_));
  XOR2X1   g09528(.A(new_n10530_), .B(new_n10501_), .Y(new_n10531_));
  XOR2X1   g09529(.A(new_n10531_), .B(new_n10500_), .Y(new_n10532_));
  XOR2X1   g09530(.A(new_n10532_), .B(new_n10467_), .Y(new_n10533_));
  XOR2X1   g09531(.A(new_n10533_), .B(new_n10466_), .Y(new_n10534_));
  XOR2X1   g09532(.A(new_n10534_), .B(new_n10403_), .Y(new_n10535_));
  XOR2X1   g09533(.A(new_n10535_), .B(new_n10402_), .Y(new_n10536_));
  XOR2X1   g09534(.A(new_n10536_), .B(new_n10272_), .Y(new_n10537_));
  XOR2X1   g09535(.A(new_n10537_), .B(new_n10270_), .Y(new_n10538_));
  XOR2X1   g09536(.A(new_n10538_), .B(new_n10010_), .Y(new_n10539_));
  NAND2X1  g09537(.A(new_n10539_), .B(new_n10007_), .Y(new_n10540_));
  OAI21X1  g09538(.A0(new_n4923_), .A1(new_n4919_), .B0(new_n5248_), .Y(new_n10541_));
  OAI21X1  g09539(.A0(new_n5246_), .A1(new_n5239_), .B0(new_n5237_), .Y(new_n10542_));
  OAI21X1  g09540(.A0(new_n10542_), .A1(new_n4919_), .B0(new_n5637_), .Y(new_n10543_));
  AND2X1   g09541(.A(new_n10543_), .B(new_n10541_), .Y(new_n10544_));
  XOR2X1   g09542(.A(new_n9232_), .B(new_n10544_), .Y(new_n10545_));
  XOR2X1   g09543(.A(new_n10005_), .B(new_n10545_), .Y(new_n10546_));
  NOR2X1   g09544(.A(new_n10546_), .B(new_n8852_), .Y(new_n10547_));
  AOI21X1  g09545(.A0(new_n8823_), .A1(new_n8810_), .B0(new_n8838_), .Y(new_n10548_));
  AOI21X1  g09546(.A0(new_n8842_), .A1(new_n5642_), .B0(new_n10548_), .Y(new_n10549_));
  OAI21X1  g09547(.A0(new_n10008_), .A1(new_n3842_), .B0(new_n3846_), .Y(new_n10550_));
  XOR2X1   g09548(.A(new_n10538_), .B(new_n10550_), .Y(new_n10551_));
  OAI21X1  g09549(.A0(new_n10006_), .A1(new_n10549_), .B0(new_n10551_), .Y(new_n10552_));
  NOR2X1   g09550(.A(new_n10552_), .B(new_n10547_), .Y(new_n10553_));
  AOI21X1  g09551(.A0(new_n10540_), .A1(new_n8850_), .B0(new_n10553_), .Y(new_n10554_));
  OR2X1    g09552(.A(new_n10005_), .B(new_n10545_), .Y(new_n10555_));
  AND2X1   g09553(.A(new_n10005_), .B(new_n10545_), .Y(new_n10556_));
  AOI21X1  g09554(.A0(new_n10555_), .A1(new_n8852_), .B0(new_n10556_), .Y(new_n10557_));
  OAI21X1  g09555(.A0(new_n8834_), .A1(new_n8769_), .B0(new_n8819_), .Y(new_n10558_));
  AOI22X1  g09556(.A0(new_n10003_), .A1(new_n9623_), .B0(new_n10558_), .B1(new_n8836_), .Y(new_n10559_));
  NOR2X1   g09557(.A(new_n10003_), .B(new_n9623_), .Y(new_n10560_));
  OR2X1    g09558(.A(new_n10560_), .B(new_n10559_), .Y(new_n10561_));
  AOI22X1  g09559(.A0(new_n10001_), .A1(new_n9818_), .B0(new_n9625_), .B1(new_n9624_), .Y(new_n10562_));
  NOR2X1   g09560(.A(new_n10001_), .B(new_n9818_), .Y(new_n10563_));
  OR2X1    g09561(.A(new_n10563_), .B(new_n10562_), .Y(new_n10564_));
  OR2X1    g09562(.A(new_n8720_), .B(new_n8740_), .Y(new_n10565_));
  OAI21X1  g09563(.A0(new_n8741_), .A1(new_n8704_), .B0(new_n8739_), .Y(new_n10566_));
  AND2X1   g09564(.A(new_n8713_), .B(new_n8678_), .Y(new_n10567_));
  AOI21X1  g09565(.A0(new_n8714_), .A1(new_n8710_), .B0(new_n8506_), .Y(new_n10568_));
  OR2X1    g09566(.A(new_n10568_), .B(new_n10567_), .Y(new_n10569_));
  XOR2X1   g09567(.A(new_n9998_), .B(new_n10569_), .Y(new_n10570_));
  AOI22X1  g09568(.A0(new_n10570_), .A1(new_n9913_), .B0(new_n10566_), .B1(new_n10565_), .Y(new_n10571_));
  NOR2X1   g09569(.A(new_n10570_), .B(new_n9913_), .Y(new_n10572_));
  OR2X1    g09570(.A(new_n10572_), .B(new_n10571_), .Y(new_n10573_));
  NOR2X1   g09571(.A(new_n9981_), .B(new_n9976_), .Y(new_n10574_));
  XOR2X1   g09572(.A(new_n9995_), .B(new_n10574_), .Y(new_n10575_));
  XOR2X1   g09573(.A(new_n10575_), .B(new_n9965_), .Y(new_n10576_));
  AOI22X1  g09574(.A0(new_n10576_), .A1(new_n9962_), .B0(new_n9915_), .B1(new_n9914_), .Y(new_n10577_));
  NOR2X1   g09575(.A(new_n10576_), .B(new_n9962_), .Y(new_n10578_));
  OR2X1    g09576(.A(new_n10578_), .B(new_n10577_), .Y(new_n10579_));
  OR2X1    g09577(.A(new_n9994_), .B(new_n9988_), .Y(new_n10580_));
  AOI22X1  g09578(.A0(new_n10580_), .A1(new_n9982_), .B0(new_n9964_), .B1(new_n9963_), .Y(new_n10581_));
  NOR4X1   g09579(.A(new_n9994_), .B(new_n9988_), .C(new_n9981_), .D(new_n9976_), .Y(new_n10582_));
  NAND3X1  g09580(.A(new_n9985_), .B(new_n9984_), .C(new_n9983_), .Y(new_n10583_));
  AOI21X1  g09581(.A0(new_n9984_), .A1(new_n9983_), .B0(new_n9985_), .Y(new_n10584_));
  AOI21X1  g09582(.A0(new_n10583_), .A1(new_n9986_), .B0(new_n10584_), .Y(new_n10585_));
  NAND3X1  g09583(.A(new_n9973_), .B(new_n9972_), .C(new_n9966_), .Y(new_n10586_));
  AOI21X1  g09584(.A0(new_n9972_), .A1(new_n9966_), .B0(new_n9973_), .Y(new_n10587_));
  AOI21X1  g09585(.A0(new_n10586_), .A1(new_n9974_), .B0(new_n10587_), .Y(new_n10588_));
  XOR2X1   g09586(.A(new_n10588_), .B(new_n10585_), .Y(new_n10589_));
  OAI21X1  g09587(.A0(new_n10582_), .A1(new_n10581_), .B0(new_n10589_), .Y(new_n10590_));
  AND2X1   g09588(.A(new_n8684_), .B(new_n8655_), .Y(new_n10591_));
  AOI21X1  g09589(.A0(new_n8690_), .A1(new_n8679_), .B0(new_n8583_), .Y(new_n10592_));
  OAI22X1  g09590(.A0(new_n9995_), .A1(new_n10574_), .B0(new_n10592_), .B1(new_n10591_), .Y(new_n10593_));
  AND2X1   g09591(.A(new_n8665_), .B(new_n8660_), .Y(new_n10594_));
  NOR3X1   g09592(.A(new_n9991_), .B(new_n9989_), .C(new_n10594_), .Y(new_n10595_));
  OAI21X1  g09593(.A0(new_n9989_), .A1(new_n10594_), .B0(new_n9991_), .Y(new_n10596_));
  OAI21X1  g09594(.A0(new_n10595_), .A1(new_n9992_), .B0(new_n10596_), .Y(new_n10597_));
  OR2X1    g09595(.A(new_n10588_), .B(new_n10597_), .Y(new_n10598_));
  AOI21X1  g09596(.A0(new_n10588_), .A1(new_n10597_), .B0(new_n10582_), .Y(new_n10599_));
  NAND3X1  g09597(.A(new_n10599_), .B(new_n10598_), .C(new_n10593_), .Y(new_n10600_));
  NAND2X1  g09598(.A(new_n10600_), .B(new_n10590_), .Y(new_n10601_));
  OR2X1    g09599(.A(new_n9946_), .B(new_n9940_), .Y(new_n10602_));
  OR2X1    g09600(.A(new_n9959_), .B(new_n9953_), .Y(new_n10603_));
  AOI22X1  g09601(.A0(new_n10603_), .A1(new_n10602_), .B0(new_n9928_), .B1(new_n9917_), .Y(new_n10604_));
  NOR4X1   g09602(.A(new_n9959_), .B(new_n9953_), .C(new_n9946_), .D(new_n9940_), .Y(new_n10605_));
  AND2X1   g09603(.A(new_n8750_), .B(new_n8749_), .Y(new_n10606_));
  NOR3X1   g09604(.A(new_n9956_), .B(new_n9954_), .C(new_n10606_), .Y(new_n10607_));
  OAI21X1  g09605(.A0(new_n9954_), .A1(new_n10606_), .B0(new_n9956_), .Y(new_n10608_));
  OAI21X1  g09606(.A0(new_n10607_), .A1(new_n9957_), .B0(new_n10608_), .Y(new_n10609_));
  NAND3X1  g09607(.A(new_n9937_), .B(new_n9936_), .C(new_n9930_), .Y(new_n10610_));
  AOI21X1  g09608(.A0(new_n9936_), .A1(new_n9930_), .B0(new_n9937_), .Y(new_n10611_));
  AOI21X1  g09609(.A0(new_n10610_), .A1(new_n9938_), .B0(new_n10611_), .Y(new_n10612_));
  AND2X1   g09610(.A(new_n10612_), .B(new_n10609_), .Y(new_n10613_));
  NOR2X1   g09611(.A(new_n10612_), .B(new_n10609_), .Y(new_n10614_));
  OAI22X1  g09612(.A0(new_n10614_), .A1(new_n10613_), .B0(new_n10605_), .B1(new_n10604_), .Y(new_n10615_));
  AND2X1   g09613(.A(new_n8461_), .B(new_n8503_), .Y(new_n10616_));
  AOI21X1  g09614(.A0(new_n8504_), .A1(new_n8398_), .B0(new_n8502_), .Y(new_n10617_));
  OAI22X1  g09615(.A0(new_n9960_), .A1(new_n9947_), .B0(new_n10617_), .B1(new_n10616_), .Y(new_n10618_));
  OR4X1    g09616(.A(new_n9959_), .B(new_n9953_), .C(new_n9946_), .D(new_n9940_), .Y(new_n10619_));
  NAND2X1  g09617(.A(new_n10612_), .B(new_n10609_), .Y(new_n10620_));
  OR2X1    g09618(.A(new_n10612_), .B(new_n10609_), .Y(new_n10621_));
  NAND4X1  g09619(.A(new_n10621_), .B(new_n10620_), .C(new_n10619_), .D(new_n10618_), .Y(new_n10622_));
  AND2X1   g09620(.A(new_n10622_), .B(new_n10615_), .Y(new_n10623_));
  XOR2X1   g09621(.A(new_n10623_), .B(new_n10601_), .Y(new_n10624_));
  XOR2X1   g09622(.A(new_n10624_), .B(new_n10579_), .Y(new_n10625_));
  OR2X1    g09623(.A(new_n9860_), .B(new_n9855_), .Y(new_n10626_));
  XOR2X1   g09624(.A(new_n9874_), .B(new_n10626_), .Y(new_n10627_));
  XOR2X1   g09625(.A(new_n10627_), .B(new_n9844_), .Y(new_n10628_));
  OAI22X1  g09626(.A0(new_n9911_), .A1(new_n10628_), .B0(new_n9823_), .B1(new_n9822_), .Y(new_n10629_));
  NOR2X1   g09627(.A(new_n9895_), .B(new_n9890_), .Y(new_n10630_));
  XOR2X1   g09628(.A(new_n9909_), .B(new_n10630_), .Y(new_n10631_));
  XOR2X1   g09629(.A(new_n10631_), .B(new_n9879_), .Y(new_n10632_));
  OR2X1    g09630(.A(new_n10632_), .B(new_n9876_), .Y(new_n10633_));
  AND2X1   g09631(.A(new_n10633_), .B(new_n10629_), .Y(new_n10634_));
  OR2X1    g09632(.A(new_n9908_), .B(new_n9902_), .Y(new_n10635_));
  AOI22X1  g09633(.A0(new_n10635_), .A1(new_n9896_), .B0(new_n9878_), .B1(new_n9877_), .Y(new_n10636_));
  NOR4X1   g09634(.A(new_n9908_), .B(new_n9902_), .C(new_n9895_), .D(new_n9890_), .Y(new_n10637_));
  NAND3X1  g09635(.A(new_n9899_), .B(new_n9898_), .C(new_n9897_), .Y(new_n10638_));
  AOI21X1  g09636(.A0(new_n9898_), .A1(new_n9897_), .B0(new_n9899_), .Y(new_n10639_));
  AOI21X1  g09637(.A0(new_n10638_), .A1(new_n9900_), .B0(new_n10639_), .Y(new_n10640_));
  NAND3X1  g09638(.A(new_n9887_), .B(new_n9886_), .C(new_n9880_), .Y(new_n10641_));
  AOI21X1  g09639(.A0(new_n9886_), .A1(new_n9880_), .B0(new_n9887_), .Y(new_n10642_));
  AOI21X1  g09640(.A0(new_n10641_), .A1(new_n9888_), .B0(new_n10642_), .Y(new_n10643_));
  XOR2X1   g09641(.A(new_n10643_), .B(new_n10640_), .Y(new_n10644_));
  OAI21X1  g09642(.A0(new_n10637_), .A1(new_n10636_), .B0(new_n10644_), .Y(new_n10645_));
  AND2X1   g09643(.A(new_n8137_), .B(new_n8227_), .Y(new_n10646_));
  AOI21X1  g09644(.A0(new_n8732_), .A1(new_n8110_), .B0(new_n8730_), .Y(new_n10647_));
  OAI22X1  g09645(.A0(new_n9909_), .A1(new_n10630_), .B0(new_n10647_), .B1(new_n10646_), .Y(new_n10648_));
  AND2X1   g09646(.A(new_n8221_), .B(new_n8220_), .Y(new_n10649_));
  NOR3X1   g09647(.A(new_n9905_), .B(new_n9903_), .C(new_n10649_), .Y(new_n10650_));
  OAI21X1  g09648(.A0(new_n9903_), .A1(new_n10649_), .B0(new_n9905_), .Y(new_n10651_));
  OAI21X1  g09649(.A0(new_n10650_), .A1(new_n9906_), .B0(new_n10651_), .Y(new_n10652_));
  OR2X1    g09650(.A(new_n10643_), .B(new_n10652_), .Y(new_n10653_));
  AOI21X1  g09651(.A0(new_n10643_), .A1(new_n10652_), .B0(new_n10637_), .Y(new_n10654_));
  NAND3X1  g09652(.A(new_n10654_), .B(new_n10653_), .C(new_n10648_), .Y(new_n10655_));
  NAND2X1  g09653(.A(new_n10655_), .B(new_n10645_), .Y(new_n10656_));
  OR2X1    g09654(.A(new_n9873_), .B(new_n9867_), .Y(new_n10657_));
  AOI22X1  g09655(.A0(new_n10657_), .A1(new_n10626_), .B0(new_n9843_), .B1(new_n9830_), .Y(new_n10658_));
  NOR4X1   g09656(.A(new_n9873_), .B(new_n9867_), .C(new_n9860_), .D(new_n9855_), .Y(new_n10659_));
  AOI21X1  g09657(.A0(new_n9827_), .A1(new_n9826_), .B0(new_n9870_), .Y(new_n10660_));
  AOI21X1  g09658(.A0(new_n10660_), .A1(new_n9863_), .B0(new_n9871_), .Y(new_n10661_));
  AOI21X1  g09659(.A0(new_n9863_), .A1(new_n9862_), .B0(new_n9864_), .Y(new_n10662_));
  NOR2X1   g09660(.A(new_n10662_), .B(new_n10661_), .Y(new_n10663_));
  NAND3X1  g09661(.A(new_n9852_), .B(new_n9851_), .C(new_n9845_), .Y(new_n10664_));
  AOI21X1  g09662(.A0(new_n9851_), .A1(new_n9845_), .B0(new_n9852_), .Y(new_n10665_));
  AOI21X1  g09663(.A0(new_n10664_), .A1(new_n9853_), .B0(new_n10665_), .Y(new_n10666_));
  XOR2X1   g09664(.A(new_n10666_), .B(new_n10663_), .Y(new_n10667_));
  OAI21X1  g09665(.A0(new_n10659_), .A1(new_n10658_), .B0(new_n10667_), .Y(new_n10668_));
  AND2X1   g09666(.A(new_n8284_), .B(new_n8326_), .Y(new_n10669_));
  AOI21X1  g09667(.A0(new_n8327_), .A1(new_n8259_), .B0(new_n8325_), .Y(new_n10670_));
  OAI22X1  g09668(.A0(new_n9874_), .A1(new_n9861_), .B0(new_n10670_), .B1(new_n10669_), .Y(new_n10671_));
  OR4X1    g09669(.A(new_n9873_), .B(new_n9867_), .C(new_n9860_), .D(new_n9855_), .Y(new_n10672_));
  OR2X1    g09670(.A(new_n10662_), .B(new_n10661_), .Y(new_n10673_));
  NAND2X1  g09671(.A(new_n10666_), .B(new_n10673_), .Y(new_n10674_));
  OR2X1    g09672(.A(new_n10666_), .B(new_n10673_), .Y(new_n10675_));
  NAND4X1  g09673(.A(new_n10675_), .B(new_n10674_), .C(new_n10672_), .D(new_n10671_), .Y(new_n10676_));
  AND2X1   g09674(.A(new_n10676_), .B(new_n10668_), .Y(new_n10677_));
  XOR2X1   g09675(.A(new_n10677_), .B(new_n10656_), .Y(new_n10678_));
  XOR2X1   g09676(.A(new_n10678_), .B(new_n10634_), .Y(new_n10679_));
  XOR2X1   g09677(.A(new_n10679_), .B(new_n10625_), .Y(new_n10680_));
  XOR2X1   g09678(.A(new_n10680_), .B(new_n10573_), .Y(new_n10681_));
  AND2X1   g09679(.A(new_n8796_), .B(new_n7731_), .Y(new_n10682_));
  AOI21X1  g09680(.A0(new_n8798_), .A1(new_n8792_), .B0(new_n7966_), .Y(new_n10683_));
  OR2X1    g09681(.A(new_n9632_), .B(new_n7842_), .Y(new_n10684_));
  OAI21X1  g09682(.A0(new_n9645_), .A1(new_n7876_), .B0(new_n7959_), .Y(new_n10685_));
  OAI22X1  g09683(.A0(new_n9646_), .A1(new_n7959_), .B0(new_n10685_), .B1(new_n9648_), .Y(new_n10686_));
  OAI22X1  g09684(.A0(new_n9659_), .A1(new_n9648_), .B0(new_n9646_), .B1(new_n7893_), .Y(new_n10687_));
  MX2X1    g09685(.A(new_n10687_), .B(new_n10686_), .S0(new_n7958_), .Y(new_n10688_));
  OAI21X1  g09686(.A0(new_n9634_), .A1(new_n9628_), .B0(new_n10688_), .Y(new_n10689_));
  AND2X1   g09687(.A(new_n10689_), .B(new_n10684_), .Y(new_n10690_));
  XOR2X1   g09688(.A(new_n9729_), .B(new_n10690_), .Y(new_n10691_));
  OR2X1    g09689(.A(new_n7578_), .B(new_n7739_), .Y(new_n10692_));
  OAI21X1  g09690(.A0(new_n8793_), .A1(new_n7548_), .B0(new_n8791_), .Y(new_n10693_));
  AND2X1   g09691(.A(new_n10693_), .B(new_n10692_), .Y(new_n10694_));
  XOR2X1   g09692(.A(new_n9815_), .B(new_n10694_), .Y(new_n10695_));
  OAI22X1  g09693(.A0(new_n10695_), .A1(new_n10691_), .B0(new_n10683_), .B1(new_n10682_), .Y(new_n10696_));
  OR2X1    g09694(.A(new_n9816_), .B(new_n9730_), .Y(new_n10697_));
  AND2X1   g09695(.A(new_n10697_), .B(new_n10696_), .Y(new_n10698_));
  NOR2X1   g09696(.A(new_n9798_), .B(new_n9793_), .Y(new_n10699_));
  XOR2X1   g09697(.A(new_n9812_), .B(new_n10699_), .Y(new_n10700_));
  XOR2X1   g09698(.A(new_n10700_), .B(new_n9782_), .Y(new_n10701_));
  AOI22X1  g09699(.A0(new_n10701_), .A1(new_n9779_), .B0(new_n10693_), .B1(new_n10692_), .Y(new_n10702_));
  NOR2X1   g09700(.A(new_n10701_), .B(new_n9779_), .Y(new_n10703_));
  OR2X1    g09701(.A(new_n10703_), .B(new_n10702_), .Y(new_n10704_));
  OR2X1    g09702(.A(new_n9811_), .B(new_n9805_), .Y(new_n10705_));
  AOI22X1  g09703(.A0(new_n10705_), .A1(new_n9799_), .B0(new_n9781_), .B1(new_n9780_), .Y(new_n10706_));
  NOR4X1   g09704(.A(new_n9811_), .B(new_n9805_), .C(new_n9798_), .D(new_n9793_), .Y(new_n10707_));
  NAND3X1  g09705(.A(new_n9802_), .B(new_n9801_), .C(new_n9800_), .Y(new_n10708_));
  AOI21X1  g09706(.A0(new_n9801_), .A1(new_n9800_), .B0(new_n9802_), .Y(new_n10709_));
  AOI21X1  g09707(.A0(new_n10708_), .A1(new_n9803_), .B0(new_n10709_), .Y(new_n10710_));
  NAND3X1  g09708(.A(new_n9790_), .B(new_n9789_), .C(new_n9783_), .Y(new_n10711_));
  AOI21X1  g09709(.A0(new_n9789_), .A1(new_n9783_), .B0(new_n9790_), .Y(new_n10712_));
  AOI21X1  g09710(.A0(new_n10711_), .A1(new_n9791_), .B0(new_n10712_), .Y(new_n10713_));
  XOR2X1   g09711(.A(new_n10713_), .B(new_n10710_), .Y(new_n10714_));
  OAI21X1  g09712(.A0(new_n10707_), .A1(new_n10706_), .B0(new_n10714_), .Y(new_n10715_));
  AND2X1   g09713(.A(new_n7560_), .B(new_n7531_), .Y(new_n10716_));
  AOI21X1  g09714(.A0(new_n7566_), .A1(new_n7555_), .B0(new_n7459_), .Y(new_n10717_));
  OAI22X1  g09715(.A0(new_n9812_), .A1(new_n10699_), .B0(new_n10717_), .B1(new_n10716_), .Y(new_n10718_));
  AND2X1   g09716(.A(new_n7541_), .B(new_n7536_), .Y(new_n10719_));
  NOR3X1   g09717(.A(new_n9808_), .B(new_n9806_), .C(new_n10719_), .Y(new_n10720_));
  OAI21X1  g09718(.A0(new_n9806_), .A1(new_n10719_), .B0(new_n9808_), .Y(new_n10721_));
  OAI21X1  g09719(.A0(new_n10720_), .A1(new_n9809_), .B0(new_n10721_), .Y(new_n10722_));
  OR2X1    g09720(.A(new_n10713_), .B(new_n10722_), .Y(new_n10723_));
  AOI21X1  g09721(.A0(new_n10713_), .A1(new_n10722_), .B0(new_n10707_), .Y(new_n10724_));
  NAND3X1  g09722(.A(new_n10724_), .B(new_n10723_), .C(new_n10718_), .Y(new_n10725_));
  NAND2X1  g09723(.A(new_n10725_), .B(new_n10715_), .Y(new_n10726_));
  OR2X1    g09724(.A(new_n9763_), .B(new_n9757_), .Y(new_n10727_));
  OR2X1    g09725(.A(new_n9776_), .B(new_n9770_), .Y(new_n10728_));
  AOI22X1  g09726(.A0(new_n10728_), .A1(new_n10727_), .B0(new_n9745_), .B1(new_n9734_), .Y(new_n10729_));
  NOR4X1   g09727(.A(new_n9776_), .B(new_n9770_), .C(new_n9763_), .D(new_n9757_), .Y(new_n10730_));
  AND2X1   g09728(.A(new_n8783_), .B(new_n8782_), .Y(new_n10731_));
  NOR3X1   g09729(.A(new_n9773_), .B(new_n9771_), .C(new_n10731_), .Y(new_n10732_));
  OAI21X1  g09730(.A0(new_n9771_), .A1(new_n10731_), .B0(new_n9773_), .Y(new_n10733_));
  OAI21X1  g09731(.A0(new_n10732_), .A1(new_n9774_), .B0(new_n10733_), .Y(new_n10734_));
  NAND3X1  g09732(.A(new_n9754_), .B(new_n9753_), .C(new_n9747_), .Y(new_n10735_));
  AOI21X1  g09733(.A0(new_n9753_), .A1(new_n9747_), .B0(new_n9754_), .Y(new_n10736_));
  AOI21X1  g09734(.A0(new_n10735_), .A1(new_n9755_), .B0(new_n10736_), .Y(new_n10737_));
  AND2X1   g09735(.A(new_n10737_), .B(new_n10734_), .Y(new_n10738_));
  NOR2X1   g09736(.A(new_n10737_), .B(new_n10734_), .Y(new_n10739_));
  OAI22X1  g09737(.A0(new_n10739_), .A1(new_n10738_), .B0(new_n10730_), .B1(new_n10729_), .Y(new_n10740_));
  AND2X1   g09738(.A(new_n7337_), .B(new_n7379_), .Y(new_n10741_));
  AOI21X1  g09739(.A0(new_n7380_), .A1(new_n7274_), .B0(new_n7378_), .Y(new_n10742_));
  OAI22X1  g09740(.A0(new_n9777_), .A1(new_n9764_), .B0(new_n10742_), .B1(new_n10741_), .Y(new_n10743_));
  OR4X1    g09741(.A(new_n9776_), .B(new_n9770_), .C(new_n9763_), .D(new_n9757_), .Y(new_n10744_));
  NAND2X1  g09742(.A(new_n10737_), .B(new_n10734_), .Y(new_n10745_));
  OR2X1    g09743(.A(new_n10737_), .B(new_n10734_), .Y(new_n10746_));
  NAND4X1  g09744(.A(new_n10746_), .B(new_n10745_), .C(new_n10744_), .D(new_n10743_), .Y(new_n10747_));
  AND2X1   g09745(.A(new_n10747_), .B(new_n10740_), .Y(new_n10748_));
  XOR2X1   g09746(.A(new_n10748_), .B(new_n10726_), .Y(new_n10749_));
  XOR2X1   g09747(.A(new_n10749_), .B(new_n10704_), .Y(new_n10750_));
  OR2X1    g09748(.A(new_n9677_), .B(new_n9672_), .Y(new_n10751_));
  XOR2X1   g09749(.A(new_n9691_), .B(new_n10751_), .Y(new_n10752_));
  XOR2X1   g09750(.A(new_n10752_), .B(new_n9661_), .Y(new_n10753_));
  OAI22X1  g09751(.A0(new_n9728_), .A1(new_n10753_), .B0(new_n9640_), .B1(new_n9639_), .Y(new_n10754_));
  NOR2X1   g09752(.A(new_n9712_), .B(new_n9707_), .Y(new_n10755_));
  XOR2X1   g09753(.A(new_n9726_), .B(new_n10755_), .Y(new_n10756_));
  XOR2X1   g09754(.A(new_n10756_), .B(new_n9696_), .Y(new_n10757_));
  OR2X1    g09755(.A(new_n10757_), .B(new_n9693_), .Y(new_n10758_));
  AND2X1   g09756(.A(new_n10758_), .B(new_n10754_), .Y(new_n10759_));
  OR2X1    g09757(.A(new_n9725_), .B(new_n9719_), .Y(new_n10760_));
  AOI22X1  g09758(.A0(new_n10760_), .A1(new_n9713_), .B0(new_n9695_), .B1(new_n9694_), .Y(new_n10761_));
  NOR4X1   g09759(.A(new_n9725_), .B(new_n9719_), .C(new_n9712_), .D(new_n9707_), .Y(new_n10762_));
  AOI21X1  g09760(.A0(new_n7846_), .A1(new_n7845_), .B0(new_n9722_), .Y(new_n10763_));
  AOI21X1  g09761(.A0(new_n10763_), .A1(new_n9715_), .B0(new_n9723_), .Y(new_n10764_));
  AOI21X1  g09762(.A0(new_n9715_), .A1(new_n9714_), .B0(new_n9716_), .Y(new_n10765_));
  NOR2X1   g09763(.A(new_n10765_), .B(new_n10764_), .Y(new_n10766_));
  NAND3X1  g09764(.A(new_n9704_), .B(new_n9703_), .C(new_n9697_), .Y(new_n10767_));
  AOI21X1  g09765(.A0(new_n9703_), .A1(new_n9697_), .B0(new_n9704_), .Y(new_n10768_));
  AOI21X1  g09766(.A0(new_n10767_), .A1(new_n9705_), .B0(new_n10768_), .Y(new_n10769_));
  XOR2X1   g09767(.A(new_n10769_), .B(new_n10766_), .Y(new_n10770_));
  OAI21X1  g09768(.A0(new_n10762_), .A1(new_n10761_), .B0(new_n10770_), .Y(new_n10771_));
  AND2X1   g09769(.A(new_n7838_), .B(new_n7860_), .Y(new_n10772_));
  AOI21X1  g09770(.A0(new_n9629_), .A1(new_n7813_), .B0(new_n7859_), .Y(new_n10773_));
  OAI22X1  g09771(.A0(new_n9726_), .A1(new_n10755_), .B0(new_n10773_), .B1(new_n10772_), .Y(new_n10774_));
  OR2X1    g09772(.A(new_n10765_), .B(new_n10764_), .Y(new_n10775_));
  OR2X1    g09773(.A(new_n10769_), .B(new_n10775_), .Y(new_n10776_));
  AOI21X1  g09774(.A0(new_n10769_), .A1(new_n10775_), .B0(new_n10762_), .Y(new_n10777_));
  NAND3X1  g09775(.A(new_n10777_), .B(new_n10776_), .C(new_n10774_), .Y(new_n10778_));
  NAND2X1  g09776(.A(new_n10778_), .B(new_n10771_), .Y(new_n10779_));
  OR2X1    g09777(.A(new_n9690_), .B(new_n9684_), .Y(new_n10780_));
  AOI22X1  g09778(.A0(new_n10780_), .A1(new_n10751_), .B0(new_n9660_), .B1(new_n9647_), .Y(new_n10781_));
  NOR4X1   g09779(.A(new_n9690_), .B(new_n9684_), .C(new_n9677_), .D(new_n9672_), .Y(new_n10782_));
  AOI21X1  g09780(.A0(new_n9644_), .A1(new_n9643_), .B0(new_n9687_), .Y(new_n10783_));
  AOI21X1  g09781(.A0(new_n10783_), .A1(new_n9680_), .B0(new_n9688_), .Y(new_n10784_));
  AOI21X1  g09782(.A0(new_n9680_), .A1(new_n9679_), .B0(new_n9681_), .Y(new_n10785_));
  NOR2X1   g09783(.A(new_n10785_), .B(new_n10784_), .Y(new_n10786_));
  NAND3X1  g09784(.A(new_n9669_), .B(new_n9668_), .C(new_n9662_), .Y(new_n10787_));
  AOI21X1  g09785(.A0(new_n9668_), .A1(new_n9662_), .B0(new_n9669_), .Y(new_n10788_));
  AOI21X1  g09786(.A0(new_n10787_), .A1(new_n9670_), .B0(new_n10788_), .Y(new_n10789_));
  XOR2X1   g09787(.A(new_n10789_), .B(new_n10786_), .Y(new_n10790_));
  OAI21X1  g09788(.A0(new_n10782_), .A1(new_n10781_), .B0(new_n10790_), .Y(new_n10791_));
  AND2X1   g09789(.A(new_n7917_), .B(new_n7959_), .Y(new_n10792_));
  AOI21X1  g09790(.A0(new_n7960_), .A1(new_n7892_), .B0(new_n7958_), .Y(new_n10793_));
  OAI22X1  g09791(.A0(new_n9691_), .A1(new_n9678_), .B0(new_n10793_), .B1(new_n10792_), .Y(new_n10794_));
  OR4X1    g09792(.A(new_n9690_), .B(new_n9684_), .C(new_n9677_), .D(new_n9672_), .Y(new_n10795_));
  OR2X1    g09793(.A(new_n10785_), .B(new_n10784_), .Y(new_n10796_));
  NAND2X1  g09794(.A(new_n10789_), .B(new_n10796_), .Y(new_n10797_));
  OR2X1    g09795(.A(new_n10789_), .B(new_n10796_), .Y(new_n10798_));
  NAND4X1  g09796(.A(new_n10798_), .B(new_n10797_), .C(new_n10795_), .D(new_n10794_), .Y(new_n10799_));
  AND2X1   g09797(.A(new_n10799_), .B(new_n10791_), .Y(new_n10800_));
  XOR2X1   g09798(.A(new_n10800_), .B(new_n10779_), .Y(new_n10801_));
  XOR2X1   g09799(.A(new_n10801_), .B(new_n10759_), .Y(new_n10802_));
  XOR2X1   g09800(.A(new_n10802_), .B(new_n10750_), .Y(new_n10803_));
  XOR2X1   g09801(.A(new_n10803_), .B(new_n10698_), .Y(new_n10804_));
  XOR2X1   g09802(.A(new_n10804_), .B(new_n10681_), .Y(new_n10805_));
  XOR2X1   g09803(.A(new_n10805_), .B(new_n10564_), .Y(new_n10806_));
  AND2X1   g09804(.A(new_n6734_), .B(new_n6713_), .Y(new_n10807_));
  AOI21X1  g09805(.A0(new_n7207_), .A1(new_n6413_), .B0(new_n7206_), .Y(new_n10808_));
  AND2X1   g09806(.A(new_n6980_), .B(new_n6948_), .Y(new_n10809_));
  AOI21X1  g09807(.A0(new_n7204_), .A1(new_n6946_), .B0(new_n7203_), .Y(new_n10810_));
  OR2X1    g09808(.A(new_n10810_), .B(new_n10809_), .Y(new_n10811_));
  XOR2X1   g09809(.A(new_n9437_), .B(new_n10811_), .Y(new_n10812_));
  OR2X1    g09810(.A(new_n6718_), .B(new_n6376_), .Y(new_n10813_));
  OAI21X1  g09811(.A0(new_n6719_), .A1(new_n6715_), .B0(new_n6013_), .Y(new_n10814_));
  AND2X1   g09812(.A(new_n10814_), .B(new_n10813_), .Y(new_n10815_));
  XOR2X1   g09813(.A(new_n9620_), .B(new_n10815_), .Y(new_n10816_));
  OAI22X1  g09814(.A0(new_n10816_), .A1(new_n10812_), .B0(new_n10808_), .B1(new_n10807_), .Y(new_n10817_));
  OR2X1    g09815(.A(new_n9621_), .B(new_n9438_), .Y(new_n10818_));
  AND2X1   g09816(.A(new_n10818_), .B(new_n10817_), .Y(new_n10819_));
  AND2X1   g09817(.A(new_n6369_), .B(new_n6408_), .Y(new_n10820_));
  AOI21X1  g09818(.A0(new_n6716_), .A1(new_n6350_), .B0(new_n6407_), .Y(new_n10821_));
  OR2X1    g09819(.A(new_n10821_), .B(new_n10820_), .Y(new_n10822_));
  XOR2X1   g09820(.A(new_n9618_), .B(new_n10822_), .Y(new_n10823_));
  AOI22X1  g09821(.A0(new_n10823_), .A1(new_n9533_), .B0(new_n10814_), .B1(new_n10813_), .Y(new_n10824_));
  NOR2X1   g09822(.A(new_n10823_), .B(new_n9533_), .Y(new_n10825_));
  OR2X1    g09823(.A(new_n10825_), .B(new_n10824_), .Y(new_n10826_));
  NOR2X1   g09824(.A(new_n9601_), .B(new_n9596_), .Y(new_n10827_));
  XOR2X1   g09825(.A(new_n9615_), .B(new_n10827_), .Y(new_n10828_));
  XOR2X1   g09826(.A(new_n10828_), .B(new_n9585_), .Y(new_n10829_));
  AOI22X1  g09827(.A0(new_n10829_), .A1(new_n9582_), .B0(new_n9535_), .B1(new_n9534_), .Y(new_n10830_));
  NOR2X1   g09828(.A(new_n10829_), .B(new_n9582_), .Y(new_n10831_));
  OR2X1    g09829(.A(new_n10831_), .B(new_n10830_), .Y(new_n10832_));
  OR2X1    g09830(.A(new_n9614_), .B(new_n9608_), .Y(new_n10833_));
  AOI22X1  g09831(.A0(new_n10833_), .A1(new_n9602_), .B0(new_n9584_), .B1(new_n9583_), .Y(new_n10834_));
  NOR4X1   g09832(.A(new_n9614_), .B(new_n9608_), .C(new_n9601_), .D(new_n9596_), .Y(new_n10835_));
  NAND3X1  g09833(.A(new_n9605_), .B(new_n9604_), .C(new_n9603_), .Y(new_n10836_));
  AOI21X1  g09834(.A0(new_n9604_), .A1(new_n9603_), .B0(new_n9605_), .Y(new_n10837_));
  AOI21X1  g09835(.A0(new_n10836_), .A1(new_n9606_), .B0(new_n10837_), .Y(new_n10838_));
  NAND3X1  g09836(.A(new_n9593_), .B(new_n9592_), .C(new_n9586_), .Y(new_n10839_));
  AOI21X1  g09837(.A0(new_n9592_), .A1(new_n9586_), .B0(new_n9593_), .Y(new_n10840_));
  AOI21X1  g09838(.A0(new_n10839_), .A1(new_n9594_), .B0(new_n10840_), .Y(new_n10841_));
  XOR2X1   g09839(.A(new_n10841_), .B(new_n10838_), .Y(new_n10842_));
  OAI21X1  g09840(.A0(new_n10835_), .A1(new_n10834_), .B0(new_n10842_), .Y(new_n10843_));
  AND2X1   g09841(.A(new_n6348_), .B(new_n6366_), .Y(new_n10844_));
  AOI21X1  g09842(.A0(new_n6386_), .A1(new_n6321_), .B0(new_n6384_), .Y(new_n10845_));
  OAI22X1  g09843(.A0(new_n9615_), .A1(new_n10827_), .B0(new_n10845_), .B1(new_n10844_), .Y(new_n10846_));
  AND2X1   g09844(.A(new_n6360_), .B(new_n6359_), .Y(new_n10847_));
  NOR3X1   g09845(.A(new_n9611_), .B(new_n9609_), .C(new_n10847_), .Y(new_n10848_));
  OAI21X1  g09846(.A0(new_n9609_), .A1(new_n10847_), .B0(new_n9611_), .Y(new_n10849_));
  OAI21X1  g09847(.A0(new_n10848_), .A1(new_n9612_), .B0(new_n10849_), .Y(new_n10850_));
  OR2X1    g09848(.A(new_n10841_), .B(new_n10850_), .Y(new_n10851_));
  AOI21X1  g09849(.A0(new_n10841_), .A1(new_n10850_), .B0(new_n10835_), .Y(new_n10852_));
  NAND3X1  g09850(.A(new_n10852_), .B(new_n10851_), .C(new_n10846_), .Y(new_n10853_));
  NAND2X1  g09851(.A(new_n10853_), .B(new_n10843_), .Y(new_n10854_));
  OR2X1    g09852(.A(new_n9566_), .B(new_n9560_), .Y(new_n10855_));
  OR2X1    g09853(.A(new_n9579_), .B(new_n9573_), .Y(new_n10856_));
  AOI22X1  g09854(.A0(new_n10856_), .A1(new_n10855_), .B0(new_n9548_), .B1(new_n9537_), .Y(new_n10857_));
  NOR4X1   g09855(.A(new_n9579_), .B(new_n9573_), .C(new_n9566_), .D(new_n9560_), .Y(new_n10858_));
  AND2X1   g09856(.A(new_n6130_), .B(new_n6126_), .Y(new_n10859_));
  NOR3X1   g09857(.A(new_n9576_), .B(new_n9574_), .C(new_n10859_), .Y(new_n10860_));
  OAI21X1  g09858(.A0(new_n9574_), .A1(new_n10859_), .B0(new_n9576_), .Y(new_n10861_));
  OAI21X1  g09859(.A0(new_n10860_), .A1(new_n9577_), .B0(new_n10861_), .Y(new_n10862_));
  NAND3X1  g09860(.A(new_n9557_), .B(new_n9556_), .C(new_n9550_), .Y(new_n10863_));
  AOI21X1  g09861(.A0(new_n9556_), .A1(new_n9550_), .B0(new_n9557_), .Y(new_n10864_));
  AOI21X1  g09862(.A0(new_n10863_), .A1(new_n9558_), .B0(new_n10864_), .Y(new_n10865_));
  AND2X1   g09863(.A(new_n10865_), .B(new_n10862_), .Y(new_n10866_));
  NOR2X1   g09864(.A(new_n10865_), .B(new_n10862_), .Y(new_n10867_));
  OAI22X1  g09865(.A0(new_n10867_), .A1(new_n10866_), .B0(new_n10858_), .B1(new_n10857_), .Y(new_n10868_));
  AND2X1   g09866(.A(new_n6403_), .B(new_n6121_), .Y(new_n10869_));
  AOI21X1  g09867(.A0(new_n6405_), .A1(new_n6392_), .B0(new_n6176_), .Y(new_n10870_));
  OAI22X1  g09868(.A0(new_n9580_), .A1(new_n9567_), .B0(new_n10870_), .B1(new_n10869_), .Y(new_n10871_));
  OR4X1    g09869(.A(new_n9579_), .B(new_n9573_), .C(new_n9566_), .D(new_n9560_), .Y(new_n10872_));
  NAND2X1  g09870(.A(new_n10865_), .B(new_n10862_), .Y(new_n10873_));
  OR2X1    g09871(.A(new_n10865_), .B(new_n10862_), .Y(new_n10874_));
  NAND4X1  g09872(.A(new_n10874_), .B(new_n10873_), .C(new_n10872_), .D(new_n10871_), .Y(new_n10875_));
  AND2X1   g09873(.A(new_n10875_), .B(new_n10868_), .Y(new_n10876_));
  XOR2X1   g09874(.A(new_n10876_), .B(new_n10854_), .Y(new_n10877_));
  XOR2X1   g09875(.A(new_n10877_), .B(new_n10832_), .Y(new_n10878_));
  OR2X1    g09876(.A(new_n9480_), .B(new_n9475_), .Y(new_n10879_));
  XOR2X1   g09877(.A(new_n9494_), .B(new_n10879_), .Y(new_n10880_));
  XOR2X1   g09878(.A(new_n10880_), .B(new_n9464_), .Y(new_n10881_));
  OAI22X1  g09879(.A0(new_n9531_), .A1(new_n10881_), .B0(new_n9443_), .B1(new_n9442_), .Y(new_n10882_));
  NOR2X1   g09880(.A(new_n9515_), .B(new_n9510_), .Y(new_n10883_));
  XOR2X1   g09881(.A(new_n9529_), .B(new_n10883_), .Y(new_n10884_));
  XOR2X1   g09882(.A(new_n10884_), .B(new_n9499_), .Y(new_n10885_));
  OR2X1    g09883(.A(new_n10885_), .B(new_n9496_), .Y(new_n10886_));
  AND2X1   g09884(.A(new_n10886_), .B(new_n10882_), .Y(new_n10887_));
  OR2X1    g09885(.A(new_n9528_), .B(new_n9522_), .Y(new_n10888_));
  AOI22X1  g09886(.A0(new_n10888_), .A1(new_n9516_), .B0(new_n9498_), .B1(new_n9497_), .Y(new_n10889_));
  NOR4X1   g09887(.A(new_n9528_), .B(new_n9522_), .C(new_n9515_), .D(new_n9510_), .Y(new_n10890_));
  NAND3X1  g09888(.A(new_n9519_), .B(new_n9518_), .C(new_n9517_), .Y(new_n10891_));
  AOI21X1  g09889(.A0(new_n9518_), .A1(new_n9517_), .B0(new_n9519_), .Y(new_n10892_));
  AOI21X1  g09890(.A0(new_n10891_), .A1(new_n9520_), .B0(new_n10892_), .Y(new_n10893_));
  NAND3X1  g09891(.A(new_n9507_), .B(new_n9506_), .C(new_n9500_), .Y(new_n10894_));
  AOI21X1  g09892(.A0(new_n9506_), .A1(new_n9500_), .B0(new_n9507_), .Y(new_n10895_));
  AOI21X1  g09893(.A0(new_n10894_), .A1(new_n9508_), .B0(new_n10895_), .Y(new_n10896_));
  XOR2X1   g09894(.A(new_n10896_), .B(new_n10893_), .Y(new_n10897_));
  OAI21X1  g09895(.A0(new_n10890_), .A1(new_n10889_), .B0(new_n10897_), .Y(new_n10898_));
  AND2X1   g09896(.A(new_n5892_), .B(new_n5791_), .Y(new_n10899_));
  AOI21X1  g09897(.A0(new_n5898_), .A1(new_n5887_), .B0(new_n5719_), .Y(new_n10900_));
  OAI22X1  g09898(.A0(new_n9529_), .A1(new_n10883_), .B0(new_n10900_), .B1(new_n10899_), .Y(new_n10901_));
  AND2X1   g09899(.A(new_n5801_), .B(new_n5796_), .Y(new_n10902_));
  NOR3X1   g09900(.A(new_n9525_), .B(new_n9523_), .C(new_n10902_), .Y(new_n10903_));
  OAI21X1  g09901(.A0(new_n9523_), .A1(new_n10902_), .B0(new_n9525_), .Y(new_n10904_));
  OAI21X1  g09902(.A0(new_n10903_), .A1(new_n9526_), .B0(new_n10904_), .Y(new_n10905_));
  OR2X1    g09903(.A(new_n10896_), .B(new_n10905_), .Y(new_n10906_));
  AOI21X1  g09904(.A0(new_n10896_), .A1(new_n10905_), .B0(new_n10890_), .Y(new_n10907_));
  NAND3X1  g09905(.A(new_n10907_), .B(new_n10906_), .C(new_n10901_), .Y(new_n10908_));
  NAND2X1  g09906(.A(new_n10908_), .B(new_n10898_), .Y(new_n10909_));
  OR2X1    g09907(.A(new_n9493_), .B(new_n9487_), .Y(new_n10910_));
  AOI22X1  g09908(.A0(new_n10910_), .A1(new_n10879_), .B0(new_n9463_), .B1(new_n9450_), .Y(new_n10911_));
  NOR4X1   g09909(.A(new_n9493_), .B(new_n9487_), .C(new_n9480_), .D(new_n9475_), .Y(new_n10912_));
  AOI21X1  g09910(.A0(new_n9447_), .A1(new_n9446_), .B0(new_n9490_), .Y(new_n10913_));
  AOI21X1  g09911(.A0(new_n10913_), .A1(new_n9483_), .B0(new_n9491_), .Y(new_n10914_));
  AOI21X1  g09912(.A0(new_n9483_), .A1(new_n9482_), .B0(new_n9484_), .Y(new_n10915_));
  NOR2X1   g09913(.A(new_n10915_), .B(new_n10914_), .Y(new_n10916_));
  NAND3X1  g09914(.A(new_n9472_), .B(new_n9471_), .C(new_n9465_), .Y(new_n10917_));
  AOI21X1  g09915(.A0(new_n9471_), .A1(new_n9465_), .B0(new_n9472_), .Y(new_n10918_));
  AOI21X1  g09916(.A0(new_n10917_), .A1(new_n9473_), .B0(new_n10918_), .Y(new_n10919_));
  XOR2X1   g09917(.A(new_n10919_), .B(new_n10916_), .Y(new_n10920_));
  OAI21X1  g09918(.A0(new_n10912_), .A1(new_n10911_), .B0(new_n10920_), .Y(new_n10921_));
  AND2X1   g09919(.A(new_n5964_), .B(new_n6006_), .Y(new_n10922_));
  AOI21X1  g09920(.A0(new_n6007_), .A1(new_n5939_), .B0(new_n6005_), .Y(new_n10923_));
  OAI22X1  g09921(.A0(new_n9494_), .A1(new_n9481_), .B0(new_n10923_), .B1(new_n10922_), .Y(new_n10924_));
  OR4X1    g09922(.A(new_n9493_), .B(new_n9487_), .C(new_n9480_), .D(new_n9475_), .Y(new_n10925_));
  OR2X1    g09923(.A(new_n10915_), .B(new_n10914_), .Y(new_n10926_));
  NAND2X1  g09924(.A(new_n10919_), .B(new_n10926_), .Y(new_n10927_));
  OR2X1    g09925(.A(new_n10919_), .B(new_n10926_), .Y(new_n10928_));
  NAND4X1  g09926(.A(new_n10928_), .B(new_n10927_), .C(new_n10925_), .D(new_n10924_), .Y(new_n10929_));
  AND2X1   g09927(.A(new_n10929_), .B(new_n10921_), .Y(new_n10930_));
  XOR2X1   g09928(.A(new_n10930_), .B(new_n10909_), .Y(new_n10931_));
  XOR2X1   g09929(.A(new_n10931_), .B(new_n10887_), .Y(new_n10932_));
  XOR2X1   g09930(.A(new_n10932_), .B(new_n10878_), .Y(new_n10933_));
  XOR2X1   g09931(.A(new_n10933_), .B(new_n10826_), .Y(new_n10934_));
  OR2X1    g09932(.A(new_n9253_), .B(new_n7079_), .Y(new_n10935_));
  OAI21X1  g09933(.A0(new_n9266_), .A1(new_n7113_), .B0(new_n7196_), .Y(new_n10936_));
  OAI22X1  g09934(.A0(new_n9267_), .A1(new_n7196_), .B0(new_n10936_), .B1(new_n9269_), .Y(new_n10937_));
  OAI22X1  g09935(.A0(new_n9280_), .A1(new_n9269_), .B0(new_n9267_), .B1(new_n7130_), .Y(new_n10938_));
  MX2X1    g09936(.A(new_n10938_), .B(new_n10937_), .S0(new_n7195_), .Y(new_n10939_));
  OAI21X1  g09937(.A0(new_n9255_), .A1(new_n9249_), .B0(new_n10939_), .Y(new_n10940_));
  AND2X1   g09938(.A(new_n10940_), .B(new_n10935_), .Y(new_n10941_));
  XOR2X1   g09939(.A(new_n9350_), .B(new_n10941_), .Y(new_n10942_));
  OR2X1    g09940(.A(new_n6953_), .B(new_n6923_), .Y(new_n10943_));
  OAI21X1  g09941(.A0(new_n6954_), .A1(new_n6950_), .B0(new_n6824_), .Y(new_n10944_));
  AND2X1   g09942(.A(new_n10944_), .B(new_n10943_), .Y(new_n10945_));
  XOR2X1   g09943(.A(new_n9435_), .B(new_n10945_), .Y(new_n10946_));
  OAI22X1  g09944(.A0(new_n10946_), .A1(new_n10942_), .B0(new_n10810_), .B1(new_n10809_), .Y(new_n10947_));
  OR2X1    g09945(.A(new_n9436_), .B(new_n9351_), .Y(new_n10948_));
  AND2X1   g09946(.A(new_n10948_), .B(new_n10947_), .Y(new_n10949_));
  NOR2X1   g09947(.A(new_n9418_), .B(new_n9413_), .Y(new_n10950_));
  XOR2X1   g09948(.A(new_n9432_), .B(new_n10950_), .Y(new_n10951_));
  XOR2X1   g09949(.A(new_n10951_), .B(new_n9402_), .Y(new_n10952_));
  AOI22X1  g09950(.A0(new_n10952_), .A1(new_n9399_), .B0(new_n10944_), .B1(new_n10943_), .Y(new_n10953_));
  NOR2X1   g09951(.A(new_n10952_), .B(new_n9399_), .Y(new_n10954_));
  OR2X1    g09952(.A(new_n10954_), .B(new_n10953_), .Y(new_n10955_));
  OR2X1    g09953(.A(new_n9431_), .B(new_n9425_), .Y(new_n10956_));
  AOI22X1  g09954(.A0(new_n10956_), .A1(new_n9419_), .B0(new_n9401_), .B1(new_n9400_), .Y(new_n10957_));
  NOR4X1   g09955(.A(new_n9431_), .B(new_n9425_), .C(new_n9418_), .D(new_n9413_), .Y(new_n10958_));
  AOI21X1  g09956(.A0(new_n6927_), .A1(new_n6926_), .B0(new_n9428_), .Y(new_n10959_));
  AOI21X1  g09957(.A0(new_n10959_), .A1(new_n9421_), .B0(new_n9429_), .Y(new_n10960_));
  AOI21X1  g09958(.A0(new_n9421_), .A1(new_n9420_), .B0(new_n9422_), .Y(new_n10961_));
  NOR2X1   g09959(.A(new_n10961_), .B(new_n10960_), .Y(new_n10962_));
  NAND3X1  g09960(.A(new_n9410_), .B(new_n9409_), .C(new_n9403_), .Y(new_n10963_));
  AOI21X1  g09961(.A0(new_n9409_), .A1(new_n9403_), .B0(new_n9410_), .Y(new_n10964_));
  AOI21X1  g09962(.A0(new_n10963_), .A1(new_n9411_), .B0(new_n10964_), .Y(new_n10965_));
  XOR2X1   g09963(.A(new_n10965_), .B(new_n10962_), .Y(new_n10966_));
  OAI21X1  g09964(.A0(new_n10958_), .A1(new_n10957_), .B0(new_n10966_), .Y(new_n10967_));
  AND2X1   g09965(.A(new_n6919_), .B(new_n6941_), .Y(new_n10968_));
  AOI21X1  g09966(.A0(new_n6951_), .A1(new_n6894_), .B0(new_n6940_), .Y(new_n10969_));
  OAI22X1  g09967(.A0(new_n9432_), .A1(new_n10950_), .B0(new_n10969_), .B1(new_n10968_), .Y(new_n10970_));
  OR2X1    g09968(.A(new_n10961_), .B(new_n10960_), .Y(new_n10971_));
  OR2X1    g09969(.A(new_n10965_), .B(new_n10971_), .Y(new_n10972_));
  AOI21X1  g09970(.A0(new_n10965_), .A1(new_n10971_), .B0(new_n10958_), .Y(new_n10973_));
  NAND3X1  g09971(.A(new_n10973_), .B(new_n10972_), .C(new_n10970_), .Y(new_n10974_));
  NAND2X1  g09972(.A(new_n10974_), .B(new_n10967_), .Y(new_n10975_));
  OR2X1    g09973(.A(new_n9383_), .B(new_n9378_), .Y(new_n10976_));
  OR2X1    g09974(.A(new_n9396_), .B(new_n9390_), .Y(new_n10977_));
  AOI22X1  g09975(.A0(new_n10977_), .A1(new_n10976_), .B0(new_n9366_), .B1(new_n9355_), .Y(new_n10978_));
  NOR4X1   g09976(.A(new_n9396_), .B(new_n9390_), .C(new_n9383_), .D(new_n9378_), .Y(new_n10979_));
  AOI21X1  g09977(.A0(new_n6774_), .A1(new_n6772_), .B0(new_n9393_), .Y(new_n10980_));
  AOI21X1  g09978(.A0(new_n10980_), .A1(new_n9386_), .B0(new_n9394_), .Y(new_n10981_));
  AOI21X1  g09979(.A0(new_n9386_), .A1(new_n9385_), .B0(new_n9387_), .Y(new_n10982_));
  NOR2X1   g09980(.A(new_n10982_), .B(new_n10981_), .Y(new_n10983_));
  NAND3X1  g09981(.A(new_n9375_), .B(new_n9374_), .C(new_n9368_), .Y(new_n10984_));
  AOI21X1  g09982(.A0(new_n9374_), .A1(new_n9368_), .B0(new_n9375_), .Y(new_n10985_));
  AOI21X1  g09983(.A0(new_n10984_), .A1(new_n9376_), .B0(new_n10985_), .Y(new_n10986_));
  XOR2X1   g09984(.A(new_n10986_), .B(new_n10983_), .Y(new_n10987_));
  OAI21X1  g09985(.A0(new_n10979_), .A1(new_n10978_), .B0(new_n10987_), .Y(new_n10988_));
  AND2X1   g09986(.A(new_n6972_), .B(new_n6764_), .Y(new_n10989_));
  AOI21X1  g09987(.A0(new_n6974_), .A1(new_n6957_), .B0(new_n6820_), .Y(new_n10990_));
  OAI22X1  g09988(.A0(new_n9397_), .A1(new_n9384_), .B0(new_n10990_), .B1(new_n10989_), .Y(new_n10991_));
  OR4X1    g09989(.A(new_n9396_), .B(new_n9390_), .C(new_n9383_), .D(new_n9378_), .Y(new_n10992_));
  OR2X1    g09990(.A(new_n10982_), .B(new_n10981_), .Y(new_n10993_));
  NAND2X1  g09991(.A(new_n10986_), .B(new_n10993_), .Y(new_n10994_));
  OR2X1    g09992(.A(new_n10986_), .B(new_n10993_), .Y(new_n10995_));
  NAND4X1  g09993(.A(new_n10995_), .B(new_n10994_), .C(new_n10992_), .D(new_n10991_), .Y(new_n10996_));
  AND2X1   g09994(.A(new_n10996_), .B(new_n10988_), .Y(new_n10997_));
  XOR2X1   g09995(.A(new_n10997_), .B(new_n10975_), .Y(new_n10998_));
  XOR2X1   g09996(.A(new_n10998_), .B(new_n10955_), .Y(new_n10999_));
  OR2X1    g09997(.A(new_n9298_), .B(new_n9293_), .Y(new_n11000_));
  XOR2X1   g09998(.A(new_n9312_), .B(new_n11000_), .Y(new_n11001_));
  XOR2X1   g09999(.A(new_n11001_), .B(new_n9282_), .Y(new_n11002_));
  OAI22X1  g10000(.A0(new_n9349_), .A1(new_n11002_), .B0(new_n9261_), .B1(new_n9260_), .Y(new_n11003_));
  NOR2X1   g10001(.A(new_n9333_), .B(new_n9328_), .Y(new_n11004_));
  XOR2X1   g10002(.A(new_n9347_), .B(new_n11004_), .Y(new_n11005_));
  XOR2X1   g10003(.A(new_n11005_), .B(new_n9317_), .Y(new_n11006_));
  OR2X1    g10004(.A(new_n11006_), .B(new_n9314_), .Y(new_n11007_));
  AND2X1   g10005(.A(new_n11007_), .B(new_n11003_), .Y(new_n11008_));
  OR2X1    g10006(.A(new_n9346_), .B(new_n9340_), .Y(new_n11009_));
  AOI22X1  g10007(.A0(new_n11009_), .A1(new_n9334_), .B0(new_n9316_), .B1(new_n9315_), .Y(new_n11010_));
  NOR4X1   g10008(.A(new_n9346_), .B(new_n9340_), .C(new_n9333_), .D(new_n9328_), .Y(new_n11011_));
  AOI21X1  g10009(.A0(new_n7083_), .A1(new_n7082_), .B0(new_n9343_), .Y(new_n11012_));
  AOI21X1  g10010(.A0(new_n11012_), .A1(new_n9336_), .B0(new_n9344_), .Y(new_n11013_));
  AOI21X1  g10011(.A0(new_n9336_), .A1(new_n9335_), .B0(new_n9337_), .Y(new_n11014_));
  NOR2X1   g10012(.A(new_n11014_), .B(new_n11013_), .Y(new_n11015_));
  NAND3X1  g10013(.A(new_n9325_), .B(new_n9324_), .C(new_n9318_), .Y(new_n11016_));
  AOI21X1  g10014(.A0(new_n9324_), .A1(new_n9318_), .B0(new_n9325_), .Y(new_n11017_));
  AOI21X1  g10015(.A0(new_n11016_), .A1(new_n9326_), .B0(new_n11017_), .Y(new_n11018_));
  XOR2X1   g10016(.A(new_n11018_), .B(new_n11015_), .Y(new_n11019_));
  OAI21X1  g10017(.A0(new_n11011_), .A1(new_n11010_), .B0(new_n11019_), .Y(new_n11020_));
  AND2X1   g10018(.A(new_n7076_), .B(new_n7097_), .Y(new_n11021_));
  AOI21X1  g10019(.A0(new_n9250_), .A1(new_n7051_), .B0(new_n7096_), .Y(new_n11022_));
  OAI22X1  g10020(.A0(new_n9347_), .A1(new_n11004_), .B0(new_n11022_), .B1(new_n11021_), .Y(new_n11023_));
  OR2X1    g10021(.A(new_n11014_), .B(new_n11013_), .Y(new_n11024_));
  OR2X1    g10022(.A(new_n11018_), .B(new_n11024_), .Y(new_n11025_));
  AOI21X1  g10023(.A0(new_n11018_), .A1(new_n11024_), .B0(new_n11011_), .Y(new_n11026_));
  NAND3X1  g10024(.A(new_n11026_), .B(new_n11025_), .C(new_n11023_), .Y(new_n11027_));
  NAND2X1  g10025(.A(new_n11027_), .B(new_n11020_), .Y(new_n11028_));
  OR2X1    g10026(.A(new_n9311_), .B(new_n9305_), .Y(new_n11029_));
  AOI22X1  g10027(.A0(new_n11029_), .A1(new_n11000_), .B0(new_n9281_), .B1(new_n9268_), .Y(new_n11030_));
  NOR4X1   g10028(.A(new_n9311_), .B(new_n9305_), .C(new_n9298_), .D(new_n9293_), .Y(new_n11031_));
  AOI21X1  g10029(.A0(new_n9265_), .A1(new_n9264_), .B0(new_n9308_), .Y(new_n11032_));
  AOI21X1  g10030(.A0(new_n11032_), .A1(new_n9301_), .B0(new_n9309_), .Y(new_n11033_));
  AOI21X1  g10031(.A0(new_n9301_), .A1(new_n9300_), .B0(new_n9302_), .Y(new_n11034_));
  NOR2X1   g10032(.A(new_n11034_), .B(new_n11033_), .Y(new_n11035_));
  NAND3X1  g10033(.A(new_n9290_), .B(new_n9289_), .C(new_n9283_), .Y(new_n11036_));
  AOI21X1  g10034(.A0(new_n9289_), .A1(new_n9283_), .B0(new_n9290_), .Y(new_n11037_));
  AOI21X1  g10035(.A0(new_n11036_), .A1(new_n9291_), .B0(new_n11037_), .Y(new_n11038_));
  XOR2X1   g10036(.A(new_n11038_), .B(new_n11035_), .Y(new_n11039_));
  OAI21X1  g10037(.A0(new_n11031_), .A1(new_n11030_), .B0(new_n11039_), .Y(new_n11040_));
  AND2X1   g10038(.A(new_n7154_), .B(new_n7196_), .Y(new_n11041_));
  AOI21X1  g10039(.A0(new_n7197_), .A1(new_n7129_), .B0(new_n7195_), .Y(new_n11042_));
  OAI22X1  g10040(.A0(new_n9312_), .A1(new_n9299_), .B0(new_n11042_), .B1(new_n11041_), .Y(new_n11043_));
  OR4X1    g10041(.A(new_n9311_), .B(new_n9305_), .C(new_n9298_), .D(new_n9293_), .Y(new_n11044_));
  OR2X1    g10042(.A(new_n11034_), .B(new_n11033_), .Y(new_n11045_));
  NAND2X1  g10043(.A(new_n11038_), .B(new_n11045_), .Y(new_n11046_));
  OR2X1    g10044(.A(new_n11038_), .B(new_n11045_), .Y(new_n11047_));
  NAND4X1  g10045(.A(new_n11047_), .B(new_n11046_), .C(new_n11044_), .D(new_n11043_), .Y(new_n11048_));
  AND2X1   g10046(.A(new_n11048_), .B(new_n11040_), .Y(new_n11049_));
  XOR2X1   g10047(.A(new_n11049_), .B(new_n11028_), .Y(new_n11050_));
  XOR2X1   g10048(.A(new_n11050_), .B(new_n11008_), .Y(new_n11051_));
  XOR2X1   g10049(.A(new_n11051_), .B(new_n10999_), .Y(new_n11052_));
  XOR2X1   g10050(.A(new_n11052_), .B(new_n10949_), .Y(new_n11053_));
  XOR2X1   g10051(.A(new_n11053_), .B(new_n10934_), .Y(new_n11054_));
  XOR2X1   g10052(.A(new_n11054_), .B(new_n10819_), .Y(new_n11055_));
  XOR2X1   g10053(.A(new_n11055_), .B(new_n10806_), .Y(new_n11056_));
  XOR2X1   g10054(.A(new_n11056_), .B(new_n10561_), .Y(new_n11057_));
  NOR3X1   g10055(.A(new_n5607_), .B(new_n5614_), .C(new_n5611_), .Y(new_n11058_));
  OAI21X1  g10056(.A0(new_n11058_), .A1(new_n5618_), .B0(new_n5620_), .Y(new_n11059_));
  XOR2X1   g10057(.A(new_n9223_), .B(new_n11059_), .Y(new_n11060_));
  XOR2X1   g10058(.A(new_n11060_), .B(new_n9163_), .Y(new_n11061_));
  XOR2X1   g10059(.A(new_n11061_), .B(new_n9103_), .Y(new_n11062_));
  AOI22X1  g10060(.A0(new_n9231_), .A1(new_n11062_), .B0(new_n10543_), .B1(new_n10541_), .Y(new_n11063_));
  AOI21X1  g10061(.A0(new_n9100_), .A1(new_n8857_), .B0(new_n11062_), .Y(new_n11064_));
  AND2X1   g10062(.A(new_n11064_), .B(new_n9101_), .Y(new_n11065_));
  OR2X1    g10063(.A(new_n11065_), .B(new_n11063_), .Y(new_n11066_));
  XOR2X1   g10064(.A(new_n9018_), .B(new_n8860_), .Y(new_n11067_));
  OAI22X1  g10065(.A0(new_n11067_), .A1(new_n9085_), .B0(new_n9229_), .B1(new_n9228_), .Y(new_n11068_));
  AND2X1   g10066(.A(new_n9018_), .B(new_n8860_), .Y(new_n11069_));
  OAI21X1  g10067(.A0(new_n9018_), .A1(new_n8860_), .B0(new_n9085_), .Y(new_n11070_));
  OR2X1    g10068(.A(new_n11070_), .B(new_n11069_), .Y(new_n11071_));
  AND2X1   g10069(.A(new_n11071_), .B(new_n11068_), .Y(new_n11072_));
  OAI22X1  g10070(.A0(new_n9017_), .A1(new_n8931_), .B0(new_n8859_), .B1(new_n8858_), .Y(new_n11073_));
  NAND2X1  g10071(.A(new_n9017_), .B(new_n8931_), .Y(new_n11074_));
  AND2X1   g10072(.A(new_n11074_), .B(new_n11073_), .Y(new_n11075_));
  AND2X1   g10073(.A(new_n4869_), .B(new_n4828_), .Y(new_n11076_));
  AOI21X1  g10074(.A0(new_n4870_), .A1(new_n4866_), .B0(new_n4656_), .Y(new_n11077_));
  OR2X1    g10075(.A(new_n8964_), .B(new_n8958_), .Y(new_n11078_));
  XOR2X1   g10076(.A(new_n8978_), .B(new_n11078_), .Y(new_n11079_));
  XOR2X1   g10077(.A(new_n11079_), .B(new_n8947_), .Y(new_n11080_));
  OAI22X1  g10078(.A0(new_n9015_), .A1(new_n11080_), .B0(new_n11077_), .B1(new_n11076_), .Y(new_n11081_));
  NOR2X1   g10079(.A(new_n8999_), .B(new_n8994_), .Y(new_n11082_));
  XOR2X1   g10080(.A(new_n9013_), .B(new_n11082_), .Y(new_n11083_));
  XOR2X1   g10081(.A(new_n11083_), .B(new_n8983_), .Y(new_n11084_));
  OR2X1    g10082(.A(new_n11084_), .B(new_n8980_), .Y(new_n11085_));
  AND2X1   g10083(.A(new_n11085_), .B(new_n11081_), .Y(new_n11086_));
  OR2X1    g10084(.A(new_n9012_), .B(new_n9006_), .Y(new_n11087_));
  AOI22X1  g10085(.A0(new_n11087_), .A1(new_n9000_), .B0(new_n8982_), .B1(new_n8981_), .Y(new_n11088_));
  NOR4X1   g10086(.A(new_n9012_), .B(new_n9006_), .C(new_n8999_), .D(new_n8994_), .Y(new_n11089_));
  NAND3X1  g10087(.A(new_n9003_), .B(new_n9002_), .C(new_n9001_), .Y(new_n11090_));
  AOI21X1  g10088(.A0(new_n9002_), .A1(new_n9001_), .B0(new_n9003_), .Y(new_n11091_));
  AOI21X1  g10089(.A0(new_n11090_), .A1(new_n9004_), .B0(new_n11091_), .Y(new_n11092_));
  NAND3X1  g10090(.A(new_n8991_), .B(new_n8990_), .C(new_n8984_), .Y(new_n11093_));
  AOI21X1  g10091(.A0(new_n8990_), .A1(new_n8984_), .B0(new_n8991_), .Y(new_n11094_));
  AOI21X1  g10092(.A0(new_n11093_), .A1(new_n8992_), .B0(new_n11094_), .Y(new_n11095_));
  XOR2X1   g10093(.A(new_n11095_), .B(new_n11092_), .Y(new_n11096_));
  OAI21X1  g10094(.A0(new_n11089_), .A1(new_n11088_), .B0(new_n11096_), .Y(new_n11097_));
  AND2X1   g10095(.A(new_n4834_), .B(new_n4805_), .Y(new_n11098_));
  AOI21X1  g10096(.A0(new_n4840_), .A1(new_n4829_), .B0(new_n4733_), .Y(new_n11099_));
  OAI22X1  g10097(.A0(new_n9013_), .A1(new_n11082_), .B0(new_n11099_), .B1(new_n11098_), .Y(new_n11100_));
  AND2X1   g10098(.A(new_n4815_), .B(new_n4810_), .Y(new_n11101_));
  NOR3X1   g10099(.A(new_n9009_), .B(new_n9007_), .C(new_n11101_), .Y(new_n11102_));
  OAI21X1  g10100(.A0(new_n9007_), .A1(new_n11101_), .B0(new_n9009_), .Y(new_n11103_));
  OAI21X1  g10101(.A0(new_n11102_), .A1(new_n9010_), .B0(new_n11103_), .Y(new_n11104_));
  OR2X1    g10102(.A(new_n11095_), .B(new_n11104_), .Y(new_n11105_));
  AOI21X1  g10103(.A0(new_n11095_), .A1(new_n11104_), .B0(new_n11089_), .Y(new_n11106_));
  NAND3X1  g10104(.A(new_n11106_), .B(new_n11105_), .C(new_n11100_), .Y(new_n11107_));
  NAND2X1  g10105(.A(new_n11107_), .B(new_n11097_), .Y(new_n11108_));
  OR2X1    g10106(.A(new_n8977_), .B(new_n8971_), .Y(new_n11109_));
  AOI22X1  g10107(.A0(new_n11109_), .A1(new_n11078_), .B0(new_n8946_), .B1(new_n8935_), .Y(new_n11110_));
  NOR4X1   g10108(.A(new_n8977_), .B(new_n8971_), .C(new_n8964_), .D(new_n8958_), .Y(new_n11111_));
  AND2X1   g10109(.A(new_n4900_), .B(new_n4899_), .Y(new_n11112_));
  NOR3X1   g10110(.A(new_n8974_), .B(new_n8972_), .C(new_n11112_), .Y(new_n11113_));
  OAI21X1  g10111(.A0(new_n8972_), .A1(new_n11112_), .B0(new_n8974_), .Y(new_n11114_));
  OAI21X1  g10112(.A0(new_n11113_), .A1(new_n8975_), .B0(new_n11114_), .Y(new_n11115_));
  NAND3X1  g10113(.A(new_n8955_), .B(new_n8954_), .C(new_n8948_), .Y(new_n11116_));
  AOI21X1  g10114(.A0(new_n8954_), .A1(new_n8948_), .B0(new_n8955_), .Y(new_n11117_));
  AOI21X1  g10115(.A0(new_n11116_), .A1(new_n8956_), .B0(new_n11117_), .Y(new_n11118_));
  AND2X1   g10116(.A(new_n11118_), .B(new_n11115_), .Y(new_n11119_));
  NOR2X1   g10117(.A(new_n11118_), .B(new_n11115_), .Y(new_n11120_));
  OAI22X1  g10118(.A0(new_n11120_), .A1(new_n11119_), .B0(new_n11111_), .B1(new_n11110_), .Y(new_n11121_));
  AND2X1   g10119(.A(new_n4611_), .B(new_n4653_), .Y(new_n11122_));
  AOI21X1  g10120(.A0(new_n4654_), .A1(new_n4548_), .B0(new_n4652_), .Y(new_n11123_));
  OAI22X1  g10121(.A0(new_n8978_), .A1(new_n8965_), .B0(new_n11123_), .B1(new_n11122_), .Y(new_n11124_));
  OR4X1    g10122(.A(new_n8977_), .B(new_n8971_), .C(new_n8964_), .D(new_n8958_), .Y(new_n11125_));
  NAND2X1  g10123(.A(new_n11118_), .B(new_n11115_), .Y(new_n11126_));
  OR2X1    g10124(.A(new_n11118_), .B(new_n11115_), .Y(new_n11127_));
  NAND4X1  g10125(.A(new_n11127_), .B(new_n11126_), .C(new_n11125_), .D(new_n11124_), .Y(new_n11128_));
  AND2X1   g10126(.A(new_n11128_), .B(new_n11121_), .Y(new_n11129_));
  XOR2X1   g10127(.A(new_n11129_), .B(new_n11108_), .Y(new_n11130_));
  XOR2X1   g10128(.A(new_n11130_), .B(new_n11086_), .Y(new_n11131_));
  NOR2X1   g10129(.A(new_n8913_), .B(new_n8907_), .Y(new_n11132_));
  XOR2X1   g10130(.A(new_n8927_), .B(new_n11132_), .Y(new_n11133_));
  XOR2X1   g10131(.A(new_n11133_), .B(new_n8898_), .Y(new_n11134_));
  AOI22X1  g10132(.A0(new_n11134_), .A1(new_n8895_), .B0(new_n8862_), .B1(new_n8861_), .Y(new_n11135_));
  NOR2X1   g10133(.A(new_n8928_), .B(new_n8898_), .Y(new_n11136_));
  AND2X1   g10134(.A(new_n8928_), .B(new_n8898_), .Y(new_n11137_));
  NOR3X1   g10135(.A(new_n11137_), .B(new_n11136_), .C(new_n8895_), .Y(new_n11138_));
  OR2X1    g10136(.A(new_n11138_), .B(new_n11135_), .Y(new_n11139_));
  AND2X1   g10137(.A(new_n8876_), .B(new_n8871_), .Y(new_n11140_));
  AOI21X1  g10138(.A0(new_n8866_), .A1(new_n8864_), .B0(new_n11140_), .Y(new_n11141_));
  NAND3X1  g10139(.A(new_n11140_), .B(new_n8866_), .C(new_n8864_), .Y(new_n11142_));
  AOI21X1  g10140(.A0(new_n11142_), .A1(new_n8878_), .B0(new_n11141_), .Y(new_n11143_));
  AOI21X1  g10141(.A0(new_n8873_), .A1(new_n8872_), .B0(new_n8870_), .Y(new_n11144_));
  INVX1    g10142(.A(new_n11144_), .Y(new_n11145_));
  OR2X1    g10143(.A(new_n8881_), .B(new_n8880_), .Y(new_n11146_));
  NOR3X1   g10144(.A(new_n11146_), .B(new_n8891_), .C(new_n8888_), .Y(new_n11147_));
  OAI21X1  g10145(.A0(new_n11147_), .A1(new_n8883_), .B0(new_n11145_), .Y(new_n11148_));
  OAI22X1  g10146(.A0(new_n11148_), .A1(new_n11141_), .B0(new_n11145_), .B1(new_n11143_), .Y(new_n11149_));
  OAI22X1  g10147(.A0(new_n8927_), .A1(new_n11132_), .B0(new_n8897_), .B1(new_n8896_), .Y(new_n11150_));
  OR4X1    g10148(.A(new_n8926_), .B(new_n8920_), .C(new_n8913_), .D(new_n8907_), .Y(new_n11151_));
  AND2X1   g10149(.A(new_n4427_), .B(new_n4426_), .Y(new_n11152_));
  NOR3X1   g10150(.A(new_n8923_), .B(new_n8921_), .C(new_n11152_), .Y(new_n11153_));
  OAI21X1  g10151(.A0(new_n8921_), .A1(new_n11152_), .B0(new_n8923_), .Y(new_n11154_));
  OAI21X1  g10152(.A0(new_n11153_), .A1(new_n8924_), .B0(new_n11154_), .Y(new_n11155_));
  NAND3X1  g10153(.A(new_n8904_), .B(new_n8903_), .C(new_n8901_), .Y(new_n11156_));
  AOI21X1  g10154(.A0(new_n8903_), .A1(new_n8901_), .B0(new_n8904_), .Y(new_n11157_));
  AOI21X1  g10155(.A0(new_n11156_), .A1(new_n8905_), .B0(new_n11157_), .Y(new_n11158_));
  XOR2X1   g10156(.A(new_n11158_), .B(new_n11155_), .Y(new_n11159_));
  AOI21X1  g10157(.A0(new_n11151_), .A1(new_n11150_), .B0(new_n11159_), .Y(new_n11160_));
  OR2X1    g10158(.A(new_n11158_), .B(new_n11155_), .Y(new_n11161_));
  NOR4X1   g10159(.A(new_n8926_), .B(new_n8920_), .C(new_n8913_), .D(new_n8907_), .Y(new_n11162_));
  AOI21X1  g10160(.A0(new_n11158_), .A1(new_n11155_), .B0(new_n11162_), .Y(new_n11163_));
  AND2X1   g10161(.A(new_n11163_), .B(new_n11161_), .Y(new_n11164_));
  AOI21X1  g10162(.A0(new_n11164_), .A1(new_n11150_), .B0(new_n11160_), .Y(new_n11165_));
  XOR2X1   g10163(.A(new_n11165_), .B(new_n11149_), .Y(new_n11166_));
  XOR2X1   g10164(.A(new_n11166_), .B(new_n11139_), .Y(new_n11167_));
  XOR2X1   g10165(.A(new_n11167_), .B(new_n11131_), .Y(new_n11168_));
  NAND2X1  g10166(.A(new_n11168_), .B(new_n11075_), .Y(new_n11169_));
  OR2X1    g10167(.A(new_n11077_), .B(new_n11076_), .Y(new_n11170_));
  XOR2X1   g10168(.A(new_n9016_), .B(new_n11170_), .Y(new_n11171_));
  AOI22X1  g10169(.A0(new_n11171_), .A1(new_n9096_), .B0(new_n9087_), .B1(new_n9086_), .Y(new_n11172_));
  AND2X1   g10170(.A(new_n9017_), .B(new_n8931_), .Y(new_n11173_));
  OR2X1    g10171(.A(new_n11173_), .B(new_n11172_), .Y(new_n11174_));
  XOR2X1   g10172(.A(new_n11168_), .B(new_n11174_), .Y(new_n11175_));
  OR2X1    g10173(.A(new_n4183_), .B(new_n4179_), .Y(new_n11176_));
  AOI22X1  g10174(.A0(new_n9083_), .A1(new_n9050_), .B0(new_n11176_), .B1(new_n9020_), .Y(new_n11177_));
  NOR2X1   g10175(.A(new_n9083_), .B(new_n9050_), .Y(new_n11178_));
  NOR2X1   g10176(.A(new_n11178_), .B(new_n11177_), .Y(new_n11179_));
  OR2X1    g10177(.A(new_n9065_), .B(new_n9060_), .Y(new_n11180_));
  OR2X1    g10178(.A(new_n9080_), .B(new_n9075_), .Y(new_n11181_));
  AOI21X1  g10179(.A0(new_n11181_), .A1(new_n11180_), .B0(new_n9052_), .Y(new_n11182_));
  NOR4X1   g10180(.A(new_n9080_), .B(new_n9075_), .C(new_n9065_), .D(new_n9060_), .Y(new_n11183_));
  AOI21X1  g10181(.A0(new_n3987_), .A1(new_n3984_), .B0(new_n9071_), .Y(new_n11184_));
  OAI21X1  g10182(.A0(new_n9067_), .A1(new_n3947_), .B0(new_n11184_), .Y(new_n11185_));
  AND2X1   g10183(.A(new_n11185_), .B(new_n9073_), .Y(new_n11186_));
  AND2X1   g10184(.A(new_n9071_), .B(new_n9070_), .Y(new_n11187_));
  OR2X1    g10185(.A(new_n11187_), .B(new_n11186_), .Y(new_n11188_));
  NAND3X1  g10186(.A(new_n9055_), .B(new_n9053_), .C(new_n3917_), .Y(new_n11189_));
  AOI21X1  g10187(.A0(new_n9053_), .A1(new_n3917_), .B0(new_n9055_), .Y(new_n11190_));
  AOI21X1  g10188(.A0(new_n11189_), .A1(new_n9058_), .B0(new_n11190_), .Y(new_n11191_));
  AND2X1   g10189(.A(new_n11191_), .B(new_n11188_), .Y(new_n11192_));
  NOR2X1   g10190(.A(new_n11191_), .B(new_n11188_), .Y(new_n11193_));
  OAI22X1  g10191(.A0(new_n11193_), .A1(new_n11192_), .B0(new_n11183_), .B1(new_n11182_), .Y(new_n11194_));
  AND2X1   g10192(.A(new_n4006_), .B(new_n3919_), .Y(new_n11195_));
  OAI22X1  g10193(.A0(new_n9081_), .A1(new_n9066_), .B0(new_n11195_), .B1(new_n9051_), .Y(new_n11196_));
  OR4X1    g10194(.A(new_n9080_), .B(new_n9075_), .C(new_n9065_), .D(new_n9060_), .Y(new_n11197_));
  NAND2X1  g10195(.A(new_n11191_), .B(new_n11188_), .Y(new_n11198_));
  OR2X1    g10196(.A(new_n11191_), .B(new_n11188_), .Y(new_n11199_));
  NAND4X1  g10197(.A(new_n11199_), .B(new_n11198_), .C(new_n11197_), .D(new_n11196_), .Y(new_n11200_));
  NAND2X1  g10198(.A(new_n11200_), .B(new_n11194_), .Y(new_n11201_));
  NOR2X1   g10199(.A(new_n9048_), .B(new_n9036_), .Y(new_n11202_));
  AND2X1   g10200(.A(new_n9030_), .B(new_n9025_), .Y(new_n11203_));
  AND2X1   g10201(.A(new_n9042_), .B(new_n9038_), .Y(new_n11204_));
  OR4X1    g10202(.A(new_n9047_), .B(new_n11204_), .C(new_n9035_), .D(new_n11203_), .Y(new_n11205_));
  OAI21X1  g10203(.A0(new_n11202_), .A1(new_n9023_), .B0(new_n11205_), .Y(new_n11206_));
  OAI21X1  g10204(.A0(new_n4127_), .A1(new_n4126_), .B0(new_n9044_), .Y(new_n11207_));
  OAI21X1  g10205(.A0(new_n11207_), .A1(new_n9037_), .B0(new_n9041_), .Y(new_n11208_));
  OAI21X1  g10206(.A0(new_n9037_), .A1(new_n4128_), .B0(new_n9040_), .Y(new_n11209_));
  AND2X1   g10207(.A(new_n11209_), .B(new_n11208_), .Y(new_n11210_));
  OAI21X1  g10208(.A0(new_n4168_), .A1(new_n4163_), .B0(new_n9032_), .Y(new_n11211_));
  OAI21X1  g10209(.A0(new_n11211_), .A1(new_n9024_), .B0(new_n9029_), .Y(new_n11212_));
  OAI21X1  g10210(.A0(new_n9024_), .A1(new_n4169_), .B0(new_n9027_), .Y(new_n11213_));
  AND2X1   g10211(.A(new_n11213_), .B(new_n11212_), .Y(new_n11214_));
  XOR2X1   g10212(.A(new_n11214_), .B(new_n11210_), .Y(new_n11215_));
  NAND2X1  g10213(.A(new_n11215_), .B(new_n11206_), .Y(new_n11216_));
  NOR2X1   g10214(.A(new_n11202_), .B(new_n9023_), .Y(new_n11217_));
  NOR4X1   g10215(.A(new_n9047_), .B(new_n11204_), .C(new_n9035_), .D(new_n11203_), .Y(new_n11218_));
  NAND2X1  g10216(.A(new_n11209_), .B(new_n11208_), .Y(new_n11219_));
  AND2X1   g10217(.A(new_n11214_), .B(new_n11219_), .Y(new_n11220_));
  NOR2X1   g10218(.A(new_n11214_), .B(new_n11219_), .Y(new_n11221_));
  OR4X1    g10219(.A(new_n11221_), .B(new_n11220_), .C(new_n11218_), .D(new_n11217_), .Y(new_n11222_));
  AND2X1   g10220(.A(new_n11222_), .B(new_n11216_), .Y(new_n11223_));
  XOR2X1   g10221(.A(new_n11223_), .B(new_n11201_), .Y(new_n11224_));
  XOR2X1   g10222(.A(new_n11224_), .B(new_n11179_), .Y(new_n11225_));
  AOI22X1  g10223(.A0(new_n11084_), .A1(new_n8980_), .B0(new_n8933_), .B1(new_n8932_), .Y(new_n11226_));
  NOR2X1   g10224(.A(new_n11084_), .B(new_n8980_), .Y(new_n11227_));
  OR2X1    g10225(.A(new_n11227_), .B(new_n11226_), .Y(new_n11228_));
  XOR2X1   g10226(.A(new_n11130_), .B(new_n11228_), .Y(new_n11229_));
  XOR2X1   g10227(.A(new_n11167_), .B(new_n11229_), .Y(new_n11230_));
  AOI21X1  g10228(.A0(new_n11230_), .A1(new_n11174_), .B0(new_n11225_), .Y(new_n11231_));
  AOI22X1  g10229(.A0(new_n11231_), .A1(new_n11169_), .B0(new_n11225_), .B1(new_n11175_), .Y(new_n11232_));
  AND2X1   g10230(.A(new_n11232_), .B(new_n11072_), .Y(new_n11233_));
  XOR2X1   g10231(.A(new_n11232_), .B(new_n11072_), .Y(new_n11234_));
  NAND2X1  g10232(.A(new_n9224_), .B(new_n9163_), .Y(new_n11235_));
  AND2X1   g10233(.A(new_n11235_), .B(new_n9103_), .Y(new_n11236_));
  NOR2X1   g10234(.A(new_n9224_), .B(new_n9163_), .Y(new_n11237_));
  OR2X1    g10235(.A(new_n11237_), .B(new_n11236_), .Y(new_n11238_));
  NAND2X1  g10236(.A(new_n9222_), .B(new_n9194_), .Y(new_n11239_));
  AND2X1   g10237(.A(new_n11239_), .B(new_n11059_), .Y(new_n11240_));
  NOR2X1   g10238(.A(new_n9222_), .B(new_n9194_), .Y(new_n11241_));
  OR2X1    g10239(.A(new_n11241_), .B(new_n11240_), .Y(new_n11242_));
  OAI21X1  g10240(.A0(new_n5603_), .A1(new_n5552_), .B0(new_n5613_), .Y(new_n11243_));
  OR2X1    g10241(.A(new_n9220_), .B(new_n9208_), .Y(new_n11244_));
  AND2X1   g10242(.A(new_n9202_), .B(new_n9197_), .Y(new_n11245_));
  AND2X1   g10243(.A(new_n9214_), .B(new_n9210_), .Y(new_n11246_));
  NOR4X1   g10244(.A(new_n9219_), .B(new_n11246_), .C(new_n9207_), .D(new_n11245_), .Y(new_n11247_));
  AOI21X1  g10245(.A0(new_n11244_), .A1(new_n11243_), .B0(new_n11247_), .Y(new_n11248_));
  OAI21X1  g10246(.A0(new_n5584_), .A1(new_n5579_), .B0(new_n9216_), .Y(new_n11249_));
  OAI21X1  g10247(.A0(new_n11249_), .A1(new_n9209_), .B0(new_n9213_), .Y(new_n11250_));
  OAI21X1  g10248(.A0(new_n9209_), .A1(new_n5597_), .B0(new_n9212_), .Y(new_n11251_));
  NAND2X1  g10249(.A(new_n11251_), .B(new_n11250_), .Y(new_n11252_));
  OAI21X1  g10250(.A0(new_n5549_), .A1(new_n5547_), .B0(new_n9204_), .Y(new_n11253_));
  OR2X1    g10251(.A(new_n11253_), .B(new_n9196_), .Y(new_n11254_));
  AOI22X1  g10252(.A0(new_n11254_), .A1(new_n9201_), .B0(new_n9199_), .B1(new_n9197_), .Y(new_n11255_));
  XOR2X1   g10253(.A(new_n11255_), .B(new_n11252_), .Y(new_n11256_));
  OR2X1    g10254(.A(new_n11256_), .B(new_n11248_), .Y(new_n11257_));
  NAND2X1  g10255(.A(new_n11244_), .B(new_n11243_), .Y(new_n11258_));
  OR4X1    g10256(.A(new_n9219_), .B(new_n11246_), .C(new_n9207_), .D(new_n11245_), .Y(new_n11259_));
  NAND2X1  g10257(.A(new_n11255_), .B(new_n11252_), .Y(new_n11260_));
  OR2X1    g10258(.A(new_n11255_), .B(new_n11252_), .Y(new_n11261_));
  NAND4X1  g10259(.A(new_n11261_), .B(new_n11260_), .C(new_n11259_), .D(new_n11258_), .Y(new_n11262_));
  NAND2X1  g10260(.A(new_n11262_), .B(new_n11257_), .Y(new_n11263_));
  NOR2X1   g10261(.A(new_n9192_), .B(new_n9180_), .Y(new_n11264_));
  AND2X1   g10262(.A(new_n9174_), .B(new_n9169_), .Y(new_n11265_));
  AND2X1   g10263(.A(new_n9186_), .B(new_n9182_), .Y(new_n11266_));
  OR4X1    g10264(.A(new_n9191_), .B(new_n11266_), .C(new_n9179_), .D(new_n11265_), .Y(new_n11267_));
  OAI21X1  g10265(.A0(new_n11264_), .A1(new_n9167_), .B0(new_n11267_), .Y(new_n11268_));
  OAI21X1  g10266(.A0(new_n5472_), .A1(new_n5471_), .B0(new_n9188_), .Y(new_n11269_));
  OAI21X1  g10267(.A0(new_n11269_), .A1(new_n9181_), .B0(new_n9185_), .Y(new_n11270_));
  OAI21X1  g10268(.A0(new_n9181_), .A1(new_n5473_), .B0(new_n9184_), .Y(new_n11271_));
  AND2X1   g10269(.A(new_n11271_), .B(new_n11270_), .Y(new_n11272_));
  OAI21X1  g10270(.A0(new_n5509_), .A1(new_n5507_), .B0(new_n9176_), .Y(new_n11273_));
  OR2X1    g10271(.A(new_n11273_), .B(new_n9168_), .Y(new_n11274_));
  AOI22X1  g10272(.A0(new_n11274_), .A1(new_n9173_), .B0(new_n9171_), .B1(new_n9169_), .Y(new_n11275_));
  XOR2X1   g10273(.A(new_n11275_), .B(new_n11272_), .Y(new_n11276_));
  NAND2X1  g10274(.A(new_n11276_), .B(new_n11268_), .Y(new_n11277_));
  OR2X1    g10275(.A(new_n11264_), .B(new_n9167_), .Y(new_n11278_));
  NAND2X1  g10276(.A(new_n11271_), .B(new_n11270_), .Y(new_n11279_));
  NAND2X1  g10277(.A(new_n11275_), .B(new_n11279_), .Y(new_n11280_));
  OR2X1    g10278(.A(new_n11275_), .B(new_n11279_), .Y(new_n11281_));
  NAND4X1  g10279(.A(new_n11281_), .B(new_n11280_), .C(new_n11267_), .D(new_n11278_), .Y(new_n11282_));
  AND2X1   g10280(.A(new_n11282_), .B(new_n11277_), .Y(new_n11283_));
  XOR2X1   g10281(.A(new_n11283_), .B(new_n11263_), .Y(new_n11284_));
  XOR2X1   g10282(.A(new_n11284_), .B(new_n11242_), .Y(new_n11285_));
  OAI21X1  g10283(.A0(new_n5432_), .A1(new_n5632_), .B0(new_n5634_), .Y(new_n11286_));
  NAND2X1  g10284(.A(new_n9161_), .B(new_n9133_), .Y(new_n11287_));
  NOR2X1   g10285(.A(new_n9161_), .B(new_n9133_), .Y(new_n11288_));
  AOI21X1  g10286(.A0(new_n11287_), .A1(new_n11286_), .B0(new_n11288_), .Y(new_n11289_));
  OAI21X1  g10287(.A0(new_n5332_), .A1(new_n5281_), .B0(new_n5342_), .Y(new_n11290_));
  OR2X1    g10288(.A(new_n9159_), .B(new_n9147_), .Y(new_n11291_));
  AND2X1   g10289(.A(new_n9141_), .B(new_n9136_), .Y(new_n11292_));
  AND2X1   g10290(.A(new_n9153_), .B(new_n9149_), .Y(new_n11293_));
  NOR4X1   g10291(.A(new_n9158_), .B(new_n11293_), .C(new_n9146_), .D(new_n11292_), .Y(new_n11294_));
  AOI21X1  g10292(.A0(new_n11291_), .A1(new_n11290_), .B0(new_n11294_), .Y(new_n11295_));
  OAI21X1  g10293(.A0(new_n5313_), .A1(new_n5308_), .B0(new_n9155_), .Y(new_n11296_));
  OAI21X1  g10294(.A0(new_n11296_), .A1(new_n9148_), .B0(new_n9152_), .Y(new_n11297_));
  OAI21X1  g10295(.A0(new_n9148_), .A1(new_n5326_), .B0(new_n9151_), .Y(new_n11298_));
  NAND2X1  g10296(.A(new_n11298_), .B(new_n11297_), .Y(new_n11299_));
  OAI21X1  g10297(.A0(new_n5278_), .A1(new_n5276_), .B0(new_n9143_), .Y(new_n11300_));
  OR2X1    g10298(.A(new_n11300_), .B(new_n9135_), .Y(new_n11301_));
  AOI22X1  g10299(.A0(new_n11301_), .A1(new_n9140_), .B0(new_n9138_), .B1(new_n9136_), .Y(new_n11302_));
  XOR2X1   g10300(.A(new_n11302_), .B(new_n11299_), .Y(new_n11303_));
  OR2X1    g10301(.A(new_n11303_), .B(new_n11295_), .Y(new_n11304_));
  NAND2X1  g10302(.A(new_n11291_), .B(new_n11290_), .Y(new_n11305_));
  OR4X1    g10303(.A(new_n9158_), .B(new_n11293_), .C(new_n9146_), .D(new_n11292_), .Y(new_n11306_));
  NAND2X1  g10304(.A(new_n11302_), .B(new_n11299_), .Y(new_n11307_));
  OR2X1    g10305(.A(new_n11302_), .B(new_n11299_), .Y(new_n11308_));
  NAND4X1  g10306(.A(new_n11308_), .B(new_n11307_), .C(new_n11306_), .D(new_n11305_), .Y(new_n11309_));
  NAND2X1  g10307(.A(new_n11309_), .B(new_n11304_), .Y(new_n11310_));
  NOR2X1   g10308(.A(new_n9131_), .B(new_n9119_), .Y(new_n11311_));
  AND2X1   g10309(.A(new_n9113_), .B(new_n9108_), .Y(new_n11312_));
  AND2X1   g10310(.A(new_n9125_), .B(new_n9121_), .Y(new_n11313_));
  OR4X1    g10311(.A(new_n9130_), .B(new_n11313_), .C(new_n9118_), .D(new_n11312_), .Y(new_n11314_));
  OAI21X1  g10312(.A0(new_n11311_), .A1(new_n9106_), .B0(new_n11314_), .Y(new_n11315_));
  OAI21X1  g10313(.A0(new_n5383_), .A1(new_n5382_), .B0(new_n9127_), .Y(new_n11316_));
  OAI21X1  g10314(.A0(new_n11316_), .A1(new_n9120_), .B0(new_n9124_), .Y(new_n11317_));
  OAI21X1  g10315(.A0(new_n9120_), .A1(new_n5384_), .B0(new_n9123_), .Y(new_n11318_));
  AND2X1   g10316(.A(new_n11318_), .B(new_n11317_), .Y(new_n11319_));
  OAI21X1  g10317(.A0(new_n5420_), .A1(new_n5418_), .B0(new_n9115_), .Y(new_n11320_));
  OR2X1    g10318(.A(new_n11320_), .B(new_n9107_), .Y(new_n11321_));
  AOI22X1  g10319(.A0(new_n11321_), .A1(new_n9112_), .B0(new_n9110_), .B1(new_n9108_), .Y(new_n11322_));
  XOR2X1   g10320(.A(new_n11322_), .B(new_n11319_), .Y(new_n11323_));
  NAND2X1  g10321(.A(new_n11323_), .B(new_n11315_), .Y(new_n11324_));
  OR2X1    g10322(.A(new_n11311_), .B(new_n9106_), .Y(new_n11325_));
  NAND2X1  g10323(.A(new_n11318_), .B(new_n11317_), .Y(new_n11326_));
  NAND2X1  g10324(.A(new_n11322_), .B(new_n11326_), .Y(new_n11327_));
  OR2X1    g10325(.A(new_n11322_), .B(new_n11326_), .Y(new_n11328_));
  NAND4X1  g10326(.A(new_n11328_), .B(new_n11327_), .C(new_n11314_), .D(new_n11325_), .Y(new_n11329_));
  AND2X1   g10327(.A(new_n11329_), .B(new_n11324_), .Y(new_n11330_));
  XOR2X1   g10328(.A(new_n11330_), .B(new_n11310_), .Y(new_n11331_));
  XOR2X1   g10329(.A(new_n11331_), .B(new_n11289_), .Y(new_n11332_));
  XOR2X1   g10330(.A(new_n11332_), .B(new_n11285_), .Y(new_n11333_));
  XOR2X1   g10331(.A(new_n11333_), .B(new_n11238_), .Y(new_n11334_));
  OAI21X1  g10332(.A0(new_n11232_), .A1(new_n11072_), .B0(new_n11334_), .Y(new_n11335_));
  OAI22X1  g10333(.A0(new_n11335_), .A1(new_n11233_), .B0(new_n11334_), .B1(new_n11234_), .Y(new_n11336_));
  XOR2X1   g10334(.A(new_n11336_), .B(new_n11066_), .Y(new_n11337_));
  XOR2X1   g10335(.A(new_n11337_), .B(new_n11057_), .Y(new_n11338_));
  AND2X1   g10336(.A(new_n11338_), .B(new_n10557_), .Y(new_n11339_));
  NOR2X1   g10337(.A(new_n10005_), .B(new_n10545_), .Y(new_n11340_));
  NAND2X1  g10338(.A(new_n10005_), .B(new_n10545_), .Y(new_n11341_));
  OAI21X1  g10339(.A0(new_n11340_), .A1(new_n10549_), .B0(new_n11341_), .Y(new_n11342_));
  XOR2X1   g10340(.A(new_n11338_), .B(new_n11342_), .Y(new_n11343_));
  AOI22X1  g10341(.A0(new_n10537_), .A1(new_n10270_), .B0(new_n10009_), .B1(new_n3846_), .Y(new_n11344_));
  NOR2X1   g10342(.A(new_n10537_), .B(new_n10270_), .Y(new_n11345_));
  OR2X1    g10343(.A(new_n11345_), .B(new_n11344_), .Y(new_n11346_));
  AOI21X1  g10344(.A0(new_n10535_), .A1(new_n10402_), .B0(new_n10272_), .Y(new_n11347_));
  NOR2X1   g10345(.A(new_n10535_), .B(new_n10402_), .Y(new_n11348_));
  OR2X1    g10346(.A(new_n11348_), .B(new_n11347_), .Y(new_n11349_));
  AOI21X1  g10347(.A0(new_n2406_), .A1(new_n2393_), .B0(new_n2395_), .Y(new_n11350_));
  OAI21X1  g10348(.A0(new_n2384_), .A1(new_n2372_), .B0(new_n2374_), .Y(new_n11351_));
  XOR2X1   g10349(.A(new_n10532_), .B(new_n11351_), .Y(new_n11352_));
  AOI21X1  g10350(.A0(new_n11352_), .A1(new_n10466_), .B0(new_n11350_), .Y(new_n11353_));
  NOR2X1   g10351(.A(new_n11352_), .B(new_n10466_), .Y(new_n11354_));
  OR2X1    g10352(.A(new_n11354_), .B(new_n11353_), .Y(new_n11355_));
  OAI21X1  g10353(.A0(new_n2352_), .A1(new_n2265_), .B0(new_n2366_), .Y(new_n11356_));
  XOR2X1   g10354(.A(new_n10530_), .B(new_n11356_), .Y(new_n11357_));
  AOI21X1  g10355(.A0(new_n11357_), .A1(new_n10500_), .B0(new_n10467_), .Y(new_n11358_));
  NOR2X1   g10356(.A(new_n11357_), .B(new_n10500_), .Y(new_n11359_));
  OR2X1    g10357(.A(new_n11359_), .B(new_n11358_), .Y(new_n11360_));
  OAI22X1  g10358(.A0(new_n10528_), .A1(new_n10523_), .B0(new_n10513_), .B1(new_n10508_), .Y(new_n11361_));
  NOR4X1   g10359(.A(new_n10528_), .B(new_n10523_), .C(new_n10513_), .D(new_n10508_), .Y(new_n11362_));
  AOI21X1  g10360(.A0(new_n11361_), .A1(new_n11356_), .B0(new_n11362_), .Y(new_n11363_));
  AOI21X1  g10361(.A0(new_n2334_), .A1(new_n2332_), .B0(new_n10519_), .Y(new_n11364_));
  OAI21X1  g10362(.A0(new_n10515_), .A1(new_n2293_), .B0(new_n11364_), .Y(new_n11365_));
  AND2X1   g10363(.A(new_n11365_), .B(new_n10521_), .Y(new_n11366_));
  AND2X1   g10364(.A(new_n10519_), .B(new_n10518_), .Y(new_n11367_));
  OR2X1    g10365(.A(new_n11367_), .B(new_n11366_), .Y(new_n11368_));
  NAND3X1  g10366(.A(new_n10504_), .B(new_n10502_), .C(new_n2263_), .Y(new_n11369_));
  AOI21X1  g10367(.A0(new_n10502_), .A1(new_n2263_), .B0(new_n10504_), .Y(new_n11370_));
  AOI21X1  g10368(.A0(new_n11369_), .A1(new_n10506_), .B0(new_n11370_), .Y(new_n11371_));
  XOR2X1   g10369(.A(new_n11371_), .B(new_n11368_), .Y(new_n11372_));
  OR2X1    g10370(.A(new_n11372_), .B(new_n11363_), .Y(new_n11373_));
  NAND2X1  g10371(.A(new_n11361_), .B(new_n11356_), .Y(new_n11374_));
  OR2X1    g10372(.A(new_n11371_), .B(new_n11368_), .Y(new_n11375_));
  AOI21X1  g10373(.A0(new_n11371_), .A1(new_n11368_), .B0(new_n11362_), .Y(new_n11376_));
  NAND3X1  g10374(.A(new_n11376_), .B(new_n11375_), .C(new_n11374_), .Y(new_n11377_));
  NAND2X1  g10375(.A(new_n11377_), .B(new_n11373_), .Y(new_n11378_));
  AND2X1   g10376(.A(new_n10477_), .B(new_n10472_), .Y(new_n11379_));
  OR2X1    g10377(.A(new_n10482_), .B(new_n11379_), .Y(new_n11380_));
  OR2X1    g10378(.A(new_n10497_), .B(new_n10492_), .Y(new_n11381_));
  AOI21X1  g10379(.A0(new_n11381_), .A1(new_n11380_), .B0(new_n10470_), .Y(new_n11382_));
  NOR4X1   g10380(.A(new_n10497_), .B(new_n10492_), .C(new_n10482_), .D(new_n11379_), .Y(new_n11383_));
  AOI21X1  g10381(.A0(new_n2107_), .A1(new_n2105_), .B0(new_n10488_), .Y(new_n11384_));
  OAI21X1  g10382(.A0(new_n10484_), .A1(new_n2066_), .B0(new_n11384_), .Y(new_n11385_));
  AOI22X1  g10383(.A0(new_n11385_), .A1(new_n10490_), .B0(new_n10488_), .B1(new_n10487_), .Y(new_n11386_));
  OAI21X1  g10384(.A0(new_n2185_), .A1(new_n2182_), .B0(new_n10479_), .Y(new_n11387_));
  OAI21X1  g10385(.A0(new_n11387_), .A1(new_n10471_), .B0(new_n10476_), .Y(new_n11388_));
  OAI21X1  g10386(.A0(new_n10471_), .A1(new_n2186_), .B0(new_n10474_), .Y(new_n11389_));
  NAND2X1  g10387(.A(new_n11389_), .B(new_n11388_), .Y(new_n11390_));
  INVX1    g10388(.A(new_n11390_), .Y(new_n11391_));
  XOR2X1   g10389(.A(new_n11391_), .B(new_n11386_), .Y(new_n11392_));
  OAI21X1  g10390(.A0(new_n11383_), .A1(new_n11382_), .B0(new_n11392_), .Y(new_n11393_));
  AND2X1   g10391(.A(new_n2191_), .B(new_n10468_), .Y(new_n11394_));
  OAI22X1  g10392(.A0(new_n10498_), .A1(new_n10483_), .B0(new_n11394_), .B1(new_n10469_), .Y(new_n11395_));
  OR4X1    g10393(.A(new_n10497_), .B(new_n10492_), .C(new_n10482_), .D(new_n11379_), .Y(new_n11396_));
  OR2X1    g10394(.A(new_n11390_), .B(new_n11386_), .Y(new_n11397_));
  NAND2X1  g10395(.A(new_n11390_), .B(new_n11386_), .Y(new_n11398_));
  NAND4X1  g10396(.A(new_n11398_), .B(new_n11397_), .C(new_n11396_), .D(new_n11395_), .Y(new_n11399_));
  AND2X1   g10397(.A(new_n11399_), .B(new_n11393_), .Y(new_n11400_));
  XOR2X1   g10398(.A(new_n11400_), .B(new_n11378_), .Y(new_n11401_));
  XOR2X1   g10399(.A(new_n11401_), .B(new_n11360_), .Y(new_n11402_));
  NOR3X1   g10400(.A(new_n1986_), .B(new_n1991_), .C(new_n1988_), .Y(new_n11403_));
  OAI21X1  g10401(.A0(new_n11403_), .A1(new_n2030_), .B0(new_n2032_), .Y(new_n11404_));
  XOR2X1   g10402(.A(new_n10432_), .B(new_n11404_), .Y(new_n11405_));
  OAI21X1  g10403(.A0(new_n10464_), .A1(new_n11405_), .B0(new_n10404_), .Y(new_n11406_));
  OAI21X1  g10404(.A0(new_n1853_), .A1(new_n1766_), .B0(new_n1941_), .Y(new_n11407_));
  XOR2X1   g10405(.A(new_n10463_), .B(new_n11407_), .Y(new_n11408_));
  OR2X1    g10406(.A(new_n11408_), .B(new_n10433_), .Y(new_n11409_));
  AND2X1   g10407(.A(new_n11409_), .B(new_n11406_), .Y(new_n11410_));
  OAI22X1  g10408(.A0(new_n10461_), .A1(new_n10456_), .B0(new_n10446_), .B1(new_n10441_), .Y(new_n11411_));
  NOR4X1   g10409(.A(new_n10461_), .B(new_n10456_), .C(new_n10446_), .D(new_n10441_), .Y(new_n11412_));
  AOI21X1  g10410(.A0(new_n11411_), .A1(new_n11407_), .B0(new_n11412_), .Y(new_n11413_));
  AOI21X1  g10411(.A0(new_n1835_), .A1(new_n1833_), .B0(new_n10452_), .Y(new_n11414_));
  OAI21X1  g10412(.A0(new_n10448_), .A1(new_n1794_), .B0(new_n11414_), .Y(new_n11415_));
  AND2X1   g10413(.A(new_n11415_), .B(new_n10454_), .Y(new_n11416_));
  AND2X1   g10414(.A(new_n10452_), .B(new_n10451_), .Y(new_n11417_));
  OR2X1    g10415(.A(new_n11417_), .B(new_n11416_), .Y(new_n11418_));
  NAND3X1  g10416(.A(new_n10437_), .B(new_n10435_), .C(new_n1764_), .Y(new_n11419_));
  AOI21X1  g10417(.A0(new_n10435_), .A1(new_n1764_), .B0(new_n10437_), .Y(new_n11420_));
  AOI21X1  g10418(.A0(new_n11419_), .A1(new_n10439_), .B0(new_n11420_), .Y(new_n11421_));
  XOR2X1   g10419(.A(new_n11421_), .B(new_n11418_), .Y(new_n11422_));
  OR2X1    g10420(.A(new_n11422_), .B(new_n11413_), .Y(new_n11423_));
  NAND2X1  g10421(.A(new_n11411_), .B(new_n11407_), .Y(new_n11424_));
  OR2X1    g10422(.A(new_n11421_), .B(new_n11418_), .Y(new_n11425_));
  AOI21X1  g10423(.A0(new_n11421_), .A1(new_n11418_), .B0(new_n11412_), .Y(new_n11426_));
  NAND3X1  g10424(.A(new_n11426_), .B(new_n11425_), .C(new_n11424_), .Y(new_n11427_));
  NAND2X1  g10425(.A(new_n11427_), .B(new_n11423_), .Y(new_n11428_));
  NOR2X1   g10426(.A(new_n10431_), .B(new_n10419_), .Y(new_n11429_));
  AND2X1   g10427(.A(new_n10413_), .B(new_n10408_), .Y(new_n11430_));
  AND2X1   g10428(.A(new_n10425_), .B(new_n10421_), .Y(new_n11431_));
  OR4X1    g10429(.A(new_n10430_), .B(new_n11431_), .C(new_n10418_), .D(new_n11430_), .Y(new_n11432_));
  OAI21X1  g10430(.A0(new_n11429_), .A1(new_n10406_), .B0(new_n11432_), .Y(new_n11433_));
  OAI21X1  g10431(.A0(new_n1982_), .A1(new_n1981_), .B0(new_n10427_), .Y(new_n11434_));
  OAI21X1  g10432(.A0(new_n11434_), .A1(new_n10420_), .B0(new_n10424_), .Y(new_n11435_));
  OAI21X1  g10433(.A0(new_n10420_), .A1(new_n1983_), .B0(new_n10423_), .Y(new_n11436_));
  NAND2X1  g10434(.A(new_n11436_), .B(new_n11435_), .Y(new_n11437_));
  OAI21X1  g10435(.A0(new_n2023_), .A1(new_n2018_), .B0(new_n10415_), .Y(new_n11438_));
  OAI21X1  g10436(.A0(new_n11438_), .A1(new_n10407_), .B0(new_n10412_), .Y(new_n11439_));
  OAI21X1  g10437(.A0(new_n10407_), .A1(new_n2024_), .B0(new_n10410_), .Y(new_n11440_));
  AND2X1   g10438(.A(new_n11440_), .B(new_n11439_), .Y(new_n11441_));
  AND2X1   g10439(.A(new_n11441_), .B(new_n11437_), .Y(new_n11442_));
  NOR2X1   g10440(.A(new_n11441_), .B(new_n11437_), .Y(new_n11443_));
  OR2X1    g10441(.A(new_n11443_), .B(new_n11442_), .Y(new_n11444_));
  NAND2X1  g10442(.A(new_n11444_), .B(new_n11433_), .Y(new_n11445_));
  NOR4X1   g10443(.A(new_n10430_), .B(new_n11431_), .C(new_n10418_), .D(new_n11430_), .Y(new_n11446_));
  NOR3X1   g10444(.A(new_n11443_), .B(new_n11442_), .C(new_n11446_), .Y(new_n11447_));
  OAI21X1  g10445(.A0(new_n11429_), .A1(new_n10406_), .B0(new_n11447_), .Y(new_n11448_));
  AND2X1   g10446(.A(new_n11448_), .B(new_n11445_), .Y(new_n11449_));
  XOR2X1   g10447(.A(new_n11449_), .B(new_n11428_), .Y(new_n11450_));
  XOR2X1   g10448(.A(new_n11450_), .B(new_n11410_), .Y(new_n11451_));
  XOR2X1   g10449(.A(new_n11451_), .B(new_n11402_), .Y(new_n11452_));
  XOR2X1   g10450(.A(new_n11452_), .B(new_n11355_), .Y(new_n11453_));
  OAI21X1  g10451(.A0(new_n1692_), .A1(new_n2416_), .B0(new_n2418_), .Y(new_n11454_));
  AOI21X1  g10452(.A0(new_n2413_), .A1(new_n1687_), .B0(new_n1689_), .Y(new_n11455_));
  XOR2X1   g10453(.A(new_n10332_), .B(new_n11455_), .Y(new_n11456_));
  AOI21X1  g10454(.A0(new_n1500_), .A1(new_n1336_), .B0(new_n1338_), .Y(new_n11457_));
  XOR2X1   g10455(.A(new_n10399_), .B(new_n11457_), .Y(new_n11458_));
  OAI21X1  g10456(.A0(new_n11458_), .A1(new_n11456_), .B0(new_n11454_), .Y(new_n11459_));
  OR2X1    g10457(.A(new_n10400_), .B(new_n10333_), .Y(new_n11460_));
  AND2X1   g10458(.A(new_n11460_), .B(new_n11459_), .Y(new_n11461_));
  OAI21X1  g10459(.A0(new_n1329_), .A1(new_n1313_), .B0(new_n1316_), .Y(new_n11462_));
  XOR2X1   g10460(.A(new_n10397_), .B(new_n11462_), .Y(new_n11463_));
  AOI21X1  g10461(.A0(new_n11463_), .A1(new_n10367_), .B0(new_n11457_), .Y(new_n11464_));
  NOR2X1   g10462(.A(new_n11463_), .B(new_n10367_), .Y(new_n11465_));
  OR2X1    g10463(.A(new_n11465_), .B(new_n11464_), .Y(new_n11466_));
  OAI22X1  g10464(.A0(new_n10395_), .A1(new_n10390_), .B0(new_n10380_), .B1(new_n10375_), .Y(new_n11467_));
  NOR4X1   g10465(.A(new_n10395_), .B(new_n10390_), .C(new_n10380_), .D(new_n10375_), .Y(new_n11468_));
  AOI21X1  g10466(.A0(new_n11467_), .A1(new_n11462_), .B0(new_n11468_), .Y(new_n11469_));
  AOI21X1  g10467(.A0(new_n1296_), .A1(new_n1294_), .B0(new_n10386_), .Y(new_n11470_));
  OAI21X1  g10468(.A0(new_n10382_), .A1(new_n1255_), .B0(new_n11470_), .Y(new_n11471_));
  AND2X1   g10469(.A(new_n11471_), .B(new_n10388_), .Y(new_n11472_));
  AND2X1   g10470(.A(new_n10386_), .B(new_n10385_), .Y(new_n11473_));
  OR2X1    g10471(.A(new_n11473_), .B(new_n11472_), .Y(new_n11474_));
  NAND3X1  g10472(.A(new_n10371_), .B(new_n10369_), .C(new_n1225_), .Y(new_n11475_));
  AOI21X1  g10473(.A0(new_n10369_), .A1(new_n1225_), .B0(new_n10371_), .Y(new_n11476_));
  AOI21X1  g10474(.A0(new_n11475_), .A1(new_n10373_), .B0(new_n11476_), .Y(new_n11477_));
  XOR2X1   g10475(.A(new_n11477_), .B(new_n11474_), .Y(new_n11478_));
  OR2X1    g10476(.A(new_n11478_), .B(new_n11469_), .Y(new_n11479_));
  NAND2X1  g10477(.A(new_n11467_), .B(new_n11462_), .Y(new_n11480_));
  OR2X1    g10478(.A(new_n11477_), .B(new_n11474_), .Y(new_n11481_));
  AOI21X1  g10479(.A0(new_n11477_), .A1(new_n11474_), .B0(new_n11468_), .Y(new_n11482_));
  NAND3X1  g10480(.A(new_n11482_), .B(new_n11481_), .C(new_n11480_), .Y(new_n11483_));
  NAND2X1  g10481(.A(new_n11483_), .B(new_n11479_), .Y(new_n11484_));
  AND2X1   g10482(.A(new_n10344_), .B(new_n10339_), .Y(new_n11485_));
  OR2X1    g10483(.A(new_n10349_), .B(new_n11485_), .Y(new_n11486_));
  OR2X1    g10484(.A(new_n10364_), .B(new_n10359_), .Y(new_n11487_));
  AOI21X1  g10485(.A0(new_n11487_), .A1(new_n11486_), .B0(new_n10337_), .Y(new_n11488_));
  NOR4X1   g10486(.A(new_n10364_), .B(new_n10359_), .C(new_n10349_), .D(new_n11485_), .Y(new_n11489_));
  AOI21X1  g10487(.A0(new_n1071_), .A1(new_n1069_), .B0(new_n10355_), .Y(new_n11490_));
  OAI21X1  g10488(.A0(new_n10351_), .A1(new_n1030_), .B0(new_n11490_), .Y(new_n11491_));
  AOI22X1  g10489(.A0(new_n11491_), .A1(new_n10357_), .B0(new_n10355_), .B1(new_n10354_), .Y(new_n11492_));
  OAI21X1  g10490(.A0(new_n1149_), .A1(new_n1146_), .B0(new_n10346_), .Y(new_n11493_));
  OAI21X1  g10491(.A0(new_n11493_), .A1(new_n10338_), .B0(new_n10343_), .Y(new_n11494_));
  OAI21X1  g10492(.A0(new_n10338_), .A1(new_n1150_), .B0(new_n10341_), .Y(new_n11495_));
  NAND2X1  g10493(.A(new_n11495_), .B(new_n11494_), .Y(new_n11496_));
  INVX1    g10494(.A(new_n11496_), .Y(new_n11497_));
  XOR2X1   g10495(.A(new_n11497_), .B(new_n11492_), .Y(new_n11498_));
  OAI21X1  g10496(.A0(new_n11489_), .A1(new_n11488_), .B0(new_n11498_), .Y(new_n11499_));
  AND2X1   g10497(.A(new_n1155_), .B(new_n10335_), .Y(new_n11500_));
  OAI22X1  g10498(.A0(new_n10365_), .A1(new_n10350_), .B0(new_n11500_), .B1(new_n10336_), .Y(new_n11501_));
  OR4X1    g10499(.A(new_n10364_), .B(new_n10359_), .C(new_n10349_), .D(new_n11485_), .Y(new_n11502_));
  OR2X1    g10500(.A(new_n11496_), .B(new_n11492_), .Y(new_n11503_));
  NAND2X1  g10501(.A(new_n11496_), .B(new_n11492_), .Y(new_n11504_));
  NAND4X1  g10502(.A(new_n11504_), .B(new_n11503_), .C(new_n11502_), .D(new_n11501_), .Y(new_n11505_));
  AND2X1   g10503(.A(new_n11505_), .B(new_n11499_), .Y(new_n11506_));
  XOR2X1   g10504(.A(new_n11506_), .B(new_n11484_), .Y(new_n11507_));
  XOR2X1   g10505(.A(new_n11507_), .B(new_n11466_), .Y(new_n11508_));
  AOI21X1  g10506(.A0(new_n1597_), .A1(new_n1587_), .B0(new_n1589_), .Y(new_n11509_));
  XOR2X1   g10507(.A(new_n10330_), .B(new_n11509_), .Y(new_n11510_));
  NAND2X1  g10508(.A(new_n11510_), .B(new_n10303_), .Y(new_n11511_));
  NOR2X1   g10509(.A(new_n11510_), .B(new_n10303_), .Y(new_n11512_));
  AOI21X1  g10510(.A0(new_n11511_), .A1(new_n10274_), .B0(new_n11512_), .Y(new_n11513_));
  OR2X1    g10511(.A(new_n10329_), .B(new_n10317_), .Y(new_n11514_));
  AND2X1   g10512(.A(new_n10311_), .B(new_n10306_), .Y(new_n11515_));
  AND2X1   g10513(.A(new_n10323_), .B(new_n10319_), .Y(new_n11516_));
  NOR4X1   g10514(.A(new_n10328_), .B(new_n11516_), .C(new_n10316_), .D(new_n11515_), .Y(new_n11517_));
  AOI21X1  g10515(.A0(new_n11514_), .A1(new_n10304_), .B0(new_n11517_), .Y(new_n11518_));
  OAI21X1  g10516(.A0(new_n1569_), .A1(new_n1564_), .B0(new_n10325_), .Y(new_n11519_));
  OAI21X1  g10517(.A0(new_n11519_), .A1(new_n10318_), .B0(new_n10322_), .Y(new_n11520_));
  OAI21X1  g10518(.A0(new_n10318_), .A1(new_n1582_), .B0(new_n10321_), .Y(new_n11521_));
  NAND2X1  g10519(.A(new_n11521_), .B(new_n11520_), .Y(new_n11522_));
  OAI21X1  g10520(.A0(new_n1534_), .A1(new_n1532_), .B0(new_n10313_), .Y(new_n11523_));
  OR2X1    g10521(.A(new_n11523_), .B(new_n10305_), .Y(new_n11524_));
  AOI22X1  g10522(.A0(new_n11524_), .A1(new_n10310_), .B0(new_n10308_), .B1(new_n10306_), .Y(new_n11525_));
  XOR2X1   g10523(.A(new_n11525_), .B(new_n11522_), .Y(new_n11526_));
  OR2X1    g10524(.A(new_n11526_), .B(new_n11518_), .Y(new_n11527_));
  NAND2X1  g10525(.A(new_n11514_), .B(new_n10304_), .Y(new_n11528_));
  OR4X1    g10526(.A(new_n10328_), .B(new_n11516_), .C(new_n10316_), .D(new_n11515_), .Y(new_n11529_));
  NAND2X1  g10527(.A(new_n11525_), .B(new_n11522_), .Y(new_n11530_));
  OR2X1    g10528(.A(new_n11525_), .B(new_n11522_), .Y(new_n11531_));
  NAND4X1  g10529(.A(new_n11531_), .B(new_n11530_), .C(new_n11529_), .D(new_n11528_), .Y(new_n11532_));
  NAND2X1  g10530(.A(new_n11532_), .B(new_n11527_), .Y(new_n11533_));
  NOR2X1   g10531(.A(new_n10301_), .B(new_n10289_), .Y(new_n11534_));
  AND2X1   g10532(.A(new_n10283_), .B(new_n10278_), .Y(new_n11535_));
  AND2X1   g10533(.A(new_n10295_), .B(new_n10291_), .Y(new_n11536_));
  OR4X1    g10534(.A(new_n10300_), .B(new_n11536_), .C(new_n10288_), .D(new_n11535_), .Y(new_n11537_));
  OAI21X1  g10535(.A0(new_n11534_), .A1(new_n10276_), .B0(new_n11537_), .Y(new_n11538_));
  OAI21X1  g10536(.A0(new_n1639_), .A1(new_n1638_), .B0(new_n10297_), .Y(new_n11539_));
  OAI21X1  g10537(.A0(new_n11539_), .A1(new_n10290_), .B0(new_n10294_), .Y(new_n11540_));
  OAI21X1  g10538(.A0(new_n10290_), .A1(new_n1640_), .B0(new_n10293_), .Y(new_n11541_));
  AND2X1   g10539(.A(new_n11541_), .B(new_n11540_), .Y(new_n11542_));
  OAI21X1  g10540(.A0(new_n1676_), .A1(new_n1674_), .B0(new_n10285_), .Y(new_n11543_));
  OR2X1    g10541(.A(new_n11543_), .B(new_n10277_), .Y(new_n11544_));
  AOI22X1  g10542(.A0(new_n11544_), .A1(new_n10282_), .B0(new_n10280_), .B1(new_n10278_), .Y(new_n11545_));
  XOR2X1   g10543(.A(new_n11545_), .B(new_n11542_), .Y(new_n11546_));
  NAND2X1  g10544(.A(new_n11546_), .B(new_n11538_), .Y(new_n11547_));
  OR2X1    g10545(.A(new_n11534_), .B(new_n10276_), .Y(new_n11548_));
  NAND2X1  g10546(.A(new_n11541_), .B(new_n11540_), .Y(new_n11549_));
  NAND2X1  g10547(.A(new_n11545_), .B(new_n11549_), .Y(new_n11550_));
  OR2X1    g10548(.A(new_n11545_), .B(new_n11549_), .Y(new_n11551_));
  NAND4X1  g10549(.A(new_n11551_), .B(new_n11550_), .C(new_n11537_), .D(new_n11548_), .Y(new_n11552_));
  AND2X1   g10550(.A(new_n11552_), .B(new_n11547_), .Y(new_n11553_));
  XOR2X1   g10551(.A(new_n11553_), .B(new_n11533_), .Y(new_n11554_));
  XOR2X1   g10552(.A(new_n11554_), .B(new_n11513_), .Y(new_n11555_));
  XOR2X1   g10553(.A(new_n11555_), .B(new_n11508_), .Y(new_n11556_));
  XOR2X1   g10554(.A(new_n11556_), .B(new_n11461_), .Y(new_n11557_));
  XOR2X1   g10555(.A(new_n11557_), .B(new_n11453_), .Y(new_n11558_));
  XOR2X1   g10556(.A(new_n11558_), .B(new_n11349_), .Y(new_n11559_));
  NOR3X1   g10557(.A(new_n3440_), .B(new_n3447_), .C(new_n3444_), .Y(new_n11560_));
  OAI21X1  g10558(.A0(new_n11560_), .A1(new_n3838_), .B0(new_n3840_), .Y(new_n11561_));
  OAI21X1  g10559(.A0(new_n10016_), .A1(new_n3834_), .B0(new_n3836_), .Y(new_n11562_));
  XOR2X1   g10560(.A(new_n10144_), .B(new_n11562_), .Y(new_n11563_));
  AOI21X1  g10561(.A0(new_n3445_), .A1(new_n3435_), .B0(new_n3437_), .Y(new_n11564_));
  XOR2X1   g10562(.A(new_n10267_), .B(new_n11564_), .Y(new_n11565_));
  OAI21X1  g10563(.A0(new_n11565_), .A1(new_n11563_), .B0(new_n11561_), .Y(new_n11566_));
  OR2X1    g10564(.A(new_n10268_), .B(new_n10145_), .Y(new_n11567_));
  AND2X1   g10565(.A(new_n11567_), .B(new_n11566_), .Y(new_n11568_));
  OAI21X1  g10566(.A0(new_n3426_), .A1(new_n3415_), .B0(new_n3417_), .Y(new_n11569_));
  XOR2X1   g10567(.A(new_n10265_), .B(new_n11569_), .Y(new_n11570_));
  AND2X1   g10568(.A(new_n11570_), .B(new_n10206_), .Y(new_n11571_));
  OR2X1    g10569(.A(new_n11570_), .B(new_n10206_), .Y(new_n11572_));
  OAI21X1  g10570(.A0(new_n11571_), .A1(new_n11564_), .B0(new_n11572_), .Y(new_n11573_));
  AOI21X1  g10571(.A0(new_n3409_), .A1(new_n3400_), .B0(new_n3402_), .Y(new_n11574_));
  XOR2X1   g10572(.A(new_n10263_), .B(new_n11574_), .Y(new_n11575_));
  NAND2X1  g10573(.A(new_n11575_), .B(new_n10236_), .Y(new_n11576_));
  AND2X1   g10574(.A(new_n11576_), .B(new_n11569_), .Y(new_n11577_));
  NOR2X1   g10575(.A(new_n11575_), .B(new_n10236_), .Y(new_n11578_));
  OR2X1    g10576(.A(new_n11578_), .B(new_n11577_), .Y(new_n11579_));
  OR2X1    g10577(.A(new_n10262_), .B(new_n10250_), .Y(new_n11580_));
  AND2X1   g10578(.A(new_n10244_), .B(new_n10239_), .Y(new_n11581_));
  AND2X1   g10579(.A(new_n10256_), .B(new_n10252_), .Y(new_n11582_));
  NOR4X1   g10580(.A(new_n10261_), .B(new_n11582_), .C(new_n10249_), .D(new_n11581_), .Y(new_n11583_));
  AOI21X1  g10581(.A0(new_n11580_), .A1(new_n10237_), .B0(new_n11583_), .Y(new_n11584_));
  OAI21X1  g10582(.A0(new_n3382_), .A1(new_n3377_), .B0(new_n10258_), .Y(new_n11585_));
  OAI21X1  g10583(.A0(new_n11585_), .A1(new_n10251_), .B0(new_n10255_), .Y(new_n11586_));
  OAI21X1  g10584(.A0(new_n10251_), .A1(new_n3395_), .B0(new_n10254_), .Y(new_n11587_));
  NAND2X1  g10585(.A(new_n11587_), .B(new_n11586_), .Y(new_n11588_));
  OAI21X1  g10586(.A0(new_n3347_), .A1(new_n3345_), .B0(new_n10246_), .Y(new_n11589_));
  OR2X1    g10587(.A(new_n11589_), .B(new_n10238_), .Y(new_n11590_));
  AOI22X1  g10588(.A0(new_n11590_), .A1(new_n10243_), .B0(new_n10241_), .B1(new_n10239_), .Y(new_n11591_));
  XOR2X1   g10589(.A(new_n11591_), .B(new_n11588_), .Y(new_n11592_));
  OR2X1    g10590(.A(new_n11592_), .B(new_n11584_), .Y(new_n11593_));
  NAND2X1  g10591(.A(new_n11580_), .B(new_n10237_), .Y(new_n11594_));
  OR4X1    g10592(.A(new_n10261_), .B(new_n11582_), .C(new_n10249_), .D(new_n11581_), .Y(new_n11595_));
  NAND2X1  g10593(.A(new_n11591_), .B(new_n11588_), .Y(new_n11596_));
  OR2X1    g10594(.A(new_n11591_), .B(new_n11588_), .Y(new_n11597_));
  NAND4X1  g10595(.A(new_n11597_), .B(new_n11596_), .C(new_n11595_), .D(new_n11594_), .Y(new_n11598_));
  NAND2X1  g10596(.A(new_n11598_), .B(new_n11593_), .Y(new_n11599_));
  NOR2X1   g10597(.A(new_n10234_), .B(new_n10222_), .Y(new_n11600_));
  AND2X1   g10598(.A(new_n10216_), .B(new_n10211_), .Y(new_n11601_));
  AND2X1   g10599(.A(new_n10228_), .B(new_n10224_), .Y(new_n11602_));
  OR4X1    g10600(.A(new_n10233_), .B(new_n11602_), .C(new_n10221_), .D(new_n11601_), .Y(new_n11603_));
  OAI21X1  g10601(.A0(new_n11600_), .A1(new_n10209_), .B0(new_n11603_), .Y(new_n11604_));
  OAI21X1  g10602(.A0(new_n3269_), .A1(new_n3268_), .B0(new_n10230_), .Y(new_n11605_));
  OAI21X1  g10603(.A0(new_n11605_), .A1(new_n10223_), .B0(new_n10227_), .Y(new_n11606_));
  OAI21X1  g10604(.A0(new_n10223_), .A1(new_n3270_), .B0(new_n10226_), .Y(new_n11607_));
  AND2X1   g10605(.A(new_n11607_), .B(new_n11606_), .Y(new_n11608_));
  OAI21X1  g10606(.A0(new_n3307_), .A1(new_n3305_), .B0(new_n10218_), .Y(new_n11609_));
  OR2X1    g10607(.A(new_n11609_), .B(new_n10210_), .Y(new_n11610_));
  AOI22X1  g10608(.A0(new_n11610_), .A1(new_n10215_), .B0(new_n10213_), .B1(new_n10211_), .Y(new_n11611_));
  XOR2X1   g10609(.A(new_n11611_), .B(new_n11608_), .Y(new_n11612_));
  NAND2X1  g10610(.A(new_n11612_), .B(new_n11604_), .Y(new_n11613_));
  OR2X1    g10611(.A(new_n11600_), .B(new_n10209_), .Y(new_n11614_));
  NAND2X1  g10612(.A(new_n11607_), .B(new_n11606_), .Y(new_n11615_));
  NAND2X1  g10613(.A(new_n11611_), .B(new_n11615_), .Y(new_n11616_));
  OR2X1    g10614(.A(new_n11611_), .B(new_n11615_), .Y(new_n11617_));
  NAND4X1  g10615(.A(new_n11617_), .B(new_n11616_), .C(new_n11603_), .D(new_n11614_), .Y(new_n11618_));
  AND2X1   g10616(.A(new_n11618_), .B(new_n11613_), .Y(new_n11619_));
  XOR2X1   g10617(.A(new_n11619_), .B(new_n11599_), .Y(new_n11620_));
  XOR2X1   g10618(.A(new_n11620_), .B(new_n11579_), .Y(new_n11621_));
  OAI21X1  g10619(.A0(new_n3432_), .A1(new_n3228_), .B0(new_n3230_), .Y(new_n11622_));
  NAND2X1  g10620(.A(new_n10204_), .B(new_n10176_), .Y(new_n11623_));
  NOR2X1   g10621(.A(new_n10204_), .B(new_n10176_), .Y(new_n11624_));
  AOI21X1  g10622(.A0(new_n11623_), .A1(new_n11622_), .B0(new_n11624_), .Y(new_n11625_));
  OAI21X1  g10623(.A0(new_n3129_), .A1(new_n3078_), .B0(new_n3139_), .Y(new_n11626_));
  OR2X1    g10624(.A(new_n10202_), .B(new_n10190_), .Y(new_n11627_));
  AND2X1   g10625(.A(new_n10184_), .B(new_n10179_), .Y(new_n11628_));
  AND2X1   g10626(.A(new_n10196_), .B(new_n10192_), .Y(new_n11629_));
  NOR4X1   g10627(.A(new_n10201_), .B(new_n11629_), .C(new_n10189_), .D(new_n11628_), .Y(new_n11630_));
  AOI21X1  g10628(.A0(new_n11627_), .A1(new_n11626_), .B0(new_n11630_), .Y(new_n11631_));
  OAI21X1  g10629(.A0(new_n3110_), .A1(new_n3105_), .B0(new_n10198_), .Y(new_n11632_));
  OAI21X1  g10630(.A0(new_n11632_), .A1(new_n10191_), .B0(new_n10195_), .Y(new_n11633_));
  OAI21X1  g10631(.A0(new_n10191_), .A1(new_n3123_), .B0(new_n10194_), .Y(new_n11634_));
  NAND2X1  g10632(.A(new_n11634_), .B(new_n11633_), .Y(new_n11635_));
  OAI21X1  g10633(.A0(new_n3075_), .A1(new_n3073_), .B0(new_n10186_), .Y(new_n11636_));
  OR2X1    g10634(.A(new_n11636_), .B(new_n10178_), .Y(new_n11637_));
  AOI22X1  g10635(.A0(new_n11637_), .A1(new_n10183_), .B0(new_n10181_), .B1(new_n10179_), .Y(new_n11638_));
  XOR2X1   g10636(.A(new_n11638_), .B(new_n11635_), .Y(new_n11639_));
  OR2X1    g10637(.A(new_n11639_), .B(new_n11631_), .Y(new_n11640_));
  NAND2X1  g10638(.A(new_n11627_), .B(new_n11626_), .Y(new_n11641_));
  OR4X1    g10639(.A(new_n10201_), .B(new_n11629_), .C(new_n10189_), .D(new_n11628_), .Y(new_n11642_));
  NAND2X1  g10640(.A(new_n11638_), .B(new_n11635_), .Y(new_n11643_));
  OR2X1    g10641(.A(new_n11638_), .B(new_n11635_), .Y(new_n11644_));
  NAND4X1  g10642(.A(new_n11644_), .B(new_n11643_), .C(new_n11642_), .D(new_n11641_), .Y(new_n11645_));
  NAND2X1  g10643(.A(new_n11645_), .B(new_n11640_), .Y(new_n11646_));
  NOR2X1   g10644(.A(new_n10174_), .B(new_n10162_), .Y(new_n11647_));
  AND2X1   g10645(.A(new_n10156_), .B(new_n10151_), .Y(new_n11648_));
  AND2X1   g10646(.A(new_n10168_), .B(new_n10164_), .Y(new_n11649_));
  OR4X1    g10647(.A(new_n10173_), .B(new_n11649_), .C(new_n10161_), .D(new_n11648_), .Y(new_n11650_));
  OAI21X1  g10648(.A0(new_n11647_), .A1(new_n10149_), .B0(new_n11650_), .Y(new_n11651_));
  OAI21X1  g10649(.A0(new_n3180_), .A1(new_n3179_), .B0(new_n10170_), .Y(new_n11652_));
  OAI21X1  g10650(.A0(new_n11652_), .A1(new_n10163_), .B0(new_n10167_), .Y(new_n11653_));
  OAI21X1  g10651(.A0(new_n10163_), .A1(new_n3181_), .B0(new_n10166_), .Y(new_n11654_));
  AND2X1   g10652(.A(new_n11654_), .B(new_n11653_), .Y(new_n11655_));
  OAI21X1  g10653(.A0(new_n3217_), .A1(new_n3215_), .B0(new_n10158_), .Y(new_n11656_));
  OR2X1    g10654(.A(new_n11656_), .B(new_n10150_), .Y(new_n11657_));
  AOI22X1  g10655(.A0(new_n11657_), .A1(new_n10155_), .B0(new_n10153_), .B1(new_n10151_), .Y(new_n11658_));
  XOR2X1   g10656(.A(new_n11658_), .B(new_n11655_), .Y(new_n11659_));
  NAND2X1  g10657(.A(new_n11659_), .B(new_n11651_), .Y(new_n11660_));
  OR2X1    g10658(.A(new_n11647_), .B(new_n10149_), .Y(new_n11661_));
  NAND2X1  g10659(.A(new_n11654_), .B(new_n11653_), .Y(new_n11662_));
  NAND2X1  g10660(.A(new_n11658_), .B(new_n11662_), .Y(new_n11663_));
  OR2X1    g10661(.A(new_n11658_), .B(new_n11662_), .Y(new_n11664_));
  NAND4X1  g10662(.A(new_n11664_), .B(new_n11663_), .C(new_n11650_), .D(new_n11661_), .Y(new_n11665_));
  AND2X1   g10663(.A(new_n11665_), .B(new_n11660_), .Y(new_n11666_));
  XOR2X1   g10664(.A(new_n11666_), .B(new_n11646_), .Y(new_n11667_));
  XOR2X1   g10665(.A(new_n11667_), .B(new_n11625_), .Y(new_n11668_));
  XOR2X1   g10666(.A(new_n11668_), .B(new_n11621_), .Y(new_n11669_));
  XOR2X1   g10667(.A(new_n11669_), .B(new_n11573_), .Y(new_n11670_));
  AOI21X1  g10668(.A0(new_n3831_), .A1(new_n10011_), .B0(new_n10013_), .Y(new_n11671_));
  XOR2X1   g10669(.A(new_n10082_), .B(new_n11671_), .Y(new_n11672_));
  AOI21X1  g10670(.A0(new_n3642_), .A1(new_n3633_), .B0(new_n3635_), .Y(new_n11673_));
  XOR2X1   g10671(.A(new_n10142_), .B(new_n11673_), .Y(new_n11674_));
  OAI21X1  g10672(.A0(new_n11674_), .A1(new_n11672_), .B0(new_n11562_), .Y(new_n11675_));
  OR2X1    g10673(.A(new_n10143_), .B(new_n10083_), .Y(new_n11676_));
  AND2X1   g10674(.A(new_n11676_), .B(new_n11675_), .Y(new_n11677_));
  AOI21X1  g10675(.A0(new_n3618_), .A1(new_n3565_), .B0(new_n3629_), .Y(new_n11678_));
  XOR2X1   g10676(.A(new_n10140_), .B(new_n11678_), .Y(new_n11679_));
  NAND2X1  g10677(.A(new_n11679_), .B(new_n10113_), .Y(new_n11680_));
  AND2X1   g10678(.A(new_n11680_), .B(new_n10084_), .Y(new_n11681_));
  NOR2X1   g10679(.A(new_n11679_), .B(new_n10113_), .Y(new_n11682_));
  OR2X1    g10680(.A(new_n11682_), .B(new_n11681_), .Y(new_n11683_));
  OR2X1    g10681(.A(new_n10139_), .B(new_n10127_), .Y(new_n11684_));
  AND2X1   g10682(.A(new_n10121_), .B(new_n10116_), .Y(new_n11685_));
  AND2X1   g10683(.A(new_n10133_), .B(new_n10129_), .Y(new_n11686_));
  NOR4X1   g10684(.A(new_n10138_), .B(new_n11686_), .C(new_n10126_), .D(new_n11685_), .Y(new_n11687_));
  AOI21X1  g10685(.A0(new_n11684_), .A1(new_n10114_), .B0(new_n11687_), .Y(new_n11688_));
  OAI21X1  g10686(.A0(new_n3602_), .A1(new_n3601_), .B0(new_n10135_), .Y(new_n11689_));
  OAI21X1  g10687(.A0(new_n11689_), .A1(new_n10128_), .B0(new_n10132_), .Y(new_n11690_));
  OAI21X1  g10688(.A0(new_n10128_), .A1(new_n3603_), .B0(new_n10131_), .Y(new_n11691_));
  NAND2X1  g10689(.A(new_n11691_), .B(new_n11690_), .Y(new_n11692_));
  OAI21X1  g10690(.A0(new_n3562_), .A1(new_n3560_), .B0(new_n10123_), .Y(new_n11693_));
  OR2X1    g10691(.A(new_n11693_), .B(new_n10115_), .Y(new_n11694_));
  AOI22X1  g10692(.A0(new_n11694_), .A1(new_n10120_), .B0(new_n10118_), .B1(new_n10116_), .Y(new_n11695_));
  XOR2X1   g10693(.A(new_n11695_), .B(new_n11692_), .Y(new_n11696_));
  OR2X1    g10694(.A(new_n11696_), .B(new_n11688_), .Y(new_n11697_));
  NAND2X1  g10695(.A(new_n11684_), .B(new_n10114_), .Y(new_n11698_));
  OR4X1    g10696(.A(new_n10138_), .B(new_n11686_), .C(new_n10126_), .D(new_n11685_), .Y(new_n11699_));
  NAND2X1  g10697(.A(new_n11695_), .B(new_n11692_), .Y(new_n11700_));
  OR2X1    g10698(.A(new_n11695_), .B(new_n11692_), .Y(new_n11701_));
  NAND4X1  g10699(.A(new_n11701_), .B(new_n11700_), .C(new_n11699_), .D(new_n11698_), .Y(new_n11702_));
  NAND2X1  g10700(.A(new_n11702_), .B(new_n11697_), .Y(new_n11703_));
  NOR2X1   g10701(.A(new_n10111_), .B(new_n10099_), .Y(new_n11704_));
  AND2X1   g10702(.A(new_n10093_), .B(new_n10088_), .Y(new_n11705_));
  AND2X1   g10703(.A(new_n10105_), .B(new_n10101_), .Y(new_n11706_));
  OR4X1    g10704(.A(new_n10110_), .B(new_n11706_), .C(new_n10098_), .D(new_n11705_), .Y(new_n11707_));
  OAI21X1  g10705(.A0(new_n11704_), .A1(new_n10086_), .B0(new_n11707_), .Y(new_n11708_));
  OAI21X1  g10706(.A0(new_n3487_), .A1(new_n3486_), .B0(new_n10107_), .Y(new_n11709_));
  OAI21X1  g10707(.A0(new_n11709_), .A1(new_n10100_), .B0(new_n10104_), .Y(new_n11710_));
  OAI21X1  g10708(.A0(new_n10100_), .A1(new_n3488_), .B0(new_n10103_), .Y(new_n11711_));
  AND2X1   g10709(.A(new_n11711_), .B(new_n11710_), .Y(new_n11712_));
  OAI21X1  g10710(.A0(new_n3524_), .A1(new_n3522_), .B0(new_n10095_), .Y(new_n11713_));
  OR2X1    g10711(.A(new_n11713_), .B(new_n10087_), .Y(new_n11714_));
  AOI22X1  g10712(.A0(new_n11714_), .A1(new_n10092_), .B0(new_n10090_), .B1(new_n10088_), .Y(new_n11715_));
  XOR2X1   g10713(.A(new_n11715_), .B(new_n11712_), .Y(new_n11716_));
  NAND2X1  g10714(.A(new_n11716_), .B(new_n11708_), .Y(new_n11717_));
  OR2X1    g10715(.A(new_n11704_), .B(new_n10086_), .Y(new_n11718_));
  NAND2X1  g10716(.A(new_n11711_), .B(new_n11710_), .Y(new_n11719_));
  NAND2X1  g10717(.A(new_n11715_), .B(new_n11719_), .Y(new_n11720_));
  OR2X1    g10718(.A(new_n11715_), .B(new_n11719_), .Y(new_n11721_));
  NAND4X1  g10719(.A(new_n11721_), .B(new_n11720_), .C(new_n11707_), .D(new_n11718_), .Y(new_n11722_));
  AND2X1   g10720(.A(new_n11722_), .B(new_n11717_), .Y(new_n11723_));
  XOR2X1   g10721(.A(new_n11723_), .B(new_n11703_), .Y(new_n11724_));
  XOR2X1   g10722(.A(new_n11724_), .B(new_n11683_), .Y(new_n11725_));
  OR2X1    g10723(.A(new_n10038_), .B(new_n10033_), .Y(new_n11726_));
  XOR2X1   g10724(.A(new_n10051_), .B(new_n11726_), .Y(new_n11727_));
  XOR2X1   g10725(.A(new_n11727_), .B(new_n10025_), .Y(new_n11728_));
  OAI21X1  g10726(.A0(new_n10081_), .A1(new_n11728_), .B0(new_n10023_), .Y(new_n11729_));
  AOI21X1  g10727(.A0(new_n3738_), .A1(new_n3728_), .B0(new_n3730_), .Y(new_n11730_));
  XOR2X1   g10728(.A(new_n10080_), .B(new_n11730_), .Y(new_n11731_));
  OR2X1    g10729(.A(new_n11731_), .B(new_n10053_), .Y(new_n11732_));
  AND2X1   g10730(.A(new_n11732_), .B(new_n11729_), .Y(new_n11733_));
  OR2X1    g10731(.A(new_n10079_), .B(new_n10067_), .Y(new_n11734_));
  AND2X1   g10732(.A(new_n10061_), .B(new_n10056_), .Y(new_n11735_));
  AND2X1   g10733(.A(new_n10073_), .B(new_n10069_), .Y(new_n11736_));
  NOR4X1   g10734(.A(new_n10078_), .B(new_n11736_), .C(new_n10066_), .D(new_n11735_), .Y(new_n11737_));
  AOI21X1  g10735(.A0(new_n11734_), .A1(new_n10054_), .B0(new_n11737_), .Y(new_n11738_));
  OAI21X1  g10736(.A0(new_n3711_), .A1(new_n3706_), .B0(new_n10075_), .Y(new_n11739_));
  OAI21X1  g10737(.A0(new_n11739_), .A1(new_n10068_), .B0(new_n10072_), .Y(new_n11740_));
  OAI21X1  g10738(.A0(new_n10068_), .A1(new_n3723_), .B0(new_n10071_), .Y(new_n11741_));
  NAND2X1  g10739(.A(new_n11741_), .B(new_n11740_), .Y(new_n11742_));
  OAI21X1  g10740(.A0(new_n3676_), .A1(new_n3674_), .B0(new_n10063_), .Y(new_n11743_));
  OR2X1    g10741(.A(new_n11743_), .B(new_n10055_), .Y(new_n11744_));
  AOI22X1  g10742(.A0(new_n11744_), .A1(new_n10060_), .B0(new_n10058_), .B1(new_n10056_), .Y(new_n11745_));
  XOR2X1   g10743(.A(new_n11745_), .B(new_n11742_), .Y(new_n11746_));
  OR2X1    g10744(.A(new_n11746_), .B(new_n11738_), .Y(new_n11747_));
  NAND2X1  g10745(.A(new_n11734_), .B(new_n10054_), .Y(new_n11748_));
  OR4X1    g10746(.A(new_n10078_), .B(new_n11736_), .C(new_n10066_), .D(new_n11735_), .Y(new_n11749_));
  NAND2X1  g10747(.A(new_n11745_), .B(new_n11742_), .Y(new_n11750_));
  OR2X1    g10748(.A(new_n11745_), .B(new_n11742_), .Y(new_n11751_));
  NAND4X1  g10749(.A(new_n11751_), .B(new_n11750_), .C(new_n11749_), .D(new_n11748_), .Y(new_n11752_));
  NAND2X1  g10750(.A(new_n11752_), .B(new_n11747_), .Y(new_n11753_));
  AND2X1   g10751(.A(new_n10045_), .B(new_n10041_), .Y(new_n11754_));
  OR2X1    g10752(.A(new_n10050_), .B(new_n11754_), .Y(new_n11755_));
  AOI21X1  g10753(.A0(new_n11755_), .A1(new_n11726_), .B0(new_n10025_), .Y(new_n11756_));
  NOR4X1   g10754(.A(new_n10050_), .B(new_n11754_), .C(new_n10038_), .D(new_n10033_), .Y(new_n11757_));
  OAI21X1  g10755(.A0(new_n3776_), .A1(new_n3775_), .B0(new_n10047_), .Y(new_n11758_));
  OAI21X1  g10756(.A0(new_n11758_), .A1(new_n10040_), .B0(new_n10044_), .Y(new_n11759_));
  OAI21X1  g10757(.A0(new_n10040_), .A1(new_n3777_), .B0(new_n10043_), .Y(new_n11760_));
  AND2X1   g10758(.A(new_n11760_), .B(new_n11759_), .Y(new_n11761_));
  NAND3X1  g10759(.A(new_n10029_), .B(new_n10027_), .C(new_n10026_), .Y(new_n11762_));
  AOI21X1  g10760(.A0(new_n10027_), .A1(new_n10026_), .B0(new_n10029_), .Y(new_n11763_));
  AOI21X1  g10761(.A0(new_n11762_), .A1(new_n10031_), .B0(new_n11763_), .Y(new_n11764_));
  XOR2X1   g10762(.A(new_n11764_), .B(new_n11761_), .Y(new_n11765_));
  OAI21X1  g10763(.A0(new_n11757_), .A1(new_n11756_), .B0(new_n11765_), .Y(new_n11766_));
  AND2X1   g10764(.A(new_n3827_), .B(new_n3822_), .Y(new_n11767_));
  OAI22X1  g10765(.A0(new_n10051_), .A1(new_n10039_), .B0(new_n11767_), .B1(new_n10024_), .Y(new_n11768_));
  OR4X1    g10766(.A(new_n10050_), .B(new_n11754_), .C(new_n10038_), .D(new_n10033_), .Y(new_n11769_));
  NAND2X1  g10767(.A(new_n11760_), .B(new_n11759_), .Y(new_n11770_));
  NAND2X1  g10768(.A(new_n11764_), .B(new_n11770_), .Y(new_n11771_));
  OR2X1    g10769(.A(new_n11764_), .B(new_n11770_), .Y(new_n11772_));
  NAND4X1  g10770(.A(new_n11772_), .B(new_n11771_), .C(new_n11769_), .D(new_n11768_), .Y(new_n11773_));
  AND2X1   g10771(.A(new_n11773_), .B(new_n11766_), .Y(new_n11774_));
  XOR2X1   g10772(.A(new_n11774_), .B(new_n11753_), .Y(new_n11775_));
  XOR2X1   g10773(.A(new_n11775_), .B(new_n11733_), .Y(new_n11776_));
  XOR2X1   g10774(.A(new_n11776_), .B(new_n11725_), .Y(new_n11777_));
  XOR2X1   g10775(.A(new_n11777_), .B(new_n11677_), .Y(new_n11778_));
  XOR2X1   g10776(.A(new_n11778_), .B(new_n11670_), .Y(new_n11779_));
  XOR2X1   g10777(.A(new_n11779_), .B(new_n11568_), .Y(new_n11780_));
  XOR2X1   g10778(.A(new_n11780_), .B(new_n11559_), .Y(new_n11781_));
  XOR2X1   g10779(.A(new_n11781_), .B(new_n11346_), .Y(new_n11782_));
  AND2X1   g10780(.A(new_n11782_), .B(new_n11343_), .Y(new_n11783_));
  XOR2X1   g10781(.A(new_n10269_), .B(new_n11561_), .Y(new_n11784_));
  NOR3X1   g10782(.A(new_n2401_), .B(new_n2408_), .C(new_n2405_), .Y(new_n11785_));
  OAI21X1  g10783(.A0(new_n11785_), .A1(new_n2420_), .B0(new_n2422_), .Y(new_n11786_));
  XOR2X1   g10784(.A(new_n10536_), .B(new_n11786_), .Y(new_n11787_));
  OAI21X1  g10785(.A0(new_n11787_), .A1(new_n11784_), .B0(new_n10550_), .Y(new_n11788_));
  OR2X1    g10786(.A(new_n10537_), .B(new_n10270_), .Y(new_n11789_));
  AND2X1   g10787(.A(new_n11789_), .B(new_n11788_), .Y(new_n11790_));
  XOR2X1   g10788(.A(new_n11781_), .B(new_n11790_), .Y(new_n11791_));
  OAI21X1  g10789(.A0(new_n11338_), .A1(new_n10557_), .B0(new_n11791_), .Y(new_n11792_));
  OAI22X1  g10790(.A0(new_n11792_), .A1(new_n11339_), .B0(new_n11783_), .B1(new_n10554_), .Y(new_n11793_));
  OR2X1    g10791(.A(new_n10808_), .B(new_n10807_), .Y(new_n11794_));
  XOR2X1   g10792(.A(new_n9622_), .B(new_n11794_), .Y(new_n11795_));
  AND2X1   g10793(.A(new_n8802_), .B(new_n8747_), .Y(new_n11796_));
  AOI21X1  g10794(.A0(new_n8806_), .A1(new_n8805_), .B0(new_n8800_), .Y(new_n11797_));
  OR2X1    g10795(.A(new_n11797_), .B(new_n11796_), .Y(new_n11798_));
  XOR2X1   g10796(.A(new_n10002_), .B(new_n11798_), .Y(new_n11799_));
  OAI22X1  g10797(.A0(new_n11799_), .A1(new_n11795_), .B0(new_n9234_), .B1(new_n8822_), .Y(new_n11800_));
  OR2X1    g10798(.A(new_n10003_), .B(new_n9623_), .Y(new_n11801_));
  AND2X1   g10799(.A(new_n11801_), .B(new_n11800_), .Y(new_n11802_));
  XOR2X1   g10800(.A(new_n11056_), .B(new_n11802_), .Y(new_n11803_));
  NOR2X1   g10801(.A(new_n11337_), .B(new_n11803_), .Y(new_n11804_));
  NAND2X1  g10802(.A(new_n11337_), .B(new_n11803_), .Y(new_n11805_));
  OAI21X1  g10803(.A0(new_n11804_), .A1(new_n10557_), .B0(new_n11805_), .Y(new_n11806_));
  XOR2X1   g10804(.A(new_n9100_), .B(new_n8857_), .Y(new_n11807_));
  OAI22X1  g10805(.A0(new_n11807_), .A1(new_n9226_), .B0(new_n8853_), .B1(new_n5640_), .Y(new_n11808_));
  NAND2X1  g10806(.A(new_n11064_), .B(new_n9101_), .Y(new_n11809_));
  INVX1    g10807(.A(new_n9021_), .Y(new_n11810_));
  XOR2X1   g10808(.A(new_n9084_), .B(new_n11810_), .Y(new_n11811_));
  AOI22X1  g10809(.A0(new_n9099_), .A1(new_n11811_), .B0(new_n8856_), .B1(new_n8855_), .Y(new_n11812_));
  NOR2X1   g10810(.A(new_n11070_), .B(new_n11069_), .Y(new_n11813_));
  OR2X1    g10811(.A(new_n11813_), .B(new_n11812_), .Y(new_n11814_));
  XOR2X1   g10812(.A(new_n11232_), .B(new_n11814_), .Y(new_n11815_));
  AOI22X1  g10813(.A0(new_n11334_), .A1(new_n11815_), .B0(new_n11809_), .B1(new_n11808_), .Y(new_n11816_));
  AOI21X1  g10814(.A0(new_n11235_), .A1(new_n9103_), .B0(new_n11237_), .Y(new_n11817_));
  XOR2X1   g10815(.A(new_n11333_), .B(new_n11817_), .Y(new_n11818_));
  OAI21X1  g10816(.A0(new_n11232_), .A1(new_n11072_), .B0(new_n11818_), .Y(new_n11819_));
  NOR2X1   g10817(.A(new_n11819_), .B(new_n11233_), .Y(new_n11820_));
  OR2X1    g10818(.A(new_n11820_), .B(new_n11816_), .Y(new_n11821_));
  OR2X1    g10819(.A(new_n11178_), .B(new_n11177_), .Y(new_n11822_));
  XOR2X1   g10820(.A(new_n11224_), .B(new_n11822_), .Y(new_n11823_));
  AOI22X1  g10821(.A0(new_n11823_), .A1(new_n11175_), .B0(new_n11071_), .B1(new_n11068_), .Y(new_n11824_));
  AND2X1   g10822(.A(new_n11168_), .B(new_n11075_), .Y(new_n11825_));
  OAI21X1  g10823(.A0(new_n11168_), .A1(new_n11075_), .B0(new_n11225_), .Y(new_n11826_));
  NOR2X1   g10824(.A(new_n11826_), .B(new_n11825_), .Y(new_n11827_));
  OR2X1    g10825(.A(new_n11827_), .B(new_n11824_), .Y(new_n11828_));
  NOR2X1   g10826(.A(new_n8894_), .B(new_n8885_), .Y(new_n11829_));
  OAI22X1  g10827(.A0(new_n8929_), .A1(new_n11829_), .B0(new_n9094_), .B1(new_n9089_), .Y(new_n11830_));
  OR4X1    g10828(.A(new_n11137_), .B(new_n11136_), .C(new_n8894_), .D(new_n8885_), .Y(new_n11831_));
  AND2X1   g10829(.A(new_n11831_), .B(new_n11830_), .Y(new_n11832_));
  XOR2X1   g10830(.A(new_n11166_), .B(new_n11832_), .Y(new_n11833_));
  OAI22X1  g10831(.A0(new_n11833_), .A1(new_n11131_), .B0(new_n11173_), .B1(new_n11172_), .Y(new_n11834_));
  OR2X1    g10832(.A(new_n11167_), .B(new_n11229_), .Y(new_n11835_));
  AND2X1   g10833(.A(new_n11835_), .B(new_n11834_), .Y(new_n11836_));
  AND2X1   g10834(.A(new_n11151_), .B(new_n11150_), .Y(new_n11837_));
  NAND3X1  g10835(.A(new_n11163_), .B(new_n11161_), .C(new_n11150_), .Y(new_n11838_));
  OAI21X1  g10836(.A0(new_n11159_), .A1(new_n11837_), .B0(new_n11838_), .Y(new_n11839_));
  OR2X1    g10837(.A(new_n11839_), .B(new_n11149_), .Y(new_n11840_));
  OAI21X1  g10838(.A0(new_n8891_), .A1(new_n8888_), .B0(new_n11146_), .Y(new_n11841_));
  OAI21X1  g10839(.A0(new_n11147_), .A1(new_n8883_), .B0(new_n11841_), .Y(new_n11842_));
  AOI21X1  g10840(.A0(new_n11142_), .A1(new_n8878_), .B0(new_n11144_), .Y(new_n11843_));
  AOI22X1  g10841(.A0(new_n11843_), .A1(new_n11841_), .B0(new_n11144_), .B1(new_n11842_), .Y(new_n11844_));
  OAI22X1  g10842(.A0(new_n11165_), .A1(new_n11844_), .B0(new_n11138_), .B1(new_n11135_), .Y(new_n11845_));
  OR2X1    g10843(.A(new_n11145_), .B(new_n11143_), .Y(new_n11846_));
  AND2X1   g10844(.A(new_n4266_), .B(new_n4265_), .Y(new_n11847_));
  NOR3X1   g10845(.A(new_n8910_), .B(new_n8908_), .C(new_n11847_), .Y(new_n11848_));
  OAI21X1  g10846(.A0(new_n8908_), .A1(new_n11847_), .B0(new_n8910_), .Y(new_n11849_));
  OAI21X1  g10847(.A0(new_n11848_), .A1(new_n8911_), .B0(new_n11849_), .Y(new_n11850_));
  NOR2X1   g10848(.A(new_n11850_), .B(new_n11155_), .Y(new_n11851_));
  AOI21X1  g10849(.A0(new_n11151_), .A1(new_n11150_), .B0(new_n11851_), .Y(new_n11852_));
  NAND2X1  g10850(.A(new_n11850_), .B(new_n11155_), .Y(new_n11853_));
  OAI21X1  g10851(.A0(new_n11145_), .A1(new_n11143_), .B0(new_n11853_), .Y(new_n11854_));
  AND2X1   g10852(.A(new_n11850_), .B(new_n11155_), .Y(new_n11855_));
  NOR2X1   g10853(.A(new_n11855_), .B(new_n11852_), .Y(new_n11856_));
  OAI22X1  g10854(.A0(new_n11856_), .A1(new_n11846_), .B0(new_n11854_), .B1(new_n11852_), .Y(new_n11857_));
  AOI21X1  g10855(.A0(new_n11845_), .A1(new_n11840_), .B0(new_n11857_), .Y(new_n11858_));
  AND2X1   g10856(.A(new_n11165_), .B(new_n11844_), .Y(new_n11859_));
  AOI22X1  g10857(.A0(new_n11839_), .A1(new_n11149_), .B0(new_n11831_), .B1(new_n11830_), .Y(new_n11860_));
  AND2X1   g10858(.A(new_n11144_), .B(new_n11842_), .Y(new_n11861_));
  OR2X1    g10859(.A(new_n11851_), .B(new_n11837_), .Y(new_n11862_));
  AOI21X1  g10860(.A0(new_n11144_), .A1(new_n11842_), .B0(new_n11855_), .Y(new_n11863_));
  OR2X1    g10861(.A(new_n11855_), .B(new_n11852_), .Y(new_n11864_));
  AOI22X1  g10862(.A0(new_n11864_), .A1(new_n11861_), .B0(new_n11863_), .B1(new_n11862_), .Y(new_n11865_));
  NOR3X1   g10863(.A(new_n11865_), .B(new_n11860_), .C(new_n11859_), .Y(new_n11866_));
  OR2X1    g10864(.A(new_n11866_), .B(new_n11858_), .Y(new_n11867_));
  AOI22X1  g10865(.A0(new_n11128_), .A1(new_n11121_), .B0(new_n11107_), .B1(new_n11097_), .Y(new_n11868_));
  AOI21X1  g10866(.A0(new_n11085_), .A1(new_n11081_), .B0(new_n11868_), .Y(new_n11869_));
  AOI22X1  g10867(.A0(new_n11127_), .A1(new_n11126_), .B0(new_n11125_), .B1(new_n11124_), .Y(new_n11870_));
  NAND3X1  g10868(.A(new_n11128_), .B(new_n11107_), .C(new_n11097_), .Y(new_n11871_));
  NOR2X1   g10869(.A(new_n11871_), .B(new_n11870_), .Y(new_n11872_));
  OR4X1    g10870(.A(new_n9012_), .B(new_n9006_), .C(new_n8999_), .D(new_n8994_), .Y(new_n11873_));
  AOI22X1  g10871(.A0(new_n11095_), .A1(new_n11092_), .B0(new_n11873_), .B1(new_n11100_), .Y(new_n11874_));
  NOR2X1   g10872(.A(new_n11095_), .B(new_n11092_), .Y(new_n11875_));
  NOR2X1   g10873(.A(new_n11875_), .B(new_n11874_), .Y(new_n11876_));
  OR2X1    g10874(.A(new_n11113_), .B(new_n8975_), .Y(new_n11877_));
  AND2X1   g10875(.A(new_n11114_), .B(new_n11877_), .Y(new_n11878_));
  AOI22X1  g10876(.A0(new_n11118_), .A1(new_n11878_), .B0(new_n11125_), .B1(new_n11124_), .Y(new_n11879_));
  AOI21X1  g10877(.A0(new_n11114_), .A1(new_n11877_), .B0(new_n11118_), .Y(new_n11880_));
  OR2X1    g10878(.A(new_n11880_), .B(new_n11879_), .Y(new_n11881_));
  NOR2X1   g10879(.A(new_n11881_), .B(new_n11876_), .Y(new_n11882_));
  AND2X1   g10880(.A(new_n11881_), .B(new_n11876_), .Y(new_n11883_));
  OAI22X1  g10881(.A0(new_n11883_), .A1(new_n11882_), .B0(new_n11872_), .B1(new_n11869_), .Y(new_n11884_));
  AND2X1   g10882(.A(new_n11107_), .B(new_n11097_), .Y(new_n11885_));
  OAI22X1  g10883(.A0(new_n11129_), .A1(new_n11885_), .B0(new_n11227_), .B1(new_n11226_), .Y(new_n11886_));
  NAND4X1  g10884(.A(new_n11128_), .B(new_n11121_), .C(new_n11107_), .D(new_n11097_), .Y(new_n11887_));
  OR2X1    g10885(.A(new_n11881_), .B(new_n11876_), .Y(new_n11888_));
  NAND2X1  g10886(.A(new_n11881_), .B(new_n11876_), .Y(new_n11889_));
  NAND4X1  g10887(.A(new_n11889_), .B(new_n11888_), .C(new_n11887_), .D(new_n11886_), .Y(new_n11890_));
  AND2X1   g10888(.A(new_n11890_), .B(new_n11884_), .Y(new_n11891_));
  XOR2X1   g10889(.A(new_n11891_), .B(new_n11867_), .Y(new_n11892_));
  NOR2X1   g10890(.A(new_n11892_), .B(new_n11836_), .Y(new_n11893_));
  AOI22X1  g10891(.A0(new_n11199_), .A1(new_n11198_), .B0(new_n11197_), .B1(new_n11196_), .Y(new_n11894_));
  NOR4X1   g10892(.A(new_n11193_), .B(new_n11192_), .C(new_n11183_), .D(new_n11182_), .Y(new_n11895_));
  AND2X1   g10893(.A(new_n11215_), .B(new_n11206_), .Y(new_n11896_));
  NOR4X1   g10894(.A(new_n11221_), .B(new_n11220_), .C(new_n11218_), .D(new_n11217_), .Y(new_n11897_));
  OAI22X1  g10895(.A0(new_n11897_), .A1(new_n11896_), .B0(new_n11895_), .B1(new_n11894_), .Y(new_n11898_));
  AND2X1   g10896(.A(new_n11898_), .B(new_n11822_), .Y(new_n11899_));
  OAI21X1  g10897(.A0(new_n11178_), .A1(new_n11177_), .B0(new_n11898_), .Y(new_n11900_));
  NAND4X1  g10898(.A(new_n11222_), .B(new_n11216_), .C(new_n11200_), .D(new_n11194_), .Y(new_n11901_));
  AND2X1   g10899(.A(new_n11901_), .B(new_n11900_), .Y(new_n11902_));
  AOI22X1  g10900(.A0(new_n11185_), .A1(new_n9073_), .B0(new_n9071_), .B1(new_n9070_), .Y(new_n11903_));
  AOI22X1  g10901(.A0(new_n11191_), .A1(new_n11903_), .B0(new_n11197_), .B1(new_n11196_), .Y(new_n11904_));
  NOR2X1   g10902(.A(new_n11191_), .B(new_n11903_), .Y(new_n11905_));
  NOR2X1   g10903(.A(new_n11905_), .B(new_n11904_), .Y(new_n11906_));
  NAND4X1  g10904(.A(new_n11213_), .B(new_n11212_), .C(new_n11209_), .D(new_n11208_), .Y(new_n11907_));
  AND2X1   g10905(.A(new_n11907_), .B(new_n11206_), .Y(new_n11908_));
  OR2X1    g10906(.A(new_n11214_), .B(new_n11210_), .Y(new_n11909_));
  INVX1    g10907(.A(new_n11909_), .Y(new_n11910_));
  OR2X1    g10908(.A(new_n11910_), .B(new_n11908_), .Y(new_n11911_));
  XOR2X1   g10909(.A(new_n11911_), .B(new_n11906_), .Y(new_n11912_));
  AOI21X1  g10910(.A0(new_n11907_), .A1(new_n11206_), .B0(new_n11910_), .Y(new_n11913_));
  NOR3X1   g10911(.A(new_n11913_), .B(new_n11905_), .C(new_n11904_), .Y(new_n11914_));
  OAI21X1  g10912(.A0(new_n11911_), .A1(new_n11906_), .B0(new_n11901_), .Y(new_n11915_));
  OR2X1    g10913(.A(new_n11915_), .B(new_n11914_), .Y(new_n11916_));
  OAI22X1  g10914(.A0(new_n11916_), .A1(new_n11899_), .B0(new_n11912_), .B1(new_n11902_), .Y(new_n11917_));
  AOI22X1  g10915(.A0(new_n11167_), .A1(new_n11229_), .B0(new_n11074_), .B1(new_n11073_), .Y(new_n11918_));
  NOR2X1   g10916(.A(new_n11167_), .B(new_n11229_), .Y(new_n11919_));
  OR2X1    g10917(.A(new_n11919_), .B(new_n11918_), .Y(new_n11920_));
  NAND2X1  g10918(.A(new_n11890_), .B(new_n11884_), .Y(new_n11921_));
  XOR2X1   g10919(.A(new_n11921_), .B(new_n11867_), .Y(new_n11922_));
  OAI21X1  g10920(.A0(new_n11922_), .A1(new_n11920_), .B0(new_n11917_), .Y(new_n11923_));
  XOR2X1   g10921(.A(new_n11892_), .B(new_n11836_), .Y(new_n11924_));
  OAI22X1  g10922(.A0(new_n11924_), .A1(new_n11917_), .B0(new_n11923_), .B1(new_n11893_), .Y(new_n11925_));
  AND2X1   g10923(.A(new_n11925_), .B(new_n11828_), .Y(new_n11926_));
  AND2X1   g10924(.A(new_n11287_), .B(new_n11286_), .Y(new_n11927_));
  OR2X1    g10925(.A(new_n11288_), .B(new_n11927_), .Y(new_n11928_));
  XOR2X1   g10926(.A(new_n11331_), .B(new_n11928_), .Y(new_n11929_));
  AOI21X1  g10927(.A0(new_n11929_), .A1(new_n11285_), .B0(new_n11817_), .Y(new_n11930_));
  AOI21X1  g10928(.A0(new_n11239_), .A1(new_n11059_), .B0(new_n11241_), .Y(new_n11931_));
  XOR2X1   g10929(.A(new_n11284_), .B(new_n11931_), .Y(new_n11932_));
  AND2X1   g10930(.A(new_n11332_), .B(new_n11932_), .Y(new_n11933_));
  OR2X1    g10931(.A(new_n11933_), .B(new_n11930_), .Y(new_n11934_));
  AOI22X1  g10932(.A0(new_n11329_), .A1(new_n11324_), .B0(new_n11309_), .B1(new_n11304_), .Y(new_n11935_));
  NAND4X1  g10933(.A(new_n11329_), .B(new_n11324_), .C(new_n11309_), .D(new_n11304_), .Y(new_n11936_));
  OAI21X1  g10934(.A0(new_n11935_), .A1(new_n11289_), .B0(new_n11936_), .Y(new_n11937_));
  AND2X1   g10935(.A(new_n11298_), .B(new_n11297_), .Y(new_n11938_));
  AOI21X1  g10936(.A0(new_n11302_), .A1(new_n11938_), .B0(new_n11295_), .Y(new_n11939_));
  NOR2X1   g10937(.A(new_n11302_), .B(new_n11938_), .Y(new_n11940_));
  OR2X1    g10938(.A(new_n11940_), .B(new_n11939_), .Y(new_n11941_));
  NAND2X1  g10939(.A(new_n11322_), .B(new_n11319_), .Y(new_n11942_));
  AND2X1   g10940(.A(new_n11942_), .B(new_n11315_), .Y(new_n11943_));
  NOR2X1   g10941(.A(new_n11322_), .B(new_n11319_), .Y(new_n11944_));
  OR2X1    g10942(.A(new_n11944_), .B(new_n11943_), .Y(new_n11945_));
  XOR2X1   g10943(.A(new_n11945_), .B(new_n11941_), .Y(new_n11946_));
  NAND2X1  g10944(.A(new_n11946_), .B(new_n11937_), .Y(new_n11947_));
  NOR2X1   g10945(.A(new_n11935_), .B(new_n11289_), .Y(new_n11948_));
  NAND3X1  g10946(.A(new_n11329_), .B(new_n11309_), .C(new_n11304_), .Y(new_n11949_));
  AOI21X1  g10947(.A0(new_n11323_), .A1(new_n11315_), .B0(new_n11949_), .Y(new_n11950_));
  AOI21X1  g10948(.A0(new_n11942_), .A1(new_n11315_), .B0(new_n11944_), .Y(new_n11951_));
  AND2X1   g10949(.A(new_n11951_), .B(new_n11941_), .Y(new_n11952_));
  NOR3X1   g10950(.A(new_n11951_), .B(new_n11940_), .C(new_n11939_), .Y(new_n11953_));
  OR4X1    g10951(.A(new_n11953_), .B(new_n11952_), .C(new_n11950_), .D(new_n11948_), .Y(new_n11954_));
  NAND2X1  g10952(.A(new_n11954_), .B(new_n11947_), .Y(new_n11955_));
  AOI22X1  g10953(.A0(new_n11282_), .A1(new_n11277_), .B0(new_n11262_), .B1(new_n11257_), .Y(new_n11956_));
  NAND4X1  g10954(.A(new_n11282_), .B(new_n11277_), .C(new_n11262_), .D(new_n11257_), .Y(new_n11957_));
  OAI21X1  g10955(.A0(new_n11956_), .A1(new_n11931_), .B0(new_n11957_), .Y(new_n11958_));
  AND2X1   g10956(.A(new_n11251_), .B(new_n11250_), .Y(new_n11959_));
  AOI21X1  g10957(.A0(new_n11255_), .A1(new_n11959_), .B0(new_n11248_), .Y(new_n11960_));
  NOR2X1   g10958(.A(new_n11255_), .B(new_n11959_), .Y(new_n11961_));
  OR2X1    g10959(.A(new_n11961_), .B(new_n11960_), .Y(new_n11962_));
  NAND2X1  g10960(.A(new_n11275_), .B(new_n11272_), .Y(new_n11963_));
  AND2X1   g10961(.A(new_n11963_), .B(new_n11268_), .Y(new_n11964_));
  NOR2X1   g10962(.A(new_n11275_), .B(new_n11272_), .Y(new_n11965_));
  OR2X1    g10963(.A(new_n11965_), .B(new_n11964_), .Y(new_n11966_));
  XOR2X1   g10964(.A(new_n11966_), .B(new_n11962_), .Y(new_n11967_));
  NAND2X1  g10965(.A(new_n11967_), .B(new_n11958_), .Y(new_n11968_));
  NOR2X1   g10966(.A(new_n11956_), .B(new_n11931_), .Y(new_n11969_));
  NAND3X1  g10967(.A(new_n11282_), .B(new_n11262_), .C(new_n11257_), .Y(new_n11970_));
  AOI21X1  g10968(.A0(new_n11276_), .A1(new_n11268_), .B0(new_n11970_), .Y(new_n11971_));
  AOI21X1  g10969(.A0(new_n11963_), .A1(new_n11268_), .B0(new_n11965_), .Y(new_n11972_));
  AND2X1   g10970(.A(new_n11972_), .B(new_n11962_), .Y(new_n11973_));
  NOR3X1   g10971(.A(new_n11972_), .B(new_n11961_), .C(new_n11960_), .Y(new_n11974_));
  OR4X1    g10972(.A(new_n11974_), .B(new_n11973_), .C(new_n11971_), .D(new_n11969_), .Y(new_n11975_));
  AND2X1   g10973(.A(new_n11975_), .B(new_n11968_), .Y(new_n11976_));
  XOR2X1   g10974(.A(new_n11976_), .B(new_n11955_), .Y(new_n11977_));
  XOR2X1   g10975(.A(new_n11977_), .B(new_n11934_), .Y(new_n11978_));
  OAI21X1  g10976(.A0(new_n11925_), .A1(new_n11828_), .B0(new_n11978_), .Y(new_n11979_));
  XOR2X1   g10977(.A(new_n11925_), .B(new_n11828_), .Y(new_n11980_));
  OAI22X1  g10978(.A0(new_n11980_), .A1(new_n11978_), .B0(new_n11979_), .B1(new_n11926_), .Y(new_n11981_));
  XOR2X1   g10979(.A(new_n11981_), .B(new_n11821_), .Y(new_n11982_));
  OR2X1    g10980(.A(new_n10683_), .B(new_n10682_), .Y(new_n11983_));
  XOR2X1   g10981(.A(new_n9817_), .B(new_n11983_), .Y(new_n11984_));
  AND2X1   g10982(.A(new_n10566_), .B(new_n10565_), .Y(new_n11985_));
  XOR2X1   g10983(.A(new_n10000_), .B(new_n11985_), .Y(new_n11986_));
  OAI22X1  g10984(.A0(new_n11986_), .A1(new_n11984_), .B0(new_n11797_), .B1(new_n11796_), .Y(new_n11987_));
  OR2X1    g10985(.A(new_n10001_), .B(new_n9818_), .Y(new_n11988_));
  AND2X1   g10986(.A(new_n11988_), .B(new_n11987_), .Y(new_n11989_));
  XOR2X1   g10987(.A(new_n10805_), .B(new_n11989_), .Y(new_n11990_));
  OAI22X1  g10988(.A0(new_n11055_), .A1(new_n11990_), .B0(new_n10560_), .B1(new_n10559_), .Y(new_n11991_));
  NAND2X1  g10989(.A(new_n11055_), .B(new_n11990_), .Y(new_n11992_));
  AND2X1   g10990(.A(new_n11992_), .B(new_n11991_), .Y(new_n11993_));
  AOI22X1  g10991(.A0(new_n9436_), .A1(new_n9351_), .B0(new_n9258_), .B1(new_n9248_), .Y(new_n11994_));
  NOR2X1   g10992(.A(new_n9436_), .B(new_n9351_), .Y(new_n11995_));
  OR2X1    g10993(.A(new_n11995_), .B(new_n11994_), .Y(new_n11996_));
  XOR2X1   g10994(.A(new_n11052_), .B(new_n11996_), .Y(new_n11997_));
  AOI22X1  g10995(.A0(new_n11997_), .A1(new_n10934_), .B0(new_n10818_), .B1(new_n10817_), .Y(new_n11998_));
  OR2X1    g10996(.A(new_n5910_), .B(new_n6010_), .Y(new_n11999_));
  OAI21X1  g10997(.A0(new_n9448_), .A1(new_n5923_), .B0(new_n6006_), .Y(new_n12000_));
  OAI22X1  g10998(.A0(new_n9449_), .A1(new_n6006_), .B0(new_n12000_), .B1(new_n9451_), .Y(new_n12001_));
  OAI22X1  g10999(.A0(new_n9462_), .A1(new_n9451_), .B0(new_n9449_), .B1(new_n5940_), .Y(new_n12002_));
  MX2X1    g11000(.A(new_n12002_), .B(new_n12001_), .S0(new_n6005_), .Y(new_n12003_));
  OAI21X1  g11001(.A0(new_n6011_), .A1(new_n5808_), .B0(new_n12003_), .Y(new_n12004_));
  AND2X1   g11002(.A(new_n12004_), .B(new_n11999_), .Y(new_n12005_));
  XOR2X1   g11003(.A(new_n9532_), .B(new_n12005_), .Y(new_n12006_));
  OAI22X1  g11004(.A0(new_n9619_), .A1(new_n12006_), .B0(new_n9440_), .B1(new_n9439_), .Y(new_n12007_));
  OR2X1    g11005(.A(new_n10823_), .B(new_n9533_), .Y(new_n12008_));
  AND2X1   g11006(.A(new_n12008_), .B(new_n12007_), .Y(new_n12009_));
  XOR2X1   g11007(.A(new_n10933_), .B(new_n12009_), .Y(new_n12010_));
  AND2X1   g11008(.A(new_n11053_), .B(new_n12010_), .Y(new_n12011_));
  OR2X1    g11009(.A(new_n12011_), .B(new_n11998_), .Y(new_n12012_));
  AOI22X1  g11010(.A0(new_n11006_), .A1(new_n9314_), .B0(new_n10940_), .B1(new_n10935_), .Y(new_n12013_));
  NOR2X1   g11011(.A(new_n11006_), .B(new_n9314_), .Y(new_n12014_));
  OR2X1    g11012(.A(new_n12014_), .B(new_n12013_), .Y(new_n12015_));
  XOR2X1   g11013(.A(new_n11050_), .B(new_n12015_), .Y(new_n12016_));
  AOI22X1  g11014(.A0(new_n12016_), .A1(new_n10999_), .B0(new_n10948_), .B1(new_n10947_), .Y(new_n12017_));
  XOR2X1   g11015(.A(new_n9397_), .B(new_n10976_), .Y(new_n12018_));
  XOR2X1   g11016(.A(new_n12018_), .B(new_n9367_), .Y(new_n12019_));
  OAI22X1  g11017(.A0(new_n9434_), .A1(new_n12019_), .B0(new_n9353_), .B1(new_n9352_), .Y(new_n12020_));
  OR2X1    g11018(.A(new_n10952_), .B(new_n9399_), .Y(new_n12021_));
  AND2X1   g11019(.A(new_n12021_), .B(new_n12020_), .Y(new_n12022_));
  XOR2X1   g11020(.A(new_n10998_), .B(new_n12022_), .Y(new_n12023_));
  AND2X1   g11021(.A(new_n11051_), .B(new_n12023_), .Y(new_n12024_));
  OR2X1    g11022(.A(new_n12024_), .B(new_n12017_), .Y(new_n12025_));
  AOI22X1  g11023(.A0(new_n11048_), .A1(new_n11040_), .B0(new_n11027_), .B1(new_n11020_), .Y(new_n12026_));
  AOI21X1  g11024(.A0(new_n11007_), .A1(new_n11003_), .B0(new_n12026_), .Y(new_n12027_));
  AOI22X1  g11025(.A0(new_n11047_), .A1(new_n11046_), .B0(new_n11044_), .B1(new_n11043_), .Y(new_n12028_));
  NAND3X1  g11026(.A(new_n11048_), .B(new_n11027_), .C(new_n11020_), .Y(new_n12029_));
  NOR2X1   g11027(.A(new_n12029_), .B(new_n12028_), .Y(new_n12030_));
  OR4X1    g11028(.A(new_n9346_), .B(new_n9340_), .C(new_n9333_), .D(new_n9328_), .Y(new_n12031_));
  AOI22X1  g11029(.A0(new_n11018_), .A1(new_n11015_), .B0(new_n12031_), .B1(new_n11023_), .Y(new_n12032_));
  NOR2X1   g11030(.A(new_n11018_), .B(new_n11015_), .Y(new_n12033_));
  OR2X1    g11031(.A(new_n12033_), .B(new_n12032_), .Y(new_n12034_));
  AOI22X1  g11032(.A0(new_n11038_), .A1(new_n11035_), .B0(new_n11044_), .B1(new_n11043_), .Y(new_n12035_));
  NOR2X1   g11033(.A(new_n11038_), .B(new_n11035_), .Y(new_n12036_));
  OR2X1    g11034(.A(new_n12036_), .B(new_n12035_), .Y(new_n12037_));
  XOR2X1   g11035(.A(new_n12037_), .B(new_n12034_), .Y(new_n12038_));
  OAI21X1  g11036(.A0(new_n12030_), .A1(new_n12027_), .B0(new_n12038_), .Y(new_n12039_));
  AND2X1   g11037(.A(new_n11027_), .B(new_n11020_), .Y(new_n12040_));
  OAI22X1  g11038(.A0(new_n11049_), .A1(new_n12040_), .B0(new_n12014_), .B1(new_n12013_), .Y(new_n12041_));
  NAND4X1  g11039(.A(new_n11048_), .B(new_n11040_), .C(new_n11027_), .D(new_n11020_), .Y(new_n12042_));
  NOR2X1   g11040(.A(new_n12036_), .B(new_n12035_), .Y(new_n12043_));
  NAND2X1  g11041(.A(new_n12043_), .B(new_n12034_), .Y(new_n12044_));
  OR2X1    g11042(.A(new_n12043_), .B(new_n12034_), .Y(new_n12045_));
  NAND4X1  g11043(.A(new_n12045_), .B(new_n12044_), .C(new_n12042_), .D(new_n12041_), .Y(new_n12046_));
  NAND2X1  g11044(.A(new_n12046_), .B(new_n12039_), .Y(new_n12047_));
  AOI22X1  g11045(.A0(new_n10996_), .A1(new_n10988_), .B0(new_n10974_), .B1(new_n10967_), .Y(new_n12048_));
  AOI21X1  g11046(.A0(new_n12021_), .A1(new_n12020_), .B0(new_n12048_), .Y(new_n12049_));
  AOI22X1  g11047(.A0(new_n10995_), .A1(new_n10994_), .B0(new_n10992_), .B1(new_n10991_), .Y(new_n12050_));
  NAND3X1  g11048(.A(new_n10996_), .B(new_n10974_), .C(new_n10967_), .Y(new_n12051_));
  NOR2X1   g11049(.A(new_n12051_), .B(new_n12050_), .Y(new_n12052_));
  OR4X1    g11050(.A(new_n9431_), .B(new_n9425_), .C(new_n9418_), .D(new_n9413_), .Y(new_n12053_));
  AOI22X1  g11051(.A0(new_n10965_), .A1(new_n10962_), .B0(new_n12053_), .B1(new_n10970_), .Y(new_n12054_));
  NOR2X1   g11052(.A(new_n10965_), .B(new_n10962_), .Y(new_n12055_));
  OR2X1    g11053(.A(new_n12055_), .B(new_n12054_), .Y(new_n12056_));
  AOI22X1  g11054(.A0(new_n10986_), .A1(new_n10983_), .B0(new_n10992_), .B1(new_n10991_), .Y(new_n12057_));
  NOR2X1   g11055(.A(new_n10986_), .B(new_n10983_), .Y(new_n12058_));
  OR2X1    g11056(.A(new_n12058_), .B(new_n12057_), .Y(new_n12059_));
  XOR2X1   g11057(.A(new_n12059_), .B(new_n12056_), .Y(new_n12060_));
  OAI21X1  g11058(.A0(new_n12052_), .A1(new_n12049_), .B0(new_n12060_), .Y(new_n12061_));
  AND2X1   g11059(.A(new_n10974_), .B(new_n10967_), .Y(new_n12062_));
  OAI22X1  g11060(.A0(new_n10997_), .A1(new_n12062_), .B0(new_n10954_), .B1(new_n10953_), .Y(new_n12063_));
  NAND4X1  g11061(.A(new_n10996_), .B(new_n10988_), .C(new_n10974_), .D(new_n10967_), .Y(new_n12064_));
  NOR2X1   g11062(.A(new_n12058_), .B(new_n12057_), .Y(new_n12065_));
  NAND2X1  g11063(.A(new_n12065_), .B(new_n12056_), .Y(new_n12066_));
  OR2X1    g11064(.A(new_n12065_), .B(new_n12056_), .Y(new_n12067_));
  NAND4X1  g11065(.A(new_n12067_), .B(new_n12066_), .C(new_n12064_), .D(new_n12063_), .Y(new_n12068_));
  AND2X1   g11066(.A(new_n12068_), .B(new_n12061_), .Y(new_n12069_));
  XOR2X1   g11067(.A(new_n12069_), .B(new_n12047_), .Y(new_n12070_));
  XOR2X1   g11068(.A(new_n12070_), .B(new_n12025_), .Y(new_n12071_));
  XOR2X1   g11069(.A(new_n9580_), .B(new_n10855_), .Y(new_n12072_));
  XOR2X1   g11070(.A(new_n12072_), .B(new_n9549_), .Y(new_n12073_));
  OAI22X1  g11071(.A0(new_n9617_), .A1(new_n12073_), .B0(new_n10821_), .B1(new_n10820_), .Y(new_n12074_));
  OR2X1    g11072(.A(new_n10829_), .B(new_n9582_), .Y(new_n12075_));
  AND2X1   g11073(.A(new_n12075_), .B(new_n12074_), .Y(new_n12076_));
  XOR2X1   g11074(.A(new_n10877_), .B(new_n12076_), .Y(new_n12077_));
  OAI22X1  g11075(.A0(new_n10932_), .A1(new_n12077_), .B0(new_n10825_), .B1(new_n10824_), .Y(new_n12078_));
  NAND2X1  g11076(.A(new_n10932_), .B(new_n12077_), .Y(new_n12079_));
  AND2X1   g11077(.A(new_n12079_), .B(new_n12078_), .Y(new_n12080_));
  AOI22X1  g11078(.A0(new_n10929_), .A1(new_n10921_), .B0(new_n10908_), .B1(new_n10898_), .Y(new_n12081_));
  AOI21X1  g11079(.A0(new_n10886_), .A1(new_n10882_), .B0(new_n12081_), .Y(new_n12082_));
  AOI22X1  g11080(.A0(new_n10928_), .A1(new_n10927_), .B0(new_n10925_), .B1(new_n10924_), .Y(new_n12083_));
  NAND3X1  g11081(.A(new_n10929_), .B(new_n10908_), .C(new_n10898_), .Y(new_n12084_));
  NOR2X1   g11082(.A(new_n12084_), .B(new_n12083_), .Y(new_n12085_));
  OR4X1    g11083(.A(new_n9528_), .B(new_n9522_), .C(new_n9515_), .D(new_n9510_), .Y(new_n12086_));
  AOI22X1  g11084(.A0(new_n10896_), .A1(new_n10893_), .B0(new_n12086_), .B1(new_n10901_), .Y(new_n12087_));
  NOR2X1   g11085(.A(new_n10896_), .B(new_n10893_), .Y(new_n12088_));
  NOR2X1   g11086(.A(new_n12088_), .B(new_n12087_), .Y(new_n12089_));
  AOI22X1  g11087(.A0(new_n10919_), .A1(new_n10916_), .B0(new_n10925_), .B1(new_n10924_), .Y(new_n12090_));
  NOR2X1   g11088(.A(new_n10919_), .B(new_n10916_), .Y(new_n12091_));
  OR2X1    g11089(.A(new_n12091_), .B(new_n12090_), .Y(new_n12092_));
  NOR2X1   g11090(.A(new_n12092_), .B(new_n12089_), .Y(new_n12093_));
  AND2X1   g11091(.A(new_n12092_), .B(new_n12089_), .Y(new_n12094_));
  OAI22X1  g11092(.A0(new_n12094_), .A1(new_n12093_), .B0(new_n12085_), .B1(new_n12082_), .Y(new_n12095_));
  AOI22X1  g11093(.A0(new_n10885_), .A1(new_n9496_), .B0(new_n12004_), .B1(new_n11999_), .Y(new_n12096_));
  NOR2X1   g11094(.A(new_n10885_), .B(new_n9496_), .Y(new_n12097_));
  AND2X1   g11095(.A(new_n10908_), .B(new_n10898_), .Y(new_n12098_));
  OAI22X1  g11096(.A0(new_n10930_), .A1(new_n12098_), .B0(new_n12097_), .B1(new_n12096_), .Y(new_n12099_));
  NAND4X1  g11097(.A(new_n10929_), .B(new_n10921_), .C(new_n10908_), .D(new_n10898_), .Y(new_n12100_));
  OR2X1    g11098(.A(new_n12092_), .B(new_n12089_), .Y(new_n12101_));
  NAND2X1  g11099(.A(new_n12092_), .B(new_n12089_), .Y(new_n12102_));
  NAND4X1  g11100(.A(new_n12102_), .B(new_n12101_), .C(new_n12100_), .D(new_n12099_), .Y(new_n12103_));
  NAND2X1  g11101(.A(new_n12103_), .B(new_n12095_), .Y(new_n12104_));
  AOI22X1  g11102(.A0(new_n10875_), .A1(new_n10868_), .B0(new_n10853_), .B1(new_n10843_), .Y(new_n12105_));
  AOI21X1  g11103(.A0(new_n12075_), .A1(new_n12074_), .B0(new_n12105_), .Y(new_n12106_));
  AOI22X1  g11104(.A0(new_n10874_), .A1(new_n10873_), .B0(new_n10872_), .B1(new_n10871_), .Y(new_n12107_));
  NAND3X1  g11105(.A(new_n10875_), .B(new_n10853_), .C(new_n10843_), .Y(new_n12108_));
  NOR2X1   g11106(.A(new_n12108_), .B(new_n12107_), .Y(new_n12109_));
  OR4X1    g11107(.A(new_n9614_), .B(new_n9608_), .C(new_n9601_), .D(new_n9596_), .Y(new_n12110_));
  AOI22X1  g11108(.A0(new_n10841_), .A1(new_n10838_), .B0(new_n12110_), .B1(new_n10846_), .Y(new_n12111_));
  NOR2X1   g11109(.A(new_n10841_), .B(new_n10838_), .Y(new_n12112_));
  NOR2X1   g11110(.A(new_n12112_), .B(new_n12111_), .Y(new_n12113_));
  OR2X1    g11111(.A(new_n10860_), .B(new_n9577_), .Y(new_n12114_));
  AND2X1   g11112(.A(new_n10861_), .B(new_n12114_), .Y(new_n12115_));
  AOI22X1  g11113(.A0(new_n10865_), .A1(new_n12115_), .B0(new_n10872_), .B1(new_n10871_), .Y(new_n12116_));
  AOI21X1  g11114(.A0(new_n10861_), .A1(new_n12114_), .B0(new_n10865_), .Y(new_n12117_));
  OR2X1    g11115(.A(new_n12117_), .B(new_n12116_), .Y(new_n12118_));
  NOR2X1   g11116(.A(new_n12118_), .B(new_n12113_), .Y(new_n12119_));
  AND2X1   g11117(.A(new_n12118_), .B(new_n12113_), .Y(new_n12120_));
  OAI22X1  g11118(.A0(new_n12120_), .A1(new_n12119_), .B0(new_n12109_), .B1(new_n12106_), .Y(new_n12121_));
  AND2X1   g11119(.A(new_n10853_), .B(new_n10843_), .Y(new_n12122_));
  OAI22X1  g11120(.A0(new_n10876_), .A1(new_n12122_), .B0(new_n10831_), .B1(new_n10830_), .Y(new_n12123_));
  NAND4X1  g11121(.A(new_n10875_), .B(new_n10868_), .C(new_n10853_), .D(new_n10843_), .Y(new_n12124_));
  OR2X1    g11122(.A(new_n12118_), .B(new_n12113_), .Y(new_n12125_));
  NAND2X1  g11123(.A(new_n12118_), .B(new_n12113_), .Y(new_n12126_));
  NAND4X1  g11124(.A(new_n12126_), .B(new_n12125_), .C(new_n12124_), .D(new_n12123_), .Y(new_n12127_));
  AND2X1   g11125(.A(new_n12127_), .B(new_n12121_), .Y(new_n12128_));
  XOR2X1   g11126(.A(new_n12128_), .B(new_n12104_), .Y(new_n12129_));
  XOR2X1   g11127(.A(new_n12129_), .B(new_n12080_), .Y(new_n12130_));
  XOR2X1   g11128(.A(new_n12130_), .B(new_n12071_), .Y(new_n12131_));
  XOR2X1   g11129(.A(new_n12131_), .B(new_n12012_), .Y(new_n12132_));
  OR2X1    g11130(.A(new_n8735_), .B(new_n8217_), .Y(new_n12133_));
  OAI21X1  g11131(.A0(new_n9828_), .A1(new_n8243_), .B0(new_n8326_), .Y(new_n12134_));
  OAI22X1  g11132(.A0(new_n9829_), .A1(new_n8326_), .B0(new_n12134_), .B1(new_n9831_), .Y(new_n12135_));
  OAI22X1  g11133(.A0(new_n9842_), .A1(new_n9831_), .B0(new_n9829_), .B1(new_n8260_), .Y(new_n12136_));
  MX2X1    g11134(.A(new_n12136_), .B(new_n12135_), .S0(new_n8325_), .Y(new_n12137_));
  OAI21X1  g11135(.A0(new_n8737_), .A1(new_n8731_), .B0(new_n12137_), .Y(new_n12138_));
  AND2X1   g11136(.A(new_n12138_), .B(new_n12133_), .Y(new_n12139_));
  XOR2X1   g11137(.A(new_n9912_), .B(new_n12139_), .Y(new_n12140_));
  OAI22X1  g11138(.A0(new_n9999_), .A1(new_n12140_), .B0(new_n9820_), .B1(new_n9819_), .Y(new_n12141_));
  OR2X1    g11139(.A(new_n10570_), .B(new_n9913_), .Y(new_n12142_));
  AND2X1   g11140(.A(new_n12142_), .B(new_n12141_), .Y(new_n12143_));
  XOR2X1   g11141(.A(new_n10680_), .B(new_n12143_), .Y(new_n12144_));
  OAI22X1  g11142(.A0(new_n10804_), .A1(new_n12144_), .B0(new_n10563_), .B1(new_n10562_), .Y(new_n12145_));
  NAND2X1  g11143(.A(new_n10804_), .B(new_n12144_), .Y(new_n12146_));
  AND2X1   g11144(.A(new_n12146_), .B(new_n12145_), .Y(new_n12147_));
  AOI22X1  g11145(.A0(new_n10757_), .A1(new_n9693_), .B0(new_n10689_), .B1(new_n10684_), .Y(new_n12148_));
  NOR2X1   g11146(.A(new_n10757_), .B(new_n9693_), .Y(new_n12149_));
  OR2X1    g11147(.A(new_n12149_), .B(new_n12148_), .Y(new_n12150_));
  XOR2X1   g11148(.A(new_n10801_), .B(new_n12150_), .Y(new_n12151_));
  AOI22X1  g11149(.A0(new_n12151_), .A1(new_n10750_), .B0(new_n10697_), .B1(new_n10696_), .Y(new_n12152_));
  XOR2X1   g11150(.A(new_n9777_), .B(new_n10727_), .Y(new_n12153_));
  XOR2X1   g11151(.A(new_n12153_), .B(new_n9746_), .Y(new_n12154_));
  OAI22X1  g11152(.A0(new_n9814_), .A1(new_n12154_), .B0(new_n9732_), .B1(new_n9731_), .Y(new_n12155_));
  OR2X1    g11153(.A(new_n10701_), .B(new_n9779_), .Y(new_n12156_));
  AND2X1   g11154(.A(new_n12156_), .B(new_n12155_), .Y(new_n12157_));
  XOR2X1   g11155(.A(new_n10749_), .B(new_n12157_), .Y(new_n12158_));
  AND2X1   g11156(.A(new_n10802_), .B(new_n12158_), .Y(new_n12159_));
  OR2X1    g11157(.A(new_n12159_), .B(new_n12152_), .Y(new_n12160_));
  AOI22X1  g11158(.A0(new_n10799_), .A1(new_n10791_), .B0(new_n10778_), .B1(new_n10771_), .Y(new_n12161_));
  AOI21X1  g11159(.A0(new_n10758_), .A1(new_n10754_), .B0(new_n12161_), .Y(new_n12162_));
  AOI22X1  g11160(.A0(new_n10798_), .A1(new_n10797_), .B0(new_n10795_), .B1(new_n10794_), .Y(new_n12163_));
  NAND3X1  g11161(.A(new_n10799_), .B(new_n10778_), .C(new_n10771_), .Y(new_n12164_));
  NOR2X1   g11162(.A(new_n12164_), .B(new_n12163_), .Y(new_n12165_));
  OR4X1    g11163(.A(new_n9725_), .B(new_n9719_), .C(new_n9712_), .D(new_n9707_), .Y(new_n12166_));
  AOI22X1  g11164(.A0(new_n10769_), .A1(new_n10766_), .B0(new_n12166_), .B1(new_n10774_), .Y(new_n12167_));
  NOR2X1   g11165(.A(new_n10769_), .B(new_n10766_), .Y(new_n12168_));
  OR2X1    g11166(.A(new_n12168_), .B(new_n12167_), .Y(new_n12169_));
  AOI22X1  g11167(.A0(new_n10789_), .A1(new_n10786_), .B0(new_n10795_), .B1(new_n10794_), .Y(new_n12170_));
  NOR2X1   g11168(.A(new_n10789_), .B(new_n10786_), .Y(new_n12171_));
  OR2X1    g11169(.A(new_n12171_), .B(new_n12170_), .Y(new_n12172_));
  XOR2X1   g11170(.A(new_n12172_), .B(new_n12169_), .Y(new_n12173_));
  OAI21X1  g11171(.A0(new_n12165_), .A1(new_n12162_), .B0(new_n12173_), .Y(new_n12174_));
  NOR2X1   g11172(.A(new_n12171_), .B(new_n12170_), .Y(new_n12175_));
  AND2X1   g11173(.A(new_n12175_), .B(new_n12169_), .Y(new_n12176_));
  NOR2X1   g11174(.A(new_n12175_), .B(new_n12169_), .Y(new_n12177_));
  OR4X1    g11175(.A(new_n12177_), .B(new_n12176_), .C(new_n12165_), .D(new_n12162_), .Y(new_n12178_));
  NAND2X1  g11176(.A(new_n12178_), .B(new_n12174_), .Y(new_n12179_));
  AOI22X1  g11177(.A0(new_n10747_), .A1(new_n10740_), .B0(new_n10725_), .B1(new_n10715_), .Y(new_n12180_));
  AOI21X1  g11178(.A0(new_n12156_), .A1(new_n12155_), .B0(new_n12180_), .Y(new_n12181_));
  AOI22X1  g11179(.A0(new_n10746_), .A1(new_n10745_), .B0(new_n10744_), .B1(new_n10743_), .Y(new_n12182_));
  NAND3X1  g11180(.A(new_n10747_), .B(new_n10725_), .C(new_n10715_), .Y(new_n12183_));
  NOR2X1   g11181(.A(new_n12183_), .B(new_n12182_), .Y(new_n12184_));
  OR4X1    g11182(.A(new_n9811_), .B(new_n9805_), .C(new_n9798_), .D(new_n9793_), .Y(new_n12185_));
  AOI22X1  g11183(.A0(new_n10713_), .A1(new_n10710_), .B0(new_n12185_), .B1(new_n10718_), .Y(new_n12186_));
  NOR2X1   g11184(.A(new_n10713_), .B(new_n10710_), .Y(new_n12187_));
  NOR2X1   g11185(.A(new_n12187_), .B(new_n12186_), .Y(new_n12188_));
  OR2X1    g11186(.A(new_n10732_), .B(new_n9774_), .Y(new_n12189_));
  AND2X1   g11187(.A(new_n10733_), .B(new_n12189_), .Y(new_n12190_));
  AOI22X1  g11188(.A0(new_n10737_), .A1(new_n12190_), .B0(new_n10744_), .B1(new_n10743_), .Y(new_n12191_));
  AOI21X1  g11189(.A0(new_n10733_), .A1(new_n12189_), .B0(new_n10737_), .Y(new_n12192_));
  OR2X1    g11190(.A(new_n12192_), .B(new_n12191_), .Y(new_n12193_));
  NOR2X1   g11191(.A(new_n12193_), .B(new_n12188_), .Y(new_n12194_));
  AND2X1   g11192(.A(new_n12193_), .B(new_n12188_), .Y(new_n12195_));
  OAI22X1  g11193(.A0(new_n12195_), .A1(new_n12194_), .B0(new_n12184_), .B1(new_n12181_), .Y(new_n12196_));
  AND2X1   g11194(.A(new_n10725_), .B(new_n10715_), .Y(new_n12197_));
  OAI22X1  g11195(.A0(new_n10748_), .A1(new_n12197_), .B0(new_n10703_), .B1(new_n10702_), .Y(new_n12198_));
  NAND4X1  g11196(.A(new_n10747_), .B(new_n10740_), .C(new_n10725_), .D(new_n10715_), .Y(new_n12199_));
  OR2X1    g11197(.A(new_n12193_), .B(new_n12188_), .Y(new_n12200_));
  NAND2X1  g11198(.A(new_n12193_), .B(new_n12188_), .Y(new_n12201_));
  NAND4X1  g11199(.A(new_n12201_), .B(new_n12200_), .C(new_n12199_), .D(new_n12198_), .Y(new_n12202_));
  AND2X1   g11200(.A(new_n12202_), .B(new_n12196_), .Y(new_n12203_));
  XOR2X1   g11201(.A(new_n12203_), .B(new_n12179_), .Y(new_n12204_));
  XOR2X1   g11202(.A(new_n12204_), .B(new_n12160_), .Y(new_n12205_));
  XOR2X1   g11203(.A(new_n9960_), .B(new_n10602_), .Y(new_n12206_));
  XOR2X1   g11204(.A(new_n12206_), .B(new_n9929_), .Y(new_n12207_));
  OAI22X1  g11205(.A0(new_n9997_), .A1(new_n12207_), .B0(new_n10568_), .B1(new_n10567_), .Y(new_n12208_));
  OR2X1    g11206(.A(new_n10576_), .B(new_n9962_), .Y(new_n12209_));
  AND2X1   g11207(.A(new_n12209_), .B(new_n12208_), .Y(new_n12210_));
  XOR2X1   g11208(.A(new_n10624_), .B(new_n12210_), .Y(new_n12211_));
  OAI22X1  g11209(.A0(new_n10679_), .A1(new_n12211_), .B0(new_n10572_), .B1(new_n10571_), .Y(new_n12212_));
  NAND2X1  g11210(.A(new_n10679_), .B(new_n12211_), .Y(new_n12213_));
  AND2X1   g11211(.A(new_n12213_), .B(new_n12212_), .Y(new_n12214_));
  AOI22X1  g11212(.A0(new_n10676_), .A1(new_n10668_), .B0(new_n10655_), .B1(new_n10645_), .Y(new_n12215_));
  AOI21X1  g11213(.A0(new_n10633_), .A1(new_n10629_), .B0(new_n12215_), .Y(new_n12216_));
  AOI22X1  g11214(.A0(new_n10675_), .A1(new_n10674_), .B0(new_n10672_), .B1(new_n10671_), .Y(new_n12217_));
  NAND3X1  g11215(.A(new_n10676_), .B(new_n10655_), .C(new_n10645_), .Y(new_n12218_));
  NOR2X1   g11216(.A(new_n12218_), .B(new_n12217_), .Y(new_n12219_));
  OR4X1    g11217(.A(new_n9908_), .B(new_n9902_), .C(new_n9895_), .D(new_n9890_), .Y(new_n12220_));
  AOI22X1  g11218(.A0(new_n10643_), .A1(new_n10640_), .B0(new_n12220_), .B1(new_n10648_), .Y(new_n12221_));
  NOR2X1   g11219(.A(new_n10643_), .B(new_n10640_), .Y(new_n12222_));
  NOR2X1   g11220(.A(new_n12222_), .B(new_n12221_), .Y(new_n12223_));
  AOI22X1  g11221(.A0(new_n10666_), .A1(new_n10663_), .B0(new_n10672_), .B1(new_n10671_), .Y(new_n12224_));
  NOR2X1   g11222(.A(new_n10666_), .B(new_n10663_), .Y(new_n12225_));
  OR2X1    g11223(.A(new_n12225_), .B(new_n12224_), .Y(new_n12226_));
  NOR2X1   g11224(.A(new_n12226_), .B(new_n12223_), .Y(new_n12227_));
  AND2X1   g11225(.A(new_n12226_), .B(new_n12223_), .Y(new_n12228_));
  OAI22X1  g11226(.A0(new_n12228_), .A1(new_n12227_), .B0(new_n12219_), .B1(new_n12216_), .Y(new_n12229_));
  AOI22X1  g11227(.A0(new_n10632_), .A1(new_n9876_), .B0(new_n12138_), .B1(new_n12133_), .Y(new_n12230_));
  NOR2X1   g11228(.A(new_n10632_), .B(new_n9876_), .Y(new_n12231_));
  AND2X1   g11229(.A(new_n10655_), .B(new_n10645_), .Y(new_n12232_));
  OAI22X1  g11230(.A0(new_n10677_), .A1(new_n12232_), .B0(new_n12231_), .B1(new_n12230_), .Y(new_n12233_));
  NAND4X1  g11231(.A(new_n10676_), .B(new_n10668_), .C(new_n10655_), .D(new_n10645_), .Y(new_n12234_));
  OR2X1    g11232(.A(new_n12226_), .B(new_n12223_), .Y(new_n12235_));
  NAND2X1  g11233(.A(new_n12226_), .B(new_n12223_), .Y(new_n12236_));
  NAND4X1  g11234(.A(new_n12236_), .B(new_n12235_), .C(new_n12234_), .D(new_n12233_), .Y(new_n12237_));
  NAND2X1  g11235(.A(new_n12237_), .B(new_n12229_), .Y(new_n12238_));
  AOI22X1  g11236(.A0(new_n10622_), .A1(new_n10615_), .B0(new_n10600_), .B1(new_n10590_), .Y(new_n12239_));
  AOI21X1  g11237(.A0(new_n12209_), .A1(new_n12208_), .B0(new_n12239_), .Y(new_n12240_));
  AOI22X1  g11238(.A0(new_n10621_), .A1(new_n10620_), .B0(new_n10619_), .B1(new_n10618_), .Y(new_n12241_));
  NAND3X1  g11239(.A(new_n10622_), .B(new_n10600_), .C(new_n10590_), .Y(new_n12242_));
  NOR2X1   g11240(.A(new_n12242_), .B(new_n12241_), .Y(new_n12243_));
  OR4X1    g11241(.A(new_n9994_), .B(new_n9988_), .C(new_n9981_), .D(new_n9976_), .Y(new_n12244_));
  AOI22X1  g11242(.A0(new_n10588_), .A1(new_n10585_), .B0(new_n12244_), .B1(new_n10593_), .Y(new_n12245_));
  NOR2X1   g11243(.A(new_n10588_), .B(new_n10585_), .Y(new_n12246_));
  NOR2X1   g11244(.A(new_n12246_), .B(new_n12245_), .Y(new_n12247_));
  OR2X1    g11245(.A(new_n10607_), .B(new_n9957_), .Y(new_n12248_));
  AND2X1   g11246(.A(new_n10608_), .B(new_n12248_), .Y(new_n12249_));
  AOI22X1  g11247(.A0(new_n10612_), .A1(new_n12249_), .B0(new_n10619_), .B1(new_n10618_), .Y(new_n12250_));
  AOI21X1  g11248(.A0(new_n10608_), .A1(new_n12248_), .B0(new_n10612_), .Y(new_n12251_));
  OR2X1    g11249(.A(new_n12251_), .B(new_n12250_), .Y(new_n12252_));
  NOR2X1   g11250(.A(new_n12252_), .B(new_n12247_), .Y(new_n12253_));
  AND2X1   g11251(.A(new_n12252_), .B(new_n12247_), .Y(new_n12254_));
  OAI22X1  g11252(.A0(new_n12254_), .A1(new_n12253_), .B0(new_n12243_), .B1(new_n12240_), .Y(new_n12255_));
  AND2X1   g11253(.A(new_n10600_), .B(new_n10590_), .Y(new_n12256_));
  OAI22X1  g11254(.A0(new_n10623_), .A1(new_n12256_), .B0(new_n10578_), .B1(new_n10577_), .Y(new_n12257_));
  NAND4X1  g11255(.A(new_n10622_), .B(new_n10615_), .C(new_n10600_), .D(new_n10590_), .Y(new_n12258_));
  OR2X1    g11256(.A(new_n12252_), .B(new_n12247_), .Y(new_n12259_));
  NAND2X1  g11257(.A(new_n12252_), .B(new_n12247_), .Y(new_n12260_));
  NAND4X1  g11258(.A(new_n12260_), .B(new_n12259_), .C(new_n12258_), .D(new_n12257_), .Y(new_n12261_));
  AND2X1   g11259(.A(new_n12261_), .B(new_n12255_), .Y(new_n12262_));
  XOR2X1   g11260(.A(new_n12262_), .B(new_n12238_), .Y(new_n12263_));
  XOR2X1   g11261(.A(new_n12263_), .B(new_n12214_), .Y(new_n12264_));
  XOR2X1   g11262(.A(new_n12264_), .B(new_n12205_), .Y(new_n12265_));
  XOR2X1   g11263(.A(new_n12265_), .B(new_n12147_), .Y(new_n12266_));
  XOR2X1   g11264(.A(new_n12266_), .B(new_n12132_), .Y(new_n12267_));
  XOR2X1   g11265(.A(new_n12267_), .B(new_n11993_), .Y(new_n12268_));
  XOR2X1   g11266(.A(new_n12268_), .B(new_n11982_), .Y(new_n12269_));
  OR2X1    g11267(.A(new_n12269_), .B(new_n11806_), .Y(new_n12270_));
  OR2X1    g11268(.A(new_n11337_), .B(new_n11803_), .Y(new_n12271_));
  AND2X1   g11269(.A(new_n11337_), .B(new_n11803_), .Y(new_n12272_));
  AOI21X1  g11270(.A0(new_n12271_), .A1(new_n11342_), .B0(new_n12272_), .Y(new_n12273_));
  XOR2X1   g11271(.A(new_n12269_), .B(new_n12273_), .Y(new_n12274_));
  AOI21X1  g11272(.A0(new_n10268_), .A1(new_n10145_), .B0(new_n10021_), .Y(new_n12275_));
  NOR2X1   g11273(.A(new_n10268_), .B(new_n10145_), .Y(new_n12276_));
  OR2X1    g11274(.A(new_n12276_), .B(new_n12275_), .Y(new_n12277_));
  XOR2X1   g11275(.A(new_n11779_), .B(new_n12277_), .Y(new_n12278_));
  AOI22X1  g11276(.A0(new_n12278_), .A1(new_n11559_), .B0(new_n11789_), .B1(new_n11788_), .Y(new_n12279_));
  XOR2X1   g11277(.A(new_n10401_), .B(new_n11454_), .Y(new_n12280_));
  XOR2X1   g11278(.A(new_n10534_), .B(new_n11350_), .Y(new_n12281_));
  OAI21X1  g11279(.A0(new_n12281_), .A1(new_n12280_), .B0(new_n11786_), .Y(new_n12282_));
  OR2X1    g11280(.A(new_n10535_), .B(new_n10402_), .Y(new_n12283_));
  AND2X1   g11281(.A(new_n12283_), .B(new_n12282_), .Y(new_n12284_));
  XOR2X1   g11282(.A(new_n11558_), .B(new_n12284_), .Y(new_n12285_));
  AND2X1   g11283(.A(new_n11780_), .B(new_n12285_), .Y(new_n12286_));
  OR2X1    g11284(.A(new_n12286_), .B(new_n12279_), .Y(new_n12287_));
  AOI21X1  g11285(.A0(new_n10143_), .A1(new_n10083_), .B0(new_n10022_), .Y(new_n12288_));
  NOR2X1   g11286(.A(new_n10143_), .B(new_n10083_), .Y(new_n12289_));
  OR2X1    g11287(.A(new_n12289_), .B(new_n12288_), .Y(new_n12290_));
  XOR2X1   g11288(.A(new_n11777_), .B(new_n12290_), .Y(new_n12291_));
  AOI22X1  g11289(.A0(new_n12291_), .A1(new_n11670_), .B0(new_n11567_), .B1(new_n11566_), .Y(new_n12292_));
  NAND2X1  g11290(.A(new_n11570_), .B(new_n10206_), .Y(new_n12293_));
  NOR2X1   g11291(.A(new_n11570_), .B(new_n10206_), .Y(new_n12294_));
  AOI21X1  g11292(.A0(new_n12293_), .A1(new_n10146_), .B0(new_n12294_), .Y(new_n12295_));
  XOR2X1   g11293(.A(new_n11669_), .B(new_n12295_), .Y(new_n12296_));
  AND2X1   g11294(.A(new_n11778_), .B(new_n12296_), .Y(new_n12297_));
  OR2X1    g11295(.A(new_n12297_), .B(new_n12292_), .Y(new_n12298_));
  AOI21X1  g11296(.A0(new_n11731_), .A1(new_n10053_), .B0(new_n11671_), .Y(new_n12299_));
  NOR2X1   g11297(.A(new_n11731_), .B(new_n10053_), .Y(new_n12300_));
  OR2X1    g11298(.A(new_n12300_), .B(new_n12299_), .Y(new_n12301_));
  XOR2X1   g11299(.A(new_n11775_), .B(new_n12301_), .Y(new_n12302_));
  AOI22X1  g11300(.A0(new_n12302_), .A1(new_n11725_), .B0(new_n11676_), .B1(new_n11675_), .Y(new_n12303_));
  AOI21X1  g11301(.A0(new_n11680_), .A1(new_n10084_), .B0(new_n11682_), .Y(new_n12304_));
  XOR2X1   g11302(.A(new_n11724_), .B(new_n12304_), .Y(new_n12305_));
  AND2X1   g11303(.A(new_n11776_), .B(new_n12305_), .Y(new_n12306_));
  OR2X1    g11304(.A(new_n12306_), .B(new_n12303_), .Y(new_n12307_));
  AOI22X1  g11305(.A0(new_n11773_), .A1(new_n11766_), .B0(new_n11752_), .B1(new_n11747_), .Y(new_n12308_));
  AOI21X1  g11306(.A0(new_n11732_), .A1(new_n11729_), .B0(new_n12308_), .Y(new_n12309_));
  AOI22X1  g11307(.A0(new_n11772_), .A1(new_n11771_), .B0(new_n11769_), .B1(new_n11768_), .Y(new_n12310_));
  NAND3X1  g11308(.A(new_n11773_), .B(new_n11752_), .C(new_n11747_), .Y(new_n12311_));
  NOR2X1   g11309(.A(new_n12311_), .B(new_n12310_), .Y(new_n12312_));
  AND2X1   g11310(.A(new_n11741_), .B(new_n11740_), .Y(new_n12313_));
  AOI21X1  g11311(.A0(new_n11745_), .A1(new_n12313_), .B0(new_n11738_), .Y(new_n12314_));
  NOR2X1   g11312(.A(new_n11745_), .B(new_n12313_), .Y(new_n12315_));
  OR2X1    g11313(.A(new_n12315_), .B(new_n12314_), .Y(new_n12316_));
  AOI22X1  g11314(.A0(new_n11764_), .A1(new_n11761_), .B0(new_n11769_), .B1(new_n11768_), .Y(new_n12317_));
  NOR2X1   g11315(.A(new_n11764_), .B(new_n11761_), .Y(new_n12318_));
  OR2X1    g11316(.A(new_n12318_), .B(new_n12317_), .Y(new_n12319_));
  XOR2X1   g11317(.A(new_n12319_), .B(new_n12316_), .Y(new_n12320_));
  OAI21X1  g11318(.A0(new_n12312_), .A1(new_n12309_), .B0(new_n12320_), .Y(new_n12321_));
  NOR2X1   g11319(.A(new_n12318_), .B(new_n12317_), .Y(new_n12322_));
  AND2X1   g11320(.A(new_n12322_), .B(new_n12316_), .Y(new_n12323_));
  NOR2X1   g11321(.A(new_n12322_), .B(new_n12316_), .Y(new_n12324_));
  OR4X1    g11322(.A(new_n12324_), .B(new_n12323_), .C(new_n12312_), .D(new_n12309_), .Y(new_n12325_));
  NAND2X1  g11323(.A(new_n12325_), .B(new_n12321_), .Y(new_n12326_));
  AOI22X1  g11324(.A0(new_n11722_), .A1(new_n11717_), .B0(new_n11702_), .B1(new_n11697_), .Y(new_n12327_));
  NAND4X1  g11325(.A(new_n11722_), .B(new_n11717_), .C(new_n11702_), .D(new_n11697_), .Y(new_n12328_));
  OAI21X1  g11326(.A0(new_n12327_), .A1(new_n12304_), .B0(new_n12328_), .Y(new_n12329_));
  AND2X1   g11327(.A(new_n11691_), .B(new_n11690_), .Y(new_n12330_));
  AOI21X1  g11328(.A0(new_n11695_), .A1(new_n12330_), .B0(new_n11688_), .Y(new_n12331_));
  NOR2X1   g11329(.A(new_n11695_), .B(new_n12330_), .Y(new_n12332_));
  OR2X1    g11330(.A(new_n12332_), .B(new_n12331_), .Y(new_n12333_));
  NAND2X1  g11331(.A(new_n11715_), .B(new_n11712_), .Y(new_n12334_));
  AND2X1   g11332(.A(new_n12334_), .B(new_n11708_), .Y(new_n12335_));
  NOR2X1   g11333(.A(new_n11715_), .B(new_n11712_), .Y(new_n12336_));
  OR2X1    g11334(.A(new_n12336_), .B(new_n12335_), .Y(new_n12337_));
  XOR2X1   g11335(.A(new_n12337_), .B(new_n12333_), .Y(new_n12338_));
  NAND2X1  g11336(.A(new_n12338_), .B(new_n12329_), .Y(new_n12339_));
  OR2X1    g11337(.A(new_n12327_), .B(new_n12304_), .Y(new_n12340_));
  AOI21X1  g11338(.A0(new_n12334_), .A1(new_n11708_), .B0(new_n12336_), .Y(new_n12341_));
  OAI21X1  g11339(.A0(new_n12332_), .A1(new_n12331_), .B0(new_n12341_), .Y(new_n12342_));
  OR2X1    g11340(.A(new_n12341_), .B(new_n12333_), .Y(new_n12343_));
  NAND4X1  g11341(.A(new_n12343_), .B(new_n12342_), .C(new_n12328_), .D(new_n12340_), .Y(new_n12344_));
  AND2X1   g11342(.A(new_n12344_), .B(new_n12339_), .Y(new_n12345_));
  XOR2X1   g11343(.A(new_n12345_), .B(new_n12326_), .Y(new_n12346_));
  XOR2X1   g11344(.A(new_n12346_), .B(new_n12307_), .Y(new_n12347_));
  AOI21X1  g11345(.A0(new_n11576_), .A1(new_n11569_), .B0(new_n11578_), .Y(new_n12348_));
  XOR2X1   g11346(.A(new_n11620_), .B(new_n12348_), .Y(new_n12349_));
  OAI21X1  g11347(.A0(new_n11668_), .A1(new_n12349_), .B0(new_n11573_), .Y(new_n12350_));
  NAND2X1  g11348(.A(new_n11668_), .B(new_n12349_), .Y(new_n12351_));
  AND2X1   g11349(.A(new_n12351_), .B(new_n12350_), .Y(new_n12352_));
  AOI22X1  g11350(.A0(new_n11665_), .A1(new_n11660_), .B0(new_n11645_), .B1(new_n11640_), .Y(new_n12353_));
  NAND4X1  g11351(.A(new_n11665_), .B(new_n11660_), .C(new_n11645_), .D(new_n11640_), .Y(new_n12354_));
  OAI21X1  g11352(.A0(new_n12353_), .A1(new_n11625_), .B0(new_n12354_), .Y(new_n12355_));
  AND2X1   g11353(.A(new_n11634_), .B(new_n11633_), .Y(new_n12356_));
  AOI21X1  g11354(.A0(new_n11638_), .A1(new_n12356_), .B0(new_n11631_), .Y(new_n12357_));
  NOR2X1   g11355(.A(new_n11638_), .B(new_n12356_), .Y(new_n12358_));
  OR2X1    g11356(.A(new_n12358_), .B(new_n12357_), .Y(new_n12359_));
  NAND2X1  g11357(.A(new_n11658_), .B(new_n11655_), .Y(new_n12360_));
  AND2X1   g11358(.A(new_n12360_), .B(new_n11651_), .Y(new_n12361_));
  NOR2X1   g11359(.A(new_n11658_), .B(new_n11655_), .Y(new_n12362_));
  OR2X1    g11360(.A(new_n12362_), .B(new_n12361_), .Y(new_n12363_));
  XOR2X1   g11361(.A(new_n12363_), .B(new_n12359_), .Y(new_n12364_));
  NAND2X1  g11362(.A(new_n12364_), .B(new_n12355_), .Y(new_n12365_));
  NOR2X1   g11363(.A(new_n12353_), .B(new_n11625_), .Y(new_n12366_));
  NAND3X1  g11364(.A(new_n11665_), .B(new_n11645_), .C(new_n11640_), .Y(new_n12367_));
  AOI21X1  g11365(.A0(new_n11659_), .A1(new_n11651_), .B0(new_n12367_), .Y(new_n12368_));
  AOI21X1  g11366(.A0(new_n12360_), .A1(new_n11651_), .B0(new_n12362_), .Y(new_n12369_));
  AND2X1   g11367(.A(new_n12369_), .B(new_n12359_), .Y(new_n12370_));
  NOR3X1   g11368(.A(new_n12369_), .B(new_n12358_), .C(new_n12357_), .Y(new_n12371_));
  OR4X1    g11369(.A(new_n12371_), .B(new_n12370_), .C(new_n12368_), .D(new_n12366_), .Y(new_n12372_));
  NAND2X1  g11370(.A(new_n12372_), .B(new_n12365_), .Y(new_n12373_));
  AOI22X1  g11371(.A0(new_n11618_), .A1(new_n11613_), .B0(new_n11598_), .B1(new_n11593_), .Y(new_n12374_));
  NAND4X1  g11372(.A(new_n11618_), .B(new_n11613_), .C(new_n11598_), .D(new_n11593_), .Y(new_n12375_));
  OAI21X1  g11373(.A0(new_n12374_), .A1(new_n12348_), .B0(new_n12375_), .Y(new_n12376_));
  AND2X1   g11374(.A(new_n11587_), .B(new_n11586_), .Y(new_n12377_));
  AOI21X1  g11375(.A0(new_n11591_), .A1(new_n12377_), .B0(new_n11584_), .Y(new_n12378_));
  NOR2X1   g11376(.A(new_n11591_), .B(new_n12377_), .Y(new_n12379_));
  OR2X1    g11377(.A(new_n12379_), .B(new_n12378_), .Y(new_n12380_));
  NAND2X1  g11378(.A(new_n11611_), .B(new_n11608_), .Y(new_n12381_));
  AND2X1   g11379(.A(new_n12381_), .B(new_n11604_), .Y(new_n12382_));
  NOR2X1   g11380(.A(new_n11611_), .B(new_n11608_), .Y(new_n12383_));
  OR2X1    g11381(.A(new_n12383_), .B(new_n12382_), .Y(new_n12384_));
  XOR2X1   g11382(.A(new_n12384_), .B(new_n12380_), .Y(new_n12385_));
  NAND2X1  g11383(.A(new_n12385_), .B(new_n12376_), .Y(new_n12386_));
  NOR2X1   g11384(.A(new_n12374_), .B(new_n12348_), .Y(new_n12387_));
  NAND3X1  g11385(.A(new_n11618_), .B(new_n11598_), .C(new_n11593_), .Y(new_n12388_));
  AOI21X1  g11386(.A0(new_n11612_), .A1(new_n11604_), .B0(new_n12388_), .Y(new_n12389_));
  AOI21X1  g11387(.A0(new_n12381_), .A1(new_n11604_), .B0(new_n12383_), .Y(new_n12390_));
  AND2X1   g11388(.A(new_n12390_), .B(new_n12380_), .Y(new_n12391_));
  NOR3X1   g11389(.A(new_n12390_), .B(new_n12379_), .C(new_n12378_), .Y(new_n12392_));
  OR4X1    g11390(.A(new_n12392_), .B(new_n12391_), .C(new_n12389_), .D(new_n12387_), .Y(new_n12393_));
  AND2X1   g11391(.A(new_n12393_), .B(new_n12386_), .Y(new_n12394_));
  XOR2X1   g11392(.A(new_n12394_), .B(new_n12373_), .Y(new_n12395_));
  XOR2X1   g11393(.A(new_n12395_), .B(new_n12352_), .Y(new_n12396_));
  XOR2X1   g11394(.A(new_n12396_), .B(new_n12347_), .Y(new_n12397_));
  XOR2X1   g11395(.A(new_n12397_), .B(new_n12298_), .Y(new_n12398_));
  AOI21X1  g11396(.A0(new_n2035_), .A1(new_n2389_), .B0(new_n2391_), .Y(new_n12399_));
  XOR2X1   g11397(.A(new_n10465_), .B(new_n12399_), .Y(new_n12400_));
  OAI21X1  g11398(.A0(new_n10533_), .A1(new_n12400_), .B0(new_n10403_), .Y(new_n12401_));
  OR2X1    g11399(.A(new_n11352_), .B(new_n10466_), .Y(new_n12402_));
  AND2X1   g11400(.A(new_n12402_), .B(new_n12401_), .Y(new_n12403_));
  XOR2X1   g11401(.A(new_n11452_), .B(new_n12403_), .Y(new_n12404_));
  OAI22X1  g11402(.A0(new_n11557_), .A1(new_n12404_), .B0(new_n11348_), .B1(new_n11347_), .Y(new_n12405_));
  NAND2X1  g11403(.A(new_n11557_), .B(new_n12404_), .Y(new_n12406_));
  AND2X1   g11404(.A(new_n12406_), .B(new_n12405_), .Y(new_n12407_));
  AND2X1   g11405(.A(new_n11511_), .B(new_n10274_), .Y(new_n12408_));
  OR2X1    g11406(.A(new_n11512_), .B(new_n12408_), .Y(new_n12409_));
  XOR2X1   g11407(.A(new_n11554_), .B(new_n12409_), .Y(new_n12410_));
  AOI22X1  g11408(.A0(new_n12410_), .A1(new_n11508_), .B0(new_n11460_), .B1(new_n11459_), .Y(new_n12411_));
  XOR2X1   g11409(.A(new_n10365_), .B(new_n11486_), .Y(new_n12412_));
  XOR2X1   g11410(.A(new_n12412_), .B(new_n10337_), .Y(new_n12413_));
  OAI21X1  g11411(.A0(new_n10398_), .A1(new_n12413_), .B0(new_n10334_), .Y(new_n12414_));
  OR2X1    g11412(.A(new_n11463_), .B(new_n10367_), .Y(new_n12415_));
  AND2X1   g11413(.A(new_n12415_), .B(new_n12414_), .Y(new_n12416_));
  XOR2X1   g11414(.A(new_n11507_), .B(new_n12416_), .Y(new_n12417_));
  AND2X1   g11415(.A(new_n11555_), .B(new_n12417_), .Y(new_n12418_));
  OR2X1    g11416(.A(new_n12418_), .B(new_n12411_), .Y(new_n12419_));
  AOI22X1  g11417(.A0(new_n11552_), .A1(new_n11547_), .B0(new_n11532_), .B1(new_n11527_), .Y(new_n12420_));
  NAND4X1  g11418(.A(new_n11552_), .B(new_n11547_), .C(new_n11532_), .D(new_n11527_), .Y(new_n12421_));
  OAI21X1  g11419(.A0(new_n12420_), .A1(new_n11513_), .B0(new_n12421_), .Y(new_n12422_));
  AND2X1   g11420(.A(new_n11521_), .B(new_n11520_), .Y(new_n12423_));
  AOI21X1  g11421(.A0(new_n11525_), .A1(new_n12423_), .B0(new_n11518_), .Y(new_n12424_));
  NOR2X1   g11422(.A(new_n11525_), .B(new_n12423_), .Y(new_n12425_));
  OR2X1    g11423(.A(new_n12425_), .B(new_n12424_), .Y(new_n12426_));
  NAND2X1  g11424(.A(new_n11545_), .B(new_n11542_), .Y(new_n12427_));
  AND2X1   g11425(.A(new_n12427_), .B(new_n11538_), .Y(new_n12428_));
  NOR2X1   g11426(.A(new_n11545_), .B(new_n11542_), .Y(new_n12429_));
  OR2X1    g11427(.A(new_n12429_), .B(new_n12428_), .Y(new_n12430_));
  XOR2X1   g11428(.A(new_n12430_), .B(new_n12426_), .Y(new_n12431_));
  NAND2X1  g11429(.A(new_n12431_), .B(new_n12422_), .Y(new_n12432_));
  NOR2X1   g11430(.A(new_n12420_), .B(new_n11513_), .Y(new_n12433_));
  NAND3X1  g11431(.A(new_n11552_), .B(new_n11532_), .C(new_n11527_), .Y(new_n12434_));
  AOI21X1  g11432(.A0(new_n11546_), .A1(new_n11538_), .B0(new_n12434_), .Y(new_n12435_));
  AOI21X1  g11433(.A0(new_n12427_), .A1(new_n11538_), .B0(new_n12429_), .Y(new_n12436_));
  AND2X1   g11434(.A(new_n12436_), .B(new_n12426_), .Y(new_n12437_));
  NOR3X1   g11435(.A(new_n12436_), .B(new_n12425_), .C(new_n12424_), .Y(new_n12438_));
  OR4X1    g11436(.A(new_n12438_), .B(new_n12437_), .C(new_n12435_), .D(new_n12433_), .Y(new_n12439_));
  NAND2X1  g11437(.A(new_n12439_), .B(new_n12432_), .Y(new_n12440_));
  AOI22X1  g11438(.A0(new_n11505_), .A1(new_n11499_), .B0(new_n11483_), .B1(new_n11479_), .Y(new_n12441_));
  AOI21X1  g11439(.A0(new_n12415_), .A1(new_n12414_), .B0(new_n12441_), .Y(new_n12442_));
  AOI22X1  g11440(.A0(new_n11504_), .A1(new_n11503_), .B0(new_n11502_), .B1(new_n11501_), .Y(new_n12443_));
  NAND3X1  g11441(.A(new_n11505_), .B(new_n11483_), .C(new_n11479_), .Y(new_n12444_));
  NOR2X1   g11442(.A(new_n12444_), .B(new_n12443_), .Y(new_n12445_));
  AOI22X1  g11443(.A0(new_n11471_), .A1(new_n10388_), .B0(new_n10386_), .B1(new_n10385_), .Y(new_n12446_));
  AOI21X1  g11444(.A0(new_n11477_), .A1(new_n12446_), .B0(new_n11469_), .Y(new_n12447_));
  NOR2X1   g11445(.A(new_n11477_), .B(new_n12446_), .Y(new_n12448_));
  NOR2X1   g11446(.A(new_n12448_), .B(new_n12447_), .Y(new_n12449_));
  AOI22X1  g11447(.A0(new_n11497_), .A1(new_n11492_), .B0(new_n11502_), .B1(new_n11501_), .Y(new_n12450_));
  AOI21X1  g11448(.A0(new_n11495_), .A1(new_n11494_), .B0(new_n11492_), .Y(new_n12451_));
  OR2X1    g11449(.A(new_n12451_), .B(new_n12450_), .Y(new_n12452_));
  NOR2X1   g11450(.A(new_n12452_), .B(new_n12449_), .Y(new_n12453_));
  AND2X1   g11451(.A(new_n12452_), .B(new_n12449_), .Y(new_n12454_));
  OAI22X1  g11452(.A0(new_n12454_), .A1(new_n12453_), .B0(new_n12445_), .B1(new_n12442_), .Y(new_n12455_));
  AND2X1   g11453(.A(new_n11483_), .B(new_n11479_), .Y(new_n12456_));
  OAI22X1  g11454(.A0(new_n11506_), .A1(new_n12456_), .B0(new_n11465_), .B1(new_n11464_), .Y(new_n12457_));
  NAND4X1  g11455(.A(new_n11505_), .B(new_n11499_), .C(new_n11483_), .D(new_n11479_), .Y(new_n12458_));
  OR2X1    g11456(.A(new_n12452_), .B(new_n12449_), .Y(new_n12459_));
  NAND2X1  g11457(.A(new_n12452_), .B(new_n12449_), .Y(new_n12460_));
  NAND4X1  g11458(.A(new_n12460_), .B(new_n12459_), .C(new_n12458_), .D(new_n12457_), .Y(new_n12461_));
  AND2X1   g11459(.A(new_n12461_), .B(new_n12455_), .Y(new_n12462_));
  XOR2X1   g11460(.A(new_n12462_), .B(new_n12440_), .Y(new_n12463_));
  XOR2X1   g11461(.A(new_n12463_), .B(new_n12419_), .Y(new_n12464_));
  XOR2X1   g11462(.A(new_n10498_), .B(new_n11380_), .Y(new_n12465_));
  XOR2X1   g11463(.A(new_n12465_), .B(new_n10470_), .Y(new_n12466_));
  OAI21X1  g11464(.A0(new_n10531_), .A1(new_n12466_), .B0(new_n11351_), .Y(new_n12467_));
  OR2X1    g11465(.A(new_n11357_), .B(new_n10500_), .Y(new_n12468_));
  AND2X1   g11466(.A(new_n12468_), .B(new_n12467_), .Y(new_n12469_));
  XOR2X1   g11467(.A(new_n11401_), .B(new_n12469_), .Y(new_n12470_));
  OAI22X1  g11468(.A0(new_n11451_), .A1(new_n12470_), .B0(new_n11354_), .B1(new_n11353_), .Y(new_n12471_));
  NAND2X1  g11469(.A(new_n11451_), .B(new_n12470_), .Y(new_n12472_));
  AND2X1   g11470(.A(new_n12472_), .B(new_n12471_), .Y(new_n12473_));
  AOI22X1  g11471(.A0(new_n11448_), .A1(new_n11445_), .B0(new_n11427_), .B1(new_n11423_), .Y(new_n12474_));
  AOI21X1  g11472(.A0(new_n11409_), .A1(new_n11406_), .B0(new_n12474_), .Y(new_n12475_));
  NAND3X1  g11473(.A(new_n11448_), .B(new_n11427_), .C(new_n11423_), .Y(new_n12476_));
  AOI21X1  g11474(.A0(new_n11444_), .A1(new_n11433_), .B0(new_n12476_), .Y(new_n12477_));
  AOI22X1  g11475(.A0(new_n11415_), .A1(new_n10454_), .B0(new_n10452_), .B1(new_n10451_), .Y(new_n12478_));
  AOI21X1  g11476(.A0(new_n11421_), .A1(new_n12478_), .B0(new_n11413_), .Y(new_n12479_));
  NOR2X1   g11477(.A(new_n11421_), .B(new_n12478_), .Y(new_n12480_));
  NOR2X1   g11478(.A(new_n12480_), .B(new_n12479_), .Y(new_n12481_));
  NAND4X1  g11479(.A(new_n11440_), .B(new_n11439_), .C(new_n11436_), .D(new_n11435_), .Y(new_n12482_));
  AND2X1   g11480(.A(new_n12482_), .B(new_n11433_), .Y(new_n12483_));
  AOI22X1  g11481(.A0(new_n11440_), .A1(new_n11439_), .B0(new_n11436_), .B1(new_n11435_), .Y(new_n12484_));
  OR2X1    g11482(.A(new_n12484_), .B(new_n12483_), .Y(new_n12485_));
  NOR2X1   g11483(.A(new_n12485_), .B(new_n12481_), .Y(new_n12486_));
  AOI21X1  g11484(.A0(new_n12482_), .A1(new_n11433_), .B0(new_n12484_), .Y(new_n12487_));
  NOR3X1   g11485(.A(new_n12487_), .B(new_n12480_), .C(new_n12479_), .Y(new_n12488_));
  OAI22X1  g11486(.A0(new_n12488_), .A1(new_n12486_), .B0(new_n12477_), .B1(new_n12475_), .Y(new_n12489_));
  AOI21X1  g11487(.A0(new_n11408_), .A1(new_n10433_), .B0(new_n12399_), .Y(new_n12490_));
  NOR2X1   g11488(.A(new_n11408_), .B(new_n10433_), .Y(new_n12491_));
  AND2X1   g11489(.A(new_n11427_), .B(new_n11423_), .Y(new_n12492_));
  OAI22X1  g11490(.A0(new_n11449_), .A1(new_n12492_), .B0(new_n12491_), .B1(new_n12490_), .Y(new_n12493_));
  NAND4X1  g11491(.A(new_n11448_), .B(new_n11445_), .C(new_n11427_), .D(new_n11423_), .Y(new_n12494_));
  OAI21X1  g11492(.A0(new_n12480_), .A1(new_n12479_), .B0(new_n12487_), .Y(new_n12495_));
  NAND2X1  g11493(.A(new_n12485_), .B(new_n12481_), .Y(new_n12496_));
  NAND4X1  g11494(.A(new_n12496_), .B(new_n12495_), .C(new_n12494_), .D(new_n12493_), .Y(new_n12497_));
  NAND2X1  g11495(.A(new_n12497_), .B(new_n12489_), .Y(new_n12498_));
  AOI22X1  g11496(.A0(new_n11399_), .A1(new_n11393_), .B0(new_n11377_), .B1(new_n11373_), .Y(new_n12499_));
  AOI21X1  g11497(.A0(new_n12468_), .A1(new_n12467_), .B0(new_n12499_), .Y(new_n12500_));
  AOI22X1  g11498(.A0(new_n11398_), .A1(new_n11397_), .B0(new_n11396_), .B1(new_n11395_), .Y(new_n12501_));
  NAND3X1  g11499(.A(new_n11399_), .B(new_n11377_), .C(new_n11373_), .Y(new_n12502_));
  NOR2X1   g11500(.A(new_n12502_), .B(new_n12501_), .Y(new_n12503_));
  AOI22X1  g11501(.A0(new_n11365_), .A1(new_n10521_), .B0(new_n10519_), .B1(new_n10518_), .Y(new_n12504_));
  AOI21X1  g11502(.A0(new_n11371_), .A1(new_n12504_), .B0(new_n11363_), .Y(new_n12505_));
  NOR2X1   g11503(.A(new_n11371_), .B(new_n12504_), .Y(new_n12506_));
  NOR2X1   g11504(.A(new_n12506_), .B(new_n12505_), .Y(new_n12507_));
  AOI22X1  g11505(.A0(new_n11391_), .A1(new_n11386_), .B0(new_n11396_), .B1(new_n11395_), .Y(new_n12508_));
  AOI21X1  g11506(.A0(new_n11389_), .A1(new_n11388_), .B0(new_n11386_), .Y(new_n12509_));
  OR2X1    g11507(.A(new_n12509_), .B(new_n12508_), .Y(new_n12510_));
  NOR2X1   g11508(.A(new_n12510_), .B(new_n12507_), .Y(new_n12511_));
  AND2X1   g11509(.A(new_n12510_), .B(new_n12507_), .Y(new_n12512_));
  OAI22X1  g11510(.A0(new_n12512_), .A1(new_n12511_), .B0(new_n12503_), .B1(new_n12500_), .Y(new_n12513_));
  AND2X1   g11511(.A(new_n11377_), .B(new_n11373_), .Y(new_n12514_));
  OAI22X1  g11512(.A0(new_n11400_), .A1(new_n12514_), .B0(new_n11359_), .B1(new_n11358_), .Y(new_n12515_));
  NAND4X1  g11513(.A(new_n11399_), .B(new_n11393_), .C(new_n11377_), .D(new_n11373_), .Y(new_n12516_));
  OR2X1    g11514(.A(new_n12510_), .B(new_n12507_), .Y(new_n12517_));
  NAND2X1  g11515(.A(new_n12510_), .B(new_n12507_), .Y(new_n12518_));
  NAND4X1  g11516(.A(new_n12518_), .B(new_n12517_), .C(new_n12516_), .D(new_n12515_), .Y(new_n12519_));
  AND2X1   g11517(.A(new_n12519_), .B(new_n12513_), .Y(new_n12520_));
  XOR2X1   g11518(.A(new_n12520_), .B(new_n12498_), .Y(new_n12521_));
  XOR2X1   g11519(.A(new_n12521_), .B(new_n12473_), .Y(new_n12522_));
  XOR2X1   g11520(.A(new_n12522_), .B(new_n12464_), .Y(new_n12523_));
  XOR2X1   g11521(.A(new_n12523_), .B(new_n12407_), .Y(new_n12524_));
  XOR2X1   g11522(.A(new_n12524_), .B(new_n12398_), .Y(new_n12525_));
  XOR2X1   g11523(.A(new_n12525_), .B(new_n12287_), .Y(new_n12526_));
  NAND2X1  g11524(.A(new_n12526_), .B(new_n12274_), .Y(new_n12527_));
  AOI21X1  g11525(.A0(new_n12269_), .A1(new_n11806_), .B0(new_n12526_), .Y(new_n12528_));
  AOI22X1  g11526(.A0(new_n12528_), .A1(new_n12270_), .B0(new_n12527_), .B1(new_n11793_), .Y(new_n12529_));
  OR2X1    g11527(.A(new_n12268_), .B(new_n11982_), .Y(new_n12530_));
  AND2X1   g11528(.A(new_n12268_), .B(new_n11982_), .Y(new_n12531_));
  AOI21X1  g11529(.A0(new_n12530_), .A1(new_n11806_), .B0(new_n12531_), .Y(new_n12532_));
  AOI22X1  g11530(.A0(new_n9816_), .A1(new_n9730_), .B0(new_n9637_), .B1(new_n9627_), .Y(new_n12533_));
  NOR2X1   g11531(.A(new_n9816_), .B(new_n9730_), .Y(new_n12534_));
  OR2X1    g11532(.A(new_n12534_), .B(new_n12533_), .Y(new_n12535_));
  XOR2X1   g11533(.A(new_n10803_), .B(new_n12535_), .Y(new_n12536_));
  AOI22X1  g11534(.A0(new_n12536_), .A1(new_n10681_), .B0(new_n11988_), .B1(new_n11987_), .Y(new_n12537_));
  AND2X1   g11535(.A(new_n10804_), .B(new_n12144_), .Y(new_n12538_));
  OR2X1    g11536(.A(new_n12538_), .B(new_n12537_), .Y(new_n12539_));
  XOR2X1   g11537(.A(new_n12265_), .B(new_n12539_), .Y(new_n12540_));
  AOI22X1  g11538(.A0(new_n12540_), .A1(new_n12132_), .B0(new_n11992_), .B1(new_n11991_), .Y(new_n12541_));
  NOR2X1   g11539(.A(new_n12540_), .B(new_n12132_), .Y(new_n12542_));
  OR2X1    g11540(.A(new_n12542_), .B(new_n12541_), .Y(new_n12543_));
  OR2X1    g11541(.A(new_n12231_), .B(new_n12230_), .Y(new_n12544_));
  XOR2X1   g11542(.A(new_n10678_), .B(new_n12544_), .Y(new_n12545_));
  AOI22X1  g11543(.A0(new_n12545_), .A1(new_n10625_), .B0(new_n12142_), .B1(new_n12141_), .Y(new_n12546_));
  AND2X1   g11544(.A(new_n10679_), .B(new_n12211_), .Y(new_n12547_));
  OR2X1    g11545(.A(new_n12547_), .B(new_n12546_), .Y(new_n12548_));
  XOR2X1   g11546(.A(new_n12263_), .B(new_n12548_), .Y(new_n12549_));
  AOI22X1  g11547(.A0(new_n12549_), .A1(new_n12205_), .B0(new_n12146_), .B1(new_n12145_), .Y(new_n12550_));
  NOR2X1   g11548(.A(new_n12549_), .B(new_n12205_), .Y(new_n12551_));
  OR2X1    g11549(.A(new_n12551_), .B(new_n12550_), .Y(new_n12552_));
  AOI22X1  g11550(.A0(new_n12261_), .A1(new_n12255_), .B0(new_n12237_), .B1(new_n12229_), .Y(new_n12553_));
  AOI21X1  g11551(.A0(new_n12213_), .A1(new_n12212_), .B0(new_n12553_), .Y(new_n12554_));
  AOI22X1  g11552(.A0(new_n12236_), .A1(new_n12235_), .B0(new_n12234_), .B1(new_n12233_), .Y(new_n12555_));
  NOR4X1   g11553(.A(new_n12228_), .B(new_n12227_), .C(new_n12219_), .D(new_n12216_), .Y(new_n12556_));
  AOI22X1  g11554(.A0(new_n12260_), .A1(new_n12259_), .B0(new_n12258_), .B1(new_n12257_), .Y(new_n12557_));
  NOR4X1   g11555(.A(new_n12254_), .B(new_n12253_), .C(new_n12243_), .D(new_n12240_), .Y(new_n12558_));
  NOR4X1   g11556(.A(new_n12558_), .B(new_n12557_), .C(new_n12556_), .D(new_n12555_), .Y(new_n12559_));
  OR4X1    g11557(.A(new_n12251_), .B(new_n12250_), .C(new_n12246_), .D(new_n12245_), .Y(new_n12560_));
  OAI21X1  g11558(.A0(new_n12243_), .A1(new_n12240_), .B0(new_n12560_), .Y(new_n12561_));
  OAI22X1  g11559(.A0(new_n12251_), .A1(new_n12250_), .B0(new_n12246_), .B1(new_n12245_), .Y(new_n12562_));
  AND2X1   g11560(.A(new_n12562_), .B(new_n12561_), .Y(new_n12563_));
  OR4X1    g11561(.A(new_n12225_), .B(new_n12224_), .C(new_n12222_), .D(new_n12221_), .Y(new_n12564_));
  OAI21X1  g11562(.A0(new_n12219_), .A1(new_n12216_), .B0(new_n12564_), .Y(new_n12565_));
  OAI22X1  g11563(.A0(new_n12225_), .A1(new_n12224_), .B0(new_n12222_), .B1(new_n12221_), .Y(new_n12566_));
  AND2X1   g11564(.A(new_n12566_), .B(new_n12565_), .Y(new_n12567_));
  XOR2X1   g11565(.A(new_n12567_), .B(new_n12563_), .Y(new_n12568_));
  OAI21X1  g11566(.A0(new_n12559_), .A1(new_n12554_), .B0(new_n12568_), .Y(new_n12569_));
  OAI22X1  g11567(.A0(new_n12558_), .A1(new_n12557_), .B0(new_n12556_), .B1(new_n12555_), .Y(new_n12570_));
  OAI21X1  g11568(.A0(new_n12547_), .A1(new_n12546_), .B0(new_n12570_), .Y(new_n12571_));
  NAND2X1  g11569(.A(new_n12562_), .B(new_n12561_), .Y(new_n12572_));
  OR2X1    g11570(.A(new_n12567_), .B(new_n12572_), .Y(new_n12573_));
  AOI21X1  g11571(.A0(new_n12567_), .A1(new_n12572_), .B0(new_n12559_), .Y(new_n12574_));
  NAND3X1  g11572(.A(new_n12574_), .B(new_n12573_), .C(new_n12571_), .Y(new_n12575_));
  NAND2X1  g11573(.A(new_n12575_), .B(new_n12569_), .Y(new_n12576_));
  OAI22X1  g11574(.A0(new_n10802_), .A1(new_n12158_), .B0(new_n12534_), .B1(new_n12533_), .Y(new_n12577_));
  NAND2X1  g11575(.A(new_n10802_), .B(new_n12158_), .Y(new_n12578_));
  AOI22X1  g11576(.A0(new_n12202_), .A1(new_n12196_), .B0(new_n12178_), .B1(new_n12174_), .Y(new_n12579_));
  AOI21X1  g11577(.A0(new_n12578_), .A1(new_n12577_), .B0(new_n12579_), .Y(new_n12580_));
  AOI22X1  g11578(.A0(new_n12201_), .A1(new_n12200_), .B0(new_n12199_), .B1(new_n12198_), .Y(new_n12581_));
  NAND3X1  g11579(.A(new_n12202_), .B(new_n12178_), .C(new_n12174_), .Y(new_n12582_));
  NOR2X1   g11580(.A(new_n12582_), .B(new_n12581_), .Y(new_n12583_));
  OR4X1    g11581(.A(new_n12192_), .B(new_n12191_), .C(new_n12187_), .D(new_n12186_), .Y(new_n12584_));
  OAI21X1  g11582(.A0(new_n12184_), .A1(new_n12181_), .B0(new_n12584_), .Y(new_n12585_));
  OAI22X1  g11583(.A0(new_n12192_), .A1(new_n12191_), .B0(new_n12187_), .B1(new_n12186_), .Y(new_n12586_));
  AND2X1   g11584(.A(new_n12586_), .B(new_n12585_), .Y(new_n12587_));
  OR4X1    g11585(.A(new_n12171_), .B(new_n12170_), .C(new_n12168_), .D(new_n12167_), .Y(new_n12588_));
  OAI21X1  g11586(.A0(new_n12165_), .A1(new_n12162_), .B0(new_n12588_), .Y(new_n12589_));
  OAI22X1  g11587(.A0(new_n12171_), .A1(new_n12170_), .B0(new_n12168_), .B1(new_n12167_), .Y(new_n12590_));
  AND2X1   g11588(.A(new_n12590_), .B(new_n12589_), .Y(new_n12591_));
  XOR2X1   g11589(.A(new_n12591_), .B(new_n12587_), .Y(new_n12592_));
  OAI21X1  g11590(.A0(new_n12583_), .A1(new_n12580_), .B0(new_n12592_), .Y(new_n12593_));
  AND2X1   g11591(.A(new_n12178_), .B(new_n12174_), .Y(new_n12594_));
  OAI22X1  g11592(.A0(new_n12203_), .A1(new_n12594_), .B0(new_n12159_), .B1(new_n12152_), .Y(new_n12595_));
  NAND4X1  g11593(.A(new_n12202_), .B(new_n12196_), .C(new_n12178_), .D(new_n12174_), .Y(new_n12596_));
  NAND2X1  g11594(.A(new_n12586_), .B(new_n12585_), .Y(new_n12597_));
  NAND2X1  g11595(.A(new_n12591_), .B(new_n12597_), .Y(new_n12598_));
  OR2X1    g11596(.A(new_n12591_), .B(new_n12597_), .Y(new_n12599_));
  NAND4X1  g11597(.A(new_n12599_), .B(new_n12598_), .C(new_n12596_), .D(new_n12595_), .Y(new_n12600_));
  AND2X1   g11598(.A(new_n12600_), .B(new_n12593_), .Y(new_n12601_));
  XOR2X1   g11599(.A(new_n12601_), .B(new_n12576_), .Y(new_n12602_));
  XOR2X1   g11600(.A(new_n12602_), .B(new_n12552_), .Y(new_n12603_));
  OAI22X1  g11601(.A0(new_n11051_), .A1(new_n12023_), .B0(new_n11995_), .B1(new_n11994_), .Y(new_n12604_));
  NAND2X1  g11602(.A(new_n11051_), .B(new_n12023_), .Y(new_n12605_));
  AND2X1   g11603(.A(new_n12605_), .B(new_n12604_), .Y(new_n12606_));
  XOR2X1   g11604(.A(new_n12070_), .B(new_n12606_), .Y(new_n12607_));
  OAI22X1  g11605(.A0(new_n12130_), .A1(new_n12607_), .B0(new_n12011_), .B1(new_n11998_), .Y(new_n12608_));
  OR2X1    g11606(.A(new_n12097_), .B(new_n12096_), .Y(new_n12609_));
  XOR2X1   g11607(.A(new_n10931_), .B(new_n12609_), .Y(new_n12610_));
  AOI22X1  g11608(.A0(new_n12610_), .A1(new_n10878_), .B0(new_n12008_), .B1(new_n12007_), .Y(new_n12611_));
  AND2X1   g11609(.A(new_n10932_), .B(new_n12077_), .Y(new_n12612_));
  OR2X1    g11610(.A(new_n12612_), .B(new_n12611_), .Y(new_n12613_));
  XOR2X1   g11611(.A(new_n12129_), .B(new_n12613_), .Y(new_n12614_));
  OR2X1    g11612(.A(new_n12614_), .B(new_n12071_), .Y(new_n12615_));
  AND2X1   g11613(.A(new_n12615_), .B(new_n12608_), .Y(new_n12616_));
  AOI22X1  g11614(.A0(new_n12127_), .A1(new_n12121_), .B0(new_n12103_), .B1(new_n12095_), .Y(new_n12617_));
  AOI21X1  g11615(.A0(new_n12079_), .A1(new_n12078_), .B0(new_n12617_), .Y(new_n12618_));
  AOI22X1  g11616(.A0(new_n12102_), .A1(new_n12101_), .B0(new_n12100_), .B1(new_n12099_), .Y(new_n12619_));
  NOR4X1   g11617(.A(new_n12094_), .B(new_n12093_), .C(new_n12085_), .D(new_n12082_), .Y(new_n12620_));
  AOI22X1  g11618(.A0(new_n12126_), .A1(new_n12125_), .B0(new_n12124_), .B1(new_n12123_), .Y(new_n12621_));
  NOR4X1   g11619(.A(new_n12120_), .B(new_n12119_), .C(new_n12109_), .D(new_n12106_), .Y(new_n12622_));
  NOR4X1   g11620(.A(new_n12622_), .B(new_n12621_), .C(new_n12620_), .D(new_n12619_), .Y(new_n12623_));
  OR4X1    g11621(.A(new_n12117_), .B(new_n12116_), .C(new_n12112_), .D(new_n12111_), .Y(new_n12624_));
  OAI21X1  g11622(.A0(new_n12109_), .A1(new_n12106_), .B0(new_n12624_), .Y(new_n12625_));
  OAI22X1  g11623(.A0(new_n12117_), .A1(new_n12116_), .B0(new_n12112_), .B1(new_n12111_), .Y(new_n12626_));
  AND2X1   g11624(.A(new_n12626_), .B(new_n12625_), .Y(new_n12627_));
  OR4X1    g11625(.A(new_n12091_), .B(new_n12090_), .C(new_n12088_), .D(new_n12087_), .Y(new_n12628_));
  OAI21X1  g11626(.A0(new_n12085_), .A1(new_n12082_), .B0(new_n12628_), .Y(new_n12629_));
  OAI22X1  g11627(.A0(new_n12091_), .A1(new_n12090_), .B0(new_n12088_), .B1(new_n12087_), .Y(new_n12630_));
  AND2X1   g11628(.A(new_n12630_), .B(new_n12629_), .Y(new_n12631_));
  XOR2X1   g11629(.A(new_n12631_), .B(new_n12627_), .Y(new_n12632_));
  OAI21X1  g11630(.A0(new_n12623_), .A1(new_n12618_), .B0(new_n12632_), .Y(new_n12633_));
  OAI22X1  g11631(.A0(new_n12622_), .A1(new_n12621_), .B0(new_n12620_), .B1(new_n12619_), .Y(new_n12634_));
  OAI21X1  g11632(.A0(new_n12612_), .A1(new_n12611_), .B0(new_n12634_), .Y(new_n12635_));
  NAND2X1  g11633(.A(new_n12626_), .B(new_n12625_), .Y(new_n12636_));
  OR2X1    g11634(.A(new_n12631_), .B(new_n12636_), .Y(new_n12637_));
  AOI21X1  g11635(.A0(new_n12631_), .A1(new_n12636_), .B0(new_n12623_), .Y(new_n12638_));
  NAND3X1  g11636(.A(new_n12638_), .B(new_n12637_), .C(new_n12635_), .Y(new_n12639_));
  NAND2X1  g11637(.A(new_n12639_), .B(new_n12633_), .Y(new_n12640_));
  AOI22X1  g11638(.A0(new_n12068_), .A1(new_n12061_), .B0(new_n12046_), .B1(new_n12039_), .Y(new_n12641_));
  AOI21X1  g11639(.A0(new_n12605_), .A1(new_n12604_), .B0(new_n12641_), .Y(new_n12642_));
  AOI22X1  g11640(.A0(new_n12067_), .A1(new_n12066_), .B0(new_n12064_), .B1(new_n12063_), .Y(new_n12643_));
  NAND3X1  g11641(.A(new_n12068_), .B(new_n12046_), .C(new_n12039_), .Y(new_n12644_));
  NOR2X1   g11642(.A(new_n12644_), .B(new_n12643_), .Y(new_n12645_));
  OR4X1    g11643(.A(new_n12058_), .B(new_n12057_), .C(new_n12055_), .D(new_n12054_), .Y(new_n12646_));
  OAI21X1  g11644(.A0(new_n12052_), .A1(new_n12049_), .B0(new_n12646_), .Y(new_n12647_));
  OAI22X1  g11645(.A0(new_n12058_), .A1(new_n12057_), .B0(new_n12055_), .B1(new_n12054_), .Y(new_n12648_));
  AND2X1   g11646(.A(new_n12648_), .B(new_n12647_), .Y(new_n12649_));
  NOR4X1   g11647(.A(new_n12036_), .B(new_n12035_), .C(new_n12033_), .D(new_n12032_), .Y(new_n12650_));
  AOI21X1  g11648(.A0(new_n12042_), .A1(new_n12041_), .B0(new_n12650_), .Y(new_n12651_));
  AOI21X1  g11649(.A0(new_n12037_), .A1(new_n12034_), .B0(new_n12651_), .Y(new_n12652_));
  XOR2X1   g11650(.A(new_n12652_), .B(new_n12649_), .Y(new_n12653_));
  OAI21X1  g11651(.A0(new_n12645_), .A1(new_n12642_), .B0(new_n12653_), .Y(new_n12654_));
  AND2X1   g11652(.A(new_n12046_), .B(new_n12039_), .Y(new_n12655_));
  OAI22X1  g11653(.A0(new_n12069_), .A1(new_n12655_), .B0(new_n12024_), .B1(new_n12017_), .Y(new_n12656_));
  NAND4X1  g11654(.A(new_n12068_), .B(new_n12061_), .C(new_n12046_), .D(new_n12039_), .Y(new_n12657_));
  NAND2X1  g11655(.A(new_n12648_), .B(new_n12647_), .Y(new_n12658_));
  NAND2X1  g11656(.A(new_n12652_), .B(new_n12658_), .Y(new_n12659_));
  OR2X1    g11657(.A(new_n12652_), .B(new_n12658_), .Y(new_n12660_));
  NAND4X1  g11658(.A(new_n12660_), .B(new_n12659_), .C(new_n12657_), .D(new_n12656_), .Y(new_n12661_));
  AND2X1   g11659(.A(new_n12661_), .B(new_n12654_), .Y(new_n12662_));
  XOR2X1   g11660(.A(new_n12662_), .B(new_n12640_), .Y(new_n12663_));
  XOR2X1   g11661(.A(new_n12663_), .B(new_n12616_), .Y(new_n12664_));
  XOR2X1   g11662(.A(new_n12664_), .B(new_n12603_), .Y(new_n12665_));
  XOR2X1   g11663(.A(new_n12665_), .B(new_n12543_), .Y(new_n12666_));
  OAI22X1  g11664(.A0(new_n11818_), .A1(new_n11234_), .B0(new_n11065_), .B1(new_n11063_), .Y(new_n12667_));
  OR2X1    g11665(.A(new_n11819_), .B(new_n11233_), .Y(new_n12668_));
  XOR2X1   g11666(.A(new_n11168_), .B(new_n11075_), .Y(new_n12669_));
  OAI22X1  g11667(.A0(new_n11225_), .A1(new_n12669_), .B0(new_n11813_), .B1(new_n11812_), .Y(new_n12670_));
  OR2X1    g11668(.A(new_n11826_), .B(new_n11825_), .Y(new_n12671_));
  AND2X1   g11669(.A(new_n12671_), .B(new_n12670_), .Y(new_n12672_));
  XOR2X1   g11670(.A(new_n11925_), .B(new_n12672_), .Y(new_n12673_));
  AOI22X1  g11671(.A0(new_n12673_), .A1(new_n11978_), .B0(new_n12668_), .B1(new_n12667_), .Y(new_n12674_));
  OAI22X1  g11672(.A0(new_n11332_), .A1(new_n11932_), .B0(new_n11237_), .B1(new_n11236_), .Y(new_n12675_));
  NAND2X1  g11673(.A(new_n11332_), .B(new_n11932_), .Y(new_n12676_));
  AND2X1   g11674(.A(new_n12676_), .B(new_n12675_), .Y(new_n12677_));
  XOR2X1   g11675(.A(new_n11977_), .B(new_n12677_), .Y(new_n12678_));
  OAI21X1  g11676(.A0(new_n11925_), .A1(new_n11828_), .B0(new_n12678_), .Y(new_n12679_));
  NOR2X1   g11677(.A(new_n12679_), .B(new_n11926_), .Y(new_n12680_));
  OR2X1    g11678(.A(new_n12680_), .B(new_n12674_), .Y(new_n12681_));
  XOR2X1   g11679(.A(new_n11892_), .B(new_n11920_), .Y(new_n12682_));
  AOI22X1  g11680(.A0(new_n12682_), .A1(new_n11917_), .B0(new_n12671_), .B1(new_n12670_), .Y(new_n12683_));
  AOI21X1  g11681(.A0(new_n11901_), .A1(new_n11900_), .B0(new_n11912_), .Y(new_n12684_));
  NOR2X1   g11682(.A(new_n11915_), .B(new_n11914_), .Y(new_n12685_));
  AOI21X1  g11683(.A0(new_n12685_), .A1(new_n11900_), .B0(new_n12684_), .Y(new_n12686_));
  OAI21X1  g11684(.A0(new_n11922_), .A1(new_n11920_), .B0(new_n12686_), .Y(new_n12687_));
  NOR2X1   g11685(.A(new_n12687_), .B(new_n11893_), .Y(new_n12688_));
  AOI22X1  g11686(.A0(new_n11889_), .A1(new_n11888_), .B0(new_n11887_), .B1(new_n11886_), .Y(new_n12689_));
  NOR4X1   g11687(.A(new_n11883_), .B(new_n11882_), .C(new_n11872_), .D(new_n11869_), .Y(new_n12690_));
  OAI22X1  g11688(.A0(new_n12690_), .A1(new_n12689_), .B0(new_n11866_), .B1(new_n11858_), .Y(new_n12691_));
  OAI21X1  g11689(.A0(new_n11919_), .A1(new_n11918_), .B0(new_n12691_), .Y(new_n12692_));
  OR4X1    g11690(.A(new_n12690_), .B(new_n12689_), .C(new_n11866_), .D(new_n11858_), .Y(new_n12693_));
  NOR4X1   g11691(.A(new_n11880_), .B(new_n11879_), .C(new_n11875_), .D(new_n11874_), .Y(new_n12694_));
  AOI21X1  g11692(.A0(new_n11887_), .A1(new_n11886_), .B0(new_n12694_), .Y(new_n12695_));
  OAI22X1  g11693(.A0(new_n11880_), .A1(new_n11879_), .B0(new_n11875_), .B1(new_n11874_), .Y(new_n12696_));
  INVX1    g11694(.A(new_n12696_), .Y(new_n12697_));
  NOR2X1   g11695(.A(new_n12697_), .B(new_n12695_), .Y(new_n12698_));
  AND2X1   g11696(.A(new_n11864_), .B(new_n11861_), .Y(new_n12699_));
  AOI22X1  g11697(.A0(new_n11863_), .A1(new_n11862_), .B0(new_n11845_), .B1(new_n11840_), .Y(new_n12700_));
  OR2X1    g11698(.A(new_n12700_), .B(new_n12699_), .Y(new_n12701_));
  XOR2X1   g11699(.A(new_n12701_), .B(new_n12698_), .Y(new_n12702_));
  AOI21X1  g11700(.A0(new_n12693_), .A1(new_n12692_), .B0(new_n12702_), .Y(new_n12703_));
  AOI22X1  g11701(.A0(new_n11921_), .A1(new_n11867_), .B0(new_n11835_), .B1(new_n11834_), .Y(new_n12704_));
  NOR4X1   g11702(.A(new_n12690_), .B(new_n12689_), .C(new_n11866_), .D(new_n11858_), .Y(new_n12705_));
  NOR2X1   g11703(.A(new_n12701_), .B(new_n12698_), .Y(new_n12706_));
  AND2X1   g11704(.A(new_n12701_), .B(new_n12698_), .Y(new_n12707_));
  NOR4X1   g11705(.A(new_n12707_), .B(new_n12706_), .C(new_n12705_), .D(new_n12704_), .Y(new_n12708_));
  NOR4X1   g11706(.A(new_n11910_), .B(new_n11908_), .C(new_n11905_), .D(new_n11904_), .Y(new_n12709_));
  OAI22X1  g11707(.A0(new_n12709_), .A1(new_n11902_), .B0(new_n11913_), .B1(new_n11906_), .Y(new_n12710_));
  NOR3X1   g11708(.A(new_n12710_), .B(new_n12708_), .C(new_n12703_), .Y(new_n12711_));
  OAI22X1  g11709(.A0(new_n12707_), .A1(new_n12706_), .B0(new_n12705_), .B1(new_n12704_), .Y(new_n12712_));
  OR4X1    g11710(.A(new_n12707_), .B(new_n12706_), .C(new_n12705_), .D(new_n12704_), .Y(new_n12713_));
  AOI21X1  g11711(.A0(new_n11901_), .A1(new_n11900_), .B0(new_n12709_), .Y(new_n12714_));
  NOR2X1   g11712(.A(new_n11913_), .B(new_n11906_), .Y(new_n12715_));
  NOR2X1   g11713(.A(new_n12715_), .B(new_n12714_), .Y(new_n12716_));
  AOI21X1  g11714(.A0(new_n12713_), .A1(new_n12712_), .B0(new_n12716_), .Y(new_n12717_));
  OAI22X1  g11715(.A0(new_n12717_), .A1(new_n12711_), .B0(new_n12688_), .B1(new_n12683_), .Y(new_n12718_));
  OR4X1    g11716(.A(new_n12717_), .B(new_n12711_), .C(new_n12688_), .D(new_n12683_), .Y(new_n12719_));
  AND2X1   g11717(.A(new_n12719_), .B(new_n12718_), .Y(new_n12720_));
  AND2X1   g11718(.A(new_n11946_), .B(new_n11937_), .Y(new_n12721_));
  NOR4X1   g11719(.A(new_n11953_), .B(new_n11952_), .C(new_n11950_), .D(new_n11948_), .Y(new_n12722_));
  AND2X1   g11720(.A(new_n11967_), .B(new_n11958_), .Y(new_n12723_));
  NOR4X1   g11721(.A(new_n11974_), .B(new_n11973_), .C(new_n11971_), .D(new_n11969_), .Y(new_n12724_));
  OAI22X1  g11722(.A0(new_n12724_), .A1(new_n12723_), .B0(new_n12722_), .B1(new_n12721_), .Y(new_n12725_));
  OAI21X1  g11723(.A0(new_n11933_), .A1(new_n11930_), .B0(new_n12725_), .Y(new_n12726_));
  NAND4X1  g11724(.A(new_n11975_), .B(new_n11968_), .C(new_n11954_), .D(new_n11947_), .Y(new_n12727_));
  OR4X1    g11725(.A(new_n11965_), .B(new_n11964_), .C(new_n11961_), .D(new_n11960_), .Y(new_n12728_));
  AND2X1   g11726(.A(new_n12728_), .B(new_n11958_), .Y(new_n12729_));
  AND2X1   g11727(.A(new_n11966_), .B(new_n11962_), .Y(new_n12730_));
  OR2X1    g11728(.A(new_n12730_), .B(new_n12729_), .Y(new_n12731_));
  OR4X1    g11729(.A(new_n11944_), .B(new_n11943_), .C(new_n11940_), .D(new_n11939_), .Y(new_n12732_));
  AND2X1   g11730(.A(new_n11945_), .B(new_n11941_), .Y(new_n12733_));
  AOI21X1  g11731(.A0(new_n12732_), .A1(new_n11937_), .B0(new_n12733_), .Y(new_n12734_));
  XOR2X1   g11732(.A(new_n12734_), .B(new_n12731_), .Y(new_n12735_));
  AOI21X1  g11733(.A0(new_n12727_), .A1(new_n12726_), .B0(new_n12735_), .Y(new_n12736_));
  AOI22X1  g11734(.A0(new_n11975_), .A1(new_n11968_), .B0(new_n11954_), .B1(new_n11947_), .Y(new_n12737_));
  AOI21X1  g11735(.A0(new_n12676_), .A1(new_n12675_), .B0(new_n12737_), .Y(new_n12738_));
  NOR4X1   g11736(.A(new_n12724_), .B(new_n12723_), .C(new_n12722_), .D(new_n12721_), .Y(new_n12739_));
  AOI21X1  g11737(.A0(new_n12728_), .A1(new_n11958_), .B0(new_n12730_), .Y(new_n12740_));
  AND2X1   g11738(.A(new_n12732_), .B(new_n11937_), .Y(new_n12741_));
  NOR3X1   g11739(.A(new_n12733_), .B(new_n12741_), .C(new_n12740_), .Y(new_n12742_));
  NOR3X1   g11740(.A(new_n12734_), .B(new_n12730_), .C(new_n12729_), .Y(new_n12743_));
  NOR4X1   g11741(.A(new_n12743_), .B(new_n12742_), .C(new_n12739_), .D(new_n12738_), .Y(new_n12744_));
  OR2X1    g11742(.A(new_n12744_), .B(new_n12736_), .Y(new_n12745_));
  NAND3X1  g11743(.A(new_n12745_), .B(new_n12719_), .C(new_n12718_), .Y(new_n12746_));
  OAI21X1  g11744(.A0(new_n12745_), .A1(new_n12720_), .B0(new_n12746_), .Y(new_n12747_));
  XOR2X1   g11745(.A(new_n12747_), .B(new_n12681_), .Y(new_n12748_));
  XOR2X1   g11746(.A(new_n12748_), .B(new_n12666_), .Y(new_n12749_));
  AND2X1   g11747(.A(new_n12749_), .B(new_n12532_), .Y(new_n12750_));
  XOR2X1   g11748(.A(new_n12749_), .B(new_n12532_), .Y(new_n12751_));
  OAI22X1  g11749(.A0(new_n11778_), .A1(new_n12296_), .B0(new_n12276_), .B1(new_n12275_), .Y(new_n12752_));
  NAND2X1  g11750(.A(new_n11778_), .B(new_n12296_), .Y(new_n12753_));
  AND2X1   g11751(.A(new_n12753_), .B(new_n12752_), .Y(new_n12754_));
  XOR2X1   g11752(.A(new_n12397_), .B(new_n12754_), .Y(new_n12755_));
  OAI22X1  g11753(.A0(new_n12524_), .A1(new_n12755_), .B0(new_n12286_), .B1(new_n12279_), .Y(new_n12756_));
  AOI21X1  g11754(.A0(new_n10400_), .A1(new_n10333_), .B0(new_n10273_), .Y(new_n12757_));
  NOR2X1   g11755(.A(new_n10400_), .B(new_n10333_), .Y(new_n12758_));
  OR2X1    g11756(.A(new_n12758_), .B(new_n12757_), .Y(new_n12759_));
  XOR2X1   g11757(.A(new_n11556_), .B(new_n12759_), .Y(new_n12760_));
  AOI22X1  g11758(.A0(new_n12760_), .A1(new_n11453_), .B0(new_n12283_), .B1(new_n12282_), .Y(new_n12761_));
  AND2X1   g11759(.A(new_n11557_), .B(new_n12404_), .Y(new_n12762_));
  OR2X1    g11760(.A(new_n12762_), .B(new_n12761_), .Y(new_n12763_));
  XOR2X1   g11761(.A(new_n12523_), .B(new_n12763_), .Y(new_n12764_));
  OR2X1    g11762(.A(new_n12764_), .B(new_n12398_), .Y(new_n12765_));
  AND2X1   g11763(.A(new_n12765_), .B(new_n12756_), .Y(new_n12766_));
  OR2X1    g11764(.A(new_n12491_), .B(new_n12490_), .Y(new_n12767_));
  XOR2X1   g11765(.A(new_n11450_), .B(new_n12767_), .Y(new_n12768_));
  AOI22X1  g11766(.A0(new_n12768_), .A1(new_n11402_), .B0(new_n12402_), .B1(new_n12401_), .Y(new_n12769_));
  AND2X1   g11767(.A(new_n11451_), .B(new_n12470_), .Y(new_n12770_));
  OR2X1    g11768(.A(new_n12770_), .B(new_n12769_), .Y(new_n12771_));
  XOR2X1   g11769(.A(new_n12521_), .B(new_n12771_), .Y(new_n12772_));
  AOI22X1  g11770(.A0(new_n12772_), .A1(new_n12464_), .B0(new_n12406_), .B1(new_n12405_), .Y(new_n12773_));
  NOR2X1   g11771(.A(new_n12772_), .B(new_n12464_), .Y(new_n12774_));
  OR2X1    g11772(.A(new_n12774_), .B(new_n12773_), .Y(new_n12775_));
  AOI22X1  g11773(.A0(new_n12519_), .A1(new_n12513_), .B0(new_n12497_), .B1(new_n12489_), .Y(new_n12776_));
  AOI21X1  g11774(.A0(new_n12472_), .A1(new_n12471_), .B0(new_n12776_), .Y(new_n12777_));
  AOI22X1  g11775(.A0(new_n12496_), .A1(new_n12495_), .B0(new_n12494_), .B1(new_n12493_), .Y(new_n12778_));
  NOR4X1   g11776(.A(new_n12488_), .B(new_n12486_), .C(new_n12477_), .D(new_n12475_), .Y(new_n12779_));
  AOI22X1  g11777(.A0(new_n12518_), .A1(new_n12517_), .B0(new_n12516_), .B1(new_n12515_), .Y(new_n12780_));
  NOR4X1   g11778(.A(new_n12512_), .B(new_n12511_), .C(new_n12503_), .D(new_n12500_), .Y(new_n12781_));
  NOR4X1   g11779(.A(new_n12781_), .B(new_n12780_), .C(new_n12779_), .D(new_n12778_), .Y(new_n12782_));
  OR4X1    g11780(.A(new_n12509_), .B(new_n12508_), .C(new_n12506_), .D(new_n12505_), .Y(new_n12783_));
  OAI21X1  g11781(.A0(new_n12503_), .A1(new_n12500_), .B0(new_n12783_), .Y(new_n12784_));
  OAI22X1  g11782(.A0(new_n12509_), .A1(new_n12508_), .B0(new_n12506_), .B1(new_n12505_), .Y(new_n12785_));
  AND2X1   g11783(.A(new_n12785_), .B(new_n12784_), .Y(new_n12786_));
  OR4X1    g11784(.A(new_n12484_), .B(new_n12483_), .C(new_n12480_), .D(new_n12479_), .Y(new_n12787_));
  OAI21X1  g11785(.A0(new_n12477_), .A1(new_n12475_), .B0(new_n12787_), .Y(new_n12788_));
  OAI22X1  g11786(.A0(new_n12484_), .A1(new_n12483_), .B0(new_n12480_), .B1(new_n12479_), .Y(new_n12789_));
  AND2X1   g11787(.A(new_n12789_), .B(new_n12788_), .Y(new_n12790_));
  XOR2X1   g11788(.A(new_n12790_), .B(new_n12786_), .Y(new_n12791_));
  OAI21X1  g11789(.A0(new_n12782_), .A1(new_n12777_), .B0(new_n12791_), .Y(new_n12792_));
  OAI22X1  g11790(.A0(new_n12781_), .A1(new_n12780_), .B0(new_n12779_), .B1(new_n12778_), .Y(new_n12793_));
  OAI21X1  g11791(.A0(new_n12770_), .A1(new_n12769_), .B0(new_n12793_), .Y(new_n12794_));
  NAND2X1  g11792(.A(new_n12785_), .B(new_n12784_), .Y(new_n12795_));
  OR2X1    g11793(.A(new_n12790_), .B(new_n12795_), .Y(new_n12796_));
  AOI21X1  g11794(.A0(new_n12790_), .A1(new_n12795_), .B0(new_n12782_), .Y(new_n12797_));
  NAND3X1  g11795(.A(new_n12797_), .B(new_n12796_), .C(new_n12794_), .Y(new_n12798_));
  NAND2X1  g11796(.A(new_n12798_), .B(new_n12792_), .Y(new_n12799_));
  OAI22X1  g11797(.A0(new_n11555_), .A1(new_n12417_), .B0(new_n12758_), .B1(new_n12757_), .Y(new_n12800_));
  NAND2X1  g11798(.A(new_n11555_), .B(new_n12417_), .Y(new_n12801_));
  AOI22X1  g11799(.A0(new_n12461_), .A1(new_n12455_), .B0(new_n12439_), .B1(new_n12432_), .Y(new_n12802_));
  AOI21X1  g11800(.A0(new_n12801_), .A1(new_n12800_), .B0(new_n12802_), .Y(new_n12803_));
  AND2X1   g11801(.A(new_n12431_), .B(new_n12422_), .Y(new_n12804_));
  NOR4X1   g11802(.A(new_n12438_), .B(new_n12437_), .C(new_n12435_), .D(new_n12433_), .Y(new_n12805_));
  AOI22X1  g11803(.A0(new_n12460_), .A1(new_n12459_), .B0(new_n12458_), .B1(new_n12457_), .Y(new_n12806_));
  NOR4X1   g11804(.A(new_n12454_), .B(new_n12453_), .C(new_n12445_), .D(new_n12442_), .Y(new_n12807_));
  NOR4X1   g11805(.A(new_n12807_), .B(new_n12806_), .C(new_n12805_), .D(new_n12804_), .Y(new_n12808_));
  OR4X1    g11806(.A(new_n12451_), .B(new_n12450_), .C(new_n12448_), .D(new_n12447_), .Y(new_n12809_));
  OAI21X1  g11807(.A0(new_n12445_), .A1(new_n12442_), .B0(new_n12809_), .Y(new_n12810_));
  OAI22X1  g11808(.A0(new_n12451_), .A1(new_n12450_), .B0(new_n12448_), .B1(new_n12447_), .Y(new_n12811_));
  AND2X1   g11809(.A(new_n12811_), .B(new_n12810_), .Y(new_n12812_));
  OR4X1    g11810(.A(new_n12429_), .B(new_n12428_), .C(new_n12425_), .D(new_n12424_), .Y(new_n12813_));
  AOI22X1  g11811(.A0(new_n12813_), .A1(new_n12422_), .B0(new_n12430_), .B1(new_n12426_), .Y(new_n12814_));
  XOR2X1   g11812(.A(new_n12814_), .B(new_n12812_), .Y(new_n12815_));
  OAI21X1  g11813(.A0(new_n12808_), .A1(new_n12803_), .B0(new_n12815_), .Y(new_n12816_));
  OAI22X1  g11814(.A0(new_n12807_), .A1(new_n12806_), .B0(new_n12805_), .B1(new_n12804_), .Y(new_n12817_));
  OAI21X1  g11815(.A0(new_n12418_), .A1(new_n12411_), .B0(new_n12817_), .Y(new_n12818_));
  NAND4X1  g11816(.A(new_n12461_), .B(new_n12455_), .C(new_n12439_), .D(new_n12432_), .Y(new_n12819_));
  NAND2X1  g11817(.A(new_n12811_), .B(new_n12810_), .Y(new_n12820_));
  NAND2X1  g11818(.A(new_n12814_), .B(new_n12820_), .Y(new_n12821_));
  OR2X1    g11819(.A(new_n12814_), .B(new_n12820_), .Y(new_n12822_));
  NAND4X1  g11820(.A(new_n12822_), .B(new_n12821_), .C(new_n12819_), .D(new_n12818_), .Y(new_n12823_));
  AND2X1   g11821(.A(new_n12823_), .B(new_n12816_), .Y(new_n12824_));
  XOR2X1   g11822(.A(new_n12824_), .B(new_n12799_), .Y(new_n12825_));
  XOR2X1   g11823(.A(new_n12825_), .B(new_n12775_), .Y(new_n12826_));
  OAI22X1  g11824(.A0(new_n11776_), .A1(new_n12305_), .B0(new_n12289_), .B1(new_n12288_), .Y(new_n12827_));
  NAND2X1  g11825(.A(new_n11776_), .B(new_n12305_), .Y(new_n12828_));
  AND2X1   g11826(.A(new_n12828_), .B(new_n12827_), .Y(new_n12829_));
  XOR2X1   g11827(.A(new_n12346_), .B(new_n12829_), .Y(new_n12830_));
  OAI22X1  g11828(.A0(new_n12396_), .A1(new_n12830_), .B0(new_n12297_), .B1(new_n12292_), .Y(new_n12831_));
  AND2X1   g11829(.A(new_n11623_), .B(new_n11622_), .Y(new_n12832_));
  OR2X1    g11830(.A(new_n11624_), .B(new_n12832_), .Y(new_n12833_));
  XOR2X1   g11831(.A(new_n11667_), .B(new_n12833_), .Y(new_n12834_));
  AOI21X1  g11832(.A0(new_n12834_), .A1(new_n11621_), .B0(new_n12295_), .Y(new_n12835_));
  AND2X1   g11833(.A(new_n11668_), .B(new_n12349_), .Y(new_n12836_));
  OR2X1    g11834(.A(new_n12836_), .B(new_n12835_), .Y(new_n12837_));
  XOR2X1   g11835(.A(new_n12395_), .B(new_n12837_), .Y(new_n12838_));
  OR2X1    g11836(.A(new_n12838_), .B(new_n12347_), .Y(new_n12839_));
  AND2X1   g11837(.A(new_n12839_), .B(new_n12831_), .Y(new_n12840_));
  AOI22X1  g11838(.A0(new_n12393_), .A1(new_n12386_), .B0(new_n12372_), .B1(new_n12365_), .Y(new_n12841_));
  AOI21X1  g11839(.A0(new_n12351_), .A1(new_n12350_), .B0(new_n12841_), .Y(new_n12842_));
  AND2X1   g11840(.A(new_n12364_), .B(new_n12355_), .Y(new_n12843_));
  NOR4X1   g11841(.A(new_n12371_), .B(new_n12370_), .C(new_n12368_), .D(new_n12366_), .Y(new_n12844_));
  AND2X1   g11842(.A(new_n12385_), .B(new_n12376_), .Y(new_n12845_));
  NOR4X1   g11843(.A(new_n12392_), .B(new_n12391_), .C(new_n12389_), .D(new_n12387_), .Y(new_n12846_));
  NOR4X1   g11844(.A(new_n12846_), .B(new_n12845_), .C(new_n12844_), .D(new_n12843_), .Y(new_n12847_));
  OR4X1    g11845(.A(new_n12383_), .B(new_n12382_), .C(new_n12379_), .D(new_n12378_), .Y(new_n12848_));
  AOI22X1  g11846(.A0(new_n12848_), .A1(new_n12376_), .B0(new_n12384_), .B1(new_n12380_), .Y(new_n12849_));
  OR4X1    g11847(.A(new_n12362_), .B(new_n12361_), .C(new_n12358_), .D(new_n12357_), .Y(new_n12850_));
  AOI22X1  g11848(.A0(new_n12850_), .A1(new_n12355_), .B0(new_n12363_), .B1(new_n12359_), .Y(new_n12851_));
  XOR2X1   g11849(.A(new_n12851_), .B(new_n12849_), .Y(new_n12852_));
  OAI21X1  g11850(.A0(new_n12847_), .A1(new_n12842_), .B0(new_n12852_), .Y(new_n12853_));
  OAI22X1  g11851(.A0(new_n12846_), .A1(new_n12845_), .B0(new_n12844_), .B1(new_n12843_), .Y(new_n12854_));
  OAI21X1  g11852(.A0(new_n12836_), .A1(new_n12835_), .B0(new_n12854_), .Y(new_n12855_));
  NAND2X1  g11853(.A(new_n12848_), .B(new_n12376_), .Y(new_n12856_));
  OAI22X1  g11854(.A0(new_n12383_), .A1(new_n12382_), .B0(new_n12379_), .B1(new_n12378_), .Y(new_n12857_));
  NAND2X1  g11855(.A(new_n12857_), .B(new_n12856_), .Y(new_n12858_));
  OR2X1    g11856(.A(new_n12851_), .B(new_n12858_), .Y(new_n12859_));
  AOI21X1  g11857(.A0(new_n12851_), .A1(new_n12858_), .B0(new_n12847_), .Y(new_n12860_));
  NAND3X1  g11858(.A(new_n12860_), .B(new_n12859_), .C(new_n12855_), .Y(new_n12861_));
  NAND2X1  g11859(.A(new_n12861_), .B(new_n12853_), .Y(new_n12862_));
  AOI22X1  g11860(.A0(new_n12344_), .A1(new_n12339_), .B0(new_n12325_), .B1(new_n12321_), .Y(new_n12863_));
  AOI21X1  g11861(.A0(new_n12828_), .A1(new_n12827_), .B0(new_n12863_), .Y(new_n12864_));
  NAND3X1  g11862(.A(new_n12344_), .B(new_n12325_), .C(new_n12321_), .Y(new_n12865_));
  AOI21X1  g11863(.A0(new_n12338_), .A1(new_n12329_), .B0(new_n12865_), .Y(new_n12866_));
  OR4X1    g11864(.A(new_n12336_), .B(new_n12335_), .C(new_n12332_), .D(new_n12331_), .Y(new_n12867_));
  AOI22X1  g11865(.A0(new_n12867_), .A1(new_n12329_), .B0(new_n12337_), .B1(new_n12333_), .Y(new_n12868_));
  OR4X1    g11866(.A(new_n12318_), .B(new_n12317_), .C(new_n12315_), .D(new_n12314_), .Y(new_n12869_));
  OAI21X1  g11867(.A0(new_n12312_), .A1(new_n12309_), .B0(new_n12869_), .Y(new_n12870_));
  OAI22X1  g11868(.A0(new_n12318_), .A1(new_n12317_), .B0(new_n12315_), .B1(new_n12314_), .Y(new_n12871_));
  AND2X1   g11869(.A(new_n12871_), .B(new_n12870_), .Y(new_n12872_));
  XOR2X1   g11870(.A(new_n12872_), .B(new_n12868_), .Y(new_n12873_));
  OAI21X1  g11871(.A0(new_n12866_), .A1(new_n12864_), .B0(new_n12873_), .Y(new_n12874_));
  AND2X1   g11872(.A(new_n12325_), .B(new_n12321_), .Y(new_n12875_));
  OAI22X1  g11873(.A0(new_n12345_), .A1(new_n12875_), .B0(new_n12306_), .B1(new_n12303_), .Y(new_n12876_));
  NAND4X1  g11874(.A(new_n12344_), .B(new_n12339_), .C(new_n12325_), .D(new_n12321_), .Y(new_n12877_));
  NAND2X1  g11875(.A(new_n12867_), .B(new_n12329_), .Y(new_n12878_));
  OAI22X1  g11876(.A0(new_n12336_), .A1(new_n12335_), .B0(new_n12332_), .B1(new_n12331_), .Y(new_n12879_));
  NAND2X1  g11877(.A(new_n12879_), .B(new_n12878_), .Y(new_n12880_));
  NAND2X1  g11878(.A(new_n12872_), .B(new_n12880_), .Y(new_n12881_));
  OR2X1    g11879(.A(new_n12872_), .B(new_n12880_), .Y(new_n12882_));
  NAND4X1  g11880(.A(new_n12882_), .B(new_n12881_), .C(new_n12877_), .D(new_n12876_), .Y(new_n12883_));
  AND2X1   g11881(.A(new_n12883_), .B(new_n12874_), .Y(new_n12884_));
  XOR2X1   g11882(.A(new_n12884_), .B(new_n12862_), .Y(new_n12885_));
  XOR2X1   g11883(.A(new_n12885_), .B(new_n12840_), .Y(new_n12886_));
  XOR2X1   g11884(.A(new_n12886_), .B(new_n12826_), .Y(new_n12887_));
  XOR2X1   g11885(.A(new_n12887_), .B(new_n12766_), .Y(new_n12888_));
  NOR2X1   g11886(.A(new_n12888_), .B(new_n12751_), .Y(new_n12889_));
  OAI21X1  g11887(.A0(new_n12749_), .A1(new_n12532_), .B0(new_n12888_), .Y(new_n12890_));
  OAI22X1  g11888(.A0(new_n12890_), .A1(new_n12750_), .B0(new_n12889_), .B1(new_n12529_), .Y(new_n12891_));
  NOR2X1   g11889(.A(new_n12268_), .B(new_n11982_), .Y(new_n12892_));
  NAND2X1  g11890(.A(new_n12268_), .B(new_n11982_), .Y(new_n12893_));
  OAI21X1  g11891(.A0(new_n12892_), .A1(new_n12273_), .B0(new_n12893_), .Y(new_n12894_));
  AOI22X1  g11892(.A0(new_n9621_), .A1(new_n9438_), .B0(new_n9246_), .B1(new_n9236_), .Y(new_n12895_));
  NOR2X1   g11893(.A(new_n9621_), .B(new_n9438_), .Y(new_n12896_));
  OR2X1    g11894(.A(new_n12896_), .B(new_n12895_), .Y(new_n12897_));
  XOR2X1   g11895(.A(new_n11054_), .B(new_n12897_), .Y(new_n12898_));
  AOI22X1  g11896(.A0(new_n12898_), .A1(new_n10806_), .B0(new_n11801_), .B1(new_n11800_), .Y(new_n12899_));
  AND2X1   g11897(.A(new_n11055_), .B(new_n11990_), .Y(new_n12900_));
  OAI22X1  g11898(.A0(new_n11053_), .A1(new_n12010_), .B0(new_n12896_), .B1(new_n12895_), .Y(new_n12901_));
  NAND2X1  g11899(.A(new_n11053_), .B(new_n12010_), .Y(new_n12902_));
  AND2X1   g11900(.A(new_n12902_), .B(new_n12901_), .Y(new_n12903_));
  XOR2X1   g11901(.A(new_n12131_), .B(new_n12903_), .Y(new_n12904_));
  OAI22X1  g11902(.A0(new_n12266_), .A1(new_n12904_), .B0(new_n12900_), .B1(new_n12899_), .Y(new_n12905_));
  OR2X1    g11903(.A(new_n12540_), .B(new_n12132_), .Y(new_n12906_));
  AND2X1   g11904(.A(new_n12906_), .B(new_n12905_), .Y(new_n12907_));
  XOR2X1   g11905(.A(new_n12665_), .B(new_n12907_), .Y(new_n12908_));
  OR2X1    g11906(.A(new_n12748_), .B(new_n12908_), .Y(new_n12909_));
  AND2X1   g11907(.A(new_n12748_), .B(new_n12908_), .Y(new_n12910_));
  AOI21X1  g11908(.A0(new_n12909_), .A1(new_n12894_), .B0(new_n12910_), .Y(new_n12911_));
  NOR2X1   g11909(.A(new_n12744_), .B(new_n12736_), .Y(new_n12912_));
  OAI22X1  g11910(.A0(new_n12912_), .A1(new_n12720_), .B0(new_n12680_), .B1(new_n12674_), .Y(new_n12913_));
  NAND3X1  g11911(.A(new_n12912_), .B(new_n12719_), .C(new_n12718_), .Y(new_n12914_));
  AND2X1   g11912(.A(new_n12914_), .B(new_n12913_), .Y(new_n12915_));
  OR4X1    g11913(.A(new_n12733_), .B(new_n12741_), .C(new_n12730_), .D(new_n12729_), .Y(new_n12916_));
  OAI21X1  g11914(.A0(new_n12739_), .A1(new_n12738_), .B0(new_n12916_), .Y(new_n12917_));
  OR2X1    g11915(.A(new_n12734_), .B(new_n12740_), .Y(new_n12918_));
  NAND2X1  g11916(.A(new_n12918_), .B(new_n12917_), .Y(new_n12919_));
  OAI21X1  g11917(.A0(new_n12708_), .A1(new_n12703_), .B0(new_n12716_), .Y(new_n12920_));
  OAI21X1  g11918(.A0(new_n12688_), .A1(new_n12683_), .B0(new_n12920_), .Y(new_n12921_));
  NAND3X1  g11919(.A(new_n12710_), .B(new_n12713_), .C(new_n12712_), .Y(new_n12922_));
  OR4X1    g11920(.A(new_n12700_), .B(new_n12697_), .C(new_n12695_), .D(new_n12699_), .Y(new_n12923_));
  OAI21X1  g11921(.A0(new_n12705_), .A1(new_n12704_), .B0(new_n12923_), .Y(new_n12924_));
  OAI22X1  g11922(.A0(new_n12700_), .A1(new_n12699_), .B0(new_n12697_), .B1(new_n12695_), .Y(new_n12925_));
  NAND2X1  g11923(.A(new_n12925_), .B(new_n12924_), .Y(new_n12926_));
  AOI21X1  g11924(.A0(new_n12922_), .A1(new_n12921_), .B0(new_n12926_), .Y(new_n12927_));
  OAI22X1  g11925(.A0(new_n11924_), .A1(new_n12686_), .B0(new_n11827_), .B1(new_n11824_), .Y(new_n12928_));
  OR2X1    g11926(.A(new_n12687_), .B(new_n11893_), .Y(new_n12929_));
  AOI21X1  g11927(.A0(new_n12713_), .A1(new_n12712_), .B0(new_n12710_), .Y(new_n12930_));
  AOI21X1  g11928(.A0(new_n12929_), .A1(new_n12928_), .B0(new_n12930_), .Y(new_n12931_));
  NOR3X1   g11929(.A(new_n12716_), .B(new_n12708_), .C(new_n12703_), .Y(new_n12932_));
  AND2X1   g11930(.A(new_n12925_), .B(new_n12924_), .Y(new_n12933_));
  NOR3X1   g11931(.A(new_n12933_), .B(new_n12932_), .C(new_n12931_), .Y(new_n12934_));
  OAI21X1  g11932(.A0(new_n12934_), .A1(new_n12927_), .B0(new_n12919_), .Y(new_n12935_));
  AND2X1   g11933(.A(new_n12918_), .B(new_n12917_), .Y(new_n12936_));
  OAI21X1  g11934(.A0(new_n12932_), .A1(new_n12931_), .B0(new_n12933_), .Y(new_n12937_));
  NAND3X1  g11935(.A(new_n12926_), .B(new_n12922_), .C(new_n12921_), .Y(new_n12938_));
  NAND3X1  g11936(.A(new_n12938_), .B(new_n12937_), .C(new_n12936_), .Y(new_n12939_));
  AND2X1   g11937(.A(new_n12939_), .B(new_n12935_), .Y(new_n12940_));
  XOR2X1   g11938(.A(new_n12940_), .B(new_n12915_), .Y(new_n12941_));
  AND2X1   g11939(.A(new_n12578_), .B(new_n12577_), .Y(new_n12942_));
  XOR2X1   g11940(.A(new_n12204_), .B(new_n12942_), .Y(new_n12943_));
  OAI22X1  g11941(.A0(new_n12264_), .A1(new_n12943_), .B0(new_n12538_), .B1(new_n12537_), .Y(new_n12944_));
  OR2X1    g11942(.A(new_n12549_), .B(new_n12205_), .Y(new_n12945_));
  AND2X1   g11943(.A(new_n12945_), .B(new_n12944_), .Y(new_n12946_));
  XOR2X1   g11944(.A(new_n12602_), .B(new_n12946_), .Y(new_n12947_));
  OAI22X1  g11945(.A0(new_n12664_), .A1(new_n12947_), .B0(new_n12542_), .B1(new_n12541_), .Y(new_n12948_));
  NAND2X1  g11946(.A(new_n12664_), .B(new_n12947_), .Y(new_n12949_));
  AND2X1   g11947(.A(new_n12949_), .B(new_n12948_), .Y(new_n12950_));
  AOI22X1  g11948(.A0(new_n12661_), .A1(new_n12654_), .B0(new_n12639_), .B1(new_n12633_), .Y(new_n12951_));
  AOI21X1  g11949(.A0(new_n12615_), .A1(new_n12608_), .B0(new_n12951_), .Y(new_n12952_));
  AOI22X1  g11950(.A0(new_n12660_), .A1(new_n12659_), .B0(new_n12657_), .B1(new_n12656_), .Y(new_n12953_));
  NAND3X1  g11951(.A(new_n12661_), .B(new_n12639_), .C(new_n12633_), .Y(new_n12954_));
  NOR2X1   g11952(.A(new_n12954_), .B(new_n12953_), .Y(new_n12955_));
  NAND4X1  g11953(.A(new_n12127_), .B(new_n12121_), .C(new_n12103_), .D(new_n12095_), .Y(new_n12956_));
  AND2X1   g11954(.A(new_n12630_), .B(new_n12626_), .Y(new_n12957_));
  AND2X1   g11955(.A(new_n12957_), .B(new_n12625_), .Y(new_n12958_));
  AOI22X1  g11956(.A0(new_n12958_), .A1(new_n12629_), .B0(new_n12956_), .B1(new_n12635_), .Y(new_n12959_));
  AOI22X1  g11957(.A0(new_n12630_), .A1(new_n12629_), .B0(new_n12626_), .B1(new_n12625_), .Y(new_n12960_));
  NOR2X1   g11958(.A(new_n12960_), .B(new_n12959_), .Y(new_n12961_));
  AOI22X1  g11959(.A0(new_n12059_), .A1(new_n12056_), .B0(new_n12037_), .B1(new_n12034_), .Y(new_n12962_));
  NAND2X1  g11960(.A(new_n12962_), .B(new_n12647_), .Y(new_n12963_));
  OAI22X1  g11961(.A0(new_n12963_), .A1(new_n12651_), .B0(new_n12645_), .B1(new_n12642_), .Y(new_n12964_));
  OAI21X1  g11962(.A0(new_n12652_), .A1(new_n12649_), .B0(new_n12964_), .Y(new_n12965_));
  NOR2X1   g11963(.A(new_n12965_), .B(new_n12961_), .Y(new_n12966_));
  AND2X1   g11964(.A(new_n12965_), .B(new_n12961_), .Y(new_n12967_));
  OAI22X1  g11965(.A0(new_n12967_), .A1(new_n12966_), .B0(new_n12955_), .B1(new_n12952_), .Y(new_n12968_));
  AOI22X1  g11966(.A0(new_n12614_), .A1(new_n12071_), .B0(new_n12902_), .B1(new_n12901_), .Y(new_n12969_));
  NOR2X1   g11967(.A(new_n12614_), .B(new_n12071_), .Y(new_n12970_));
  AND2X1   g11968(.A(new_n12639_), .B(new_n12633_), .Y(new_n12971_));
  OAI22X1  g11969(.A0(new_n12662_), .A1(new_n12971_), .B0(new_n12970_), .B1(new_n12969_), .Y(new_n12972_));
  NAND4X1  g11970(.A(new_n12661_), .B(new_n12654_), .C(new_n12639_), .D(new_n12633_), .Y(new_n12973_));
  OR2X1    g11971(.A(new_n12965_), .B(new_n12961_), .Y(new_n12974_));
  NAND2X1  g11972(.A(new_n12965_), .B(new_n12961_), .Y(new_n12975_));
  NAND4X1  g11973(.A(new_n12975_), .B(new_n12974_), .C(new_n12973_), .D(new_n12972_), .Y(new_n12976_));
  NAND2X1  g11974(.A(new_n12976_), .B(new_n12968_), .Y(new_n12977_));
  AOI22X1  g11975(.A0(new_n12600_), .A1(new_n12593_), .B0(new_n12575_), .B1(new_n12569_), .Y(new_n12978_));
  AOI21X1  g11976(.A0(new_n12945_), .A1(new_n12944_), .B0(new_n12978_), .Y(new_n12979_));
  AOI22X1  g11977(.A0(new_n12599_), .A1(new_n12598_), .B0(new_n12596_), .B1(new_n12595_), .Y(new_n12980_));
  NAND3X1  g11978(.A(new_n12600_), .B(new_n12575_), .C(new_n12569_), .Y(new_n12981_));
  NOR2X1   g11979(.A(new_n12981_), .B(new_n12980_), .Y(new_n12982_));
  NAND4X1  g11980(.A(new_n12261_), .B(new_n12255_), .C(new_n12237_), .D(new_n12229_), .Y(new_n12983_));
  AND2X1   g11981(.A(new_n12566_), .B(new_n12562_), .Y(new_n12984_));
  AND2X1   g11982(.A(new_n12984_), .B(new_n12561_), .Y(new_n12985_));
  AOI22X1  g11983(.A0(new_n12985_), .A1(new_n12565_), .B0(new_n12983_), .B1(new_n12571_), .Y(new_n12986_));
  AOI22X1  g11984(.A0(new_n12566_), .A1(new_n12565_), .B0(new_n12562_), .B1(new_n12561_), .Y(new_n12987_));
  NOR2X1   g11985(.A(new_n12987_), .B(new_n12986_), .Y(new_n12988_));
  AND2X1   g11986(.A(new_n12590_), .B(new_n12586_), .Y(new_n12989_));
  AND2X1   g11987(.A(new_n12989_), .B(new_n12585_), .Y(new_n12990_));
  AOI22X1  g11988(.A0(new_n12990_), .A1(new_n12589_), .B0(new_n12596_), .B1(new_n12595_), .Y(new_n12991_));
  AOI22X1  g11989(.A0(new_n12590_), .A1(new_n12589_), .B0(new_n12586_), .B1(new_n12585_), .Y(new_n12992_));
  OR2X1    g11990(.A(new_n12992_), .B(new_n12991_), .Y(new_n12993_));
  NOR2X1   g11991(.A(new_n12993_), .B(new_n12988_), .Y(new_n12994_));
  AND2X1   g11992(.A(new_n12993_), .B(new_n12988_), .Y(new_n12995_));
  OAI22X1  g11993(.A0(new_n12995_), .A1(new_n12994_), .B0(new_n12982_), .B1(new_n12979_), .Y(new_n12996_));
  AND2X1   g11994(.A(new_n12575_), .B(new_n12569_), .Y(new_n12997_));
  OAI22X1  g11995(.A0(new_n12601_), .A1(new_n12997_), .B0(new_n12551_), .B1(new_n12550_), .Y(new_n12998_));
  NAND4X1  g11996(.A(new_n12600_), .B(new_n12593_), .C(new_n12575_), .D(new_n12569_), .Y(new_n12999_));
  OR2X1    g11997(.A(new_n12993_), .B(new_n12988_), .Y(new_n13000_));
  NAND2X1  g11998(.A(new_n12993_), .B(new_n12988_), .Y(new_n13001_));
  NAND4X1  g11999(.A(new_n13001_), .B(new_n13000_), .C(new_n12999_), .D(new_n12998_), .Y(new_n13002_));
  AND2X1   g12000(.A(new_n13002_), .B(new_n12996_), .Y(new_n13003_));
  XOR2X1   g12001(.A(new_n13003_), .B(new_n12977_), .Y(new_n13004_));
  XOR2X1   g12002(.A(new_n13004_), .B(new_n12950_), .Y(new_n13005_));
  XOR2X1   g12003(.A(new_n13005_), .B(new_n12941_), .Y(new_n13006_));
  XOR2X1   g12004(.A(new_n13006_), .B(new_n12911_), .Y(new_n13007_));
  OAI22X1  g12005(.A0(new_n11780_), .A1(new_n12285_), .B0(new_n11345_), .B1(new_n11344_), .Y(new_n13008_));
  NAND2X1  g12006(.A(new_n11780_), .B(new_n12285_), .Y(new_n13009_));
  AOI22X1  g12007(.A0(new_n12764_), .A1(new_n12398_), .B0(new_n13009_), .B1(new_n13008_), .Y(new_n13010_));
  NOR2X1   g12008(.A(new_n12764_), .B(new_n12398_), .Y(new_n13011_));
  AND2X1   g12009(.A(new_n12801_), .B(new_n12800_), .Y(new_n13012_));
  XOR2X1   g12010(.A(new_n12463_), .B(new_n13012_), .Y(new_n13013_));
  OAI22X1  g12011(.A0(new_n12522_), .A1(new_n13013_), .B0(new_n12762_), .B1(new_n12761_), .Y(new_n13014_));
  OR2X1    g12012(.A(new_n12772_), .B(new_n12464_), .Y(new_n13015_));
  AND2X1   g12013(.A(new_n13015_), .B(new_n13014_), .Y(new_n13016_));
  XOR2X1   g12014(.A(new_n12825_), .B(new_n13016_), .Y(new_n13017_));
  OAI22X1  g12015(.A0(new_n12886_), .A1(new_n13017_), .B0(new_n13011_), .B1(new_n13010_), .Y(new_n13018_));
  NAND2X1  g12016(.A(new_n12886_), .B(new_n13017_), .Y(new_n13019_));
  AND2X1   g12017(.A(new_n13019_), .B(new_n13018_), .Y(new_n13020_));
  AOI22X1  g12018(.A0(new_n12883_), .A1(new_n12874_), .B0(new_n12861_), .B1(new_n12853_), .Y(new_n13021_));
  AOI21X1  g12019(.A0(new_n12839_), .A1(new_n12831_), .B0(new_n13021_), .Y(new_n13022_));
  AOI22X1  g12020(.A0(new_n12882_), .A1(new_n12881_), .B0(new_n12877_), .B1(new_n12876_), .Y(new_n13023_));
  NAND3X1  g12021(.A(new_n12883_), .B(new_n12861_), .C(new_n12853_), .Y(new_n13024_));
  NOR2X1   g12022(.A(new_n13024_), .B(new_n13023_), .Y(new_n13025_));
  NAND4X1  g12023(.A(new_n12393_), .B(new_n12386_), .C(new_n12372_), .D(new_n12365_), .Y(new_n13026_));
  NAND2X1  g12024(.A(new_n12850_), .B(new_n12355_), .Y(new_n13027_));
  AOI22X1  g12025(.A0(new_n12384_), .A1(new_n12380_), .B0(new_n12363_), .B1(new_n12359_), .Y(new_n13028_));
  AND2X1   g12026(.A(new_n13028_), .B(new_n12856_), .Y(new_n13029_));
  AOI22X1  g12027(.A0(new_n13029_), .A1(new_n13027_), .B0(new_n13026_), .B1(new_n12855_), .Y(new_n13030_));
  NOR2X1   g12028(.A(new_n12851_), .B(new_n12849_), .Y(new_n13031_));
  OR2X1    g12029(.A(new_n13031_), .B(new_n13030_), .Y(new_n13032_));
  NAND2X1  g12030(.A(new_n12871_), .B(new_n12879_), .Y(new_n13033_));
  AOI21X1  g12031(.A0(new_n12867_), .A1(new_n12329_), .B0(new_n13033_), .Y(new_n13034_));
  AOI22X1  g12032(.A0(new_n13034_), .A1(new_n12870_), .B0(new_n12877_), .B1(new_n12876_), .Y(new_n13035_));
  AOI21X1  g12033(.A0(new_n12871_), .A1(new_n12870_), .B0(new_n12868_), .Y(new_n13036_));
  OR2X1    g12034(.A(new_n13036_), .B(new_n13035_), .Y(new_n13037_));
  XOR2X1   g12035(.A(new_n13037_), .B(new_n13032_), .Y(new_n13038_));
  OAI21X1  g12036(.A0(new_n13025_), .A1(new_n13022_), .B0(new_n13038_), .Y(new_n13039_));
  AOI22X1  g12037(.A0(new_n12838_), .A1(new_n12347_), .B0(new_n12753_), .B1(new_n12752_), .Y(new_n13040_));
  NOR2X1   g12038(.A(new_n12838_), .B(new_n12347_), .Y(new_n13041_));
  AND2X1   g12039(.A(new_n12861_), .B(new_n12853_), .Y(new_n13042_));
  OAI22X1  g12040(.A0(new_n12884_), .A1(new_n13042_), .B0(new_n13041_), .B1(new_n13040_), .Y(new_n13043_));
  NAND4X1  g12041(.A(new_n12883_), .B(new_n12874_), .C(new_n12861_), .D(new_n12853_), .Y(new_n13044_));
  NOR2X1   g12042(.A(new_n13036_), .B(new_n13035_), .Y(new_n13045_));
  NAND2X1  g12043(.A(new_n13045_), .B(new_n13032_), .Y(new_n13046_));
  OR2X1    g12044(.A(new_n13045_), .B(new_n13032_), .Y(new_n13047_));
  NAND4X1  g12045(.A(new_n13047_), .B(new_n13046_), .C(new_n13044_), .D(new_n13043_), .Y(new_n13048_));
  NAND2X1  g12046(.A(new_n13048_), .B(new_n13039_), .Y(new_n13049_));
  AOI22X1  g12047(.A0(new_n12823_), .A1(new_n12816_), .B0(new_n12798_), .B1(new_n12792_), .Y(new_n13050_));
  AOI21X1  g12048(.A0(new_n13015_), .A1(new_n13014_), .B0(new_n13050_), .Y(new_n13051_));
  AOI22X1  g12049(.A0(new_n12822_), .A1(new_n12821_), .B0(new_n12819_), .B1(new_n12818_), .Y(new_n13052_));
  NAND3X1  g12050(.A(new_n12823_), .B(new_n12798_), .C(new_n12792_), .Y(new_n13053_));
  NOR2X1   g12051(.A(new_n13053_), .B(new_n13052_), .Y(new_n13054_));
  NAND4X1  g12052(.A(new_n12519_), .B(new_n12513_), .C(new_n12497_), .D(new_n12489_), .Y(new_n13055_));
  AND2X1   g12053(.A(new_n12789_), .B(new_n12785_), .Y(new_n13056_));
  AND2X1   g12054(.A(new_n13056_), .B(new_n12784_), .Y(new_n13057_));
  AOI22X1  g12055(.A0(new_n13057_), .A1(new_n12788_), .B0(new_n13055_), .B1(new_n12794_), .Y(new_n13058_));
  AOI22X1  g12056(.A0(new_n12789_), .A1(new_n12788_), .B0(new_n12785_), .B1(new_n12784_), .Y(new_n13059_));
  NOR2X1   g12057(.A(new_n13059_), .B(new_n13058_), .Y(new_n13060_));
  NAND2X1  g12058(.A(new_n12813_), .B(new_n12422_), .Y(new_n13061_));
  OAI22X1  g12059(.A0(new_n12429_), .A1(new_n12428_), .B0(new_n12425_), .B1(new_n12424_), .Y(new_n13062_));
  AND2X1   g12060(.A(new_n13062_), .B(new_n12811_), .Y(new_n13063_));
  AND2X1   g12061(.A(new_n13063_), .B(new_n12810_), .Y(new_n13064_));
  AOI22X1  g12062(.A0(new_n13064_), .A1(new_n13061_), .B0(new_n12819_), .B1(new_n12818_), .Y(new_n13065_));
  AOI21X1  g12063(.A0(new_n12811_), .A1(new_n12810_), .B0(new_n12814_), .Y(new_n13066_));
  OR2X1    g12064(.A(new_n13066_), .B(new_n13065_), .Y(new_n13067_));
  NOR2X1   g12065(.A(new_n13067_), .B(new_n13060_), .Y(new_n13068_));
  AND2X1   g12066(.A(new_n13067_), .B(new_n13060_), .Y(new_n13069_));
  OAI22X1  g12067(.A0(new_n13069_), .A1(new_n13068_), .B0(new_n13054_), .B1(new_n13051_), .Y(new_n13070_));
  AND2X1   g12068(.A(new_n12798_), .B(new_n12792_), .Y(new_n13071_));
  OAI22X1  g12069(.A0(new_n12824_), .A1(new_n13071_), .B0(new_n12774_), .B1(new_n12773_), .Y(new_n13072_));
  NAND4X1  g12070(.A(new_n12823_), .B(new_n12816_), .C(new_n12798_), .D(new_n12792_), .Y(new_n13073_));
  OR2X1    g12071(.A(new_n13067_), .B(new_n13060_), .Y(new_n13074_));
  NAND2X1  g12072(.A(new_n13067_), .B(new_n13060_), .Y(new_n13075_));
  NAND4X1  g12073(.A(new_n13075_), .B(new_n13074_), .C(new_n13073_), .D(new_n13072_), .Y(new_n13076_));
  AND2X1   g12074(.A(new_n13076_), .B(new_n13070_), .Y(new_n13077_));
  XOR2X1   g12075(.A(new_n13077_), .B(new_n13049_), .Y(new_n13078_));
  XOR2X1   g12076(.A(new_n13078_), .B(new_n13020_), .Y(new_n13079_));
  OR2X1    g12077(.A(new_n13079_), .B(new_n13007_), .Y(new_n13080_));
  OAI21X1  g12078(.A0(new_n13006_), .A1(new_n12911_), .B0(new_n13079_), .Y(new_n13081_));
  AOI21X1  g12079(.A0(new_n13006_), .A1(new_n12911_), .B0(new_n13081_), .Y(new_n13082_));
  AOI21X1  g12080(.A0(new_n13080_), .A1(new_n12891_), .B0(new_n13082_), .Y(new_n13083_));
  OAI22X1  g12081(.A0(new_n11980_), .A1(new_n12678_), .B0(new_n11820_), .B1(new_n11816_), .Y(new_n13084_));
  OR2X1    g12082(.A(new_n12679_), .B(new_n11926_), .Y(new_n13085_));
  AOI21X1  g12083(.A0(new_n12719_), .A1(new_n12718_), .B0(new_n12912_), .Y(new_n13086_));
  AOI21X1  g12084(.A0(new_n13085_), .A1(new_n13084_), .B0(new_n13086_), .Y(new_n13087_));
  AND2X1   g12085(.A(new_n12912_), .B(new_n12718_), .Y(new_n13088_));
  AND2X1   g12086(.A(new_n13088_), .B(new_n12719_), .Y(new_n13089_));
  OR2X1    g12087(.A(new_n13089_), .B(new_n13087_), .Y(new_n13090_));
  XOR2X1   g12088(.A(new_n12940_), .B(new_n13090_), .Y(new_n13091_));
  NOR2X1   g12089(.A(new_n13005_), .B(new_n13091_), .Y(new_n13092_));
  NAND2X1  g12090(.A(new_n13005_), .B(new_n13091_), .Y(new_n13093_));
  OAI21X1  g12091(.A0(new_n13092_), .A1(new_n12911_), .B0(new_n13093_), .Y(new_n13094_));
  AOI21X1  g12092(.A0(new_n12938_), .A1(new_n12937_), .B0(new_n12936_), .Y(new_n13095_));
  NOR3X1   g12093(.A(new_n12934_), .B(new_n12927_), .C(new_n12919_), .Y(new_n13096_));
  AOI21X1  g12094(.A0(new_n12914_), .A1(new_n12913_), .B0(new_n13096_), .Y(new_n13097_));
  AOI21X1  g12095(.A0(new_n12922_), .A1(new_n12921_), .B0(new_n12933_), .Y(new_n13098_));
  OAI21X1  g12096(.A0(new_n13097_), .A1(new_n13095_), .B0(new_n13098_), .Y(new_n13099_));
  OR2X1    g12097(.A(new_n13098_), .B(new_n13095_), .Y(new_n13100_));
  OR2X1    g12098(.A(new_n13100_), .B(new_n13097_), .Y(new_n13101_));
  AOI22X1  g12099(.A0(new_n13002_), .A1(new_n12996_), .B0(new_n12976_), .B1(new_n12968_), .Y(new_n13102_));
  AOI21X1  g12100(.A0(new_n12949_), .A1(new_n12948_), .B0(new_n13102_), .Y(new_n13103_));
  AOI22X1  g12101(.A0(new_n12975_), .A1(new_n12974_), .B0(new_n12973_), .B1(new_n12972_), .Y(new_n13104_));
  NOR4X1   g12102(.A(new_n12967_), .B(new_n12966_), .C(new_n12955_), .D(new_n12952_), .Y(new_n13105_));
  AOI22X1  g12103(.A0(new_n13001_), .A1(new_n13000_), .B0(new_n12999_), .B1(new_n12998_), .Y(new_n13106_));
  NOR4X1   g12104(.A(new_n12995_), .B(new_n12994_), .C(new_n12982_), .D(new_n12979_), .Y(new_n13107_));
  NOR4X1   g12105(.A(new_n13107_), .B(new_n13106_), .C(new_n13105_), .D(new_n13104_), .Y(new_n13108_));
  OR4X1    g12106(.A(new_n12992_), .B(new_n12991_), .C(new_n12987_), .D(new_n12986_), .Y(new_n13109_));
  OAI21X1  g12107(.A0(new_n12982_), .A1(new_n12979_), .B0(new_n13109_), .Y(new_n13110_));
  OAI22X1  g12108(.A0(new_n12992_), .A1(new_n12991_), .B0(new_n12987_), .B1(new_n12986_), .Y(new_n13111_));
  NAND2X1  g12109(.A(new_n13111_), .B(new_n13110_), .Y(new_n13112_));
  INVX1    g12110(.A(new_n12964_), .Y(new_n13113_));
  OAI22X1  g12111(.A0(new_n12652_), .A1(new_n12649_), .B0(new_n12631_), .B1(new_n12627_), .Y(new_n13114_));
  OR2X1    g12112(.A(new_n13114_), .B(new_n12959_), .Y(new_n13115_));
  OAI22X1  g12113(.A0(new_n13115_), .A1(new_n13113_), .B0(new_n12955_), .B1(new_n12952_), .Y(new_n13116_));
  OAI21X1  g12114(.A0(new_n12960_), .A1(new_n12959_), .B0(new_n12965_), .Y(new_n13117_));
  AND2X1   g12115(.A(new_n13117_), .B(new_n13116_), .Y(new_n13118_));
  AND2X1   g12116(.A(new_n13118_), .B(new_n13112_), .Y(new_n13119_));
  NOR2X1   g12117(.A(new_n13118_), .B(new_n13112_), .Y(new_n13120_));
  OAI22X1  g12118(.A0(new_n13120_), .A1(new_n13119_), .B0(new_n13108_), .B1(new_n13103_), .Y(new_n13121_));
  OR2X1    g12119(.A(new_n12970_), .B(new_n12969_), .Y(new_n13122_));
  XOR2X1   g12120(.A(new_n12663_), .B(new_n13122_), .Y(new_n13123_));
  AOI22X1  g12121(.A0(new_n13123_), .A1(new_n12603_), .B0(new_n12906_), .B1(new_n12905_), .Y(new_n13124_));
  AND2X1   g12122(.A(new_n12664_), .B(new_n12947_), .Y(new_n13125_));
  OAI22X1  g12123(.A0(new_n13107_), .A1(new_n13106_), .B0(new_n13105_), .B1(new_n13104_), .Y(new_n13126_));
  OAI21X1  g12124(.A0(new_n13125_), .A1(new_n13124_), .B0(new_n13126_), .Y(new_n13127_));
  NAND4X1  g12125(.A(new_n13002_), .B(new_n12996_), .C(new_n12976_), .D(new_n12968_), .Y(new_n13128_));
  NAND2X1  g12126(.A(new_n13118_), .B(new_n13112_), .Y(new_n13129_));
  OR2X1    g12127(.A(new_n13118_), .B(new_n13112_), .Y(new_n13130_));
  NAND4X1  g12128(.A(new_n13130_), .B(new_n13129_), .C(new_n13128_), .D(new_n13127_), .Y(new_n13131_));
  AOI22X1  g12129(.A0(new_n13131_), .A1(new_n13121_), .B0(new_n13101_), .B1(new_n13099_), .Y(new_n13132_));
  OAI21X1  g12130(.A0(new_n13089_), .A1(new_n13087_), .B0(new_n12939_), .Y(new_n13133_));
  INVX1    g12131(.A(new_n13098_), .Y(new_n13134_));
  AOI21X1  g12132(.A0(new_n13133_), .A1(new_n12935_), .B0(new_n13134_), .Y(new_n13135_));
  NOR2X1   g12133(.A(new_n13100_), .B(new_n13097_), .Y(new_n13136_));
  AOI22X1  g12134(.A0(new_n13130_), .A1(new_n13129_), .B0(new_n13128_), .B1(new_n13127_), .Y(new_n13137_));
  NOR4X1   g12135(.A(new_n13120_), .B(new_n13119_), .C(new_n13108_), .D(new_n13103_), .Y(new_n13138_));
  NOR4X1   g12136(.A(new_n13138_), .B(new_n13137_), .C(new_n13136_), .D(new_n13135_), .Y(new_n13139_));
  NOR2X1   g12137(.A(new_n13139_), .B(new_n13132_), .Y(new_n13140_));
  XOR2X1   g12138(.A(new_n13140_), .B(new_n13094_), .Y(new_n13141_));
  OR2X1    g12139(.A(new_n13041_), .B(new_n13040_), .Y(new_n13142_));
  XOR2X1   g12140(.A(new_n12885_), .B(new_n13142_), .Y(new_n13143_));
  AOI22X1  g12141(.A0(new_n13143_), .A1(new_n12826_), .B0(new_n12765_), .B1(new_n12756_), .Y(new_n13144_));
  AND2X1   g12142(.A(new_n12886_), .B(new_n13017_), .Y(new_n13145_));
  AND2X1   g12143(.A(new_n13048_), .B(new_n13039_), .Y(new_n13146_));
  OAI22X1  g12144(.A0(new_n13077_), .A1(new_n13146_), .B0(new_n13145_), .B1(new_n13144_), .Y(new_n13147_));
  NAND4X1  g12145(.A(new_n13076_), .B(new_n13070_), .C(new_n13048_), .D(new_n13039_), .Y(new_n13148_));
  OR4X1    g12146(.A(new_n13066_), .B(new_n13065_), .C(new_n13059_), .D(new_n13058_), .Y(new_n13149_));
  OAI21X1  g12147(.A0(new_n13054_), .A1(new_n13051_), .B0(new_n13149_), .Y(new_n13150_));
  OAI22X1  g12148(.A0(new_n13066_), .A1(new_n13065_), .B0(new_n13059_), .B1(new_n13058_), .Y(new_n13151_));
  NAND2X1  g12149(.A(new_n13151_), .B(new_n13150_), .Y(new_n13152_));
  NOR4X1   g12150(.A(new_n13036_), .B(new_n13035_), .C(new_n13031_), .D(new_n13030_), .Y(new_n13153_));
  AOI21X1  g12151(.A0(new_n13044_), .A1(new_n13043_), .B0(new_n13153_), .Y(new_n13154_));
  AND2X1   g12152(.A(new_n13037_), .B(new_n13032_), .Y(new_n13155_));
  NOR2X1   g12153(.A(new_n13155_), .B(new_n13154_), .Y(new_n13156_));
  XOR2X1   g12154(.A(new_n13156_), .B(new_n13152_), .Y(new_n13157_));
  AOI21X1  g12155(.A0(new_n13148_), .A1(new_n13147_), .B0(new_n13157_), .Y(new_n13158_));
  AOI22X1  g12156(.A0(new_n13076_), .A1(new_n13070_), .B0(new_n13048_), .B1(new_n13039_), .Y(new_n13159_));
  AOI21X1  g12157(.A0(new_n13019_), .A1(new_n13018_), .B0(new_n13159_), .Y(new_n13160_));
  AOI22X1  g12158(.A0(new_n13075_), .A1(new_n13074_), .B0(new_n13073_), .B1(new_n13072_), .Y(new_n13161_));
  NAND3X1  g12159(.A(new_n13076_), .B(new_n13048_), .C(new_n13039_), .Y(new_n13162_));
  NOR2X1   g12160(.A(new_n13162_), .B(new_n13161_), .Y(new_n13163_));
  AND2X1   g12161(.A(new_n13156_), .B(new_n13152_), .Y(new_n13164_));
  NOR2X1   g12162(.A(new_n13156_), .B(new_n13152_), .Y(new_n13165_));
  NOR4X1   g12163(.A(new_n13165_), .B(new_n13164_), .C(new_n13163_), .D(new_n13160_), .Y(new_n13166_));
  NOR2X1   g12164(.A(new_n13166_), .B(new_n13158_), .Y(new_n13167_));
  NOR2X1   g12165(.A(new_n13167_), .B(new_n13141_), .Y(new_n13168_));
  OR2X1    g12166(.A(new_n13168_), .B(new_n13083_), .Y(new_n13169_));
  AND2X1   g12167(.A(new_n13140_), .B(new_n13094_), .Y(new_n13170_));
  NOR2X1   g12168(.A(new_n13140_), .B(new_n13094_), .Y(new_n13171_));
  OR4X1    g12169(.A(new_n13166_), .B(new_n13158_), .C(new_n13171_), .D(new_n13170_), .Y(new_n13172_));
  NOR2X1   g12170(.A(new_n12748_), .B(new_n12908_), .Y(new_n13173_));
  NAND2X1  g12171(.A(new_n12748_), .B(new_n12908_), .Y(new_n13174_));
  OAI21X1  g12172(.A0(new_n13173_), .A1(new_n12532_), .B0(new_n13174_), .Y(new_n13175_));
  OR2X1    g12173(.A(new_n13005_), .B(new_n13091_), .Y(new_n13176_));
  AND2X1   g12174(.A(new_n13005_), .B(new_n13091_), .Y(new_n13177_));
  AOI21X1  g12175(.A0(new_n13176_), .A1(new_n13175_), .B0(new_n13177_), .Y(new_n13178_));
  OR4X1    g12176(.A(new_n13138_), .B(new_n13137_), .C(new_n13136_), .D(new_n13135_), .Y(new_n13179_));
  OAI21X1  g12177(.A0(new_n13132_), .A1(new_n13178_), .B0(new_n13179_), .Y(new_n13180_));
  AND2X1   g12178(.A(new_n13117_), .B(new_n13111_), .Y(new_n13181_));
  NAND3X1  g12179(.A(new_n13181_), .B(new_n13116_), .C(new_n13110_), .Y(new_n13182_));
  OAI21X1  g12180(.A0(new_n13108_), .A1(new_n13103_), .B0(new_n13182_), .Y(new_n13183_));
  AOI22X1  g12181(.A0(new_n13117_), .A1(new_n13116_), .B0(new_n13111_), .B1(new_n13110_), .Y(new_n13184_));
  INVX1    g12182(.A(new_n13184_), .Y(new_n13185_));
  NAND3X1  g12183(.A(new_n13185_), .B(new_n13183_), .C(new_n13099_), .Y(new_n13186_));
  AND2X1   g12184(.A(new_n13181_), .B(new_n13110_), .Y(new_n13187_));
  AOI22X1  g12185(.A0(new_n13187_), .A1(new_n13116_), .B0(new_n13128_), .B1(new_n13127_), .Y(new_n13188_));
  OAI21X1  g12186(.A0(new_n13184_), .A1(new_n13188_), .B0(new_n13135_), .Y(new_n13189_));
  AND2X1   g12187(.A(new_n13189_), .B(new_n13186_), .Y(new_n13190_));
  NAND2X1  g12188(.A(new_n13190_), .B(new_n13180_), .Y(new_n13191_));
  AOI21X1  g12189(.A0(new_n13189_), .A1(new_n13186_), .B0(new_n13139_), .Y(new_n13192_));
  OAI21X1  g12190(.A0(new_n13132_), .A1(new_n13178_), .B0(new_n13192_), .Y(new_n13193_));
  INVX1    g12191(.A(new_n13155_), .Y(new_n13194_));
  NAND3X1  g12192(.A(new_n13194_), .B(new_n13151_), .C(new_n13150_), .Y(new_n13195_));
  OAI22X1  g12193(.A0(new_n13195_), .A1(new_n13154_), .B0(new_n13163_), .B1(new_n13160_), .Y(new_n13196_));
  OAI21X1  g12194(.A0(new_n13155_), .A1(new_n13154_), .B0(new_n13152_), .Y(new_n13197_));
  AND2X1   g12195(.A(new_n13197_), .B(new_n13196_), .Y(new_n13198_));
  INVX1    g12196(.A(new_n13198_), .Y(new_n13199_));
  AOI21X1  g12197(.A0(new_n13193_), .A1(new_n13191_), .B0(new_n13199_), .Y(new_n13200_));
  AOI21X1  g12198(.A0(new_n13172_), .A1(new_n13169_), .B0(new_n13200_), .Y(new_n13201_));
  AND2X1   g12199(.A(new_n13190_), .B(new_n13180_), .Y(new_n13202_));
  OR2X1    g12200(.A(new_n13132_), .B(new_n13178_), .Y(new_n13203_));
  AND2X1   g12201(.A(new_n13192_), .B(new_n13203_), .Y(new_n13204_));
  NOR3X1   g12202(.A(new_n13198_), .B(new_n13204_), .C(new_n13202_), .Y(new_n13205_));
  INVX1    g12203(.A(new_n13189_), .Y(new_n13206_));
  AOI21X1  g12204(.A0(new_n13186_), .A1(new_n13180_), .B0(new_n13206_), .Y(new_n13207_));
  OAI21X1  g12205(.A0(new_n13205_), .A1(new_n13201_), .B0(new_n13207_), .Y(new_n13208_));
  OR2X1    g12206(.A(new_n13207_), .B(new_n13205_), .Y(new_n13209_));
  OR2X1    g12207(.A(new_n13209_), .B(new_n13201_), .Y(new_n13210_));
  AND2X1   g12208(.A(new_n13210_), .B(new_n13208_), .Y(new_n13211_));
  NOR3X1   g12209(.A(new_n8838_), .B(new_n8837_), .C(new_n8833_), .Y(new_n13212_));
  AOI21X1  g12210(.A0(new_n8823_), .A1(new_n8810_), .B0(new_n8829_), .Y(new_n13213_));
  OAI21X1  g12211(.A0(new_n13213_), .A1(new_n13212_), .B0(new_n8841_), .Y(new_n13214_));
  OAI21X1  g12212(.A0(new_n10548_), .A1(new_n8851_), .B0(new_n5642_), .Y(new_n13215_));
  INVX1    g12213(.A(new_n8847_), .Y(new_n13216_));
  NAND3X1  g12214(.A(new_n13216_), .B(new_n13215_), .C(new_n13214_), .Y(new_n13217_));
  AOI21X1  g12215(.A0(new_n13215_), .A1(new_n13214_), .B0(new_n13216_), .Y(new_n13218_));
  AOI21X1  g12216(.A0(new_n13217_), .A1(new_n3848_), .B0(new_n13218_), .Y(new_n13219_));
  OR2X1    g12217(.A(new_n10546_), .B(new_n8852_), .Y(new_n13220_));
  AOI21X1  g12218(.A0(new_n10546_), .A1(new_n8852_), .B0(new_n10551_), .Y(new_n13221_));
  AOI22X1  g12219(.A0(new_n13221_), .A1(new_n13220_), .B0(new_n10551_), .B1(new_n10007_), .Y(new_n13222_));
  INVX1    g12220(.A(new_n8845_), .Y(new_n13223_));
  AOI21X1  g12221(.A0(new_n8828_), .A1(new_n8824_), .B0(new_n8845_), .Y(new_n13224_));
  OAI21X1  g12222(.A0(new_n8828_), .A1(new_n8824_), .B0(new_n13224_), .Y(new_n13225_));
  OAI21X1  g12223(.A0(new_n8846_), .A1(new_n13223_), .B0(new_n13225_), .Y(new_n13226_));
  AND2X1   g12224(.A(new_n13226_), .B(\A[1000] ), .Y(new_n13227_));
  OAI21X1  g12225(.A0(new_n13222_), .A1(new_n13219_), .B0(new_n13227_), .Y(new_n13228_));
  XOR2X1   g12226(.A(new_n10546_), .B(new_n8852_), .Y(new_n13229_));
  OAI21X1  g12227(.A0(new_n10006_), .A1(new_n10549_), .B0(new_n10539_), .Y(new_n13230_));
  OAI22X1  g12228(.A0(new_n13230_), .A1(new_n10547_), .B0(new_n10539_), .B1(new_n13229_), .Y(new_n13231_));
  NAND3X1  g12229(.A(new_n8847_), .B(new_n13215_), .C(new_n13214_), .Y(new_n13232_));
  OAI21X1  g12230(.A0(new_n8844_), .A1(new_n8840_), .B0(new_n13216_), .Y(new_n13233_));
  AOI21X1  g12231(.A0(new_n13233_), .A1(new_n13232_), .B0(new_n3848_), .Y(new_n13234_));
  AOI21X1  g12232(.A0(new_n8849_), .A1(new_n13217_), .B0(new_n3849_), .Y(new_n13235_));
  OAI22X1  g12233(.A0(new_n13235_), .A1(new_n13234_), .B0(new_n13231_), .B1(new_n8850_), .Y(new_n13236_));
  NOR2X1   g12234(.A(new_n13236_), .B(new_n13228_), .Y(new_n13237_));
  AND2X1   g12235(.A(new_n10539_), .B(new_n10007_), .Y(new_n13238_));
  OAI22X1  g12236(.A0(new_n10552_), .A1(new_n10547_), .B0(new_n13238_), .B1(new_n13219_), .Y(new_n13239_));
  XOR2X1   g12237(.A(new_n11338_), .B(new_n10557_), .Y(new_n13240_));
  OAI21X1  g12238(.A0(new_n11338_), .A1(new_n10557_), .B0(new_n11782_), .Y(new_n13241_));
  OAI22X1  g12239(.A0(new_n13241_), .A1(new_n11339_), .B0(new_n11782_), .B1(new_n13240_), .Y(new_n13242_));
  XOR2X1   g12240(.A(new_n13242_), .B(new_n13239_), .Y(new_n13243_));
  AND2X1   g12241(.A(new_n13243_), .B(new_n13237_), .Y(new_n13244_));
  NAND2X1  g12242(.A(new_n11782_), .B(new_n11343_), .Y(new_n13245_));
  NOR2X1   g12243(.A(new_n11792_), .B(new_n11339_), .Y(new_n13246_));
  AOI21X1  g12244(.A0(new_n13245_), .A1(new_n13239_), .B0(new_n13246_), .Y(new_n13247_));
  AND2X1   g12245(.A(new_n13009_), .B(new_n13008_), .Y(new_n13248_));
  XOR2X1   g12246(.A(new_n12525_), .B(new_n13248_), .Y(new_n13249_));
  AOI21X1  g12247(.A0(new_n12269_), .A1(new_n11806_), .B0(new_n13249_), .Y(new_n13250_));
  AOI22X1  g12248(.A0(new_n13250_), .A1(new_n12270_), .B0(new_n13249_), .B1(new_n12274_), .Y(new_n13251_));
  XOR2X1   g12249(.A(new_n13251_), .B(new_n13247_), .Y(new_n13252_));
  AND2X1   g12250(.A(new_n13252_), .B(new_n13244_), .Y(new_n13253_));
  NAND2X1  g12251(.A(new_n12749_), .B(new_n12532_), .Y(new_n13254_));
  XOR2X1   g12252(.A(new_n12749_), .B(new_n12894_), .Y(new_n13255_));
  XOR2X1   g12253(.A(new_n12748_), .B(new_n12908_), .Y(new_n13256_));
  AOI21X1  g12254(.A0(new_n13256_), .A1(new_n12894_), .B0(new_n12888_), .Y(new_n13257_));
  AOI22X1  g12255(.A0(new_n13257_), .A1(new_n13254_), .B0(new_n12888_), .B1(new_n13255_), .Y(new_n13258_));
  XOR2X1   g12256(.A(new_n13258_), .B(new_n12529_), .Y(new_n13259_));
  NAND2X1  g12257(.A(new_n13259_), .B(new_n13253_), .Y(new_n13260_));
  NAND2X1  g12258(.A(new_n13006_), .B(new_n12911_), .Y(new_n13261_));
  XOR2X1   g12259(.A(new_n13006_), .B(new_n13175_), .Y(new_n13262_));
  XOR2X1   g12260(.A(new_n13005_), .B(new_n13091_), .Y(new_n13263_));
  AOI21X1  g12261(.A0(new_n13263_), .A1(new_n13175_), .B0(new_n13079_), .Y(new_n13264_));
  AOI22X1  g12262(.A0(new_n13264_), .A1(new_n13261_), .B0(new_n13079_), .B1(new_n13262_), .Y(new_n13265_));
  XOR2X1   g12263(.A(new_n13265_), .B(new_n12891_), .Y(new_n13266_));
  OR2X1    g12264(.A(new_n13266_), .B(new_n13260_), .Y(new_n13267_));
  OR2X1    g12265(.A(new_n13140_), .B(new_n13094_), .Y(new_n13268_));
  XOR2X1   g12266(.A(new_n13140_), .B(new_n13178_), .Y(new_n13269_));
  AOI21X1  g12267(.A0(new_n13140_), .A1(new_n13094_), .B0(new_n13167_), .Y(new_n13270_));
  AOI22X1  g12268(.A0(new_n13270_), .A1(new_n13268_), .B0(new_n13167_), .B1(new_n13269_), .Y(new_n13271_));
  XOR2X1   g12269(.A(new_n13271_), .B(new_n13083_), .Y(new_n13272_));
  INVX1    g12270(.A(new_n13272_), .Y(new_n13273_));
  NOR2X1   g12271(.A(new_n13168_), .B(new_n13083_), .Y(new_n13274_));
  NOR4X1   g12272(.A(new_n13166_), .B(new_n13158_), .C(new_n13171_), .D(new_n13170_), .Y(new_n13275_));
  AOI21X1  g12273(.A0(new_n13193_), .A1(new_n13191_), .B0(new_n13198_), .Y(new_n13276_));
  NOR3X1   g12274(.A(new_n13199_), .B(new_n13204_), .C(new_n13202_), .Y(new_n13277_));
  NOR4X1   g12275(.A(new_n13277_), .B(new_n13276_), .C(new_n13275_), .D(new_n13274_), .Y(new_n13278_));
  OAI21X1  g12276(.A0(new_n13204_), .A1(new_n13202_), .B0(new_n13199_), .Y(new_n13279_));
  NAND3X1  g12277(.A(new_n13198_), .B(new_n13193_), .C(new_n13191_), .Y(new_n13280_));
  AOI22X1  g12278(.A0(new_n13280_), .A1(new_n13279_), .B0(new_n13172_), .B1(new_n13169_), .Y(new_n13281_));
  NOR4X1   g12279(.A(new_n13281_), .B(new_n13278_), .C(new_n13273_), .D(new_n13267_), .Y(new_n13282_));
  AND2X1   g12280(.A(new_n13259_), .B(new_n13253_), .Y(new_n13283_));
  XOR2X1   g12281(.A(new_n13222_), .B(new_n13219_), .Y(new_n13284_));
  INVX1    g12282(.A(new_n13227_), .Y(new_n13285_));
  NOR3X1   g12283(.A(new_n13216_), .B(new_n8844_), .C(new_n8840_), .Y(new_n13286_));
  AOI21X1  g12284(.A0(new_n13215_), .A1(new_n13214_), .B0(new_n8847_), .Y(new_n13287_));
  OAI21X1  g12285(.A0(new_n13287_), .A1(new_n13286_), .B0(new_n3849_), .Y(new_n13288_));
  OAI21X1  g12286(.A0(new_n13218_), .A1(new_n8848_), .B0(new_n3848_), .Y(new_n13289_));
  AOI21X1  g12287(.A0(new_n13289_), .A1(new_n13288_), .B0(new_n13285_), .Y(new_n13290_));
  OAI22X1  g12288(.A0(new_n13290_), .A1(new_n13284_), .B0(new_n13236_), .B1(new_n13228_), .Y(new_n13291_));
  NAND3X1  g12289(.A(new_n13289_), .B(new_n13288_), .C(new_n13227_), .Y(new_n13292_));
  OAI21X1  g12290(.A0(new_n13235_), .A1(new_n13234_), .B0(new_n13285_), .Y(new_n13293_));
  NAND3X1  g12291(.A(new_n13293_), .B(new_n13292_), .C(new_n13291_), .Y(new_n13294_));
  XOR2X1   g12292(.A(new_n13243_), .B(new_n13237_), .Y(new_n13295_));
  NAND2X1  g12293(.A(new_n13295_), .B(new_n13294_), .Y(new_n13296_));
  XOR2X1   g12294(.A(new_n13251_), .B(new_n11793_), .Y(new_n13297_));
  XOR2X1   g12295(.A(new_n13297_), .B(new_n13244_), .Y(new_n13298_));
  AND2X1   g12296(.A(new_n13298_), .B(new_n13296_), .Y(new_n13299_));
  NOR2X1   g12297(.A(new_n13259_), .B(new_n13253_), .Y(new_n13300_));
  OR4X1    g12298(.A(new_n13300_), .B(new_n13299_), .C(new_n13266_), .D(new_n13283_), .Y(new_n13301_));
  XOR2X1   g12299(.A(new_n13272_), .B(new_n13267_), .Y(new_n13302_));
  OR2X1    g12300(.A(new_n13302_), .B(new_n13301_), .Y(new_n13303_));
  NOR2X1   g12301(.A(new_n13266_), .B(new_n13260_), .Y(new_n13304_));
  AND2X1   g12302(.A(new_n13272_), .B(new_n13304_), .Y(new_n13305_));
  NOR2X1   g12303(.A(new_n13281_), .B(new_n13278_), .Y(new_n13306_));
  NOR2X1   g12304(.A(new_n13306_), .B(new_n13305_), .Y(new_n13307_));
  NOR4X1   g12305(.A(new_n13307_), .B(new_n13303_), .C(new_n13282_), .D(new_n13211_), .Y(new_n13308_));
  NOR2X1   g12306(.A(new_n13205_), .B(new_n13201_), .Y(new_n13309_));
  OR2X1    g12307(.A(new_n13281_), .B(new_n13278_), .Y(new_n13310_));
  NOR4X1   g12308(.A(new_n13310_), .B(new_n13273_), .C(new_n13267_), .D(new_n13211_), .Y(new_n13311_));
  NOR3X1   g12309(.A(new_n13311_), .B(new_n13207_), .C(new_n13309_), .Y(new_n13312_));
  OAI21X1  g12310(.A0(new_n13207_), .A1(new_n13309_), .B0(new_n13282_), .Y(new_n13313_));
  NOR2X1   g12311(.A(new_n13313_), .B(new_n13211_), .Y(new_n13314_));
  OR4X1    g12312(.A(new_n13278_), .B(new_n13273_), .C(new_n13267_), .D(new_n13207_), .Y(new_n13315_));
  NOR4X1   g12313(.A(new_n13315_), .B(new_n13281_), .C(new_n13211_), .D(new_n13309_), .Y(new_n13316_));
  NOR4X1   g12314(.A(new_n13316_), .B(new_n13314_), .C(new_n13312_), .D(new_n13308_), .Y(new_n13317_));
  XOR2X1   g12315(.A(new_n13282_), .B(new_n13211_), .Y(new_n13318_));
  XOR2X1   g12316(.A(new_n13306_), .B(new_n13305_), .Y(new_n13319_));
  XOR2X1   g12317(.A(new_n13302_), .B(new_n13301_), .Y(new_n13320_));
  NOR2X1   g12318(.A(new_n13290_), .B(new_n13284_), .Y(new_n13321_));
  NOR2X1   g12319(.A(new_n13321_), .B(new_n13237_), .Y(new_n13322_));
  NAND2X1  g12320(.A(new_n13293_), .B(new_n13292_), .Y(new_n13323_));
  INVX1    g12321(.A(new_n13226_), .Y(new_n13324_));
  AND2X1   g12322(.A(new_n13225_), .B(\A[1000] ), .Y(new_n13325_));
  OAI21X1  g12323(.A0(new_n8846_), .A1(new_n13223_), .B0(new_n13325_), .Y(new_n13326_));
  OAI21X1  g12324(.A0(new_n13324_), .A1(\A[1000] ), .B0(new_n13326_), .Y(new_n13327_));
  MX2X1    g12325(.A(new_n13327_), .B(new_n13322_), .S0(new_n13323_), .Y(new_n13328_));
  MX2X1    g12326(.A(new_n13295_), .B(new_n13328_), .S0(new_n13294_), .Y(new_n13329_));
  AND2X1   g12327(.A(new_n13329_), .B(new_n13296_), .Y(new_n13330_));
  NOR2X1   g12328(.A(new_n13298_), .B(new_n13296_), .Y(new_n13331_));
  NAND2X1  g12329(.A(new_n13252_), .B(new_n13244_), .Y(new_n13332_));
  XOR2X1   g12330(.A(new_n13259_), .B(new_n13332_), .Y(new_n13333_));
  XOR2X1   g12331(.A(new_n13333_), .B(new_n13299_), .Y(new_n13334_));
  NOR3X1   g12332(.A(new_n13334_), .B(new_n13331_), .C(new_n13330_), .Y(new_n13335_));
  OR4X1    g12333(.A(new_n13335_), .B(new_n13300_), .C(new_n13299_), .D(new_n13283_), .Y(new_n13337_));
  OR2X1    g12334(.A(new_n13333_), .B(new_n13299_), .Y(new_n13338_));
  XOR2X1   g12335(.A(new_n13266_), .B(new_n13260_), .Y(new_n13339_));
  AND2X1   g12336(.A(new_n13339_), .B(new_n13338_), .Y(new_n13340_));
  INVX1    g12337(.A(new_n13340_), .Y(new_n13341_));
  NAND2X1  g12338(.A(new_n13341_), .B(new_n13337_), .Y(new_n13342_));
  AND2X1   g12339(.A(new_n13342_), .B(new_n13320_), .Y(new_n13343_));
  NOR2X1   g12340(.A(new_n13272_), .B(new_n13304_), .Y(new_n13344_));
  NOR4X1   g12341(.A(new_n13344_), .B(new_n13301_), .C(new_n13310_), .D(new_n13305_), .Y(new_n13345_));
  NOR3X1   g12342(.A(new_n13335_), .B(new_n13333_), .C(new_n13299_), .Y(new_n13346_));
  NOR3X1   g12343(.A(new_n13340_), .B(new_n13346_), .C(new_n13320_), .Y(new_n13347_));
  OAI21X1  g12344(.A0(new_n13347_), .A1(new_n13302_), .B0(new_n13345_), .Y(new_n13348_));
  OAI21X1  g12345(.A0(new_n13348_), .A1(new_n13343_), .B0(new_n13319_), .Y(new_n13349_));
  NOR4X1   g12346(.A(new_n13307_), .B(new_n13303_), .C(new_n13282_), .D(new_n13211_), .Y(new_n13352_));
  AOI21X1  g12347(.A0(new_n13352_), .A1(new_n13349_), .B0(new_n13318_), .Y(new_n13353_));
  INVX1    g12348(.A(new_n13319_), .Y(new_n13354_));
  NOR4X1   g12349(.A(new_n13349_), .B(new_n13308_), .C(new_n13354_), .D(new_n13303_), .Y(new_n13355_));
  NOR3X1   g12350(.A(new_n13355_), .B(new_n13353_), .C(new_n13308_), .Y(new_n13356_));
  OAI21X1  g12351(.A0(new_n13313_), .A1(new_n13211_), .B0(new_n13345_), .Y(new_n13357_));
  NOR3X1   g12352(.A(new_n13357_), .B(new_n13312_), .C(new_n13318_), .Y(new_n13358_));
  OAI21X1  g12353(.A0(new_n13358_), .A1(new_n13356_), .B0(new_n13317_), .Y(maj));
endmodule


