//Converted to Combinational , Module name: b06 , Timestamp: 2018-11-27T15:20:53.240910 
module b06 ( EQL, CONT_EQL, STATE_REG_2_, STATE_REG_1_, STATE_REG_0_, CC_MUX_REG_2_, CC_MUX_REG_1_, USCITE_REG_2_, USCITE_REG_1_, ENABLE_COUNT_REG, ACKOUT_REG, n21, n26, n31 );
input EQL, CONT_EQL, STATE_REG_2_, STATE_REG_1_, STATE_REG_0_;
output CC_MUX_REG_2_, CC_MUX_REG_1_, USCITE_REG_2_, USCITE_REG_1_, ENABLE_COUNT_REG, ACKOUT_REG, n21, n26, n31;
wire n35, n36_1, n37, n38, n39, n40_1, n42, n43, n44_1, n45, n47, n48_1, n49, n50, n51_1, n53, n55, n57, n58, CC_MUX_REG_2__1, CC_MUX_REG_1__1, USCITE_REG_2__1, USCITE_REG_1__1, ENABLE_COUNT_REG_1;
INVX1    g00(.A(STATE_REG_0_), .Y(n35));
NAND2X1  g01(.A(STATE_REG_1_), .B(STATE_REG_2_), .Y(CC_MUX_REG_2__1));
NOR2X1   g02(.A(CC_MUX_REG_2__1), .B(n35), .Y(n37));
INVX1    g03(.A(EQL), .Y(n38));
INVX1    g04(.A(STATE_REG_2_), .Y(n39));
NAND4X1  g05(.A(STATE_REG_1_), .B(n39), .C(n38), .D(n35), .Y(CC_MUX_REG_1__1));
OAI21X1  g06(.A0(n37), .A1(CONT_EQL), .B0(CC_MUX_REG_1__1), .Y(ACKOUT_REG));
NOR2X1   g07(.A(STATE_REG_0_), .B(STATE_REG_1_), .Y(n42));
OAI21X1  g08(.A0(n42), .A1(EQL), .B0(STATE_REG_2_), .Y(n43));
INVX1    g09(.A(STATE_REG_1_), .Y(USCITE_REG_2__1));
NAND3X1  g10(.A(STATE_REG_0_), .B(USCITE_REG_2__1), .C(n39), .Y(n45));
OAI21X1  g11(.A0(n45), .A1(EQL), .B0(n43), .Y(n21));
NAND2X1  g12(.A(STATE_REG_1_), .B(EQL), .Y(n47));
NAND3X1  g13(.A(STATE_REG_0_), .B(n39), .C(EQL), .Y(USCITE_REG_1__1));
NAND4X1  g14(.A(USCITE_REG_2__1), .B(STATE_REG_2_), .C(n38), .D(n35), .Y(n49));
OR2X1    g15(.A(STATE_REG_0_), .B(STATE_REG_2_), .Y(n50));
OR2X1    g16(.A(n50), .B(USCITE_REG_2__1), .Y(ENABLE_COUNT_REG_1));
NAND4X1  g17(.A(n49), .B(USCITE_REG_1__1), .C(n47), .D(ENABLE_COUNT_REG_1), .Y(n26));
MX2X1    g18(.A(n35), .B(n50), .S0(USCITE_REG_2__1), .Y(n53));
OAI21X1  g19(.A0(n42), .A1(EQL), .B0(n53), .Y(n31));
OR2X1    g20(.A(n47), .B(STATE_REG_0_), .Y(n55));
NAND3X1  g21(.A(n55), .B(n45), .C(n43), .Y(CC_MUX_REG_2_));
OAI21X1  g22(.A0(STATE_REG_0_), .A1(n38), .B0(STATE_REG_1_), .Y(n57));
AOI22X1  g23(.A0(USCITE_REG_2__1), .A1(EQL), .B0(STATE_REG_2_), .B1(STATE_REG_0_), .Y(n58));
NAND3X1  g24(.A(n58), .B(n57), .C(n50), .Y(CC_MUX_REG_1_));
OAI21X1  g25(.A0(n47), .A1(n39), .B0(n49), .Y(USCITE_REG_2_));
NAND3X1  g26(.A(n53), .B(CC_MUX_REG_2__1), .C(EQL), .Y(USCITE_REG_1_));
OAI21X1  g27(.A0(n37), .A1(CONT_EQL), .B0(CC_MUX_REG_1__1), .Y(ENABLE_COUNT_REG));
endmodule
