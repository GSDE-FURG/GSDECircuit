//Converted to Combinational (Partial output: n7417) , Module name: s38584_n7417 , Timestamp: 2018-12-03T15:51:18.036961 
module s38584_n7417 ( g35, g2070, g2084, g1246, g1996, g1087, g1061, g979, g4180, g1211, g1205, g1216, g1221, g1171, g1183, g956, g2145, g2130, g2138, g947, g134, g209, g1193, g969, g1008, g691, n7417 );
input g35, g2070, g2084, g1246, g1996, g1087, g1061, g979, g4180, g1211, g1205, g1216, g1221, g1171, g1183, g956, g2145, g2130, g2138, g947, g134, g209, g1193, g969, g1008, g691;
output n7417;
wire n10785, n8497, n10784, n6085, n10782, n10783, n6081, n6084, n10781, n5528, n6080, n6082, n6083_1, n5524, n4664, n4665, n6079, n5246_1, n5752, n5269_1, n5519, n5245, n5518, n4709, n5517, n4707_1, n4708, n5516_1;
MX2X1    g6131(.A(g2070), .B(n10785), .S0(g35), .Y(n7417));
MX2X1    g6130(.A(g2084), .B(n10784), .S0(n8497), .Y(n10785));
INVX1    g3850(.A(n6085), .Y(n8497));
XOR2X1   g6129(.A(n10783), .B(n10782), .Y(n10784));
AND2X1   g1445(.A(n6084), .B(n6081), .Y(n6085));
MX2X1    g6127(.A(n10781), .B(g1246), .S0(n6084), .Y(n10782));
OAI21X1  g6128(.A0(g1996), .A1(g2070), .B0(g2084), .Y(n10783));
OAI21X1  g1441(.A0(n6080), .A1(n5528), .B0(g1087), .Y(n6081));
NOR2X1   g1444(.A(n6083_1), .B(n6082), .Y(n6084));
NOR2X1   g6126(.A(n6082), .B(n5524), .Y(n10781));
INVX1    g0888(.A(n4664), .Y(n5528));
NAND4X1  g1440(.A(g979), .B(n6079), .C(n4665), .D(g1061), .Y(n6080));
NAND2X1  g1442(.A(n5752), .B(n5246_1), .Y(n6082));
NOR2X1   g1443(.A(n5519), .B(n5269_1), .Y(n6083_1));
INVX1    g0884(.A(g4180), .Y(n5524));
NOR4X1   g0044(.A(g1221), .B(g1216), .C(g1205), .D(g1211), .Y(n4664));
INVX1    g0045(.A(g1171), .Y(n4665));
INVX1    g1439(.A(g1183), .Y(n6079));
NAND2X1  g0606(.A(n5245), .B(g956), .Y(n5246_1));
INVX1    g1112(.A(n5518), .Y(n5752));
INVX1    g0629(.A(g2145), .Y(n5269_1));
NAND2X1  g0879(.A(g2138), .B(g2130), .Y(n5519));
INVX1    g0605(.A(g947), .Y(n5245));
AOI21X1  g0878(.A0(n5517), .A1(n4709), .B0(g134), .Y(n5518));
NOR2X1   g0089(.A(n4708), .B(n4707_1), .Y(n4709));
NOR2X1   g0877(.A(n5516_1), .B(g209), .Y(n5517));
INVX1    g0087(.A(g1193), .Y(n4707_1));
NOR2X1   g0088(.A(g1008), .B(g969), .Y(n4708));
INVX1    g0876(.A(g691), .Y(n5516_1));

endmodule
