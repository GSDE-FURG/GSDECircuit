//Converted to Combinational (Partial output: n906) , Module name: s35932_n906 , Timestamp: 2018-12-03T15:51:08.497314 
module s35932_n906 ( RESET, TM1, TM0, WX499, WX723, WX851, WX2016, WX2144, WX659, WX787, WX1952, WX2080, WX853, WX855, WX857, WX859, WX861, WX863, WX865, WX867, WX869, WX837, WX871, WX839, WX873, WX841, WX875, WX843, WX877, WX845, WX879, WX847, WX881, WX849, WX883, WX885, WX887, WX889, WX891, WX893, WX895, WX897, WX899, n906 );
input RESET, TM1, TM0, WX499, WX723, WX851, WX2016, WX2144, WX659, WX787, WX1952, WX2080, WX853, WX855, WX857, WX859, WX861, WX863, WX865, WX867, WX869, WX837, WX871, WX839, WX873, WX841, WX875, WX843, WX877, WX845, WX879, WX847, WX881, WX849, WX883, WX885, WX887, WX889, WX891, WX893, WX895, WX897, WX899;
output n906;
wire n5827, n5923, n5922, n5920, n5539, n5600, n5921_1, n5918, n5913, n5597, n5599, n5915, n5917, CRC_OUT_9_24, n5596_1, n5598, n5914, n5916_1, n6360, CRC_OUT_9_23, n6358, CRC_OUT_9_22, n6356, CRC_OUT_9_21, n6354_1, CRC_OUT_9_20, n6352, CRC_OUT_9_19, n6350, CRC_OUT_9_18, n6348, CRC_OUT_9_17, n6346, CRC_OUT_9_16, n6344_1, CRC_OUT_9_15, n6343, n6341, CRC_OUT_9_31, CRC_OUT_9_14, n6374_1, n6339_1, CRC_OUT_9_30, CRC_OUT_9_13, n6372, n6337, CRC_OUT_9_29, CRC_OUT_9_12, n6370, n6335, CRC_OUT_9_28, CRC_OUT_9_11, n6368, n6333, CRC_OUT_9_27, CRC_OUT_9_10, n6332, n6366, n6330, CRC_OUT_9_26, CRC_OUT_9_9, n6364_1, n6328, CRC_OUT_9_25, CRC_OUT_9_8, n6362, n6326, CRC_OUT_9_7, n6324_1, CRC_OUT_9_6, n6322, CRC_OUT_9_5, n6320, CRC_OUT_9_4, n6318, CRC_OUT_9_3, n6317, n6315, CRC_OUT_9_2, n6313, CRC_OUT_9_1, n6311, CRC_OUT_9_0, n6309_1;
NOR2X1   g0377(.A(n5923), .B(n5827), .Y(n906));
INVX1    g0288(.A(RESET), .Y(n5827));
MX2X1    g0376(.A(n5920), .B(n5922), .S0(TM1), .Y(n5923));
MX2X1    g0375(.A(n5921_1), .B(n5600), .S0(n5539), .Y(n5922));
MX2X1    g0373(.A(n5913), .B(n5918), .S0(n5539), .Y(n5920));
INVX1    g0000(.A(TM0), .Y(n5539));
XOR2X1   g0061(.A(n5599), .B(n5597), .Y(n5600));
INVX1    g0374(.A(WX499), .Y(n5921_1));
XOR2X1   g0372(.A(n5917), .B(n5915), .Y(n5918));
INVX1    g0367(.A(CRC_OUT_9_24), .Y(n5913));
XOR2X1   g0058(.A(n5596_1), .B(WX723), .Y(n5597));
XOR2X1   g0060(.A(WX851), .B(n5598), .Y(n5599));
XOR2X1   g0369(.A(n5914), .B(WX2016), .Y(n5915));
XOR2X1   g0371(.A(WX2144), .B(n5916_1), .Y(n5917));
NOR2X1   g0790(.A(n6360), .B(n5827), .Y(CRC_OUT_9_24));
XOR2X1   g0057(.A(WX659), .B(TM1), .Y(n5596_1));
INVX1    g0059(.A(WX787), .Y(n5598));
XOR2X1   g0368(.A(WX1952), .B(TM1), .Y(n5914));
INVX1    g0370(.A(WX2080), .Y(n5916_1));
XOR2X1   g0789(.A(CRC_OUT_9_23), .B(WX851), .Y(n6360));
NOR2X1   g0788(.A(n6358), .B(n5827), .Y(CRC_OUT_9_23));
XOR2X1   g0787(.A(CRC_OUT_9_22), .B(WX853), .Y(n6358));
NOR2X1   g0786(.A(n6356), .B(n5827), .Y(CRC_OUT_9_22));
XOR2X1   g0785(.A(CRC_OUT_9_21), .B(WX855), .Y(n6356));
NOR2X1   g0784(.A(n6354_1), .B(n5827), .Y(CRC_OUT_9_21));
XOR2X1   g0783(.A(CRC_OUT_9_20), .B(WX857), .Y(n6354_1));
NOR2X1   g0782(.A(n6352), .B(n5827), .Y(CRC_OUT_9_20));
XOR2X1   g0781(.A(CRC_OUT_9_19), .B(WX859), .Y(n6352));
NOR2X1   g0780(.A(n6350), .B(n5827), .Y(CRC_OUT_9_19));
XOR2X1   g0779(.A(CRC_OUT_9_18), .B(WX861), .Y(n6350));
NOR2X1   g0778(.A(n6348), .B(n5827), .Y(CRC_OUT_9_18));
XOR2X1   g0777(.A(CRC_OUT_9_17), .B(WX863), .Y(n6348));
NOR2X1   g0776(.A(n6346), .B(n5827), .Y(CRC_OUT_9_17));
XOR2X1   g0775(.A(CRC_OUT_9_16), .B(WX865), .Y(n6346));
NOR2X1   g0774(.A(n6344_1), .B(n5827), .Y(CRC_OUT_9_16));
XOR2X1   g0773(.A(n6343), .B(CRC_OUT_9_15), .Y(n6344_1));
NOR2X1   g0771(.A(n6341), .B(n5827), .Y(CRC_OUT_9_15));
XOR2X1   g0772(.A(CRC_OUT_9_31), .B(WX867), .Y(n6343));
XOR2X1   g0770(.A(CRC_OUT_9_14), .B(WX869), .Y(n6341));
NOR2X1   g0804(.A(n6374_1), .B(n5827), .Y(CRC_OUT_9_31));
NOR2X1   g0769(.A(n6339_1), .B(n5827), .Y(CRC_OUT_9_14));
XOR2X1   g0803(.A(CRC_OUT_9_30), .B(WX837), .Y(n6374_1));
XOR2X1   g0768(.A(CRC_OUT_9_13), .B(WX871), .Y(n6339_1));
NOR2X1   g0802(.A(n6372), .B(n5827), .Y(CRC_OUT_9_30));
NOR2X1   g0767(.A(n6337), .B(n5827), .Y(CRC_OUT_9_13));
XOR2X1   g0801(.A(CRC_OUT_9_29), .B(WX839), .Y(n6372));
XOR2X1   g0766(.A(CRC_OUT_9_12), .B(WX873), .Y(n6337));
NOR2X1   g0800(.A(n6370), .B(n5827), .Y(CRC_OUT_9_29));
NOR2X1   g0765(.A(n6335), .B(n5827), .Y(CRC_OUT_9_12));
XOR2X1   g0799(.A(CRC_OUT_9_28), .B(WX841), .Y(n6370));
XOR2X1   g0764(.A(CRC_OUT_9_11), .B(WX875), .Y(n6335));
NOR2X1   g0798(.A(n6368), .B(n5827), .Y(CRC_OUT_9_28));
NOR2X1   g0763(.A(n6333), .B(n5827), .Y(CRC_OUT_9_11));
XOR2X1   g0797(.A(CRC_OUT_9_27), .B(WX843), .Y(n6368));
XOR2X1   g0762(.A(n6332), .B(CRC_OUT_9_10), .Y(n6333));
NOR2X1   g0796(.A(n6366), .B(n5827), .Y(CRC_OUT_9_27));
NOR2X1   g0760(.A(n6330), .B(n5827), .Y(CRC_OUT_9_10));
XOR2X1   g0761(.A(CRC_OUT_9_31), .B(WX877), .Y(n6332));
XOR2X1   g0795(.A(CRC_OUT_9_26), .B(WX845), .Y(n6366));
XOR2X1   g0759(.A(CRC_OUT_9_9), .B(WX879), .Y(n6330));
NOR2X1   g0794(.A(n6364_1), .B(n5827), .Y(CRC_OUT_9_26));
NOR2X1   g0758(.A(n6328), .B(n5827), .Y(CRC_OUT_9_9));
XOR2X1   g0793(.A(CRC_OUT_9_25), .B(WX847), .Y(n6364_1));
XOR2X1   g0757(.A(CRC_OUT_9_8), .B(WX881), .Y(n6328));
NOR2X1   g0792(.A(n6362), .B(n5827), .Y(CRC_OUT_9_25));
NOR2X1   g0756(.A(n6326), .B(n5827), .Y(CRC_OUT_9_8));
XOR2X1   g0791(.A(CRC_OUT_9_24), .B(WX849), .Y(n6362));
XOR2X1   g0755(.A(CRC_OUT_9_7), .B(WX883), .Y(n6326));
NOR2X1   g0754(.A(n6324_1), .B(n5827), .Y(CRC_OUT_9_7));
XOR2X1   g0753(.A(CRC_OUT_9_6), .B(WX885), .Y(n6324_1));
NOR2X1   g0752(.A(n6322), .B(n5827), .Y(CRC_OUT_9_6));
XOR2X1   g0751(.A(CRC_OUT_9_5), .B(WX887), .Y(n6322));
NOR2X1   g0750(.A(n6320), .B(n5827), .Y(CRC_OUT_9_5));
XOR2X1   g0749(.A(CRC_OUT_9_4), .B(WX889), .Y(n6320));
NOR2X1   g0748(.A(n6318), .B(n5827), .Y(CRC_OUT_9_4));
XOR2X1   g0747(.A(n6317), .B(CRC_OUT_9_3), .Y(n6318));
NOR2X1   g0745(.A(n6315), .B(n5827), .Y(CRC_OUT_9_3));
XOR2X1   g0746(.A(CRC_OUT_9_31), .B(WX891), .Y(n6317));
XOR2X1   g0744(.A(CRC_OUT_9_2), .B(WX893), .Y(n6315));
NOR2X1   g0743(.A(n6313), .B(n5827), .Y(CRC_OUT_9_2));
XOR2X1   g0742(.A(CRC_OUT_9_1), .B(WX895), .Y(n6313));
NOR2X1   g0741(.A(n6311), .B(n5827), .Y(CRC_OUT_9_1));
XOR2X1   g0740(.A(CRC_OUT_9_0), .B(WX897), .Y(n6311));
NOR2X1   g0739(.A(n6309_1), .B(n5827), .Y(CRC_OUT_9_0));
XOR2X1   g0738(.A(CRC_OUT_9_31), .B(WX899), .Y(n6309_1));

endmodule
