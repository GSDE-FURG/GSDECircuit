// Benchmark "top" written by ABC on Mon Sep 21 03:35:54 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] ,
    \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] ,
    \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] ,
    \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] ,
    \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] ,
    \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] ,
    \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] ,
    \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] ,
    \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] ,
    \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] ,
    \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] ,
    \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] ,
    \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] ,
    \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] ,
    \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] ,
    \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] ,
    \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] ,
    \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] ,
    \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] ,
    \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] ,
    \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] ,
    \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127] , cOut  );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] ,
    \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] ,
    \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] ,
    \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] ,
    \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] ,
    \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] ,
    \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] ,
    \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] ,
    \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] ,
    \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] ,
    \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] ,
    \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] ,
    \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] ,
    \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] ,
    \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] ,
    \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] ,
    \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] ,
    \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] ,
    \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] ,
    \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] ,
    \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] ,
    \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] ,
    \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] ,
    \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] ,
    \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] , cOut;
  wire new_n387_, new_n388_, new_n389_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n403_, new_n404_, new_n405_, new_n407_, new_n408_,
    new_n409_, new_n410_, new_n411_, new_n412_, new_n413_, new_n415_,
    new_n416_, new_n417_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n427_, new_n428_, new_n429_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n439_, new_n440_, new_n441_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n451_,
    new_n452_, new_n453_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n463_, new_n464_, new_n465_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n475_, new_n476_, new_n477_, new_n479_, new_n480_,
    new_n481_, new_n482_, new_n483_, new_n484_, new_n485_, new_n487_,
    new_n488_, new_n489_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n499_, new_n500_, new_n501_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n511_, new_n512_, new_n513_, new_n515_, new_n516_,
    new_n517_, new_n518_, new_n519_, new_n520_, new_n521_, new_n523_,
    new_n524_, new_n525_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n535_, new_n536_, new_n537_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n547_, new_n548_, new_n549_, new_n551_, new_n552_,
    new_n553_, new_n554_, new_n555_, new_n556_, new_n557_, new_n559_,
    new_n560_, new_n561_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n571_, new_n572_, new_n573_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n583_, new_n584_, new_n585_, new_n587_, new_n588_,
    new_n589_, new_n590_, new_n591_, new_n592_, new_n593_, new_n595_,
    new_n596_, new_n597_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n607_, new_n608_, new_n609_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n619_, new_n620_, new_n621_, new_n623_, new_n624_,
    new_n625_, new_n626_, new_n627_, new_n628_, new_n629_, new_n631_,
    new_n632_, new_n633_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n643_, new_n644_, new_n645_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n655_, new_n656_, new_n657_, new_n659_, new_n660_,
    new_n661_, new_n662_, new_n663_, new_n664_, new_n665_, new_n667_,
    new_n668_, new_n669_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n679_, new_n680_, new_n681_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n691_, new_n692_, new_n693_, new_n695_, new_n696_,
    new_n697_, new_n698_, new_n699_, new_n700_, new_n701_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n715_, new_n716_, new_n717_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n727_, new_n728_, new_n729_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n739_,
    new_n740_, new_n741_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n751_, new_n752_, new_n753_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n763_, new_n764_, new_n765_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n775_,
    new_n776_, new_n777_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n787_, new_n788_, new_n789_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n799_, new_n800_, new_n801_, new_n803_, new_n804_,
    new_n805_, new_n806_, new_n807_, new_n808_, new_n809_, new_n811_,
    new_n812_, new_n813_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n823_, new_n824_, new_n825_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n835_, new_n836_, new_n837_, new_n839_, new_n840_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n847_,
    new_n848_, new_n849_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n859_, new_n860_, new_n861_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n871_, new_n872_, new_n873_, new_n875_, new_n876_,
    new_n877_, new_n878_, new_n879_, new_n880_, new_n881_, new_n883_,
    new_n884_, new_n885_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n895_, new_n896_, new_n897_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n907_, new_n908_, new_n909_, new_n911_, new_n912_,
    new_n913_, new_n914_, new_n915_, new_n916_, new_n917_, new_n919_,
    new_n920_, new_n921_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n931_, new_n932_, new_n933_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n943_, new_n944_, new_n945_, new_n947_, new_n948_,
    new_n949_, new_n950_, new_n951_, new_n952_, new_n953_, new_n955_,
    new_n956_, new_n957_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n967_, new_n968_, new_n969_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n979_, new_n980_, new_n981_, new_n983_, new_n984_,
    new_n985_, new_n986_, new_n987_, new_n988_, new_n989_, new_n991_,
    new_n992_, new_n993_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1003_, new_n1004_, new_n1005_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1015_, new_n1016_, new_n1017_, new_n1019_, new_n1020_,
    new_n1021_, new_n1022_, new_n1023_, new_n1024_, new_n1025_, new_n1027_,
    new_n1028_, new_n1029_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1039_, new_n1040_, new_n1041_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1051_, new_n1052_, new_n1053_, new_n1055_, new_n1056_,
    new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_, new_n1063_,
    new_n1064_, new_n1065_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1075_, new_n1076_, new_n1077_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1087_, new_n1088_, new_n1089_, new_n1091_, new_n1092_,
    new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_, new_n1099_,
    new_n1100_, new_n1101_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1111_, new_n1112_, new_n1113_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1123_, new_n1124_, new_n1125_, new_n1127_, new_n1128_,
    new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_, new_n1135_,
    new_n1136_, new_n1137_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1146_, new_n1147_;
  XOR2X1   g000(.A(\b[0] ), .B(\a[0] ), .Y(\f[0] ));
  NAND2X1  g001(.A(\b[0] ), .B(\a[0] ), .Y(new_n387_));
  INVX1    g002(.A(new_n387_), .Y(new_n388_));
  XOR2X1   g003(.A(\b[1] ), .B(\a[1] ), .Y(new_n389_));
  XOR2X1   g004(.A(new_n389_), .B(new_n388_), .Y(\f[1] ));
  NOR2X1   g005(.A(\b[1] ), .B(\a[1] ), .Y(new_n391_));
  NAND2X1  g006(.A(\b[1] ), .B(\a[1] ), .Y(new_n392_));
  OAI21X1  g007(.A0(new_n391_), .A1(new_n387_), .B0(new_n392_), .Y(new_n393_));
  XOR2X1   g008(.A(\b[2] ), .B(\a[2] ), .Y(new_n394_));
  XOR2X1   g009(.A(new_n394_), .B(new_n393_), .Y(\f[2] ));
  OR2X1    g010(.A(\b[2] ), .B(\a[2] ), .Y(new_n396_));
  AND2X1   g011(.A(\b[2] ), .B(\a[2] ), .Y(new_n397_));
  AOI21X1  g012(.A0(new_n396_), .A1(new_n393_), .B0(new_n397_), .Y(new_n398_));
  NOR2X1   g013(.A(\b[3] ), .B(\a[3] ), .Y(new_n399_));
  AND2X1   g014(.A(\b[3] ), .B(\a[3] ), .Y(new_n400_));
  OR2X1    g015(.A(new_n400_), .B(new_n399_), .Y(new_n401_));
  XOR2X1   g016(.A(new_n401_), .B(new_n398_), .Y(\f[3] ));
  INVX1    g017(.A(new_n400_), .Y(new_n403_));
  OAI21X1  g018(.A0(new_n399_), .A1(new_n398_), .B0(new_n403_), .Y(new_n404_));
  XOR2X1   g019(.A(\b[4] ), .B(\a[4] ), .Y(new_n405_));
  XOR2X1   g020(.A(new_n405_), .B(new_n404_), .Y(\f[4] ));
  NOR2X1   g021(.A(\b[4] ), .B(\a[4] ), .Y(new_n407_));
  INVX1    g022(.A(new_n407_), .Y(new_n408_));
  AND2X1   g023(.A(\b[4] ), .B(\a[4] ), .Y(new_n409_));
  AOI21X1  g024(.A0(new_n408_), .A1(new_n404_), .B0(new_n409_), .Y(new_n410_));
  NOR2X1   g025(.A(\b[5] ), .B(\a[5] ), .Y(new_n411_));
  AND2X1   g026(.A(\b[5] ), .B(\a[5] ), .Y(new_n412_));
  OR2X1    g027(.A(new_n412_), .B(new_n411_), .Y(new_n413_));
  XOR2X1   g028(.A(new_n413_), .B(new_n410_), .Y(\f[5] ));
  INVX1    g029(.A(new_n412_), .Y(new_n415_));
  OAI21X1  g030(.A0(new_n411_), .A1(new_n410_), .B0(new_n415_), .Y(new_n416_));
  XOR2X1   g031(.A(\b[6] ), .B(\a[6] ), .Y(new_n417_));
  XOR2X1   g032(.A(new_n417_), .B(new_n416_), .Y(\f[6] ));
  NOR2X1   g033(.A(\b[6] ), .B(\a[6] ), .Y(new_n419_));
  INVX1    g034(.A(new_n419_), .Y(new_n420_));
  AND2X1   g035(.A(\b[6] ), .B(\a[6] ), .Y(new_n421_));
  AOI21X1  g036(.A0(new_n420_), .A1(new_n416_), .B0(new_n421_), .Y(new_n422_));
  NOR2X1   g037(.A(\b[7] ), .B(\a[7] ), .Y(new_n423_));
  AND2X1   g038(.A(\b[7] ), .B(\a[7] ), .Y(new_n424_));
  OR2X1    g039(.A(new_n424_), .B(new_n423_), .Y(new_n425_));
  XOR2X1   g040(.A(new_n425_), .B(new_n422_), .Y(\f[7] ));
  INVX1    g041(.A(new_n424_), .Y(new_n427_));
  OAI21X1  g042(.A0(new_n423_), .A1(new_n422_), .B0(new_n427_), .Y(new_n428_));
  XOR2X1   g043(.A(\b[8] ), .B(\a[8] ), .Y(new_n429_));
  XOR2X1   g044(.A(new_n429_), .B(new_n428_), .Y(\f[8] ));
  NOR2X1   g045(.A(\b[8] ), .B(\a[8] ), .Y(new_n431_));
  INVX1    g046(.A(new_n431_), .Y(new_n432_));
  AND2X1   g047(.A(\b[8] ), .B(\a[8] ), .Y(new_n433_));
  AOI21X1  g048(.A0(new_n432_), .A1(new_n428_), .B0(new_n433_), .Y(new_n434_));
  NOR2X1   g049(.A(\b[9] ), .B(\a[9] ), .Y(new_n435_));
  AND2X1   g050(.A(\b[9] ), .B(\a[9] ), .Y(new_n436_));
  OR2X1    g051(.A(new_n436_), .B(new_n435_), .Y(new_n437_));
  XOR2X1   g052(.A(new_n437_), .B(new_n434_), .Y(\f[9] ));
  INVX1    g053(.A(new_n436_), .Y(new_n439_));
  OAI21X1  g054(.A0(new_n435_), .A1(new_n434_), .B0(new_n439_), .Y(new_n440_));
  XOR2X1   g055(.A(\b[10] ), .B(\a[10] ), .Y(new_n441_));
  XOR2X1   g056(.A(new_n441_), .B(new_n440_), .Y(\f[10] ));
  NOR2X1   g057(.A(\b[10] ), .B(\a[10] ), .Y(new_n443_));
  INVX1    g058(.A(new_n443_), .Y(new_n444_));
  AND2X1   g059(.A(\b[10] ), .B(\a[10] ), .Y(new_n445_));
  AOI21X1  g060(.A0(new_n444_), .A1(new_n440_), .B0(new_n445_), .Y(new_n446_));
  NOR2X1   g061(.A(\b[11] ), .B(\a[11] ), .Y(new_n447_));
  AND2X1   g062(.A(\b[11] ), .B(\a[11] ), .Y(new_n448_));
  OR2X1    g063(.A(new_n448_), .B(new_n447_), .Y(new_n449_));
  XOR2X1   g064(.A(new_n449_), .B(new_n446_), .Y(\f[11] ));
  INVX1    g065(.A(new_n448_), .Y(new_n451_));
  OAI21X1  g066(.A0(new_n447_), .A1(new_n446_), .B0(new_n451_), .Y(new_n452_));
  XOR2X1   g067(.A(\b[12] ), .B(\a[12] ), .Y(new_n453_));
  XOR2X1   g068(.A(new_n453_), .B(new_n452_), .Y(\f[12] ));
  NOR2X1   g069(.A(\b[12] ), .B(\a[12] ), .Y(new_n455_));
  INVX1    g070(.A(new_n455_), .Y(new_n456_));
  AND2X1   g071(.A(\b[12] ), .B(\a[12] ), .Y(new_n457_));
  AOI21X1  g072(.A0(new_n456_), .A1(new_n452_), .B0(new_n457_), .Y(new_n458_));
  NOR2X1   g073(.A(\b[13] ), .B(\a[13] ), .Y(new_n459_));
  AND2X1   g074(.A(\b[13] ), .B(\a[13] ), .Y(new_n460_));
  OR2X1    g075(.A(new_n460_), .B(new_n459_), .Y(new_n461_));
  XOR2X1   g076(.A(new_n461_), .B(new_n458_), .Y(\f[13] ));
  INVX1    g077(.A(new_n460_), .Y(new_n463_));
  OAI21X1  g078(.A0(new_n459_), .A1(new_n458_), .B0(new_n463_), .Y(new_n464_));
  XOR2X1   g079(.A(\b[14] ), .B(\a[14] ), .Y(new_n465_));
  XOR2X1   g080(.A(new_n465_), .B(new_n464_), .Y(\f[14] ));
  NOR2X1   g081(.A(\b[14] ), .B(\a[14] ), .Y(new_n467_));
  INVX1    g082(.A(new_n467_), .Y(new_n468_));
  AND2X1   g083(.A(\b[14] ), .B(\a[14] ), .Y(new_n469_));
  AOI21X1  g084(.A0(new_n468_), .A1(new_n464_), .B0(new_n469_), .Y(new_n470_));
  NOR2X1   g085(.A(\b[15] ), .B(\a[15] ), .Y(new_n471_));
  AND2X1   g086(.A(\b[15] ), .B(\a[15] ), .Y(new_n472_));
  OR2X1    g087(.A(new_n472_), .B(new_n471_), .Y(new_n473_));
  XOR2X1   g088(.A(new_n473_), .B(new_n470_), .Y(\f[15] ));
  INVX1    g089(.A(new_n472_), .Y(new_n475_));
  OAI21X1  g090(.A0(new_n471_), .A1(new_n470_), .B0(new_n475_), .Y(new_n476_));
  XOR2X1   g091(.A(\b[16] ), .B(\a[16] ), .Y(new_n477_));
  XOR2X1   g092(.A(new_n477_), .B(new_n476_), .Y(\f[16] ));
  NOR2X1   g093(.A(\b[16] ), .B(\a[16] ), .Y(new_n479_));
  INVX1    g094(.A(new_n479_), .Y(new_n480_));
  AND2X1   g095(.A(\b[16] ), .B(\a[16] ), .Y(new_n481_));
  AOI21X1  g096(.A0(new_n480_), .A1(new_n476_), .B0(new_n481_), .Y(new_n482_));
  NOR2X1   g097(.A(\b[17] ), .B(\a[17] ), .Y(new_n483_));
  AND2X1   g098(.A(\b[17] ), .B(\a[17] ), .Y(new_n484_));
  OR2X1    g099(.A(new_n484_), .B(new_n483_), .Y(new_n485_));
  XOR2X1   g100(.A(new_n485_), .B(new_n482_), .Y(\f[17] ));
  INVX1    g101(.A(new_n484_), .Y(new_n487_));
  OAI21X1  g102(.A0(new_n483_), .A1(new_n482_), .B0(new_n487_), .Y(new_n488_));
  XOR2X1   g103(.A(\b[18] ), .B(\a[18] ), .Y(new_n489_));
  XOR2X1   g104(.A(new_n489_), .B(new_n488_), .Y(\f[18] ));
  NOR2X1   g105(.A(\b[18] ), .B(\a[18] ), .Y(new_n491_));
  INVX1    g106(.A(new_n491_), .Y(new_n492_));
  AND2X1   g107(.A(\b[18] ), .B(\a[18] ), .Y(new_n493_));
  AOI21X1  g108(.A0(new_n492_), .A1(new_n488_), .B0(new_n493_), .Y(new_n494_));
  NOR2X1   g109(.A(\b[19] ), .B(\a[19] ), .Y(new_n495_));
  AND2X1   g110(.A(\b[19] ), .B(\a[19] ), .Y(new_n496_));
  OR2X1    g111(.A(new_n496_), .B(new_n495_), .Y(new_n497_));
  XOR2X1   g112(.A(new_n497_), .B(new_n494_), .Y(\f[19] ));
  INVX1    g113(.A(new_n496_), .Y(new_n499_));
  OAI21X1  g114(.A0(new_n495_), .A1(new_n494_), .B0(new_n499_), .Y(new_n500_));
  XOR2X1   g115(.A(\b[20] ), .B(\a[20] ), .Y(new_n501_));
  XOR2X1   g116(.A(new_n501_), .B(new_n500_), .Y(\f[20] ));
  NOR2X1   g117(.A(\b[20] ), .B(\a[20] ), .Y(new_n503_));
  INVX1    g118(.A(new_n503_), .Y(new_n504_));
  AND2X1   g119(.A(\b[20] ), .B(\a[20] ), .Y(new_n505_));
  AOI21X1  g120(.A0(new_n504_), .A1(new_n500_), .B0(new_n505_), .Y(new_n506_));
  NOR2X1   g121(.A(\b[21] ), .B(\a[21] ), .Y(new_n507_));
  AND2X1   g122(.A(\b[21] ), .B(\a[21] ), .Y(new_n508_));
  OR2X1    g123(.A(new_n508_), .B(new_n507_), .Y(new_n509_));
  XOR2X1   g124(.A(new_n509_), .B(new_n506_), .Y(\f[21] ));
  INVX1    g125(.A(new_n508_), .Y(new_n511_));
  OAI21X1  g126(.A0(new_n507_), .A1(new_n506_), .B0(new_n511_), .Y(new_n512_));
  XOR2X1   g127(.A(\b[22] ), .B(\a[22] ), .Y(new_n513_));
  XOR2X1   g128(.A(new_n513_), .B(new_n512_), .Y(\f[22] ));
  NOR2X1   g129(.A(\b[22] ), .B(\a[22] ), .Y(new_n515_));
  INVX1    g130(.A(new_n515_), .Y(new_n516_));
  AND2X1   g131(.A(\b[22] ), .B(\a[22] ), .Y(new_n517_));
  AOI21X1  g132(.A0(new_n516_), .A1(new_n512_), .B0(new_n517_), .Y(new_n518_));
  NOR2X1   g133(.A(\b[23] ), .B(\a[23] ), .Y(new_n519_));
  AND2X1   g134(.A(\b[23] ), .B(\a[23] ), .Y(new_n520_));
  OR2X1    g135(.A(new_n520_), .B(new_n519_), .Y(new_n521_));
  XOR2X1   g136(.A(new_n521_), .B(new_n518_), .Y(\f[23] ));
  INVX1    g137(.A(new_n520_), .Y(new_n523_));
  OAI21X1  g138(.A0(new_n519_), .A1(new_n518_), .B0(new_n523_), .Y(new_n524_));
  XOR2X1   g139(.A(\b[24] ), .B(\a[24] ), .Y(new_n525_));
  XOR2X1   g140(.A(new_n525_), .B(new_n524_), .Y(\f[24] ));
  NOR2X1   g141(.A(\b[24] ), .B(\a[24] ), .Y(new_n527_));
  INVX1    g142(.A(new_n527_), .Y(new_n528_));
  AND2X1   g143(.A(\b[24] ), .B(\a[24] ), .Y(new_n529_));
  AOI21X1  g144(.A0(new_n528_), .A1(new_n524_), .B0(new_n529_), .Y(new_n530_));
  NOR2X1   g145(.A(\b[25] ), .B(\a[25] ), .Y(new_n531_));
  AND2X1   g146(.A(\b[25] ), .B(\a[25] ), .Y(new_n532_));
  OR2X1    g147(.A(new_n532_), .B(new_n531_), .Y(new_n533_));
  XOR2X1   g148(.A(new_n533_), .B(new_n530_), .Y(\f[25] ));
  INVX1    g149(.A(new_n532_), .Y(new_n535_));
  OAI21X1  g150(.A0(new_n531_), .A1(new_n530_), .B0(new_n535_), .Y(new_n536_));
  XOR2X1   g151(.A(\b[26] ), .B(\a[26] ), .Y(new_n537_));
  XOR2X1   g152(.A(new_n537_), .B(new_n536_), .Y(\f[26] ));
  NOR2X1   g153(.A(\b[26] ), .B(\a[26] ), .Y(new_n539_));
  INVX1    g154(.A(new_n539_), .Y(new_n540_));
  AND2X1   g155(.A(\b[26] ), .B(\a[26] ), .Y(new_n541_));
  AOI21X1  g156(.A0(new_n540_), .A1(new_n536_), .B0(new_n541_), .Y(new_n542_));
  NOR2X1   g157(.A(\b[27] ), .B(\a[27] ), .Y(new_n543_));
  AND2X1   g158(.A(\b[27] ), .B(\a[27] ), .Y(new_n544_));
  OR2X1    g159(.A(new_n544_), .B(new_n543_), .Y(new_n545_));
  XOR2X1   g160(.A(new_n545_), .B(new_n542_), .Y(\f[27] ));
  INVX1    g161(.A(new_n544_), .Y(new_n547_));
  OAI21X1  g162(.A0(new_n543_), .A1(new_n542_), .B0(new_n547_), .Y(new_n548_));
  XOR2X1   g163(.A(\b[28] ), .B(\a[28] ), .Y(new_n549_));
  XOR2X1   g164(.A(new_n549_), .B(new_n548_), .Y(\f[28] ));
  NOR2X1   g165(.A(\b[28] ), .B(\a[28] ), .Y(new_n551_));
  INVX1    g166(.A(new_n551_), .Y(new_n552_));
  AND2X1   g167(.A(\b[28] ), .B(\a[28] ), .Y(new_n553_));
  AOI21X1  g168(.A0(new_n552_), .A1(new_n548_), .B0(new_n553_), .Y(new_n554_));
  NOR2X1   g169(.A(\b[29] ), .B(\a[29] ), .Y(new_n555_));
  AND2X1   g170(.A(\b[29] ), .B(\a[29] ), .Y(new_n556_));
  OR2X1    g171(.A(new_n556_), .B(new_n555_), .Y(new_n557_));
  XOR2X1   g172(.A(new_n557_), .B(new_n554_), .Y(\f[29] ));
  INVX1    g173(.A(new_n556_), .Y(new_n559_));
  OAI21X1  g174(.A0(new_n555_), .A1(new_n554_), .B0(new_n559_), .Y(new_n560_));
  XOR2X1   g175(.A(\b[30] ), .B(\a[30] ), .Y(new_n561_));
  XOR2X1   g176(.A(new_n561_), .B(new_n560_), .Y(\f[30] ));
  NOR2X1   g177(.A(\b[30] ), .B(\a[30] ), .Y(new_n563_));
  INVX1    g178(.A(new_n563_), .Y(new_n564_));
  AND2X1   g179(.A(\b[30] ), .B(\a[30] ), .Y(new_n565_));
  AOI21X1  g180(.A0(new_n564_), .A1(new_n560_), .B0(new_n565_), .Y(new_n566_));
  NOR2X1   g181(.A(\b[31] ), .B(\a[31] ), .Y(new_n567_));
  AND2X1   g182(.A(\b[31] ), .B(\a[31] ), .Y(new_n568_));
  OR2X1    g183(.A(new_n568_), .B(new_n567_), .Y(new_n569_));
  XOR2X1   g184(.A(new_n569_), .B(new_n566_), .Y(\f[31] ));
  INVX1    g185(.A(new_n568_), .Y(new_n571_));
  OAI21X1  g186(.A0(new_n567_), .A1(new_n566_), .B0(new_n571_), .Y(new_n572_));
  XOR2X1   g187(.A(\b[32] ), .B(\a[32] ), .Y(new_n573_));
  XOR2X1   g188(.A(new_n573_), .B(new_n572_), .Y(\f[32] ));
  NOR2X1   g189(.A(\b[32] ), .B(\a[32] ), .Y(new_n575_));
  INVX1    g190(.A(new_n575_), .Y(new_n576_));
  AND2X1   g191(.A(\b[32] ), .B(\a[32] ), .Y(new_n577_));
  AOI21X1  g192(.A0(new_n576_), .A1(new_n572_), .B0(new_n577_), .Y(new_n578_));
  NOR2X1   g193(.A(\b[33] ), .B(\a[33] ), .Y(new_n579_));
  AND2X1   g194(.A(\b[33] ), .B(\a[33] ), .Y(new_n580_));
  OR2X1    g195(.A(new_n580_), .B(new_n579_), .Y(new_n581_));
  XOR2X1   g196(.A(new_n581_), .B(new_n578_), .Y(\f[33] ));
  INVX1    g197(.A(new_n580_), .Y(new_n583_));
  OAI21X1  g198(.A0(new_n579_), .A1(new_n578_), .B0(new_n583_), .Y(new_n584_));
  XOR2X1   g199(.A(\b[34] ), .B(\a[34] ), .Y(new_n585_));
  XOR2X1   g200(.A(new_n585_), .B(new_n584_), .Y(\f[34] ));
  NOR2X1   g201(.A(\b[34] ), .B(\a[34] ), .Y(new_n587_));
  INVX1    g202(.A(new_n587_), .Y(new_n588_));
  AND2X1   g203(.A(\b[34] ), .B(\a[34] ), .Y(new_n589_));
  AOI21X1  g204(.A0(new_n588_), .A1(new_n584_), .B0(new_n589_), .Y(new_n590_));
  NOR2X1   g205(.A(\b[35] ), .B(\a[35] ), .Y(new_n591_));
  AND2X1   g206(.A(\b[35] ), .B(\a[35] ), .Y(new_n592_));
  OR2X1    g207(.A(new_n592_), .B(new_n591_), .Y(new_n593_));
  XOR2X1   g208(.A(new_n593_), .B(new_n590_), .Y(\f[35] ));
  INVX1    g209(.A(new_n592_), .Y(new_n595_));
  OAI21X1  g210(.A0(new_n591_), .A1(new_n590_), .B0(new_n595_), .Y(new_n596_));
  XOR2X1   g211(.A(\b[36] ), .B(\a[36] ), .Y(new_n597_));
  XOR2X1   g212(.A(new_n597_), .B(new_n596_), .Y(\f[36] ));
  NOR2X1   g213(.A(\b[36] ), .B(\a[36] ), .Y(new_n599_));
  INVX1    g214(.A(new_n599_), .Y(new_n600_));
  AND2X1   g215(.A(\b[36] ), .B(\a[36] ), .Y(new_n601_));
  AOI21X1  g216(.A0(new_n600_), .A1(new_n596_), .B0(new_n601_), .Y(new_n602_));
  NOR2X1   g217(.A(\b[37] ), .B(\a[37] ), .Y(new_n603_));
  AND2X1   g218(.A(\b[37] ), .B(\a[37] ), .Y(new_n604_));
  OR2X1    g219(.A(new_n604_), .B(new_n603_), .Y(new_n605_));
  XOR2X1   g220(.A(new_n605_), .B(new_n602_), .Y(\f[37] ));
  INVX1    g221(.A(new_n604_), .Y(new_n607_));
  OAI21X1  g222(.A0(new_n603_), .A1(new_n602_), .B0(new_n607_), .Y(new_n608_));
  XOR2X1   g223(.A(\b[38] ), .B(\a[38] ), .Y(new_n609_));
  XOR2X1   g224(.A(new_n609_), .B(new_n608_), .Y(\f[38] ));
  NOR2X1   g225(.A(\b[38] ), .B(\a[38] ), .Y(new_n611_));
  INVX1    g226(.A(new_n611_), .Y(new_n612_));
  AND2X1   g227(.A(\b[38] ), .B(\a[38] ), .Y(new_n613_));
  AOI21X1  g228(.A0(new_n612_), .A1(new_n608_), .B0(new_n613_), .Y(new_n614_));
  NOR2X1   g229(.A(\b[39] ), .B(\a[39] ), .Y(new_n615_));
  AND2X1   g230(.A(\b[39] ), .B(\a[39] ), .Y(new_n616_));
  OR2X1    g231(.A(new_n616_), .B(new_n615_), .Y(new_n617_));
  XOR2X1   g232(.A(new_n617_), .B(new_n614_), .Y(\f[39] ));
  INVX1    g233(.A(new_n616_), .Y(new_n619_));
  OAI21X1  g234(.A0(new_n615_), .A1(new_n614_), .B0(new_n619_), .Y(new_n620_));
  XOR2X1   g235(.A(\b[40] ), .B(\a[40] ), .Y(new_n621_));
  XOR2X1   g236(.A(new_n621_), .B(new_n620_), .Y(\f[40] ));
  NOR2X1   g237(.A(\b[40] ), .B(\a[40] ), .Y(new_n623_));
  INVX1    g238(.A(new_n623_), .Y(new_n624_));
  AND2X1   g239(.A(\b[40] ), .B(\a[40] ), .Y(new_n625_));
  AOI21X1  g240(.A0(new_n624_), .A1(new_n620_), .B0(new_n625_), .Y(new_n626_));
  NOR2X1   g241(.A(\b[41] ), .B(\a[41] ), .Y(new_n627_));
  AND2X1   g242(.A(\b[41] ), .B(\a[41] ), .Y(new_n628_));
  OR2X1    g243(.A(new_n628_), .B(new_n627_), .Y(new_n629_));
  XOR2X1   g244(.A(new_n629_), .B(new_n626_), .Y(\f[41] ));
  INVX1    g245(.A(new_n628_), .Y(new_n631_));
  OAI21X1  g246(.A0(new_n627_), .A1(new_n626_), .B0(new_n631_), .Y(new_n632_));
  XOR2X1   g247(.A(\b[42] ), .B(\a[42] ), .Y(new_n633_));
  XOR2X1   g248(.A(new_n633_), .B(new_n632_), .Y(\f[42] ));
  NOR2X1   g249(.A(\b[42] ), .B(\a[42] ), .Y(new_n635_));
  INVX1    g250(.A(new_n635_), .Y(new_n636_));
  AND2X1   g251(.A(\b[42] ), .B(\a[42] ), .Y(new_n637_));
  AOI21X1  g252(.A0(new_n636_), .A1(new_n632_), .B0(new_n637_), .Y(new_n638_));
  NOR2X1   g253(.A(\b[43] ), .B(\a[43] ), .Y(new_n639_));
  AND2X1   g254(.A(\b[43] ), .B(\a[43] ), .Y(new_n640_));
  OR2X1    g255(.A(new_n640_), .B(new_n639_), .Y(new_n641_));
  XOR2X1   g256(.A(new_n641_), .B(new_n638_), .Y(\f[43] ));
  INVX1    g257(.A(new_n640_), .Y(new_n643_));
  OAI21X1  g258(.A0(new_n639_), .A1(new_n638_), .B0(new_n643_), .Y(new_n644_));
  XOR2X1   g259(.A(\b[44] ), .B(\a[44] ), .Y(new_n645_));
  XOR2X1   g260(.A(new_n645_), .B(new_n644_), .Y(\f[44] ));
  NOR2X1   g261(.A(\b[44] ), .B(\a[44] ), .Y(new_n647_));
  INVX1    g262(.A(new_n647_), .Y(new_n648_));
  AND2X1   g263(.A(\b[44] ), .B(\a[44] ), .Y(new_n649_));
  AOI21X1  g264(.A0(new_n648_), .A1(new_n644_), .B0(new_n649_), .Y(new_n650_));
  NOR2X1   g265(.A(\b[45] ), .B(\a[45] ), .Y(new_n651_));
  AND2X1   g266(.A(\b[45] ), .B(\a[45] ), .Y(new_n652_));
  OR2X1    g267(.A(new_n652_), .B(new_n651_), .Y(new_n653_));
  XOR2X1   g268(.A(new_n653_), .B(new_n650_), .Y(\f[45] ));
  INVX1    g269(.A(new_n652_), .Y(new_n655_));
  OAI21X1  g270(.A0(new_n651_), .A1(new_n650_), .B0(new_n655_), .Y(new_n656_));
  XOR2X1   g271(.A(\b[46] ), .B(\a[46] ), .Y(new_n657_));
  XOR2X1   g272(.A(new_n657_), .B(new_n656_), .Y(\f[46] ));
  NOR2X1   g273(.A(\b[46] ), .B(\a[46] ), .Y(new_n659_));
  INVX1    g274(.A(new_n659_), .Y(new_n660_));
  AND2X1   g275(.A(\b[46] ), .B(\a[46] ), .Y(new_n661_));
  AOI21X1  g276(.A0(new_n660_), .A1(new_n656_), .B0(new_n661_), .Y(new_n662_));
  NOR2X1   g277(.A(\b[47] ), .B(\a[47] ), .Y(new_n663_));
  AND2X1   g278(.A(\b[47] ), .B(\a[47] ), .Y(new_n664_));
  OR2X1    g279(.A(new_n664_), .B(new_n663_), .Y(new_n665_));
  XOR2X1   g280(.A(new_n665_), .B(new_n662_), .Y(\f[47] ));
  INVX1    g281(.A(new_n664_), .Y(new_n667_));
  OAI21X1  g282(.A0(new_n663_), .A1(new_n662_), .B0(new_n667_), .Y(new_n668_));
  XOR2X1   g283(.A(\b[48] ), .B(\a[48] ), .Y(new_n669_));
  XOR2X1   g284(.A(new_n669_), .B(new_n668_), .Y(\f[48] ));
  NOR2X1   g285(.A(\b[48] ), .B(\a[48] ), .Y(new_n671_));
  INVX1    g286(.A(new_n671_), .Y(new_n672_));
  AND2X1   g287(.A(\b[48] ), .B(\a[48] ), .Y(new_n673_));
  AOI21X1  g288(.A0(new_n672_), .A1(new_n668_), .B0(new_n673_), .Y(new_n674_));
  NOR2X1   g289(.A(\b[49] ), .B(\a[49] ), .Y(new_n675_));
  AND2X1   g290(.A(\b[49] ), .B(\a[49] ), .Y(new_n676_));
  OR2X1    g291(.A(new_n676_), .B(new_n675_), .Y(new_n677_));
  XOR2X1   g292(.A(new_n677_), .B(new_n674_), .Y(\f[49] ));
  INVX1    g293(.A(new_n676_), .Y(new_n679_));
  OAI21X1  g294(.A0(new_n675_), .A1(new_n674_), .B0(new_n679_), .Y(new_n680_));
  XOR2X1   g295(.A(\b[50] ), .B(\a[50] ), .Y(new_n681_));
  XOR2X1   g296(.A(new_n681_), .B(new_n680_), .Y(\f[50] ));
  NOR2X1   g297(.A(\b[50] ), .B(\a[50] ), .Y(new_n683_));
  INVX1    g298(.A(new_n683_), .Y(new_n684_));
  AND2X1   g299(.A(\b[50] ), .B(\a[50] ), .Y(new_n685_));
  AOI21X1  g300(.A0(new_n684_), .A1(new_n680_), .B0(new_n685_), .Y(new_n686_));
  NOR2X1   g301(.A(\b[51] ), .B(\a[51] ), .Y(new_n687_));
  AND2X1   g302(.A(\b[51] ), .B(\a[51] ), .Y(new_n688_));
  OR2X1    g303(.A(new_n688_), .B(new_n687_), .Y(new_n689_));
  XOR2X1   g304(.A(new_n689_), .B(new_n686_), .Y(\f[51] ));
  INVX1    g305(.A(new_n688_), .Y(new_n691_));
  OAI21X1  g306(.A0(new_n687_), .A1(new_n686_), .B0(new_n691_), .Y(new_n692_));
  XOR2X1   g307(.A(\b[52] ), .B(\a[52] ), .Y(new_n693_));
  XOR2X1   g308(.A(new_n693_), .B(new_n692_), .Y(\f[52] ));
  NOR2X1   g309(.A(\b[52] ), .B(\a[52] ), .Y(new_n695_));
  INVX1    g310(.A(new_n695_), .Y(new_n696_));
  AND2X1   g311(.A(\b[52] ), .B(\a[52] ), .Y(new_n697_));
  AOI21X1  g312(.A0(new_n696_), .A1(new_n692_), .B0(new_n697_), .Y(new_n698_));
  NOR2X1   g313(.A(\b[53] ), .B(\a[53] ), .Y(new_n699_));
  AND2X1   g314(.A(\b[53] ), .B(\a[53] ), .Y(new_n700_));
  OR2X1    g315(.A(new_n700_), .B(new_n699_), .Y(new_n701_));
  XOR2X1   g316(.A(new_n701_), .B(new_n698_), .Y(\f[53] ));
  INVX1    g317(.A(new_n700_), .Y(new_n703_));
  OAI21X1  g318(.A0(new_n699_), .A1(new_n698_), .B0(new_n703_), .Y(new_n704_));
  XOR2X1   g319(.A(\b[54] ), .B(\a[54] ), .Y(new_n705_));
  XOR2X1   g320(.A(new_n705_), .B(new_n704_), .Y(\f[54] ));
  NOR2X1   g321(.A(\b[54] ), .B(\a[54] ), .Y(new_n707_));
  INVX1    g322(.A(new_n707_), .Y(new_n708_));
  AND2X1   g323(.A(\b[54] ), .B(\a[54] ), .Y(new_n709_));
  AOI21X1  g324(.A0(new_n708_), .A1(new_n704_), .B0(new_n709_), .Y(new_n710_));
  NOR2X1   g325(.A(\b[55] ), .B(\a[55] ), .Y(new_n711_));
  AND2X1   g326(.A(\b[55] ), .B(\a[55] ), .Y(new_n712_));
  OR2X1    g327(.A(new_n712_), .B(new_n711_), .Y(new_n713_));
  XOR2X1   g328(.A(new_n713_), .B(new_n710_), .Y(\f[55] ));
  INVX1    g329(.A(new_n712_), .Y(new_n715_));
  OAI21X1  g330(.A0(new_n711_), .A1(new_n710_), .B0(new_n715_), .Y(new_n716_));
  XOR2X1   g331(.A(\b[56] ), .B(\a[56] ), .Y(new_n717_));
  XOR2X1   g332(.A(new_n717_), .B(new_n716_), .Y(\f[56] ));
  NOR2X1   g333(.A(\b[56] ), .B(\a[56] ), .Y(new_n719_));
  INVX1    g334(.A(new_n719_), .Y(new_n720_));
  AND2X1   g335(.A(\b[56] ), .B(\a[56] ), .Y(new_n721_));
  AOI21X1  g336(.A0(new_n720_), .A1(new_n716_), .B0(new_n721_), .Y(new_n722_));
  NOR2X1   g337(.A(\b[57] ), .B(\a[57] ), .Y(new_n723_));
  AND2X1   g338(.A(\b[57] ), .B(\a[57] ), .Y(new_n724_));
  OR2X1    g339(.A(new_n724_), .B(new_n723_), .Y(new_n725_));
  XOR2X1   g340(.A(new_n725_), .B(new_n722_), .Y(\f[57] ));
  INVX1    g341(.A(new_n724_), .Y(new_n727_));
  OAI21X1  g342(.A0(new_n723_), .A1(new_n722_), .B0(new_n727_), .Y(new_n728_));
  XOR2X1   g343(.A(\b[58] ), .B(\a[58] ), .Y(new_n729_));
  XOR2X1   g344(.A(new_n729_), .B(new_n728_), .Y(\f[58] ));
  NOR2X1   g345(.A(\b[58] ), .B(\a[58] ), .Y(new_n731_));
  INVX1    g346(.A(new_n731_), .Y(new_n732_));
  AND2X1   g347(.A(\b[58] ), .B(\a[58] ), .Y(new_n733_));
  AOI21X1  g348(.A0(new_n732_), .A1(new_n728_), .B0(new_n733_), .Y(new_n734_));
  NOR2X1   g349(.A(\b[59] ), .B(\a[59] ), .Y(new_n735_));
  AND2X1   g350(.A(\b[59] ), .B(\a[59] ), .Y(new_n736_));
  OR2X1    g351(.A(new_n736_), .B(new_n735_), .Y(new_n737_));
  XOR2X1   g352(.A(new_n737_), .B(new_n734_), .Y(\f[59] ));
  INVX1    g353(.A(new_n736_), .Y(new_n739_));
  OAI21X1  g354(.A0(new_n735_), .A1(new_n734_), .B0(new_n739_), .Y(new_n740_));
  XOR2X1   g355(.A(\b[60] ), .B(\a[60] ), .Y(new_n741_));
  XOR2X1   g356(.A(new_n741_), .B(new_n740_), .Y(\f[60] ));
  NOR2X1   g357(.A(\b[60] ), .B(\a[60] ), .Y(new_n743_));
  INVX1    g358(.A(new_n743_), .Y(new_n744_));
  AND2X1   g359(.A(\b[60] ), .B(\a[60] ), .Y(new_n745_));
  AOI21X1  g360(.A0(new_n744_), .A1(new_n740_), .B0(new_n745_), .Y(new_n746_));
  NOR2X1   g361(.A(\b[61] ), .B(\a[61] ), .Y(new_n747_));
  AND2X1   g362(.A(\b[61] ), .B(\a[61] ), .Y(new_n748_));
  OR2X1    g363(.A(new_n748_), .B(new_n747_), .Y(new_n749_));
  XOR2X1   g364(.A(new_n749_), .B(new_n746_), .Y(\f[61] ));
  INVX1    g365(.A(new_n748_), .Y(new_n751_));
  OAI21X1  g366(.A0(new_n747_), .A1(new_n746_), .B0(new_n751_), .Y(new_n752_));
  XOR2X1   g367(.A(\b[62] ), .B(\a[62] ), .Y(new_n753_));
  XOR2X1   g368(.A(new_n753_), .B(new_n752_), .Y(\f[62] ));
  NOR2X1   g369(.A(\b[62] ), .B(\a[62] ), .Y(new_n755_));
  INVX1    g370(.A(new_n755_), .Y(new_n756_));
  AND2X1   g371(.A(\b[62] ), .B(\a[62] ), .Y(new_n757_));
  AOI21X1  g372(.A0(new_n756_), .A1(new_n752_), .B0(new_n757_), .Y(new_n758_));
  NOR2X1   g373(.A(\b[63] ), .B(\a[63] ), .Y(new_n759_));
  AND2X1   g374(.A(\b[63] ), .B(\a[63] ), .Y(new_n760_));
  OR2X1    g375(.A(new_n760_), .B(new_n759_), .Y(new_n761_));
  XOR2X1   g376(.A(new_n761_), .B(new_n758_), .Y(\f[63] ));
  INVX1    g377(.A(new_n760_), .Y(new_n763_));
  OAI21X1  g378(.A0(new_n759_), .A1(new_n758_), .B0(new_n763_), .Y(new_n764_));
  XOR2X1   g379(.A(\b[64] ), .B(\a[64] ), .Y(new_n765_));
  XOR2X1   g380(.A(new_n765_), .B(new_n764_), .Y(\f[64] ));
  NOR2X1   g381(.A(\b[64] ), .B(\a[64] ), .Y(new_n767_));
  INVX1    g382(.A(new_n767_), .Y(new_n768_));
  AND2X1   g383(.A(\b[64] ), .B(\a[64] ), .Y(new_n769_));
  AOI21X1  g384(.A0(new_n768_), .A1(new_n764_), .B0(new_n769_), .Y(new_n770_));
  NOR2X1   g385(.A(\b[65] ), .B(\a[65] ), .Y(new_n771_));
  AND2X1   g386(.A(\b[65] ), .B(\a[65] ), .Y(new_n772_));
  OR2X1    g387(.A(new_n772_), .B(new_n771_), .Y(new_n773_));
  XOR2X1   g388(.A(new_n773_), .B(new_n770_), .Y(\f[65] ));
  INVX1    g389(.A(new_n772_), .Y(new_n775_));
  OAI21X1  g390(.A0(new_n771_), .A1(new_n770_), .B0(new_n775_), .Y(new_n776_));
  XOR2X1   g391(.A(\b[66] ), .B(\a[66] ), .Y(new_n777_));
  XOR2X1   g392(.A(new_n777_), .B(new_n776_), .Y(\f[66] ));
  NOR2X1   g393(.A(\b[66] ), .B(\a[66] ), .Y(new_n779_));
  INVX1    g394(.A(new_n779_), .Y(new_n780_));
  AND2X1   g395(.A(\b[66] ), .B(\a[66] ), .Y(new_n781_));
  AOI21X1  g396(.A0(new_n780_), .A1(new_n776_), .B0(new_n781_), .Y(new_n782_));
  NOR2X1   g397(.A(\b[67] ), .B(\a[67] ), .Y(new_n783_));
  AND2X1   g398(.A(\b[67] ), .B(\a[67] ), .Y(new_n784_));
  OR2X1    g399(.A(new_n784_), .B(new_n783_), .Y(new_n785_));
  XOR2X1   g400(.A(new_n785_), .B(new_n782_), .Y(\f[67] ));
  INVX1    g401(.A(new_n784_), .Y(new_n787_));
  OAI21X1  g402(.A0(new_n783_), .A1(new_n782_), .B0(new_n787_), .Y(new_n788_));
  XOR2X1   g403(.A(\b[68] ), .B(\a[68] ), .Y(new_n789_));
  XOR2X1   g404(.A(new_n789_), .B(new_n788_), .Y(\f[68] ));
  NOR2X1   g405(.A(\b[68] ), .B(\a[68] ), .Y(new_n791_));
  INVX1    g406(.A(new_n791_), .Y(new_n792_));
  AND2X1   g407(.A(\b[68] ), .B(\a[68] ), .Y(new_n793_));
  AOI21X1  g408(.A0(new_n792_), .A1(new_n788_), .B0(new_n793_), .Y(new_n794_));
  NOR2X1   g409(.A(\b[69] ), .B(\a[69] ), .Y(new_n795_));
  AND2X1   g410(.A(\b[69] ), .B(\a[69] ), .Y(new_n796_));
  OR2X1    g411(.A(new_n796_), .B(new_n795_), .Y(new_n797_));
  XOR2X1   g412(.A(new_n797_), .B(new_n794_), .Y(\f[69] ));
  INVX1    g413(.A(new_n796_), .Y(new_n799_));
  OAI21X1  g414(.A0(new_n795_), .A1(new_n794_), .B0(new_n799_), .Y(new_n800_));
  XOR2X1   g415(.A(\b[70] ), .B(\a[70] ), .Y(new_n801_));
  XOR2X1   g416(.A(new_n801_), .B(new_n800_), .Y(\f[70] ));
  NOR2X1   g417(.A(\b[70] ), .B(\a[70] ), .Y(new_n803_));
  INVX1    g418(.A(new_n803_), .Y(new_n804_));
  AND2X1   g419(.A(\b[70] ), .B(\a[70] ), .Y(new_n805_));
  AOI21X1  g420(.A0(new_n804_), .A1(new_n800_), .B0(new_n805_), .Y(new_n806_));
  NOR2X1   g421(.A(\b[71] ), .B(\a[71] ), .Y(new_n807_));
  AND2X1   g422(.A(\b[71] ), .B(\a[71] ), .Y(new_n808_));
  OR2X1    g423(.A(new_n808_), .B(new_n807_), .Y(new_n809_));
  XOR2X1   g424(.A(new_n809_), .B(new_n806_), .Y(\f[71] ));
  INVX1    g425(.A(new_n808_), .Y(new_n811_));
  OAI21X1  g426(.A0(new_n807_), .A1(new_n806_), .B0(new_n811_), .Y(new_n812_));
  XOR2X1   g427(.A(\b[72] ), .B(\a[72] ), .Y(new_n813_));
  XOR2X1   g428(.A(new_n813_), .B(new_n812_), .Y(\f[72] ));
  NOR2X1   g429(.A(\b[72] ), .B(\a[72] ), .Y(new_n815_));
  INVX1    g430(.A(new_n815_), .Y(new_n816_));
  AND2X1   g431(.A(\b[72] ), .B(\a[72] ), .Y(new_n817_));
  AOI21X1  g432(.A0(new_n816_), .A1(new_n812_), .B0(new_n817_), .Y(new_n818_));
  NOR2X1   g433(.A(\b[73] ), .B(\a[73] ), .Y(new_n819_));
  AND2X1   g434(.A(\b[73] ), .B(\a[73] ), .Y(new_n820_));
  OR2X1    g435(.A(new_n820_), .B(new_n819_), .Y(new_n821_));
  XOR2X1   g436(.A(new_n821_), .B(new_n818_), .Y(\f[73] ));
  INVX1    g437(.A(new_n820_), .Y(new_n823_));
  OAI21X1  g438(.A0(new_n819_), .A1(new_n818_), .B0(new_n823_), .Y(new_n824_));
  XOR2X1   g439(.A(\b[74] ), .B(\a[74] ), .Y(new_n825_));
  XOR2X1   g440(.A(new_n825_), .B(new_n824_), .Y(\f[74] ));
  NOR2X1   g441(.A(\b[74] ), .B(\a[74] ), .Y(new_n827_));
  INVX1    g442(.A(new_n827_), .Y(new_n828_));
  AND2X1   g443(.A(\b[74] ), .B(\a[74] ), .Y(new_n829_));
  AOI21X1  g444(.A0(new_n828_), .A1(new_n824_), .B0(new_n829_), .Y(new_n830_));
  NOR2X1   g445(.A(\b[75] ), .B(\a[75] ), .Y(new_n831_));
  AND2X1   g446(.A(\b[75] ), .B(\a[75] ), .Y(new_n832_));
  OR2X1    g447(.A(new_n832_), .B(new_n831_), .Y(new_n833_));
  XOR2X1   g448(.A(new_n833_), .B(new_n830_), .Y(\f[75] ));
  INVX1    g449(.A(new_n832_), .Y(new_n835_));
  OAI21X1  g450(.A0(new_n831_), .A1(new_n830_), .B0(new_n835_), .Y(new_n836_));
  XOR2X1   g451(.A(\b[76] ), .B(\a[76] ), .Y(new_n837_));
  XOR2X1   g452(.A(new_n837_), .B(new_n836_), .Y(\f[76] ));
  NOR2X1   g453(.A(\b[76] ), .B(\a[76] ), .Y(new_n839_));
  INVX1    g454(.A(new_n839_), .Y(new_n840_));
  AND2X1   g455(.A(\b[76] ), .B(\a[76] ), .Y(new_n841_));
  AOI21X1  g456(.A0(new_n840_), .A1(new_n836_), .B0(new_n841_), .Y(new_n842_));
  NOR2X1   g457(.A(\b[77] ), .B(\a[77] ), .Y(new_n843_));
  AND2X1   g458(.A(\b[77] ), .B(\a[77] ), .Y(new_n844_));
  OR2X1    g459(.A(new_n844_), .B(new_n843_), .Y(new_n845_));
  XOR2X1   g460(.A(new_n845_), .B(new_n842_), .Y(\f[77] ));
  INVX1    g461(.A(new_n844_), .Y(new_n847_));
  OAI21X1  g462(.A0(new_n843_), .A1(new_n842_), .B0(new_n847_), .Y(new_n848_));
  XOR2X1   g463(.A(\b[78] ), .B(\a[78] ), .Y(new_n849_));
  XOR2X1   g464(.A(new_n849_), .B(new_n848_), .Y(\f[78] ));
  NOR2X1   g465(.A(\b[78] ), .B(\a[78] ), .Y(new_n851_));
  INVX1    g466(.A(new_n851_), .Y(new_n852_));
  AND2X1   g467(.A(\b[78] ), .B(\a[78] ), .Y(new_n853_));
  AOI21X1  g468(.A0(new_n852_), .A1(new_n848_), .B0(new_n853_), .Y(new_n854_));
  NOR2X1   g469(.A(\b[79] ), .B(\a[79] ), .Y(new_n855_));
  AND2X1   g470(.A(\b[79] ), .B(\a[79] ), .Y(new_n856_));
  OR2X1    g471(.A(new_n856_), .B(new_n855_), .Y(new_n857_));
  XOR2X1   g472(.A(new_n857_), .B(new_n854_), .Y(\f[79] ));
  INVX1    g473(.A(new_n856_), .Y(new_n859_));
  OAI21X1  g474(.A0(new_n855_), .A1(new_n854_), .B0(new_n859_), .Y(new_n860_));
  XOR2X1   g475(.A(\b[80] ), .B(\a[80] ), .Y(new_n861_));
  XOR2X1   g476(.A(new_n861_), .B(new_n860_), .Y(\f[80] ));
  NOR2X1   g477(.A(\b[80] ), .B(\a[80] ), .Y(new_n863_));
  INVX1    g478(.A(new_n863_), .Y(new_n864_));
  AND2X1   g479(.A(\b[80] ), .B(\a[80] ), .Y(new_n865_));
  AOI21X1  g480(.A0(new_n864_), .A1(new_n860_), .B0(new_n865_), .Y(new_n866_));
  NOR2X1   g481(.A(\b[81] ), .B(\a[81] ), .Y(new_n867_));
  AND2X1   g482(.A(\b[81] ), .B(\a[81] ), .Y(new_n868_));
  OR2X1    g483(.A(new_n868_), .B(new_n867_), .Y(new_n869_));
  XOR2X1   g484(.A(new_n869_), .B(new_n866_), .Y(\f[81] ));
  INVX1    g485(.A(new_n868_), .Y(new_n871_));
  OAI21X1  g486(.A0(new_n867_), .A1(new_n866_), .B0(new_n871_), .Y(new_n872_));
  XOR2X1   g487(.A(\b[82] ), .B(\a[82] ), .Y(new_n873_));
  XOR2X1   g488(.A(new_n873_), .B(new_n872_), .Y(\f[82] ));
  NOR2X1   g489(.A(\b[82] ), .B(\a[82] ), .Y(new_n875_));
  INVX1    g490(.A(new_n875_), .Y(new_n876_));
  AND2X1   g491(.A(\b[82] ), .B(\a[82] ), .Y(new_n877_));
  AOI21X1  g492(.A0(new_n876_), .A1(new_n872_), .B0(new_n877_), .Y(new_n878_));
  NOR2X1   g493(.A(\b[83] ), .B(\a[83] ), .Y(new_n879_));
  AND2X1   g494(.A(\b[83] ), .B(\a[83] ), .Y(new_n880_));
  OR2X1    g495(.A(new_n880_), .B(new_n879_), .Y(new_n881_));
  XOR2X1   g496(.A(new_n881_), .B(new_n878_), .Y(\f[83] ));
  INVX1    g497(.A(new_n880_), .Y(new_n883_));
  OAI21X1  g498(.A0(new_n879_), .A1(new_n878_), .B0(new_n883_), .Y(new_n884_));
  XOR2X1   g499(.A(\b[84] ), .B(\a[84] ), .Y(new_n885_));
  XOR2X1   g500(.A(new_n885_), .B(new_n884_), .Y(\f[84] ));
  NOR2X1   g501(.A(\b[84] ), .B(\a[84] ), .Y(new_n887_));
  INVX1    g502(.A(new_n887_), .Y(new_n888_));
  AND2X1   g503(.A(\b[84] ), .B(\a[84] ), .Y(new_n889_));
  AOI21X1  g504(.A0(new_n888_), .A1(new_n884_), .B0(new_n889_), .Y(new_n890_));
  NOR2X1   g505(.A(\b[85] ), .B(\a[85] ), .Y(new_n891_));
  AND2X1   g506(.A(\b[85] ), .B(\a[85] ), .Y(new_n892_));
  OR2X1    g507(.A(new_n892_), .B(new_n891_), .Y(new_n893_));
  XOR2X1   g508(.A(new_n893_), .B(new_n890_), .Y(\f[85] ));
  INVX1    g509(.A(new_n892_), .Y(new_n895_));
  OAI21X1  g510(.A0(new_n891_), .A1(new_n890_), .B0(new_n895_), .Y(new_n896_));
  XOR2X1   g511(.A(\b[86] ), .B(\a[86] ), .Y(new_n897_));
  XOR2X1   g512(.A(new_n897_), .B(new_n896_), .Y(\f[86] ));
  NOR2X1   g513(.A(\b[86] ), .B(\a[86] ), .Y(new_n899_));
  INVX1    g514(.A(new_n899_), .Y(new_n900_));
  AND2X1   g515(.A(\b[86] ), .B(\a[86] ), .Y(new_n901_));
  AOI21X1  g516(.A0(new_n900_), .A1(new_n896_), .B0(new_n901_), .Y(new_n902_));
  NOR2X1   g517(.A(\b[87] ), .B(\a[87] ), .Y(new_n903_));
  AND2X1   g518(.A(\b[87] ), .B(\a[87] ), .Y(new_n904_));
  OR2X1    g519(.A(new_n904_), .B(new_n903_), .Y(new_n905_));
  XOR2X1   g520(.A(new_n905_), .B(new_n902_), .Y(\f[87] ));
  INVX1    g521(.A(new_n904_), .Y(new_n907_));
  OAI21X1  g522(.A0(new_n903_), .A1(new_n902_), .B0(new_n907_), .Y(new_n908_));
  XOR2X1   g523(.A(\b[88] ), .B(\a[88] ), .Y(new_n909_));
  XOR2X1   g524(.A(new_n909_), .B(new_n908_), .Y(\f[88] ));
  NOR2X1   g525(.A(\b[88] ), .B(\a[88] ), .Y(new_n911_));
  INVX1    g526(.A(new_n911_), .Y(new_n912_));
  AND2X1   g527(.A(\b[88] ), .B(\a[88] ), .Y(new_n913_));
  AOI21X1  g528(.A0(new_n912_), .A1(new_n908_), .B0(new_n913_), .Y(new_n914_));
  NOR2X1   g529(.A(\b[89] ), .B(\a[89] ), .Y(new_n915_));
  AND2X1   g530(.A(\b[89] ), .B(\a[89] ), .Y(new_n916_));
  OR2X1    g531(.A(new_n916_), .B(new_n915_), .Y(new_n917_));
  XOR2X1   g532(.A(new_n917_), .B(new_n914_), .Y(\f[89] ));
  INVX1    g533(.A(new_n916_), .Y(new_n919_));
  OAI21X1  g534(.A0(new_n915_), .A1(new_n914_), .B0(new_n919_), .Y(new_n920_));
  XOR2X1   g535(.A(\b[90] ), .B(\a[90] ), .Y(new_n921_));
  XOR2X1   g536(.A(new_n921_), .B(new_n920_), .Y(\f[90] ));
  NOR2X1   g537(.A(\b[90] ), .B(\a[90] ), .Y(new_n923_));
  INVX1    g538(.A(new_n923_), .Y(new_n924_));
  AND2X1   g539(.A(\b[90] ), .B(\a[90] ), .Y(new_n925_));
  AOI21X1  g540(.A0(new_n924_), .A1(new_n920_), .B0(new_n925_), .Y(new_n926_));
  NOR2X1   g541(.A(\b[91] ), .B(\a[91] ), .Y(new_n927_));
  AND2X1   g542(.A(\b[91] ), .B(\a[91] ), .Y(new_n928_));
  OR2X1    g543(.A(new_n928_), .B(new_n927_), .Y(new_n929_));
  XOR2X1   g544(.A(new_n929_), .B(new_n926_), .Y(\f[91] ));
  INVX1    g545(.A(new_n928_), .Y(new_n931_));
  OAI21X1  g546(.A0(new_n927_), .A1(new_n926_), .B0(new_n931_), .Y(new_n932_));
  XOR2X1   g547(.A(\b[92] ), .B(\a[92] ), .Y(new_n933_));
  XOR2X1   g548(.A(new_n933_), .B(new_n932_), .Y(\f[92] ));
  NOR2X1   g549(.A(\b[92] ), .B(\a[92] ), .Y(new_n935_));
  INVX1    g550(.A(new_n935_), .Y(new_n936_));
  AND2X1   g551(.A(\b[92] ), .B(\a[92] ), .Y(new_n937_));
  AOI21X1  g552(.A0(new_n936_), .A1(new_n932_), .B0(new_n937_), .Y(new_n938_));
  NOR2X1   g553(.A(\b[93] ), .B(\a[93] ), .Y(new_n939_));
  AND2X1   g554(.A(\b[93] ), .B(\a[93] ), .Y(new_n940_));
  OR2X1    g555(.A(new_n940_), .B(new_n939_), .Y(new_n941_));
  XOR2X1   g556(.A(new_n941_), .B(new_n938_), .Y(\f[93] ));
  INVX1    g557(.A(new_n940_), .Y(new_n943_));
  OAI21X1  g558(.A0(new_n939_), .A1(new_n938_), .B0(new_n943_), .Y(new_n944_));
  XOR2X1   g559(.A(\b[94] ), .B(\a[94] ), .Y(new_n945_));
  XOR2X1   g560(.A(new_n945_), .B(new_n944_), .Y(\f[94] ));
  NOR2X1   g561(.A(\b[94] ), .B(\a[94] ), .Y(new_n947_));
  INVX1    g562(.A(new_n947_), .Y(new_n948_));
  AND2X1   g563(.A(\b[94] ), .B(\a[94] ), .Y(new_n949_));
  AOI21X1  g564(.A0(new_n948_), .A1(new_n944_), .B0(new_n949_), .Y(new_n950_));
  NOR2X1   g565(.A(\b[95] ), .B(\a[95] ), .Y(new_n951_));
  AND2X1   g566(.A(\b[95] ), .B(\a[95] ), .Y(new_n952_));
  OR2X1    g567(.A(new_n952_), .B(new_n951_), .Y(new_n953_));
  XOR2X1   g568(.A(new_n953_), .B(new_n950_), .Y(\f[95] ));
  INVX1    g569(.A(new_n952_), .Y(new_n955_));
  OAI21X1  g570(.A0(new_n951_), .A1(new_n950_), .B0(new_n955_), .Y(new_n956_));
  XOR2X1   g571(.A(\b[96] ), .B(\a[96] ), .Y(new_n957_));
  XOR2X1   g572(.A(new_n957_), .B(new_n956_), .Y(\f[96] ));
  NOR2X1   g573(.A(\b[96] ), .B(\a[96] ), .Y(new_n959_));
  INVX1    g574(.A(new_n959_), .Y(new_n960_));
  AND2X1   g575(.A(\b[96] ), .B(\a[96] ), .Y(new_n961_));
  AOI21X1  g576(.A0(new_n960_), .A1(new_n956_), .B0(new_n961_), .Y(new_n962_));
  NOR2X1   g577(.A(\b[97] ), .B(\a[97] ), .Y(new_n963_));
  AND2X1   g578(.A(\b[97] ), .B(\a[97] ), .Y(new_n964_));
  OR2X1    g579(.A(new_n964_), .B(new_n963_), .Y(new_n965_));
  XOR2X1   g580(.A(new_n965_), .B(new_n962_), .Y(\f[97] ));
  INVX1    g581(.A(new_n964_), .Y(new_n967_));
  OAI21X1  g582(.A0(new_n963_), .A1(new_n962_), .B0(new_n967_), .Y(new_n968_));
  XOR2X1   g583(.A(\b[98] ), .B(\a[98] ), .Y(new_n969_));
  XOR2X1   g584(.A(new_n969_), .B(new_n968_), .Y(\f[98] ));
  NOR2X1   g585(.A(\b[98] ), .B(\a[98] ), .Y(new_n971_));
  INVX1    g586(.A(new_n971_), .Y(new_n972_));
  AND2X1   g587(.A(\b[98] ), .B(\a[98] ), .Y(new_n973_));
  AOI21X1  g588(.A0(new_n972_), .A1(new_n968_), .B0(new_n973_), .Y(new_n974_));
  NOR2X1   g589(.A(\b[99] ), .B(\a[99] ), .Y(new_n975_));
  AND2X1   g590(.A(\b[99] ), .B(\a[99] ), .Y(new_n976_));
  OR2X1    g591(.A(new_n976_), .B(new_n975_), .Y(new_n977_));
  XOR2X1   g592(.A(new_n977_), .B(new_n974_), .Y(\f[99] ));
  INVX1    g593(.A(new_n976_), .Y(new_n979_));
  OAI21X1  g594(.A0(new_n975_), .A1(new_n974_), .B0(new_n979_), .Y(new_n980_));
  XOR2X1   g595(.A(\b[100] ), .B(\a[100] ), .Y(new_n981_));
  XOR2X1   g596(.A(new_n981_), .B(new_n980_), .Y(\f[100] ));
  NOR2X1   g597(.A(\b[100] ), .B(\a[100] ), .Y(new_n983_));
  INVX1    g598(.A(new_n983_), .Y(new_n984_));
  AND2X1   g599(.A(\b[100] ), .B(\a[100] ), .Y(new_n985_));
  AOI21X1  g600(.A0(new_n984_), .A1(new_n980_), .B0(new_n985_), .Y(new_n986_));
  NOR2X1   g601(.A(\b[101] ), .B(\a[101] ), .Y(new_n987_));
  AND2X1   g602(.A(\b[101] ), .B(\a[101] ), .Y(new_n988_));
  OR2X1    g603(.A(new_n988_), .B(new_n987_), .Y(new_n989_));
  XOR2X1   g604(.A(new_n989_), .B(new_n986_), .Y(\f[101] ));
  INVX1    g605(.A(new_n988_), .Y(new_n991_));
  OAI21X1  g606(.A0(new_n987_), .A1(new_n986_), .B0(new_n991_), .Y(new_n992_));
  XOR2X1   g607(.A(\b[102] ), .B(\a[102] ), .Y(new_n993_));
  XOR2X1   g608(.A(new_n993_), .B(new_n992_), .Y(\f[102] ));
  NOR2X1   g609(.A(\b[102] ), .B(\a[102] ), .Y(new_n995_));
  INVX1    g610(.A(new_n995_), .Y(new_n996_));
  AND2X1   g611(.A(\b[102] ), .B(\a[102] ), .Y(new_n997_));
  AOI21X1  g612(.A0(new_n996_), .A1(new_n992_), .B0(new_n997_), .Y(new_n998_));
  NOR2X1   g613(.A(\b[103] ), .B(\a[103] ), .Y(new_n999_));
  AND2X1   g614(.A(\b[103] ), .B(\a[103] ), .Y(new_n1000_));
  OR2X1    g615(.A(new_n1000_), .B(new_n999_), .Y(new_n1001_));
  XOR2X1   g616(.A(new_n1001_), .B(new_n998_), .Y(\f[103] ));
  INVX1    g617(.A(new_n1000_), .Y(new_n1003_));
  OAI21X1  g618(.A0(new_n999_), .A1(new_n998_), .B0(new_n1003_), .Y(new_n1004_));
  XOR2X1   g619(.A(\b[104] ), .B(\a[104] ), .Y(new_n1005_));
  XOR2X1   g620(.A(new_n1005_), .B(new_n1004_), .Y(\f[104] ));
  NOR2X1   g621(.A(\b[104] ), .B(\a[104] ), .Y(new_n1007_));
  INVX1    g622(.A(new_n1007_), .Y(new_n1008_));
  AND2X1   g623(.A(\b[104] ), .B(\a[104] ), .Y(new_n1009_));
  AOI21X1  g624(.A0(new_n1008_), .A1(new_n1004_), .B0(new_n1009_), .Y(new_n1010_));
  NOR2X1   g625(.A(\b[105] ), .B(\a[105] ), .Y(new_n1011_));
  AND2X1   g626(.A(\b[105] ), .B(\a[105] ), .Y(new_n1012_));
  OR2X1    g627(.A(new_n1012_), .B(new_n1011_), .Y(new_n1013_));
  XOR2X1   g628(.A(new_n1013_), .B(new_n1010_), .Y(\f[105] ));
  INVX1    g629(.A(new_n1012_), .Y(new_n1015_));
  OAI21X1  g630(.A0(new_n1011_), .A1(new_n1010_), .B0(new_n1015_), .Y(new_n1016_));
  XOR2X1   g631(.A(\b[106] ), .B(\a[106] ), .Y(new_n1017_));
  XOR2X1   g632(.A(new_n1017_), .B(new_n1016_), .Y(\f[106] ));
  NOR2X1   g633(.A(\b[106] ), .B(\a[106] ), .Y(new_n1019_));
  INVX1    g634(.A(new_n1019_), .Y(new_n1020_));
  AND2X1   g635(.A(\b[106] ), .B(\a[106] ), .Y(new_n1021_));
  AOI21X1  g636(.A0(new_n1020_), .A1(new_n1016_), .B0(new_n1021_), .Y(new_n1022_));
  NOR2X1   g637(.A(\b[107] ), .B(\a[107] ), .Y(new_n1023_));
  AND2X1   g638(.A(\b[107] ), .B(\a[107] ), .Y(new_n1024_));
  OR2X1    g639(.A(new_n1024_), .B(new_n1023_), .Y(new_n1025_));
  XOR2X1   g640(.A(new_n1025_), .B(new_n1022_), .Y(\f[107] ));
  INVX1    g641(.A(new_n1024_), .Y(new_n1027_));
  OAI21X1  g642(.A0(new_n1023_), .A1(new_n1022_), .B0(new_n1027_), .Y(new_n1028_));
  XOR2X1   g643(.A(\b[108] ), .B(\a[108] ), .Y(new_n1029_));
  XOR2X1   g644(.A(new_n1029_), .B(new_n1028_), .Y(\f[108] ));
  NOR2X1   g645(.A(\b[108] ), .B(\a[108] ), .Y(new_n1031_));
  INVX1    g646(.A(new_n1031_), .Y(new_n1032_));
  AND2X1   g647(.A(\b[108] ), .B(\a[108] ), .Y(new_n1033_));
  AOI21X1  g648(.A0(new_n1032_), .A1(new_n1028_), .B0(new_n1033_), .Y(new_n1034_));
  NOR2X1   g649(.A(\b[109] ), .B(\a[109] ), .Y(new_n1035_));
  AND2X1   g650(.A(\b[109] ), .B(\a[109] ), .Y(new_n1036_));
  OR2X1    g651(.A(new_n1036_), .B(new_n1035_), .Y(new_n1037_));
  XOR2X1   g652(.A(new_n1037_), .B(new_n1034_), .Y(\f[109] ));
  INVX1    g653(.A(new_n1036_), .Y(new_n1039_));
  OAI21X1  g654(.A0(new_n1035_), .A1(new_n1034_), .B0(new_n1039_), .Y(new_n1040_));
  XOR2X1   g655(.A(\b[110] ), .B(\a[110] ), .Y(new_n1041_));
  XOR2X1   g656(.A(new_n1041_), .B(new_n1040_), .Y(\f[110] ));
  NOR2X1   g657(.A(\b[110] ), .B(\a[110] ), .Y(new_n1043_));
  INVX1    g658(.A(new_n1043_), .Y(new_n1044_));
  AND2X1   g659(.A(\b[110] ), .B(\a[110] ), .Y(new_n1045_));
  AOI21X1  g660(.A0(new_n1044_), .A1(new_n1040_), .B0(new_n1045_), .Y(new_n1046_));
  NOR2X1   g661(.A(\b[111] ), .B(\a[111] ), .Y(new_n1047_));
  AND2X1   g662(.A(\b[111] ), .B(\a[111] ), .Y(new_n1048_));
  OR2X1    g663(.A(new_n1048_), .B(new_n1047_), .Y(new_n1049_));
  XOR2X1   g664(.A(new_n1049_), .B(new_n1046_), .Y(\f[111] ));
  INVX1    g665(.A(new_n1048_), .Y(new_n1051_));
  OAI21X1  g666(.A0(new_n1047_), .A1(new_n1046_), .B0(new_n1051_), .Y(new_n1052_));
  XOR2X1   g667(.A(\b[112] ), .B(\a[112] ), .Y(new_n1053_));
  XOR2X1   g668(.A(new_n1053_), .B(new_n1052_), .Y(\f[112] ));
  NOR2X1   g669(.A(\b[112] ), .B(\a[112] ), .Y(new_n1055_));
  INVX1    g670(.A(new_n1055_), .Y(new_n1056_));
  AND2X1   g671(.A(\b[112] ), .B(\a[112] ), .Y(new_n1057_));
  AOI21X1  g672(.A0(new_n1056_), .A1(new_n1052_), .B0(new_n1057_), .Y(new_n1058_));
  NOR2X1   g673(.A(\b[113] ), .B(\a[113] ), .Y(new_n1059_));
  AND2X1   g674(.A(\b[113] ), .B(\a[113] ), .Y(new_n1060_));
  OR2X1    g675(.A(new_n1060_), .B(new_n1059_), .Y(new_n1061_));
  XOR2X1   g676(.A(new_n1061_), .B(new_n1058_), .Y(\f[113] ));
  INVX1    g677(.A(new_n1060_), .Y(new_n1063_));
  OAI21X1  g678(.A0(new_n1059_), .A1(new_n1058_), .B0(new_n1063_), .Y(new_n1064_));
  XOR2X1   g679(.A(\b[114] ), .B(\a[114] ), .Y(new_n1065_));
  XOR2X1   g680(.A(new_n1065_), .B(new_n1064_), .Y(\f[114] ));
  NOR2X1   g681(.A(\b[114] ), .B(\a[114] ), .Y(new_n1067_));
  INVX1    g682(.A(new_n1067_), .Y(new_n1068_));
  AND2X1   g683(.A(\b[114] ), .B(\a[114] ), .Y(new_n1069_));
  AOI21X1  g684(.A0(new_n1068_), .A1(new_n1064_), .B0(new_n1069_), .Y(new_n1070_));
  NOR2X1   g685(.A(\b[115] ), .B(\a[115] ), .Y(new_n1071_));
  AND2X1   g686(.A(\b[115] ), .B(\a[115] ), .Y(new_n1072_));
  OR2X1    g687(.A(new_n1072_), .B(new_n1071_), .Y(new_n1073_));
  XOR2X1   g688(.A(new_n1073_), .B(new_n1070_), .Y(\f[115] ));
  INVX1    g689(.A(new_n1072_), .Y(new_n1075_));
  OAI21X1  g690(.A0(new_n1071_), .A1(new_n1070_), .B0(new_n1075_), .Y(new_n1076_));
  XOR2X1   g691(.A(\b[116] ), .B(\a[116] ), .Y(new_n1077_));
  XOR2X1   g692(.A(new_n1077_), .B(new_n1076_), .Y(\f[116] ));
  NOR2X1   g693(.A(\b[116] ), .B(\a[116] ), .Y(new_n1079_));
  INVX1    g694(.A(new_n1079_), .Y(new_n1080_));
  AND2X1   g695(.A(\b[116] ), .B(\a[116] ), .Y(new_n1081_));
  AOI21X1  g696(.A0(new_n1080_), .A1(new_n1076_), .B0(new_n1081_), .Y(new_n1082_));
  NOR2X1   g697(.A(\b[117] ), .B(\a[117] ), .Y(new_n1083_));
  AND2X1   g698(.A(\b[117] ), .B(\a[117] ), .Y(new_n1084_));
  OR2X1    g699(.A(new_n1084_), .B(new_n1083_), .Y(new_n1085_));
  XOR2X1   g700(.A(new_n1085_), .B(new_n1082_), .Y(\f[117] ));
  INVX1    g701(.A(new_n1084_), .Y(new_n1087_));
  OAI21X1  g702(.A0(new_n1083_), .A1(new_n1082_), .B0(new_n1087_), .Y(new_n1088_));
  XOR2X1   g703(.A(\b[118] ), .B(\a[118] ), .Y(new_n1089_));
  XOR2X1   g704(.A(new_n1089_), .B(new_n1088_), .Y(\f[118] ));
  NOR2X1   g705(.A(\b[118] ), .B(\a[118] ), .Y(new_n1091_));
  INVX1    g706(.A(new_n1091_), .Y(new_n1092_));
  AND2X1   g707(.A(\b[118] ), .B(\a[118] ), .Y(new_n1093_));
  AOI21X1  g708(.A0(new_n1092_), .A1(new_n1088_), .B0(new_n1093_), .Y(new_n1094_));
  NOR2X1   g709(.A(\b[119] ), .B(\a[119] ), .Y(new_n1095_));
  AND2X1   g710(.A(\b[119] ), .B(\a[119] ), .Y(new_n1096_));
  OR2X1    g711(.A(new_n1096_), .B(new_n1095_), .Y(new_n1097_));
  XOR2X1   g712(.A(new_n1097_), .B(new_n1094_), .Y(\f[119] ));
  INVX1    g713(.A(new_n1096_), .Y(new_n1099_));
  OAI21X1  g714(.A0(new_n1095_), .A1(new_n1094_), .B0(new_n1099_), .Y(new_n1100_));
  XOR2X1   g715(.A(\b[120] ), .B(\a[120] ), .Y(new_n1101_));
  XOR2X1   g716(.A(new_n1101_), .B(new_n1100_), .Y(\f[120] ));
  NOR2X1   g717(.A(\b[120] ), .B(\a[120] ), .Y(new_n1103_));
  INVX1    g718(.A(new_n1103_), .Y(new_n1104_));
  AND2X1   g719(.A(\b[120] ), .B(\a[120] ), .Y(new_n1105_));
  AOI21X1  g720(.A0(new_n1104_), .A1(new_n1100_), .B0(new_n1105_), .Y(new_n1106_));
  NOR2X1   g721(.A(\b[121] ), .B(\a[121] ), .Y(new_n1107_));
  AND2X1   g722(.A(\b[121] ), .B(\a[121] ), .Y(new_n1108_));
  OR2X1    g723(.A(new_n1108_), .B(new_n1107_), .Y(new_n1109_));
  XOR2X1   g724(.A(new_n1109_), .B(new_n1106_), .Y(\f[121] ));
  INVX1    g725(.A(new_n1108_), .Y(new_n1111_));
  OAI21X1  g726(.A0(new_n1107_), .A1(new_n1106_), .B0(new_n1111_), .Y(new_n1112_));
  XOR2X1   g727(.A(\b[122] ), .B(\a[122] ), .Y(new_n1113_));
  XOR2X1   g728(.A(new_n1113_), .B(new_n1112_), .Y(\f[122] ));
  NOR2X1   g729(.A(\b[122] ), .B(\a[122] ), .Y(new_n1115_));
  INVX1    g730(.A(new_n1115_), .Y(new_n1116_));
  AND2X1   g731(.A(\b[122] ), .B(\a[122] ), .Y(new_n1117_));
  AOI21X1  g732(.A0(new_n1116_), .A1(new_n1112_), .B0(new_n1117_), .Y(new_n1118_));
  NOR2X1   g733(.A(\b[123] ), .B(\a[123] ), .Y(new_n1119_));
  AND2X1   g734(.A(\b[123] ), .B(\a[123] ), .Y(new_n1120_));
  OR2X1    g735(.A(new_n1120_), .B(new_n1119_), .Y(new_n1121_));
  XOR2X1   g736(.A(new_n1121_), .B(new_n1118_), .Y(\f[123] ));
  INVX1    g737(.A(new_n1120_), .Y(new_n1123_));
  OAI21X1  g738(.A0(new_n1119_), .A1(new_n1118_), .B0(new_n1123_), .Y(new_n1124_));
  XOR2X1   g739(.A(\b[124] ), .B(\a[124] ), .Y(new_n1125_));
  XOR2X1   g740(.A(new_n1125_), .B(new_n1124_), .Y(\f[124] ));
  NOR2X1   g741(.A(\b[124] ), .B(\a[124] ), .Y(new_n1127_));
  INVX1    g742(.A(new_n1127_), .Y(new_n1128_));
  AND2X1   g743(.A(\b[124] ), .B(\a[124] ), .Y(new_n1129_));
  AOI21X1  g744(.A0(new_n1128_), .A1(new_n1124_), .B0(new_n1129_), .Y(new_n1130_));
  NOR2X1   g745(.A(\b[125] ), .B(\a[125] ), .Y(new_n1131_));
  AND2X1   g746(.A(\b[125] ), .B(\a[125] ), .Y(new_n1132_));
  OR2X1    g747(.A(new_n1132_), .B(new_n1131_), .Y(new_n1133_));
  XOR2X1   g748(.A(new_n1133_), .B(new_n1130_), .Y(\f[125] ));
  INVX1    g749(.A(new_n1132_), .Y(new_n1135_));
  OAI21X1  g750(.A0(new_n1131_), .A1(new_n1130_), .B0(new_n1135_), .Y(new_n1136_));
  XOR2X1   g751(.A(\b[126] ), .B(\a[126] ), .Y(new_n1137_));
  XOR2X1   g752(.A(new_n1137_), .B(new_n1136_), .Y(\f[126] ));
  NOR2X1   g753(.A(\b[126] ), .B(\a[126] ), .Y(new_n1139_));
  INVX1    g754(.A(new_n1139_), .Y(new_n1140_));
  AND2X1   g755(.A(\b[126] ), .B(\a[126] ), .Y(new_n1141_));
  AOI21X1  g756(.A0(new_n1140_), .A1(new_n1136_), .B0(new_n1141_), .Y(new_n1142_));
  INVX1    g757(.A(\a[127] ), .Y(new_n1143_));
  XOR2X1   g758(.A(\b[127] ), .B(new_n1143_), .Y(new_n1144_));
  XOR2X1   g759(.A(new_n1144_), .B(new_n1142_), .Y(\f[127] ));
  NOR2X1   g760(.A(\b[127] ), .B(\a[127] ), .Y(new_n1146_));
  NAND2X1  g761(.A(\b[127] ), .B(\a[127] ), .Y(new_n1147_));
  OAI21X1  g762(.A0(new_n1146_), .A1(new_n1142_), .B0(new_n1147_), .Y(cOut));
endmodule


