// Benchmark "top" written by ABC on Mon Sep 21 03:42:05 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] ,
    \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] ,
    \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] ,
    \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] ,
    \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \b[0] ,
    \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] ,
    \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] ,
    \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] ,
    \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] ,
    \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] ,
    \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] ,
    \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] ,
    \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ,
    \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] ,
    \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] ,
    \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] ,
    \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] ,
    \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] ,
    \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] ,
    \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] ,
    \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] ,
    \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] ,
    \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] ,
    \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] ,
    \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] ,
    \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] ,
    \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] ,
    \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] ,
    \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] ,
    \f[125] , \f[126] , \f[127]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] ,
    \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] ,
    \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] ,
    \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] ,
    \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] ,
    \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] ,
    \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] ,
    \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] ,
    \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] ,
    \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] ,
    \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] ,
    \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] ;
  output \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] ,
    \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] ,
    \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] ,
    \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] ,
    \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] ,
    \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] ,
    \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] ,
    \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] ,
    \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] ,
    \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] ,
    \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] ,
    \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] ,
    \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] ,
    \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] ,
    \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] ,
    \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] ,
    \f[124] , \f[125] , \f[126] , \f[127] ;
  wire new_n257_, new_n258_, new_n259_, new_n260_, new_n262_, new_n263_,
    new_n264_, new_n265_, new_n266_, new_n267_, new_n268_, new_n269_,
    new_n270_, new_n272_, new_n273_, new_n274_, new_n275_, new_n276_,
    new_n277_, new_n278_, new_n279_, new_n280_, new_n281_, new_n282_,
    new_n283_, new_n284_, new_n285_, new_n286_, new_n287_, new_n288_,
    new_n289_, new_n291_, new_n292_, new_n293_, new_n294_, new_n295_,
    new_n296_, new_n297_, new_n298_, new_n299_, new_n300_, new_n301_,
    new_n302_, new_n303_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n385_, new_n386_, new_n387_, new_n388_, new_n389_,
    new_n390_, new_n391_, new_n392_, new_n393_, new_n394_, new_n395_,
    new_n396_, new_n397_, new_n398_, new_n399_, new_n400_, new_n401_,
    new_n402_, new_n403_, new_n404_, new_n405_, new_n406_, new_n407_,
    new_n408_, new_n409_, new_n410_, new_n411_, new_n412_, new_n413_,
    new_n414_, new_n415_, new_n416_, new_n417_, new_n418_, new_n419_,
    new_n420_, new_n421_, new_n422_, new_n423_, new_n424_, new_n425_,
    new_n426_, new_n428_, new_n429_, new_n430_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n437_, new_n438_,
    new_n439_, new_n440_, new_n441_, new_n442_, new_n443_, new_n444_,
    new_n445_, new_n446_, new_n447_, new_n448_, new_n449_, new_n450_,
    new_n451_, new_n452_, new_n453_, new_n454_, new_n455_, new_n456_,
    new_n457_, new_n458_, new_n459_, new_n460_, new_n461_, new_n463_,
    new_n464_, new_n465_, new_n466_, new_n467_, new_n468_, new_n469_,
    new_n470_, new_n471_, new_n472_, new_n473_, new_n474_, new_n475_,
    new_n476_, new_n477_, new_n478_, new_n479_, new_n480_, new_n481_,
    new_n482_, new_n483_, new_n484_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n491_, new_n492_, new_n493_,
    new_n494_, new_n495_, new_n496_, new_n497_, new_n498_, new_n499_,
    new_n500_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n644_, new_n645_, new_n646_, new_n647_,
    new_n648_, new_n649_, new_n650_, new_n651_, new_n652_, new_n653_,
    new_n654_, new_n655_, new_n656_, new_n657_, new_n658_, new_n659_,
    new_n660_, new_n661_, new_n662_, new_n663_, new_n664_, new_n665_,
    new_n666_, new_n667_, new_n668_, new_n669_, new_n670_, new_n671_,
    new_n672_, new_n673_, new_n674_, new_n675_, new_n676_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n683_,
    new_n684_, new_n685_, new_n686_, new_n687_, new_n688_, new_n689_,
    new_n690_, new_n691_, new_n692_, new_n693_, new_n694_, new_n695_,
    new_n696_, new_n697_, new_n698_, new_n699_, new_n700_, new_n701_,
    new_n702_, new_n703_, new_n704_, new_n705_, new_n706_, new_n707_,
    new_n708_, new_n709_, new_n710_, new_n711_, new_n712_, new_n713_,
    new_n714_, new_n715_, new_n716_, new_n717_, new_n718_, new_n719_,
    new_n720_, new_n721_, new_n722_, new_n723_, new_n724_, new_n725_,
    new_n726_, new_n728_, new_n729_, new_n730_, new_n731_, new_n732_,
    new_n733_, new_n734_, new_n735_, new_n736_, new_n737_, new_n738_,
    new_n739_, new_n740_, new_n741_, new_n742_, new_n743_, new_n744_,
    new_n745_, new_n746_, new_n747_, new_n748_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n760_, new_n761_, new_n762_,
    new_n763_, new_n764_, new_n765_, new_n766_, new_n767_, new_n768_,
    new_n769_, new_n770_, new_n771_, new_n772_, new_n773_, new_n774_,
    new_n775_, new_n776_, new_n777_, new_n778_, new_n779_, new_n780_,
    new_n781_, new_n782_, new_n783_, new_n784_, new_n786_, new_n787_,
    new_n788_, new_n789_, new_n790_, new_n791_, new_n792_, new_n793_,
    new_n794_, new_n795_, new_n796_, new_n797_, new_n798_, new_n799_,
    new_n800_, new_n801_, new_n802_, new_n803_, new_n804_, new_n805_,
    new_n806_, new_n807_, new_n808_, new_n809_, new_n810_, new_n811_,
    new_n812_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n821_, new_n822_, new_n823_,
    new_n824_, new_n825_, new_n826_, new_n827_, new_n828_, new_n829_,
    new_n830_, new_n831_, new_n832_, new_n833_, new_n834_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1052_, new_n1053_, new_n1054_, new_n1055_,
    new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_, new_n1061_,
    new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_, new_n1067_,
    new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_, new_n1073_,
    new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_, new_n1079_,
    new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_, new_n1085_,
    new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_, new_n1091_,
    new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_, new_n1097_,
    new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_, new_n1103_,
    new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_, new_n1109_,
    new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_, new_n1115_,
    new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_, new_n1121_,
    new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_, new_n1127_,
    new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_, new_n1133_,
    new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_, new_n1139_,
    new_n1141_, new_n1142_, new_n1143_, new_n1144_, new_n1145_, new_n1146_,
    new_n1147_, new_n1148_, new_n1149_, new_n1150_, new_n1151_, new_n1152_,
    new_n1153_, new_n1154_, new_n1155_, new_n1156_, new_n1157_, new_n1158_,
    new_n1159_, new_n1160_, new_n1161_, new_n1162_, new_n1163_, new_n1164_,
    new_n1165_, new_n1166_, new_n1167_, new_n1168_, new_n1169_, new_n1170_,
    new_n1171_, new_n1172_, new_n1173_, new_n1174_, new_n1175_, new_n1176_,
    new_n1177_, new_n1178_, new_n1179_, new_n1180_, new_n1181_, new_n1182_,
    new_n1183_, new_n1184_, new_n1185_, new_n1186_, new_n1187_, new_n1188_,
    new_n1189_, new_n1190_, new_n1191_, new_n1192_, new_n1193_, new_n1194_,
    new_n1195_, new_n1196_, new_n1197_, new_n1198_, new_n1199_, new_n1200_,
    new_n1201_, new_n1202_, new_n1203_, new_n1204_, new_n1205_, new_n1206_,
    new_n1207_, new_n1208_, new_n1209_, new_n1210_, new_n1211_, new_n1212_,
    new_n1213_, new_n1214_, new_n1215_, new_n1216_, new_n1217_, new_n1218_,
    new_n1219_, new_n1220_, new_n1221_, new_n1222_, new_n1223_, new_n1224_,
    new_n1225_, new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_,
    new_n1232_, new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_,
    new_n1238_, new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_,
    new_n1244_, new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_,
    new_n1250_, new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_,
    new_n1256_, new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_,
    new_n1262_, new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_,
    new_n1268_, new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_,
    new_n1274_, new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_,
    new_n1280_, new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_,
    new_n1286_, new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_,
    new_n1292_, new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_,
    new_n1298_, new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_,
    new_n1304_, new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1582_, new_n1583_,
    new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_, new_n1589_,
    new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_, new_n1595_,
    new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_, new_n1601_,
    new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_, new_n1607_,
    new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_, new_n1613_,
    new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_, new_n1619_,
    new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_, new_n1625_,
    new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_, new_n1631_,
    new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_, new_n1637_,
    new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_, new_n1643_,
    new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_, new_n1649_,
    new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_, new_n1655_,
    new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_, new_n1661_,
    new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_, new_n1667_,
    new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_, new_n1673_,
    new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_, new_n1679_,
    new_n1680_, new_n1681_, new_n1682_, new_n1684_, new_n1685_, new_n1686_,
    new_n1687_, new_n1688_, new_n1689_, new_n1690_, new_n1691_, new_n1692_,
    new_n1693_, new_n1694_, new_n1695_, new_n1696_, new_n1697_, new_n1698_,
    new_n1699_, new_n1700_, new_n1701_, new_n1702_, new_n1703_, new_n1704_,
    new_n1705_, new_n1706_, new_n1707_, new_n1708_, new_n1709_, new_n1710_,
    new_n1711_, new_n1712_, new_n1713_, new_n1714_, new_n1715_, new_n1716_,
    new_n1717_, new_n1718_, new_n1719_, new_n1720_, new_n1721_, new_n1722_,
    new_n1723_, new_n1724_, new_n1725_, new_n1726_, new_n1727_, new_n1728_,
    new_n1729_, new_n1730_, new_n1731_, new_n1732_, new_n1733_, new_n1734_,
    new_n1735_, new_n1736_, new_n1737_, new_n1738_, new_n1739_, new_n1740_,
    new_n1741_, new_n1742_, new_n1743_, new_n1744_, new_n1745_, new_n1746_,
    new_n1747_, new_n1748_, new_n1749_, new_n1750_, new_n1751_, new_n1752_,
    new_n1753_, new_n1754_, new_n1755_, new_n1756_, new_n1757_, new_n1758_,
    new_n1759_, new_n1760_, new_n1761_, new_n1762_, new_n1763_, new_n1764_,
    new_n1765_, new_n1766_, new_n1767_, new_n1768_, new_n1769_, new_n1770_,
    new_n1771_, new_n1772_, new_n1773_, new_n1774_, new_n1775_, new_n1776_,
    new_n1777_, new_n1778_, new_n1779_, new_n1780_, new_n1781_, new_n1782_,
    new_n1783_, new_n1784_, new_n1785_, new_n1786_, new_n1787_, new_n1788_,
    new_n1790_, new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_,
    new_n1796_, new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_,
    new_n1802_, new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_,
    new_n1808_, new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_,
    new_n1814_, new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_,
    new_n1820_, new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_,
    new_n1826_, new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_,
    new_n1832_, new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_,
    new_n1838_, new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_,
    new_n1844_, new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_,
    new_n1850_, new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_,
    new_n1856_, new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_,
    new_n1862_, new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_,
    new_n1868_, new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_,
    new_n1874_, new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_,
    new_n1880_, new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_,
    new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_,
    new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_,
    new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_, new_n2230_,
    new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_, new_n2236_,
    new_n2237_, new_n2238_, new_n2239_, new_n2241_, new_n2242_, new_n2243_,
    new_n2244_, new_n2245_, new_n2246_, new_n2247_, new_n2248_, new_n2249_,
    new_n2250_, new_n2251_, new_n2252_, new_n2253_, new_n2254_, new_n2255_,
    new_n2256_, new_n2257_, new_n2258_, new_n2259_, new_n2260_, new_n2261_,
    new_n2262_, new_n2263_, new_n2264_, new_n2265_, new_n2266_, new_n2267_,
    new_n2268_, new_n2269_, new_n2270_, new_n2271_, new_n2272_, new_n2273_,
    new_n2274_, new_n2275_, new_n2276_, new_n2277_, new_n2278_, new_n2279_,
    new_n2280_, new_n2281_, new_n2282_, new_n2283_, new_n2284_, new_n2285_,
    new_n2286_, new_n2287_, new_n2288_, new_n2289_, new_n2290_, new_n2291_,
    new_n2292_, new_n2293_, new_n2294_, new_n2295_, new_n2296_, new_n2297_,
    new_n2298_, new_n2299_, new_n2300_, new_n2301_, new_n2302_, new_n2303_,
    new_n2304_, new_n2305_, new_n2306_, new_n2307_, new_n2308_, new_n2309_,
    new_n2310_, new_n2311_, new_n2312_, new_n2313_, new_n2314_, new_n2315_,
    new_n2316_, new_n2317_, new_n2318_, new_n2319_, new_n2320_, new_n2321_,
    new_n2322_, new_n2323_, new_n2324_, new_n2325_, new_n2326_, new_n2327_,
    new_n2328_, new_n2329_, new_n2330_, new_n2331_, new_n2332_, new_n2333_,
    new_n2334_, new_n2335_, new_n2336_, new_n2337_, new_n2338_, new_n2339_,
    new_n2340_, new_n2341_, new_n2342_, new_n2343_, new_n2344_, new_n2345_,
    new_n2346_, new_n2347_, new_n2348_, new_n2349_, new_n2350_, new_n2351_,
    new_n2352_, new_n2353_, new_n2354_, new_n2355_, new_n2356_, new_n2357_,
    new_n2358_, new_n2359_, new_n2360_, new_n2361_, new_n2362_, new_n2363_,
    new_n2364_, new_n2365_, new_n2366_, new_n2367_, new_n2368_, new_n2370_,
    new_n2371_, new_n2372_, new_n2373_, new_n2374_, new_n2375_, new_n2376_,
    new_n2377_, new_n2378_, new_n2379_, new_n2380_, new_n2381_, new_n2382_,
    new_n2383_, new_n2384_, new_n2385_, new_n2386_, new_n2387_, new_n2388_,
    new_n2389_, new_n2390_, new_n2391_, new_n2392_, new_n2393_, new_n2394_,
    new_n2395_, new_n2396_, new_n2397_, new_n2398_, new_n2399_, new_n2400_,
    new_n2401_, new_n2402_, new_n2403_, new_n2404_, new_n2405_, new_n2406_,
    new_n2407_, new_n2408_, new_n2409_, new_n2410_, new_n2411_, new_n2412_,
    new_n2413_, new_n2414_, new_n2415_, new_n2416_, new_n2417_, new_n2418_,
    new_n2419_, new_n2420_, new_n2421_, new_n2422_, new_n2423_, new_n2424_,
    new_n2425_, new_n2426_, new_n2427_, new_n2428_, new_n2429_, new_n2430_,
    new_n2431_, new_n2432_, new_n2433_, new_n2434_, new_n2435_, new_n2436_,
    new_n2437_, new_n2438_, new_n2439_, new_n2440_, new_n2441_, new_n2442_,
    new_n2443_, new_n2444_, new_n2445_, new_n2446_, new_n2447_, new_n2448_,
    new_n2449_, new_n2450_, new_n2451_, new_n2452_, new_n2453_, new_n2454_,
    new_n2455_, new_n2456_, new_n2457_, new_n2458_, new_n2459_, new_n2460_,
    new_n2461_, new_n2462_, new_n2463_, new_n2464_, new_n2465_, new_n2466_,
    new_n2467_, new_n2468_, new_n2469_, new_n2470_, new_n2471_, new_n2472_,
    new_n2473_, new_n2474_, new_n2475_, new_n2476_, new_n2477_, new_n2478_,
    new_n2479_, new_n2480_, new_n2481_, new_n2482_, new_n2483_, new_n2484_,
    new_n2485_, new_n2486_, new_n2487_, new_n2488_, new_n2489_, new_n2490_,
    new_n2491_, new_n2492_, new_n2493_, new_n2494_, new_n2495_, new_n2496_,
    new_n2497_, new_n2498_, new_n2499_, new_n2500_, new_n2501_, new_n2502_,
    new_n2503_, new_n2504_, new_n2505_, new_n2506_, new_n2507_, new_n2508_,
    new_n2509_, new_n2510_, new_n2511_, new_n2513_, new_n2514_, new_n2515_,
    new_n2516_, new_n2517_, new_n2518_, new_n2519_, new_n2520_, new_n2521_,
    new_n2522_, new_n2523_, new_n2524_, new_n2525_, new_n2526_, new_n2527_,
    new_n2528_, new_n2529_, new_n2530_, new_n2531_, new_n2532_, new_n2533_,
    new_n2534_, new_n2535_, new_n2536_, new_n2537_, new_n2538_, new_n2539_,
    new_n2540_, new_n2541_, new_n2542_, new_n2543_, new_n2544_, new_n2545_,
    new_n2546_, new_n2547_, new_n2548_, new_n2549_, new_n2550_, new_n2551_,
    new_n2552_, new_n2553_, new_n2554_, new_n2555_, new_n2556_, new_n2557_,
    new_n2558_, new_n2559_, new_n2560_, new_n2561_, new_n2562_, new_n2563_,
    new_n2564_, new_n2565_, new_n2566_, new_n2567_, new_n2568_, new_n2569_,
    new_n2570_, new_n2571_, new_n2572_, new_n2573_, new_n2574_, new_n2575_,
    new_n2576_, new_n2577_, new_n2578_, new_n2579_, new_n2580_, new_n2581_,
    new_n2582_, new_n2583_, new_n2584_, new_n2585_, new_n2586_, new_n2587_,
    new_n2588_, new_n2589_, new_n2590_, new_n2591_, new_n2592_, new_n2593_,
    new_n2594_, new_n2595_, new_n2596_, new_n2597_, new_n2598_, new_n2599_,
    new_n2600_, new_n2601_, new_n2602_, new_n2603_, new_n2604_, new_n2605_,
    new_n2606_, new_n2607_, new_n2608_, new_n2609_, new_n2610_, new_n2611_,
    new_n2612_, new_n2613_, new_n2614_, new_n2615_, new_n2616_, new_n2617_,
    new_n2618_, new_n2619_, new_n2620_, new_n2622_, new_n2623_, new_n2624_,
    new_n2625_, new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_,
    new_n2631_, new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_,
    new_n2637_, new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_,
    new_n2643_, new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_,
    new_n2649_, new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_,
    new_n2655_, new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_,
    new_n2661_, new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_,
    new_n2667_, new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_,
    new_n2673_, new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_,
    new_n2679_, new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_,
    new_n2685_, new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_,
    new_n2691_, new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_,
    new_n2697_, new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_,
    new_n2703_, new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_,
    new_n2709_, new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_,
    new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_,
    new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_,
    new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_,
    new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_,
    new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_,
    new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_,
    new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_,
    new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_,
    new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_,
    new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_,
    new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_,
    new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_,
    new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_,
    new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_,
    new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_,
    new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_,
    new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_,
    new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_,
    new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_, new_n3089_,
    new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_, new_n3095_,
    new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_, new_n3101_,
    new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_, new_n3107_,
    new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_, new_n3113_,
    new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_, new_n3119_,
    new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_, new_n3125_,
    new_n3126_, new_n3127_, new_n3128_, new_n3129_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_, new_n3168_,
    new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_, new_n3174_,
    new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_, new_n3180_,
    new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_, new_n3186_,
    new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_, new_n3192_,
    new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_, new_n3198_,
    new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_, new_n3204_,
    new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_, new_n3210_,
    new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_, new_n3216_,
    new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_, new_n3222_,
    new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_, new_n3228_,
    new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_, new_n3234_,
    new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_, new_n3240_,
    new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_, new_n3246_,
    new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_, new_n3252_,
    new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_, new_n3258_,
    new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_, new_n3264_,
    new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_, new_n3270_,
    new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_, new_n3276_,
    new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_, new_n3282_,
    new_n3283_, new_n3284_, new_n3286_, new_n3287_, new_n3288_, new_n3289_,
    new_n3290_, new_n3291_, new_n3292_, new_n3293_, new_n3294_, new_n3295_,
    new_n3296_, new_n3297_, new_n3298_, new_n3299_, new_n3300_, new_n3301_,
    new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_, new_n3307_,
    new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_, new_n3313_,
    new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_, new_n3319_,
    new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_, new_n3325_,
    new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_, new_n3331_,
    new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_, new_n3337_,
    new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_, new_n3343_,
    new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_, new_n3361_,
    new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_,
    new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_,
    new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_, new_n3379_,
    new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_, new_n3385_,
    new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_, new_n3391_,
    new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_, new_n3397_,
    new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_, new_n3403_,
    new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_, new_n3409_,
    new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_, new_n3415_,
    new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_,
    new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_,
    new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_,
    new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_,
    new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_,
    new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_,
    new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_,
    new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_,
    new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_,
    new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_,
    new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_,
    new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_,
    new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_,
    new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_,
    new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_,
    new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_,
    new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_,
    new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_,
    new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_,
    new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_,
    new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_,
    new_n3555_, new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3730_,
    new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_, new_n3736_,
    new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_, new_n3742_,
    new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_, new_n3748_,
    new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_, new_n3754_,
    new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_, new_n3760_,
    new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_, new_n3766_,
    new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_, new_n3772_,
    new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_, new_n3778_,
    new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_, new_n3784_,
    new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_, new_n3790_,
    new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_, new_n3796_,
    new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_, new_n3802_,
    new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_, new_n3808_,
    new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_, new_n3814_,
    new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_, new_n3820_,
    new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_, new_n3826_,
    new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_, new_n3832_,
    new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_, new_n3838_,
    new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_, new_n3844_,
    new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_, new_n3850_,
    new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_, new_n3856_,
    new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_,
    new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_,
    new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_, new_n3875_,
    new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_, new_n3881_,
    new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_, new_n3887_,
    new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_, new_n3893_,
    new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_, new_n3899_,
    new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_, new_n3905_,
    new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_, new_n3911_,
    new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_, new_n3917_,
    new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_, new_n3923_,
    new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_, new_n3929_,
    new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_, new_n3935_,
    new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_, new_n3941_,
    new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_, new_n3947_,
    new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_, new_n3953_,
    new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_, new_n3959_,
    new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_, new_n3965_,
    new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_, new_n3971_,
    new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_, new_n3977_,
    new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_, new_n3983_,
    new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_, new_n3989_,
    new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_, new_n3995_,
    new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_, new_n4001_,
    new_n4002_, new_n4003_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4029_, new_n4030_, new_n4031_, new_n4032_,
    new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_, new_n4038_,
    new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_, new_n4044_,
    new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_, new_n4050_,
    new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_, new_n4056_,
    new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_, new_n4062_,
    new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_, new_n4068_,
    new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_, new_n4074_,
    new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_, new_n4080_,
    new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_, new_n4086_,
    new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_, new_n4092_,
    new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_, new_n4098_,
    new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_, new_n4104_,
    new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_, new_n4110_,
    new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_, new_n4116_,
    new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_, new_n4122_,
    new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_, new_n4128_,
    new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_, new_n4134_,
    new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_, new_n4140_,
    new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_, new_n4146_,
    new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_, new_n4152_,
    new_n4153_, new_n4154_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4185_, new_n4186_, new_n4187_, new_n4188_, new_n4189_,
    new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_, new_n4195_,
    new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_, new_n4201_,
    new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_, new_n4207_,
    new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_, new_n4213_,
    new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_, new_n4219_,
    new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_, new_n4225_,
    new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_, new_n4231_,
    new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_, new_n4237_,
    new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_, new_n4243_,
    new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_, new_n4249_,
    new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_, new_n4255_,
    new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_, new_n4261_,
    new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_, new_n4267_,
    new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_, new_n4273_,
    new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_, new_n4279_,
    new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_, new_n4285_,
    new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_, new_n4291_,
    new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_, new_n4297_,
    new_n4298_, new_n4299_, new_n4300_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4346_,
    new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_,
    new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_,
    new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_,
    new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_,
    new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_,
    new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_,
    new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_,
    new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_,
    new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_,
    new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_,
    new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_,
    new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_,
    new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_,
    new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_,
    new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_,
    new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_,
    new_n4443_, new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_,
    new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_,
    new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_,
    new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_,
    new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_,
    new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_,
    new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_,
    new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_,
    new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4519_, new_n4520_, new_n4521_,
    new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_,
    new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_,
    new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_,
    new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_,
    new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_,
    new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_,
    new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4686_, new_n4687_, new_n4688_, new_n4689_, new_n4690_,
    new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_, new_n4696_,
    new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_, new_n4702_,
    new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_, new_n4708_,
    new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_, new_n4714_,
    new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_, new_n4720_,
    new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_, new_n4726_,
    new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_, new_n4732_,
    new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_, new_n4738_,
    new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_, new_n4744_,
    new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_, new_n4750_,
    new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_,
    new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_,
    new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_,
    new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_,
    new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_,
    new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_,
    new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4846_, new_n4847_,
    new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_, new_n4853_,
    new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_, new_n4859_,
    new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_, new_n4865_,
    new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_, new_n4871_,
    new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_, new_n4877_,
    new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_, new_n4883_,
    new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_, new_n4889_,
    new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_, new_n4895_,
    new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_, new_n4901_,
    new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_, new_n4907_,
    new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_, new_n4913_,
    new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_, new_n4919_,
    new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_, new_n4925_,
    new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_, new_n4931_,
    new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_, new_n4937_,
    new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_, new_n4943_,
    new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_, new_n4949_,
    new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_, new_n4955_,
    new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_, new_n4961_,
    new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_, new_n4967_,
    new_n4968_, new_n4969_, new_n4970_, new_n4971_, new_n4972_, new_n4973_,
    new_n4974_, new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_,
    new_n4980_, new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_,
    new_n4986_, new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_,
    new_n4992_, new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_,
    new_n4998_, new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_,
    new_n5004_, new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_,
    new_n5010_, new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_,
    new_n5016_, new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_,
    new_n5022_, new_n5023_, new_n5024_, new_n5025_, new_n5026_, new_n5027_,
    new_n5028_, new_n5029_, new_n5030_, new_n5031_, new_n5032_, new_n5033_,
    new_n5034_, new_n5035_, new_n5036_, new_n5037_, new_n5038_, new_n5039_,
    new_n5040_, new_n5041_, new_n5042_, new_n5043_, new_n5044_, new_n5046_,
    new_n5047_, new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_,
    new_n5053_, new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_,
    new_n5059_, new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_,
    new_n5065_, new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_,
    new_n5071_, new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_,
    new_n5077_, new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_,
    new_n5083_, new_n5084_, new_n5085_, new_n5086_, new_n5087_, new_n5088_,
    new_n5089_, new_n5090_, new_n5091_, new_n5092_, new_n5093_, new_n5094_,
    new_n5095_, new_n5096_, new_n5097_, new_n5098_, new_n5099_, new_n5100_,
    new_n5101_, new_n5102_, new_n5103_, new_n5104_, new_n5105_, new_n5106_,
    new_n5107_, new_n5108_, new_n5109_, new_n5110_, new_n5111_, new_n5112_,
    new_n5113_, new_n5114_, new_n5115_, new_n5116_, new_n5117_, new_n5118_,
    new_n5119_, new_n5120_, new_n5121_, new_n5122_, new_n5123_, new_n5124_,
    new_n5125_, new_n5126_, new_n5127_, new_n5128_, new_n5129_, new_n5130_,
    new_n5131_, new_n5132_, new_n5133_, new_n5134_, new_n5135_, new_n5136_,
    new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_, new_n5142_,
    new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_, new_n5148_,
    new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_, new_n5154_,
    new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_, new_n5160_,
    new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_, new_n5166_,
    new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_, new_n5172_,
    new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_, new_n5178_,
    new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_, new_n5184_,
    new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_, new_n5190_,
    new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_, new_n5196_,
    new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_, new_n5202_,
    new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_, new_n5208_,
    new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5214_, new_n5215_,
    new_n5216_, new_n5217_, new_n5218_, new_n5219_, new_n5220_, new_n5221_,
    new_n5222_, new_n5223_, new_n5224_, new_n5225_, new_n5226_, new_n5227_,
    new_n5228_, new_n5229_, new_n5230_, new_n5231_, new_n5232_, new_n5233_,
    new_n5234_, new_n5235_, new_n5236_, new_n5237_, new_n5238_, new_n5239_,
    new_n5240_, new_n5241_, new_n5242_, new_n5243_, new_n5244_, new_n5245_,
    new_n5246_, new_n5247_, new_n5248_, new_n5249_, new_n5250_, new_n5251_,
    new_n5252_, new_n5253_, new_n5254_, new_n5255_, new_n5256_, new_n5257_,
    new_n5258_, new_n5259_, new_n5260_, new_n5261_, new_n5262_, new_n5263_,
    new_n5264_, new_n5265_, new_n5266_, new_n5267_, new_n5268_, new_n5269_,
    new_n5270_, new_n5271_, new_n5272_, new_n5273_, new_n5274_, new_n5275_,
    new_n5276_, new_n5277_, new_n5278_, new_n5279_, new_n5280_, new_n5281_,
    new_n5282_, new_n5283_, new_n5284_, new_n5285_, new_n5286_, new_n5287_,
    new_n5288_, new_n5289_, new_n5290_, new_n5291_, new_n5292_, new_n5293_,
    new_n5294_, new_n5295_, new_n5296_, new_n5297_, new_n5298_, new_n5299_,
    new_n5300_, new_n5301_, new_n5302_, new_n5303_, new_n5304_, new_n5305_,
    new_n5306_, new_n5307_, new_n5308_, new_n5309_, new_n5310_, new_n5311_,
    new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_, new_n5317_,
    new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_, new_n5323_,
    new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_, new_n5329_,
    new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_, new_n5335_,
    new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_, new_n5341_,
    new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_, new_n5347_,
    new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_, new_n5353_,
    new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_, new_n5359_,
    new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_, new_n5365_,
    new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_, new_n5371_,
    new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_, new_n5377_,
    new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_, new_n5383_,
    new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_, new_n5389_,
    new_n5390_, new_n5391_, new_n5393_, new_n5394_, new_n5395_, new_n5396_,
    new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_,
    new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_,
    new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_,
    new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_,
    new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_,
    new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_,
    new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_,
    new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_,
    new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_,
    new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_,
    new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_,
    new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_,
    new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_,
    new_n5475_, new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_,
    new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_,
    new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_,
    new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_,
    new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_,
    new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_,
    new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_,
    new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_,
    new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_,
    new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_,
    new_n5535_, new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_,
    new_n5541_, new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_,
    new_n5547_, new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_,
    new_n5553_, new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_,
    new_n5559_, new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_,
    new_n5565_, new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_,
    new_n5571_, new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_,
    new_n5577_, new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_,
    new_n5583_, new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_,
    new_n5589_, new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_,
    new_n5595_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_,
    new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_,
    new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_,
    new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_,
    new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_,
    new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_,
    new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_,
    new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_,
    new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_,
    new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_,
    new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_,
    new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_,
    new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_,
    new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_,
    new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_,
    new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_,
    new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_,
    new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_,
    new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_,
    new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_,
    new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_,
    new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_,
    new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_,
    new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_,
    new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_,
    new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_,
    new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_,
    new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_,
    new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_,
    new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_,
    new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_,
    new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_,
    new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_,
    new_n5800_, new_n5802_, new_n5803_, new_n5804_, new_n5805_, new_n5806_,
    new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_, new_n5812_,
    new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_, new_n5818_,
    new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_, new_n5824_,
    new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_, new_n5830_,
    new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_, new_n5836_,
    new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_, new_n5842_,
    new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_, new_n5848_,
    new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_, new_n5854_,
    new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_, new_n5860_,
    new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_, new_n5866_,
    new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_, new_n5872_,
    new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_, new_n5878_,
    new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_, new_n5884_,
    new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_, new_n5890_,
    new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_, new_n5896_,
    new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_, new_n5902_,
    new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_, new_n5908_,
    new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_, new_n5914_,
    new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_, new_n5920_,
    new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_, new_n5926_,
    new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_, new_n5932_,
    new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_, new_n5938_,
    new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_, new_n5944_,
    new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_, new_n5950_,
    new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_, new_n5956_,
    new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_, new_n5962_,
    new_n5963_, new_n5964_, new_n5966_, new_n5967_, new_n5968_, new_n5969_,
    new_n5970_, new_n5971_, new_n5972_, new_n5973_, new_n5974_, new_n5975_,
    new_n5976_, new_n5977_, new_n5978_, new_n5979_, new_n5980_, new_n5981_,
    new_n5982_, new_n5983_, new_n5984_, new_n5985_, new_n5986_, new_n5987_,
    new_n5988_, new_n5989_, new_n5990_, new_n5991_, new_n5992_, new_n5993_,
    new_n5994_, new_n5995_, new_n5996_, new_n5997_, new_n5998_, new_n5999_,
    new_n6000_, new_n6001_, new_n6002_, new_n6003_, new_n6004_, new_n6005_,
    new_n6006_, new_n6007_, new_n6008_, new_n6009_, new_n6010_, new_n6011_,
    new_n6012_, new_n6013_, new_n6014_, new_n6015_, new_n6016_, new_n6017_,
    new_n6018_, new_n6019_, new_n6020_, new_n6021_, new_n6022_, new_n6023_,
    new_n6024_, new_n6025_, new_n6026_, new_n6027_, new_n6028_, new_n6029_,
    new_n6030_, new_n6031_, new_n6032_, new_n6033_, new_n6034_, new_n6035_,
    new_n6036_, new_n6037_, new_n6038_, new_n6039_, new_n6040_, new_n6041_,
    new_n6042_, new_n6043_, new_n6044_, new_n6045_, new_n6046_, new_n6047_,
    new_n6048_, new_n6049_, new_n6050_, new_n6051_, new_n6052_, new_n6053_,
    new_n6054_, new_n6055_, new_n6056_, new_n6057_, new_n6058_, new_n6059_,
    new_n6060_, new_n6061_, new_n6062_, new_n6063_, new_n6064_, new_n6065_,
    new_n6066_, new_n6067_, new_n6068_, new_n6069_, new_n6070_, new_n6071_,
    new_n6072_, new_n6073_, new_n6074_, new_n6075_, new_n6076_, new_n6077_,
    new_n6078_, new_n6079_, new_n6080_, new_n6081_, new_n6082_, new_n6083_,
    new_n6084_, new_n6085_, new_n6086_, new_n6087_, new_n6088_, new_n6089_,
    new_n6090_, new_n6091_, new_n6092_, new_n6093_, new_n6094_, new_n6095_,
    new_n6096_, new_n6097_, new_n6098_, new_n6099_, new_n6100_, new_n6101_,
    new_n6102_, new_n6103_, new_n6104_, new_n6105_, new_n6106_, new_n6107_,
    new_n6108_, new_n6109_, new_n6110_, new_n6111_, new_n6112_, new_n6113_,
    new_n6114_, new_n6115_, new_n6116_, new_n6117_, new_n6118_, new_n6119_,
    new_n6120_, new_n6121_, new_n6122_, new_n6123_, new_n6124_, new_n6125_,
    new_n6126_, new_n6127_, new_n6128_, new_n6129_, new_n6130_, new_n6131_,
    new_n6132_, new_n6133_, new_n6134_, new_n6135_, new_n6136_, new_n6137_,
    new_n6138_, new_n6139_, new_n6140_, new_n6141_, new_n6142_, new_n6143_,
    new_n6144_, new_n6145_, new_n6146_, new_n6147_, new_n6148_, new_n6149_,
    new_n6150_, new_n6151_, new_n6152_, new_n6153_, new_n6154_, new_n6155_,
    new_n6156_, new_n6158_, new_n6159_, new_n6160_, new_n6161_, new_n6162_,
    new_n6163_, new_n6164_, new_n6165_, new_n6166_, new_n6167_, new_n6168_,
    new_n6169_, new_n6170_, new_n6171_, new_n6172_, new_n6173_, new_n6174_,
    new_n6175_, new_n6176_, new_n6177_, new_n6178_, new_n6179_, new_n6180_,
    new_n6181_, new_n6182_, new_n6183_, new_n6184_, new_n6185_, new_n6186_,
    new_n6187_, new_n6188_, new_n6189_, new_n6190_, new_n6191_, new_n6192_,
    new_n6193_, new_n6194_, new_n6195_, new_n6196_, new_n6197_, new_n6198_,
    new_n6199_, new_n6200_, new_n6201_, new_n6202_, new_n6203_, new_n6204_,
    new_n6205_, new_n6206_, new_n6207_, new_n6208_, new_n6209_, new_n6210_,
    new_n6211_, new_n6212_, new_n6213_, new_n6214_, new_n6215_, new_n6216_,
    new_n6217_, new_n6218_, new_n6219_, new_n6220_, new_n6221_, new_n6222_,
    new_n6223_, new_n6224_, new_n6225_, new_n6226_, new_n6227_, new_n6228_,
    new_n6229_, new_n6230_, new_n6231_, new_n6232_, new_n6233_, new_n6234_,
    new_n6235_, new_n6236_, new_n6237_, new_n6238_, new_n6239_, new_n6240_,
    new_n6241_, new_n6242_, new_n6243_, new_n6244_, new_n6245_, new_n6246_,
    new_n6247_, new_n6248_, new_n6249_, new_n6250_, new_n6251_, new_n6252_,
    new_n6253_, new_n6254_, new_n6255_, new_n6256_, new_n6257_, new_n6258_,
    new_n6259_, new_n6260_, new_n6261_, new_n6262_, new_n6263_, new_n6264_,
    new_n6265_, new_n6266_, new_n6267_, new_n6268_, new_n6269_, new_n6270_,
    new_n6271_, new_n6272_, new_n6273_, new_n6274_, new_n6275_, new_n6276_,
    new_n6277_, new_n6278_, new_n6279_, new_n6280_, new_n6281_, new_n6282_,
    new_n6283_, new_n6284_, new_n6285_, new_n6286_, new_n6287_, new_n6288_,
    new_n6289_, new_n6290_, new_n6291_, new_n6292_, new_n6293_, new_n6294_,
    new_n6295_, new_n6296_, new_n6297_, new_n6298_, new_n6299_, new_n6300_,
    new_n6301_, new_n6302_, new_n6303_, new_n6304_, new_n6305_, new_n6306_,
    new_n6307_, new_n6308_, new_n6309_, new_n6310_, new_n6311_, new_n6312_,
    new_n6313_, new_n6314_, new_n6315_, new_n6316_, new_n6317_, new_n6318_,
    new_n6319_, new_n6320_, new_n6321_, new_n6322_, new_n6323_, new_n6324_,
    new_n6325_, new_n6326_, new_n6327_, new_n6328_, new_n6329_, new_n6330_,
    new_n6331_, new_n6332_, new_n6333_, new_n6334_, new_n6335_, new_n6336_,
    new_n6337_, new_n6338_, new_n6339_, new_n6340_, new_n6341_, new_n6342_,
    new_n6343_, new_n6344_, new_n6345_, new_n6346_, new_n6347_, new_n6348_,
    new_n6349_, new_n6350_, new_n6352_, new_n6353_, new_n6354_, new_n6355_,
    new_n6356_, new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_,
    new_n6362_, new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_,
    new_n6368_, new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_,
    new_n6374_, new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_,
    new_n6380_, new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_,
    new_n6386_, new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_,
    new_n6392_, new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_,
    new_n6398_, new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_,
    new_n6404_, new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_,
    new_n6410_, new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_,
    new_n6416_, new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_,
    new_n6422_, new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_,
    new_n6428_, new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_,
    new_n6434_, new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_,
    new_n6440_, new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_,
    new_n6446_, new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_,
    new_n6452_, new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_,
    new_n6458_, new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_,
    new_n6464_, new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_,
    new_n6470_, new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_,
    new_n6476_, new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_,
    new_n6482_, new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_,
    new_n6488_, new_n6489_, new_n6490_, new_n6491_, new_n6492_, new_n6493_,
    new_n6494_, new_n6495_, new_n6496_, new_n6497_, new_n6498_, new_n6499_,
    new_n6500_, new_n6501_, new_n6502_, new_n6503_, new_n6504_, new_n6505_,
    new_n6506_, new_n6507_, new_n6508_, new_n6509_, new_n6510_, new_n6511_,
    new_n6512_, new_n6513_, new_n6514_, new_n6515_, new_n6516_, new_n6517_,
    new_n6518_, new_n6519_, new_n6520_, new_n6521_, new_n6522_, new_n6523_,
    new_n6524_, new_n6525_, new_n6526_, new_n6527_, new_n6528_, new_n6529_,
    new_n6530_, new_n6531_, new_n6532_, new_n6534_, new_n6535_, new_n6536_,
    new_n6537_, new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_,
    new_n6543_, new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_,
    new_n6549_, new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_,
    new_n6555_, new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_,
    new_n6561_, new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_,
    new_n6567_, new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_,
    new_n6573_, new_n6574_, new_n6575_, new_n6576_, new_n6577_, new_n6578_,
    new_n6579_, new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_,
    new_n6585_, new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_,
    new_n6591_, new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_,
    new_n6597_, new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_,
    new_n6603_, new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_,
    new_n6609_, new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_,
    new_n6615_, new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_,
    new_n6621_, new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_,
    new_n6627_, new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_,
    new_n6633_, new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_,
    new_n6639_, new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_,
    new_n6645_, new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_,
    new_n6651_, new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_,
    new_n6657_, new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_,
    new_n6663_, new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_,
    new_n6669_, new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_,
    new_n6675_, new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_,
    new_n6681_, new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_,
    new_n6687_, new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_,
    new_n6693_, new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_,
    new_n6699_, new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_,
    new_n6705_, new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_,
    new_n6711_, new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_,
    new_n6717_, new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_,
    new_n6723_, new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_,
    new_n6729_, new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_,
    new_n6735_, new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_,
    new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_,
    new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_,
    new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_,
    new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_,
    new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_,
    new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_,
    new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_,
    new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_,
    new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_,
    new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_,
    new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_,
    new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_,
    new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_,
    new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_,
    new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_,
    new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_,
    new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_,
    new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_,
    new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_,
    new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6867_,
    new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_,
    new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_,
    new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_,
    new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_,
    new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_,
    new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_,
    new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_,
    new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_,
    new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_,
    new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_,
    new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_,
    new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_,
    new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_, new_n6946_,
    new_n6947_, new_n6948_, new_n6949_, new_n6950_, new_n6951_, new_n6952_,
    new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_, new_n6958_,
    new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_, new_n6964_,
    new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_, new_n6970_,
    new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_, new_n6976_,
    new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_, new_n6982_,
    new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_, new_n6988_,
    new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_, new_n6994_,
    new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_, new_n7000_,
    new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_, new_n7006_,
    new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_, new_n7012_,
    new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_, new_n7018_,
    new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_, new_n7024_,
    new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_, new_n7030_,
    new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_, new_n7036_,
    new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_, new_n7042_,
    new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_, new_n7048_,
    new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_, new_n7054_,
    new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_, new_n7060_,
    new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_, new_n7066_,
    new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_, new_n7072_,
    new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_, new_n7078_,
    new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_, new_n7084_,
    new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_, new_n7090_,
    new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_, new_n7096_,
    new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_, new_n7102_,
    new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_, new_n7108_,
    new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_, new_n7114_,
    new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_, new_n7120_,
    new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_, new_n7126_,
    new_n7127_, new_n7128_, new_n7129_, new_n7131_, new_n7132_, new_n7133_,
    new_n7134_, new_n7135_, new_n7136_, new_n7137_, new_n7138_, new_n7139_,
    new_n7140_, new_n7141_, new_n7142_, new_n7143_, new_n7144_, new_n7145_,
    new_n7146_, new_n7147_, new_n7148_, new_n7149_, new_n7150_, new_n7151_,
    new_n7152_, new_n7153_, new_n7154_, new_n7155_, new_n7156_, new_n7157_,
    new_n7158_, new_n7159_, new_n7160_, new_n7161_, new_n7162_, new_n7163_,
    new_n7164_, new_n7165_, new_n7166_, new_n7167_, new_n7168_, new_n7169_,
    new_n7170_, new_n7171_, new_n7172_, new_n7173_, new_n7174_, new_n7175_,
    new_n7176_, new_n7177_, new_n7178_, new_n7179_, new_n7180_, new_n7181_,
    new_n7182_, new_n7183_, new_n7184_, new_n7185_, new_n7186_, new_n7187_,
    new_n7188_, new_n7189_, new_n7190_, new_n7191_, new_n7192_, new_n7193_,
    new_n7194_, new_n7195_, new_n7196_, new_n7197_, new_n7198_, new_n7199_,
    new_n7200_, new_n7201_, new_n7202_, new_n7203_, new_n7204_, new_n7205_,
    new_n7206_, new_n7207_, new_n7208_, new_n7209_, new_n7210_, new_n7211_,
    new_n7212_, new_n7213_, new_n7214_, new_n7215_, new_n7216_, new_n7217_,
    new_n7218_, new_n7219_, new_n7220_, new_n7221_, new_n7222_, new_n7223_,
    new_n7224_, new_n7225_, new_n7226_, new_n7227_, new_n7228_, new_n7229_,
    new_n7230_, new_n7231_, new_n7232_, new_n7233_, new_n7234_, new_n7235_,
    new_n7236_, new_n7237_, new_n7238_, new_n7239_, new_n7240_, new_n7241_,
    new_n7242_, new_n7243_, new_n7244_, new_n7245_, new_n7246_, new_n7247_,
    new_n7248_, new_n7249_, new_n7250_, new_n7251_, new_n7252_, new_n7253_,
    new_n7254_, new_n7255_, new_n7256_, new_n7257_, new_n7258_, new_n7259_,
    new_n7260_, new_n7261_, new_n7262_, new_n7263_, new_n7264_, new_n7265_,
    new_n7266_, new_n7267_, new_n7268_, new_n7269_, new_n7270_, new_n7271_,
    new_n7272_, new_n7273_, new_n7274_, new_n7275_, new_n7276_, new_n7277_,
    new_n7278_, new_n7279_, new_n7280_, new_n7281_, new_n7282_, new_n7283_,
    new_n7284_, new_n7285_, new_n7286_, new_n7287_, new_n7288_, new_n7289_,
    new_n7290_, new_n7291_, new_n7292_, new_n7293_, new_n7294_, new_n7295_,
    new_n7296_, new_n7297_, new_n7298_, new_n7299_, new_n7300_, new_n7301_,
    new_n7302_, new_n7303_, new_n7304_, new_n7305_, new_n7306_, new_n7307_,
    new_n7308_, new_n7309_, new_n7310_, new_n7311_, new_n7312_, new_n7313_,
    new_n7314_, new_n7315_, new_n7316_, new_n7317_, new_n7318_, new_n7319_,
    new_n7320_, new_n7321_, new_n7322_, new_n7323_, new_n7324_, new_n7325_,
    new_n7326_, new_n7327_, new_n7328_, new_n7329_, new_n7330_, new_n7331_,
    new_n7332_, new_n7333_, new_n7334_, new_n7335_, new_n7336_, new_n7337_,
    new_n7338_, new_n7339_, new_n7340_, new_n7341_, new_n7342_, new_n7343_,
    new_n7344_, new_n7345_, new_n7346_, new_n7347_, new_n7348_, new_n7349_,
    new_n7350_, new_n7351_, new_n7353_, new_n7354_, new_n7355_, new_n7356_,
    new_n7357_, new_n7358_, new_n7359_, new_n7360_, new_n7361_, new_n7362_,
    new_n7363_, new_n7364_, new_n7365_, new_n7366_, new_n7367_, new_n7368_,
    new_n7369_, new_n7370_, new_n7371_, new_n7372_, new_n7373_, new_n7374_,
    new_n7375_, new_n7376_, new_n7377_, new_n7378_, new_n7379_, new_n7380_,
    new_n7381_, new_n7382_, new_n7383_, new_n7384_, new_n7385_, new_n7386_,
    new_n7387_, new_n7388_, new_n7389_, new_n7390_, new_n7391_, new_n7392_,
    new_n7393_, new_n7394_, new_n7395_, new_n7396_, new_n7397_, new_n7398_,
    new_n7399_, new_n7400_, new_n7401_, new_n7402_, new_n7403_, new_n7404_,
    new_n7405_, new_n7406_, new_n7407_, new_n7408_, new_n7409_, new_n7410_,
    new_n7411_, new_n7412_, new_n7413_, new_n7414_, new_n7415_, new_n7416_,
    new_n7417_, new_n7418_, new_n7419_, new_n7420_, new_n7421_, new_n7422_,
    new_n7423_, new_n7424_, new_n7425_, new_n7426_, new_n7427_, new_n7428_,
    new_n7429_, new_n7430_, new_n7431_, new_n7432_, new_n7433_, new_n7434_,
    new_n7435_, new_n7436_, new_n7437_, new_n7438_, new_n7439_, new_n7440_,
    new_n7441_, new_n7442_, new_n7443_, new_n7444_, new_n7445_, new_n7446_,
    new_n7447_, new_n7448_, new_n7449_, new_n7450_, new_n7451_, new_n7452_,
    new_n7453_, new_n7454_, new_n7455_, new_n7456_, new_n7457_, new_n7458_,
    new_n7459_, new_n7460_, new_n7461_, new_n7462_, new_n7463_, new_n7464_,
    new_n7465_, new_n7466_, new_n7467_, new_n7468_, new_n7469_, new_n7470_,
    new_n7471_, new_n7472_, new_n7473_, new_n7474_, new_n7475_, new_n7476_,
    new_n7477_, new_n7478_, new_n7479_, new_n7480_, new_n7481_, new_n7482_,
    new_n7483_, new_n7484_, new_n7485_, new_n7486_, new_n7487_, new_n7488_,
    new_n7489_, new_n7490_, new_n7491_, new_n7492_, new_n7493_, new_n7494_,
    new_n7495_, new_n7496_, new_n7497_, new_n7498_, new_n7499_, new_n7500_,
    new_n7501_, new_n7502_, new_n7503_, new_n7504_, new_n7505_, new_n7506_,
    new_n7507_, new_n7508_, new_n7509_, new_n7510_, new_n7511_, new_n7512_,
    new_n7513_, new_n7514_, new_n7515_, new_n7516_, new_n7517_, new_n7518_,
    new_n7519_, new_n7520_, new_n7521_, new_n7522_, new_n7523_, new_n7524_,
    new_n7525_, new_n7526_, new_n7527_, new_n7528_, new_n7529_, new_n7530_,
    new_n7531_, new_n7532_, new_n7533_, new_n7534_, new_n7535_, new_n7536_,
    new_n7537_, new_n7538_, new_n7539_, new_n7540_, new_n7541_, new_n7542_,
    new_n7543_, new_n7544_, new_n7545_, new_n7546_, new_n7547_, new_n7548_,
    new_n7549_, new_n7550_, new_n7551_, new_n7552_, new_n7553_, new_n7554_,
    new_n7555_, new_n7556_, new_n7557_, new_n7558_, new_n7559_, new_n7560_,
    new_n7561_, new_n7562_, new_n7563_, new_n7564_, new_n7565_, new_n7567_,
    new_n7568_, new_n7569_, new_n7570_, new_n7571_, new_n7572_, new_n7573_,
    new_n7574_, new_n7575_, new_n7576_, new_n7577_, new_n7578_, new_n7579_,
    new_n7580_, new_n7581_, new_n7582_, new_n7583_, new_n7584_, new_n7585_,
    new_n7586_, new_n7587_, new_n7588_, new_n7589_, new_n7590_, new_n7591_,
    new_n7592_, new_n7593_, new_n7594_, new_n7595_, new_n7596_, new_n7597_,
    new_n7598_, new_n7599_, new_n7600_, new_n7601_, new_n7602_, new_n7603_,
    new_n7604_, new_n7605_, new_n7606_, new_n7607_, new_n7608_, new_n7609_,
    new_n7610_, new_n7611_, new_n7612_, new_n7613_, new_n7614_, new_n7615_,
    new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_, new_n7621_,
    new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_, new_n7627_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7681_,
    new_n7682_, new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_,
    new_n7688_, new_n7689_, new_n7690_, new_n7691_, new_n7692_, new_n7693_,
    new_n7694_, new_n7695_, new_n7696_, new_n7697_, new_n7698_, new_n7699_,
    new_n7700_, new_n7701_, new_n7702_, new_n7703_, new_n7704_, new_n7705_,
    new_n7706_, new_n7707_, new_n7708_, new_n7709_, new_n7710_, new_n7711_,
    new_n7712_, new_n7713_, new_n7714_, new_n7715_, new_n7716_, new_n7717_,
    new_n7718_, new_n7719_, new_n7720_, new_n7721_, new_n7722_, new_n7723_,
    new_n7724_, new_n7725_, new_n7726_, new_n7727_, new_n7728_, new_n7729_,
    new_n7730_, new_n7731_, new_n7732_, new_n7733_, new_n7734_, new_n7735_,
    new_n7736_, new_n7737_, new_n7738_, new_n7739_, new_n7740_, new_n7741_,
    new_n7742_, new_n7743_, new_n7744_, new_n7745_, new_n7746_, new_n7747_,
    new_n7748_, new_n7749_, new_n7750_, new_n7751_, new_n7752_, new_n7753_,
    new_n7754_, new_n7755_, new_n7756_, new_n7757_, new_n7758_, new_n7759_,
    new_n7760_, new_n7761_, new_n7763_, new_n7764_, new_n7765_, new_n7766_,
    new_n7767_, new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_,
    new_n7773_, new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_,
    new_n7779_, new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_,
    new_n7785_, new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_,
    new_n7791_, new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_,
    new_n7797_, new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_,
    new_n7803_, new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_,
    new_n7809_, new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_,
    new_n7815_, new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_,
    new_n7821_, new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_,
    new_n7827_, new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_,
    new_n7833_, new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_,
    new_n7839_, new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_,
    new_n7845_, new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_,
    new_n7851_, new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_,
    new_n7857_, new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_,
    new_n7863_, new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_,
    new_n7869_, new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_,
    new_n7875_, new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_,
    new_n7881_, new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_,
    new_n7887_, new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_,
    new_n7893_, new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_,
    new_n7899_, new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_,
    new_n7905_, new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_,
    new_n7911_, new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_,
    new_n7917_, new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_,
    new_n7923_, new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_,
    new_n7929_, new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_,
    new_n7935_, new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_,
    new_n7941_, new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_,
    new_n7947_, new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_,
    new_n7953_, new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_,
    new_n7959_, new_n7960_, new_n7961_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_,
    new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_,
    new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_,
    new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_,
    new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_,
    new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_,
    new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_,
    new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_,
    new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_,
    new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_,
    new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_,
    new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_,
    new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_,
    new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_,
    new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_,
    new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_,
    new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_,
    new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_,
    new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_,
    new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_,
    new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_,
    new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_,
    new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_,
    new_n8170_, new_n8171_, new_n8172_, new_n8174_, new_n8175_, new_n8176_,
    new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_, new_n8182_,
    new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_, new_n8188_,
    new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_, new_n8194_,
    new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_, new_n8200_,
    new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_, new_n8206_,
    new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_, new_n8212_,
    new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_, new_n8218_,
    new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_,
    new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_, new_n8230_,
    new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_, new_n8236_,
    new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_, new_n8242_,
    new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_, new_n8248_,
    new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_, new_n8254_,
    new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_, new_n8260_,
    new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_, new_n8266_,
    new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_, new_n8272_,
    new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_, new_n8278_,
    new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_, new_n8284_,
    new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_, new_n8290_,
    new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_, new_n8296_,
    new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_, new_n8302_,
    new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_, new_n8308_,
    new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_, new_n8314_,
    new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_, new_n8320_,
    new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_, new_n8326_,
    new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_, new_n8332_,
    new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_, new_n8338_,
    new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_, new_n8344_,
    new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_, new_n8350_,
    new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8364_, new_n8365_, new_n8366_, new_n8367_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8374_, new_n8375_,
    new_n8376_, new_n8377_, new_n8378_, new_n8379_, new_n8380_, new_n8381_,
    new_n8382_, new_n8383_, new_n8384_, new_n8385_, new_n8386_, new_n8387_,
    new_n8388_, new_n8389_, new_n8390_, new_n8391_, new_n8392_, new_n8393_,
    new_n8394_, new_n8395_, new_n8396_, new_n8397_, new_n8398_, new_n8399_,
    new_n8400_, new_n8401_, new_n8402_, new_n8403_, new_n8404_, new_n8405_,
    new_n8406_, new_n8407_, new_n8408_, new_n8409_, new_n8410_, new_n8411_,
    new_n8412_, new_n8413_, new_n8414_, new_n8415_, new_n8416_, new_n8417_,
    new_n8418_, new_n8419_, new_n8420_, new_n8421_, new_n8422_, new_n8423_,
    new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_, new_n8429_,
    new_n8430_, new_n8431_, new_n8432_, new_n8433_, new_n8434_, new_n8435_,
    new_n8436_, new_n8437_, new_n8438_, new_n8439_, new_n8440_, new_n8441_,
    new_n8442_, new_n8443_, new_n8444_, new_n8445_, new_n8446_, new_n8447_,
    new_n8448_, new_n8449_, new_n8450_, new_n8451_, new_n8452_, new_n8453_,
    new_n8454_, new_n8455_, new_n8456_, new_n8457_, new_n8458_, new_n8459_,
    new_n8460_, new_n8461_, new_n8462_, new_n8463_, new_n8464_, new_n8465_,
    new_n8466_, new_n8467_, new_n8468_, new_n8469_, new_n8470_, new_n8471_,
    new_n8472_, new_n8473_, new_n8474_, new_n8475_, new_n8476_, new_n8477_,
    new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_, new_n8483_,
    new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8488_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8497_, new_n8498_, new_n8499_, new_n8500_, new_n8501_,
    new_n8502_, new_n8503_, new_n8504_, new_n8505_, new_n8506_, new_n8507_,
    new_n8508_, new_n8509_, new_n8510_, new_n8511_, new_n8512_, new_n8513_,
    new_n8514_, new_n8515_, new_n8516_, new_n8517_, new_n8518_, new_n8519_,
    new_n8520_, new_n8521_, new_n8522_, new_n8523_, new_n8524_, new_n8525_,
    new_n8526_, new_n8527_, new_n8528_, new_n8529_, new_n8530_, new_n8531_,
    new_n8532_, new_n8533_, new_n8534_, new_n8535_, new_n8536_, new_n8537_,
    new_n8538_, new_n8539_, new_n8540_, new_n8541_, new_n8542_, new_n8543_,
    new_n8544_, new_n8545_, new_n8546_, new_n8547_, new_n8548_, new_n8549_,
    new_n8550_, new_n8551_, new_n8552_, new_n8553_, new_n8554_, new_n8555_,
    new_n8556_, new_n8557_, new_n8558_, new_n8559_, new_n8560_, new_n8561_,
    new_n8562_, new_n8563_, new_n8564_, new_n8565_, new_n8566_, new_n8567_,
    new_n8568_, new_n8569_, new_n8570_, new_n8572_, new_n8573_, new_n8574_,
    new_n8575_, new_n8576_, new_n8577_, new_n8578_, new_n8579_, new_n8580_,
    new_n8581_, new_n8582_, new_n8583_, new_n8584_, new_n8585_, new_n8586_,
    new_n8587_, new_n8588_, new_n8589_, new_n8590_, new_n8591_, new_n8592_,
    new_n8593_, new_n8594_, new_n8595_, new_n8596_, new_n8597_, new_n8598_,
    new_n8599_, new_n8600_, new_n8601_, new_n8602_, new_n8603_, new_n8604_,
    new_n8605_, new_n8606_, new_n8607_, new_n8608_, new_n8609_, new_n8610_,
    new_n8611_, new_n8612_, new_n8613_, new_n8614_, new_n8615_, new_n8616_,
    new_n8617_, new_n8618_, new_n8619_, new_n8620_, new_n8621_, new_n8622_,
    new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_, new_n8628_,
    new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_, new_n8634_,
    new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_, new_n8640_,
    new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_, new_n8646_,
    new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_, new_n8652_,
    new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_, new_n8658_,
    new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_, new_n8664_,
    new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_, new_n8670_,
    new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_, new_n8676_,
    new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_, new_n8682_,
    new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_, new_n8688_,
    new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_, new_n8694_,
    new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_, new_n8700_,
    new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_, new_n8706_,
    new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_, new_n8712_,
    new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_, new_n8718_,
    new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_, new_n8724_,
    new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_, new_n8730_,
    new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_, new_n8736_,
    new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_, new_n8742_,
    new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_, new_n8748_,
    new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_, new_n8754_,
    new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_, new_n8760_,
    new_n8761_, new_n8762_, new_n8763_, new_n8765_, new_n8766_, new_n8767_,
    new_n8768_, new_n8769_, new_n8770_, new_n8771_, new_n8772_, new_n8773_,
    new_n8774_, new_n8775_, new_n8776_, new_n8777_, new_n8778_, new_n8779_,
    new_n8780_, new_n8781_, new_n8782_, new_n8783_, new_n8784_, new_n8785_,
    new_n8786_, new_n8787_, new_n8788_, new_n8789_, new_n8790_, new_n8791_,
    new_n8792_, new_n8793_, new_n8794_, new_n8795_, new_n8796_, new_n8797_,
    new_n8798_, new_n8799_, new_n8800_, new_n8801_, new_n8802_, new_n8803_,
    new_n8804_, new_n8805_, new_n8806_, new_n8807_, new_n8808_, new_n8809_,
    new_n8810_, new_n8811_, new_n8812_, new_n8813_, new_n8814_, new_n8815_,
    new_n8816_, new_n8817_, new_n8818_, new_n8819_, new_n8820_, new_n8821_,
    new_n8822_, new_n8823_, new_n8824_, new_n8825_, new_n8826_, new_n8827_,
    new_n8828_, new_n8829_, new_n8830_, new_n8831_, new_n8832_, new_n8833_,
    new_n8834_, new_n8835_, new_n8836_, new_n8837_, new_n8838_, new_n8839_,
    new_n8840_, new_n8841_, new_n8842_, new_n8843_, new_n8844_, new_n8845_,
    new_n8846_, new_n8847_, new_n8848_, new_n8849_, new_n8850_, new_n8851_,
    new_n8852_, new_n8853_, new_n8854_, new_n8855_, new_n8856_, new_n8857_,
    new_n8858_, new_n8859_, new_n8860_, new_n8861_, new_n8862_, new_n8863_,
    new_n8864_, new_n8865_, new_n8866_, new_n8867_, new_n8868_, new_n8869_,
    new_n8870_, new_n8871_, new_n8872_, new_n8873_, new_n8874_, new_n8875_,
    new_n8876_, new_n8877_, new_n8878_, new_n8879_, new_n8880_, new_n8881_,
    new_n8882_, new_n8883_, new_n8884_, new_n8885_, new_n8886_, new_n8887_,
    new_n8888_, new_n8889_, new_n8890_, new_n8891_, new_n8892_, new_n8893_,
    new_n8894_, new_n8895_, new_n8896_, new_n8897_, new_n8898_, new_n8899_,
    new_n8900_, new_n8901_, new_n8902_, new_n8903_, new_n8904_, new_n8905_,
    new_n8906_, new_n8907_, new_n8908_, new_n8909_, new_n8910_, new_n8911_,
    new_n8912_, new_n8913_, new_n8914_, new_n8915_, new_n8916_, new_n8917_,
    new_n8918_, new_n8919_, new_n8920_, new_n8921_, new_n8922_, new_n8923_,
    new_n8924_, new_n8925_, new_n8926_, new_n8927_, new_n8928_, new_n8929_,
    new_n8930_, new_n8931_, new_n8932_, new_n8933_, new_n8934_, new_n8935_,
    new_n8936_, new_n8937_, new_n8938_, new_n8939_, new_n8940_, new_n8941_,
    new_n8942_, new_n8943_, new_n8944_, new_n8945_, new_n8946_, new_n8947_,
    new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_, new_n8953_,
    new_n8954_, new_n8955_, new_n8957_, new_n8958_, new_n8959_, new_n8960_,
    new_n8961_, new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_,
    new_n8967_, new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_,
    new_n8973_, new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_,
    new_n8979_, new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_,
    new_n8985_, new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_,
    new_n8991_, new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_,
    new_n8997_, new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_,
    new_n9003_, new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_,
    new_n9009_, new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_,
    new_n9015_, new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_,
    new_n9021_, new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_,
    new_n9027_, new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_,
    new_n9033_, new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_,
    new_n9039_, new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_,
    new_n9045_, new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_,
    new_n9051_, new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_,
    new_n9057_, new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_,
    new_n9063_, new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_,
    new_n9069_, new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_,
    new_n9075_, new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_,
    new_n9081_, new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_,
    new_n9087_, new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_,
    new_n9093_, new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_,
    new_n9099_, new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_,
    new_n9105_, new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_,
    new_n9111_, new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_,
    new_n9117_, new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_,
    new_n9123_, new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_,
    new_n9129_, new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_,
    new_n9135_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_,
    new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_,
    new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_,
    new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_,
    new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_,
    new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_,
    new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_,
    new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9331_, new_n9332_, new_n9333_, new_n9334_,
    new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_, new_n9340_,
    new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_, new_n9346_,
    new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_, new_n9352_,
    new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_, new_n9358_,
    new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_, new_n9364_,
    new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_, new_n9370_,
    new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_, new_n9376_,
    new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_, new_n9382_,
    new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_, new_n9388_,
    new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_, new_n9394_,
    new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_, new_n9400_,
    new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_, new_n9406_,
    new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_, new_n9412_,
    new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_, new_n9418_,
    new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_, new_n9424_,
    new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_, new_n9430_,
    new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_, new_n9436_,
    new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_, new_n9442_,
    new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_, new_n9454_,
    new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_, new_n9460_,
    new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_, new_n9466_,
    new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_, new_n9472_,
    new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_, new_n9478_,
    new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_, new_n9484_,
    new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9490_,
    new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_, new_n9496_,
    new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_, new_n9502_,
    new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9508_, new_n9509_,
    new_n9510_, new_n9511_, new_n9512_, new_n9513_, new_n9514_, new_n9515_,
    new_n9516_, new_n9517_, new_n9518_, new_n9519_, new_n9520_, new_n9521_,
    new_n9522_, new_n9523_, new_n9524_, new_n9525_, new_n9526_, new_n9527_,
    new_n9528_, new_n9529_, new_n9530_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9535_, new_n9536_, new_n9537_, new_n9538_, new_n9539_,
    new_n9540_, new_n9541_, new_n9542_, new_n9543_, new_n9544_, new_n9545_,
    new_n9546_, new_n9547_, new_n9548_, new_n9549_, new_n9550_, new_n9551_,
    new_n9552_, new_n9553_, new_n9554_, new_n9555_, new_n9556_, new_n9557_,
    new_n9558_, new_n9559_, new_n9560_, new_n9561_, new_n9562_, new_n9563_,
    new_n9564_, new_n9565_, new_n9566_, new_n9567_, new_n9568_, new_n9569_,
    new_n9570_, new_n9571_, new_n9572_, new_n9573_, new_n9574_, new_n9575_,
    new_n9576_, new_n9577_, new_n9578_, new_n9579_, new_n9580_, new_n9581_,
    new_n9582_, new_n9583_, new_n9584_, new_n9585_, new_n9586_, new_n9587_,
    new_n9588_, new_n9589_, new_n9590_, new_n9591_, new_n9592_, new_n9593_,
    new_n9594_, new_n9595_, new_n9596_, new_n9597_, new_n9598_, new_n9599_,
    new_n9600_, new_n9601_, new_n9602_, new_n9603_, new_n9604_, new_n9605_,
    new_n9606_, new_n9607_, new_n9608_, new_n9609_, new_n9610_, new_n9611_,
    new_n9612_, new_n9613_, new_n9614_, new_n9615_, new_n9616_, new_n9617_,
    new_n9618_, new_n9619_, new_n9620_, new_n9621_, new_n9622_, new_n9623_,
    new_n9624_, new_n9625_, new_n9626_, new_n9627_, new_n9628_, new_n9629_,
    new_n9630_, new_n9631_, new_n9632_, new_n9633_, new_n9634_, new_n9635_,
    new_n9636_, new_n9637_, new_n9638_, new_n9639_, new_n9640_, new_n9641_,
    new_n9642_, new_n9643_, new_n9644_, new_n9645_, new_n9646_, new_n9647_,
    new_n9648_, new_n9649_, new_n9650_, new_n9651_, new_n9652_, new_n9653_,
    new_n9654_, new_n9655_, new_n9656_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9662_, new_n9663_, new_n9664_, new_n9665_,
    new_n9666_, new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_,
    new_n9672_, new_n9673_, new_n9674_, new_n9675_, new_n9676_, new_n9677_,
    new_n9678_, new_n9679_, new_n9680_, new_n9681_, new_n9682_, new_n9683_,
    new_n9684_, new_n9685_, new_n9687_, new_n9688_, new_n9689_, new_n9690_,
    new_n9691_, new_n9692_, new_n9693_, new_n9694_, new_n9695_, new_n9696_,
    new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_, new_n9702_,
    new_n9703_, new_n9704_, new_n9705_, new_n9706_, new_n9707_, new_n9708_,
    new_n9709_, new_n9710_, new_n9711_, new_n9712_, new_n9713_, new_n9714_,
    new_n9715_, new_n9716_, new_n9717_, new_n9718_, new_n9719_, new_n9720_,
    new_n9721_, new_n9722_, new_n9723_, new_n9724_, new_n9725_, new_n9726_,
    new_n9727_, new_n9728_, new_n9729_, new_n9730_, new_n9731_, new_n9732_,
    new_n9733_, new_n9734_, new_n9735_, new_n9736_, new_n9737_, new_n9738_,
    new_n9739_, new_n9740_, new_n9741_, new_n9742_, new_n9743_, new_n9744_,
    new_n9745_, new_n9746_, new_n9747_, new_n9748_, new_n9749_, new_n9750_,
    new_n9751_, new_n9752_, new_n9753_, new_n9754_, new_n9755_, new_n9756_,
    new_n9757_, new_n9758_, new_n9759_, new_n9760_, new_n9761_, new_n9762_,
    new_n9763_, new_n9764_, new_n9765_, new_n9766_, new_n9767_, new_n9768_,
    new_n9769_, new_n9770_, new_n9771_, new_n9772_, new_n9773_, new_n9774_,
    new_n9775_, new_n9776_, new_n9777_, new_n9778_, new_n9779_, new_n9780_,
    new_n9781_, new_n9782_, new_n9783_, new_n9784_, new_n9785_, new_n9786_,
    new_n9787_, new_n9788_, new_n9789_, new_n9790_, new_n9791_, new_n9792_,
    new_n9793_, new_n9794_, new_n9795_, new_n9796_, new_n9797_, new_n9798_,
    new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_, new_n9804_,
    new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_, new_n9810_,
    new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_, new_n9816_,
    new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_, new_n9822_,
    new_n9823_, new_n9824_, new_n9825_, new_n9826_, new_n9827_, new_n9828_,
    new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_,
    new_n9835_, new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_,
    new_n9841_, new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_,
    new_n9847_, new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_,
    new_n9853_, new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10026_, new_n10027_,
    new_n10028_, new_n10029_, new_n10030_, new_n10031_, new_n10032_,
    new_n10033_, new_n10034_, new_n10036_, new_n10037_, new_n10038_,
    new_n10039_, new_n10040_, new_n10041_, new_n10042_, new_n10043_,
    new_n10044_, new_n10045_, new_n10046_, new_n10047_, new_n10048_,
    new_n10049_, new_n10050_, new_n10051_, new_n10052_, new_n10053_,
    new_n10054_, new_n10055_, new_n10056_, new_n10057_, new_n10058_,
    new_n10059_, new_n10060_, new_n10061_, new_n10062_, new_n10063_,
    new_n10064_, new_n10065_, new_n10066_, new_n10067_, new_n10068_,
    new_n10069_, new_n10070_, new_n10071_, new_n10072_, new_n10073_,
    new_n10074_, new_n10075_, new_n10076_, new_n10077_, new_n10078_,
    new_n10079_, new_n10080_, new_n10081_, new_n10082_, new_n10083_,
    new_n10084_, new_n10085_, new_n10086_, new_n10087_, new_n10088_,
    new_n10089_, new_n10090_, new_n10091_, new_n10092_, new_n10093_,
    new_n10094_, new_n10095_, new_n10096_, new_n10097_, new_n10098_,
    new_n10099_, new_n10100_, new_n10101_, new_n10102_, new_n10103_,
    new_n10104_, new_n10105_, new_n10106_, new_n10107_, new_n10108_,
    new_n10109_, new_n10110_, new_n10111_, new_n10112_, new_n10113_,
    new_n10114_, new_n10115_, new_n10116_, new_n10117_, new_n10118_,
    new_n10119_, new_n10120_, new_n10121_, new_n10122_, new_n10123_,
    new_n10124_, new_n10125_, new_n10126_, new_n10127_, new_n10128_,
    new_n10129_, new_n10130_, new_n10131_, new_n10132_, new_n10133_,
    new_n10134_, new_n10135_, new_n10136_, new_n10137_, new_n10138_,
    new_n10139_, new_n10140_, new_n10141_, new_n10142_, new_n10143_,
    new_n10144_, new_n10145_, new_n10146_, new_n10147_, new_n10148_,
    new_n10149_, new_n10150_, new_n10151_, new_n10152_, new_n10153_,
    new_n10154_, new_n10155_, new_n10156_, new_n10157_, new_n10158_,
    new_n10159_, new_n10160_, new_n10161_, new_n10162_, new_n10163_,
    new_n10164_, new_n10165_, new_n10166_, new_n10167_, new_n10168_,
    new_n10169_, new_n10170_, new_n10171_, new_n10172_, new_n10173_,
    new_n10174_, new_n10175_, new_n10176_, new_n10177_, new_n10178_,
    new_n10179_, new_n10180_, new_n10181_, new_n10182_, new_n10183_,
    new_n10184_, new_n10185_, new_n10186_, new_n10187_, new_n10188_,
    new_n10189_, new_n10190_, new_n10191_, new_n10192_, new_n10193_,
    new_n10194_, new_n10195_, new_n10196_, new_n10197_, new_n10198_,
    new_n10199_, new_n10200_, new_n10201_, new_n10202_, new_n10203_,
    new_n10204_, new_n10205_, new_n10206_, new_n10207_, new_n10208_,
    new_n10209_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10541_,
    new_n10542_, new_n10543_, new_n10544_, new_n10545_, new_n10546_,
    new_n10547_, new_n10548_, new_n10549_, new_n10550_, new_n10551_,
    new_n10552_, new_n10553_, new_n10554_, new_n10555_, new_n10556_,
    new_n10557_, new_n10558_, new_n10559_, new_n10560_, new_n10561_,
    new_n10562_, new_n10563_, new_n10564_, new_n10565_, new_n10566_,
    new_n10567_, new_n10568_, new_n10569_, new_n10570_, new_n10571_,
    new_n10572_, new_n10573_, new_n10574_, new_n10575_, new_n10576_,
    new_n10577_, new_n10578_, new_n10579_, new_n10580_, new_n10581_,
    new_n10582_, new_n10583_, new_n10584_, new_n10585_, new_n10586_,
    new_n10587_, new_n10588_, new_n10589_, new_n10590_, new_n10591_,
    new_n10592_, new_n10593_, new_n10594_, new_n10595_, new_n10596_,
    new_n10597_, new_n10598_, new_n10599_, new_n10600_, new_n10601_,
    new_n10602_, new_n10603_, new_n10604_, new_n10605_, new_n10606_,
    new_n10607_, new_n10608_, new_n10609_, new_n10610_, new_n10611_,
    new_n10612_, new_n10613_, new_n10614_, new_n10615_, new_n10616_,
    new_n10617_, new_n10618_, new_n10619_, new_n10620_, new_n10621_,
    new_n10622_, new_n10623_, new_n10624_, new_n10625_, new_n10626_,
    new_n10627_, new_n10628_, new_n10629_, new_n10630_, new_n10631_,
    new_n10632_, new_n10633_, new_n10634_, new_n10635_, new_n10636_,
    new_n10637_, new_n10638_, new_n10639_, new_n10640_, new_n10641_,
    new_n10642_, new_n10643_, new_n10644_, new_n10645_, new_n10646_,
    new_n10647_, new_n10648_, new_n10649_, new_n10650_, new_n10651_,
    new_n10652_, new_n10653_, new_n10654_, new_n10655_, new_n10656_,
    new_n10657_, new_n10658_, new_n10659_, new_n10660_, new_n10661_,
    new_n10662_, new_n10663_, new_n10664_, new_n10665_, new_n10666_,
    new_n10667_, new_n10668_, new_n10669_, new_n10670_, new_n10671_,
    new_n10672_, new_n10673_, new_n10674_, new_n10675_, new_n10676_,
    new_n10677_, new_n10678_, new_n10679_, new_n10680_, new_n10681_,
    new_n10682_, new_n10683_, new_n10684_, new_n10685_, new_n10686_,
    new_n10687_, new_n10688_, new_n10689_, new_n10690_, new_n10691_,
    new_n10692_, new_n10693_, new_n10694_, new_n10695_, new_n10696_,
    new_n10697_, new_n10698_, new_n10699_, new_n10700_, new_n10702_,
    new_n10703_, new_n10704_, new_n10705_, new_n10706_, new_n10707_,
    new_n10708_, new_n10709_, new_n10710_, new_n10711_, new_n10712_,
    new_n10713_, new_n10714_, new_n10715_, new_n10716_, new_n10717_,
    new_n10718_, new_n10719_, new_n10720_, new_n10721_, new_n10722_,
    new_n10723_, new_n10724_, new_n10725_, new_n10726_, new_n10727_,
    new_n10728_, new_n10729_, new_n10730_, new_n10731_, new_n10732_,
    new_n10733_, new_n10734_, new_n10735_, new_n10736_, new_n10737_,
    new_n10738_, new_n10739_, new_n10740_, new_n10741_, new_n10742_,
    new_n10743_, new_n10744_, new_n10745_, new_n10746_, new_n10747_,
    new_n10748_, new_n10749_, new_n10750_, new_n10751_, new_n10752_,
    new_n10753_, new_n10754_, new_n10755_, new_n10756_, new_n10757_,
    new_n10758_, new_n10759_, new_n10760_, new_n10761_, new_n10762_,
    new_n10763_, new_n10764_, new_n10765_, new_n10766_, new_n10767_,
    new_n10768_, new_n10769_, new_n10770_, new_n10771_, new_n10772_,
    new_n10773_, new_n10774_, new_n10775_, new_n10776_, new_n10777_,
    new_n10778_, new_n10779_, new_n10780_, new_n10781_, new_n10782_,
    new_n10783_, new_n10784_, new_n10785_, new_n10786_, new_n10787_,
    new_n10788_, new_n10789_, new_n10790_, new_n10791_, new_n10792_,
    new_n10793_, new_n10794_, new_n10795_, new_n10796_, new_n10797_,
    new_n10798_, new_n10799_, new_n10800_, new_n10801_, new_n10802_,
    new_n10803_, new_n10804_, new_n10805_, new_n10806_, new_n10807_,
    new_n10808_, new_n10809_, new_n10810_, new_n10811_, new_n10812_,
    new_n10813_, new_n10814_, new_n10815_, new_n10816_, new_n10817_,
    new_n10818_, new_n10819_, new_n10820_, new_n10821_, new_n10822_,
    new_n10823_, new_n10824_, new_n10825_, new_n10826_, new_n10827_,
    new_n10828_, new_n10829_, new_n10830_, new_n10831_, new_n10832_,
    new_n10833_, new_n10834_, new_n10835_, new_n10836_, new_n10837_,
    new_n10838_, new_n10839_, new_n10840_, new_n10841_, new_n10842_,
    new_n10843_, new_n10844_, new_n10845_, new_n10846_, new_n10847_,
    new_n10848_, new_n10849_, new_n10850_, new_n10851_, new_n10852_,
    new_n10853_, new_n10854_, new_n10855_, new_n10856_, new_n10857_,
    new_n10859_, new_n10860_, new_n10861_, new_n10862_, new_n10863_,
    new_n10864_, new_n10865_, new_n10866_, new_n10867_, new_n10868_,
    new_n10869_, new_n10870_, new_n10871_, new_n10872_, new_n10873_,
    new_n10874_, new_n10875_, new_n10876_, new_n10877_, new_n10878_,
    new_n10879_, new_n10880_, new_n10881_, new_n10882_, new_n10883_,
    new_n10884_, new_n10885_, new_n10886_, new_n10887_, new_n10888_,
    new_n10889_, new_n10890_, new_n10891_, new_n10892_, new_n10893_,
    new_n10894_, new_n10895_, new_n10896_, new_n10897_, new_n10898_,
    new_n10899_, new_n10900_, new_n10901_, new_n10902_, new_n10903_,
    new_n10904_, new_n10905_, new_n10906_, new_n10907_, new_n10908_,
    new_n10909_, new_n10910_, new_n10911_, new_n10912_, new_n10913_,
    new_n10914_, new_n10915_, new_n10916_, new_n10917_, new_n10918_,
    new_n10919_, new_n10920_, new_n10921_, new_n10922_, new_n10923_,
    new_n10924_, new_n10925_, new_n10926_, new_n10927_, new_n10928_,
    new_n10929_, new_n10930_, new_n10931_, new_n10932_, new_n10933_,
    new_n10934_, new_n10935_, new_n10936_, new_n10937_, new_n10938_,
    new_n10939_, new_n10940_, new_n10941_, new_n10942_, new_n10943_,
    new_n10944_, new_n10945_, new_n10946_, new_n10947_, new_n10948_,
    new_n10949_, new_n10950_, new_n10951_, new_n10952_, new_n10953_,
    new_n10954_, new_n10955_, new_n10956_, new_n10957_, new_n10958_,
    new_n10959_, new_n10960_, new_n10961_, new_n10962_, new_n10963_,
    new_n10964_, new_n10965_, new_n10966_, new_n10967_, new_n10968_,
    new_n10969_, new_n10970_, new_n10971_, new_n10972_, new_n10973_,
    new_n10974_, new_n10975_, new_n10976_, new_n10977_, new_n10978_,
    new_n10979_, new_n10980_, new_n10981_, new_n10982_, new_n10983_,
    new_n10984_, new_n10985_, new_n10986_, new_n10987_, new_n10988_,
    new_n10989_, new_n10990_, new_n10991_, new_n10992_, new_n10993_,
    new_n10994_, new_n10995_, new_n10996_, new_n10997_, new_n10998_,
    new_n10999_, new_n11000_, new_n11001_, new_n11002_, new_n11003_,
    new_n11004_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11050_, new_n11051_, new_n11052_, new_n11053_, new_n11054_,
    new_n11055_, new_n11056_, new_n11057_, new_n11058_, new_n11059_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11073_, new_n11074_,
    new_n11075_, new_n11076_, new_n11077_, new_n11078_, new_n11079_,
    new_n11080_, new_n11081_, new_n11082_, new_n11083_, new_n11084_,
    new_n11085_, new_n11086_, new_n11087_, new_n11088_, new_n11089_,
    new_n11090_, new_n11091_, new_n11092_, new_n11093_, new_n11094_,
    new_n11095_, new_n11096_, new_n11097_, new_n11098_, new_n11099_,
    new_n11100_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11106_, new_n11107_, new_n11108_, new_n11109_,
    new_n11110_, new_n11111_, new_n11112_, new_n11113_, new_n11114_,
    new_n11115_, new_n11116_, new_n11117_, new_n11118_, new_n11119_,
    new_n11120_, new_n11121_, new_n11122_, new_n11123_, new_n11124_,
    new_n11125_, new_n11126_, new_n11127_, new_n11128_, new_n11129_,
    new_n11130_, new_n11131_, new_n11132_, new_n11133_, new_n11134_,
    new_n11135_, new_n11136_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11146_, new_n11147_, new_n11148_, new_n11149_,
    new_n11150_, new_n11151_, new_n11152_, new_n11153_, new_n11154_,
    new_n11155_, new_n11156_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11166_, new_n11167_, new_n11168_, new_n11169_, new_n11170_,
    new_n11171_, new_n11172_, new_n11173_, new_n11174_, new_n11175_,
    new_n11176_, new_n11177_, new_n11178_, new_n11179_, new_n11180_,
    new_n11181_, new_n11182_, new_n11183_, new_n11184_, new_n11185_,
    new_n11186_, new_n11187_, new_n11188_, new_n11189_, new_n11190_,
    new_n11191_, new_n11192_, new_n11193_, new_n11194_, new_n11195_,
    new_n11196_, new_n11197_, new_n11198_, new_n11199_, new_n11200_,
    new_n11201_, new_n11202_, new_n11203_, new_n11204_, new_n11205_,
    new_n11206_, new_n11207_, new_n11208_, new_n11209_, new_n11210_,
    new_n11211_, new_n11212_, new_n11213_, new_n11214_, new_n11215_,
    new_n11216_, new_n11217_, new_n11218_, new_n11219_, new_n11220_,
    new_n11221_, new_n11222_, new_n11223_, new_n11224_, new_n11225_,
    new_n11226_, new_n11227_, new_n11228_, new_n11229_, new_n11230_,
    new_n11231_, new_n11232_, new_n11233_, new_n11234_, new_n11235_,
    new_n11236_, new_n11237_, new_n11238_, new_n11239_, new_n11240_,
    new_n11241_, new_n11242_, new_n11243_, new_n11244_, new_n11245_,
    new_n11246_, new_n11247_, new_n11248_, new_n11249_, new_n11250_,
    new_n11251_, new_n11252_, new_n11253_, new_n11254_, new_n11255_,
    new_n11256_, new_n11257_, new_n11258_, new_n11259_, new_n11260_,
    new_n11261_, new_n11262_, new_n11263_, new_n11264_, new_n11265_,
    new_n11266_, new_n11267_, new_n11268_, new_n11269_, new_n11270_,
    new_n11271_, new_n11272_, new_n11273_, new_n11274_, new_n11275_,
    new_n11276_, new_n11277_, new_n11278_, new_n11279_, new_n11280_,
    new_n11281_, new_n11282_, new_n11283_, new_n11284_, new_n11285_,
    new_n11286_, new_n11287_, new_n11288_, new_n11289_, new_n11290_,
    new_n11291_, new_n11292_, new_n11293_, new_n11294_, new_n11295_,
    new_n11296_, new_n11298_, new_n11299_, new_n11300_, new_n11301_,
    new_n11302_, new_n11303_, new_n11304_, new_n11305_, new_n11306_,
    new_n11307_, new_n11308_, new_n11309_, new_n11310_, new_n11311_,
    new_n11312_, new_n11313_, new_n11314_, new_n11315_, new_n11316_,
    new_n11317_, new_n11318_, new_n11319_, new_n11320_, new_n11321_,
    new_n11322_, new_n11323_, new_n11324_, new_n11325_, new_n11326_,
    new_n11327_, new_n11328_, new_n11329_, new_n11330_, new_n11331_,
    new_n11332_, new_n11333_, new_n11334_, new_n11335_, new_n11336_,
    new_n11337_, new_n11338_, new_n11339_, new_n11340_, new_n11341_,
    new_n11342_, new_n11343_, new_n11344_, new_n11345_, new_n11346_,
    new_n11347_, new_n11348_, new_n11349_, new_n11350_, new_n11351_,
    new_n11352_, new_n11353_, new_n11354_, new_n11355_, new_n11356_,
    new_n11357_, new_n11358_, new_n11359_, new_n11360_, new_n11361_,
    new_n11362_, new_n11363_, new_n11364_, new_n11365_, new_n11366_,
    new_n11367_, new_n11368_, new_n11369_, new_n11370_, new_n11371_,
    new_n11372_, new_n11373_, new_n11374_, new_n11375_, new_n11376_,
    new_n11377_, new_n11378_, new_n11379_, new_n11380_, new_n11381_,
    new_n11382_, new_n11383_, new_n11384_, new_n11385_, new_n11386_,
    new_n11387_, new_n11388_, new_n11389_, new_n11390_, new_n11391_,
    new_n11392_, new_n11393_, new_n11394_, new_n11395_, new_n11396_,
    new_n11397_, new_n11398_, new_n11399_, new_n11400_, new_n11401_,
    new_n11402_, new_n11403_, new_n11404_, new_n11405_, new_n11406_,
    new_n11407_, new_n11408_, new_n11409_, new_n11410_, new_n11411_,
    new_n11412_, new_n11413_, new_n11414_, new_n11415_, new_n11416_,
    new_n11417_, new_n11418_, new_n11419_, new_n11420_, new_n11421_,
    new_n11422_, new_n11423_, new_n11424_, new_n11425_, new_n11426_,
    new_n11427_, new_n11428_, new_n11429_, new_n11430_, new_n11431_,
    new_n11432_, new_n11433_, new_n11434_, new_n11435_, new_n11436_,
    new_n11437_, new_n11438_, new_n11439_, new_n11441_, new_n11442_,
    new_n11443_, new_n11444_, new_n11445_, new_n11446_, new_n11447_,
    new_n11448_, new_n11449_, new_n11450_, new_n11451_, new_n11452_,
    new_n11453_, new_n11454_, new_n11455_, new_n11456_, new_n11457_,
    new_n11458_, new_n11459_, new_n11460_, new_n11461_, new_n11462_,
    new_n11463_, new_n11464_, new_n11465_, new_n11466_, new_n11467_,
    new_n11468_, new_n11469_, new_n11470_, new_n11471_, new_n11472_,
    new_n11473_, new_n11474_, new_n11475_, new_n11476_, new_n11477_,
    new_n11478_, new_n11479_, new_n11480_, new_n11481_, new_n11482_,
    new_n11483_, new_n11484_, new_n11485_, new_n11486_, new_n11487_,
    new_n11488_, new_n11489_, new_n11490_, new_n11491_, new_n11492_,
    new_n11493_, new_n11494_, new_n11495_, new_n11496_, new_n11497_,
    new_n11498_, new_n11499_, new_n11500_, new_n11501_, new_n11502_,
    new_n11503_, new_n11504_, new_n11505_, new_n11506_, new_n11507_,
    new_n11508_, new_n11509_, new_n11510_, new_n11511_, new_n11512_,
    new_n11513_, new_n11514_, new_n11515_, new_n11516_, new_n11517_,
    new_n11518_, new_n11519_, new_n11520_, new_n11521_, new_n11522_,
    new_n11523_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11554_, new_n11555_, new_n11556_, new_n11557_,
    new_n11558_, new_n11559_, new_n11560_, new_n11561_, new_n11562_,
    new_n11563_, new_n11564_, new_n11565_, new_n11566_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11576_, new_n11577_, new_n11578_,
    new_n11579_, new_n11580_, new_n11581_, new_n11582_, new_n11583_,
    new_n11584_, new_n11585_, new_n11586_, new_n11587_, new_n11588_,
    new_n11589_, new_n11590_, new_n11591_, new_n11592_, new_n11593_,
    new_n11594_, new_n11595_, new_n11596_, new_n11597_, new_n11598_,
    new_n11599_, new_n11600_, new_n11601_, new_n11602_, new_n11603_,
    new_n11604_, new_n11605_, new_n11606_, new_n11607_, new_n11608_,
    new_n11609_, new_n11610_, new_n11611_, new_n11612_, new_n11613_,
    new_n11614_, new_n11615_, new_n11616_, new_n11617_, new_n11618_,
    new_n11619_, new_n11620_, new_n11621_, new_n11622_, new_n11623_,
    new_n11624_, new_n11625_, new_n11626_, new_n11627_, new_n11628_,
    new_n11629_, new_n11630_, new_n11631_, new_n11632_, new_n11633_,
    new_n11634_, new_n11635_, new_n11636_, new_n11637_, new_n11638_,
    new_n11639_, new_n11640_, new_n11641_, new_n11642_, new_n11643_,
    new_n11644_, new_n11645_, new_n11646_, new_n11647_, new_n11648_,
    new_n11649_, new_n11650_, new_n11651_, new_n11652_, new_n11653_,
    new_n11654_, new_n11655_, new_n11656_, new_n11657_, new_n11658_,
    new_n11659_, new_n11660_, new_n11661_, new_n11662_, new_n11663_,
    new_n11664_, new_n11665_, new_n11666_, new_n11667_, new_n11668_,
    new_n11669_, new_n11670_, new_n11671_, new_n11672_, new_n11673_,
    new_n11674_, new_n11675_, new_n11676_, new_n11677_, new_n11678_,
    new_n11679_, new_n11680_, new_n11681_, new_n11682_, new_n11683_,
    new_n11684_, new_n11685_, new_n11686_, new_n11687_, new_n11688_,
    new_n11689_, new_n11690_, new_n11691_, new_n11692_, new_n11693_,
    new_n11694_, new_n11695_, new_n11696_, new_n11697_, new_n11698_,
    new_n11699_, new_n11700_, new_n11701_, new_n11702_, new_n11703_,
    new_n11704_, new_n11705_, new_n11706_, new_n11707_, new_n11709_,
    new_n11710_, new_n11711_, new_n11712_, new_n11713_, new_n11714_,
    new_n11715_, new_n11716_, new_n11717_, new_n11718_, new_n11719_,
    new_n11720_, new_n11721_, new_n11722_, new_n11723_, new_n11724_,
    new_n11725_, new_n11726_, new_n11727_, new_n11728_, new_n11729_,
    new_n11730_, new_n11731_, new_n11732_, new_n11733_, new_n11734_,
    new_n11735_, new_n11736_, new_n11737_, new_n11738_, new_n11739_,
    new_n11740_, new_n11741_, new_n11742_, new_n11743_, new_n11744_,
    new_n11745_, new_n11746_, new_n11747_, new_n11748_, new_n11749_,
    new_n11750_, new_n11751_, new_n11752_, new_n11753_, new_n11754_,
    new_n11755_, new_n11756_, new_n11757_, new_n11758_, new_n11759_,
    new_n11760_, new_n11761_, new_n11762_, new_n11763_, new_n11764_,
    new_n11765_, new_n11766_, new_n11767_, new_n11768_, new_n11769_,
    new_n11770_, new_n11771_, new_n11772_, new_n11773_, new_n11774_,
    new_n11775_, new_n11776_, new_n11777_, new_n11778_, new_n11779_,
    new_n11780_, new_n11781_, new_n11782_, new_n11783_, new_n11784_,
    new_n11785_, new_n11786_, new_n11787_, new_n11788_, new_n11789_,
    new_n11790_, new_n11791_, new_n11792_, new_n11793_, new_n11794_,
    new_n11795_, new_n11796_, new_n11797_, new_n11798_, new_n11799_,
    new_n11800_, new_n11801_, new_n11802_, new_n11803_, new_n11804_,
    new_n11805_, new_n11806_, new_n11807_, new_n11808_, new_n11809_,
    new_n11810_, new_n11811_, new_n11812_, new_n11813_, new_n11814_,
    new_n11815_, new_n11816_, new_n11817_, new_n11818_, new_n11819_,
    new_n11820_, new_n11821_, new_n11822_, new_n11823_, new_n11824_,
    new_n11825_, new_n11826_, new_n11827_, new_n11828_, new_n11829_,
    new_n11830_, new_n11831_, new_n11832_, new_n11833_, new_n11834_,
    new_n11835_, new_n11836_, new_n11837_, new_n11838_, new_n11839_,
    new_n11840_, new_n11841_, new_n11842_, new_n11843_, new_n11844_,
    new_n11845_, new_n11846_, new_n11848_, new_n11849_, new_n11850_,
    new_n11851_, new_n11852_, new_n11853_, new_n11854_, new_n11855_,
    new_n11856_, new_n11857_, new_n11858_, new_n11859_, new_n11860_,
    new_n11861_, new_n11862_, new_n11863_, new_n11864_, new_n11865_,
    new_n11866_, new_n11867_, new_n11868_, new_n11869_, new_n11870_,
    new_n11871_, new_n11872_, new_n11873_, new_n11874_, new_n11875_,
    new_n11876_, new_n11877_, new_n11878_, new_n11879_, new_n11880_,
    new_n11881_, new_n11882_, new_n11883_, new_n11884_, new_n11885_,
    new_n11886_, new_n11887_, new_n11888_, new_n11889_, new_n11890_,
    new_n11891_, new_n11892_, new_n11893_, new_n11894_, new_n11895_,
    new_n11896_, new_n11897_, new_n11898_, new_n11899_, new_n11900_,
    new_n11901_, new_n11902_, new_n11903_, new_n11904_, new_n11905_,
    new_n11906_, new_n11907_, new_n11908_, new_n11909_, new_n11910_,
    new_n11911_, new_n11912_, new_n11913_, new_n11914_, new_n11915_,
    new_n11916_, new_n11917_, new_n11918_, new_n11919_, new_n11920_,
    new_n11921_, new_n11922_, new_n11923_, new_n11924_, new_n11925_,
    new_n11926_, new_n11927_, new_n11928_, new_n11929_, new_n11930_,
    new_n11931_, new_n11932_, new_n11933_, new_n11934_, new_n11935_,
    new_n11936_, new_n11937_, new_n11938_, new_n11939_, new_n11940_,
    new_n11941_, new_n11942_, new_n11943_, new_n11944_, new_n11945_,
    new_n11946_, new_n11947_, new_n11948_, new_n11949_, new_n11950_,
    new_n11951_, new_n11952_, new_n11953_, new_n11954_, new_n11955_,
    new_n11956_, new_n11957_, new_n11958_, new_n11959_, new_n11960_,
    new_n11961_, new_n11962_, new_n11963_, new_n11964_, new_n11965_,
    new_n11966_, new_n11967_, new_n11968_, new_n11969_, new_n11970_,
    new_n11971_, new_n11972_, new_n11973_, new_n11974_, new_n11975_,
    new_n11977_, new_n11978_, new_n11979_, new_n11980_, new_n11981_,
    new_n11982_, new_n11983_, new_n11984_, new_n11985_, new_n11986_,
    new_n11987_, new_n11988_, new_n11989_, new_n11990_, new_n11991_,
    new_n11992_, new_n11993_, new_n11994_, new_n11995_, new_n11996_,
    new_n11997_, new_n11998_, new_n11999_, new_n12000_, new_n12001_,
    new_n12002_, new_n12003_, new_n12004_, new_n12005_, new_n12006_,
    new_n12007_, new_n12008_, new_n12009_, new_n12010_, new_n12011_,
    new_n12012_, new_n12013_, new_n12014_, new_n12015_, new_n12016_,
    new_n12017_, new_n12018_, new_n12019_, new_n12020_, new_n12021_,
    new_n12022_, new_n12023_, new_n12024_, new_n12025_, new_n12026_,
    new_n12027_, new_n12028_, new_n12029_, new_n12030_, new_n12031_,
    new_n12032_, new_n12033_, new_n12034_, new_n12035_, new_n12036_,
    new_n12037_, new_n12038_, new_n12039_, new_n12040_, new_n12041_,
    new_n12042_, new_n12043_, new_n12044_, new_n12045_, new_n12046_,
    new_n12047_, new_n12048_, new_n12049_, new_n12050_, new_n12051_,
    new_n12052_, new_n12053_, new_n12054_, new_n12055_, new_n12056_,
    new_n12057_, new_n12058_, new_n12059_, new_n12060_, new_n12061_,
    new_n12062_, new_n12063_, new_n12064_, new_n12065_, new_n12066_,
    new_n12067_, new_n12068_, new_n12069_, new_n12070_, new_n12071_,
    new_n12072_, new_n12073_, new_n12074_, new_n12075_, new_n12076_,
    new_n12077_, new_n12078_, new_n12079_, new_n12080_, new_n12081_,
    new_n12082_, new_n12083_, new_n12084_, new_n12085_, new_n12086_,
    new_n12087_, new_n12088_, new_n12089_, new_n12090_, new_n12091_,
    new_n12092_, new_n12093_, new_n12094_, new_n12095_, new_n12096_,
    new_n12097_, new_n12098_, new_n12099_, new_n12101_, new_n12102_,
    new_n12103_, new_n12104_, new_n12105_, new_n12106_, new_n12107_,
    new_n12108_, new_n12109_, new_n12110_, new_n12111_, new_n12112_,
    new_n12113_, new_n12114_, new_n12115_, new_n12116_, new_n12117_,
    new_n12118_, new_n12119_, new_n12120_, new_n12121_, new_n12122_,
    new_n12123_, new_n12124_, new_n12125_, new_n12126_, new_n12127_,
    new_n12128_, new_n12129_, new_n12130_, new_n12131_, new_n12132_,
    new_n12133_, new_n12134_, new_n12135_, new_n12136_, new_n12137_,
    new_n12138_, new_n12139_, new_n12140_, new_n12141_, new_n12142_,
    new_n12143_, new_n12144_, new_n12145_, new_n12146_, new_n12147_,
    new_n12148_, new_n12149_, new_n12150_, new_n12151_, new_n12152_,
    new_n12153_, new_n12154_, new_n12155_, new_n12156_, new_n12157_,
    new_n12158_, new_n12159_, new_n12160_, new_n12161_, new_n12162_,
    new_n12163_, new_n12164_, new_n12165_, new_n12166_, new_n12167_,
    new_n12168_, new_n12169_, new_n12170_, new_n12171_, new_n12172_,
    new_n12173_, new_n12174_, new_n12175_, new_n12176_, new_n12177_,
    new_n12178_, new_n12179_, new_n12180_, new_n12181_, new_n12182_,
    new_n12183_, new_n12184_, new_n12185_, new_n12186_, new_n12187_,
    new_n12188_, new_n12189_, new_n12190_, new_n12191_, new_n12192_,
    new_n12193_, new_n12194_, new_n12195_, new_n12196_, new_n12197_,
    new_n12198_, new_n12199_, new_n12200_, new_n12201_, new_n12202_,
    new_n12203_, new_n12204_, new_n12205_, new_n12206_, new_n12207_,
    new_n12208_, new_n12209_, new_n12210_, new_n12211_, new_n12212_,
    new_n12213_, new_n12214_, new_n12215_, new_n12216_, new_n12217_,
    new_n12218_, new_n12219_, new_n12220_, new_n12221_, new_n12222_,
    new_n12223_, new_n12224_, new_n12225_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12254_, new_n12255_, new_n12256_, new_n12257_, new_n12258_,
    new_n12259_, new_n12260_, new_n12261_, new_n12262_, new_n12263_,
    new_n12264_, new_n12265_, new_n12266_, new_n12267_, new_n12268_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12280_, new_n12281_, new_n12282_, new_n12283_,
    new_n12284_, new_n12285_, new_n12286_, new_n12287_, new_n12288_,
    new_n12289_, new_n12290_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12296_, new_n12297_, new_n12298_,
    new_n12299_, new_n12300_, new_n12301_, new_n12302_, new_n12303_,
    new_n12304_, new_n12305_, new_n12306_, new_n12307_, new_n12308_,
    new_n12309_, new_n12310_, new_n12311_, new_n12312_, new_n12313_,
    new_n12314_, new_n12315_, new_n12316_, new_n12317_, new_n12318_,
    new_n12319_, new_n12320_, new_n12321_, new_n12322_, new_n12323_,
    new_n12324_, new_n12325_, new_n12326_, new_n12327_, new_n12328_,
    new_n12329_, new_n12330_, new_n12331_, new_n12332_, new_n12333_,
    new_n12334_, new_n12335_, new_n12336_, new_n12337_, new_n12338_,
    new_n12339_, new_n12340_, new_n12341_, new_n12342_, new_n12343_,
    new_n12344_, new_n12345_, new_n12346_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12470_,
    new_n12471_, new_n12472_, new_n12473_, new_n12474_, new_n12475_,
    new_n12476_, new_n12477_, new_n12478_, new_n12479_, new_n12480_,
    new_n12481_, new_n12482_, new_n12483_, new_n12484_, new_n12485_,
    new_n12486_, new_n12487_, new_n12488_, new_n12489_, new_n12490_,
    new_n12491_, new_n12492_, new_n12493_, new_n12494_, new_n12495_,
    new_n12496_, new_n12497_, new_n12498_, new_n12499_, new_n12500_,
    new_n12501_, new_n12502_, new_n12503_, new_n12504_, new_n12505_,
    new_n12506_, new_n12507_, new_n12508_, new_n12509_, new_n12510_,
    new_n12511_, new_n12512_, new_n12513_, new_n12514_, new_n12515_,
    new_n12516_, new_n12517_, new_n12518_, new_n12519_, new_n12520_,
    new_n12521_, new_n12522_, new_n12523_, new_n12524_, new_n12525_,
    new_n12526_, new_n12527_, new_n12528_, new_n12529_, new_n12530_,
    new_n12531_, new_n12532_, new_n12533_, new_n12534_, new_n12535_,
    new_n12536_, new_n12537_, new_n12538_, new_n12539_, new_n12540_,
    new_n12541_, new_n12542_, new_n12543_, new_n12544_, new_n12545_,
    new_n12546_, new_n12547_, new_n12548_, new_n12549_, new_n12550_,
    new_n12551_, new_n12552_, new_n12553_, new_n12554_, new_n12555_,
    new_n12556_, new_n12557_, new_n12558_, new_n12559_, new_n12560_,
    new_n12561_, new_n12562_, new_n12563_, new_n12564_, new_n12565_,
    new_n12566_, new_n12567_, new_n12568_, new_n12569_, new_n12570_,
    new_n12571_, new_n12572_, new_n12573_, new_n12574_, new_n12575_,
    new_n12576_, new_n12577_, new_n12578_, new_n12579_, new_n12580_,
    new_n12582_, new_n12583_, new_n12584_, new_n12585_, new_n12586_,
    new_n12587_, new_n12588_, new_n12589_, new_n12590_, new_n12591_,
    new_n12592_, new_n12593_, new_n12594_, new_n12595_, new_n12596_,
    new_n12597_, new_n12598_, new_n12599_, new_n12600_, new_n12601_,
    new_n12602_, new_n12603_, new_n12604_, new_n12605_, new_n12606_,
    new_n12607_, new_n12608_, new_n12609_, new_n12610_, new_n12611_,
    new_n12612_, new_n12613_, new_n12614_, new_n12615_, new_n12616_,
    new_n12617_, new_n12618_, new_n12619_, new_n12620_, new_n12621_,
    new_n12622_, new_n12623_, new_n12624_, new_n12625_, new_n12626_,
    new_n12627_, new_n12628_, new_n12629_, new_n12630_, new_n12631_,
    new_n12632_, new_n12633_, new_n12634_, new_n12635_, new_n12636_,
    new_n12637_, new_n12638_, new_n12639_, new_n12640_, new_n12641_,
    new_n12642_, new_n12643_, new_n12644_, new_n12645_, new_n12646_,
    new_n12647_, new_n12648_, new_n12649_, new_n12650_, new_n12651_,
    new_n12652_, new_n12653_, new_n12654_, new_n12655_, new_n12656_,
    new_n12657_, new_n12658_, new_n12659_, new_n12660_, new_n12661_,
    new_n12662_, new_n12663_, new_n12664_, new_n12665_, new_n12666_,
    new_n12667_, new_n12668_, new_n12669_, new_n12670_, new_n12671_,
    new_n12672_, new_n12673_, new_n12674_, new_n12675_, new_n12676_,
    new_n12677_, new_n12678_, new_n12679_, new_n12680_, new_n12681_,
    new_n12682_, new_n12683_, new_n12684_, new_n12685_, new_n12686_,
    new_n12687_, new_n12689_, new_n12690_, new_n12691_, new_n12692_,
    new_n12693_, new_n12694_, new_n12695_, new_n12696_, new_n12697_,
    new_n12698_, new_n12699_, new_n12700_, new_n12701_, new_n12702_,
    new_n12703_, new_n12704_, new_n12705_, new_n12706_, new_n12707_,
    new_n12708_, new_n12709_, new_n12710_, new_n12711_, new_n12712_,
    new_n12713_, new_n12714_, new_n12715_, new_n12716_, new_n12717_,
    new_n12718_, new_n12719_, new_n12720_, new_n12721_, new_n12722_,
    new_n12723_, new_n12724_, new_n12725_, new_n12726_, new_n12727_,
    new_n12728_, new_n12729_, new_n12730_, new_n12731_, new_n12732_,
    new_n12733_, new_n12734_, new_n12735_, new_n12736_, new_n12737_,
    new_n12738_, new_n12739_, new_n12740_, new_n12741_, new_n12742_,
    new_n12743_, new_n12744_, new_n12745_, new_n12746_, new_n12747_,
    new_n12748_, new_n12749_, new_n12750_, new_n12751_, new_n12752_,
    new_n12753_, new_n12754_, new_n12755_, new_n12756_, new_n12757_,
    new_n12758_, new_n12759_, new_n12760_, new_n12761_, new_n12762_,
    new_n12763_, new_n12764_, new_n12765_, new_n12766_, new_n12767_,
    new_n12768_, new_n12769_, new_n12770_, new_n12771_, new_n12772_,
    new_n12773_, new_n12774_, new_n12775_, new_n12776_, new_n12777_,
    new_n12778_, new_n12779_, new_n12780_, new_n12781_, new_n12782_,
    new_n12783_, new_n12784_, new_n12785_, new_n12786_, new_n12787_,
    new_n12788_, new_n12789_, new_n12790_, new_n12791_, new_n12792_,
    new_n12793_, new_n12794_, new_n12795_, new_n12796_, new_n12797_,
    new_n12798_, new_n12799_, new_n12800_, new_n12802_, new_n12803_,
    new_n12804_, new_n12805_, new_n12806_, new_n12807_, new_n12808_,
    new_n12809_, new_n12810_, new_n12811_, new_n12812_, new_n12813_,
    new_n12814_, new_n12815_, new_n12816_, new_n12817_, new_n12818_,
    new_n12819_, new_n12820_, new_n12821_, new_n12822_, new_n12823_,
    new_n12824_, new_n12825_, new_n12826_, new_n12827_, new_n12828_,
    new_n12829_, new_n12830_, new_n12831_, new_n12832_, new_n12833_,
    new_n12834_, new_n12835_, new_n12836_, new_n12837_, new_n12838_,
    new_n12839_, new_n12840_, new_n12841_, new_n12842_, new_n12843_,
    new_n12844_, new_n12845_, new_n12846_, new_n12847_, new_n12848_,
    new_n12849_, new_n12850_, new_n12851_, new_n12852_, new_n12853_,
    new_n12854_, new_n12855_, new_n12856_, new_n12857_, new_n12858_,
    new_n12859_, new_n12860_, new_n12861_, new_n12862_, new_n12863_,
    new_n12864_, new_n12865_, new_n12866_, new_n12867_, new_n12868_,
    new_n12869_, new_n12870_, new_n12871_, new_n12872_, new_n12873_,
    new_n12874_, new_n12875_, new_n12876_, new_n12877_, new_n12878_,
    new_n12879_, new_n12880_, new_n12881_, new_n12882_, new_n12883_,
    new_n12884_, new_n12885_, new_n12886_, new_n12887_, new_n12888_,
    new_n12889_, new_n12890_, new_n12891_, new_n12892_, new_n12893_,
    new_n12894_, new_n12895_, new_n12896_, new_n12897_, new_n12898_,
    new_n12899_, new_n12900_, new_n12901_, new_n12902_, new_n12903_,
    new_n12904_, new_n12905_, new_n12906_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13006_, new_n13007_, new_n13008_, new_n13009_, new_n13010_,
    new_n13011_, new_n13012_, new_n13013_, new_n13014_, new_n13015_,
    new_n13016_, new_n13017_, new_n13018_, new_n13019_, new_n13020_,
    new_n13021_, new_n13022_, new_n13023_, new_n13024_, new_n13025_,
    new_n13026_, new_n13027_, new_n13028_, new_n13029_, new_n13030_,
    new_n13031_, new_n13032_, new_n13033_, new_n13034_, new_n13035_,
    new_n13036_, new_n13037_, new_n13038_, new_n13039_, new_n13040_,
    new_n13041_, new_n13042_, new_n13043_, new_n13044_, new_n13045_,
    new_n13046_, new_n13047_, new_n13048_, new_n13049_, new_n13050_,
    new_n13051_, new_n13052_, new_n13053_, new_n13054_, new_n13055_,
    new_n13056_, new_n13057_, new_n13058_, new_n13059_, new_n13060_,
    new_n13061_, new_n13062_, new_n13063_, new_n13064_, new_n13065_,
    new_n13066_, new_n13067_, new_n13068_, new_n13069_, new_n13070_,
    new_n13071_, new_n13072_, new_n13073_, new_n13074_, new_n13075_,
    new_n13076_, new_n13077_, new_n13078_, new_n13079_, new_n13080_,
    new_n13081_, new_n13082_, new_n13083_, new_n13084_, new_n13085_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13111_,
    new_n13112_, new_n13113_, new_n13114_, new_n13115_, new_n13116_,
    new_n13117_, new_n13118_, new_n13119_, new_n13120_, new_n13121_,
    new_n13122_, new_n13123_, new_n13124_, new_n13125_, new_n13126_,
    new_n13127_, new_n13128_, new_n13129_, new_n13130_, new_n13131_,
    new_n13132_, new_n13133_, new_n13134_, new_n13135_, new_n13136_,
    new_n13137_, new_n13138_, new_n13139_, new_n13140_, new_n13141_,
    new_n13142_, new_n13143_, new_n13144_, new_n13145_, new_n13146_,
    new_n13147_, new_n13148_, new_n13149_, new_n13150_, new_n13151_,
    new_n13152_, new_n13153_, new_n13154_, new_n13155_, new_n13156_,
    new_n13157_, new_n13158_, new_n13159_, new_n13160_, new_n13161_,
    new_n13162_, new_n13163_, new_n13164_, new_n13165_, new_n13166_,
    new_n13167_, new_n13168_, new_n13169_, new_n13170_, new_n13171_,
    new_n13172_, new_n13173_, new_n13174_, new_n13175_, new_n13176_,
    new_n13177_, new_n13178_, new_n13179_, new_n13180_, new_n13181_,
    new_n13182_, new_n13183_, new_n13184_, new_n13185_, new_n13186_,
    new_n13187_, new_n13188_, new_n13189_, new_n13190_, new_n13191_,
    new_n13192_, new_n13193_, new_n13194_, new_n13195_, new_n13196_,
    new_n13197_, new_n13198_, new_n13199_, new_n13200_, new_n13202_,
    new_n13203_, new_n13204_, new_n13205_, new_n13206_, new_n13207_,
    new_n13208_, new_n13209_, new_n13210_, new_n13211_, new_n13212_,
    new_n13213_, new_n13214_, new_n13215_, new_n13216_, new_n13217_,
    new_n13218_, new_n13219_, new_n13220_, new_n13221_, new_n13222_,
    new_n13223_, new_n13224_, new_n13225_, new_n13226_, new_n13227_,
    new_n13228_, new_n13229_, new_n13230_, new_n13231_, new_n13232_,
    new_n13233_, new_n13234_, new_n13235_, new_n13236_, new_n13237_,
    new_n13238_, new_n13239_, new_n13240_, new_n13241_, new_n13242_,
    new_n13243_, new_n13244_, new_n13245_, new_n13246_, new_n13247_,
    new_n13248_, new_n13249_, new_n13250_, new_n13251_, new_n13252_,
    new_n13253_, new_n13254_, new_n13255_, new_n13256_, new_n13257_,
    new_n13258_, new_n13259_, new_n13260_, new_n13261_, new_n13262_,
    new_n13263_, new_n13264_, new_n13265_, new_n13266_, new_n13267_,
    new_n13268_, new_n13269_, new_n13270_, new_n13271_, new_n13272_,
    new_n13273_, new_n13274_, new_n13275_, new_n13276_, new_n13277_,
    new_n13278_, new_n13279_, new_n13280_, new_n13281_, new_n13282_,
    new_n13283_, new_n13284_, new_n13285_, new_n13286_, new_n13287_,
    new_n13288_, new_n13290_, new_n13291_, new_n13292_, new_n13293_,
    new_n13294_, new_n13295_, new_n13296_, new_n13297_, new_n13298_,
    new_n13299_, new_n13300_, new_n13301_, new_n13302_, new_n13303_,
    new_n13304_, new_n13305_, new_n13306_, new_n13307_, new_n13308_,
    new_n13309_, new_n13310_, new_n13311_, new_n13312_, new_n13313_,
    new_n13314_, new_n13315_, new_n13316_, new_n13317_, new_n13318_,
    new_n13319_, new_n13320_, new_n13321_, new_n13322_, new_n13323_,
    new_n13324_, new_n13325_, new_n13326_, new_n13327_, new_n13328_,
    new_n13329_, new_n13330_, new_n13331_, new_n13332_, new_n13333_,
    new_n13334_, new_n13335_, new_n13336_, new_n13337_, new_n13338_,
    new_n13339_, new_n13340_, new_n13341_, new_n13342_, new_n13343_,
    new_n13344_, new_n13345_, new_n13346_, new_n13347_, new_n13348_,
    new_n13349_, new_n13350_, new_n13351_, new_n13352_, new_n13353_,
    new_n13354_, new_n13355_, new_n13356_, new_n13357_, new_n13358_,
    new_n13359_, new_n13360_, new_n13361_, new_n13362_, new_n13363_,
    new_n13364_, new_n13365_, new_n13366_, new_n13367_, new_n13368_,
    new_n13369_, new_n13370_, new_n13371_, new_n13372_, new_n13373_,
    new_n13374_, new_n13375_, new_n13376_, new_n13377_, new_n13378_,
    new_n13379_, new_n13380_, new_n13382_, new_n13383_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13396_, new_n13397_, new_n13398_, new_n13399_,
    new_n13400_, new_n13401_, new_n13402_, new_n13403_, new_n13404_,
    new_n13405_, new_n13406_, new_n13407_, new_n13408_, new_n13409_,
    new_n13410_, new_n13411_, new_n13412_, new_n13413_, new_n13414_,
    new_n13415_, new_n13416_, new_n13417_, new_n13418_, new_n13419_,
    new_n13420_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13425_, new_n13426_, new_n13427_, new_n13428_, new_n13429_,
    new_n13430_, new_n13431_, new_n13432_, new_n13433_, new_n13434_,
    new_n13435_, new_n13436_, new_n13437_, new_n13438_, new_n13439_,
    new_n13440_, new_n13441_, new_n13442_, new_n13443_, new_n13444_,
    new_n13445_, new_n13446_, new_n13447_, new_n13448_, new_n13449_,
    new_n13450_, new_n13451_, new_n13452_, new_n13453_, new_n13454_,
    new_n13455_, new_n13456_, new_n13457_, new_n13458_, new_n13459_,
    new_n13460_, new_n13461_, new_n13462_, new_n13463_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13537_, new_n13538_, new_n13539_, new_n13540_,
    new_n13541_, new_n13542_, new_n13543_, new_n13544_, new_n13545_,
    new_n13546_, new_n13547_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13633_, new_n13634_, new_n13635_, new_n13636_, new_n13637_,
    new_n13638_, new_n13639_, new_n13640_, new_n13641_, new_n13642_,
    new_n13643_, new_n13644_, new_n13645_, new_n13646_, new_n13647_,
    new_n13648_, new_n13649_, new_n13650_, new_n13651_, new_n13652_,
    new_n13653_, new_n13654_, new_n13655_, new_n13656_, new_n13657_,
    new_n13658_, new_n13659_, new_n13660_, new_n13661_, new_n13662_,
    new_n13663_, new_n13664_, new_n13665_, new_n13666_, new_n13667_,
    new_n13668_, new_n13669_, new_n13670_, new_n13671_, new_n13672_,
    new_n13673_, new_n13674_, new_n13675_, new_n13676_, new_n13677_,
    new_n13678_, new_n13679_, new_n13680_, new_n13681_, new_n13682_,
    new_n13683_, new_n13684_, new_n13685_, new_n13686_, new_n13687_,
    new_n13688_, new_n13689_, new_n13690_, new_n13691_, new_n13692_,
    new_n13693_, new_n13694_, new_n13695_, new_n13696_, new_n13697_,
    new_n13698_, new_n13699_, new_n13700_, new_n13701_, new_n13702_,
    new_n13703_, new_n13704_, new_n13705_, new_n13707_, new_n13708_,
    new_n13709_, new_n13710_, new_n13711_, new_n13712_, new_n13713_,
    new_n13714_, new_n13715_, new_n13716_, new_n13717_, new_n13718_,
    new_n13719_, new_n13720_, new_n13721_, new_n13722_, new_n13723_,
    new_n13724_, new_n13725_, new_n13726_, new_n13727_, new_n13728_,
    new_n13729_, new_n13730_, new_n13731_, new_n13732_, new_n13733_,
    new_n13734_, new_n13735_, new_n13736_, new_n13737_, new_n13738_,
    new_n13739_, new_n13740_, new_n13741_, new_n13742_, new_n13743_,
    new_n13744_, new_n13745_, new_n13746_, new_n13747_, new_n13748_,
    new_n13749_, new_n13750_, new_n13751_, new_n13752_, new_n13753_,
    new_n13754_, new_n13755_, new_n13756_, new_n13757_, new_n13758_,
    new_n13759_, new_n13760_, new_n13761_, new_n13762_, new_n13763_,
    new_n13764_, new_n13765_, new_n13766_, new_n13767_, new_n13768_,
    new_n13769_, new_n13770_, new_n13771_, new_n13772_, new_n13773_,
    new_n13774_, new_n13775_, new_n13776_, new_n13777_, new_n13778_,
    new_n13780_, new_n13781_, new_n13782_, new_n13783_, new_n13784_,
    new_n13785_, new_n13786_, new_n13787_, new_n13788_, new_n13789_,
    new_n13790_, new_n13791_, new_n13792_, new_n13793_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13799_,
    new_n13800_, new_n13801_, new_n13802_, new_n13803_, new_n13804_,
    new_n13805_, new_n13806_, new_n13807_, new_n13808_, new_n13809_,
    new_n13810_, new_n13811_, new_n13812_, new_n13813_, new_n13814_,
    new_n13815_, new_n13816_, new_n13817_, new_n13818_, new_n13819_,
    new_n13820_, new_n13821_, new_n13822_, new_n13823_, new_n13824_,
    new_n13825_, new_n13826_, new_n13827_, new_n13828_, new_n13829_,
    new_n13830_, new_n13831_, new_n13832_, new_n13833_, new_n13834_,
    new_n13835_, new_n13836_, new_n13837_, new_n13838_, new_n13839_,
    new_n13840_, new_n13841_, new_n13842_, new_n13843_, new_n13844_,
    new_n13845_, new_n13846_, new_n13847_, new_n13848_, new_n13849_,
    new_n13850_, new_n13851_, new_n13852_, new_n13854_, new_n13855_,
    new_n13856_, new_n13857_, new_n13858_, new_n13859_, new_n13860_,
    new_n13861_, new_n13862_, new_n13863_, new_n13864_, new_n13865_,
    new_n13866_, new_n13867_, new_n13868_, new_n13869_, new_n13870_,
    new_n13871_, new_n13872_, new_n13873_, new_n13874_, new_n13875_,
    new_n13876_, new_n13877_, new_n13878_, new_n13879_, new_n13880_,
    new_n13881_, new_n13882_, new_n13883_, new_n13884_, new_n13885_,
    new_n13886_, new_n13887_, new_n13888_, new_n13889_, new_n13890_,
    new_n13891_, new_n13892_, new_n13893_, new_n13894_, new_n13895_,
    new_n13896_, new_n13897_, new_n13898_, new_n13899_, new_n13900_,
    new_n13901_, new_n13902_, new_n13903_, new_n13904_, new_n13905_,
    new_n13906_, new_n13907_, new_n13908_, new_n13909_, new_n13910_,
    new_n13911_, new_n13912_, new_n13913_, new_n13914_, new_n13915_,
    new_n13916_, new_n13918_, new_n13919_, new_n13920_, new_n13921_,
    new_n13922_, new_n13923_, new_n13924_, new_n13925_, new_n13926_,
    new_n13927_, new_n13928_, new_n13929_, new_n13930_, new_n13931_,
    new_n13932_, new_n13933_, new_n13934_, new_n13935_, new_n13936_,
    new_n13937_, new_n13938_, new_n13939_, new_n13940_, new_n13941_,
    new_n13942_, new_n13943_, new_n13944_, new_n13945_, new_n13946_,
    new_n13947_, new_n13948_, new_n13949_, new_n13950_, new_n13951_,
    new_n13952_, new_n13953_, new_n13954_, new_n13955_, new_n13956_,
    new_n13957_, new_n13958_, new_n13959_, new_n13960_, new_n13961_,
    new_n13962_, new_n13963_, new_n13964_, new_n13965_, new_n13966_,
    new_n13967_, new_n13968_, new_n13969_, new_n13970_, new_n13971_,
    new_n13972_, new_n13973_, new_n13974_, new_n13975_, new_n13976_,
    new_n13977_, new_n13978_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13998_, new_n13999_, new_n14000_, new_n14001_, new_n14002_,
    new_n14003_, new_n14004_, new_n14005_, new_n14006_, new_n14007_,
    new_n14008_, new_n14009_, new_n14010_, new_n14011_, new_n14012_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14019_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14031_, new_n14032_,
    new_n14033_, new_n14034_, new_n14035_, new_n14036_, new_n14037_,
    new_n14038_, new_n14039_, new_n14040_, new_n14041_, new_n14042_,
    new_n14043_, new_n14045_, new_n14046_, new_n14047_, new_n14048_,
    new_n14049_, new_n14050_, new_n14051_, new_n14052_, new_n14053_,
    new_n14054_, new_n14055_, new_n14056_, new_n14057_, new_n14058_,
    new_n14059_, new_n14060_, new_n14061_, new_n14062_, new_n14063_,
    new_n14064_, new_n14065_, new_n14066_, new_n14067_, new_n14068_,
    new_n14069_, new_n14070_, new_n14071_, new_n14072_, new_n14073_,
    new_n14074_, new_n14075_, new_n14076_, new_n14077_, new_n14078_,
    new_n14079_, new_n14080_, new_n14081_, new_n14082_, new_n14083_,
    new_n14084_, new_n14085_, new_n14086_, new_n14087_, new_n14088_,
    new_n14089_, new_n14090_, new_n14091_, new_n14092_, new_n14093_,
    new_n14094_, new_n14095_, new_n14096_, new_n14097_, new_n14098_,
    new_n14100_, new_n14101_, new_n14102_, new_n14103_, new_n14104_,
    new_n14105_, new_n14106_, new_n14107_, new_n14108_, new_n14109_,
    new_n14110_, new_n14111_, new_n14112_, new_n14113_, new_n14114_,
    new_n14115_, new_n14116_, new_n14117_, new_n14118_, new_n14119_,
    new_n14120_, new_n14121_, new_n14122_, new_n14123_, new_n14124_,
    new_n14125_, new_n14126_, new_n14127_, new_n14128_, new_n14129_,
    new_n14130_, new_n14131_, new_n14132_, new_n14133_, new_n14134_,
    new_n14135_, new_n14136_, new_n14137_, new_n14138_, new_n14139_,
    new_n14140_, new_n14141_, new_n14142_, new_n14143_, new_n14144_,
    new_n14145_, new_n14146_, new_n14147_, new_n14148_, new_n14149_,
    new_n14150_, new_n14151_, new_n14152_, new_n14153_, new_n14154_,
    new_n14156_, new_n14157_, new_n14158_, new_n14159_, new_n14160_,
    new_n14161_, new_n14162_, new_n14163_, new_n14164_, new_n14165_,
    new_n14166_, new_n14167_, new_n14168_, new_n14169_, new_n14170_,
    new_n14171_, new_n14172_, new_n14173_, new_n14174_, new_n14175_,
    new_n14176_, new_n14177_, new_n14178_, new_n14179_, new_n14180_,
    new_n14181_, new_n14182_, new_n14183_, new_n14184_, new_n14185_,
    new_n14186_, new_n14187_, new_n14188_, new_n14189_, new_n14190_,
    new_n14191_, new_n14192_, new_n14193_, new_n14194_, new_n14195_,
    new_n14196_, new_n14197_, new_n14198_, new_n14199_, new_n14200_,
    new_n14201_, new_n14202_, new_n14203_, new_n14204_, new_n14205_,
    new_n14207_, new_n14208_, new_n14209_, new_n14210_, new_n14211_,
    new_n14212_, new_n14213_, new_n14214_, new_n14215_, new_n14216_,
    new_n14217_, new_n14218_, new_n14219_, new_n14220_, new_n14221_,
    new_n14222_, new_n14223_, new_n14224_, new_n14225_, new_n14226_,
    new_n14227_, new_n14228_, new_n14229_, new_n14230_, new_n14231_,
    new_n14232_, new_n14233_, new_n14234_, new_n14235_, new_n14236_,
    new_n14237_, new_n14238_, new_n14239_, new_n14240_, new_n14241_,
    new_n14242_, new_n14243_, new_n14244_, new_n14245_, new_n14246_,
    new_n14247_, new_n14248_, new_n14249_, new_n14250_, new_n14251_,
    new_n14252_, new_n14253_, new_n14254_, new_n14255_, new_n14256_,
    new_n14258_, new_n14259_, new_n14260_, new_n14261_, new_n14262_,
    new_n14263_, new_n14264_, new_n14265_, new_n14266_, new_n14267_,
    new_n14268_, new_n14269_, new_n14270_, new_n14271_, new_n14272_,
    new_n14273_, new_n14274_, new_n14275_, new_n14276_, new_n14277_,
    new_n14278_, new_n14279_, new_n14280_, new_n14281_, new_n14282_,
    new_n14283_, new_n14284_, new_n14285_, new_n14286_, new_n14287_,
    new_n14288_, new_n14289_, new_n14290_, new_n14291_, new_n14292_,
    new_n14293_, new_n14294_, new_n14295_, new_n14296_, new_n14297_,
    new_n14298_, new_n14299_, new_n14300_, new_n14301_, new_n14303_,
    new_n14304_, new_n14305_, new_n14306_, new_n14307_, new_n14308_,
    new_n14309_, new_n14310_, new_n14311_, new_n14312_, new_n14313_,
    new_n14314_, new_n14315_, new_n14316_, new_n14317_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14324_, new_n14325_, new_n14326_, new_n14327_, new_n14328_,
    new_n14329_, new_n14330_, new_n14331_, new_n14332_, new_n14333_,
    new_n14334_, new_n14335_, new_n14336_, new_n14337_, new_n14338_,
    new_n14339_, new_n14340_, new_n14341_, new_n14342_, new_n14343_,
    new_n14344_, new_n14345_, new_n14346_, new_n14348_, new_n14349_,
    new_n14350_, new_n14351_, new_n14352_, new_n14353_, new_n14354_,
    new_n14355_, new_n14356_, new_n14357_, new_n14358_, new_n14359_,
    new_n14360_, new_n14361_, new_n14362_, new_n14363_, new_n14364_,
    new_n14365_, new_n14366_, new_n14367_, new_n14368_, new_n14369_,
    new_n14370_, new_n14371_, new_n14372_, new_n14373_, new_n14374_,
    new_n14375_, new_n14376_, new_n14377_, new_n14378_, new_n14379_,
    new_n14380_, new_n14381_, new_n14382_, new_n14383_, new_n14385_,
    new_n14386_, new_n14387_, new_n14388_, new_n14389_, new_n14390_,
    new_n14391_, new_n14392_, new_n14393_, new_n14394_, new_n14395_,
    new_n14396_, new_n14397_, new_n14398_, new_n14399_, new_n14400_,
    new_n14401_, new_n14402_, new_n14403_, new_n14404_, new_n14405_,
    new_n14406_, new_n14407_, new_n14408_, new_n14409_, new_n14410_,
    new_n14411_, new_n14412_, new_n14413_, new_n14414_, new_n14415_,
    new_n14416_, new_n14417_, new_n14418_, new_n14419_, new_n14420_,
    new_n14421_, new_n14423_, new_n14424_, new_n14425_, new_n14426_,
    new_n14427_, new_n14428_, new_n14429_, new_n14430_, new_n14431_,
    new_n14432_, new_n14433_, new_n14434_, new_n14435_, new_n14436_,
    new_n14437_, new_n14438_, new_n14439_, new_n14440_, new_n14441_,
    new_n14442_, new_n14443_, new_n14444_, new_n14445_, new_n14446_,
    new_n14447_, new_n14448_, new_n14449_, new_n14450_, new_n14451_,
    new_n14452_, new_n14453_, new_n14454_, new_n14456_, new_n14457_,
    new_n14458_, new_n14459_, new_n14460_, new_n14461_, new_n14462_,
    new_n14463_, new_n14464_, new_n14465_, new_n14466_, new_n14467_,
    new_n14468_, new_n14469_, new_n14470_, new_n14471_, new_n14472_,
    new_n14473_, new_n14474_, new_n14475_, new_n14476_, new_n14477_,
    new_n14478_, new_n14479_, new_n14480_, new_n14481_, new_n14482_,
    new_n14483_, new_n14484_, new_n14485_, new_n14487_, new_n14488_,
    new_n14489_, new_n14490_, new_n14491_, new_n14492_, new_n14493_,
    new_n14494_, new_n14495_, new_n14496_, new_n14497_, new_n14498_,
    new_n14499_, new_n14500_, new_n14501_, new_n14502_, new_n14503_,
    new_n14504_, new_n14505_, new_n14506_, new_n14507_, new_n14508_,
    new_n14509_, new_n14510_, new_n14511_, new_n14512_, new_n14513_,
    new_n14515_, new_n14516_, new_n14517_, new_n14518_, new_n14519_,
    new_n14520_, new_n14521_, new_n14522_, new_n14523_, new_n14524_,
    new_n14525_, new_n14526_, new_n14527_, new_n14528_, new_n14529_,
    new_n14530_, new_n14531_, new_n14532_, new_n14533_, new_n14534_,
    new_n14535_, new_n14536_, new_n14537_, new_n14538_, new_n14539_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14561_,
    new_n14562_, new_n14563_, new_n14564_, new_n14565_, new_n14566_,
    new_n14567_, new_n14568_, new_n14569_, new_n14570_, new_n14571_,
    new_n14572_, new_n14573_, new_n14574_, new_n14575_, new_n14576_,
    new_n14577_, new_n14578_, new_n14579_, new_n14580_, new_n14581_,
    new_n14583_, new_n14584_, new_n14585_, new_n14586_, new_n14587_,
    new_n14588_, new_n14589_, new_n14590_, new_n14591_, new_n14592_,
    new_n14593_, new_n14594_, new_n14595_, new_n14596_, new_n14598_,
    new_n14599_, new_n14600_, new_n14601_, new_n14602_, new_n14603_,
    new_n14604_, new_n14605_, new_n14607_, new_n14608_, new_n14609_,
    new_n14610_, new_n14611_, new_n14612_;
  INVX1    g00000(.A(\a[2] ), .Y(new_n257_));
  AND2X1   g00001(.A(\b[0] ), .B(\a[0] ), .Y(new_n258_));
  OR2X1    g00002(.A(new_n258_), .B(new_n257_), .Y(new_n259_));
  OR2X1    g00003(.A(new_n258_), .B(\a[2] ), .Y(new_n260_));
  AND2X1   g00004(.A(new_n260_), .B(new_n259_), .Y(\f[0] ));
  XOR2X1   g00005(.A(\a[2] ), .B(\a[1] ), .Y(new_n262_));
  XOR2X1   g00006(.A(\b[1] ), .B(\b[0] ), .Y(new_n263_));
  NAND3X1  g00007(.A(new_n263_), .B(new_n262_), .C(\a[0] ), .Y(new_n264_));
  INVX1    g00008(.A(\a[0] ), .Y(new_n265_));
  AND2X1   g00009(.A(\a[1] ), .B(new_n265_), .Y(new_n266_));
  NOR2X1   g00010(.A(new_n262_), .B(new_n265_), .Y(new_n267_));
  AOI22X1  g00011(.A0(new_n267_), .A1(\b[1] ), .B0(new_n266_), .B1(\b[0] ), .Y(new_n268_));
  NAND2X1  g00012(.A(new_n268_), .B(new_n264_), .Y(new_n269_));
  XOR2X1   g00013(.A(new_n269_), .B(new_n257_), .Y(new_n270_));
  XOR2X1   g00014(.A(new_n270_), .B(new_n259_), .Y(\f[1] ));
  OR2X1    g00015(.A(new_n270_), .B(new_n259_), .Y(new_n272_));
  NAND2X1  g00016(.A(new_n262_), .B(\a[0] ), .Y(new_n273_));
  INVX1    g00017(.A(\b[0] ), .Y(new_n274_));
  INVX1    g00018(.A(\b[1] ), .Y(new_n275_));
  NOR3X1   g00019(.A(\b[2] ), .B(new_n275_), .C(new_n274_), .Y(new_n276_));
  INVX1    g00020(.A(\b[2] ), .Y(new_n277_));
  OR2X1    g00021(.A(new_n277_), .B(\b[1] ), .Y(new_n278_));
  OAI21X1  g00022(.A0(new_n277_), .A1(\b[0] ), .B0(\b[1] ), .Y(new_n279_));
  AND2X1   g00023(.A(new_n279_), .B(new_n278_), .Y(new_n280_));
  OR2X1    g00024(.A(new_n280_), .B(new_n276_), .Y(new_n281_));
  NOR3X1   g00025(.A(new_n257_), .B(\a[1] ), .C(\a[0] ), .Y(new_n282_));
  INVX1    g00026(.A(\a[1] ), .Y(new_n283_));
  OR2X1    g00027(.A(new_n283_), .B(\a[0] ), .Y(new_n284_));
  OR2X1    g00028(.A(new_n262_), .B(new_n265_), .Y(new_n285_));
  OAI22X1  g00029(.A0(new_n285_), .A1(new_n277_), .B0(new_n284_), .B1(new_n275_), .Y(new_n286_));
  AOI21X1  g00030(.A0(new_n282_), .A1(\b[0] ), .B0(new_n286_), .Y(new_n287_));
  OAI21X1  g00031(.A0(new_n281_), .A1(new_n273_), .B0(new_n287_), .Y(new_n288_));
  XOR2X1   g00032(.A(new_n288_), .B(new_n257_), .Y(new_n289_));
  XOR2X1   g00033(.A(new_n289_), .B(new_n272_), .Y(\f[2] ));
  NOR4X1   g00034(.A(new_n288_), .B(new_n269_), .C(new_n258_), .D(new_n257_), .Y(new_n291_));
  OAI21X1  g00035(.A0(\b[2] ), .A1(\b[0] ), .B0(\b[1] ), .Y(new_n292_));
  XOR2X1   g00036(.A(\b[3] ), .B(\b[2] ), .Y(new_n293_));
  XOR2X1   g00037(.A(new_n293_), .B(new_n292_), .Y(new_n294_));
  NOR2X1   g00038(.A(new_n294_), .B(new_n273_), .Y(new_n295_));
  NOR4X1   g00039(.A(new_n275_), .B(new_n257_), .C(\a[1] ), .D(\a[0] ), .Y(new_n296_));
  INVX1    g00040(.A(\b[3] ), .Y(new_n297_));
  OAI22X1  g00041(.A0(new_n285_), .A1(new_n297_), .B0(new_n284_), .B1(new_n277_), .Y(new_n298_));
  NOR3X1   g00042(.A(new_n298_), .B(new_n296_), .C(new_n295_), .Y(new_n299_));
  XOR2X1   g00043(.A(new_n299_), .B(new_n257_), .Y(new_n300_));
  XOR2X1   g00044(.A(\a[3] ), .B(\a[2] ), .Y(new_n301_));
  AND2X1   g00045(.A(new_n301_), .B(\b[0] ), .Y(new_n302_));
  XOR2X1   g00046(.A(new_n302_), .B(new_n300_), .Y(new_n303_));
  XOR2X1   g00047(.A(new_n303_), .B(new_n291_), .Y(\f[3] ));
  INVX1    g00048(.A(\a[5] ), .Y(new_n305_));
  OR2X1    g00049(.A(new_n302_), .B(new_n305_), .Y(new_n306_));
  XOR2X1   g00050(.A(\a[5] ), .B(\a[4] ), .Y(new_n307_));
  AND2X1   g00051(.A(new_n307_), .B(new_n301_), .Y(new_n308_));
  AND2X1   g00052(.A(new_n308_), .B(new_n263_), .Y(new_n309_));
  INVX1    g00053(.A(\a[3] ), .Y(new_n310_));
  XOR2X1   g00054(.A(\a[4] ), .B(new_n310_), .Y(new_n311_));
  NOR3X1   g00055(.A(new_n311_), .B(new_n301_), .C(new_n274_), .Y(new_n312_));
  XOR2X1   g00056(.A(\a[3] ), .B(new_n257_), .Y(new_n313_));
  NOR3X1   g00057(.A(new_n307_), .B(new_n313_), .C(new_n275_), .Y(new_n314_));
  NOR3X1   g00058(.A(new_n314_), .B(new_n312_), .C(new_n309_), .Y(new_n315_));
  XOR2X1   g00059(.A(new_n315_), .B(\a[5] ), .Y(new_n316_));
  XOR2X1   g00060(.A(new_n316_), .B(new_n306_), .Y(new_n317_));
  AND2X1   g00061(.A(new_n262_), .B(\a[0] ), .Y(new_n318_));
  NOR2X1   g00062(.A(\b[3] ), .B(\b[2] ), .Y(new_n319_));
  NAND2X1  g00063(.A(\b[3] ), .B(\b[2] ), .Y(new_n320_));
  OAI21X1  g00064(.A0(new_n319_), .A1(new_n292_), .B0(new_n320_), .Y(new_n321_));
  XOR2X1   g00065(.A(\b[4] ), .B(\b[3] ), .Y(new_n322_));
  XOR2X1   g00066(.A(new_n322_), .B(new_n321_), .Y(new_n323_));
  NAND2X1  g00067(.A(new_n323_), .B(new_n318_), .Y(new_n324_));
  INVX1    g00068(.A(\b[4] ), .Y(new_n325_));
  OAI22X1  g00069(.A0(new_n285_), .A1(new_n325_), .B0(new_n284_), .B1(new_n297_), .Y(new_n326_));
  AOI21X1  g00070(.A0(new_n282_), .A1(\b[2] ), .B0(new_n326_), .Y(new_n327_));
  NAND2X1  g00071(.A(new_n327_), .B(new_n324_), .Y(new_n328_));
  XOR2X1   g00072(.A(new_n328_), .B(new_n257_), .Y(new_n329_));
  XOR2X1   g00073(.A(new_n329_), .B(new_n317_), .Y(new_n330_));
  AND2X1   g00074(.A(new_n302_), .B(new_n300_), .Y(new_n331_));
  AOI21X1  g00075(.A0(new_n303_), .A1(new_n291_), .B0(new_n331_), .Y(new_n332_));
  XOR2X1   g00076(.A(new_n332_), .B(new_n330_), .Y(\f[4] ));
  NOR2X1   g00077(.A(new_n316_), .B(new_n306_), .Y(new_n334_));
  XOR2X1   g00078(.A(new_n305_), .B(\a[4] ), .Y(new_n335_));
  XOR2X1   g00079(.A(\a[4] ), .B(\a[3] ), .Y(new_n336_));
  NOR4X1   g00080(.A(new_n336_), .B(new_n335_), .C(new_n301_), .D(new_n274_), .Y(new_n337_));
  NOR3X1   g00081(.A(new_n307_), .B(new_n313_), .C(new_n277_), .Y(new_n338_));
  NOR3X1   g00082(.A(new_n311_), .B(new_n301_), .C(new_n275_), .Y(new_n339_));
  OR4X1    g00083(.A(new_n339_), .B(new_n338_), .C(new_n337_), .D(new_n308_), .Y(new_n340_));
  AOI21X1  g00084(.A0(new_n279_), .A1(new_n278_), .B0(new_n276_), .Y(new_n341_));
  OR4X1    g00085(.A(new_n339_), .B(new_n338_), .C(new_n337_), .D(new_n341_), .Y(new_n342_));
  AND2X1   g00086(.A(new_n342_), .B(new_n340_), .Y(new_n343_));
  XOR2X1   g00087(.A(new_n343_), .B(new_n305_), .Y(new_n344_));
  XOR2X1   g00088(.A(new_n344_), .B(new_n334_), .Y(new_n345_));
  AND2X1   g00089(.A(\b[4] ), .B(\b[3] ), .Y(new_n346_));
  AOI21X1  g00090(.A0(new_n322_), .A1(new_n321_), .B0(new_n346_), .Y(new_n347_));
  XOR2X1   g00091(.A(\b[5] ), .B(new_n325_), .Y(new_n348_));
  XOR2X1   g00092(.A(new_n348_), .B(new_n347_), .Y(new_n349_));
  INVX1    g00093(.A(new_n282_), .Y(new_n350_));
  AOI22X1  g00094(.A0(new_n267_), .A1(\b[5] ), .B0(new_n266_), .B1(\b[4] ), .Y(new_n351_));
  OAI21X1  g00095(.A0(new_n350_), .A1(new_n297_), .B0(new_n351_), .Y(new_n352_));
  AOI21X1  g00096(.A0(new_n349_), .A1(new_n318_), .B0(new_n352_), .Y(new_n353_));
  XOR2X1   g00097(.A(new_n353_), .B(\a[2] ), .Y(new_n354_));
  XOR2X1   g00098(.A(new_n354_), .B(new_n345_), .Y(new_n355_));
  XOR2X1   g00099(.A(new_n328_), .B(\a[2] ), .Y(new_n356_));
  NAND2X1  g00100(.A(new_n356_), .B(new_n317_), .Y(new_n357_));
  OAI21X1  g00101(.A0(new_n332_), .A1(new_n330_), .B0(new_n357_), .Y(new_n358_));
  XOR2X1   g00102(.A(new_n358_), .B(new_n355_), .Y(\f[5] ));
  NOR2X1   g00103(.A(new_n354_), .B(new_n345_), .Y(new_n360_));
  AOI21X1  g00104(.A0(new_n358_), .A1(new_n355_), .B0(new_n360_), .Y(new_n361_));
  OR4X1    g00105(.A(new_n343_), .B(new_n316_), .C(new_n302_), .D(new_n305_), .Y(new_n362_));
  XOR2X1   g00106(.A(\a[6] ), .B(\a[5] ), .Y(new_n363_));
  AND2X1   g00107(.A(new_n363_), .B(\b[0] ), .Y(new_n364_));
  XOR2X1   g00108(.A(new_n364_), .B(new_n362_), .Y(new_n365_));
  INVX1    g00109(.A(new_n294_), .Y(new_n366_));
  NAND3X1  g00110(.A(new_n311_), .B(new_n307_), .C(new_n313_), .Y(new_n367_));
  AND2X1   g00111(.A(new_n336_), .B(new_n313_), .Y(new_n368_));
  AND2X1   g00112(.A(new_n335_), .B(new_n301_), .Y(new_n369_));
  AOI22X1  g00113(.A0(new_n369_), .A1(\b[3] ), .B0(new_n368_), .B1(\b[2] ), .Y(new_n370_));
  OAI21X1  g00114(.A0(new_n367_), .A1(new_n275_), .B0(new_n370_), .Y(new_n371_));
  AOI21X1  g00115(.A0(new_n308_), .A1(new_n366_), .B0(new_n371_), .Y(new_n372_));
  XOR2X1   g00116(.A(new_n372_), .B(\a[5] ), .Y(new_n373_));
  XOR2X1   g00117(.A(new_n373_), .B(new_n365_), .Y(new_n374_));
  NAND2X1  g00118(.A(\b[5] ), .B(\b[4] ), .Y(new_n375_));
  OAI21X1  g00119(.A0(new_n348_), .A1(new_n347_), .B0(new_n375_), .Y(new_n376_));
  XOR2X1   g00120(.A(\b[6] ), .B(\b[5] ), .Y(new_n377_));
  XOR2X1   g00121(.A(new_n377_), .B(new_n376_), .Y(new_n378_));
  AOI22X1  g00122(.A0(new_n267_), .A1(\b[6] ), .B0(new_n266_), .B1(\b[5] ), .Y(new_n379_));
  OAI21X1  g00123(.A0(new_n350_), .A1(new_n325_), .B0(new_n379_), .Y(new_n380_));
  AOI21X1  g00124(.A0(new_n378_), .A1(new_n318_), .B0(new_n380_), .Y(new_n381_));
  XOR2X1   g00125(.A(new_n381_), .B(\a[2] ), .Y(new_n382_));
  XOR2X1   g00126(.A(new_n382_), .B(new_n374_), .Y(new_n383_));
  XOR2X1   g00127(.A(new_n383_), .B(new_n361_), .Y(\f[6] ));
  NOR4X1   g00128(.A(new_n343_), .B(new_n316_), .C(new_n302_), .D(new_n305_), .Y(new_n385_));
  XOR2X1   g00129(.A(new_n364_), .B(new_n385_), .Y(new_n386_));
  XOR2X1   g00130(.A(new_n373_), .B(new_n386_), .Y(new_n387_));
  OR2X1    g00131(.A(new_n382_), .B(new_n387_), .Y(new_n388_));
  OAI21X1  g00132(.A0(new_n383_), .A1(new_n361_), .B0(new_n388_), .Y(new_n389_));
  AND2X1   g00133(.A(\b[6] ), .B(\b[5] ), .Y(new_n390_));
  AOI21X1  g00134(.A0(new_n377_), .A1(new_n376_), .B0(new_n390_), .Y(new_n391_));
  INVX1    g00135(.A(\b[6] ), .Y(new_n392_));
  XOR2X1   g00136(.A(\b[7] ), .B(new_n392_), .Y(new_n393_));
  XOR2X1   g00137(.A(new_n393_), .B(new_n391_), .Y(new_n394_));
  INVX1    g00138(.A(\b[5] ), .Y(new_n395_));
  AOI22X1  g00139(.A0(new_n267_), .A1(\b[7] ), .B0(new_n266_), .B1(\b[6] ), .Y(new_n396_));
  OAI21X1  g00140(.A0(new_n350_), .A1(new_n395_), .B0(new_n396_), .Y(new_n397_));
  AOI21X1  g00141(.A0(new_n394_), .A1(new_n318_), .B0(new_n397_), .Y(new_n398_));
  XOR2X1   g00142(.A(new_n398_), .B(new_n257_), .Y(new_n399_));
  INVX1    g00143(.A(\a[8] ), .Y(new_n400_));
  AOI21X1  g00144(.A0(new_n363_), .A1(\b[0] ), .B0(new_n400_), .Y(new_n401_));
  INVX1    g00145(.A(new_n401_), .Y(new_n402_));
  XOR2X1   g00146(.A(\a[8] ), .B(\a[7] ), .Y(new_n403_));
  AND2X1   g00147(.A(new_n403_), .B(new_n363_), .Y(new_n404_));
  AND2X1   g00148(.A(new_n404_), .B(new_n263_), .Y(new_n405_));
  INVX1    g00149(.A(\a[6] ), .Y(new_n406_));
  XOR2X1   g00150(.A(\a[7] ), .B(new_n406_), .Y(new_n407_));
  NOR3X1   g00151(.A(new_n407_), .B(new_n363_), .C(new_n274_), .Y(new_n408_));
  XOR2X1   g00152(.A(\a[6] ), .B(new_n305_), .Y(new_n409_));
  NOR3X1   g00153(.A(new_n403_), .B(new_n409_), .C(new_n275_), .Y(new_n410_));
  NOR3X1   g00154(.A(new_n410_), .B(new_n408_), .C(new_n405_), .Y(new_n411_));
  XOR2X1   g00155(.A(new_n411_), .B(\a[8] ), .Y(new_n412_));
  XOR2X1   g00156(.A(new_n412_), .B(new_n402_), .Y(new_n413_));
  AND2X1   g00157(.A(new_n323_), .B(new_n308_), .Y(new_n414_));
  NOR4X1   g00158(.A(new_n336_), .B(new_n335_), .C(new_n301_), .D(new_n277_), .Y(new_n415_));
  NAND2X1  g00159(.A(new_n336_), .B(new_n313_), .Y(new_n416_));
  NAND3X1  g00160(.A(new_n335_), .B(new_n301_), .C(\b[4] ), .Y(new_n417_));
  OAI21X1  g00161(.A0(new_n416_), .A1(new_n297_), .B0(new_n417_), .Y(new_n418_));
  NOR3X1   g00162(.A(new_n418_), .B(new_n415_), .C(new_n414_), .Y(new_n419_));
  XOR2X1   g00163(.A(new_n419_), .B(\a[5] ), .Y(new_n420_));
  XOR2X1   g00164(.A(new_n420_), .B(new_n413_), .Y(new_n421_));
  AND2X1   g00165(.A(new_n364_), .B(new_n385_), .Y(new_n422_));
  XOR2X1   g00166(.A(new_n372_), .B(new_n305_), .Y(new_n423_));
  AOI21X1  g00167(.A0(new_n423_), .A1(new_n386_), .B0(new_n422_), .Y(new_n424_));
  XOR2X1   g00168(.A(new_n424_), .B(new_n421_), .Y(new_n425_));
  XOR2X1   g00169(.A(new_n425_), .B(new_n399_), .Y(new_n426_));
  XOR2X1   g00170(.A(new_n426_), .B(new_n389_), .Y(\f[7] ));
  NOR2X1   g00171(.A(new_n412_), .B(new_n402_), .Y(new_n428_));
  INVX1    g00172(.A(new_n404_), .Y(new_n429_));
  XOR2X1   g00173(.A(new_n400_), .B(\a[7] ), .Y(new_n430_));
  XOR2X1   g00174(.A(\a[7] ), .B(\a[6] ), .Y(new_n431_));
  NOR4X1   g00175(.A(new_n431_), .B(new_n430_), .C(new_n363_), .D(new_n274_), .Y(new_n432_));
  NOR3X1   g00176(.A(new_n403_), .B(new_n409_), .C(new_n277_), .Y(new_n433_));
  NOR3X1   g00177(.A(new_n407_), .B(new_n363_), .C(new_n275_), .Y(new_n434_));
  NOR3X1   g00178(.A(new_n434_), .B(new_n433_), .C(new_n432_), .Y(new_n435_));
  OAI21X1  g00179(.A0(new_n429_), .A1(new_n281_), .B0(new_n435_), .Y(new_n436_));
  XOR2X1   g00180(.A(new_n436_), .B(new_n400_), .Y(new_n437_));
  XOR2X1   g00181(.A(new_n437_), .B(new_n428_), .Y(new_n438_));
  AOI22X1  g00182(.A0(new_n369_), .A1(\b[5] ), .B0(new_n368_), .B1(\b[4] ), .Y(new_n439_));
  OAI21X1  g00183(.A0(new_n367_), .A1(new_n297_), .B0(new_n439_), .Y(new_n440_));
  AOI21X1  g00184(.A0(new_n349_), .A1(new_n308_), .B0(new_n440_), .Y(new_n441_));
  XOR2X1   g00185(.A(new_n441_), .B(new_n305_), .Y(new_n442_));
  XOR2X1   g00186(.A(new_n442_), .B(new_n438_), .Y(new_n443_));
  XOR2X1   g00187(.A(new_n412_), .B(new_n401_), .Y(new_n444_));
  NOR2X1   g00188(.A(new_n420_), .B(new_n444_), .Y(new_n445_));
  XOR2X1   g00189(.A(new_n420_), .B(new_n444_), .Y(new_n446_));
  NAND2X1  g00190(.A(new_n364_), .B(new_n385_), .Y(new_n447_));
  OAI21X1  g00191(.A0(new_n373_), .A1(new_n365_), .B0(new_n447_), .Y(new_n448_));
  AOI21X1  g00192(.A0(new_n448_), .A1(new_n446_), .B0(new_n445_), .Y(new_n449_));
  XOR2X1   g00193(.A(new_n449_), .B(new_n443_), .Y(new_n450_));
  NAND2X1  g00194(.A(\b[7] ), .B(\b[6] ), .Y(new_n451_));
  OAI21X1  g00195(.A0(new_n393_), .A1(new_n391_), .B0(new_n451_), .Y(new_n452_));
  XOR2X1   g00196(.A(\b[8] ), .B(\b[7] ), .Y(new_n453_));
  XOR2X1   g00197(.A(new_n453_), .B(new_n452_), .Y(new_n454_));
  AOI22X1  g00198(.A0(new_n267_), .A1(\b[8] ), .B0(new_n266_), .B1(\b[7] ), .Y(new_n455_));
  OAI21X1  g00199(.A0(new_n350_), .A1(new_n392_), .B0(new_n455_), .Y(new_n456_));
  AOI21X1  g00200(.A0(new_n454_), .A1(new_n318_), .B0(new_n456_), .Y(new_n457_));
  XOR2X1   g00201(.A(new_n457_), .B(\a[2] ), .Y(new_n458_));
  XOR2X1   g00202(.A(new_n458_), .B(new_n450_), .Y(new_n459_));
  AND2X1   g00203(.A(new_n425_), .B(new_n399_), .Y(new_n460_));
  AOI21X1  g00204(.A0(new_n426_), .A1(new_n389_), .B0(new_n460_), .Y(new_n461_));
  XOR2X1   g00205(.A(new_n461_), .B(new_n459_), .Y(\f[8] ));
  NOR4X1   g00206(.A(new_n436_), .B(new_n412_), .C(new_n364_), .D(new_n400_), .Y(new_n463_));
  XOR2X1   g00207(.A(\a[9] ), .B(\a[8] ), .Y(new_n464_));
  AND2X1   g00208(.A(new_n464_), .B(\b[0] ), .Y(new_n465_));
  XOR2X1   g00209(.A(new_n465_), .B(new_n463_), .Y(new_n466_));
  NAND3X1  g00210(.A(new_n407_), .B(new_n403_), .C(new_n409_), .Y(new_n467_));
  AND2X1   g00211(.A(new_n431_), .B(new_n409_), .Y(new_n468_));
  AND2X1   g00212(.A(new_n430_), .B(new_n363_), .Y(new_n469_));
  AOI22X1  g00213(.A0(new_n469_), .A1(\b[3] ), .B0(new_n468_), .B1(\b[2] ), .Y(new_n470_));
  OAI21X1  g00214(.A0(new_n467_), .A1(new_n275_), .B0(new_n470_), .Y(new_n471_));
  AOI21X1  g00215(.A0(new_n404_), .A1(new_n366_), .B0(new_n471_), .Y(new_n472_));
  XOR2X1   g00216(.A(new_n472_), .B(\a[8] ), .Y(new_n473_));
  XOR2X1   g00217(.A(new_n473_), .B(new_n466_), .Y(new_n474_));
  AOI22X1  g00218(.A0(new_n369_), .A1(\b[6] ), .B0(new_n368_), .B1(\b[5] ), .Y(new_n475_));
  OAI21X1  g00219(.A0(new_n367_), .A1(new_n325_), .B0(new_n475_), .Y(new_n476_));
  AOI21X1  g00220(.A0(new_n378_), .A1(new_n308_), .B0(new_n476_), .Y(new_n477_));
  XOR2X1   g00221(.A(new_n477_), .B(\a[5] ), .Y(new_n478_));
  XOR2X1   g00222(.A(new_n478_), .B(new_n474_), .Y(new_n479_));
  XOR2X1   g00223(.A(new_n441_), .B(\a[5] ), .Y(new_n480_));
  NOR2X1   g00224(.A(new_n480_), .B(new_n438_), .Y(new_n481_));
  XOR2X1   g00225(.A(new_n480_), .B(new_n438_), .Y(new_n482_));
  OR2X1    g00226(.A(new_n420_), .B(new_n444_), .Y(new_n483_));
  OAI21X1  g00227(.A0(new_n424_), .A1(new_n421_), .B0(new_n483_), .Y(new_n484_));
  AOI21X1  g00228(.A0(new_n484_), .A1(new_n482_), .B0(new_n481_), .Y(new_n485_));
  XOR2X1   g00229(.A(new_n485_), .B(new_n479_), .Y(new_n486_));
  AND2X1   g00230(.A(\b[8] ), .B(\b[7] ), .Y(new_n487_));
  AOI21X1  g00231(.A0(new_n453_), .A1(new_n452_), .B0(new_n487_), .Y(new_n488_));
  INVX1    g00232(.A(\b[8] ), .Y(new_n489_));
  XOR2X1   g00233(.A(\b[9] ), .B(new_n489_), .Y(new_n490_));
  XOR2X1   g00234(.A(new_n490_), .B(new_n488_), .Y(new_n491_));
  INVX1    g00235(.A(\b[7] ), .Y(new_n492_));
  AOI22X1  g00236(.A0(new_n267_), .A1(\b[9] ), .B0(new_n266_), .B1(\b[8] ), .Y(new_n493_));
  OAI21X1  g00237(.A0(new_n350_), .A1(new_n492_), .B0(new_n493_), .Y(new_n494_));
  AOI21X1  g00238(.A0(new_n491_), .A1(new_n318_), .B0(new_n494_), .Y(new_n495_));
  XOR2X1   g00239(.A(new_n495_), .B(\a[2] ), .Y(new_n496_));
  XOR2X1   g00240(.A(new_n496_), .B(new_n486_), .Y(new_n497_));
  XOR2X1   g00241(.A(new_n449_), .B(new_n482_), .Y(new_n498_));
  OR2X1    g00242(.A(new_n458_), .B(new_n498_), .Y(new_n499_));
  OAI21X1  g00243(.A0(new_n461_), .A1(new_n459_), .B0(new_n499_), .Y(new_n500_));
  XOR2X1   g00244(.A(new_n500_), .B(new_n497_), .Y(\f[9] ));
  NOR2X1   g00245(.A(new_n496_), .B(new_n486_), .Y(new_n502_));
  AOI21X1  g00246(.A0(new_n500_), .A1(new_n497_), .B0(new_n502_), .Y(new_n503_));
  OR4X1    g00247(.A(new_n436_), .B(new_n412_), .C(new_n364_), .D(new_n400_), .Y(new_n504_));
  XOR2X1   g00248(.A(new_n465_), .B(new_n504_), .Y(new_n505_));
  NAND2X1  g00249(.A(new_n465_), .B(new_n463_), .Y(new_n506_));
  OAI21X1  g00250(.A0(new_n473_), .A1(new_n505_), .B0(new_n506_), .Y(new_n507_));
  AND2X1   g00251(.A(new_n404_), .B(new_n323_), .Y(new_n508_));
  NOR4X1   g00252(.A(new_n431_), .B(new_n430_), .C(new_n363_), .D(new_n277_), .Y(new_n509_));
  NAND2X1  g00253(.A(new_n431_), .B(new_n409_), .Y(new_n510_));
  NAND2X1  g00254(.A(new_n430_), .B(new_n363_), .Y(new_n511_));
  OAI22X1  g00255(.A0(new_n511_), .A1(new_n325_), .B0(new_n510_), .B1(new_n297_), .Y(new_n512_));
  NOR3X1   g00256(.A(new_n512_), .B(new_n509_), .C(new_n508_), .Y(new_n513_));
  XOR2X1   g00257(.A(new_n513_), .B(new_n400_), .Y(new_n514_));
  INVX1    g00258(.A(\a[11] ), .Y(new_n515_));
  OR2X1    g00259(.A(new_n465_), .B(new_n515_), .Y(new_n516_));
  XOR2X1   g00260(.A(\a[11] ), .B(\a[10] ), .Y(new_n517_));
  AND2X1   g00261(.A(new_n517_), .B(new_n464_), .Y(new_n518_));
  AND2X1   g00262(.A(new_n518_), .B(new_n263_), .Y(new_n519_));
  INVX1    g00263(.A(\a[9] ), .Y(new_n520_));
  XOR2X1   g00264(.A(\a[10] ), .B(new_n520_), .Y(new_n521_));
  NOR3X1   g00265(.A(new_n521_), .B(new_n464_), .C(new_n274_), .Y(new_n522_));
  XOR2X1   g00266(.A(\a[9] ), .B(new_n400_), .Y(new_n523_));
  NOR3X1   g00267(.A(new_n517_), .B(new_n523_), .C(new_n275_), .Y(new_n524_));
  NOR3X1   g00268(.A(new_n524_), .B(new_n522_), .C(new_n519_), .Y(new_n525_));
  XOR2X1   g00269(.A(new_n525_), .B(\a[11] ), .Y(new_n526_));
  XOR2X1   g00270(.A(new_n526_), .B(new_n516_), .Y(new_n527_));
  XOR2X1   g00271(.A(new_n527_), .B(new_n514_), .Y(new_n528_));
  XOR2X1   g00272(.A(new_n528_), .B(new_n507_), .Y(new_n529_));
  AOI22X1  g00273(.A0(new_n369_), .A1(\b[7] ), .B0(new_n368_), .B1(\b[6] ), .Y(new_n530_));
  OAI21X1  g00274(.A0(new_n367_), .A1(new_n395_), .B0(new_n530_), .Y(new_n531_));
  AOI21X1  g00275(.A0(new_n394_), .A1(new_n308_), .B0(new_n531_), .Y(new_n532_));
  XOR2X1   g00276(.A(new_n532_), .B(\a[5] ), .Y(new_n533_));
  XOR2X1   g00277(.A(new_n533_), .B(new_n529_), .Y(new_n534_));
  NOR2X1   g00278(.A(new_n478_), .B(new_n474_), .Y(new_n535_));
  OR2X1    g00279(.A(new_n480_), .B(new_n438_), .Y(new_n536_));
  OAI21X1  g00280(.A0(new_n449_), .A1(new_n443_), .B0(new_n536_), .Y(new_n537_));
  AOI21X1  g00281(.A0(new_n537_), .A1(new_n479_), .B0(new_n535_), .Y(new_n538_));
  XOR2X1   g00282(.A(new_n538_), .B(new_n534_), .Y(new_n539_));
  NAND2X1  g00283(.A(\b[9] ), .B(\b[8] ), .Y(new_n540_));
  OAI21X1  g00284(.A0(new_n490_), .A1(new_n488_), .B0(new_n540_), .Y(new_n541_));
  XOR2X1   g00285(.A(\b[10] ), .B(\b[9] ), .Y(new_n542_));
  XOR2X1   g00286(.A(new_n542_), .B(new_n541_), .Y(new_n543_));
  AOI22X1  g00287(.A0(new_n267_), .A1(\b[10] ), .B0(new_n266_), .B1(\b[9] ), .Y(new_n544_));
  OAI21X1  g00288(.A0(new_n350_), .A1(new_n489_), .B0(new_n544_), .Y(new_n545_));
  AOI21X1  g00289(.A0(new_n543_), .A1(new_n318_), .B0(new_n545_), .Y(new_n546_));
  XOR2X1   g00290(.A(new_n546_), .B(\a[2] ), .Y(new_n547_));
  XOR2X1   g00291(.A(new_n547_), .B(new_n539_), .Y(new_n548_));
  XOR2X1   g00292(.A(new_n548_), .B(new_n503_), .Y(\f[10] ));
  XOR2X1   g00293(.A(new_n472_), .B(new_n400_), .Y(new_n550_));
  AND2X1   g00294(.A(new_n465_), .B(new_n463_), .Y(new_n551_));
  AOI21X1  g00295(.A0(new_n550_), .A1(new_n466_), .B0(new_n551_), .Y(new_n552_));
  XOR2X1   g00296(.A(new_n528_), .B(new_n552_), .Y(new_n553_));
  XOR2X1   g00297(.A(new_n533_), .B(new_n553_), .Y(new_n554_));
  XOR2X1   g00298(.A(new_n538_), .B(new_n554_), .Y(new_n555_));
  OR2X1    g00299(.A(new_n547_), .B(new_n555_), .Y(new_n556_));
  OAI21X1  g00300(.A0(new_n548_), .A1(new_n503_), .B0(new_n556_), .Y(new_n557_));
  OR2X1    g00301(.A(new_n533_), .B(new_n553_), .Y(new_n558_));
  OAI21X1  g00302(.A0(new_n538_), .A1(new_n534_), .B0(new_n558_), .Y(new_n559_));
  AOI22X1  g00303(.A0(new_n369_), .A1(\b[8] ), .B0(new_n368_), .B1(\b[7] ), .Y(new_n560_));
  OAI21X1  g00304(.A0(new_n367_), .A1(new_n392_), .B0(new_n560_), .Y(new_n561_));
  AOI21X1  g00305(.A0(new_n454_), .A1(new_n308_), .B0(new_n561_), .Y(new_n562_));
  XOR2X1   g00306(.A(new_n562_), .B(\a[5] ), .Y(new_n563_));
  AND2X1   g00307(.A(new_n527_), .B(new_n514_), .Y(new_n564_));
  AOI21X1  g00308(.A0(new_n528_), .A1(new_n507_), .B0(new_n564_), .Y(new_n565_));
  NOR2X1   g00309(.A(new_n526_), .B(new_n516_), .Y(new_n566_));
  INVX1    g00310(.A(new_n518_), .Y(new_n567_));
  XOR2X1   g00311(.A(new_n515_), .B(\a[10] ), .Y(new_n568_));
  XOR2X1   g00312(.A(\a[10] ), .B(\a[9] ), .Y(new_n569_));
  NOR4X1   g00313(.A(new_n569_), .B(new_n568_), .C(new_n464_), .D(new_n274_), .Y(new_n570_));
  NOR3X1   g00314(.A(new_n517_), .B(new_n523_), .C(new_n277_), .Y(new_n571_));
  NOR3X1   g00315(.A(new_n521_), .B(new_n464_), .C(new_n275_), .Y(new_n572_));
  NOR3X1   g00316(.A(new_n572_), .B(new_n571_), .C(new_n570_), .Y(new_n573_));
  OAI21X1  g00317(.A0(new_n567_), .A1(new_n281_), .B0(new_n573_), .Y(new_n574_));
  XOR2X1   g00318(.A(new_n574_), .B(new_n515_), .Y(new_n575_));
  XOR2X1   g00319(.A(new_n575_), .B(new_n566_), .Y(new_n576_));
  AOI22X1  g00320(.A0(new_n469_), .A1(\b[5] ), .B0(new_n468_), .B1(\b[4] ), .Y(new_n577_));
  OAI21X1  g00321(.A0(new_n467_), .A1(new_n297_), .B0(new_n577_), .Y(new_n578_));
  AOI21X1  g00322(.A0(new_n404_), .A1(new_n349_), .B0(new_n578_), .Y(new_n579_));
  XOR2X1   g00323(.A(new_n579_), .B(new_n400_), .Y(new_n580_));
  XOR2X1   g00324(.A(new_n580_), .B(new_n576_), .Y(new_n581_));
  XOR2X1   g00325(.A(new_n581_), .B(new_n565_), .Y(new_n582_));
  XOR2X1   g00326(.A(new_n582_), .B(new_n563_), .Y(new_n583_));
  XOR2X1   g00327(.A(new_n583_), .B(new_n559_), .Y(new_n584_));
  AND2X1   g00328(.A(\b[10] ), .B(\b[9] ), .Y(new_n585_));
  AOI21X1  g00329(.A0(new_n542_), .A1(new_n541_), .B0(new_n585_), .Y(new_n586_));
  INVX1    g00330(.A(\b[10] ), .Y(new_n587_));
  XOR2X1   g00331(.A(\b[11] ), .B(new_n587_), .Y(new_n588_));
  XOR2X1   g00332(.A(new_n588_), .B(new_n586_), .Y(new_n589_));
  INVX1    g00333(.A(\b[9] ), .Y(new_n590_));
  AOI22X1  g00334(.A0(new_n267_), .A1(\b[11] ), .B0(new_n266_), .B1(\b[10] ), .Y(new_n591_));
  OAI21X1  g00335(.A0(new_n350_), .A1(new_n590_), .B0(new_n591_), .Y(new_n592_));
  AOI21X1  g00336(.A0(new_n589_), .A1(new_n318_), .B0(new_n592_), .Y(new_n593_));
  XOR2X1   g00337(.A(new_n593_), .B(\a[2] ), .Y(new_n594_));
  XOR2X1   g00338(.A(new_n594_), .B(new_n584_), .Y(new_n595_));
  XOR2X1   g00339(.A(new_n595_), .B(new_n557_), .Y(\f[11] ));
  OR4X1    g00340(.A(new_n574_), .B(new_n526_), .C(new_n465_), .D(new_n515_), .Y(new_n597_));
  XOR2X1   g00341(.A(\a[12] ), .B(\a[11] ), .Y(new_n598_));
  AND2X1   g00342(.A(new_n598_), .B(\b[0] ), .Y(new_n599_));
  XOR2X1   g00343(.A(new_n599_), .B(new_n597_), .Y(new_n600_));
  NAND3X1  g00344(.A(new_n521_), .B(new_n517_), .C(new_n523_), .Y(new_n601_));
  AND2X1   g00345(.A(new_n569_), .B(new_n523_), .Y(new_n602_));
  AND2X1   g00346(.A(new_n568_), .B(new_n464_), .Y(new_n603_));
  AOI22X1  g00347(.A0(new_n603_), .A1(\b[3] ), .B0(new_n602_), .B1(\b[2] ), .Y(new_n604_));
  OAI21X1  g00348(.A0(new_n601_), .A1(new_n275_), .B0(new_n604_), .Y(new_n605_));
  AOI21X1  g00349(.A0(new_n518_), .A1(new_n366_), .B0(new_n605_), .Y(new_n606_));
  XOR2X1   g00350(.A(new_n606_), .B(\a[11] ), .Y(new_n607_));
  XOR2X1   g00351(.A(new_n607_), .B(new_n600_), .Y(new_n608_));
  AOI22X1  g00352(.A0(new_n469_), .A1(\b[6] ), .B0(new_n468_), .B1(\b[5] ), .Y(new_n609_));
  OAI21X1  g00353(.A0(new_n467_), .A1(new_n325_), .B0(new_n609_), .Y(new_n610_));
  AOI21X1  g00354(.A0(new_n404_), .A1(new_n378_), .B0(new_n610_), .Y(new_n611_));
  XOR2X1   g00355(.A(new_n611_), .B(\a[8] ), .Y(new_n612_));
  XOR2X1   g00356(.A(new_n612_), .B(new_n608_), .Y(new_n613_));
  NOR2X1   g00357(.A(new_n527_), .B(new_n514_), .Y(new_n614_));
  NAND2X1  g00358(.A(new_n527_), .B(new_n514_), .Y(new_n615_));
  OAI21X1  g00359(.A0(new_n614_), .A1(new_n552_), .B0(new_n615_), .Y(new_n616_));
  XOR2X1   g00360(.A(new_n579_), .B(\a[8] ), .Y(new_n617_));
  NOR2X1   g00361(.A(new_n617_), .B(new_n576_), .Y(new_n618_));
  XOR2X1   g00362(.A(new_n617_), .B(new_n576_), .Y(new_n619_));
  AOI21X1  g00363(.A0(new_n619_), .A1(new_n616_), .B0(new_n618_), .Y(new_n620_));
  XOR2X1   g00364(.A(new_n620_), .B(new_n613_), .Y(new_n621_));
  AOI22X1  g00365(.A0(new_n369_), .A1(\b[9] ), .B0(new_n368_), .B1(\b[8] ), .Y(new_n622_));
  OAI21X1  g00366(.A0(new_n367_), .A1(new_n492_), .B0(new_n622_), .Y(new_n623_));
  AOI21X1  g00367(.A0(new_n491_), .A1(new_n308_), .B0(new_n623_), .Y(new_n624_));
  XOR2X1   g00368(.A(new_n624_), .B(\a[5] ), .Y(new_n625_));
  XOR2X1   g00369(.A(new_n625_), .B(new_n621_), .Y(new_n626_));
  INVX1    g00370(.A(new_n563_), .Y(new_n627_));
  AND2X1   g00371(.A(new_n582_), .B(new_n627_), .Y(new_n628_));
  XOR2X1   g00372(.A(new_n582_), .B(new_n627_), .Y(new_n629_));
  AOI21X1  g00373(.A0(new_n629_), .A1(new_n559_), .B0(new_n628_), .Y(new_n630_));
  XOR2X1   g00374(.A(new_n630_), .B(new_n626_), .Y(new_n631_));
  NAND2X1  g00375(.A(\b[11] ), .B(\b[10] ), .Y(new_n632_));
  OAI21X1  g00376(.A0(new_n588_), .A1(new_n586_), .B0(new_n632_), .Y(new_n633_));
  XOR2X1   g00377(.A(\b[12] ), .B(\b[11] ), .Y(new_n634_));
  XOR2X1   g00378(.A(new_n634_), .B(new_n633_), .Y(new_n635_));
  AOI22X1  g00379(.A0(new_n267_), .A1(\b[12] ), .B0(new_n266_), .B1(\b[11] ), .Y(new_n636_));
  OAI21X1  g00380(.A0(new_n350_), .A1(new_n587_), .B0(new_n636_), .Y(new_n637_));
  AOI21X1  g00381(.A0(new_n635_), .A1(new_n318_), .B0(new_n637_), .Y(new_n638_));
  XOR2X1   g00382(.A(new_n638_), .B(\a[2] ), .Y(new_n639_));
  XOR2X1   g00383(.A(new_n639_), .B(new_n631_), .Y(new_n640_));
  NOR2X1   g00384(.A(new_n594_), .B(new_n584_), .Y(new_n641_));
  AOI21X1  g00385(.A0(new_n595_), .A1(new_n557_), .B0(new_n641_), .Y(new_n642_));
  XOR2X1   g00386(.A(new_n642_), .B(new_n640_), .Y(\f[12] ));
  NOR4X1   g00387(.A(new_n574_), .B(new_n526_), .C(new_n465_), .D(new_n515_), .Y(new_n644_));
  XOR2X1   g00388(.A(new_n599_), .B(new_n644_), .Y(new_n645_));
  XOR2X1   g00389(.A(new_n607_), .B(new_n645_), .Y(new_n646_));
  XOR2X1   g00390(.A(new_n612_), .B(new_n646_), .Y(new_n647_));
  XOR2X1   g00391(.A(new_n620_), .B(new_n647_), .Y(new_n648_));
  XOR2X1   g00392(.A(new_n625_), .B(new_n648_), .Y(new_n649_));
  XOR2X1   g00393(.A(new_n630_), .B(new_n649_), .Y(new_n650_));
  OR2X1    g00394(.A(new_n639_), .B(new_n650_), .Y(new_n651_));
  OAI21X1  g00395(.A0(new_n642_), .A1(new_n640_), .B0(new_n651_), .Y(new_n652_));
  OR2X1    g00396(.A(new_n625_), .B(new_n648_), .Y(new_n653_));
  OAI21X1  g00397(.A0(new_n630_), .A1(new_n626_), .B0(new_n653_), .Y(new_n654_));
  XOR2X1   g00398(.A(new_n606_), .B(new_n515_), .Y(new_n655_));
  AND2X1   g00399(.A(new_n599_), .B(new_n644_), .Y(new_n656_));
  AOI21X1  g00400(.A0(new_n655_), .A1(new_n645_), .B0(new_n656_), .Y(new_n657_));
  AND2X1   g00401(.A(new_n518_), .B(new_n323_), .Y(new_n658_));
  NOR4X1   g00402(.A(new_n569_), .B(new_n568_), .C(new_n464_), .D(new_n277_), .Y(new_n659_));
  NAND2X1  g00403(.A(new_n569_), .B(new_n523_), .Y(new_n660_));
  NAND2X1  g00404(.A(new_n568_), .B(new_n464_), .Y(new_n661_));
  OAI22X1  g00405(.A0(new_n661_), .A1(new_n325_), .B0(new_n660_), .B1(new_n297_), .Y(new_n662_));
  NOR3X1   g00406(.A(new_n662_), .B(new_n659_), .C(new_n658_), .Y(new_n663_));
  XOR2X1   g00407(.A(new_n663_), .B(new_n515_), .Y(new_n664_));
  INVX1    g00408(.A(\a[14] ), .Y(new_n665_));
  OR2X1    g00409(.A(new_n599_), .B(new_n665_), .Y(new_n666_));
  XOR2X1   g00410(.A(\a[14] ), .B(\a[13] ), .Y(new_n667_));
  AND2X1   g00411(.A(new_n667_), .B(new_n598_), .Y(new_n668_));
  AND2X1   g00412(.A(new_n668_), .B(new_n263_), .Y(new_n669_));
  INVX1    g00413(.A(\a[12] ), .Y(new_n670_));
  XOR2X1   g00414(.A(\a[13] ), .B(new_n670_), .Y(new_n671_));
  NOR3X1   g00415(.A(new_n671_), .B(new_n598_), .C(new_n274_), .Y(new_n672_));
  XOR2X1   g00416(.A(\a[12] ), .B(new_n515_), .Y(new_n673_));
  NOR3X1   g00417(.A(new_n667_), .B(new_n673_), .C(new_n275_), .Y(new_n674_));
  NOR3X1   g00418(.A(new_n674_), .B(new_n672_), .C(new_n669_), .Y(new_n675_));
  XOR2X1   g00419(.A(new_n675_), .B(\a[14] ), .Y(new_n676_));
  XOR2X1   g00420(.A(new_n676_), .B(new_n666_), .Y(new_n677_));
  XOR2X1   g00421(.A(new_n677_), .B(new_n664_), .Y(new_n678_));
  XOR2X1   g00422(.A(new_n678_), .B(new_n657_), .Y(new_n679_));
  AOI22X1  g00423(.A0(new_n469_), .A1(\b[7] ), .B0(new_n468_), .B1(\b[6] ), .Y(new_n680_));
  OAI21X1  g00424(.A0(new_n467_), .A1(new_n395_), .B0(new_n680_), .Y(new_n681_));
  AOI21X1  g00425(.A0(new_n404_), .A1(new_n394_), .B0(new_n681_), .Y(new_n682_));
  XOR2X1   g00426(.A(new_n682_), .B(\a[8] ), .Y(new_n683_));
  XOR2X1   g00427(.A(new_n683_), .B(new_n679_), .Y(new_n684_));
  NOR2X1   g00428(.A(new_n612_), .B(new_n646_), .Y(new_n685_));
  OR2X1    g00429(.A(new_n617_), .B(new_n576_), .Y(new_n686_));
  OAI21X1  g00430(.A0(new_n581_), .A1(new_n565_), .B0(new_n686_), .Y(new_n687_));
  AOI21X1  g00431(.A0(new_n687_), .A1(new_n647_), .B0(new_n685_), .Y(new_n688_));
  XOR2X1   g00432(.A(new_n688_), .B(new_n684_), .Y(new_n689_));
  AOI22X1  g00433(.A0(new_n369_), .A1(\b[10] ), .B0(new_n368_), .B1(\b[9] ), .Y(new_n690_));
  OAI21X1  g00434(.A0(new_n367_), .A1(new_n489_), .B0(new_n690_), .Y(new_n691_));
  AOI21X1  g00435(.A0(new_n543_), .A1(new_n308_), .B0(new_n691_), .Y(new_n692_));
  XOR2X1   g00436(.A(new_n692_), .B(\a[5] ), .Y(new_n693_));
  NOR2X1   g00437(.A(new_n693_), .B(new_n689_), .Y(new_n694_));
  AND2X1   g00438(.A(new_n693_), .B(new_n689_), .Y(new_n695_));
  OR2X1    g00439(.A(new_n695_), .B(new_n694_), .Y(new_n696_));
  NAND2X1  g00440(.A(new_n696_), .B(new_n654_), .Y(new_n697_));
  NOR2X1   g00441(.A(new_n625_), .B(new_n648_), .Y(new_n698_));
  NOR2X1   g00442(.A(new_n533_), .B(new_n553_), .Y(new_n699_));
  OR2X1    g00443(.A(new_n478_), .B(new_n474_), .Y(new_n700_));
  XOR2X1   g00444(.A(new_n473_), .B(new_n505_), .Y(new_n701_));
  XOR2X1   g00445(.A(new_n478_), .B(new_n701_), .Y(new_n702_));
  OAI21X1  g00446(.A0(new_n485_), .A1(new_n702_), .B0(new_n700_), .Y(new_n703_));
  AOI21X1  g00447(.A0(new_n703_), .A1(new_n554_), .B0(new_n699_), .Y(new_n704_));
  NAND2X1  g00448(.A(new_n582_), .B(new_n627_), .Y(new_n705_));
  OAI21X1  g00449(.A0(new_n583_), .A1(new_n704_), .B0(new_n705_), .Y(new_n706_));
  AOI21X1  g00450(.A0(new_n706_), .A1(new_n649_), .B0(new_n698_), .Y(new_n707_));
  OR2X1    g00451(.A(new_n693_), .B(new_n689_), .Y(new_n708_));
  NAND2X1  g00452(.A(new_n693_), .B(new_n689_), .Y(new_n709_));
  NAND3X1  g00453(.A(new_n709_), .B(new_n708_), .C(new_n707_), .Y(new_n710_));
  AND2X1   g00454(.A(\b[12] ), .B(\b[11] ), .Y(new_n711_));
  AOI21X1  g00455(.A0(new_n634_), .A1(new_n633_), .B0(new_n711_), .Y(new_n712_));
  INVX1    g00456(.A(\b[12] ), .Y(new_n713_));
  XOR2X1   g00457(.A(\b[13] ), .B(new_n713_), .Y(new_n714_));
  XOR2X1   g00458(.A(new_n714_), .B(new_n712_), .Y(new_n715_));
  INVX1    g00459(.A(\b[11] ), .Y(new_n716_));
  AOI22X1  g00460(.A0(new_n267_), .A1(\b[13] ), .B0(new_n266_), .B1(\b[12] ), .Y(new_n717_));
  OAI21X1  g00461(.A0(new_n350_), .A1(new_n716_), .B0(new_n717_), .Y(new_n718_));
  AOI21X1  g00462(.A0(new_n715_), .A1(new_n318_), .B0(new_n718_), .Y(new_n719_));
  XOR2X1   g00463(.A(new_n719_), .B(new_n257_), .Y(new_n720_));
  AOI21X1  g00464(.A0(new_n710_), .A1(new_n697_), .B0(new_n720_), .Y(new_n721_));
  AND2X1   g00465(.A(new_n696_), .B(new_n654_), .Y(new_n722_));
  NOR3X1   g00466(.A(new_n695_), .B(new_n694_), .C(new_n654_), .Y(new_n723_));
  XOR2X1   g00467(.A(new_n719_), .B(\a[2] ), .Y(new_n724_));
  NOR3X1   g00468(.A(new_n724_), .B(new_n723_), .C(new_n722_), .Y(new_n725_));
  OR2X1    g00469(.A(new_n725_), .B(new_n721_), .Y(new_n726_));
  XOR2X1   g00470(.A(new_n726_), .B(new_n652_), .Y(\f[13] ));
  OAI21X1  g00471(.A0(new_n725_), .A1(new_n721_), .B0(new_n652_), .Y(new_n728_));
  OAI21X1  g00472(.A0(new_n723_), .A1(new_n722_), .B0(new_n720_), .Y(new_n729_));
  AND2X1   g00473(.A(new_n729_), .B(new_n728_), .Y(new_n730_));
  NAND2X1  g00474(.A(\b[13] ), .B(\b[12] ), .Y(new_n731_));
  OAI21X1  g00475(.A0(new_n714_), .A1(new_n712_), .B0(new_n731_), .Y(new_n732_));
  XOR2X1   g00476(.A(\b[14] ), .B(\b[13] ), .Y(new_n733_));
  XOR2X1   g00477(.A(new_n733_), .B(new_n732_), .Y(new_n734_));
  AOI22X1  g00478(.A0(new_n267_), .A1(\b[14] ), .B0(new_n266_), .B1(\b[13] ), .Y(new_n735_));
  OAI21X1  g00479(.A0(new_n350_), .A1(new_n713_), .B0(new_n735_), .Y(new_n736_));
  AOI21X1  g00480(.A0(new_n734_), .A1(new_n318_), .B0(new_n736_), .Y(new_n737_));
  XOR2X1   g00481(.A(new_n737_), .B(\a[2] ), .Y(new_n738_));
  OAI21X1  g00482(.A0(new_n695_), .A1(new_n707_), .B0(new_n708_), .Y(new_n739_));
  AOI22X1  g00483(.A0(new_n369_), .A1(\b[11] ), .B0(new_n368_), .B1(\b[10] ), .Y(new_n740_));
  OAI21X1  g00484(.A0(new_n367_), .A1(new_n590_), .B0(new_n740_), .Y(new_n741_));
  AOI21X1  g00485(.A0(new_n589_), .A1(new_n308_), .B0(new_n741_), .Y(new_n742_));
  XOR2X1   g00486(.A(new_n742_), .B(new_n305_), .Y(new_n743_));
  OR2X1    g00487(.A(new_n683_), .B(new_n679_), .Y(new_n744_));
  NAND2X1  g00488(.A(new_n599_), .B(new_n644_), .Y(new_n745_));
  OAI21X1  g00489(.A0(new_n607_), .A1(new_n600_), .B0(new_n745_), .Y(new_n746_));
  XOR2X1   g00490(.A(new_n678_), .B(new_n746_), .Y(new_n747_));
  XOR2X1   g00491(.A(new_n683_), .B(new_n747_), .Y(new_n748_));
  OAI21X1  g00492(.A0(new_n688_), .A1(new_n748_), .B0(new_n744_), .Y(new_n749_));
  NOR2X1   g00493(.A(new_n676_), .B(new_n666_), .Y(new_n750_));
  INVX1    g00494(.A(new_n668_), .Y(new_n751_));
  XOR2X1   g00495(.A(new_n665_), .B(\a[13] ), .Y(new_n752_));
  XOR2X1   g00496(.A(\a[13] ), .B(\a[12] ), .Y(new_n753_));
  NOR4X1   g00497(.A(new_n753_), .B(new_n752_), .C(new_n598_), .D(new_n274_), .Y(new_n754_));
  NOR3X1   g00498(.A(new_n667_), .B(new_n673_), .C(new_n277_), .Y(new_n755_));
  NOR3X1   g00499(.A(new_n671_), .B(new_n598_), .C(new_n275_), .Y(new_n756_));
  NOR3X1   g00500(.A(new_n756_), .B(new_n755_), .C(new_n754_), .Y(new_n757_));
  OAI21X1  g00501(.A0(new_n751_), .A1(new_n281_), .B0(new_n757_), .Y(new_n758_));
  XOR2X1   g00502(.A(new_n758_), .B(new_n665_), .Y(new_n759_));
  XOR2X1   g00503(.A(new_n759_), .B(new_n750_), .Y(new_n760_));
  AOI22X1  g00504(.A0(new_n603_), .A1(\b[5] ), .B0(new_n602_), .B1(\b[4] ), .Y(new_n761_));
  OAI21X1  g00505(.A0(new_n601_), .A1(new_n297_), .B0(new_n761_), .Y(new_n762_));
  AOI21X1  g00506(.A0(new_n518_), .A1(new_n349_), .B0(new_n762_), .Y(new_n763_));
  XOR2X1   g00507(.A(new_n763_), .B(\a[11] ), .Y(new_n764_));
  NAND2X1  g00508(.A(new_n764_), .B(new_n760_), .Y(new_n765_));
  AND2X1   g00509(.A(new_n677_), .B(new_n664_), .Y(new_n766_));
  AOI21X1  g00510(.A0(new_n678_), .A1(new_n746_), .B0(new_n766_), .Y(new_n767_));
  OR2X1    g00511(.A(new_n764_), .B(new_n760_), .Y(new_n768_));
  AOI21X1  g00512(.A0(new_n765_), .A1(new_n768_), .B0(new_n767_), .Y(new_n769_));
  NOR2X1   g00513(.A(new_n677_), .B(new_n664_), .Y(new_n770_));
  NAND2X1  g00514(.A(new_n677_), .B(new_n664_), .Y(new_n771_));
  OAI21X1  g00515(.A0(new_n770_), .A1(new_n657_), .B0(new_n771_), .Y(new_n772_));
  NOR2X1   g00516(.A(new_n764_), .B(new_n760_), .Y(new_n773_));
  AOI21X1  g00517(.A0(new_n765_), .A1(new_n772_), .B0(new_n773_), .Y(new_n774_));
  AOI21X1  g00518(.A0(new_n774_), .A1(new_n765_), .B0(new_n769_), .Y(new_n775_));
  AOI22X1  g00519(.A0(new_n469_), .A1(\b[8] ), .B0(new_n468_), .B1(\b[7] ), .Y(new_n776_));
  OAI21X1  g00520(.A0(new_n467_), .A1(new_n392_), .B0(new_n776_), .Y(new_n777_));
  AOI21X1  g00521(.A0(new_n454_), .A1(new_n404_), .B0(new_n777_), .Y(new_n778_));
  XOR2X1   g00522(.A(new_n778_), .B(\a[8] ), .Y(new_n779_));
  XOR2X1   g00523(.A(new_n779_), .B(new_n775_), .Y(new_n780_));
  XOR2X1   g00524(.A(new_n780_), .B(new_n749_), .Y(new_n781_));
  XOR2X1   g00525(.A(new_n781_), .B(new_n743_), .Y(new_n782_));
  XOR2X1   g00526(.A(new_n782_), .B(new_n739_), .Y(new_n783_));
  XOR2X1   g00527(.A(new_n783_), .B(new_n738_), .Y(new_n784_));
  XOR2X1   g00528(.A(new_n784_), .B(new_n730_), .Y(\f[14] ));
  AOI21X1  g00529(.A0(new_n729_), .A1(new_n728_), .B0(new_n784_), .Y(new_n786_));
  INVX1    g00530(.A(new_n738_), .Y(new_n787_));
  AND2X1   g00531(.A(new_n783_), .B(new_n787_), .Y(new_n788_));
  OR2X1    g00532(.A(new_n788_), .B(new_n786_), .Y(new_n789_));
  AND2X1   g00533(.A(\b[14] ), .B(\b[13] ), .Y(new_n790_));
  AOI21X1  g00534(.A0(new_n733_), .A1(new_n732_), .B0(new_n790_), .Y(new_n791_));
  INVX1    g00535(.A(\b[14] ), .Y(new_n792_));
  XOR2X1   g00536(.A(\b[15] ), .B(new_n792_), .Y(new_n793_));
  XOR2X1   g00537(.A(new_n793_), .B(new_n791_), .Y(new_n794_));
  INVX1    g00538(.A(\b[13] ), .Y(new_n795_));
  AOI22X1  g00539(.A0(new_n267_), .A1(\b[15] ), .B0(new_n266_), .B1(\b[14] ), .Y(new_n796_));
  OAI21X1  g00540(.A0(new_n350_), .A1(new_n795_), .B0(new_n796_), .Y(new_n797_));
  AOI21X1  g00541(.A0(new_n794_), .A1(new_n318_), .B0(new_n797_), .Y(new_n798_));
  XOR2X1   g00542(.A(new_n798_), .B(new_n257_), .Y(new_n799_));
  AND2X1   g00543(.A(new_n781_), .B(new_n743_), .Y(new_n800_));
  AOI21X1  g00544(.A0(new_n782_), .A1(new_n739_), .B0(new_n800_), .Y(new_n801_));
  AOI22X1  g00545(.A0(new_n369_), .A1(\b[12] ), .B0(new_n368_), .B1(\b[11] ), .Y(new_n802_));
  OAI21X1  g00546(.A0(new_n367_), .A1(new_n587_), .B0(new_n802_), .Y(new_n803_));
  AOI21X1  g00547(.A0(new_n635_), .A1(new_n308_), .B0(new_n803_), .Y(new_n804_));
  XOR2X1   g00548(.A(new_n804_), .B(\a[5] ), .Y(new_n805_));
  NOR2X1   g00549(.A(new_n779_), .B(new_n775_), .Y(new_n806_));
  AOI21X1  g00550(.A0(new_n780_), .A1(new_n749_), .B0(new_n806_), .Y(new_n807_));
  AOI22X1  g00551(.A0(new_n469_), .A1(\b[9] ), .B0(new_n468_), .B1(\b[8] ), .Y(new_n808_));
  OAI21X1  g00552(.A0(new_n467_), .A1(new_n492_), .B0(new_n808_), .Y(new_n809_));
  AOI21X1  g00553(.A0(new_n491_), .A1(new_n404_), .B0(new_n809_), .Y(new_n810_));
  XOR2X1   g00554(.A(new_n810_), .B(\a[8] ), .Y(new_n811_));
  OR4X1    g00555(.A(new_n758_), .B(new_n676_), .C(new_n599_), .D(new_n665_), .Y(new_n812_));
  XOR2X1   g00556(.A(\a[15] ), .B(\a[14] ), .Y(new_n813_));
  AND2X1   g00557(.A(new_n813_), .B(\b[0] ), .Y(new_n814_));
  XOR2X1   g00558(.A(new_n814_), .B(new_n812_), .Y(new_n815_));
  NAND3X1  g00559(.A(new_n671_), .B(new_n667_), .C(new_n673_), .Y(new_n816_));
  AND2X1   g00560(.A(new_n753_), .B(new_n673_), .Y(new_n817_));
  AND2X1   g00561(.A(new_n752_), .B(new_n598_), .Y(new_n818_));
  AOI22X1  g00562(.A0(new_n818_), .A1(\b[3] ), .B0(new_n817_), .B1(\b[2] ), .Y(new_n819_));
  OAI21X1  g00563(.A0(new_n816_), .A1(new_n275_), .B0(new_n819_), .Y(new_n820_));
  AOI21X1  g00564(.A0(new_n668_), .A1(new_n366_), .B0(new_n820_), .Y(new_n821_));
  XOR2X1   g00565(.A(new_n821_), .B(\a[14] ), .Y(new_n822_));
  XOR2X1   g00566(.A(new_n822_), .B(new_n815_), .Y(new_n823_));
  AOI22X1  g00567(.A0(new_n603_), .A1(\b[6] ), .B0(new_n602_), .B1(\b[5] ), .Y(new_n824_));
  OAI21X1  g00568(.A0(new_n601_), .A1(new_n325_), .B0(new_n824_), .Y(new_n825_));
  AOI21X1  g00569(.A0(new_n518_), .A1(new_n378_), .B0(new_n825_), .Y(new_n826_));
  XOR2X1   g00570(.A(new_n826_), .B(\a[11] ), .Y(new_n827_));
  XOR2X1   g00571(.A(new_n827_), .B(new_n823_), .Y(new_n828_));
  XOR2X1   g00572(.A(new_n828_), .B(new_n774_), .Y(new_n829_));
  XOR2X1   g00573(.A(new_n829_), .B(new_n811_), .Y(new_n830_));
  XOR2X1   g00574(.A(new_n830_), .B(new_n807_), .Y(new_n831_));
  XOR2X1   g00575(.A(new_n831_), .B(new_n805_), .Y(new_n832_));
  XOR2X1   g00576(.A(new_n832_), .B(new_n801_), .Y(new_n833_));
  XOR2X1   g00577(.A(new_n833_), .B(new_n799_), .Y(new_n834_));
  XOR2X1   g00578(.A(new_n834_), .B(new_n789_), .Y(\f[15] ));
  NAND2X1  g00579(.A(new_n833_), .B(new_n799_), .Y(new_n836_));
  OAI21X1  g00580(.A0(new_n788_), .A1(new_n786_), .B0(new_n834_), .Y(new_n837_));
  AND2X1   g00581(.A(new_n837_), .B(new_n836_), .Y(new_n838_));
  NAND2X1  g00582(.A(\b[15] ), .B(\b[14] ), .Y(new_n839_));
  OAI21X1  g00583(.A0(new_n793_), .A1(new_n791_), .B0(new_n839_), .Y(new_n840_));
  XOR2X1   g00584(.A(\b[16] ), .B(\b[15] ), .Y(new_n841_));
  XOR2X1   g00585(.A(new_n841_), .B(new_n840_), .Y(new_n842_));
  AOI22X1  g00586(.A0(new_n267_), .A1(\b[16] ), .B0(new_n266_), .B1(\b[15] ), .Y(new_n843_));
  OAI21X1  g00587(.A0(new_n350_), .A1(new_n792_), .B0(new_n843_), .Y(new_n844_));
  AOI21X1  g00588(.A0(new_n842_), .A1(new_n318_), .B0(new_n844_), .Y(new_n845_));
  XOR2X1   g00589(.A(new_n845_), .B(\a[2] ), .Y(new_n846_));
  INVX1    g00590(.A(new_n805_), .Y(new_n847_));
  NAND2X1  g00591(.A(new_n831_), .B(new_n847_), .Y(new_n848_));
  OAI21X1  g00592(.A0(new_n832_), .A1(new_n801_), .B0(new_n848_), .Y(new_n849_));
  AOI22X1  g00593(.A0(new_n369_), .A1(\b[13] ), .B0(new_n368_), .B1(\b[12] ), .Y(new_n850_));
  OAI21X1  g00594(.A0(new_n367_), .A1(new_n716_), .B0(new_n850_), .Y(new_n851_));
  AOI21X1  g00595(.A0(new_n715_), .A1(new_n308_), .B0(new_n851_), .Y(new_n852_));
  XOR2X1   g00596(.A(new_n852_), .B(new_n305_), .Y(new_n853_));
  INVX1    g00597(.A(new_n811_), .Y(new_n854_));
  NAND2X1  g00598(.A(new_n829_), .B(new_n854_), .Y(new_n855_));
  OAI21X1  g00599(.A0(new_n830_), .A1(new_n807_), .B0(new_n855_), .Y(new_n856_));
  AOI22X1  g00600(.A0(new_n469_), .A1(\b[10] ), .B0(new_n468_), .B1(\b[9] ), .Y(new_n857_));
  OAI21X1  g00601(.A0(new_n467_), .A1(new_n489_), .B0(new_n857_), .Y(new_n858_));
  AOI21X1  g00602(.A0(new_n543_), .A1(new_n404_), .B0(new_n858_), .Y(new_n859_));
  XOR2X1   g00603(.A(new_n859_), .B(new_n400_), .Y(new_n860_));
  NOR4X1   g00604(.A(new_n758_), .B(new_n676_), .C(new_n599_), .D(new_n665_), .Y(new_n861_));
  XOR2X1   g00605(.A(new_n814_), .B(new_n861_), .Y(new_n862_));
  XOR2X1   g00606(.A(new_n822_), .B(new_n862_), .Y(new_n863_));
  OR2X1    g00607(.A(new_n827_), .B(new_n863_), .Y(new_n864_));
  OAI21X1  g00608(.A0(new_n828_), .A1(new_n774_), .B0(new_n864_), .Y(new_n865_));
  AOI22X1  g00609(.A0(new_n603_), .A1(\b[7] ), .B0(new_n602_), .B1(\b[6] ), .Y(new_n866_));
  OAI21X1  g00610(.A0(new_n601_), .A1(new_n395_), .B0(new_n866_), .Y(new_n867_));
  AOI21X1  g00611(.A0(new_n518_), .A1(new_n394_), .B0(new_n867_), .Y(new_n868_));
  XOR2X1   g00612(.A(new_n868_), .B(new_n515_), .Y(new_n869_));
  NAND2X1  g00613(.A(new_n814_), .B(new_n861_), .Y(new_n870_));
  OAI21X1  g00614(.A0(new_n822_), .A1(new_n815_), .B0(new_n870_), .Y(new_n871_));
  AND2X1   g00615(.A(new_n668_), .B(new_n323_), .Y(new_n872_));
  NOR4X1   g00616(.A(new_n753_), .B(new_n752_), .C(new_n598_), .D(new_n277_), .Y(new_n873_));
  NAND2X1  g00617(.A(new_n753_), .B(new_n673_), .Y(new_n874_));
  NAND2X1  g00618(.A(new_n752_), .B(new_n598_), .Y(new_n875_));
  OAI22X1  g00619(.A0(new_n875_), .A1(new_n325_), .B0(new_n874_), .B1(new_n297_), .Y(new_n876_));
  NOR3X1   g00620(.A(new_n876_), .B(new_n873_), .C(new_n872_), .Y(new_n877_));
  XOR2X1   g00621(.A(new_n877_), .B(new_n665_), .Y(new_n878_));
  INVX1    g00622(.A(\a[17] ), .Y(new_n879_));
  OR2X1    g00623(.A(new_n814_), .B(new_n879_), .Y(new_n880_));
  XOR2X1   g00624(.A(\a[17] ), .B(\a[16] ), .Y(new_n881_));
  AND2X1   g00625(.A(new_n881_), .B(new_n813_), .Y(new_n882_));
  AND2X1   g00626(.A(new_n882_), .B(new_n263_), .Y(new_n883_));
  INVX1    g00627(.A(\a[15] ), .Y(new_n884_));
  XOR2X1   g00628(.A(\a[16] ), .B(new_n884_), .Y(new_n885_));
  NOR3X1   g00629(.A(new_n885_), .B(new_n813_), .C(new_n274_), .Y(new_n886_));
  XOR2X1   g00630(.A(\a[15] ), .B(new_n665_), .Y(new_n887_));
  NOR3X1   g00631(.A(new_n881_), .B(new_n887_), .C(new_n275_), .Y(new_n888_));
  NOR3X1   g00632(.A(new_n888_), .B(new_n886_), .C(new_n883_), .Y(new_n889_));
  XOR2X1   g00633(.A(new_n889_), .B(\a[17] ), .Y(new_n890_));
  XOR2X1   g00634(.A(new_n890_), .B(new_n880_), .Y(new_n891_));
  XOR2X1   g00635(.A(new_n891_), .B(new_n878_), .Y(new_n892_));
  XOR2X1   g00636(.A(new_n892_), .B(new_n871_), .Y(new_n893_));
  XOR2X1   g00637(.A(new_n893_), .B(new_n869_), .Y(new_n894_));
  XOR2X1   g00638(.A(new_n894_), .B(new_n865_), .Y(new_n895_));
  XOR2X1   g00639(.A(new_n895_), .B(new_n860_), .Y(new_n896_));
  XOR2X1   g00640(.A(new_n896_), .B(new_n856_), .Y(new_n897_));
  XOR2X1   g00641(.A(new_n897_), .B(new_n853_), .Y(new_n898_));
  XOR2X1   g00642(.A(new_n898_), .B(new_n849_), .Y(new_n899_));
  XOR2X1   g00643(.A(new_n899_), .B(new_n846_), .Y(new_n900_));
  XOR2X1   g00644(.A(new_n900_), .B(new_n838_), .Y(\f[16] ));
  AND2X1   g00645(.A(new_n897_), .B(new_n853_), .Y(new_n902_));
  AOI21X1  g00646(.A0(new_n898_), .A1(new_n849_), .B0(new_n902_), .Y(new_n903_));
  AOI22X1  g00647(.A0(new_n369_), .A1(\b[14] ), .B0(new_n368_), .B1(\b[13] ), .Y(new_n904_));
  OAI21X1  g00648(.A0(new_n367_), .A1(new_n713_), .B0(new_n904_), .Y(new_n905_));
  AOI21X1  g00649(.A0(new_n734_), .A1(new_n308_), .B0(new_n905_), .Y(new_n906_));
  XOR2X1   g00650(.A(new_n906_), .B(new_n305_), .Y(new_n907_));
  NOR2X1   g00651(.A(new_n683_), .B(new_n679_), .Y(new_n908_));
  OR2X1    g00652(.A(new_n612_), .B(new_n646_), .Y(new_n909_));
  OAI21X1  g00653(.A0(new_n620_), .A1(new_n613_), .B0(new_n909_), .Y(new_n910_));
  AOI21X1  g00654(.A0(new_n910_), .A1(new_n684_), .B0(new_n908_), .Y(new_n911_));
  AND2X1   g00655(.A(new_n779_), .B(new_n775_), .Y(new_n912_));
  OR2X1    g00656(.A(new_n779_), .B(new_n775_), .Y(new_n913_));
  OAI21X1  g00657(.A0(new_n912_), .A1(new_n911_), .B0(new_n913_), .Y(new_n914_));
  AND2X1   g00658(.A(new_n829_), .B(new_n854_), .Y(new_n915_));
  XOR2X1   g00659(.A(new_n829_), .B(new_n854_), .Y(new_n916_));
  AOI21X1  g00660(.A0(new_n916_), .A1(new_n914_), .B0(new_n915_), .Y(new_n917_));
  NOR2X1   g00661(.A(new_n895_), .B(new_n860_), .Y(new_n918_));
  NAND2X1  g00662(.A(new_n895_), .B(new_n860_), .Y(new_n919_));
  OAI21X1  g00663(.A0(new_n918_), .A1(new_n917_), .B0(new_n919_), .Y(new_n920_));
  AOI22X1  g00664(.A0(new_n469_), .A1(\b[11] ), .B0(new_n468_), .B1(\b[10] ), .Y(new_n921_));
  OAI21X1  g00665(.A0(new_n467_), .A1(new_n590_), .B0(new_n921_), .Y(new_n922_));
  AOI21X1  g00666(.A0(new_n589_), .A1(new_n404_), .B0(new_n922_), .Y(new_n923_));
  XOR2X1   g00667(.A(new_n923_), .B(new_n400_), .Y(new_n924_));
  AND2X1   g00668(.A(new_n764_), .B(new_n760_), .Y(new_n925_));
  OAI21X1  g00669(.A0(new_n925_), .A1(new_n767_), .B0(new_n768_), .Y(new_n926_));
  NOR2X1   g00670(.A(new_n827_), .B(new_n863_), .Y(new_n927_));
  XOR2X1   g00671(.A(new_n827_), .B(new_n863_), .Y(new_n928_));
  AOI21X1  g00672(.A0(new_n928_), .A1(new_n926_), .B0(new_n927_), .Y(new_n929_));
  NOR2X1   g00673(.A(new_n893_), .B(new_n869_), .Y(new_n930_));
  NAND2X1  g00674(.A(new_n893_), .B(new_n869_), .Y(new_n931_));
  OAI21X1  g00675(.A0(new_n930_), .A1(new_n929_), .B0(new_n931_), .Y(new_n932_));
  NOR2X1   g00676(.A(new_n890_), .B(new_n880_), .Y(new_n933_));
  INVX1    g00677(.A(new_n882_), .Y(new_n934_));
  XOR2X1   g00678(.A(new_n879_), .B(\a[16] ), .Y(new_n935_));
  XOR2X1   g00679(.A(\a[16] ), .B(\a[15] ), .Y(new_n936_));
  NOR4X1   g00680(.A(new_n936_), .B(new_n935_), .C(new_n813_), .D(new_n274_), .Y(new_n937_));
  NOR3X1   g00681(.A(new_n881_), .B(new_n887_), .C(new_n277_), .Y(new_n938_));
  NOR3X1   g00682(.A(new_n885_), .B(new_n813_), .C(new_n275_), .Y(new_n939_));
  NOR3X1   g00683(.A(new_n939_), .B(new_n938_), .C(new_n937_), .Y(new_n940_));
  OAI21X1  g00684(.A0(new_n934_), .A1(new_n281_), .B0(new_n940_), .Y(new_n941_));
  XOR2X1   g00685(.A(new_n941_), .B(new_n879_), .Y(new_n942_));
  XOR2X1   g00686(.A(new_n942_), .B(new_n933_), .Y(new_n943_));
  AOI22X1  g00687(.A0(new_n818_), .A1(\b[5] ), .B0(new_n817_), .B1(\b[4] ), .Y(new_n944_));
  OAI21X1  g00688(.A0(new_n816_), .A1(new_n297_), .B0(new_n944_), .Y(new_n945_));
  AOI21X1  g00689(.A0(new_n668_), .A1(new_n349_), .B0(new_n945_), .Y(new_n946_));
  XOR2X1   g00690(.A(new_n946_), .B(\a[14] ), .Y(new_n947_));
  NAND2X1  g00691(.A(new_n947_), .B(new_n943_), .Y(new_n948_));
  AND2X1   g00692(.A(new_n891_), .B(new_n878_), .Y(new_n949_));
  AOI21X1  g00693(.A0(new_n892_), .A1(new_n871_), .B0(new_n949_), .Y(new_n950_));
  OR2X1    g00694(.A(new_n947_), .B(new_n943_), .Y(new_n951_));
  AOI21X1  g00695(.A0(new_n948_), .A1(new_n951_), .B0(new_n950_), .Y(new_n952_));
  XOR2X1   g00696(.A(new_n821_), .B(new_n665_), .Y(new_n953_));
  AND2X1   g00697(.A(new_n814_), .B(new_n861_), .Y(new_n954_));
  AOI21X1  g00698(.A0(new_n953_), .A1(new_n862_), .B0(new_n954_), .Y(new_n955_));
  NOR2X1   g00699(.A(new_n891_), .B(new_n878_), .Y(new_n956_));
  NAND2X1  g00700(.A(new_n891_), .B(new_n878_), .Y(new_n957_));
  OAI21X1  g00701(.A0(new_n956_), .A1(new_n955_), .B0(new_n957_), .Y(new_n958_));
  NOR2X1   g00702(.A(new_n947_), .B(new_n943_), .Y(new_n959_));
  AOI21X1  g00703(.A0(new_n948_), .A1(new_n958_), .B0(new_n959_), .Y(new_n960_));
  AOI21X1  g00704(.A0(new_n960_), .A1(new_n948_), .B0(new_n952_), .Y(new_n961_));
  AOI22X1  g00705(.A0(new_n603_), .A1(\b[8] ), .B0(new_n602_), .B1(\b[7] ), .Y(new_n962_));
  OAI21X1  g00706(.A0(new_n601_), .A1(new_n392_), .B0(new_n962_), .Y(new_n963_));
  AOI21X1  g00707(.A0(new_n518_), .A1(new_n454_), .B0(new_n963_), .Y(new_n964_));
  XOR2X1   g00708(.A(new_n964_), .B(\a[11] ), .Y(new_n965_));
  XOR2X1   g00709(.A(new_n965_), .B(new_n961_), .Y(new_n966_));
  XOR2X1   g00710(.A(new_n966_), .B(new_n932_), .Y(new_n967_));
  XOR2X1   g00711(.A(new_n967_), .B(new_n924_), .Y(new_n968_));
  XOR2X1   g00712(.A(new_n968_), .B(new_n920_), .Y(new_n969_));
  XOR2X1   g00713(.A(new_n969_), .B(new_n907_), .Y(new_n970_));
  XOR2X1   g00714(.A(new_n970_), .B(new_n903_), .Y(new_n971_));
  AND2X1   g00715(.A(\b[16] ), .B(\b[15] ), .Y(new_n972_));
  AOI21X1  g00716(.A0(new_n841_), .A1(new_n840_), .B0(new_n972_), .Y(new_n973_));
  INVX1    g00717(.A(\b[16] ), .Y(new_n974_));
  XOR2X1   g00718(.A(\b[17] ), .B(new_n974_), .Y(new_n975_));
  XOR2X1   g00719(.A(new_n975_), .B(new_n973_), .Y(new_n976_));
  INVX1    g00720(.A(\b[15] ), .Y(new_n977_));
  AOI22X1  g00721(.A0(new_n267_), .A1(\b[17] ), .B0(new_n266_), .B1(\b[16] ), .Y(new_n978_));
  OAI21X1  g00722(.A0(new_n350_), .A1(new_n977_), .B0(new_n978_), .Y(new_n979_));
  AOI21X1  g00723(.A0(new_n976_), .A1(new_n318_), .B0(new_n979_), .Y(new_n980_));
  XOR2X1   g00724(.A(new_n980_), .B(\a[2] ), .Y(new_n981_));
  XOR2X1   g00725(.A(new_n981_), .B(new_n971_), .Y(new_n982_));
  AOI21X1  g00726(.A0(new_n837_), .A1(new_n836_), .B0(new_n900_), .Y(new_n983_));
  INVX1    g00727(.A(new_n846_), .Y(new_n984_));
  AND2X1   g00728(.A(new_n899_), .B(new_n984_), .Y(new_n985_));
  OR2X1    g00729(.A(new_n985_), .B(new_n983_), .Y(new_n986_));
  XOR2X1   g00730(.A(new_n986_), .B(new_n982_), .Y(\f[17] ));
  NOR2X1   g00731(.A(new_n969_), .B(new_n907_), .Y(new_n988_));
  NAND2X1  g00732(.A(new_n969_), .B(new_n907_), .Y(new_n989_));
  OAI21X1  g00733(.A0(new_n988_), .A1(new_n903_), .B0(new_n989_), .Y(new_n990_));
  AOI22X1  g00734(.A0(new_n369_), .A1(\b[15] ), .B0(new_n368_), .B1(\b[14] ), .Y(new_n991_));
  OAI21X1  g00735(.A0(new_n367_), .A1(new_n795_), .B0(new_n991_), .Y(new_n992_));
  AOI21X1  g00736(.A0(new_n794_), .A1(new_n308_), .B0(new_n992_), .Y(new_n993_));
  XOR2X1   g00737(.A(new_n993_), .B(new_n305_), .Y(new_n994_));
  AND2X1   g00738(.A(new_n895_), .B(new_n860_), .Y(new_n995_));
  AOI21X1  g00739(.A0(new_n896_), .A1(new_n856_), .B0(new_n995_), .Y(new_n996_));
  NOR2X1   g00740(.A(new_n967_), .B(new_n924_), .Y(new_n997_));
  NAND2X1  g00741(.A(new_n967_), .B(new_n924_), .Y(new_n998_));
  OAI21X1  g00742(.A0(new_n997_), .A1(new_n996_), .B0(new_n998_), .Y(new_n999_));
  AOI22X1  g00743(.A0(new_n469_), .A1(\b[12] ), .B0(new_n468_), .B1(\b[11] ), .Y(new_n1000_));
  OAI21X1  g00744(.A0(new_n467_), .A1(new_n587_), .B0(new_n1000_), .Y(new_n1001_));
  AOI21X1  g00745(.A0(new_n635_), .A1(new_n404_), .B0(new_n1001_), .Y(new_n1002_));
  XOR2X1   g00746(.A(new_n1002_), .B(new_n400_), .Y(new_n1003_));
  AND2X1   g00747(.A(new_n893_), .B(new_n869_), .Y(new_n1004_));
  AOI21X1  g00748(.A0(new_n894_), .A1(new_n865_), .B0(new_n1004_), .Y(new_n1005_));
  AND2X1   g00749(.A(new_n965_), .B(new_n961_), .Y(new_n1006_));
  OR2X1    g00750(.A(new_n965_), .B(new_n961_), .Y(new_n1007_));
  OAI21X1  g00751(.A0(new_n1006_), .A1(new_n1005_), .B0(new_n1007_), .Y(new_n1008_));
  AND2X1   g00752(.A(new_n947_), .B(new_n943_), .Y(new_n1009_));
  OAI21X1  g00753(.A0(new_n1009_), .A1(new_n950_), .B0(new_n951_), .Y(new_n1010_));
  OR4X1    g00754(.A(new_n941_), .B(new_n890_), .C(new_n814_), .D(new_n879_), .Y(new_n1011_));
  XOR2X1   g00755(.A(\a[18] ), .B(\a[17] ), .Y(new_n1012_));
  AND2X1   g00756(.A(new_n1012_), .B(\b[0] ), .Y(new_n1013_));
  XOR2X1   g00757(.A(new_n1013_), .B(new_n1011_), .Y(new_n1014_));
  NAND3X1  g00758(.A(new_n885_), .B(new_n881_), .C(new_n887_), .Y(new_n1015_));
  AND2X1   g00759(.A(new_n936_), .B(new_n887_), .Y(new_n1016_));
  AND2X1   g00760(.A(new_n935_), .B(new_n813_), .Y(new_n1017_));
  AOI22X1  g00761(.A0(new_n1017_), .A1(\b[3] ), .B0(new_n1016_), .B1(\b[2] ), .Y(new_n1018_));
  OAI21X1  g00762(.A0(new_n1015_), .A1(new_n275_), .B0(new_n1018_), .Y(new_n1019_));
  AOI21X1  g00763(.A0(new_n882_), .A1(new_n366_), .B0(new_n1019_), .Y(new_n1020_));
  XOR2X1   g00764(.A(new_n1020_), .B(\a[17] ), .Y(new_n1021_));
  XOR2X1   g00765(.A(new_n1021_), .B(new_n1014_), .Y(new_n1022_));
  AOI22X1  g00766(.A0(new_n818_), .A1(\b[6] ), .B0(new_n817_), .B1(\b[5] ), .Y(new_n1023_));
  OAI21X1  g00767(.A0(new_n816_), .A1(new_n325_), .B0(new_n1023_), .Y(new_n1024_));
  AOI21X1  g00768(.A0(new_n668_), .A1(new_n378_), .B0(new_n1024_), .Y(new_n1025_));
  XOR2X1   g00769(.A(new_n1025_), .B(\a[14] ), .Y(new_n1026_));
  XOR2X1   g00770(.A(new_n1026_), .B(new_n1022_), .Y(new_n1027_));
  XOR2X1   g00771(.A(new_n1027_), .B(new_n1010_), .Y(new_n1028_));
  AOI22X1  g00772(.A0(new_n603_), .A1(\b[9] ), .B0(new_n602_), .B1(\b[8] ), .Y(new_n1029_));
  OAI21X1  g00773(.A0(new_n601_), .A1(new_n492_), .B0(new_n1029_), .Y(new_n1030_));
  AOI21X1  g00774(.A0(new_n518_), .A1(new_n491_), .B0(new_n1030_), .Y(new_n1031_));
  XOR2X1   g00775(.A(new_n1031_), .B(\a[11] ), .Y(new_n1032_));
  XOR2X1   g00776(.A(new_n1032_), .B(new_n1028_), .Y(new_n1033_));
  XOR2X1   g00777(.A(new_n1033_), .B(new_n1008_), .Y(new_n1034_));
  XOR2X1   g00778(.A(new_n1034_), .B(new_n1003_), .Y(new_n1035_));
  XOR2X1   g00779(.A(new_n1035_), .B(new_n999_), .Y(new_n1036_));
  XOR2X1   g00780(.A(new_n1036_), .B(new_n994_), .Y(new_n1037_));
  XOR2X1   g00781(.A(new_n1037_), .B(new_n990_), .Y(new_n1038_));
  NAND2X1  g00782(.A(\b[17] ), .B(\b[16] ), .Y(new_n1039_));
  OAI21X1  g00783(.A0(new_n975_), .A1(new_n973_), .B0(new_n1039_), .Y(new_n1040_));
  XOR2X1   g00784(.A(\b[18] ), .B(\b[17] ), .Y(new_n1041_));
  XOR2X1   g00785(.A(new_n1041_), .B(new_n1040_), .Y(new_n1042_));
  AOI22X1  g00786(.A0(new_n267_), .A1(\b[18] ), .B0(new_n266_), .B1(\b[17] ), .Y(new_n1043_));
  OAI21X1  g00787(.A0(new_n350_), .A1(new_n974_), .B0(new_n1043_), .Y(new_n1044_));
  AOI21X1  g00788(.A0(new_n1042_), .A1(new_n318_), .B0(new_n1044_), .Y(new_n1045_));
  XOR2X1   g00789(.A(new_n1045_), .B(\a[2] ), .Y(new_n1046_));
  XOR2X1   g00790(.A(new_n1046_), .B(new_n1038_), .Y(new_n1047_));
  OR2X1    g00791(.A(new_n981_), .B(new_n971_), .Y(new_n1048_));
  OAI21X1  g00792(.A0(new_n985_), .A1(new_n983_), .B0(new_n982_), .Y(new_n1049_));
  AND2X1   g00793(.A(new_n1049_), .B(new_n1048_), .Y(new_n1050_));
  XOR2X1   g00794(.A(new_n1050_), .B(new_n1047_), .Y(\f[18] ));
  NOR4X1   g00795(.A(new_n941_), .B(new_n890_), .C(new_n814_), .D(new_n879_), .Y(new_n1052_));
  XOR2X1   g00796(.A(new_n1013_), .B(new_n1052_), .Y(new_n1053_));
  XOR2X1   g00797(.A(new_n1021_), .B(new_n1053_), .Y(new_n1054_));
  NOR2X1   g00798(.A(new_n1026_), .B(new_n1054_), .Y(new_n1055_));
  XOR2X1   g00799(.A(new_n1026_), .B(new_n1054_), .Y(new_n1056_));
  AOI21X1  g00800(.A0(new_n1056_), .A1(new_n1010_), .B0(new_n1055_), .Y(new_n1057_));
  AOI22X1  g00801(.A0(new_n818_), .A1(\b[7] ), .B0(new_n817_), .B1(\b[6] ), .Y(new_n1058_));
  OAI21X1  g00802(.A0(new_n816_), .A1(new_n395_), .B0(new_n1058_), .Y(new_n1059_));
  AOI21X1  g00803(.A0(new_n668_), .A1(new_n394_), .B0(new_n1059_), .Y(new_n1060_));
  XOR2X1   g00804(.A(new_n1060_), .B(new_n665_), .Y(new_n1061_));
  XOR2X1   g00805(.A(new_n1020_), .B(new_n879_), .Y(new_n1062_));
  AND2X1   g00806(.A(new_n1013_), .B(new_n1052_), .Y(new_n1063_));
  AOI21X1  g00807(.A0(new_n1062_), .A1(new_n1053_), .B0(new_n1063_), .Y(new_n1064_));
  AND2X1   g00808(.A(new_n882_), .B(new_n323_), .Y(new_n1065_));
  NOR4X1   g00809(.A(new_n936_), .B(new_n935_), .C(new_n813_), .D(new_n277_), .Y(new_n1066_));
  NAND2X1  g00810(.A(new_n936_), .B(new_n887_), .Y(new_n1067_));
  NAND2X1  g00811(.A(new_n935_), .B(new_n813_), .Y(new_n1068_));
  OAI22X1  g00812(.A0(new_n1068_), .A1(new_n325_), .B0(new_n1067_), .B1(new_n297_), .Y(new_n1069_));
  NOR3X1   g00813(.A(new_n1069_), .B(new_n1066_), .C(new_n1065_), .Y(new_n1070_));
  XOR2X1   g00814(.A(new_n1070_), .B(\a[17] ), .Y(new_n1071_));
  INVX1    g00815(.A(\a[20] ), .Y(new_n1072_));
  OR2X1    g00816(.A(new_n1013_), .B(new_n1072_), .Y(new_n1073_));
  XOR2X1   g00817(.A(\a[20] ), .B(\a[19] ), .Y(new_n1074_));
  AND2X1   g00818(.A(new_n1074_), .B(new_n1012_), .Y(new_n1075_));
  XOR2X1   g00819(.A(\a[18] ), .B(new_n879_), .Y(new_n1076_));
  XOR2X1   g00820(.A(\a[19] ), .B(\a[18] ), .Y(new_n1077_));
  NAND2X1  g00821(.A(new_n1077_), .B(new_n1076_), .Y(new_n1078_));
  XOR2X1   g00822(.A(new_n1072_), .B(\a[19] ), .Y(new_n1079_));
  NAND2X1  g00823(.A(new_n1079_), .B(new_n1012_), .Y(new_n1080_));
  OAI22X1  g00824(.A0(new_n1080_), .A1(new_n275_), .B0(new_n1078_), .B1(new_n274_), .Y(new_n1081_));
  AOI21X1  g00825(.A0(new_n1075_), .A1(new_n263_), .B0(new_n1081_), .Y(new_n1082_));
  XOR2X1   g00826(.A(new_n1082_), .B(\a[20] ), .Y(new_n1083_));
  XOR2X1   g00827(.A(new_n1083_), .B(new_n1073_), .Y(new_n1084_));
  XOR2X1   g00828(.A(new_n1084_), .B(new_n1071_), .Y(new_n1085_));
  XOR2X1   g00829(.A(new_n1085_), .B(new_n1064_), .Y(new_n1086_));
  XOR2X1   g00830(.A(new_n1086_), .B(new_n1061_), .Y(new_n1087_));
  XOR2X1   g00831(.A(new_n1087_), .B(new_n1057_), .Y(new_n1088_));
  AOI22X1  g00832(.A0(new_n603_), .A1(\b[10] ), .B0(new_n602_), .B1(\b[9] ), .Y(new_n1089_));
  OAI21X1  g00833(.A0(new_n601_), .A1(new_n489_), .B0(new_n1089_), .Y(new_n1090_));
  AOI21X1  g00834(.A0(new_n543_), .A1(new_n518_), .B0(new_n1090_), .Y(new_n1091_));
  XOR2X1   g00835(.A(new_n1091_), .B(\a[11] ), .Y(new_n1092_));
  XOR2X1   g00836(.A(new_n1092_), .B(new_n1088_), .Y(new_n1093_));
  NOR2X1   g00837(.A(new_n1032_), .B(new_n1028_), .Y(new_n1094_));
  AOI21X1  g00838(.A0(new_n1033_), .A1(new_n1008_), .B0(new_n1094_), .Y(new_n1095_));
  XOR2X1   g00839(.A(new_n1095_), .B(new_n1093_), .Y(new_n1096_));
  AOI22X1  g00840(.A0(new_n469_), .A1(\b[13] ), .B0(new_n468_), .B1(\b[12] ), .Y(new_n1097_));
  OAI21X1  g00841(.A0(new_n467_), .A1(new_n716_), .B0(new_n1097_), .Y(new_n1098_));
  AOI21X1  g00842(.A0(new_n715_), .A1(new_n404_), .B0(new_n1098_), .Y(new_n1099_));
  XOR2X1   g00843(.A(new_n1099_), .B(\a[8] ), .Y(new_n1100_));
  XOR2X1   g00844(.A(new_n1100_), .B(new_n1096_), .Y(new_n1101_));
  AND2X1   g00845(.A(new_n1034_), .B(new_n1003_), .Y(new_n1102_));
  AOI21X1  g00846(.A0(new_n1035_), .A1(new_n999_), .B0(new_n1102_), .Y(new_n1103_));
  XOR2X1   g00847(.A(new_n1103_), .B(new_n1101_), .Y(new_n1104_));
  AOI22X1  g00848(.A0(new_n369_), .A1(\b[16] ), .B0(new_n368_), .B1(\b[15] ), .Y(new_n1105_));
  OAI21X1  g00849(.A0(new_n367_), .A1(new_n792_), .B0(new_n1105_), .Y(new_n1106_));
  AOI21X1  g00850(.A0(new_n842_), .A1(new_n308_), .B0(new_n1106_), .Y(new_n1107_));
  XOR2X1   g00851(.A(new_n1107_), .B(\a[5] ), .Y(new_n1108_));
  XOR2X1   g00852(.A(new_n1108_), .B(new_n1104_), .Y(new_n1109_));
  AND2X1   g00853(.A(new_n1036_), .B(new_n994_), .Y(new_n1110_));
  AOI21X1  g00854(.A0(new_n1037_), .A1(new_n990_), .B0(new_n1110_), .Y(new_n1111_));
  XOR2X1   g00855(.A(new_n1111_), .B(new_n1109_), .Y(new_n1112_));
  AND2X1   g00856(.A(\b[18] ), .B(\b[17] ), .Y(new_n1113_));
  AOI21X1  g00857(.A0(new_n1041_), .A1(new_n1040_), .B0(new_n1113_), .Y(new_n1114_));
  INVX1    g00858(.A(\b[18] ), .Y(new_n1115_));
  XOR2X1   g00859(.A(\b[19] ), .B(new_n1115_), .Y(new_n1116_));
  XOR2X1   g00860(.A(new_n1116_), .B(new_n1114_), .Y(new_n1117_));
  INVX1    g00861(.A(\b[17] ), .Y(new_n1118_));
  AOI22X1  g00862(.A0(new_n267_), .A1(\b[19] ), .B0(new_n266_), .B1(\b[18] ), .Y(new_n1119_));
  OAI21X1  g00863(.A0(new_n350_), .A1(new_n1118_), .B0(new_n1119_), .Y(new_n1120_));
  AOI21X1  g00864(.A0(new_n1117_), .A1(new_n318_), .B0(new_n1120_), .Y(new_n1121_));
  XOR2X1   g00865(.A(new_n1121_), .B(\a[2] ), .Y(new_n1122_));
  XOR2X1   g00866(.A(new_n1122_), .B(new_n1112_), .Y(new_n1123_));
  AOI21X1  g00867(.A0(new_n709_), .A1(new_n654_), .B0(new_n694_), .Y(new_n1124_));
  NOR2X1   g00868(.A(new_n781_), .B(new_n743_), .Y(new_n1125_));
  NAND2X1  g00869(.A(new_n781_), .B(new_n743_), .Y(new_n1126_));
  OAI21X1  g00870(.A0(new_n1125_), .A1(new_n1124_), .B0(new_n1126_), .Y(new_n1127_));
  AND2X1   g00871(.A(new_n831_), .B(new_n847_), .Y(new_n1128_));
  XOR2X1   g00872(.A(new_n831_), .B(new_n847_), .Y(new_n1129_));
  AOI21X1  g00873(.A0(new_n1129_), .A1(new_n1127_), .B0(new_n1128_), .Y(new_n1130_));
  NOR2X1   g00874(.A(new_n897_), .B(new_n853_), .Y(new_n1131_));
  NAND2X1  g00875(.A(new_n897_), .B(new_n853_), .Y(new_n1132_));
  OAI21X1  g00876(.A0(new_n1131_), .A1(new_n1130_), .B0(new_n1132_), .Y(new_n1133_));
  AND2X1   g00877(.A(new_n969_), .B(new_n907_), .Y(new_n1134_));
  AOI21X1  g00878(.A0(new_n970_), .A1(new_n1133_), .B0(new_n1134_), .Y(new_n1135_));
  XOR2X1   g00879(.A(new_n1037_), .B(new_n1135_), .Y(new_n1136_));
  NOR2X1   g00880(.A(new_n1046_), .B(new_n1136_), .Y(new_n1137_));
  AOI21X1  g00881(.A0(new_n1049_), .A1(new_n1048_), .B0(new_n1047_), .Y(new_n1138_));
  OR2X1    g00882(.A(new_n1138_), .B(new_n1137_), .Y(new_n1139_));
  XOR2X1   g00883(.A(new_n1139_), .B(new_n1123_), .Y(\f[19] ));
  OR2X1    g00884(.A(new_n1108_), .B(new_n1104_), .Y(new_n1141_));
  OR2X1    g00885(.A(new_n1026_), .B(new_n1054_), .Y(new_n1142_));
  OAI21X1  g00886(.A0(new_n1027_), .A1(new_n960_), .B0(new_n1142_), .Y(new_n1143_));
  XOR2X1   g00887(.A(new_n1087_), .B(new_n1143_), .Y(new_n1144_));
  XOR2X1   g00888(.A(new_n1092_), .B(new_n1144_), .Y(new_n1145_));
  XOR2X1   g00889(.A(new_n1095_), .B(new_n1145_), .Y(new_n1146_));
  XOR2X1   g00890(.A(new_n1100_), .B(new_n1146_), .Y(new_n1147_));
  XOR2X1   g00891(.A(new_n1103_), .B(new_n1147_), .Y(new_n1148_));
  XOR2X1   g00892(.A(new_n1108_), .B(new_n1148_), .Y(new_n1149_));
  OAI21X1  g00893(.A0(new_n1111_), .A1(new_n1149_), .B0(new_n1141_), .Y(new_n1150_));
  AOI22X1  g00894(.A0(new_n369_), .A1(\b[17] ), .B0(new_n368_), .B1(\b[16] ), .Y(new_n1151_));
  OAI21X1  g00895(.A0(new_n367_), .A1(new_n977_), .B0(new_n1151_), .Y(new_n1152_));
  AOI21X1  g00896(.A0(new_n976_), .A1(new_n308_), .B0(new_n1152_), .Y(new_n1153_));
  XOR2X1   g00897(.A(new_n1153_), .B(\a[5] ), .Y(new_n1154_));
  OR2X1    g00898(.A(new_n1092_), .B(new_n1088_), .Y(new_n1155_));
  OAI21X1  g00899(.A0(new_n1095_), .A1(new_n1145_), .B0(new_n1155_), .Y(new_n1156_));
  AOI22X1  g00900(.A0(new_n603_), .A1(\b[11] ), .B0(new_n602_), .B1(\b[10] ), .Y(new_n1157_));
  OAI21X1  g00901(.A0(new_n601_), .A1(new_n590_), .B0(new_n1157_), .Y(new_n1158_));
  AOI21X1  g00902(.A0(new_n589_), .A1(new_n518_), .B0(new_n1158_), .Y(new_n1159_));
  XOR2X1   g00903(.A(new_n1159_), .B(new_n515_), .Y(new_n1160_));
  NAND2X1  g00904(.A(new_n1086_), .B(new_n1061_), .Y(new_n1161_));
  NOR2X1   g00905(.A(new_n1086_), .B(new_n1061_), .Y(new_n1162_));
  OAI21X1  g00906(.A0(new_n1162_), .A1(new_n1057_), .B0(new_n1161_), .Y(new_n1163_));
  NOR2X1   g00907(.A(new_n1083_), .B(new_n1073_), .Y(new_n1164_));
  INVX1    g00908(.A(new_n1075_), .Y(new_n1165_));
  OR2X1    g00909(.A(new_n1077_), .B(new_n1012_), .Y(new_n1166_));
  NOR2X1   g00910(.A(new_n1166_), .B(new_n1079_), .Y(new_n1167_));
  OAI22X1  g00911(.A0(new_n1080_), .A1(new_n277_), .B0(new_n1078_), .B1(new_n275_), .Y(new_n1168_));
  AOI21X1  g00912(.A0(new_n1167_), .A1(\b[0] ), .B0(new_n1168_), .Y(new_n1169_));
  OAI21X1  g00913(.A0(new_n1165_), .A1(new_n281_), .B0(new_n1169_), .Y(new_n1170_));
  XOR2X1   g00914(.A(new_n1170_), .B(new_n1072_), .Y(new_n1171_));
  XOR2X1   g00915(.A(new_n1171_), .B(new_n1164_), .Y(new_n1172_));
  AOI22X1  g00916(.A0(new_n1017_), .A1(\b[5] ), .B0(new_n1016_), .B1(\b[4] ), .Y(new_n1173_));
  OAI21X1  g00917(.A0(new_n1015_), .A1(new_n297_), .B0(new_n1173_), .Y(new_n1174_));
  AOI21X1  g00918(.A0(new_n882_), .A1(new_n349_), .B0(new_n1174_), .Y(new_n1175_));
  XOR2X1   g00919(.A(new_n1175_), .B(\a[17] ), .Y(new_n1176_));
  NAND2X1  g00920(.A(new_n1176_), .B(new_n1172_), .Y(new_n1177_));
  NAND2X1  g00921(.A(new_n1013_), .B(new_n1052_), .Y(new_n1178_));
  OAI21X1  g00922(.A0(new_n1021_), .A1(new_n1014_), .B0(new_n1178_), .Y(new_n1179_));
  XOR2X1   g00923(.A(new_n1070_), .B(new_n879_), .Y(new_n1180_));
  XOR2X1   g00924(.A(new_n1084_), .B(new_n1180_), .Y(new_n1181_));
  AND2X1   g00925(.A(new_n1084_), .B(new_n1180_), .Y(new_n1182_));
  AOI21X1  g00926(.A0(new_n1181_), .A1(new_n1179_), .B0(new_n1182_), .Y(new_n1183_));
  OR2X1    g00927(.A(new_n1176_), .B(new_n1172_), .Y(new_n1184_));
  AOI21X1  g00928(.A0(new_n1177_), .A1(new_n1184_), .B0(new_n1183_), .Y(new_n1185_));
  NAND2X1  g00929(.A(new_n1084_), .B(new_n1180_), .Y(new_n1186_));
  OAI21X1  g00930(.A0(new_n1085_), .A1(new_n1064_), .B0(new_n1186_), .Y(new_n1187_));
  NOR2X1   g00931(.A(new_n1176_), .B(new_n1172_), .Y(new_n1188_));
  AOI21X1  g00932(.A0(new_n1177_), .A1(new_n1187_), .B0(new_n1188_), .Y(new_n1189_));
  AOI21X1  g00933(.A0(new_n1189_), .A1(new_n1177_), .B0(new_n1185_), .Y(new_n1190_));
  AOI22X1  g00934(.A0(new_n818_), .A1(\b[8] ), .B0(new_n817_), .B1(\b[7] ), .Y(new_n1191_));
  OAI21X1  g00935(.A0(new_n816_), .A1(new_n392_), .B0(new_n1191_), .Y(new_n1192_));
  AOI21X1  g00936(.A0(new_n668_), .A1(new_n454_), .B0(new_n1192_), .Y(new_n1193_));
  XOR2X1   g00937(.A(new_n1193_), .B(\a[14] ), .Y(new_n1194_));
  XOR2X1   g00938(.A(new_n1194_), .B(new_n1190_), .Y(new_n1195_));
  XOR2X1   g00939(.A(new_n1195_), .B(new_n1163_), .Y(new_n1196_));
  XOR2X1   g00940(.A(new_n1196_), .B(new_n1160_), .Y(new_n1197_));
  XOR2X1   g00941(.A(new_n1197_), .B(new_n1156_), .Y(new_n1198_));
  AOI22X1  g00942(.A0(new_n469_), .A1(\b[14] ), .B0(new_n468_), .B1(\b[13] ), .Y(new_n1199_));
  OAI21X1  g00943(.A0(new_n467_), .A1(new_n713_), .B0(new_n1199_), .Y(new_n1200_));
  AOI21X1  g00944(.A0(new_n734_), .A1(new_n404_), .B0(new_n1200_), .Y(new_n1201_));
  XOR2X1   g00945(.A(new_n1201_), .B(\a[8] ), .Y(new_n1202_));
  XOR2X1   g00946(.A(new_n1202_), .B(new_n1198_), .Y(new_n1203_));
  NOR2X1   g00947(.A(new_n1100_), .B(new_n1096_), .Y(new_n1204_));
  AND2X1   g00948(.A(new_n967_), .B(new_n924_), .Y(new_n1205_));
  AOI21X1  g00949(.A0(new_n968_), .A1(new_n920_), .B0(new_n1205_), .Y(new_n1206_));
  NOR2X1   g00950(.A(new_n1034_), .B(new_n1003_), .Y(new_n1207_));
  NAND2X1  g00951(.A(new_n1034_), .B(new_n1003_), .Y(new_n1208_));
  OAI21X1  g00952(.A0(new_n1207_), .A1(new_n1206_), .B0(new_n1208_), .Y(new_n1209_));
  AOI21X1  g00953(.A0(new_n1209_), .A1(new_n1101_), .B0(new_n1204_), .Y(new_n1210_));
  XOR2X1   g00954(.A(new_n1210_), .B(new_n1203_), .Y(new_n1211_));
  XOR2X1   g00955(.A(new_n1211_), .B(new_n1154_), .Y(new_n1212_));
  XOR2X1   g00956(.A(new_n1212_), .B(new_n1150_), .Y(new_n1213_));
  NAND2X1  g00957(.A(\b[19] ), .B(\b[18] ), .Y(new_n1214_));
  OAI21X1  g00958(.A0(new_n1116_), .A1(new_n1114_), .B0(new_n1214_), .Y(new_n1215_));
  XOR2X1   g00959(.A(\b[20] ), .B(\b[19] ), .Y(new_n1216_));
  XOR2X1   g00960(.A(new_n1216_), .B(new_n1215_), .Y(new_n1217_));
  AOI22X1  g00961(.A0(new_n267_), .A1(\b[20] ), .B0(new_n266_), .B1(\b[19] ), .Y(new_n1218_));
  OAI21X1  g00962(.A0(new_n350_), .A1(new_n1115_), .B0(new_n1218_), .Y(new_n1219_));
  AOI21X1  g00963(.A0(new_n1217_), .A1(new_n318_), .B0(new_n1219_), .Y(new_n1220_));
  XOR2X1   g00964(.A(new_n1220_), .B(new_n257_), .Y(new_n1221_));
  XOR2X1   g00965(.A(new_n1221_), .B(new_n1213_), .Y(new_n1222_));
  OR2X1    g00966(.A(new_n1122_), .B(new_n1112_), .Y(new_n1223_));
  OAI21X1  g00967(.A0(new_n1138_), .A1(new_n1137_), .B0(new_n1123_), .Y(new_n1224_));
  AND2X1   g00968(.A(new_n1224_), .B(new_n1223_), .Y(new_n1225_));
  XOR2X1   g00969(.A(new_n1225_), .B(new_n1222_), .Y(\f[20] ));
  INVX1    g00970(.A(new_n1202_), .Y(new_n1227_));
  AND2X1   g00971(.A(new_n1227_), .B(new_n1198_), .Y(new_n1228_));
  XOR2X1   g00972(.A(new_n1227_), .B(new_n1198_), .Y(new_n1229_));
  OR2X1    g00973(.A(new_n1100_), .B(new_n1096_), .Y(new_n1230_));
  OAI21X1  g00974(.A0(new_n1103_), .A1(new_n1147_), .B0(new_n1230_), .Y(new_n1231_));
  AOI21X1  g00975(.A0(new_n1231_), .A1(new_n1229_), .B0(new_n1228_), .Y(new_n1232_));
  AOI22X1  g00976(.A0(new_n469_), .A1(\b[15] ), .B0(new_n468_), .B1(\b[14] ), .Y(new_n1233_));
  OAI21X1  g00977(.A0(new_n467_), .A1(new_n795_), .B0(new_n1233_), .Y(new_n1234_));
  AOI21X1  g00978(.A0(new_n794_), .A1(new_n404_), .B0(new_n1234_), .Y(new_n1235_));
  XOR2X1   g00979(.A(new_n1235_), .B(new_n400_), .Y(new_n1236_));
  NOR2X1   g00980(.A(new_n1092_), .B(new_n1088_), .Y(new_n1237_));
  NOR2X1   g00981(.A(new_n965_), .B(new_n961_), .Y(new_n1238_));
  AOI21X1  g00982(.A0(new_n966_), .A1(new_n932_), .B0(new_n1238_), .Y(new_n1239_));
  OR2X1    g00983(.A(new_n1032_), .B(new_n1028_), .Y(new_n1240_));
  AND2X1   g00984(.A(new_n1032_), .B(new_n1028_), .Y(new_n1241_));
  OAI21X1  g00985(.A0(new_n1241_), .A1(new_n1239_), .B0(new_n1240_), .Y(new_n1242_));
  AOI21X1  g00986(.A0(new_n1242_), .A1(new_n1093_), .B0(new_n1237_), .Y(new_n1243_));
  NOR2X1   g00987(.A(new_n1196_), .B(new_n1160_), .Y(new_n1244_));
  NAND2X1  g00988(.A(new_n1196_), .B(new_n1160_), .Y(new_n1245_));
  OAI21X1  g00989(.A0(new_n1244_), .A1(new_n1243_), .B0(new_n1245_), .Y(new_n1246_));
  AOI22X1  g00990(.A0(new_n603_), .A1(\b[12] ), .B0(new_n602_), .B1(\b[11] ), .Y(new_n1247_));
  OAI21X1  g00991(.A0(new_n601_), .A1(new_n587_), .B0(new_n1247_), .Y(new_n1248_));
  AOI21X1  g00992(.A0(new_n635_), .A1(new_n518_), .B0(new_n1248_), .Y(new_n1249_));
  XOR2X1   g00993(.A(new_n1249_), .B(new_n515_), .Y(new_n1250_));
  AND2X1   g00994(.A(new_n1086_), .B(new_n1061_), .Y(new_n1251_));
  AOI21X1  g00995(.A0(new_n1087_), .A1(new_n1143_), .B0(new_n1251_), .Y(new_n1252_));
  AND2X1   g00996(.A(new_n1194_), .B(new_n1190_), .Y(new_n1253_));
  OR2X1    g00997(.A(new_n1194_), .B(new_n1190_), .Y(new_n1254_));
  OAI21X1  g00998(.A0(new_n1253_), .A1(new_n1252_), .B0(new_n1254_), .Y(new_n1255_));
  NOR4X1   g00999(.A(new_n1170_), .B(new_n1083_), .C(new_n1013_), .D(new_n1072_), .Y(new_n1256_));
  XOR2X1   g01000(.A(\a[21] ), .B(\a[20] ), .Y(new_n1257_));
  NAND2X1  g01001(.A(new_n1257_), .B(\b[0] ), .Y(new_n1258_));
  INVX1    g01002(.A(new_n1258_), .Y(new_n1259_));
  XOR2X1   g01003(.A(new_n1259_), .B(new_n1256_), .Y(new_n1260_));
  INVX1    g01004(.A(new_n1167_), .Y(new_n1261_));
  AND2X1   g01005(.A(new_n1077_), .B(new_n1076_), .Y(new_n1262_));
  AND2X1   g01006(.A(new_n1079_), .B(new_n1012_), .Y(new_n1263_));
  AOI22X1  g01007(.A0(new_n1263_), .A1(\b[3] ), .B0(new_n1262_), .B1(\b[2] ), .Y(new_n1264_));
  OAI21X1  g01008(.A0(new_n1261_), .A1(new_n275_), .B0(new_n1264_), .Y(new_n1265_));
  AOI21X1  g01009(.A0(new_n1075_), .A1(new_n366_), .B0(new_n1265_), .Y(new_n1266_));
  XOR2X1   g01010(.A(new_n1266_), .B(\a[20] ), .Y(new_n1267_));
  XOR2X1   g01011(.A(new_n1267_), .B(new_n1260_), .Y(new_n1268_));
  AOI22X1  g01012(.A0(new_n1017_), .A1(\b[6] ), .B0(new_n1016_), .B1(\b[5] ), .Y(new_n1269_));
  OAI21X1  g01013(.A0(new_n1015_), .A1(new_n325_), .B0(new_n1269_), .Y(new_n1270_));
  AOI21X1  g01014(.A0(new_n882_), .A1(new_n378_), .B0(new_n1270_), .Y(new_n1271_));
  XOR2X1   g01015(.A(new_n1271_), .B(\a[17] ), .Y(new_n1272_));
  XOR2X1   g01016(.A(new_n1272_), .B(new_n1268_), .Y(new_n1273_));
  XOR2X1   g01017(.A(new_n1273_), .B(new_n1189_), .Y(new_n1274_));
  AOI22X1  g01018(.A0(new_n818_), .A1(\b[9] ), .B0(new_n817_), .B1(\b[8] ), .Y(new_n1275_));
  OAI21X1  g01019(.A0(new_n816_), .A1(new_n492_), .B0(new_n1275_), .Y(new_n1276_));
  AOI21X1  g01020(.A0(new_n668_), .A1(new_n491_), .B0(new_n1276_), .Y(new_n1277_));
  XOR2X1   g01021(.A(new_n1277_), .B(\a[14] ), .Y(new_n1278_));
  XOR2X1   g01022(.A(new_n1278_), .B(new_n1274_), .Y(new_n1279_));
  XOR2X1   g01023(.A(new_n1279_), .B(new_n1255_), .Y(new_n1280_));
  XOR2X1   g01024(.A(new_n1280_), .B(new_n1250_), .Y(new_n1281_));
  XOR2X1   g01025(.A(new_n1281_), .B(new_n1246_), .Y(new_n1282_));
  XOR2X1   g01026(.A(new_n1282_), .B(new_n1236_), .Y(new_n1283_));
  XOR2X1   g01027(.A(new_n1283_), .B(new_n1232_), .Y(new_n1284_));
  AOI22X1  g01028(.A0(new_n369_), .A1(\b[18] ), .B0(new_n368_), .B1(\b[17] ), .Y(new_n1285_));
  OAI21X1  g01029(.A0(new_n367_), .A1(new_n974_), .B0(new_n1285_), .Y(new_n1286_));
  AOI21X1  g01030(.A0(new_n1042_), .A1(new_n308_), .B0(new_n1286_), .Y(new_n1287_));
  XOR2X1   g01031(.A(new_n1287_), .B(\a[5] ), .Y(new_n1288_));
  XOR2X1   g01032(.A(new_n1288_), .B(new_n1284_), .Y(new_n1289_));
  INVX1    g01033(.A(new_n1154_), .Y(new_n1290_));
  AND2X1   g01034(.A(new_n1211_), .B(new_n1290_), .Y(new_n1291_));
  XOR2X1   g01035(.A(new_n1211_), .B(new_n1290_), .Y(new_n1292_));
  AOI21X1  g01036(.A0(new_n1292_), .A1(new_n1150_), .B0(new_n1291_), .Y(new_n1293_));
  XOR2X1   g01037(.A(new_n1293_), .B(new_n1289_), .Y(new_n1294_));
  AND2X1   g01038(.A(\b[20] ), .B(\b[19] ), .Y(new_n1295_));
  AOI21X1  g01039(.A0(new_n1216_), .A1(new_n1215_), .B0(new_n1295_), .Y(new_n1296_));
  INVX1    g01040(.A(\b[20] ), .Y(new_n1297_));
  XOR2X1   g01041(.A(\b[21] ), .B(new_n1297_), .Y(new_n1298_));
  XOR2X1   g01042(.A(new_n1298_), .B(new_n1296_), .Y(new_n1299_));
  INVX1    g01043(.A(\b[19] ), .Y(new_n1300_));
  AOI22X1  g01044(.A0(new_n267_), .A1(\b[21] ), .B0(new_n266_), .B1(\b[20] ), .Y(new_n1301_));
  OAI21X1  g01045(.A0(new_n350_), .A1(new_n1300_), .B0(new_n1301_), .Y(new_n1302_));
  AOI21X1  g01046(.A0(new_n1299_), .A1(new_n318_), .B0(new_n1302_), .Y(new_n1303_));
  XOR2X1   g01047(.A(new_n1303_), .B(\a[2] ), .Y(new_n1304_));
  XOR2X1   g01048(.A(new_n1304_), .B(new_n1294_), .Y(new_n1305_));
  INVX1    g01049(.A(new_n1221_), .Y(new_n1306_));
  NOR2X1   g01050(.A(new_n1306_), .B(new_n1213_), .Y(new_n1307_));
  AOI21X1  g01051(.A0(new_n1224_), .A1(new_n1223_), .B0(new_n1222_), .Y(new_n1308_));
  OR2X1    g01052(.A(new_n1308_), .B(new_n1307_), .Y(new_n1309_));
  XOR2X1   g01053(.A(new_n1309_), .B(new_n1305_), .Y(\f[21] ));
  OR2X1    g01054(.A(new_n1304_), .B(new_n1294_), .Y(new_n1311_));
  OAI21X1  g01055(.A0(new_n1308_), .A1(new_n1307_), .B0(new_n1305_), .Y(new_n1312_));
  AND2X1   g01056(.A(new_n1312_), .B(new_n1311_), .Y(new_n1313_));
  NAND2X1  g01057(.A(new_n1227_), .B(new_n1198_), .Y(new_n1314_));
  OAI21X1  g01058(.A0(new_n1210_), .A1(new_n1203_), .B0(new_n1314_), .Y(new_n1315_));
  AND2X1   g01059(.A(new_n1282_), .B(new_n1236_), .Y(new_n1316_));
  AOI21X1  g01060(.A0(new_n1283_), .A1(new_n1315_), .B0(new_n1316_), .Y(new_n1317_));
  AOI22X1  g01061(.A0(new_n469_), .A1(\b[16] ), .B0(new_n468_), .B1(\b[15] ), .Y(new_n1318_));
  OAI21X1  g01062(.A0(new_n467_), .A1(new_n792_), .B0(new_n1318_), .Y(new_n1319_));
  AOI21X1  g01063(.A0(new_n842_), .A1(new_n404_), .B0(new_n1319_), .Y(new_n1320_));
  XOR2X1   g01064(.A(new_n1320_), .B(new_n400_), .Y(new_n1321_));
  AND2X1   g01065(.A(new_n1196_), .B(new_n1160_), .Y(new_n1322_));
  AOI21X1  g01066(.A0(new_n1197_), .A1(new_n1156_), .B0(new_n1322_), .Y(new_n1323_));
  NOR2X1   g01067(.A(new_n1280_), .B(new_n1250_), .Y(new_n1324_));
  NAND2X1  g01068(.A(new_n1280_), .B(new_n1250_), .Y(new_n1325_));
  OAI21X1  g01069(.A0(new_n1324_), .A1(new_n1323_), .B0(new_n1325_), .Y(new_n1326_));
  OR2X1    g01070(.A(new_n1272_), .B(new_n1268_), .Y(new_n1327_));
  OR4X1    g01071(.A(new_n1170_), .B(new_n1083_), .C(new_n1013_), .D(new_n1072_), .Y(new_n1328_));
  XOR2X1   g01072(.A(new_n1259_), .B(new_n1328_), .Y(new_n1329_));
  XOR2X1   g01073(.A(new_n1267_), .B(new_n1329_), .Y(new_n1330_));
  XOR2X1   g01074(.A(new_n1272_), .B(new_n1330_), .Y(new_n1331_));
  OAI21X1  g01075(.A0(new_n1331_), .A1(new_n1189_), .B0(new_n1327_), .Y(new_n1332_));
  AOI22X1  g01076(.A0(new_n1017_), .A1(\b[7] ), .B0(new_n1016_), .B1(\b[6] ), .Y(new_n1333_));
  OAI21X1  g01077(.A0(new_n1015_), .A1(new_n395_), .B0(new_n1333_), .Y(new_n1334_));
  AOI21X1  g01078(.A0(new_n882_), .A1(new_n394_), .B0(new_n1334_), .Y(new_n1335_));
  XOR2X1   g01079(.A(new_n1335_), .B(new_n879_), .Y(new_n1336_));
  XOR2X1   g01080(.A(new_n1266_), .B(new_n1072_), .Y(new_n1337_));
  AND2X1   g01081(.A(new_n1259_), .B(new_n1256_), .Y(new_n1338_));
  AOI21X1  g01082(.A0(new_n1337_), .A1(new_n1260_), .B0(new_n1338_), .Y(new_n1339_));
  AND2X1   g01083(.A(new_n1075_), .B(new_n323_), .Y(new_n1340_));
  NOR3X1   g01084(.A(new_n1166_), .B(new_n1079_), .C(new_n277_), .Y(new_n1341_));
  OAI22X1  g01085(.A0(new_n1080_), .A1(new_n325_), .B0(new_n1078_), .B1(new_n297_), .Y(new_n1342_));
  NOR3X1   g01086(.A(new_n1342_), .B(new_n1341_), .C(new_n1340_), .Y(new_n1343_));
  XOR2X1   g01087(.A(new_n1343_), .B(\a[20] ), .Y(new_n1344_));
  NAND2X1  g01088(.A(new_n1258_), .B(\a[23] ), .Y(new_n1345_));
  XOR2X1   g01089(.A(\a[23] ), .B(\a[22] ), .Y(new_n1346_));
  AND2X1   g01090(.A(new_n1346_), .B(new_n1257_), .Y(new_n1347_));
  XOR2X1   g01091(.A(\a[21] ), .B(new_n1072_), .Y(new_n1348_));
  XOR2X1   g01092(.A(\a[22] ), .B(\a[21] ), .Y(new_n1349_));
  NAND2X1  g01093(.A(new_n1349_), .B(new_n1348_), .Y(new_n1350_));
  INVX1    g01094(.A(\a[23] ), .Y(new_n1351_));
  XOR2X1   g01095(.A(new_n1351_), .B(\a[22] ), .Y(new_n1352_));
  NAND2X1  g01096(.A(new_n1352_), .B(new_n1257_), .Y(new_n1353_));
  OAI22X1  g01097(.A0(new_n1353_), .A1(new_n275_), .B0(new_n1350_), .B1(new_n274_), .Y(new_n1354_));
  AOI21X1  g01098(.A0(new_n1347_), .A1(new_n263_), .B0(new_n1354_), .Y(new_n1355_));
  XOR2X1   g01099(.A(new_n1355_), .B(\a[23] ), .Y(new_n1356_));
  XOR2X1   g01100(.A(new_n1356_), .B(new_n1345_), .Y(new_n1357_));
  XOR2X1   g01101(.A(new_n1357_), .B(new_n1344_), .Y(new_n1358_));
  XOR2X1   g01102(.A(new_n1358_), .B(new_n1339_), .Y(new_n1359_));
  XOR2X1   g01103(.A(new_n1359_), .B(new_n1336_), .Y(new_n1360_));
  AND2X1   g01104(.A(new_n1360_), .B(new_n1332_), .Y(new_n1361_));
  NOR2X1   g01105(.A(new_n1360_), .B(new_n1332_), .Y(new_n1362_));
  OR2X1    g01106(.A(new_n1362_), .B(new_n1361_), .Y(new_n1363_));
  AOI22X1  g01107(.A0(new_n818_), .A1(\b[10] ), .B0(new_n817_), .B1(\b[9] ), .Y(new_n1364_));
  OAI21X1  g01108(.A0(new_n816_), .A1(new_n489_), .B0(new_n1364_), .Y(new_n1365_));
  AOI21X1  g01109(.A0(new_n668_), .A1(new_n543_), .B0(new_n1365_), .Y(new_n1366_));
  XOR2X1   g01110(.A(new_n1366_), .B(\a[14] ), .Y(new_n1367_));
  XOR2X1   g01111(.A(new_n1367_), .B(new_n1363_), .Y(new_n1368_));
  NOR2X1   g01112(.A(new_n1278_), .B(new_n1274_), .Y(new_n1369_));
  AOI21X1  g01113(.A0(new_n1279_), .A1(new_n1255_), .B0(new_n1369_), .Y(new_n1370_));
  XOR2X1   g01114(.A(new_n1370_), .B(new_n1368_), .Y(new_n1371_));
  AOI22X1  g01115(.A0(new_n603_), .A1(\b[13] ), .B0(new_n602_), .B1(\b[12] ), .Y(new_n1372_));
  OAI21X1  g01116(.A0(new_n601_), .A1(new_n716_), .B0(new_n1372_), .Y(new_n1373_));
  AOI21X1  g01117(.A0(new_n715_), .A1(new_n518_), .B0(new_n1373_), .Y(new_n1374_));
  XOR2X1   g01118(.A(new_n1374_), .B(\a[11] ), .Y(new_n1375_));
  XOR2X1   g01119(.A(new_n1375_), .B(new_n1371_), .Y(new_n1376_));
  XOR2X1   g01120(.A(new_n1376_), .B(new_n1326_), .Y(new_n1377_));
  XOR2X1   g01121(.A(new_n1377_), .B(new_n1321_), .Y(new_n1378_));
  XOR2X1   g01122(.A(new_n1378_), .B(new_n1317_), .Y(new_n1379_));
  AOI22X1  g01123(.A0(new_n369_), .A1(\b[19] ), .B0(new_n368_), .B1(\b[18] ), .Y(new_n1380_));
  OAI21X1  g01124(.A0(new_n367_), .A1(new_n1118_), .B0(new_n1380_), .Y(new_n1381_));
  AOI21X1  g01125(.A0(new_n1117_), .A1(new_n308_), .B0(new_n1381_), .Y(new_n1382_));
  XOR2X1   g01126(.A(new_n1382_), .B(\a[5] ), .Y(new_n1383_));
  INVX1    g01127(.A(new_n1383_), .Y(new_n1384_));
  XOR2X1   g01128(.A(new_n1384_), .B(new_n1379_), .Y(new_n1385_));
  NOR2X1   g01129(.A(new_n1288_), .B(new_n1284_), .Y(new_n1386_));
  NOR2X1   g01130(.A(new_n1108_), .B(new_n1104_), .Y(new_n1387_));
  NAND2X1  g01131(.A(new_n1036_), .B(new_n994_), .Y(new_n1388_));
  NOR2X1   g01132(.A(new_n1036_), .B(new_n994_), .Y(new_n1389_));
  OAI21X1  g01133(.A0(new_n1389_), .A1(new_n1135_), .B0(new_n1388_), .Y(new_n1390_));
  AOI21X1  g01134(.A0(new_n1390_), .A1(new_n1109_), .B0(new_n1387_), .Y(new_n1391_));
  NAND2X1  g01135(.A(new_n1211_), .B(new_n1290_), .Y(new_n1392_));
  OAI21X1  g01136(.A0(new_n1212_), .A1(new_n1391_), .B0(new_n1392_), .Y(new_n1393_));
  AOI21X1  g01137(.A0(new_n1393_), .A1(new_n1289_), .B0(new_n1386_), .Y(new_n1394_));
  XOR2X1   g01138(.A(new_n1394_), .B(new_n1385_), .Y(new_n1395_));
  NAND2X1  g01139(.A(\b[21] ), .B(\b[20] ), .Y(new_n1396_));
  OAI21X1  g01140(.A0(new_n1298_), .A1(new_n1296_), .B0(new_n1396_), .Y(new_n1397_));
  XOR2X1   g01141(.A(\b[22] ), .B(\b[21] ), .Y(new_n1398_));
  XOR2X1   g01142(.A(new_n1398_), .B(new_n1397_), .Y(new_n1399_));
  AOI22X1  g01143(.A0(new_n267_), .A1(\b[22] ), .B0(new_n266_), .B1(\b[21] ), .Y(new_n1400_));
  OAI21X1  g01144(.A0(new_n350_), .A1(new_n1297_), .B0(new_n1400_), .Y(new_n1401_));
  AOI21X1  g01145(.A0(new_n1399_), .A1(new_n318_), .B0(new_n1401_), .Y(new_n1402_));
  XOR2X1   g01146(.A(new_n1402_), .B(\a[2] ), .Y(new_n1403_));
  XOR2X1   g01147(.A(new_n1403_), .B(new_n1395_), .Y(new_n1404_));
  XOR2X1   g01148(.A(new_n1404_), .B(new_n1313_), .Y(\f[22] ));
  NAND2X1  g01149(.A(new_n1377_), .B(new_n1321_), .Y(new_n1406_));
  NOR2X1   g01150(.A(new_n1377_), .B(new_n1321_), .Y(new_n1407_));
  OAI21X1  g01151(.A0(new_n1407_), .A1(new_n1317_), .B0(new_n1406_), .Y(new_n1408_));
  AOI22X1  g01152(.A0(new_n469_), .A1(\b[17] ), .B0(new_n468_), .B1(\b[16] ), .Y(new_n1409_));
  OAI21X1  g01153(.A0(new_n467_), .A1(new_n977_), .B0(new_n1409_), .Y(new_n1410_));
  AOI21X1  g01154(.A0(new_n976_), .A1(new_n404_), .B0(new_n1410_), .Y(new_n1411_));
  XOR2X1   g01155(.A(new_n1411_), .B(\a[8] ), .Y(new_n1412_));
  OR2X1    g01156(.A(new_n1367_), .B(new_n1363_), .Y(new_n1413_));
  XOR2X1   g01157(.A(new_n1360_), .B(new_n1332_), .Y(new_n1414_));
  XOR2X1   g01158(.A(new_n1367_), .B(new_n1414_), .Y(new_n1415_));
  OAI21X1  g01159(.A0(new_n1370_), .A1(new_n1415_), .B0(new_n1413_), .Y(new_n1416_));
  AOI22X1  g01160(.A0(new_n818_), .A1(\b[11] ), .B0(new_n817_), .B1(\b[10] ), .Y(new_n1417_));
  OAI21X1  g01161(.A0(new_n816_), .A1(new_n590_), .B0(new_n1417_), .Y(new_n1418_));
  AOI21X1  g01162(.A0(new_n668_), .A1(new_n589_), .B0(new_n1418_), .Y(new_n1419_));
  XOR2X1   g01163(.A(new_n1419_), .B(new_n665_), .Y(new_n1420_));
  NAND2X1  g01164(.A(new_n1359_), .B(new_n1336_), .Y(new_n1421_));
  NAND2X1  g01165(.A(new_n1360_), .B(new_n1332_), .Y(new_n1422_));
  NAND2X1  g01166(.A(new_n1422_), .B(new_n1421_), .Y(new_n1423_));
  INVX1    g01167(.A(new_n1344_), .Y(new_n1424_));
  NAND2X1  g01168(.A(new_n1357_), .B(new_n1424_), .Y(new_n1425_));
  OAI21X1  g01169(.A0(new_n1358_), .A1(new_n1339_), .B0(new_n1425_), .Y(new_n1426_));
  NOR2X1   g01170(.A(new_n1356_), .B(new_n1345_), .Y(new_n1427_));
  INVX1    g01171(.A(new_n1347_), .Y(new_n1428_));
  OR2X1    g01172(.A(new_n1349_), .B(new_n1257_), .Y(new_n1429_));
  NOR2X1   g01173(.A(new_n1429_), .B(new_n1352_), .Y(new_n1430_));
  OAI22X1  g01174(.A0(new_n1353_), .A1(new_n277_), .B0(new_n1350_), .B1(new_n275_), .Y(new_n1431_));
  AOI21X1  g01175(.A0(new_n1430_), .A1(\b[0] ), .B0(new_n1431_), .Y(new_n1432_));
  OAI21X1  g01176(.A0(new_n1428_), .A1(new_n281_), .B0(new_n1432_), .Y(new_n1433_));
  XOR2X1   g01177(.A(new_n1433_), .B(new_n1351_), .Y(new_n1434_));
  XOR2X1   g01178(.A(new_n1434_), .B(new_n1427_), .Y(new_n1435_));
  AOI22X1  g01179(.A0(new_n1263_), .A1(\b[5] ), .B0(new_n1262_), .B1(\b[4] ), .Y(new_n1436_));
  OAI21X1  g01180(.A0(new_n1261_), .A1(new_n297_), .B0(new_n1436_), .Y(new_n1437_));
  AOI21X1  g01181(.A0(new_n1075_), .A1(new_n349_), .B0(new_n1437_), .Y(new_n1438_));
  XOR2X1   g01182(.A(new_n1438_), .B(\a[20] ), .Y(new_n1439_));
  NAND2X1  g01183(.A(new_n1439_), .B(new_n1435_), .Y(new_n1440_));
  NOR2X1   g01184(.A(new_n1439_), .B(new_n1435_), .Y(new_n1441_));
  AND2X1   g01185(.A(new_n1439_), .B(new_n1435_), .Y(new_n1442_));
  OR2X1    g01186(.A(new_n1442_), .B(new_n1441_), .Y(new_n1443_));
  AOI21X1  g01187(.A0(new_n1440_), .A1(new_n1426_), .B0(new_n1441_), .Y(new_n1444_));
  AOI22X1  g01188(.A0(new_n1444_), .A1(new_n1440_), .B0(new_n1443_), .B1(new_n1426_), .Y(new_n1445_));
  AOI22X1  g01189(.A0(new_n1017_), .A1(\b[8] ), .B0(new_n1016_), .B1(\b[7] ), .Y(new_n1446_));
  OAI21X1  g01190(.A0(new_n1015_), .A1(new_n392_), .B0(new_n1446_), .Y(new_n1447_));
  AOI21X1  g01191(.A0(new_n882_), .A1(new_n454_), .B0(new_n1447_), .Y(new_n1448_));
  XOR2X1   g01192(.A(new_n1448_), .B(\a[17] ), .Y(new_n1449_));
  XOR2X1   g01193(.A(new_n1449_), .B(new_n1445_), .Y(new_n1450_));
  XOR2X1   g01194(.A(new_n1450_), .B(new_n1423_), .Y(new_n1451_));
  XOR2X1   g01195(.A(new_n1451_), .B(new_n1420_), .Y(new_n1452_));
  XOR2X1   g01196(.A(new_n1452_), .B(new_n1416_), .Y(new_n1453_));
  AOI22X1  g01197(.A0(new_n603_), .A1(\b[14] ), .B0(new_n602_), .B1(\b[13] ), .Y(new_n1454_));
  OAI21X1  g01198(.A0(new_n601_), .A1(new_n713_), .B0(new_n1454_), .Y(new_n1455_));
  AOI21X1  g01199(.A0(new_n734_), .A1(new_n518_), .B0(new_n1455_), .Y(new_n1456_));
  XOR2X1   g01200(.A(new_n1456_), .B(\a[11] ), .Y(new_n1457_));
  XOR2X1   g01201(.A(new_n1457_), .B(new_n1453_), .Y(new_n1458_));
  NOR2X1   g01202(.A(new_n1375_), .B(new_n1371_), .Y(new_n1459_));
  AOI21X1  g01203(.A0(new_n1376_), .A1(new_n1326_), .B0(new_n1459_), .Y(new_n1460_));
  XOR2X1   g01204(.A(new_n1460_), .B(new_n1458_), .Y(new_n1461_));
  XOR2X1   g01205(.A(new_n1461_), .B(new_n1412_), .Y(new_n1462_));
  XOR2X1   g01206(.A(new_n1462_), .B(new_n1408_), .Y(new_n1463_));
  AOI22X1  g01207(.A0(new_n369_), .A1(\b[20] ), .B0(new_n368_), .B1(\b[19] ), .Y(new_n1464_));
  OAI21X1  g01208(.A0(new_n367_), .A1(new_n1115_), .B0(new_n1464_), .Y(new_n1465_));
  AOI21X1  g01209(.A0(new_n1217_), .A1(new_n308_), .B0(new_n1465_), .Y(new_n1466_));
  XOR2X1   g01210(.A(new_n1466_), .B(\a[5] ), .Y(new_n1467_));
  XOR2X1   g01211(.A(new_n1467_), .B(new_n1463_), .Y(new_n1468_));
  NOR2X1   g01212(.A(new_n1383_), .B(new_n1379_), .Y(new_n1469_));
  XOR2X1   g01213(.A(new_n1383_), .B(new_n1379_), .Y(new_n1470_));
  OR2X1    g01214(.A(new_n1288_), .B(new_n1284_), .Y(new_n1471_));
  XOR2X1   g01215(.A(new_n1283_), .B(new_n1315_), .Y(new_n1472_));
  XOR2X1   g01216(.A(new_n1288_), .B(new_n1472_), .Y(new_n1473_));
  OAI21X1  g01217(.A0(new_n1293_), .A1(new_n1473_), .B0(new_n1471_), .Y(new_n1474_));
  AOI21X1  g01218(.A0(new_n1474_), .A1(new_n1470_), .B0(new_n1469_), .Y(new_n1475_));
  XOR2X1   g01219(.A(new_n1475_), .B(new_n1468_), .Y(new_n1476_));
  AND2X1   g01220(.A(\b[22] ), .B(\b[21] ), .Y(new_n1477_));
  AOI21X1  g01221(.A0(new_n1398_), .A1(new_n1397_), .B0(new_n1477_), .Y(new_n1478_));
  INVX1    g01222(.A(\b[22] ), .Y(new_n1479_));
  XOR2X1   g01223(.A(\b[23] ), .B(new_n1479_), .Y(new_n1480_));
  XOR2X1   g01224(.A(new_n1480_), .B(new_n1478_), .Y(new_n1481_));
  INVX1    g01225(.A(\b[21] ), .Y(new_n1482_));
  AOI22X1  g01226(.A0(new_n267_), .A1(\b[23] ), .B0(new_n266_), .B1(\b[22] ), .Y(new_n1483_));
  OAI21X1  g01227(.A0(new_n350_), .A1(new_n1482_), .B0(new_n1483_), .Y(new_n1484_));
  AOI21X1  g01228(.A0(new_n1481_), .A1(new_n318_), .B0(new_n1484_), .Y(new_n1485_));
  XOR2X1   g01229(.A(new_n1485_), .B(\a[2] ), .Y(new_n1486_));
  XOR2X1   g01230(.A(new_n1486_), .B(new_n1476_), .Y(new_n1487_));
  XOR2X1   g01231(.A(new_n1394_), .B(new_n1470_), .Y(new_n1488_));
  NOR2X1   g01232(.A(new_n1403_), .B(new_n1488_), .Y(new_n1489_));
  AOI21X1  g01233(.A0(new_n1312_), .A1(new_n1311_), .B0(new_n1404_), .Y(new_n1490_));
  OR2X1    g01234(.A(new_n1490_), .B(new_n1489_), .Y(new_n1491_));
  XOR2X1   g01235(.A(new_n1491_), .B(new_n1487_), .Y(\f[23] ));
  OR2X1    g01236(.A(new_n1467_), .B(new_n1463_), .Y(new_n1493_));
  NAND2X1  g01237(.A(new_n1282_), .B(new_n1236_), .Y(new_n1494_));
  NOR2X1   g01238(.A(new_n1282_), .B(new_n1236_), .Y(new_n1495_));
  OAI21X1  g01239(.A0(new_n1495_), .A1(new_n1232_), .B0(new_n1494_), .Y(new_n1496_));
  AND2X1   g01240(.A(new_n1377_), .B(new_n1321_), .Y(new_n1497_));
  AOI21X1  g01241(.A0(new_n1378_), .A1(new_n1496_), .B0(new_n1497_), .Y(new_n1498_));
  XOR2X1   g01242(.A(new_n1462_), .B(new_n1498_), .Y(new_n1499_));
  XOR2X1   g01243(.A(new_n1467_), .B(new_n1499_), .Y(new_n1500_));
  OAI21X1  g01244(.A0(new_n1475_), .A1(new_n1500_), .B0(new_n1493_), .Y(new_n1501_));
  AOI22X1  g01245(.A0(new_n369_), .A1(\b[21] ), .B0(new_n368_), .B1(\b[20] ), .Y(new_n1502_));
  OAI21X1  g01246(.A0(new_n367_), .A1(new_n1300_), .B0(new_n1502_), .Y(new_n1503_));
  AOI21X1  g01247(.A0(new_n1299_), .A1(new_n308_), .B0(new_n1503_), .Y(new_n1504_));
  XOR2X1   g01248(.A(new_n1504_), .B(\a[5] ), .Y(new_n1505_));
  INVX1    g01249(.A(new_n1412_), .Y(new_n1506_));
  NAND2X1  g01250(.A(new_n1461_), .B(new_n1506_), .Y(new_n1507_));
  OAI21X1  g01251(.A0(new_n1462_), .A1(new_n1498_), .B0(new_n1507_), .Y(new_n1508_));
  AND2X1   g01252(.A(new_n1451_), .B(new_n1420_), .Y(new_n1509_));
  AOI21X1  g01253(.A0(new_n1452_), .A1(new_n1416_), .B0(new_n1509_), .Y(new_n1510_));
  AOI22X1  g01254(.A0(new_n818_), .A1(\b[12] ), .B0(new_n817_), .B1(\b[11] ), .Y(new_n1511_));
  OAI21X1  g01255(.A0(new_n816_), .A1(new_n587_), .B0(new_n1511_), .Y(new_n1512_));
  AOI21X1  g01256(.A0(new_n668_), .A1(new_n635_), .B0(new_n1512_), .Y(new_n1513_));
  XOR2X1   g01257(.A(new_n1513_), .B(new_n665_), .Y(new_n1514_));
  AND2X1   g01258(.A(new_n1422_), .B(new_n1421_), .Y(new_n1515_));
  AND2X1   g01259(.A(new_n1449_), .B(new_n1445_), .Y(new_n1516_));
  OR2X1    g01260(.A(new_n1449_), .B(new_n1445_), .Y(new_n1517_));
  OAI21X1  g01261(.A0(new_n1516_), .A1(new_n1515_), .B0(new_n1517_), .Y(new_n1518_));
  OR4X1    g01262(.A(new_n1433_), .B(new_n1356_), .C(new_n1259_), .D(new_n1351_), .Y(new_n1519_));
  XOR2X1   g01263(.A(\a[24] ), .B(\a[23] ), .Y(new_n1520_));
  NAND2X1  g01264(.A(new_n1520_), .B(\b[0] ), .Y(new_n1521_));
  INVX1    g01265(.A(new_n1521_), .Y(new_n1522_));
  XOR2X1   g01266(.A(new_n1522_), .B(new_n1519_), .Y(new_n1523_));
  INVX1    g01267(.A(new_n1430_), .Y(new_n1524_));
  AND2X1   g01268(.A(new_n1349_), .B(new_n1348_), .Y(new_n1525_));
  AND2X1   g01269(.A(new_n1352_), .B(new_n1257_), .Y(new_n1526_));
  AOI22X1  g01270(.A0(new_n1526_), .A1(\b[3] ), .B0(new_n1525_), .B1(\b[2] ), .Y(new_n1527_));
  OAI21X1  g01271(.A0(new_n1524_), .A1(new_n275_), .B0(new_n1527_), .Y(new_n1528_));
  AOI21X1  g01272(.A0(new_n1347_), .A1(new_n366_), .B0(new_n1528_), .Y(new_n1529_));
  XOR2X1   g01273(.A(new_n1529_), .B(\a[23] ), .Y(new_n1530_));
  XOR2X1   g01274(.A(new_n1530_), .B(new_n1523_), .Y(new_n1531_));
  AOI22X1  g01275(.A0(new_n1263_), .A1(\b[6] ), .B0(new_n1262_), .B1(\b[5] ), .Y(new_n1532_));
  OAI21X1  g01276(.A0(new_n1261_), .A1(new_n325_), .B0(new_n1532_), .Y(new_n1533_));
  AOI21X1  g01277(.A0(new_n1075_), .A1(new_n378_), .B0(new_n1533_), .Y(new_n1534_));
  XOR2X1   g01278(.A(new_n1534_), .B(new_n1072_), .Y(new_n1535_));
  XOR2X1   g01279(.A(new_n1535_), .B(new_n1531_), .Y(new_n1536_));
  XOR2X1   g01280(.A(new_n1536_), .B(new_n1444_), .Y(new_n1537_));
  AOI22X1  g01281(.A0(new_n1017_), .A1(\b[9] ), .B0(new_n1016_), .B1(\b[8] ), .Y(new_n1538_));
  OAI21X1  g01282(.A0(new_n1015_), .A1(new_n492_), .B0(new_n1538_), .Y(new_n1539_));
  AOI21X1  g01283(.A0(new_n882_), .A1(new_n491_), .B0(new_n1539_), .Y(new_n1540_));
  XOR2X1   g01284(.A(new_n1540_), .B(\a[17] ), .Y(new_n1541_));
  XOR2X1   g01285(.A(new_n1541_), .B(new_n1537_), .Y(new_n1542_));
  XOR2X1   g01286(.A(new_n1542_), .B(new_n1518_), .Y(new_n1543_));
  XOR2X1   g01287(.A(new_n1543_), .B(new_n1514_), .Y(new_n1544_));
  XOR2X1   g01288(.A(new_n1544_), .B(new_n1510_), .Y(new_n1545_));
  AOI22X1  g01289(.A0(new_n603_), .A1(\b[15] ), .B0(new_n602_), .B1(\b[14] ), .Y(new_n1546_));
  OAI21X1  g01290(.A0(new_n601_), .A1(new_n795_), .B0(new_n1546_), .Y(new_n1547_));
  AOI21X1  g01291(.A0(new_n794_), .A1(new_n518_), .B0(new_n1547_), .Y(new_n1548_));
  XOR2X1   g01292(.A(new_n1548_), .B(\a[11] ), .Y(new_n1549_));
  XOR2X1   g01293(.A(new_n1549_), .B(new_n1545_), .Y(new_n1550_));
  INVX1    g01294(.A(new_n1457_), .Y(new_n1551_));
  AND2X1   g01295(.A(new_n1551_), .B(new_n1453_), .Y(new_n1552_));
  XOR2X1   g01296(.A(new_n1551_), .B(new_n1453_), .Y(new_n1553_));
  AND2X1   g01297(.A(new_n1280_), .B(new_n1250_), .Y(new_n1554_));
  AOI21X1  g01298(.A0(new_n1281_), .A1(new_n1246_), .B0(new_n1554_), .Y(new_n1555_));
  AND2X1   g01299(.A(new_n1375_), .B(new_n1371_), .Y(new_n1556_));
  OR2X1    g01300(.A(new_n1375_), .B(new_n1371_), .Y(new_n1557_));
  OAI21X1  g01301(.A0(new_n1556_), .A1(new_n1555_), .B0(new_n1557_), .Y(new_n1558_));
  AOI21X1  g01302(.A0(new_n1558_), .A1(new_n1553_), .B0(new_n1552_), .Y(new_n1559_));
  XOR2X1   g01303(.A(new_n1559_), .B(new_n1550_), .Y(new_n1560_));
  AOI22X1  g01304(.A0(new_n469_), .A1(\b[18] ), .B0(new_n468_), .B1(\b[17] ), .Y(new_n1561_));
  OAI21X1  g01305(.A0(new_n467_), .A1(new_n974_), .B0(new_n1561_), .Y(new_n1562_));
  AOI21X1  g01306(.A0(new_n1042_), .A1(new_n404_), .B0(new_n1562_), .Y(new_n1563_));
  XOR2X1   g01307(.A(new_n1563_), .B(\a[8] ), .Y(new_n1564_));
  XOR2X1   g01308(.A(new_n1564_), .B(new_n1560_), .Y(new_n1565_));
  XOR2X1   g01309(.A(new_n1565_), .B(new_n1508_), .Y(new_n1566_));
  XOR2X1   g01310(.A(new_n1566_), .B(new_n1505_), .Y(new_n1567_));
  XOR2X1   g01311(.A(new_n1567_), .B(new_n1501_), .Y(new_n1568_));
  NAND2X1  g01312(.A(\b[23] ), .B(\b[22] ), .Y(new_n1569_));
  OAI21X1  g01313(.A0(new_n1480_), .A1(new_n1478_), .B0(new_n1569_), .Y(new_n1570_));
  XOR2X1   g01314(.A(\b[24] ), .B(\b[23] ), .Y(new_n1571_));
  XOR2X1   g01315(.A(new_n1571_), .B(new_n1570_), .Y(new_n1572_));
  AOI22X1  g01316(.A0(new_n267_), .A1(\b[24] ), .B0(new_n266_), .B1(\b[23] ), .Y(new_n1573_));
  OAI21X1  g01317(.A0(new_n350_), .A1(new_n1479_), .B0(new_n1573_), .Y(new_n1574_));
  AOI21X1  g01318(.A0(new_n1572_), .A1(new_n318_), .B0(new_n1574_), .Y(new_n1575_));
  XOR2X1   g01319(.A(new_n1575_), .B(new_n257_), .Y(new_n1576_));
  XOR2X1   g01320(.A(new_n1576_), .B(new_n1568_), .Y(new_n1577_));
  OR2X1    g01321(.A(new_n1486_), .B(new_n1476_), .Y(new_n1578_));
  OAI21X1  g01322(.A0(new_n1490_), .A1(new_n1489_), .B0(new_n1487_), .Y(new_n1579_));
  AND2X1   g01323(.A(new_n1579_), .B(new_n1578_), .Y(new_n1580_));
  XOR2X1   g01324(.A(new_n1580_), .B(new_n1577_), .Y(\f[24] ));
  INVX1    g01325(.A(new_n1576_), .Y(new_n1582_));
  NOR2X1   g01326(.A(new_n1582_), .B(new_n1568_), .Y(new_n1583_));
  AOI21X1  g01327(.A0(new_n1579_), .A1(new_n1578_), .B0(new_n1577_), .Y(new_n1584_));
  OR2X1    g01328(.A(new_n1584_), .B(new_n1583_), .Y(new_n1585_));
  AND2X1   g01329(.A(\b[24] ), .B(\b[23] ), .Y(new_n1586_));
  AOI21X1  g01330(.A0(new_n1571_), .A1(new_n1570_), .B0(new_n1586_), .Y(new_n1587_));
  INVX1    g01331(.A(\b[24] ), .Y(new_n1588_));
  XOR2X1   g01332(.A(\b[25] ), .B(new_n1588_), .Y(new_n1589_));
  XOR2X1   g01333(.A(new_n1589_), .B(new_n1587_), .Y(new_n1590_));
  INVX1    g01334(.A(\b[23] ), .Y(new_n1591_));
  AOI22X1  g01335(.A0(new_n267_), .A1(\b[25] ), .B0(new_n266_), .B1(\b[24] ), .Y(new_n1592_));
  OAI21X1  g01336(.A0(new_n350_), .A1(new_n1591_), .B0(new_n1592_), .Y(new_n1593_));
  AOI21X1  g01337(.A0(new_n1590_), .A1(new_n318_), .B0(new_n1593_), .Y(new_n1594_));
  XOR2X1   g01338(.A(new_n1594_), .B(new_n257_), .Y(new_n1595_));
  INVX1    g01339(.A(new_n1505_), .Y(new_n1596_));
  AND2X1   g01340(.A(new_n1566_), .B(new_n1596_), .Y(new_n1597_));
  XOR2X1   g01341(.A(new_n1566_), .B(new_n1596_), .Y(new_n1598_));
  AOI21X1  g01342(.A0(new_n1598_), .A1(new_n1501_), .B0(new_n1597_), .Y(new_n1599_));
  NAND2X1  g01343(.A(new_n1535_), .B(new_n1531_), .Y(new_n1600_));
  XOR2X1   g01344(.A(new_n1534_), .B(\a[20] ), .Y(new_n1601_));
  XOR2X1   g01345(.A(new_n1601_), .B(new_n1531_), .Y(new_n1602_));
  OAI21X1  g01346(.A0(new_n1602_), .A1(new_n1444_), .B0(new_n1600_), .Y(new_n1603_));
  AOI22X1  g01347(.A0(new_n1263_), .A1(\b[7] ), .B0(new_n1262_), .B1(\b[6] ), .Y(new_n1604_));
  OAI21X1  g01348(.A0(new_n1261_), .A1(new_n395_), .B0(new_n1604_), .Y(new_n1605_));
  AOI21X1  g01349(.A0(new_n1075_), .A1(new_n394_), .B0(new_n1605_), .Y(new_n1606_));
  XOR2X1   g01350(.A(new_n1606_), .B(new_n1072_), .Y(new_n1607_));
  OR2X1    g01351(.A(new_n1521_), .B(new_n1519_), .Y(new_n1608_));
  OAI21X1  g01352(.A0(new_n1530_), .A1(new_n1523_), .B0(new_n1608_), .Y(new_n1609_));
  AND2X1   g01353(.A(new_n1347_), .B(new_n323_), .Y(new_n1610_));
  NOR3X1   g01354(.A(new_n1429_), .B(new_n1352_), .C(new_n277_), .Y(new_n1611_));
  OAI22X1  g01355(.A0(new_n1353_), .A1(new_n325_), .B0(new_n1350_), .B1(new_n297_), .Y(new_n1612_));
  NOR3X1   g01356(.A(new_n1612_), .B(new_n1611_), .C(new_n1610_), .Y(new_n1613_));
  XOR2X1   g01357(.A(new_n1613_), .B(new_n1351_), .Y(new_n1614_));
  NAND2X1  g01358(.A(new_n1521_), .B(\a[26] ), .Y(new_n1615_));
  XOR2X1   g01359(.A(\a[26] ), .B(\a[25] ), .Y(new_n1616_));
  AND2X1   g01360(.A(new_n1616_), .B(new_n1520_), .Y(new_n1617_));
  XOR2X1   g01361(.A(\a[24] ), .B(new_n1351_), .Y(new_n1618_));
  XOR2X1   g01362(.A(\a[25] ), .B(\a[24] ), .Y(new_n1619_));
  NAND2X1  g01363(.A(new_n1619_), .B(new_n1618_), .Y(new_n1620_));
  INVX1    g01364(.A(\a[26] ), .Y(new_n1621_));
  XOR2X1   g01365(.A(new_n1621_), .B(\a[25] ), .Y(new_n1622_));
  NAND2X1  g01366(.A(new_n1622_), .B(new_n1520_), .Y(new_n1623_));
  OAI22X1  g01367(.A0(new_n1623_), .A1(new_n275_), .B0(new_n1620_), .B1(new_n274_), .Y(new_n1624_));
  AOI21X1  g01368(.A0(new_n1617_), .A1(new_n263_), .B0(new_n1624_), .Y(new_n1625_));
  XOR2X1   g01369(.A(new_n1625_), .B(\a[26] ), .Y(new_n1626_));
  XOR2X1   g01370(.A(new_n1626_), .B(new_n1615_), .Y(new_n1627_));
  XOR2X1   g01371(.A(new_n1627_), .B(new_n1614_), .Y(new_n1628_));
  XOR2X1   g01372(.A(new_n1628_), .B(new_n1609_), .Y(new_n1629_));
  XOR2X1   g01373(.A(new_n1629_), .B(new_n1607_), .Y(new_n1630_));
  XOR2X1   g01374(.A(new_n1630_), .B(new_n1603_), .Y(new_n1631_));
  AOI22X1  g01375(.A0(new_n1017_), .A1(\b[10] ), .B0(new_n1016_), .B1(\b[9] ), .Y(new_n1632_));
  OAI21X1  g01376(.A0(new_n1015_), .A1(new_n489_), .B0(new_n1632_), .Y(new_n1633_));
  AOI21X1  g01377(.A0(new_n882_), .A1(new_n543_), .B0(new_n1633_), .Y(new_n1634_));
  XOR2X1   g01378(.A(new_n1634_), .B(\a[17] ), .Y(new_n1635_));
  XOR2X1   g01379(.A(new_n1635_), .B(new_n1631_), .Y(new_n1636_));
  NOR2X1   g01380(.A(new_n1541_), .B(new_n1537_), .Y(new_n1637_));
  AOI21X1  g01381(.A0(new_n1542_), .A1(new_n1518_), .B0(new_n1637_), .Y(new_n1638_));
  XOR2X1   g01382(.A(new_n1638_), .B(new_n1636_), .Y(new_n1639_));
  AOI22X1  g01383(.A0(new_n818_), .A1(\b[13] ), .B0(new_n817_), .B1(\b[12] ), .Y(new_n1640_));
  OAI21X1  g01384(.A0(new_n816_), .A1(new_n716_), .B0(new_n1640_), .Y(new_n1641_));
  AOI21X1  g01385(.A0(new_n715_), .A1(new_n668_), .B0(new_n1641_), .Y(new_n1642_));
  XOR2X1   g01386(.A(new_n1642_), .B(\a[14] ), .Y(new_n1643_));
  XOR2X1   g01387(.A(new_n1643_), .B(new_n1639_), .Y(new_n1644_));
  NOR3X1   g01388(.A(new_n1367_), .B(new_n1362_), .C(new_n1361_), .Y(new_n1645_));
  NOR2X1   g01389(.A(new_n1194_), .B(new_n1190_), .Y(new_n1646_));
  AOI21X1  g01390(.A0(new_n1195_), .A1(new_n1163_), .B0(new_n1646_), .Y(new_n1647_));
  OR2X1    g01391(.A(new_n1278_), .B(new_n1274_), .Y(new_n1648_));
  AND2X1   g01392(.A(new_n1278_), .B(new_n1274_), .Y(new_n1649_));
  OAI21X1  g01393(.A0(new_n1649_), .A1(new_n1647_), .B0(new_n1648_), .Y(new_n1650_));
  AOI21X1  g01394(.A0(new_n1650_), .A1(new_n1368_), .B0(new_n1645_), .Y(new_n1651_));
  NOR2X1   g01395(.A(new_n1451_), .B(new_n1420_), .Y(new_n1652_));
  NAND2X1  g01396(.A(new_n1451_), .B(new_n1420_), .Y(new_n1653_));
  OAI21X1  g01397(.A0(new_n1652_), .A1(new_n1651_), .B0(new_n1653_), .Y(new_n1654_));
  AND2X1   g01398(.A(new_n1543_), .B(new_n1514_), .Y(new_n1655_));
  AOI21X1  g01399(.A0(new_n1544_), .A1(new_n1654_), .B0(new_n1655_), .Y(new_n1656_));
  XOR2X1   g01400(.A(new_n1656_), .B(new_n1644_), .Y(new_n1657_));
  AOI22X1  g01401(.A0(new_n603_), .A1(\b[16] ), .B0(new_n602_), .B1(\b[15] ), .Y(new_n1658_));
  OAI21X1  g01402(.A0(new_n601_), .A1(new_n792_), .B0(new_n1658_), .Y(new_n1659_));
  AOI21X1  g01403(.A0(new_n842_), .A1(new_n518_), .B0(new_n1659_), .Y(new_n1660_));
  XOR2X1   g01404(.A(new_n1660_), .B(\a[11] ), .Y(new_n1661_));
  XOR2X1   g01405(.A(new_n1661_), .B(new_n1657_), .Y(new_n1662_));
  NOR2X1   g01406(.A(new_n1549_), .B(new_n1545_), .Y(new_n1663_));
  NAND2X1  g01407(.A(new_n1551_), .B(new_n1453_), .Y(new_n1664_));
  OAI21X1  g01408(.A0(new_n1460_), .A1(new_n1458_), .B0(new_n1664_), .Y(new_n1665_));
  AOI21X1  g01409(.A0(new_n1665_), .A1(new_n1550_), .B0(new_n1663_), .Y(new_n1666_));
  XOR2X1   g01410(.A(new_n1666_), .B(new_n1662_), .Y(new_n1667_));
  AOI22X1  g01411(.A0(new_n469_), .A1(\b[19] ), .B0(new_n468_), .B1(\b[18] ), .Y(new_n1668_));
  OAI21X1  g01412(.A0(new_n467_), .A1(new_n1118_), .B0(new_n1668_), .Y(new_n1669_));
  AOI21X1  g01413(.A0(new_n1117_), .A1(new_n404_), .B0(new_n1669_), .Y(new_n1670_));
  XOR2X1   g01414(.A(new_n1670_), .B(\a[8] ), .Y(new_n1671_));
  XOR2X1   g01415(.A(new_n1671_), .B(new_n1667_), .Y(new_n1672_));
  NOR2X1   g01416(.A(new_n1564_), .B(new_n1560_), .Y(new_n1673_));
  AOI21X1  g01417(.A0(new_n1565_), .A1(new_n1508_), .B0(new_n1673_), .Y(new_n1674_));
  XOR2X1   g01418(.A(new_n1674_), .B(new_n1672_), .Y(new_n1675_));
  AOI22X1  g01419(.A0(new_n369_), .A1(\b[22] ), .B0(new_n368_), .B1(\b[21] ), .Y(new_n1676_));
  OAI21X1  g01420(.A0(new_n367_), .A1(new_n1297_), .B0(new_n1676_), .Y(new_n1677_));
  AOI21X1  g01421(.A0(new_n1399_), .A1(new_n308_), .B0(new_n1677_), .Y(new_n1678_));
  XOR2X1   g01422(.A(new_n1678_), .B(\a[5] ), .Y(new_n1679_));
  XOR2X1   g01423(.A(new_n1679_), .B(new_n1675_), .Y(new_n1680_));
  XOR2X1   g01424(.A(new_n1680_), .B(new_n1599_), .Y(new_n1681_));
  XOR2X1   g01425(.A(new_n1681_), .B(new_n1595_), .Y(new_n1682_));
  XOR2X1   g01426(.A(new_n1682_), .B(new_n1585_), .Y(\f[25] ));
  NAND2X1  g01427(.A(new_n1681_), .B(new_n1595_), .Y(new_n1684_));
  OAI21X1  g01428(.A0(new_n1584_), .A1(new_n1583_), .B0(new_n1682_), .Y(new_n1685_));
  AND2X1   g01429(.A(new_n1685_), .B(new_n1684_), .Y(new_n1686_));
  NOR2X1   g01430(.A(new_n1467_), .B(new_n1463_), .Y(new_n1687_));
  OR2X1    g01431(.A(new_n1383_), .B(new_n1379_), .Y(new_n1688_));
  OAI21X1  g01432(.A0(new_n1394_), .A1(new_n1385_), .B0(new_n1688_), .Y(new_n1689_));
  AOI21X1  g01433(.A0(new_n1689_), .A1(new_n1468_), .B0(new_n1687_), .Y(new_n1690_));
  NAND2X1  g01434(.A(new_n1566_), .B(new_n1596_), .Y(new_n1691_));
  OAI21X1  g01435(.A0(new_n1567_), .A1(new_n1690_), .B0(new_n1691_), .Y(new_n1692_));
  AND2X1   g01436(.A(new_n1630_), .B(new_n1603_), .Y(new_n1693_));
  NOR2X1   g01437(.A(new_n1630_), .B(new_n1603_), .Y(new_n1694_));
  OR2X1    g01438(.A(new_n1694_), .B(new_n1693_), .Y(new_n1695_));
  XOR2X1   g01439(.A(new_n1635_), .B(new_n1695_), .Y(new_n1696_));
  XOR2X1   g01440(.A(new_n1638_), .B(new_n1696_), .Y(new_n1697_));
  XOR2X1   g01441(.A(new_n1643_), .B(new_n1697_), .Y(new_n1698_));
  XOR2X1   g01442(.A(new_n1656_), .B(new_n1698_), .Y(new_n1699_));
  XOR2X1   g01443(.A(new_n1661_), .B(new_n1699_), .Y(new_n1700_));
  XOR2X1   g01444(.A(new_n1666_), .B(new_n1700_), .Y(new_n1701_));
  XOR2X1   g01445(.A(new_n1671_), .B(new_n1701_), .Y(new_n1702_));
  XOR2X1   g01446(.A(new_n1674_), .B(new_n1702_), .Y(new_n1703_));
  XOR2X1   g01447(.A(new_n1679_), .B(new_n1703_), .Y(new_n1704_));
  NOR2X1   g01448(.A(new_n1679_), .B(new_n1703_), .Y(new_n1705_));
  AOI21X1  g01449(.A0(new_n1704_), .A1(new_n1692_), .B0(new_n1705_), .Y(new_n1706_));
  OR2X1    g01450(.A(new_n1661_), .B(new_n1699_), .Y(new_n1707_));
  OAI21X1  g01451(.A0(new_n1666_), .A1(new_n1662_), .B0(new_n1707_), .Y(new_n1708_));
  OR2X1    g01452(.A(new_n1643_), .B(new_n1697_), .Y(new_n1709_));
  OAI21X1  g01453(.A0(new_n1656_), .A1(new_n1644_), .B0(new_n1709_), .Y(new_n1710_));
  OR2X1    g01454(.A(new_n1635_), .B(new_n1695_), .Y(new_n1711_));
  OAI21X1  g01455(.A0(new_n1638_), .A1(new_n1636_), .B0(new_n1711_), .Y(new_n1712_));
  AOI22X1  g01456(.A0(new_n1017_), .A1(\b[11] ), .B0(new_n1016_), .B1(\b[10] ), .Y(new_n1713_));
  OAI21X1  g01457(.A0(new_n1015_), .A1(new_n590_), .B0(new_n1713_), .Y(new_n1714_));
  AOI21X1  g01458(.A0(new_n882_), .A1(new_n589_), .B0(new_n1714_), .Y(new_n1715_));
  XOR2X1   g01459(.A(new_n1715_), .B(new_n879_), .Y(new_n1716_));
  NAND2X1  g01460(.A(new_n1629_), .B(new_n1607_), .Y(new_n1717_));
  NAND2X1  g01461(.A(new_n1630_), .B(new_n1603_), .Y(new_n1718_));
  AND2X1   g01462(.A(new_n1718_), .B(new_n1717_), .Y(new_n1719_));
  AND2X1   g01463(.A(new_n1627_), .B(new_n1614_), .Y(new_n1720_));
  AOI21X1  g01464(.A0(new_n1628_), .A1(new_n1609_), .B0(new_n1720_), .Y(new_n1721_));
  NOR2X1   g01465(.A(new_n1626_), .B(new_n1615_), .Y(new_n1722_));
  INVX1    g01466(.A(new_n1617_), .Y(new_n1723_));
  OR2X1    g01467(.A(new_n1619_), .B(new_n1520_), .Y(new_n1724_));
  NOR2X1   g01468(.A(new_n1724_), .B(new_n1622_), .Y(new_n1725_));
  OAI22X1  g01469(.A0(new_n1623_), .A1(new_n277_), .B0(new_n1620_), .B1(new_n275_), .Y(new_n1726_));
  AOI21X1  g01470(.A0(new_n1725_), .A1(\b[0] ), .B0(new_n1726_), .Y(new_n1727_));
  OAI21X1  g01471(.A0(new_n1723_), .A1(new_n281_), .B0(new_n1727_), .Y(new_n1728_));
  XOR2X1   g01472(.A(new_n1728_), .B(new_n1621_), .Y(new_n1729_));
  XOR2X1   g01473(.A(new_n1729_), .B(new_n1722_), .Y(new_n1730_));
  AOI22X1  g01474(.A0(new_n1526_), .A1(\b[5] ), .B0(new_n1525_), .B1(\b[4] ), .Y(new_n1731_));
  OAI21X1  g01475(.A0(new_n1524_), .A1(new_n297_), .B0(new_n1731_), .Y(new_n1732_));
  AOI21X1  g01476(.A0(new_n1347_), .A1(new_n349_), .B0(new_n1732_), .Y(new_n1733_));
  XOR2X1   g01477(.A(new_n1733_), .B(\a[23] ), .Y(new_n1734_));
  AND2X1   g01478(.A(new_n1734_), .B(new_n1730_), .Y(new_n1735_));
  XOR2X1   g01479(.A(new_n1734_), .B(new_n1730_), .Y(new_n1736_));
  OR2X1    g01480(.A(new_n1734_), .B(new_n1730_), .Y(new_n1737_));
  OAI21X1  g01481(.A0(new_n1735_), .A1(new_n1721_), .B0(new_n1737_), .Y(new_n1738_));
  OAI22X1  g01482(.A0(new_n1738_), .A1(new_n1735_), .B0(new_n1736_), .B1(new_n1721_), .Y(new_n1739_));
  AOI22X1  g01483(.A0(new_n1263_), .A1(\b[8] ), .B0(new_n1262_), .B1(\b[7] ), .Y(new_n1740_));
  OAI21X1  g01484(.A0(new_n1261_), .A1(new_n392_), .B0(new_n1740_), .Y(new_n1741_));
  AOI21X1  g01485(.A0(new_n1075_), .A1(new_n454_), .B0(new_n1741_), .Y(new_n1742_));
  XOR2X1   g01486(.A(new_n1742_), .B(\a[20] ), .Y(new_n1743_));
  XOR2X1   g01487(.A(new_n1743_), .B(new_n1739_), .Y(new_n1744_));
  XOR2X1   g01488(.A(new_n1744_), .B(new_n1719_), .Y(new_n1745_));
  XOR2X1   g01489(.A(new_n1745_), .B(new_n1716_), .Y(new_n1746_));
  XOR2X1   g01490(.A(new_n1746_), .B(new_n1712_), .Y(new_n1747_));
  AOI22X1  g01491(.A0(new_n818_), .A1(\b[14] ), .B0(new_n817_), .B1(\b[13] ), .Y(new_n1748_));
  OAI21X1  g01492(.A0(new_n816_), .A1(new_n713_), .B0(new_n1748_), .Y(new_n1749_));
  AOI21X1  g01493(.A0(new_n734_), .A1(new_n668_), .B0(new_n1749_), .Y(new_n1750_));
  XOR2X1   g01494(.A(new_n1750_), .B(\a[14] ), .Y(new_n1751_));
  XOR2X1   g01495(.A(new_n1751_), .B(new_n1747_), .Y(new_n1752_));
  XOR2X1   g01496(.A(new_n1752_), .B(new_n1710_), .Y(new_n1753_));
  AOI22X1  g01497(.A0(new_n603_), .A1(\b[17] ), .B0(new_n602_), .B1(\b[16] ), .Y(new_n1754_));
  OAI21X1  g01498(.A0(new_n601_), .A1(new_n977_), .B0(new_n1754_), .Y(new_n1755_));
  AOI21X1  g01499(.A0(new_n976_), .A1(new_n518_), .B0(new_n1755_), .Y(new_n1756_));
  XOR2X1   g01500(.A(new_n1756_), .B(\a[11] ), .Y(new_n1757_));
  XOR2X1   g01501(.A(new_n1757_), .B(new_n1753_), .Y(new_n1758_));
  XOR2X1   g01502(.A(new_n1758_), .B(new_n1708_), .Y(new_n1759_));
  AOI22X1  g01503(.A0(new_n469_), .A1(\b[20] ), .B0(new_n468_), .B1(\b[19] ), .Y(new_n1760_));
  OAI21X1  g01504(.A0(new_n467_), .A1(new_n1115_), .B0(new_n1760_), .Y(new_n1761_));
  AOI21X1  g01505(.A0(new_n1217_), .A1(new_n404_), .B0(new_n1761_), .Y(new_n1762_));
  XOR2X1   g01506(.A(new_n1762_), .B(\a[8] ), .Y(new_n1763_));
  XOR2X1   g01507(.A(new_n1763_), .B(new_n1759_), .Y(new_n1764_));
  NOR2X1   g01508(.A(new_n1671_), .B(new_n1701_), .Y(new_n1765_));
  AND2X1   g01509(.A(new_n1461_), .B(new_n1506_), .Y(new_n1766_));
  XOR2X1   g01510(.A(new_n1461_), .B(new_n1506_), .Y(new_n1767_));
  AOI21X1  g01511(.A0(new_n1767_), .A1(new_n1408_), .B0(new_n1766_), .Y(new_n1768_));
  AND2X1   g01512(.A(new_n1564_), .B(new_n1560_), .Y(new_n1769_));
  OR2X1    g01513(.A(new_n1564_), .B(new_n1560_), .Y(new_n1770_));
  OAI21X1  g01514(.A0(new_n1769_), .A1(new_n1768_), .B0(new_n1770_), .Y(new_n1771_));
  AOI21X1  g01515(.A0(new_n1771_), .A1(new_n1702_), .B0(new_n1765_), .Y(new_n1772_));
  XOR2X1   g01516(.A(new_n1772_), .B(new_n1764_), .Y(new_n1773_));
  AOI22X1  g01517(.A0(new_n369_), .A1(\b[23] ), .B0(new_n368_), .B1(\b[22] ), .Y(new_n1774_));
  OAI21X1  g01518(.A0(new_n367_), .A1(new_n1482_), .B0(new_n1774_), .Y(new_n1775_));
  AOI21X1  g01519(.A0(new_n1481_), .A1(new_n308_), .B0(new_n1775_), .Y(new_n1776_));
  XOR2X1   g01520(.A(new_n1776_), .B(\a[5] ), .Y(new_n1777_));
  XOR2X1   g01521(.A(new_n1777_), .B(new_n1773_), .Y(new_n1778_));
  XOR2X1   g01522(.A(new_n1778_), .B(new_n1706_), .Y(new_n1779_));
  NAND2X1  g01523(.A(\b[25] ), .B(\b[24] ), .Y(new_n1780_));
  OAI21X1  g01524(.A0(new_n1589_), .A1(new_n1587_), .B0(new_n1780_), .Y(new_n1781_));
  XOR2X1   g01525(.A(\b[26] ), .B(\b[25] ), .Y(new_n1782_));
  XOR2X1   g01526(.A(new_n1782_), .B(new_n1781_), .Y(new_n1783_));
  AOI22X1  g01527(.A0(new_n267_), .A1(\b[26] ), .B0(new_n266_), .B1(\b[25] ), .Y(new_n1784_));
  OAI21X1  g01528(.A0(new_n350_), .A1(new_n1588_), .B0(new_n1784_), .Y(new_n1785_));
  AOI21X1  g01529(.A0(new_n1783_), .A1(new_n318_), .B0(new_n1785_), .Y(new_n1786_));
  XOR2X1   g01530(.A(new_n1786_), .B(\a[2] ), .Y(new_n1787_));
  XOR2X1   g01531(.A(new_n1787_), .B(new_n1779_), .Y(new_n1788_));
  XOR2X1   g01532(.A(new_n1788_), .B(new_n1686_), .Y(\f[26] ));
  OR2X1    g01533(.A(new_n1679_), .B(new_n1703_), .Y(new_n1790_));
  OAI21X1  g01534(.A0(new_n1680_), .A1(new_n1599_), .B0(new_n1790_), .Y(new_n1791_));
  XOR2X1   g01535(.A(new_n1778_), .B(new_n1791_), .Y(new_n1792_));
  NOR2X1   g01536(.A(new_n1787_), .B(new_n1792_), .Y(new_n1793_));
  AOI21X1  g01537(.A0(new_n1685_), .A1(new_n1684_), .B0(new_n1788_), .Y(new_n1794_));
  OR2X1    g01538(.A(new_n1794_), .B(new_n1793_), .Y(new_n1795_));
  AND2X1   g01539(.A(new_n1745_), .B(new_n1716_), .Y(new_n1796_));
  AOI21X1  g01540(.A0(new_n1746_), .A1(new_n1712_), .B0(new_n1796_), .Y(new_n1797_));
  AOI22X1  g01541(.A0(new_n1017_), .A1(\b[12] ), .B0(new_n1016_), .B1(\b[11] ), .Y(new_n1798_));
  OAI21X1  g01542(.A0(new_n1015_), .A1(new_n587_), .B0(new_n1798_), .Y(new_n1799_));
  AOI21X1  g01543(.A0(new_n882_), .A1(new_n635_), .B0(new_n1799_), .Y(new_n1800_));
  XOR2X1   g01544(.A(new_n1800_), .B(new_n879_), .Y(new_n1801_));
  OR2X1    g01545(.A(new_n1736_), .B(new_n1721_), .Y(new_n1802_));
  INVX1    g01546(.A(new_n1735_), .Y(new_n1803_));
  NAND3X1  g01547(.A(new_n1803_), .B(new_n1737_), .C(new_n1721_), .Y(new_n1804_));
  AOI21X1  g01548(.A0(new_n1804_), .A1(new_n1802_), .B0(new_n1743_), .Y(new_n1805_));
  AOI21X1  g01549(.A0(new_n1718_), .A1(new_n1717_), .B0(new_n1744_), .Y(new_n1806_));
  OR2X1    g01550(.A(new_n1806_), .B(new_n1805_), .Y(new_n1807_));
  OR4X1    g01551(.A(new_n1728_), .B(new_n1626_), .C(new_n1522_), .D(new_n1621_), .Y(new_n1808_));
  XOR2X1   g01552(.A(\a[27] ), .B(\a[26] ), .Y(new_n1809_));
  NAND2X1  g01553(.A(new_n1809_), .B(\b[0] ), .Y(new_n1810_));
  XOR2X1   g01554(.A(new_n1810_), .B(new_n1808_), .Y(new_n1811_));
  INVX1    g01555(.A(new_n1725_), .Y(new_n1812_));
  AND2X1   g01556(.A(new_n1619_), .B(new_n1618_), .Y(new_n1813_));
  AND2X1   g01557(.A(new_n1622_), .B(new_n1520_), .Y(new_n1814_));
  AOI22X1  g01558(.A0(new_n1814_), .A1(\b[3] ), .B0(new_n1813_), .B1(\b[2] ), .Y(new_n1815_));
  OAI21X1  g01559(.A0(new_n1812_), .A1(new_n275_), .B0(new_n1815_), .Y(new_n1816_));
  AOI21X1  g01560(.A0(new_n1617_), .A1(new_n366_), .B0(new_n1816_), .Y(new_n1817_));
  XOR2X1   g01561(.A(new_n1817_), .B(\a[26] ), .Y(new_n1818_));
  XOR2X1   g01562(.A(new_n1818_), .B(new_n1811_), .Y(new_n1819_));
  AOI22X1  g01563(.A0(new_n1526_), .A1(\b[6] ), .B0(new_n1525_), .B1(\b[5] ), .Y(new_n1820_));
  OAI21X1  g01564(.A0(new_n1524_), .A1(new_n325_), .B0(new_n1820_), .Y(new_n1821_));
  AOI21X1  g01565(.A0(new_n1347_), .A1(new_n378_), .B0(new_n1821_), .Y(new_n1822_));
  XOR2X1   g01566(.A(new_n1822_), .B(\a[23] ), .Y(new_n1823_));
  XOR2X1   g01567(.A(new_n1823_), .B(new_n1819_), .Y(new_n1824_));
  INVX1    g01568(.A(new_n1824_), .Y(new_n1825_));
  XOR2X1   g01569(.A(new_n1825_), .B(new_n1738_), .Y(new_n1826_));
  AOI22X1  g01570(.A0(new_n1263_), .A1(\b[9] ), .B0(new_n1262_), .B1(\b[8] ), .Y(new_n1827_));
  OAI21X1  g01571(.A0(new_n1261_), .A1(new_n492_), .B0(new_n1827_), .Y(new_n1828_));
  AOI21X1  g01572(.A0(new_n1075_), .A1(new_n491_), .B0(new_n1828_), .Y(new_n1829_));
  XOR2X1   g01573(.A(new_n1829_), .B(\a[20] ), .Y(new_n1830_));
  XOR2X1   g01574(.A(new_n1830_), .B(new_n1826_), .Y(new_n1831_));
  XOR2X1   g01575(.A(new_n1831_), .B(new_n1807_), .Y(new_n1832_));
  XOR2X1   g01576(.A(new_n1832_), .B(new_n1801_), .Y(new_n1833_));
  XOR2X1   g01577(.A(new_n1833_), .B(new_n1797_), .Y(new_n1834_));
  AOI22X1  g01578(.A0(new_n818_), .A1(\b[15] ), .B0(new_n817_), .B1(\b[14] ), .Y(new_n1835_));
  OAI21X1  g01579(.A0(new_n816_), .A1(new_n795_), .B0(new_n1835_), .Y(new_n1836_));
  AOI21X1  g01580(.A0(new_n794_), .A1(new_n668_), .B0(new_n1836_), .Y(new_n1837_));
  XOR2X1   g01581(.A(new_n1837_), .B(\a[14] ), .Y(new_n1838_));
  XOR2X1   g01582(.A(new_n1838_), .B(new_n1834_), .Y(new_n1839_));
  INVX1    g01583(.A(new_n1751_), .Y(new_n1840_));
  AND2X1   g01584(.A(new_n1840_), .B(new_n1747_), .Y(new_n1841_));
  XOR2X1   g01585(.A(new_n1840_), .B(new_n1747_), .Y(new_n1842_));
  AOI21X1  g01586(.A0(new_n1842_), .A1(new_n1710_), .B0(new_n1841_), .Y(new_n1843_));
  XOR2X1   g01587(.A(new_n1843_), .B(new_n1839_), .Y(new_n1844_));
  AOI22X1  g01588(.A0(new_n603_), .A1(\b[18] ), .B0(new_n602_), .B1(\b[17] ), .Y(new_n1845_));
  OAI21X1  g01589(.A0(new_n601_), .A1(new_n974_), .B0(new_n1845_), .Y(new_n1846_));
  AOI21X1  g01590(.A0(new_n1042_), .A1(new_n518_), .B0(new_n1846_), .Y(new_n1847_));
  XOR2X1   g01591(.A(new_n1847_), .B(\a[11] ), .Y(new_n1848_));
  XOR2X1   g01592(.A(new_n1848_), .B(new_n1844_), .Y(new_n1849_));
  NOR2X1   g01593(.A(new_n1757_), .B(new_n1753_), .Y(new_n1850_));
  AOI21X1  g01594(.A0(new_n1758_), .A1(new_n1708_), .B0(new_n1850_), .Y(new_n1851_));
  XOR2X1   g01595(.A(new_n1851_), .B(new_n1849_), .Y(new_n1852_));
  AOI22X1  g01596(.A0(new_n469_), .A1(\b[21] ), .B0(new_n468_), .B1(\b[20] ), .Y(new_n1853_));
  OAI21X1  g01597(.A0(new_n467_), .A1(new_n1300_), .B0(new_n1853_), .Y(new_n1854_));
  AOI21X1  g01598(.A0(new_n1299_), .A1(new_n404_), .B0(new_n1854_), .Y(new_n1855_));
  XOR2X1   g01599(.A(new_n1855_), .B(\a[8] ), .Y(new_n1856_));
  XOR2X1   g01600(.A(new_n1856_), .B(new_n1852_), .Y(new_n1857_));
  INVX1    g01601(.A(new_n1763_), .Y(new_n1858_));
  AND2X1   g01602(.A(new_n1858_), .B(new_n1759_), .Y(new_n1859_));
  XOR2X1   g01603(.A(new_n1858_), .B(new_n1759_), .Y(new_n1860_));
  OR2X1    g01604(.A(new_n1671_), .B(new_n1701_), .Y(new_n1861_));
  OAI21X1  g01605(.A0(new_n1674_), .A1(new_n1672_), .B0(new_n1861_), .Y(new_n1862_));
  AOI21X1  g01606(.A0(new_n1862_), .A1(new_n1860_), .B0(new_n1859_), .Y(new_n1863_));
  XOR2X1   g01607(.A(new_n1863_), .B(new_n1857_), .Y(new_n1864_));
  AOI22X1  g01608(.A0(new_n369_), .A1(\b[24] ), .B0(new_n368_), .B1(\b[23] ), .Y(new_n1865_));
  OAI21X1  g01609(.A0(new_n367_), .A1(new_n1479_), .B0(new_n1865_), .Y(new_n1866_));
  AOI21X1  g01610(.A0(new_n1572_), .A1(new_n308_), .B0(new_n1866_), .Y(new_n1867_));
  XOR2X1   g01611(.A(new_n1867_), .B(\a[5] ), .Y(new_n1868_));
  XOR2X1   g01612(.A(new_n1868_), .B(new_n1864_), .Y(new_n1869_));
  XOR2X1   g01613(.A(new_n1772_), .B(new_n1860_), .Y(new_n1870_));
  NOR2X1   g01614(.A(new_n1777_), .B(new_n1870_), .Y(new_n1871_));
  XOR2X1   g01615(.A(new_n1777_), .B(new_n1870_), .Y(new_n1872_));
  AOI21X1  g01616(.A0(new_n1872_), .A1(new_n1791_), .B0(new_n1871_), .Y(new_n1873_));
  XOR2X1   g01617(.A(new_n1873_), .B(new_n1869_), .Y(new_n1874_));
  AND2X1   g01618(.A(\b[26] ), .B(\b[25] ), .Y(new_n1875_));
  AOI21X1  g01619(.A0(new_n1782_), .A1(new_n1781_), .B0(new_n1875_), .Y(new_n1876_));
  INVX1    g01620(.A(\b[26] ), .Y(new_n1877_));
  XOR2X1   g01621(.A(\b[27] ), .B(new_n1877_), .Y(new_n1878_));
  XOR2X1   g01622(.A(new_n1878_), .B(new_n1876_), .Y(new_n1879_));
  INVX1    g01623(.A(\b[25] ), .Y(new_n1880_));
  AOI22X1  g01624(.A0(new_n267_), .A1(\b[27] ), .B0(new_n266_), .B1(\b[26] ), .Y(new_n1881_));
  OAI21X1  g01625(.A0(new_n350_), .A1(new_n1880_), .B0(new_n1881_), .Y(new_n1882_));
  AOI21X1  g01626(.A0(new_n1879_), .A1(new_n318_), .B0(new_n1882_), .Y(new_n1883_));
  XOR2X1   g01627(.A(new_n1883_), .B(\a[2] ), .Y(new_n1884_));
  XOR2X1   g01628(.A(new_n1884_), .B(new_n1874_), .Y(new_n1885_));
  XOR2X1   g01629(.A(new_n1885_), .B(new_n1795_), .Y(\f[27] ));
  OR2X1    g01630(.A(new_n1884_), .B(new_n1874_), .Y(new_n1887_));
  OAI21X1  g01631(.A0(new_n1794_), .A1(new_n1793_), .B0(new_n1885_), .Y(new_n1888_));
  AND2X1   g01632(.A(new_n1888_), .B(new_n1887_), .Y(new_n1889_));
  NOR2X1   g01633(.A(new_n1823_), .B(new_n1819_), .Y(new_n1890_));
  AOI21X1  g01634(.A0(new_n1824_), .A1(new_n1738_), .B0(new_n1890_), .Y(new_n1891_));
  AOI22X1  g01635(.A0(new_n1526_), .A1(\b[7] ), .B0(new_n1525_), .B1(\b[6] ), .Y(new_n1892_));
  OAI21X1  g01636(.A0(new_n1524_), .A1(new_n395_), .B0(new_n1892_), .Y(new_n1893_));
  AOI21X1  g01637(.A0(new_n1347_), .A1(new_n394_), .B0(new_n1893_), .Y(new_n1894_));
  XOR2X1   g01638(.A(new_n1894_), .B(\a[23] ), .Y(new_n1895_));
  INVX1    g01639(.A(new_n1810_), .Y(new_n1896_));
  XOR2X1   g01640(.A(new_n1896_), .B(new_n1808_), .Y(new_n1897_));
  OR2X1    g01641(.A(new_n1810_), .B(new_n1808_), .Y(new_n1898_));
  OAI21X1  g01642(.A0(new_n1818_), .A1(new_n1897_), .B0(new_n1898_), .Y(new_n1899_));
  AND2X1   g01643(.A(new_n1617_), .B(new_n323_), .Y(new_n1900_));
  NOR3X1   g01644(.A(new_n1724_), .B(new_n1622_), .C(new_n277_), .Y(new_n1901_));
  OAI22X1  g01645(.A0(new_n1623_), .A1(new_n325_), .B0(new_n1620_), .B1(new_n297_), .Y(new_n1902_));
  NOR3X1   g01646(.A(new_n1902_), .B(new_n1901_), .C(new_n1900_), .Y(new_n1903_));
  XOR2X1   g01647(.A(new_n1903_), .B(new_n1621_), .Y(new_n1904_));
  NAND2X1  g01648(.A(new_n1810_), .B(\a[29] ), .Y(new_n1905_));
  XOR2X1   g01649(.A(\a[29] ), .B(\a[28] ), .Y(new_n1906_));
  AND2X1   g01650(.A(new_n1906_), .B(new_n1809_), .Y(new_n1907_));
  XOR2X1   g01651(.A(\a[27] ), .B(new_n1621_), .Y(new_n1908_));
  XOR2X1   g01652(.A(\a[28] ), .B(\a[27] ), .Y(new_n1909_));
  NAND2X1  g01653(.A(new_n1909_), .B(new_n1908_), .Y(new_n1910_));
  INVX1    g01654(.A(\a[29] ), .Y(new_n1911_));
  XOR2X1   g01655(.A(new_n1911_), .B(\a[28] ), .Y(new_n1912_));
  NAND2X1  g01656(.A(new_n1912_), .B(new_n1809_), .Y(new_n1913_));
  OAI22X1  g01657(.A0(new_n1913_), .A1(new_n275_), .B0(new_n1910_), .B1(new_n274_), .Y(new_n1914_));
  AOI21X1  g01658(.A0(new_n1907_), .A1(new_n263_), .B0(new_n1914_), .Y(new_n1915_));
  XOR2X1   g01659(.A(new_n1915_), .B(\a[29] ), .Y(new_n1916_));
  XOR2X1   g01660(.A(new_n1916_), .B(new_n1905_), .Y(new_n1917_));
  XOR2X1   g01661(.A(new_n1917_), .B(new_n1904_), .Y(new_n1918_));
  XOR2X1   g01662(.A(new_n1918_), .B(new_n1899_), .Y(new_n1919_));
  XOR2X1   g01663(.A(new_n1919_), .B(new_n1895_), .Y(new_n1920_));
  XOR2X1   g01664(.A(new_n1920_), .B(new_n1891_), .Y(new_n1921_));
  AOI22X1  g01665(.A0(new_n1263_), .A1(\b[10] ), .B0(new_n1262_), .B1(\b[9] ), .Y(new_n1922_));
  OAI21X1  g01666(.A0(new_n1261_), .A1(new_n489_), .B0(new_n1922_), .Y(new_n1923_));
  AOI21X1  g01667(.A0(new_n1075_), .A1(new_n543_), .B0(new_n1923_), .Y(new_n1924_));
  XOR2X1   g01668(.A(new_n1924_), .B(\a[20] ), .Y(new_n1925_));
  XOR2X1   g01669(.A(new_n1925_), .B(new_n1921_), .Y(new_n1926_));
  OR2X1    g01670(.A(new_n1830_), .B(new_n1826_), .Y(new_n1927_));
  OAI21X1  g01671(.A0(new_n1806_), .A1(new_n1805_), .B0(new_n1831_), .Y(new_n1928_));
  AND2X1   g01672(.A(new_n1928_), .B(new_n1927_), .Y(new_n1929_));
  XOR2X1   g01673(.A(new_n1929_), .B(new_n1926_), .Y(new_n1930_));
  AOI22X1  g01674(.A0(new_n1017_), .A1(\b[13] ), .B0(new_n1016_), .B1(\b[12] ), .Y(new_n1931_));
  OAI21X1  g01675(.A0(new_n1015_), .A1(new_n716_), .B0(new_n1931_), .Y(new_n1932_));
  AOI21X1  g01676(.A0(new_n882_), .A1(new_n715_), .B0(new_n1932_), .Y(new_n1933_));
  XOR2X1   g01677(.A(new_n1933_), .B(\a[17] ), .Y(new_n1934_));
  XOR2X1   g01678(.A(new_n1934_), .B(new_n1930_), .Y(new_n1935_));
  NOR3X1   g01679(.A(new_n1635_), .B(new_n1694_), .C(new_n1693_), .Y(new_n1936_));
  NOR2X1   g01680(.A(new_n1449_), .B(new_n1445_), .Y(new_n1937_));
  AOI21X1  g01681(.A0(new_n1450_), .A1(new_n1423_), .B0(new_n1937_), .Y(new_n1938_));
  OR2X1    g01682(.A(new_n1541_), .B(new_n1537_), .Y(new_n1939_));
  AND2X1   g01683(.A(new_n1541_), .B(new_n1537_), .Y(new_n1940_));
  OAI21X1  g01684(.A0(new_n1940_), .A1(new_n1938_), .B0(new_n1939_), .Y(new_n1941_));
  AOI21X1  g01685(.A0(new_n1941_), .A1(new_n1696_), .B0(new_n1936_), .Y(new_n1942_));
  NOR2X1   g01686(.A(new_n1745_), .B(new_n1716_), .Y(new_n1943_));
  NAND2X1  g01687(.A(new_n1745_), .B(new_n1716_), .Y(new_n1944_));
  OAI21X1  g01688(.A0(new_n1943_), .A1(new_n1942_), .B0(new_n1944_), .Y(new_n1945_));
  AND2X1   g01689(.A(new_n1832_), .B(new_n1801_), .Y(new_n1946_));
  AOI21X1  g01690(.A0(new_n1833_), .A1(new_n1945_), .B0(new_n1946_), .Y(new_n1947_));
  XOR2X1   g01691(.A(new_n1947_), .B(new_n1935_), .Y(new_n1948_));
  AOI22X1  g01692(.A0(new_n818_), .A1(\b[16] ), .B0(new_n817_), .B1(\b[15] ), .Y(new_n1949_));
  OAI21X1  g01693(.A0(new_n816_), .A1(new_n792_), .B0(new_n1949_), .Y(new_n1950_));
  AOI21X1  g01694(.A0(new_n842_), .A1(new_n668_), .B0(new_n1950_), .Y(new_n1951_));
  XOR2X1   g01695(.A(new_n1951_), .B(\a[14] ), .Y(new_n1952_));
  XOR2X1   g01696(.A(new_n1952_), .B(new_n1948_), .Y(new_n1953_));
  NOR2X1   g01697(.A(new_n1838_), .B(new_n1834_), .Y(new_n1954_));
  NOR2X1   g01698(.A(new_n1643_), .B(new_n1697_), .Y(new_n1955_));
  NOR2X1   g01699(.A(new_n1543_), .B(new_n1514_), .Y(new_n1956_));
  NAND2X1  g01700(.A(new_n1543_), .B(new_n1514_), .Y(new_n1957_));
  OAI21X1  g01701(.A0(new_n1956_), .A1(new_n1510_), .B0(new_n1957_), .Y(new_n1958_));
  AOI21X1  g01702(.A0(new_n1958_), .A1(new_n1698_), .B0(new_n1955_), .Y(new_n1959_));
  NAND2X1  g01703(.A(new_n1840_), .B(new_n1747_), .Y(new_n1960_));
  OAI21X1  g01704(.A0(new_n1752_), .A1(new_n1959_), .B0(new_n1960_), .Y(new_n1961_));
  AOI21X1  g01705(.A0(new_n1961_), .A1(new_n1839_), .B0(new_n1954_), .Y(new_n1962_));
  XOR2X1   g01706(.A(new_n1962_), .B(new_n1953_), .Y(new_n1963_));
  AOI22X1  g01707(.A0(new_n603_), .A1(\b[19] ), .B0(new_n602_), .B1(\b[18] ), .Y(new_n1964_));
  OAI21X1  g01708(.A0(new_n601_), .A1(new_n1118_), .B0(new_n1964_), .Y(new_n1965_));
  AOI21X1  g01709(.A0(new_n1117_), .A1(new_n518_), .B0(new_n1965_), .Y(new_n1966_));
  XOR2X1   g01710(.A(new_n1966_), .B(\a[11] ), .Y(new_n1967_));
  XOR2X1   g01711(.A(new_n1967_), .B(new_n1963_), .Y(new_n1968_));
  NOR2X1   g01712(.A(new_n1848_), .B(new_n1844_), .Y(new_n1969_));
  NOR2X1   g01713(.A(new_n1661_), .B(new_n1699_), .Y(new_n1970_));
  OR2X1    g01714(.A(new_n1549_), .B(new_n1545_), .Y(new_n1971_));
  INVX1    g01715(.A(new_n1549_), .Y(new_n1972_));
  XOR2X1   g01716(.A(new_n1972_), .B(new_n1545_), .Y(new_n1973_));
  OAI21X1  g01717(.A0(new_n1559_), .A1(new_n1973_), .B0(new_n1971_), .Y(new_n1974_));
  AOI21X1  g01718(.A0(new_n1974_), .A1(new_n1700_), .B0(new_n1970_), .Y(new_n1975_));
  OR2X1    g01719(.A(new_n1757_), .B(new_n1753_), .Y(new_n1976_));
  AND2X1   g01720(.A(new_n1757_), .B(new_n1753_), .Y(new_n1977_));
  OAI21X1  g01721(.A0(new_n1977_), .A1(new_n1975_), .B0(new_n1976_), .Y(new_n1978_));
  AOI21X1  g01722(.A0(new_n1978_), .A1(new_n1849_), .B0(new_n1969_), .Y(new_n1979_));
  XOR2X1   g01723(.A(new_n1979_), .B(new_n1968_), .Y(new_n1980_));
  AOI22X1  g01724(.A0(new_n469_), .A1(\b[22] ), .B0(new_n468_), .B1(\b[21] ), .Y(new_n1981_));
  OAI21X1  g01725(.A0(new_n467_), .A1(new_n1297_), .B0(new_n1981_), .Y(new_n1982_));
  AOI21X1  g01726(.A0(new_n1399_), .A1(new_n404_), .B0(new_n1982_), .Y(new_n1983_));
  XOR2X1   g01727(.A(new_n1983_), .B(\a[8] ), .Y(new_n1984_));
  XOR2X1   g01728(.A(new_n1984_), .B(new_n1980_), .Y(new_n1985_));
  NOR2X1   g01729(.A(new_n1856_), .B(new_n1852_), .Y(new_n1986_));
  NAND2X1  g01730(.A(new_n1858_), .B(new_n1759_), .Y(new_n1987_));
  OAI21X1  g01731(.A0(new_n1772_), .A1(new_n1764_), .B0(new_n1987_), .Y(new_n1988_));
  AOI21X1  g01732(.A0(new_n1988_), .A1(new_n1857_), .B0(new_n1986_), .Y(new_n1989_));
  XOR2X1   g01733(.A(new_n1989_), .B(new_n1985_), .Y(new_n1990_));
  AOI22X1  g01734(.A0(new_n369_), .A1(\b[25] ), .B0(new_n368_), .B1(\b[24] ), .Y(new_n1991_));
  OAI21X1  g01735(.A0(new_n367_), .A1(new_n1591_), .B0(new_n1991_), .Y(new_n1992_));
  AOI21X1  g01736(.A0(new_n1590_), .A1(new_n308_), .B0(new_n1992_), .Y(new_n1993_));
  XOR2X1   g01737(.A(new_n1993_), .B(\a[5] ), .Y(new_n1994_));
  XOR2X1   g01738(.A(new_n1994_), .B(new_n1990_), .Y(new_n1995_));
  NOR2X1   g01739(.A(new_n1868_), .B(new_n1864_), .Y(new_n1996_));
  OR2X1    g01740(.A(new_n1777_), .B(new_n1870_), .Y(new_n1997_));
  OAI21X1  g01741(.A0(new_n1778_), .A1(new_n1706_), .B0(new_n1997_), .Y(new_n1998_));
  AOI21X1  g01742(.A0(new_n1998_), .A1(new_n1869_), .B0(new_n1996_), .Y(new_n1999_));
  XOR2X1   g01743(.A(new_n1999_), .B(new_n1995_), .Y(new_n2000_));
  NAND2X1  g01744(.A(\b[27] ), .B(\b[26] ), .Y(new_n2001_));
  OAI21X1  g01745(.A0(new_n1878_), .A1(new_n1876_), .B0(new_n2001_), .Y(new_n2002_));
  XOR2X1   g01746(.A(\b[28] ), .B(\b[27] ), .Y(new_n2003_));
  XOR2X1   g01747(.A(new_n2003_), .B(new_n2002_), .Y(new_n2004_));
  AOI22X1  g01748(.A0(new_n267_), .A1(\b[28] ), .B0(new_n266_), .B1(\b[27] ), .Y(new_n2005_));
  OAI21X1  g01749(.A0(new_n350_), .A1(new_n1877_), .B0(new_n2005_), .Y(new_n2006_));
  AOI21X1  g01750(.A0(new_n2004_), .A1(new_n318_), .B0(new_n2006_), .Y(new_n2007_));
  XOR2X1   g01751(.A(new_n2007_), .B(\a[2] ), .Y(new_n2008_));
  XOR2X1   g01752(.A(new_n2008_), .B(new_n2000_), .Y(new_n2009_));
  XOR2X1   g01753(.A(new_n2009_), .B(new_n1889_), .Y(\f[28] ));
  INVX1    g01754(.A(new_n1926_), .Y(new_n2011_));
  XOR2X1   g01755(.A(new_n1929_), .B(new_n2011_), .Y(new_n2012_));
  XOR2X1   g01756(.A(new_n1934_), .B(new_n2012_), .Y(new_n2013_));
  XOR2X1   g01757(.A(new_n1947_), .B(new_n2013_), .Y(new_n2014_));
  XOR2X1   g01758(.A(new_n1952_), .B(new_n2014_), .Y(new_n2015_));
  XOR2X1   g01759(.A(new_n1962_), .B(new_n2015_), .Y(new_n2016_));
  XOR2X1   g01760(.A(new_n1967_), .B(new_n2016_), .Y(new_n2017_));
  XOR2X1   g01761(.A(new_n1979_), .B(new_n2017_), .Y(new_n2018_));
  XOR2X1   g01762(.A(new_n1984_), .B(new_n2018_), .Y(new_n2019_));
  XOR2X1   g01763(.A(new_n1989_), .B(new_n2019_), .Y(new_n2020_));
  OR2X1    g01764(.A(new_n1994_), .B(new_n2020_), .Y(new_n2021_));
  OAI21X1  g01765(.A0(new_n1999_), .A1(new_n1995_), .B0(new_n2021_), .Y(new_n2022_));
  AOI22X1  g01766(.A0(new_n369_), .A1(\b[26] ), .B0(new_n368_), .B1(\b[25] ), .Y(new_n2023_));
  OAI21X1  g01767(.A0(new_n367_), .A1(new_n1588_), .B0(new_n2023_), .Y(new_n2024_));
  AOI21X1  g01768(.A0(new_n1783_), .A1(new_n308_), .B0(new_n2024_), .Y(new_n2025_));
  XOR2X1   g01769(.A(new_n2025_), .B(\a[5] ), .Y(new_n2026_));
  OR2X1    g01770(.A(new_n1967_), .B(new_n2016_), .Y(new_n2027_));
  OAI21X1  g01771(.A0(new_n1979_), .A1(new_n1968_), .B0(new_n2027_), .Y(new_n2028_));
  INVX1    g01772(.A(new_n1921_), .Y(new_n2029_));
  NOR2X1   g01773(.A(new_n1925_), .B(new_n2029_), .Y(new_n2030_));
  AOI21X1  g01774(.A0(new_n1928_), .A1(new_n1927_), .B0(new_n1926_), .Y(new_n2031_));
  OR2X1    g01775(.A(new_n2031_), .B(new_n2030_), .Y(new_n2032_));
  AOI22X1  g01776(.A0(new_n1263_), .A1(\b[11] ), .B0(new_n1262_), .B1(\b[10] ), .Y(new_n2033_));
  OAI21X1  g01777(.A0(new_n1261_), .A1(new_n590_), .B0(new_n2033_), .Y(new_n2034_));
  AOI21X1  g01778(.A0(new_n1075_), .A1(new_n589_), .B0(new_n2034_), .Y(new_n2035_));
  XOR2X1   g01779(.A(new_n2035_), .B(new_n1072_), .Y(new_n2036_));
  INVX1    g01780(.A(new_n1895_), .Y(new_n2037_));
  NAND2X1  g01781(.A(new_n1919_), .B(new_n2037_), .Y(new_n2038_));
  OAI21X1  g01782(.A0(new_n1920_), .A1(new_n1891_), .B0(new_n2038_), .Y(new_n2039_));
  AND2X1   g01783(.A(new_n1917_), .B(new_n1904_), .Y(new_n2040_));
  AOI21X1  g01784(.A0(new_n1918_), .A1(new_n1899_), .B0(new_n2040_), .Y(new_n2041_));
  NOR2X1   g01785(.A(new_n1916_), .B(new_n1905_), .Y(new_n2042_));
  INVX1    g01786(.A(new_n1907_), .Y(new_n2043_));
  OR2X1    g01787(.A(new_n1909_), .B(new_n1809_), .Y(new_n2044_));
  NOR2X1   g01788(.A(new_n2044_), .B(new_n1912_), .Y(new_n2045_));
  OAI22X1  g01789(.A0(new_n1913_), .A1(new_n277_), .B0(new_n1910_), .B1(new_n275_), .Y(new_n2046_));
  AOI21X1  g01790(.A0(new_n2045_), .A1(\b[0] ), .B0(new_n2046_), .Y(new_n2047_));
  OAI21X1  g01791(.A0(new_n2043_), .A1(new_n281_), .B0(new_n2047_), .Y(new_n2048_));
  XOR2X1   g01792(.A(new_n2048_), .B(new_n1911_), .Y(new_n2049_));
  XOR2X1   g01793(.A(new_n2049_), .B(new_n2042_), .Y(new_n2050_));
  AOI22X1  g01794(.A0(new_n1814_), .A1(\b[5] ), .B0(new_n1813_), .B1(\b[4] ), .Y(new_n2051_));
  OAI21X1  g01795(.A0(new_n1812_), .A1(new_n297_), .B0(new_n2051_), .Y(new_n2052_));
  AOI21X1  g01796(.A0(new_n1617_), .A1(new_n349_), .B0(new_n2052_), .Y(new_n2053_));
  XOR2X1   g01797(.A(new_n2053_), .B(\a[26] ), .Y(new_n2054_));
  XOR2X1   g01798(.A(new_n2054_), .B(new_n2050_), .Y(new_n2055_));
  OR2X1    g01799(.A(new_n2055_), .B(new_n2041_), .Y(new_n2056_));
  OR2X1    g01800(.A(new_n2054_), .B(new_n2050_), .Y(new_n2057_));
  AND2X1   g01801(.A(new_n2054_), .B(new_n2050_), .Y(new_n2058_));
  INVX1    g01802(.A(new_n2058_), .Y(new_n2059_));
  NAND3X1  g01803(.A(new_n2059_), .B(new_n2057_), .C(new_n2041_), .Y(new_n2060_));
  AND2X1   g01804(.A(new_n2060_), .B(new_n2056_), .Y(new_n2061_));
  AOI22X1  g01805(.A0(new_n1526_), .A1(\b[8] ), .B0(new_n1525_), .B1(\b[7] ), .Y(new_n2062_));
  OAI21X1  g01806(.A0(new_n1524_), .A1(new_n392_), .B0(new_n2062_), .Y(new_n2063_));
  AOI21X1  g01807(.A0(new_n1347_), .A1(new_n454_), .B0(new_n2063_), .Y(new_n2064_));
  XOR2X1   g01808(.A(new_n2064_), .B(\a[23] ), .Y(new_n2065_));
  XOR2X1   g01809(.A(new_n2065_), .B(new_n2061_), .Y(new_n2066_));
  XOR2X1   g01810(.A(new_n2066_), .B(new_n2039_), .Y(new_n2067_));
  XOR2X1   g01811(.A(new_n2067_), .B(new_n2036_), .Y(new_n2068_));
  XOR2X1   g01812(.A(new_n2068_), .B(new_n2032_), .Y(new_n2069_));
  AOI22X1  g01813(.A0(new_n1017_), .A1(\b[14] ), .B0(new_n1016_), .B1(\b[13] ), .Y(new_n2070_));
  OAI21X1  g01814(.A0(new_n1015_), .A1(new_n713_), .B0(new_n2070_), .Y(new_n2071_));
  AOI21X1  g01815(.A0(new_n882_), .A1(new_n734_), .B0(new_n2071_), .Y(new_n2072_));
  XOR2X1   g01816(.A(new_n2072_), .B(\a[17] ), .Y(new_n2073_));
  INVX1    g01817(.A(new_n2073_), .Y(new_n2074_));
  XOR2X1   g01818(.A(new_n2074_), .B(new_n2069_), .Y(new_n2075_));
  NOR2X1   g01819(.A(new_n1934_), .B(new_n2012_), .Y(new_n2076_));
  NOR2X1   g01820(.A(new_n1832_), .B(new_n1801_), .Y(new_n2077_));
  NAND2X1  g01821(.A(new_n1832_), .B(new_n1801_), .Y(new_n2078_));
  OAI21X1  g01822(.A0(new_n2077_), .A1(new_n1797_), .B0(new_n2078_), .Y(new_n2079_));
  AOI21X1  g01823(.A0(new_n2079_), .A1(new_n2013_), .B0(new_n2076_), .Y(new_n2080_));
  XOR2X1   g01824(.A(new_n2080_), .B(new_n2075_), .Y(new_n2081_));
  AOI22X1  g01825(.A0(new_n818_), .A1(\b[17] ), .B0(new_n817_), .B1(\b[16] ), .Y(new_n2082_));
  OAI21X1  g01826(.A0(new_n816_), .A1(new_n977_), .B0(new_n2082_), .Y(new_n2083_));
  AOI21X1  g01827(.A0(new_n976_), .A1(new_n668_), .B0(new_n2083_), .Y(new_n2084_));
  XOR2X1   g01828(.A(new_n2084_), .B(\a[14] ), .Y(new_n2085_));
  XOR2X1   g01829(.A(new_n2085_), .B(new_n2081_), .Y(new_n2086_));
  NOR2X1   g01830(.A(new_n1952_), .B(new_n2014_), .Y(new_n2087_));
  OR2X1    g01831(.A(new_n1838_), .B(new_n1834_), .Y(new_n2088_));
  INVX1    g01832(.A(new_n1838_), .Y(new_n2089_));
  XOR2X1   g01833(.A(new_n2089_), .B(new_n1834_), .Y(new_n2090_));
  OAI21X1  g01834(.A0(new_n1843_), .A1(new_n2090_), .B0(new_n2088_), .Y(new_n2091_));
  AOI21X1  g01835(.A0(new_n2091_), .A1(new_n2015_), .B0(new_n2087_), .Y(new_n2092_));
  XOR2X1   g01836(.A(new_n2092_), .B(new_n2086_), .Y(new_n2093_));
  AOI22X1  g01837(.A0(new_n603_), .A1(\b[20] ), .B0(new_n602_), .B1(\b[19] ), .Y(new_n2094_));
  OAI21X1  g01838(.A0(new_n601_), .A1(new_n1115_), .B0(new_n2094_), .Y(new_n2095_));
  AOI21X1  g01839(.A0(new_n1217_), .A1(new_n518_), .B0(new_n2095_), .Y(new_n2096_));
  XOR2X1   g01840(.A(new_n2096_), .B(\a[11] ), .Y(new_n2097_));
  NAND2X1  g01841(.A(new_n2097_), .B(new_n2093_), .Y(new_n2098_));
  NOR2X1   g01842(.A(new_n2097_), .B(new_n2093_), .Y(new_n2099_));
  AND2X1   g01843(.A(new_n2097_), .B(new_n2093_), .Y(new_n2100_));
  OR2X1    g01844(.A(new_n2100_), .B(new_n2099_), .Y(new_n2101_));
  AOI21X1  g01845(.A0(new_n2098_), .A1(new_n2028_), .B0(new_n2099_), .Y(new_n2102_));
  AOI22X1  g01846(.A0(new_n2102_), .A1(new_n2098_), .B0(new_n2101_), .B1(new_n2028_), .Y(new_n2103_));
  AOI22X1  g01847(.A0(new_n469_), .A1(\b[23] ), .B0(new_n468_), .B1(\b[22] ), .Y(new_n2104_));
  OAI21X1  g01848(.A0(new_n467_), .A1(new_n1482_), .B0(new_n2104_), .Y(new_n2105_));
  AOI21X1  g01849(.A0(new_n1481_), .A1(new_n404_), .B0(new_n2105_), .Y(new_n2106_));
  XOR2X1   g01850(.A(new_n2106_), .B(\a[8] ), .Y(new_n2107_));
  INVX1    g01851(.A(new_n2107_), .Y(new_n2108_));
  XOR2X1   g01852(.A(new_n2108_), .B(new_n2103_), .Y(new_n2109_));
  NOR2X1   g01853(.A(new_n1984_), .B(new_n2018_), .Y(new_n2110_));
  OR2X1    g01854(.A(new_n1856_), .B(new_n1852_), .Y(new_n2111_));
  XOR2X1   g01855(.A(new_n1843_), .B(new_n2090_), .Y(new_n2112_));
  XOR2X1   g01856(.A(new_n1848_), .B(new_n2112_), .Y(new_n2113_));
  XOR2X1   g01857(.A(new_n1851_), .B(new_n2113_), .Y(new_n2114_));
  XOR2X1   g01858(.A(new_n1856_), .B(new_n2114_), .Y(new_n2115_));
  OAI21X1  g01859(.A0(new_n1863_), .A1(new_n2115_), .B0(new_n2111_), .Y(new_n2116_));
  AOI21X1  g01860(.A0(new_n2116_), .A1(new_n2019_), .B0(new_n2110_), .Y(new_n2117_));
  XOR2X1   g01861(.A(new_n2117_), .B(new_n2109_), .Y(new_n2118_));
  XOR2X1   g01862(.A(new_n2118_), .B(new_n2026_), .Y(new_n2119_));
  XOR2X1   g01863(.A(new_n2119_), .B(new_n2022_), .Y(new_n2120_));
  AND2X1   g01864(.A(\b[28] ), .B(\b[27] ), .Y(new_n2121_));
  AOI21X1  g01865(.A0(new_n2003_), .A1(new_n2002_), .B0(new_n2121_), .Y(new_n2122_));
  XOR2X1   g01866(.A(\b[29] ), .B(\b[28] ), .Y(new_n2123_));
  INVX1    g01867(.A(new_n2123_), .Y(new_n2124_));
  XOR2X1   g01868(.A(new_n2124_), .B(new_n2122_), .Y(new_n2125_));
  INVX1    g01869(.A(\b[27] ), .Y(new_n2126_));
  AOI22X1  g01870(.A0(new_n267_), .A1(\b[29] ), .B0(new_n266_), .B1(\b[28] ), .Y(new_n2127_));
  OAI21X1  g01871(.A0(new_n350_), .A1(new_n2126_), .B0(new_n2127_), .Y(new_n2128_));
  AOI21X1  g01872(.A0(new_n2125_), .A1(new_n318_), .B0(new_n2128_), .Y(new_n2129_));
  XOR2X1   g01873(.A(new_n2129_), .B(\a[2] ), .Y(new_n2130_));
  XOR2X1   g01874(.A(new_n2130_), .B(new_n2120_), .Y(new_n2131_));
  XOR2X1   g01875(.A(new_n1994_), .B(new_n2020_), .Y(new_n2132_));
  XOR2X1   g01876(.A(new_n1999_), .B(new_n2132_), .Y(new_n2133_));
  NOR2X1   g01877(.A(new_n2008_), .B(new_n2133_), .Y(new_n2134_));
  AOI21X1  g01878(.A0(new_n1888_), .A1(new_n1887_), .B0(new_n2009_), .Y(new_n2135_));
  OR2X1    g01879(.A(new_n2135_), .B(new_n2134_), .Y(new_n2136_));
  XOR2X1   g01880(.A(new_n2136_), .B(new_n2131_), .Y(\f[29] ));
  OR2X1    g01881(.A(new_n2107_), .B(new_n2103_), .Y(new_n2138_));
  OAI21X1  g01882(.A0(new_n2117_), .A1(new_n2109_), .B0(new_n2138_), .Y(new_n2139_));
  NOR2X1   g01883(.A(new_n1967_), .B(new_n2016_), .Y(new_n2140_));
  OR2X1    g01884(.A(new_n1848_), .B(new_n1844_), .Y(new_n2141_));
  OAI21X1  g01885(.A0(new_n1851_), .A1(new_n2113_), .B0(new_n2141_), .Y(new_n2142_));
  AOI21X1  g01886(.A0(new_n2142_), .A1(new_n2017_), .B0(new_n2140_), .Y(new_n2143_));
  OR2X1    g01887(.A(new_n2097_), .B(new_n2093_), .Y(new_n2144_));
  OAI21X1  g01888(.A0(new_n2100_), .A1(new_n2143_), .B0(new_n2144_), .Y(new_n2145_));
  NAND2X1  g01889(.A(new_n2067_), .B(new_n2036_), .Y(new_n2146_));
  OAI21X1  g01890(.A0(new_n2031_), .A1(new_n2030_), .B0(new_n2068_), .Y(new_n2147_));
  AND2X1   g01891(.A(new_n2147_), .B(new_n2146_), .Y(new_n2148_));
  AOI22X1  g01892(.A0(new_n1263_), .A1(\b[12] ), .B0(new_n1262_), .B1(\b[11] ), .Y(new_n2149_));
  OAI21X1  g01893(.A0(new_n1261_), .A1(new_n587_), .B0(new_n2149_), .Y(new_n2150_));
  AOI21X1  g01894(.A0(new_n1075_), .A1(new_n635_), .B0(new_n2150_), .Y(new_n2151_));
  XOR2X1   g01895(.A(new_n2151_), .B(new_n1072_), .Y(new_n2152_));
  AOI21X1  g01896(.A0(new_n2060_), .A1(new_n2056_), .B0(new_n2065_), .Y(new_n2153_));
  AND2X1   g01897(.A(new_n2066_), .B(new_n2039_), .Y(new_n2154_));
  OR2X1    g01898(.A(new_n2154_), .B(new_n2153_), .Y(new_n2155_));
  OAI21X1  g01899(.A0(new_n2058_), .A1(new_n2041_), .B0(new_n2057_), .Y(new_n2156_));
  OR4X1    g01900(.A(new_n2048_), .B(new_n1916_), .C(new_n1896_), .D(new_n1911_), .Y(new_n2157_));
  XOR2X1   g01901(.A(\a[30] ), .B(\a[29] ), .Y(new_n2158_));
  NAND2X1  g01902(.A(new_n2158_), .B(\b[0] ), .Y(new_n2159_));
  XOR2X1   g01903(.A(new_n2159_), .B(new_n2157_), .Y(new_n2160_));
  INVX1    g01904(.A(new_n2045_), .Y(new_n2161_));
  AND2X1   g01905(.A(new_n1909_), .B(new_n1908_), .Y(new_n2162_));
  AND2X1   g01906(.A(new_n1912_), .B(new_n1809_), .Y(new_n2163_));
  AOI22X1  g01907(.A0(new_n2163_), .A1(\b[3] ), .B0(new_n2162_), .B1(\b[2] ), .Y(new_n2164_));
  OAI21X1  g01908(.A0(new_n2161_), .A1(new_n275_), .B0(new_n2164_), .Y(new_n2165_));
  AOI21X1  g01909(.A0(new_n1907_), .A1(new_n366_), .B0(new_n2165_), .Y(new_n2166_));
  XOR2X1   g01910(.A(new_n2166_), .B(\a[29] ), .Y(new_n2167_));
  XOR2X1   g01911(.A(new_n2167_), .B(new_n2160_), .Y(new_n2168_));
  AOI22X1  g01912(.A0(new_n1814_), .A1(\b[6] ), .B0(new_n1813_), .B1(\b[5] ), .Y(new_n2169_));
  OAI21X1  g01913(.A0(new_n1812_), .A1(new_n325_), .B0(new_n2169_), .Y(new_n2170_));
  AOI21X1  g01914(.A0(new_n1617_), .A1(new_n378_), .B0(new_n2170_), .Y(new_n2171_));
  XOR2X1   g01915(.A(new_n2171_), .B(\a[26] ), .Y(new_n2172_));
  XOR2X1   g01916(.A(new_n2172_), .B(new_n2168_), .Y(new_n2173_));
  INVX1    g01917(.A(new_n2173_), .Y(new_n2174_));
  XOR2X1   g01918(.A(new_n2174_), .B(new_n2156_), .Y(new_n2175_));
  AOI22X1  g01919(.A0(new_n1526_), .A1(\b[9] ), .B0(new_n1525_), .B1(\b[8] ), .Y(new_n2176_));
  OAI21X1  g01920(.A0(new_n1524_), .A1(new_n492_), .B0(new_n2176_), .Y(new_n2177_));
  AOI21X1  g01921(.A0(new_n1347_), .A1(new_n491_), .B0(new_n2177_), .Y(new_n2178_));
  XOR2X1   g01922(.A(new_n2178_), .B(\a[23] ), .Y(new_n2179_));
  XOR2X1   g01923(.A(new_n2179_), .B(new_n2175_), .Y(new_n2180_));
  XOR2X1   g01924(.A(new_n2180_), .B(new_n2155_), .Y(new_n2181_));
  XOR2X1   g01925(.A(new_n2181_), .B(new_n2152_), .Y(new_n2182_));
  XOR2X1   g01926(.A(new_n2182_), .B(new_n2148_), .Y(new_n2183_));
  AOI22X1  g01927(.A0(new_n1017_), .A1(\b[15] ), .B0(new_n1016_), .B1(\b[14] ), .Y(new_n2184_));
  OAI21X1  g01928(.A0(new_n1015_), .A1(new_n795_), .B0(new_n2184_), .Y(new_n2185_));
  AOI21X1  g01929(.A0(new_n882_), .A1(new_n794_), .B0(new_n2185_), .Y(new_n2186_));
  XOR2X1   g01930(.A(new_n2186_), .B(\a[17] ), .Y(new_n2187_));
  INVX1    g01931(.A(new_n2187_), .Y(new_n2188_));
  XOR2X1   g01932(.A(new_n2188_), .B(new_n2183_), .Y(new_n2189_));
  AND2X1   g01933(.A(new_n2074_), .B(new_n2069_), .Y(new_n2190_));
  OR2X1    g01934(.A(new_n1934_), .B(new_n2012_), .Y(new_n2191_));
  OAI21X1  g01935(.A0(new_n1947_), .A1(new_n1935_), .B0(new_n2191_), .Y(new_n2192_));
  AOI21X1  g01936(.A0(new_n2192_), .A1(new_n2075_), .B0(new_n2190_), .Y(new_n2193_));
  XOR2X1   g01937(.A(new_n2193_), .B(new_n2189_), .Y(new_n2194_));
  AOI22X1  g01938(.A0(new_n818_), .A1(\b[18] ), .B0(new_n817_), .B1(\b[17] ), .Y(new_n2195_));
  OAI21X1  g01939(.A0(new_n816_), .A1(new_n974_), .B0(new_n2195_), .Y(new_n2196_));
  AOI21X1  g01940(.A0(new_n1042_), .A1(new_n668_), .B0(new_n2196_), .Y(new_n2197_));
  XOR2X1   g01941(.A(new_n2197_), .B(\a[14] ), .Y(new_n2198_));
  XOR2X1   g01942(.A(new_n2198_), .B(new_n2194_), .Y(new_n2199_));
  NOR2X1   g01943(.A(new_n2085_), .B(new_n2081_), .Y(new_n2200_));
  OR2X1    g01944(.A(new_n1952_), .B(new_n2014_), .Y(new_n2201_));
  OAI21X1  g01945(.A0(new_n1962_), .A1(new_n1953_), .B0(new_n2201_), .Y(new_n2202_));
  AOI21X1  g01946(.A0(new_n2202_), .A1(new_n2086_), .B0(new_n2200_), .Y(new_n2203_));
  XOR2X1   g01947(.A(new_n2203_), .B(new_n2199_), .Y(new_n2204_));
  AOI22X1  g01948(.A0(new_n603_), .A1(\b[21] ), .B0(new_n602_), .B1(\b[20] ), .Y(new_n2205_));
  OAI21X1  g01949(.A0(new_n601_), .A1(new_n1300_), .B0(new_n2205_), .Y(new_n2206_));
  AOI21X1  g01950(.A0(new_n1299_), .A1(new_n518_), .B0(new_n2206_), .Y(new_n2207_));
  XOR2X1   g01951(.A(new_n2207_), .B(\a[11] ), .Y(new_n2208_));
  XOR2X1   g01952(.A(new_n2208_), .B(new_n2204_), .Y(new_n2209_));
  XOR2X1   g01953(.A(new_n2209_), .B(new_n2145_), .Y(new_n2210_));
  AOI22X1  g01954(.A0(new_n469_), .A1(\b[24] ), .B0(new_n468_), .B1(\b[23] ), .Y(new_n2211_));
  OAI21X1  g01955(.A0(new_n467_), .A1(new_n1479_), .B0(new_n2211_), .Y(new_n2212_));
  AOI21X1  g01956(.A0(new_n1572_), .A1(new_n404_), .B0(new_n2212_), .Y(new_n2213_));
  XOR2X1   g01957(.A(new_n2213_), .B(\a[8] ), .Y(new_n2214_));
  XOR2X1   g01958(.A(new_n2214_), .B(new_n2210_), .Y(new_n2215_));
  XOR2X1   g01959(.A(new_n2215_), .B(new_n2139_), .Y(new_n2216_));
  AOI22X1  g01960(.A0(new_n369_), .A1(\b[27] ), .B0(new_n368_), .B1(\b[26] ), .Y(new_n2217_));
  OAI21X1  g01961(.A0(new_n367_), .A1(new_n1880_), .B0(new_n2217_), .Y(new_n2218_));
  AOI21X1  g01962(.A0(new_n1879_), .A1(new_n308_), .B0(new_n2218_), .Y(new_n2219_));
  XOR2X1   g01963(.A(new_n2219_), .B(\a[5] ), .Y(new_n2220_));
  XOR2X1   g01964(.A(new_n2220_), .B(new_n2216_), .Y(new_n2221_));
  INVX1    g01965(.A(new_n2026_), .Y(new_n2222_));
  AND2X1   g01966(.A(new_n2118_), .B(new_n2222_), .Y(new_n2223_));
  XOR2X1   g01967(.A(new_n2118_), .B(new_n2222_), .Y(new_n2224_));
  AOI21X1  g01968(.A0(new_n2224_), .A1(new_n2022_), .B0(new_n2223_), .Y(new_n2225_));
  XOR2X1   g01969(.A(new_n2225_), .B(new_n2221_), .Y(new_n2226_));
  NAND2X1  g01970(.A(\b[29] ), .B(\b[28] ), .Y(new_n2227_));
  OAI21X1  g01971(.A0(new_n2124_), .A1(new_n2122_), .B0(new_n2227_), .Y(new_n2228_));
  XOR2X1   g01972(.A(\b[30] ), .B(\b[29] ), .Y(new_n2229_));
  XOR2X1   g01973(.A(new_n2229_), .B(new_n2228_), .Y(new_n2230_));
  INVX1    g01974(.A(\b[28] ), .Y(new_n2231_));
  AOI22X1  g01975(.A0(new_n267_), .A1(\b[30] ), .B0(new_n266_), .B1(\b[29] ), .Y(new_n2232_));
  OAI21X1  g01976(.A0(new_n350_), .A1(new_n2231_), .B0(new_n2232_), .Y(new_n2233_));
  AOI21X1  g01977(.A0(new_n2230_), .A1(new_n318_), .B0(new_n2233_), .Y(new_n2234_));
  XOR2X1   g01978(.A(new_n2234_), .B(\a[2] ), .Y(new_n2235_));
  XOR2X1   g01979(.A(new_n2235_), .B(new_n2226_), .Y(new_n2236_));
  OR2X1    g01980(.A(new_n2130_), .B(new_n2120_), .Y(new_n2237_));
  OAI21X1  g01981(.A0(new_n2135_), .A1(new_n2134_), .B0(new_n2131_), .Y(new_n2238_));
  AND2X1   g01982(.A(new_n2238_), .B(new_n2237_), .Y(new_n2239_));
  XOR2X1   g01983(.A(new_n2239_), .B(new_n2236_), .Y(\f[30] ));
  NOR2X1   g01984(.A(new_n2172_), .B(new_n2168_), .Y(new_n2241_));
  AOI21X1  g01985(.A0(new_n2173_), .A1(new_n2156_), .B0(new_n2241_), .Y(new_n2242_));
  AOI22X1  g01986(.A0(new_n1814_), .A1(\b[7] ), .B0(new_n1813_), .B1(\b[6] ), .Y(new_n2243_));
  OAI21X1  g01987(.A0(new_n1812_), .A1(new_n395_), .B0(new_n2243_), .Y(new_n2244_));
  AOI21X1  g01988(.A0(new_n1617_), .A1(new_n394_), .B0(new_n2244_), .Y(new_n2245_));
  XOR2X1   g01989(.A(new_n2245_), .B(new_n1621_), .Y(new_n2246_));
  INVX1    g01990(.A(new_n2159_), .Y(new_n2247_));
  XOR2X1   g01991(.A(new_n2247_), .B(new_n2157_), .Y(new_n2248_));
  OR2X1    g01992(.A(new_n2159_), .B(new_n2157_), .Y(new_n2249_));
  OAI21X1  g01993(.A0(new_n2167_), .A1(new_n2248_), .B0(new_n2249_), .Y(new_n2250_));
  AND2X1   g01994(.A(new_n1907_), .B(new_n323_), .Y(new_n2251_));
  NOR3X1   g01995(.A(new_n2044_), .B(new_n1912_), .C(new_n277_), .Y(new_n2252_));
  OAI22X1  g01996(.A0(new_n1913_), .A1(new_n325_), .B0(new_n1910_), .B1(new_n297_), .Y(new_n2253_));
  NOR3X1   g01997(.A(new_n2253_), .B(new_n2252_), .C(new_n2251_), .Y(new_n2254_));
  XOR2X1   g01998(.A(new_n2254_), .B(new_n1911_), .Y(new_n2255_));
  NAND2X1  g01999(.A(new_n2159_), .B(\a[32] ), .Y(new_n2256_));
  INVX1    g02000(.A(new_n2158_), .Y(new_n2257_));
  INVX1    g02001(.A(\a[32] ), .Y(new_n2258_));
  XOR2X1   g02002(.A(new_n2258_), .B(\a[31] ), .Y(new_n2259_));
  NOR2X1   g02003(.A(new_n2259_), .B(new_n2257_), .Y(new_n2260_));
  XOR2X1   g02004(.A(\a[31] ), .B(\a[30] ), .Y(new_n2261_));
  NAND2X1  g02005(.A(new_n2261_), .B(new_n2257_), .Y(new_n2262_));
  NAND2X1  g02006(.A(new_n2259_), .B(new_n2158_), .Y(new_n2263_));
  OAI22X1  g02007(.A0(new_n2263_), .A1(new_n275_), .B0(new_n2262_), .B1(new_n274_), .Y(new_n2264_));
  AOI21X1  g02008(.A0(new_n2260_), .A1(new_n263_), .B0(new_n2264_), .Y(new_n2265_));
  XOR2X1   g02009(.A(new_n2265_), .B(\a[32] ), .Y(new_n2266_));
  XOR2X1   g02010(.A(new_n2266_), .B(new_n2256_), .Y(new_n2267_));
  XOR2X1   g02011(.A(new_n2267_), .B(new_n2255_), .Y(new_n2268_));
  XOR2X1   g02012(.A(new_n2268_), .B(new_n2250_), .Y(new_n2269_));
  XOR2X1   g02013(.A(new_n2269_), .B(new_n2246_), .Y(new_n2270_));
  XOR2X1   g02014(.A(new_n2270_), .B(new_n2242_), .Y(new_n2271_));
  AOI22X1  g02015(.A0(new_n1526_), .A1(\b[10] ), .B0(new_n1525_), .B1(\b[9] ), .Y(new_n2272_));
  OAI21X1  g02016(.A0(new_n1524_), .A1(new_n489_), .B0(new_n2272_), .Y(new_n2273_));
  AOI21X1  g02017(.A0(new_n1347_), .A1(new_n543_), .B0(new_n2273_), .Y(new_n2274_));
  XOR2X1   g02018(.A(new_n2274_), .B(\a[23] ), .Y(new_n2275_));
  INVX1    g02019(.A(new_n2275_), .Y(new_n2276_));
  XOR2X1   g02020(.A(new_n2276_), .B(new_n2271_), .Y(new_n2277_));
  INVX1    g02021(.A(new_n2277_), .Y(new_n2278_));
  OR2X1    g02022(.A(new_n2179_), .B(new_n2175_), .Y(new_n2279_));
  OAI21X1  g02023(.A0(new_n2154_), .A1(new_n2153_), .B0(new_n2180_), .Y(new_n2280_));
  AND2X1   g02024(.A(new_n2280_), .B(new_n2279_), .Y(new_n2281_));
  XOR2X1   g02025(.A(new_n2281_), .B(new_n2278_), .Y(new_n2282_));
  AOI22X1  g02026(.A0(new_n1263_), .A1(\b[13] ), .B0(new_n1262_), .B1(\b[12] ), .Y(new_n2283_));
  OAI21X1  g02027(.A0(new_n1261_), .A1(new_n716_), .B0(new_n2283_), .Y(new_n2284_));
  AOI21X1  g02028(.A0(new_n1075_), .A1(new_n715_), .B0(new_n2284_), .Y(new_n2285_));
  XOR2X1   g02029(.A(new_n2285_), .B(\a[20] ), .Y(new_n2286_));
  XOR2X1   g02030(.A(new_n2286_), .B(new_n2282_), .Y(new_n2287_));
  NAND2X1  g02031(.A(new_n2147_), .B(new_n2146_), .Y(new_n2288_));
  AND2X1   g02032(.A(new_n2181_), .B(new_n2152_), .Y(new_n2289_));
  AOI21X1  g02033(.A0(new_n2182_), .A1(new_n2288_), .B0(new_n2289_), .Y(new_n2290_));
  XOR2X1   g02034(.A(new_n2290_), .B(new_n2287_), .Y(new_n2291_));
  AOI22X1  g02035(.A0(new_n1017_), .A1(\b[16] ), .B0(new_n1016_), .B1(\b[15] ), .Y(new_n2292_));
  OAI21X1  g02036(.A0(new_n1015_), .A1(new_n792_), .B0(new_n2292_), .Y(new_n2293_));
  AOI21X1  g02037(.A0(new_n882_), .A1(new_n842_), .B0(new_n2293_), .Y(new_n2294_));
  XOR2X1   g02038(.A(new_n2294_), .B(\a[17] ), .Y(new_n2295_));
  XOR2X1   g02039(.A(new_n2295_), .B(new_n2291_), .Y(new_n2296_));
  NOR2X1   g02040(.A(new_n2187_), .B(new_n2183_), .Y(new_n2297_));
  XOR2X1   g02041(.A(new_n2187_), .B(new_n2183_), .Y(new_n2298_));
  NAND2X1  g02042(.A(new_n2074_), .B(new_n2069_), .Y(new_n2299_));
  XOR2X1   g02043(.A(new_n2073_), .B(new_n2069_), .Y(new_n2300_));
  OAI21X1  g02044(.A0(new_n2080_), .A1(new_n2300_), .B0(new_n2299_), .Y(new_n2301_));
  AOI21X1  g02045(.A0(new_n2301_), .A1(new_n2298_), .B0(new_n2297_), .Y(new_n2302_));
  XOR2X1   g02046(.A(new_n2302_), .B(new_n2296_), .Y(new_n2303_));
  AOI22X1  g02047(.A0(new_n818_), .A1(\b[19] ), .B0(new_n817_), .B1(\b[18] ), .Y(new_n2304_));
  OAI21X1  g02048(.A0(new_n816_), .A1(new_n1118_), .B0(new_n2304_), .Y(new_n2305_));
  AOI21X1  g02049(.A0(new_n1117_), .A1(new_n668_), .B0(new_n2305_), .Y(new_n2306_));
  XOR2X1   g02050(.A(new_n2306_), .B(\a[14] ), .Y(new_n2307_));
  XOR2X1   g02051(.A(new_n2307_), .B(new_n2303_), .Y(new_n2308_));
  XOR2X1   g02052(.A(new_n2193_), .B(new_n2298_), .Y(new_n2309_));
  NOR2X1   g02053(.A(new_n2198_), .B(new_n2309_), .Y(new_n2310_));
  XOR2X1   g02054(.A(new_n2198_), .B(new_n2309_), .Y(new_n2311_));
  OR2X1    g02055(.A(new_n2085_), .B(new_n2081_), .Y(new_n2312_));
  XOR2X1   g02056(.A(new_n2080_), .B(new_n2300_), .Y(new_n2313_));
  XOR2X1   g02057(.A(new_n2085_), .B(new_n2313_), .Y(new_n2314_));
  OAI21X1  g02058(.A0(new_n2092_), .A1(new_n2314_), .B0(new_n2312_), .Y(new_n2315_));
  AOI21X1  g02059(.A0(new_n2315_), .A1(new_n2311_), .B0(new_n2310_), .Y(new_n2316_));
  XOR2X1   g02060(.A(new_n2316_), .B(new_n2308_), .Y(new_n2317_));
  AOI22X1  g02061(.A0(new_n603_), .A1(\b[22] ), .B0(new_n602_), .B1(\b[21] ), .Y(new_n2318_));
  OAI21X1  g02062(.A0(new_n601_), .A1(new_n1297_), .B0(new_n2318_), .Y(new_n2319_));
  AOI21X1  g02063(.A0(new_n1399_), .A1(new_n518_), .B0(new_n2319_), .Y(new_n2320_));
  XOR2X1   g02064(.A(new_n2320_), .B(\a[11] ), .Y(new_n2321_));
  XOR2X1   g02065(.A(new_n2321_), .B(new_n2317_), .Y(new_n2322_));
  XOR2X1   g02066(.A(new_n2203_), .B(new_n2311_), .Y(new_n2323_));
  NOR2X1   g02067(.A(new_n2208_), .B(new_n2323_), .Y(new_n2324_));
  XOR2X1   g02068(.A(new_n2208_), .B(new_n2323_), .Y(new_n2325_));
  AOI21X1  g02069(.A0(new_n2325_), .A1(new_n2145_), .B0(new_n2324_), .Y(new_n2326_));
  XOR2X1   g02070(.A(new_n2326_), .B(new_n2322_), .Y(new_n2327_));
  AOI22X1  g02071(.A0(new_n469_), .A1(\b[25] ), .B0(new_n468_), .B1(\b[24] ), .Y(new_n2328_));
  OAI21X1  g02072(.A0(new_n467_), .A1(new_n1591_), .B0(new_n2328_), .Y(new_n2329_));
  AOI21X1  g02073(.A0(new_n1590_), .A1(new_n404_), .B0(new_n2329_), .Y(new_n2330_));
  XOR2X1   g02074(.A(new_n2330_), .B(\a[8] ), .Y(new_n2331_));
  XOR2X1   g02075(.A(new_n2331_), .B(new_n2327_), .Y(new_n2332_));
  NOR2X1   g02076(.A(new_n2214_), .B(new_n2210_), .Y(new_n2333_));
  AOI21X1  g02077(.A0(new_n2215_), .A1(new_n2139_), .B0(new_n2333_), .Y(new_n2334_));
  XOR2X1   g02078(.A(new_n2334_), .B(new_n2332_), .Y(new_n2335_));
  AOI22X1  g02079(.A0(new_n369_), .A1(\b[28] ), .B0(new_n368_), .B1(\b[27] ), .Y(new_n2336_));
  OAI21X1  g02080(.A0(new_n367_), .A1(new_n1877_), .B0(new_n2336_), .Y(new_n2337_));
  AOI21X1  g02081(.A0(new_n2004_), .A1(new_n308_), .B0(new_n2337_), .Y(new_n2338_));
  XOR2X1   g02082(.A(new_n2338_), .B(\a[5] ), .Y(new_n2339_));
  XOR2X1   g02083(.A(new_n2339_), .B(new_n2335_), .Y(new_n2340_));
  INVX1    g02084(.A(new_n2220_), .Y(new_n2341_));
  AND2X1   g02085(.A(new_n2341_), .B(new_n2216_), .Y(new_n2342_));
  XOR2X1   g02086(.A(new_n2341_), .B(new_n2216_), .Y(new_n2343_));
  NOR2X1   g02087(.A(new_n1994_), .B(new_n2020_), .Y(new_n2344_));
  OR2X1    g02088(.A(new_n1868_), .B(new_n1864_), .Y(new_n2345_));
  XOR2X1   g02089(.A(new_n1863_), .B(new_n2115_), .Y(new_n2346_));
  XOR2X1   g02090(.A(new_n1868_), .B(new_n2346_), .Y(new_n2347_));
  OAI21X1  g02091(.A0(new_n1873_), .A1(new_n2347_), .B0(new_n2345_), .Y(new_n2348_));
  AOI21X1  g02092(.A0(new_n2348_), .A1(new_n2132_), .B0(new_n2344_), .Y(new_n2349_));
  NAND2X1  g02093(.A(new_n2118_), .B(new_n2222_), .Y(new_n2350_));
  OAI21X1  g02094(.A0(new_n2119_), .A1(new_n2349_), .B0(new_n2350_), .Y(new_n2351_));
  AOI21X1  g02095(.A0(new_n2351_), .A1(new_n2343_), .B0(new_n2342_), .Y(new_n2352_));
  XOR2X1   g02096(.A(new_n2352_), .B(new_n2340_), .Y(new_n2353_));
  AND2X1   g02097(.A(\b[30] ), .B(\b[29] ), .Y(new_n2354_));
  AOI21X1  g02098(.A0(new_n2229_), .A1(new_n2228_), .B0(new_n2354_), .Y(new_n2355_));
  INVX1    g02099(.A(\b[30] ), .Y(new_n2356_));
  XOR2X1   g02100(.A(\b[31] ), .B(new_n2356_), .Y(new_n2357_));
  XOR2X1   g02101(.A(new_n2357_), .B(new_n2355_), .Y(new_n2358_));
  INVX1    g02102(.A(\b[29] ), .Y(new_n2359_));
  AOI22X1  g02103(.A0(new_n267_), .A1(\b[31] ), .B0(new_n266_), .B1(\b[30] ), .Y(new_n2360_));
  OAI21X1  g02104(.A0(new_n350_), .A1(new_n2359_), .B0(new_n2360_), .Y(new_n2361_));
  AOI21X1  g02105(.A0(new_n2358_), .A1(new_n318_), .B0(new_n2361_), .Y(new_n2362_));
  XOR2X1   g02106(.A(new_n2362_), .B(\a[2] ), .Y(new_n2363_));
  XOR2X1   g02107(.A(new_n2363_), .B(new_n2353_), .Y(new_n2364_));
  XOR2X1   g02108(.A(new_n2225_), .B(new_n2343_), .Y(new_n2365_));
  NOR2X1   g02109(.A(new_n2235_), .B(new_n2365_), .Y(new_n2366_));
  AOI21X1  g02110(.A0(new_n2238_), .A1(new_n2237_), .B0(new_n2236_), .Y(new_n2367_));
  OR2X1    g02111(.A(new_n2367_), .B(new_n2366_), .Y(new_n2368_));
  XOR2X1   g02112(.A(new_n2368_), .B(new_n2364_), .Y(\f[31] ));
  OR2X1    g02113(.A(new_n2363_), .B(new_n2353_), .Y(new_n2370_));
  OAI21X1  g02114(.A0(new_n2367_), .A1(new_n2366_), .B0(new_n2364_), .Y(new_n2371_));
  AND2X1   g02115(.A(new_n2371_), .B(new_n2370_), .Y(new_n2372_));
  OR2X1    g02116(.A(new_n2339_), .B(new_n2335_), .Y(new_n2373_));
  OR2X1    g02117(.A(new_n2187_), .B(new_n2183_), .Y(new_n2374_));
  OAI21X1  g02118(.A0(new_n2193_), .A1(new_n2189_), .B0(new_n2374_), .Y(new_n2375_));
  XOR2X1   g02119(.A(new_n2375_), .B(new_n2296_), .Y(new_n2376_));
  XOR2X1   g02120(.A(new_n2307_), .B(new_n2376_), .Y(new_n2377_));
  XOR2X1   g02121(.A(new_n2316_), .B(new_n2377_), .Y(new_n2378_));
  XOR2X1   g02122(.A(new_n2321_), .B(new_n2378_), .Y(new_n2379_));
  XOR2X1   g02123(.A(new_n2326_), .B(new_n2379_), .Y(new_n2380_));
  XOR2X1   g02124(.A(new_n2331_), .B(new_n2380_), .Y(new_n2381_));
  XOR2X1   g02125(.A(new_n2334_), .B(new_n2381_), .Y(new_n2382_));
  XOR2X1   g02126(.A(new_n2339_), .B(new_n2382_), .Y(new_n2383_));
  OAI21X1  g02127(.A0(new_n2352_), .A1(new_n2383_), .B0(new_n2373_), .Y(new_n2384_));
  NOR2X1   g02128(.A(new_n2321_), .B(new_n2317_), .Y(new_n2385_));
  OR2X1    g02129(.A(new_n2208_), .B(new_n2323_), .Y(new_n2386_));
  OAI21X1  g02130(.A0(new_n2209_), .A1(new_n2102_), .B0(new_n2386_), .Y(new_n2387_));
  AOI21X1  g02131(.A0(new_n2387_), .A1(new_n2322_), .B0(new_n2385_), .Y(new_n2388_));
  OR2X1    g02132(.A(new_n2307_), .B(new_n2303_), .Y(new_n2389_));
  OAI21X1  g02133(.A0(new_n2316_), .A1(new_n2377_), .B0(new_n2389_), .Y(new_n2390_));
  AND2X1   g02134(.A(new_n2286_), .B(new_n2282_), .Y(new_n2391_));
  OR2X1    g02135(.A(new_n2286_), .B(new_n2282_), .Y(new_n2392_));
  OAI21X1  g02136(.A0(new_n2290_), .A1(new_n2391_), .B0(new_n2392_), .Y(new_n2393_));
  NOR2X1   g02137(.A(new_n2275_), .B(new_n2271_), .Y(new_n2394_));
  AOI21X1  g02138(.A0(new_n2280_), .A1(new_n2279_), .B0(new_n2277_), .Y(new_n2395_));
  OR2X1    g02139(.A(new_n2395_), .B(new_n2394_), .Y(new_n2396_));
  AND2X1   g02140(.A(new_n2267_), .B(new_n2255_), .Y(new_n2397_));
  AOI21X1  g02141(.A0(new_n2268_), .A1(new_n2250_), .B0(new_n2397_), .Y(new_n2398_));
  NOR2X1   g02142(.A(new_n2266_), .B(new_n2256_), .Y(new_n2399_));
  INVX1    g02143(.A(new_n2260_), .Y(new_n2400_));
  OR2X1    g02144(.A(new_n2261_), .B(new_n2158_), .Y(new_n2401_));
  NOR2X1   g02145(.A(new_n2401_), .B(new_n2259_), .Y(new_n2402_));
  OAI22X1  g02146(.A0(new_n2263_), .A1(new_n277_), .B0(new_n2262_), .B1(new_n275_), .Y(new_n2403_));
  AOI21X1  g02147(.A0(new_n2402_), .A1(\b[0] ), .B0(new_n2403_), .Y(new_n2404_));
  OAI21X1  g02148(.A0(new_n2400_), .A1(new_n281_), .B0(new_n2404_), .Y(new_n2405_));
  XOR2X1   g02149(.A(new_n2405_), .B(new_n2258_), .Y(new_n2406_));
  XOR2X1   g02150(.A(new_n2406_), .B(new_n2399_), .Y(new_n2407_));
  AOI22X1  g02151(.A0(new_n2163_), .A1(\b[5] ), .B0(new_n2162_), .B1(\b[4] ), .Y(new_n2408_));
  OAI21X1  g02152(.A0(new_n2161_), .A1(new_n297_), .B0(new_n2408_), .Y(new_n2409_));
  AOI21X1  g02153(.A0(new_n1907_), .A1(new_n349_), .B0(new_n2409_), .Y(new_n2410_));
  XOR2X1   g02154(.A(new_n2410_), .B(\a[29] ), .Y(new_n2411_));
  AND2X1   g02155(.A(new_n2411_), .B(new_n2407_), .Y(new_n2412_));
  XOR2X1   g02156(.A(new_n2411_), .B(new_n2407_), .Y(new_n2413_));
  OR2X1    g02157(.A(new_n2411_), .B(new_n2407_), .Y(new_n2414_));
  OAI21X1  g02158(.A0(new_n2412_), .A1(new_n2398_), .B0(new_n2414_), .Y(new_n2415_));
  OAI22X1  g02159(.A0(new_n2415_), .A1(new_n2412_), .B0(new_n2413_), .B1(new_n2398_), .Y(new_n2416_));
  AOI22X1  g02160(.A0(new_n1814_), .A1(\b[8] ), .B0(new_n1813_), .B1(\b[7] ), .Y(new_n2417_));
  OAI21X1  g02161(.A0(new_n1812_), .A1(new_n392_), .B0(new_n2417_), .Y(new_n2418_));
  AOI21X1  g02162(.A0(new_n1617_), .A1(new_n454_), .B0(new_n2418_), .Y(new_n2419_));
  XOR2X1   g02163(.A(new_n2419_), .B(\a[26] ), .Y(new_n2420_));
  XOR2X1   g02164(.A(new_n2420_), .B(new_n2416_), .Y(new_n2421_));
  NAND2X1  g02165(.A(new_n2269_), .B(new_n2246_), .Y(new_n2422_));
  AND2X1   g02166(.A(new_n2173_), .B(new_n2156_), .Y(new_n2423_));
  OAI21X1  g02167(.A0(new_n2423_), .A1(new_n2241_), .B0(new_n2270_), .Y(new_n2424_));
  NAND2X1  g02168(.A(new_n2424_), .B(new_n2422_), .Y(new_n2425_));
  XOR2X1   g02169(.A(new_n2425_), .B(new_n2421_), .Y(new_n2426_));
  AOI22X1  g02170(.A0(new_n1526_), .A1(\b[11] ), .B0(new_n1525_), .B1(\b[10] ), .Y(new_n2427_));
  OAI21X1  g02171(.A0(new_n1524_), .A1(new_n590_), .B0(new_n2427_), .Y(new_n2428_));
  AOI21X1  g02172(.A0(new_n1347_), .A1(new_n589_), .B0(new_n2428_), .Y(new_n2429_));
  XOR2X1   g02173(.A(new_n2429_), .B(\a[23] ), .Y(new_n2430_));
  NAND2X1  g02174(.A(new_n2430_), .B(new_n2426_), .Y(new_n2431_));
  NOR2X1   g02175(.A(new_n2430_), .B(new_n2426_), .Y(new_n2432_));
  AND2X1   g02176(.A(new_n2430_), .B(new_n2426_), .Y(new_n2433_));
  OR2X1    g02177(.A(new_n2433_), .B(new_n2432_), .Y(new_n2434_));
  AOI21X1  g02178(.A0(new_n2431_), .A1(new_n2396_), .B0(new_n2432_), .Y(new_n2435_));
  AOI22X1  g02179(.A0(new_n2435_), .A1(new_n2431_), .B0(new_n2434_), .B1(new_n2396_), .Y(new_n2436_));
  AOI22X1  g02180(.A0(new_n1263_), .A1(\b[14] ), .B0(new_n1262_), .B1(\b[13] ), .Y(new_n2437_));
  OAI21X1  g02181(.A0(new_n1261_), .A1(new_n713_), .B0(new_n2437_), .Y(new_n2438_));
  AOI21X1  g02182(.A0(new_n1075_), .A1(new_n734_), .B0(new_n2438_), .Y(new_n2439_));
  XOR2X1   g02183(.A(new_n2439_), .B(\a[20] ), .Y(new_n2440_));
  XOR2X1   g02184(.A(new_n2440_), .B(new_n2436_), .Y(new_n2441_));
  XOR2X1   g02185(.A(new_n2441_), .B(new_n2393_), .Y(new_n2442_));
  AOI22X1  g02186(.A0(new_n1017_), .A1(\b[17] ), .B0(new_n1016_), .B1(\b[16] ), .Y(new_n2443_));
  OAI21X1  g02187(.A0(new_n1015_), .A1(new_n977_), .B0(new_n2443_), .Y(new_n2444_));
  AOI21X1  g02188(.A0(new_n976_), .A1(new_n882_), .B0(new_n2444_), .Y(new_n2445_));
  XOR2X1   g02189(.A(new_n2445_), .B(\a[17] ), .Y(new_n2446_));
  INVX1    g02190(.A(new_n2446_), .Y(new_n2447_));
  XOR2X1   g02191(.A(new_n2447_), .B(new_n2442_), .Y(new_n2448_));
  NOR2X1   g02192(.A(new_n2295_), .B(new_n2291_), .Y(new_n2449_));
  AOI21X1  g02193(.A0(new_n2375_), .A1(new_n2296_), .B0(new_n2449_), .Y(new_n2450_));
  XOR2X1   g02194(.A(new_n2450_), .B(new_n2448_), .Y(new_n2451_));
  AOI22X1  g02195(.A0(new_n818_), .A1(\b[20] ), .B0(new_n817_), .B1(\b[19] ), .Y(new_n2452_));
  OAI21X1  g02196(.A0(new_n816_), .A1(new_n1115_), .B0(new_n2452_), .Y(new_n2453_));
  AOI21X1  g02197(.A0(new_n1217_), .A1(new_n668_), .B0(new_n2453_), .Y(new_n2454_));
  XOR2X1   g02198(.A(new_n2454_), .B(\a[14] ), .Y(new_n2455_));
  NOR2X1   g02199(.A(new_n2455_), .B(new_n2451_), .Y(new_n2456_));
  AND2X1   g02200(.A(new_n2455_), .B(new_n2451_), .Y(new_n2457_));
  OR2X1    g02201(.A(new_n2457_), .B(new_n2456_), .Y(new_n2458_));
  NOR3X1   g02202(.A(new_n2457_), .B(new_n2456_), .C(new_n2390_), .Y(new_n2459_));
  AOI21X1  g02203(.A0(new_n2458_), .A1(new_n2390_), .B0(new_n2459_), .Y(new_n2460_));
  AOI22X1  g02204(.A0(new_n603_), .A1(\b[23] ), .B0(new_n602_), .B1(\b[22] ), .Y(new_n2461_));
  OAI21X1  g02205(.A0(new_n601_), .A1(new_n1482_), .B0(new_n2461_), .Y(new_n2462_));
  AOI21X1  g02206(.A0(new_n1481_), .A1(new_n518_), .B0(new_n2462_), .Y(new_n2463_));
  XOR2X1   g02207(.A(new_n2463_), .B(\a[11] ), .Y(new_n2464_));
  XOR2X1   g02208(.A(new_n2464_), .B(new_n2460_), .Y(new_n2465_));
  XOR2X1   g02209(.A(new_n2465_), .B(new_n2388_), .Y(new_n2466_));
  AOI22X1  g02210(.A0(new_n469_), .A1(\b[26] ), .B0(new_n468_), .B1(\b[25] ), .Y(new_n2467_));
  OAI21X1  g02211(.A0(new_n467_), .A1(new_n1588_), .B0(new_n2467_), .Y(new_n2468_));
  AOI21X1  g02212(.A0(new_n1783_), .A1(new_n404_), .B0(new_n2468_), .Y(new_n2469_));
  XOR2X1   g02213(.A(new_n2469_), .B(\a[8] ), .Y(new_n2470_));
  XOR2X1   g02214(.A(new_n2470_), .B(new_n2466_), .Y(new_n2471_));
  NOR2X1   g02215(.A(new_n2331_), .B(new_n2327_), .Y(new_n2472_));
  NOR2X1   g02216(.A(new_n2107_), .B(new_n2103_), .Y(new_n2473_));
  XOR2X1   g02217(.A(new_n2107_), .B(new_n2103_), .Y(new_n2474_));
  OR2X1    g02218(.A(new_n1984_), .B(new_n2018_), .Y(new_n2475_));
  OAI21X1  g02219(.A0(new_n1989_), .A1(new_n1985_), .B0(new_n2475_), .Y(new_n2476_));
  AOI21X1  g02220(.A0(new_n2476_), .A1(new_n2474_), .B0(new_n2473_), .Y(new_n2477_));
  OR2X1    g02221(.A(new_n2214_), .B(new_n2210_), .Y(new_n2478_));
  AND2X1   g02222(.A(new_n2214_), .B(new_n2210_), .Y(new_n2479_));
  OAI21X1  g02223(.A0(new_n2479_), .A1(new_n2477_), .B0(new_n2478_), .Y(new_n2480_));
  AOI21X1  g02224(.A0(new_n2480_), .A1(new_n2332_), .B0(new_n2472_), .Y(new_n2481_));
  XOR2X1   g02225(.A(new_n2481_), .B(new_n2471_), .Y(new_n2482_));
  AOI22X1  g02226(.A0(new_n369_), .A1(\b[29] ), .B0(new_n368_), .B1(\b[28] ), .Y(new_n2483_));
  OAI21X1  g02227(.A0(new_n367_), .A1(new_n2126_), .B0(new_n2483_), .Y(new_n2484_));
  AOI21X1  g02228(.A0(new_n2125_), .A1(new_n308_), .B0(new_n2484_), .Y(new_n2485_));
  XOR2X1   g02229(.A(new_n2485_), .B(\a[5] ), .Y(new_n2486_));
  NOR2X1   g02230(.A(new_n2486_), .B(new_n2482_), .Y(new_n2487_));
  AND2X1   g02231(.A(new_n2486_), .B(new_n2482_), .Y(new_n2488_));
  OR2X1    g02232(.A(new_n2488_), .B(new_n2487_), .Y(new_n2489_));
  AND2X1   g02233(.A(new_n2489_), .B(new_n2384_), .Y(new_n2490_));
  NOR3X1   g02234(.A(new_n2488_), .B(new_n2487_), .C(new_n2384_), .Y(new_n2491_));
  NAND2X1  g02235(.A(\b[31] ), .B(\b[30] ), .Y(new_n2492_));
  OAI21X1  g02236(.A0(new_n2357_), .A1(new_n2355_), .B0(new_n2492_), .Y(new_n2493_));
  XOR2X1   g02237(.A(\b[32] ), .B(\b[31] ), .Y(new_n2494_));
  XOR2X1   g02238(.A(new_n2494_), .B(new_n2493_), .Y(new_n2495_));
  AOI22X1  g02239(.A0(new_n267_), .A1(\b[32] ), .B0(new_n266_), .B1(\b[31] ), .Y(new_n2496_));
  OAI21X1  g02240(.A0(new_n350_), .A1(new_n2356_), .B0(new_n2496_), .Y(new_n2497_));
  AOI21X1  g02241(.A0(new_n2495_), .A1(new_n318_), .B0(new_n2497_), .Y(new_n2498_));
  XOR2X1   g02242(.A(new_n2498_), .B(\a[2] ), .Y(new_n2499_));
  OAI21X1  g02243(.A0(new_n2491_), .A1(new_n2490_), .B0(new_n2499_), .Y(new_n2500_));
  NAND2X1  g02244(.A(new_n2489_), .B(new_n2384_), .Y(new_n2501_));
  NOR2X1   g02245(.A(new_n2339_), .B(new_n2335_), .Y(new_n2502_));
  NAND2X1  g02246(.A(new_n2341_), .B(new_n2216_), .Y(new_n2503_));
  OAI21X1  g02247(.A0(new_n2225_), .A1(new_n2221_), .B0(new_n2503_), .Y(new_n2504_));
  AOI21X1  g02248(.A0(new_n2504_), .A1(new_n2340_), .B0(new_n2502_), .Y(new_n2505_));
  OR2X1    g02249(.A(new_n2486_), .B(new_n2482_), .Y(new_n2506_));
  NAND2X1  g02250(.A(new_n2486_), .B(new_n2482_), .Y(new_n2507_));
  NAND3X1  g02251(.A(new_n2507_), .B(new_n2506_), .C(new_n2505_), .Y(new_n2508_));
  XOR2X1   g02252(.A(new_n2498_), .B(new_n257_), .Y(new_n2509_));
  NAND3X1  g02253(.A(new_n2509_), .B(new_n2508_), .C(new_n2501_), .Y(new_n2510_));
  AND2X1   g02254(.A(new_n2510_), .B(new_n2500_), .Y(new_n2511_));
  XOR2X1   g02255(.A(new_n2511_), .B(new_n2372_), .Y(\f[32] ));
  AOI22X1  g02256(.A0(new_n2510_), .A1(new_n2500_), .B0(new_n2371_), .B1(new_n2370_), .Y(new_n2513_));
  AOI21X1  g02257(.A0(new_n2508_), .A1(new_n2501_), .B0(new_n2499_), .Y(new_n2514_));
  OR2X1    g02258(.A(new_n2514_), .B(new_n2513_), .Y(new_n2515_));
  OAI21X1  g02259(.A0(new_n2488_), .A1(new_n2505_), .B0(new_n2506_), .Y(new_n2516_));
  OR2X1    g02260(.A(new_n2321_), .B(new_n2317_), .Y(new_n2517_));
  OAI21X1  g02261(.A0(new_n2326_), .A1(new_n2379_), .B0(new_n2517_), .Y(new_n2518_));
  NOR2X1   g02262(.A(new_n2464_), .B(new_n2460_), .Y(new_n2519_));
  AOI21X1  g02263(.A0(new_n2465_), .A1(new_n2518_), .B0(new_n2519_), .Y(new_n2520_));
  NOR2X1   g02264(.A(new_n2307_), .B(new_n2303_), .Y(new_n2521_));
  OR2X1    g02265(.A(new_n2198_), .B(new_n2309_), .Y(new_n2522_));
  OAI21X1  g02266(.A0(new_n2203_), .A1(new_n2199_), .B0(new_n2522_), .Y(new_n2523_));
  AOI21X1  g02267(.A0(new_n2523_), .A1(new_n2308_), .B0(new_n2521_), .Y(new_n2524_));
  OR2X1    g02268(.A(new_n2455_), .B(new_n2451_), .Y(new_n2525_));
  OAI21X1  g02269(.A0(new_n2457_), .A1(new_n2524_), .B0(new_n2525_), .Y(new_n2526_));
  NAND2X1  g02270(.A(new_n2447_), .B(new_n2442_), .Y(new_n2527_));
  XOR2X1   g02271(.A(new_n2446_), .B(new_n2442_), .Y(new_n2528_));
  OAI21X1  g02272(.A0(new_n2450_), .A1(new_n2528_), .B0(new_n2527_), .Y(new_n2529_));
  NOR2X1   g02273(.A(new_n2440_), .B(new_n2436_), .Y(new_n2530_));
  AOI21X1  g02274(.A0(new_n2441_), .A1(new_n2393_), .B0(new_n2530_), .Y(new_n2531_));
  OR2X1    g02275(.A(new_n2413_), .B(new_n2398_), .Y(new_n2532_));
  INVX1    g02276(.A(new_n2412_), .Y(new_n2533_));
  NAND3X1  g02277(.A(new_n2533_), .B(new_n2414_), .C(new_n2398_), .Y(new_n2534_));
  AOI21X1  g02278(.A0(new_n2534_), .A1(new_n2532_), .B0(new_n2420_), .Y(new_n2535_));
  AOI21X1  g02279(.A0(new_n2424_), .A1(new_n2422_), .B0(new_n2421_), .Y(new_n2536_));
  NOR2X1   g02280(.A(new_n2536_), .B(new_n2535_), .Y(new_n2537_));
  OR4X1    g02281(.A(new_n2405_), .B(new_n2266_), .C(new_n2247_), .D(new_n2258_), .Y(new_n2538_));
  XOR2X1   g02282(.A(\a[33] ), .B(\a[32] ), .Y(new_n2539_));
  NAND2X1  g02283(.A(new_n2539_), .B(\b[0] ), .Y(new_n2540_));
  INVX1    g02284(.A(new_n2540_), .Y(new_n2541_));
  XOR2X1   g02285(.A(new_n2541_), .B(new_n2538_), .Y(new_n2542_));
  INVX1    g02286(.A(new_n2402_), .Y(new_n2543_));
  INVX1    g02287(.A(new_n2262_), .Y(new_n2544_));
  INVX1    g02288(.A(new_n2263_), .Y(new_n2545_));
  AOI22X1  g02289(.A0(new_n2545_), .A1(\b[3] ), .B0(new_n2544_), .B1(\b[2] ), .Y(new_n2546_));
  OAI21X1  g02290(.A0(new_n2543_), .A1(new_n275_), .B0(new_n2546_), .Y(new_n2547_));
  AOI21X1  g02291(.A0(new_n2260_), .A1(new_n366_), .B0(new_n2547_), .Y(new_n2548_));
  XOR2X1   g02292(.A(new_n2548_), .B(\a[32] ), .Y(new_n2549_));
  XOR2X1   g02293(.A(new_n2549_), .B(new_n2542_), .Y(new_n2550_));
  AOI22X1  g02294(.A0(new_n2163_), .A1(\b[6] ), .B0(new_n2162_), .B1(\b[5] ), .Y(new_n2551_));
  OAI21X1  g02295(.A0(new_n2161_), .A1(new_n325_), .B0(new_n2551_), .Y(new_n2552_));
  AOI21X1  g02296(.A0(new_n1907_), .A1(new_n378_), .B0(new_n2552_), .Y(new_n2553_));
  XOR2X1   g02297(.A(new_n2553_), .B(\a[29] ), .Y(new_n2554_));
  XOR2X1   g02298(.A(new_n2554_), .B(new_n2550_), .Y(new_n2555_));
  XOR2X1   g02299(.A(new_n2555_), .B(new_n2415_), .Y(new_n2556_));
  AOI22X1  g02300(.A0(new_n1814_), .A1(\b[9] ), .B0(new_n1813_), .B1(\b[8] ), .Y(new_n2557_));
  OAI21X1  g02301(.A0(new_n1812_), .A1(new_n492_), .B0(new_n2557_), .Y(new_n2558_));
  AOI21X1  g02302(.A0(new_n1617_), .A1(new_n491_), .B0(new_n2558_), .Y(new_n2559_));
  XOR2X1   g02303(.A(new_n2559_), .B(\a[26] ), .Y(new_n2560_));
  XOR2X1   g02304(.A(new_n2560_), .B(new_n2556_), .Y(new_n2561_));
  XOR2X1   g02305(.A(new_n2561_), .B(new_n2537_), .Y(new_n2562_));
  AOI22X1  g02306(.A0(new_n1526_), .A1(\b[12] ), .B0(new_n1525_), .B1(\b[11] ), .Y(new_n2563_));
  OAI21X1  g02307(.A0(new_n1524_), .A1(new_n587_), .B0(new_n2563_), .Y(new_n2564_));
  AOI21X1  g02308(.A0(new_n1347_), .A1(new_n635_), .B0(new_n2564_), .Y(new_n2565_));
  XOR2X1   g02309(.A(new_n2565_), .B(\a[23] ), .Y(new_n2566_));
  XOR2X1   g02310(.A(new_n2566_), .B(new_n2562_), .Y(new_n2567_));
  XOR2X1   g02311(.A(new_n2567_), .B(new_n2435_), .Y(new_n2568_));
  AOI22X1  g02312(.A0(new_n1263_), .A1(\b[15] ), .B0(new_n1262_), .B1(\b[14] ), .Y(new_n2569_));
  OAI21X1  g02313(.A0(new_n1261_), .A1(new_n795_), .B0(new_n2569_), .Y(new_n2570_));
  AOI21X1  g02314(.A0(new_n1075_), .A1(new_n794_), .B0(new_n2570_), .Y(new_n2571_));
  XOR2X1   g02315(.A(new_n2571_), .B(\a[20] ), .Y(new_n2572_));
  XOR2X1   g02316(.A(new_n2572_), .B(new_n2568_), .Y(new_n2573_));
  XOR2X1   g02317(.A(new_n2573_), .B(new_n2531_), .Y(new_n2574_));
  AOI22X1  g02318(.A0(new_n1017_), .A1(\b[18] ), .B0(new_n1016_), .B1(\b[17] ), .Y(new_n2575_));
  OAI21X1  g02319(.A0(new_n1015_), .A1(new_n974_), .B0(new_n2575_), .Y(new_n2576_));
  AOI21X1  g02320(.A0(new_n1042_), .A1(new_n882_), .B0(new_n2576_), .Y(new_n2577_));
  XOR2X1   g02321(.A(new_n2577_), .B(\a[17] ), .Y(new_n2578_));
  XOR2X1   g02322(.A(new_n2578_), .B(new_n2574_), .Y(new_n2579_));
  XOR2X1   g02323(.A(new_n2579_), .B(new_n2529_), .Y(new_n2580_));
  AOI22X1  g02324(.A0(new_n818_), .A1(\b[21] ), .B0(new_n817_), .B1(\b[20] ), .Y(new_n2581_));
  OAI21X1  g02325(.A0(new_n816_), .A1(new_n1300_), .B0(new_n2581_), .Y(new_n2582_));
  AOI21X1  g02326(.A0(new_n1299_), .A1(new_n668_), .B0(new_n2582_), .Y(new_n2583_));
  XOR2X1   g02327(.A(new_n2583_), .B(\a[14] ), .Y(new_n2584_));
  XOR2X1   g02328(.A(new_n2584_), .B(new_n2580_), .Y(new_n2585_));
  XOR2X1   g02329(.A(new_n2585_), .B(new_n2526_), .Y(new_n2586_));
  AOI22X1  g02330(.A0(new_n603_), .A1(\b[24] ), .B0(new_n602_), .B1(\b[23] ), .Y(new_n2587_));
  OAI21X1  g02331(.A0(new_n601_), .A1(new_n1479_), .B0(new_n2587_), .Y(new_n2588_));
  AOI21X1  g02332(.A0(new_n1572_), .A1(new_n518_), .B0(new_n2588_), .Y(new_n2589_));
  XOR2X1   g02333(.A(new_n2589_), .B(\a[11] ), .Y(new_n2590_));
  XOR2X1   g02334(.A(new_n2590_), .B(new_n2586_), .Y(new_n2591_));
  XOR2X1   g02335(.A(new_n2591_), .B(new_n2520_), .Y(new_n2592_));
  AOI22X1  g02336(.A0(new_n469_), .A1(\b[27] ), .B0(new_n468_), .B1(\b[26] ), .Y(new_n2593_));
  OAI21X1  g02337(.A0(new_n467_), .A1(new_n1880_), .B0(new_n2593_), .Y(new_n2594_));
  AOI21X1  g02338(.A0(new_n1879_), .A1(new_n404_), .B0(new_n2594_), .Y(new_n2595_));
  XOR2X1   g02339(.A(new_n2595_), .B(\a[8] ), .Y(new_n2596_));
  INVX1    g02340(.A(new_n2596_), .Y(new_n2597_));
  XOR2X1   g02341(.A(new_n2597_), .B(new_n2592_), .Y(new_n2598_));
  NOR2X1   g02342(.A(new_n2470_), .B(new_n2466_), .Y(new_n2599_));
  OR2X1    g02343(.A(new_n2331_), .B(new_n2327_), .Y(new_n2600_));
  OAI21X1  g02344(.A0(new_n2334_), .A1(new_n2381_), .B0(new_n2600_), .Y(new_n2601_));
  AOI21X1  g02345(.A0(new_n2601_), .A1(new_n2471_), .B0(new_n2599_), .Y(new_n2602_));
  XOR2X1   g02346(.A(new_n2602_), .B(new_n2598_), .Y(new_n2603_));
  AOI22X1  g02347(.A0(new_n369_), .A1(\b[30] ), .B0(new_n368_), .B1(\b[29] ), .Y(new_n2604_));
  OAI21X1  g02348(.A0(new_n367_), .A1(new_n2231_), .B0(new_n2604_), .Y(new_n2605_));
  AOI21X1  g02349(.A0(new_n2230_), .A1(new_n308_), .B0(new_n2605_), .Y(new_n2606_));
  XOR2X1   g02350(.A(new_n2606_), .B(\a[5] ), .Y(new_n2607_));
  XOR2X1   g02351(.A(new_n2607_), .B(new_n2603_), .Y(new_n2608_));
  XOR2X1   g02352(.A(new_n2608_), .B(new_n2516_), .Y(new_n2609_));
  AND2X1   g02353(.A(\b[32] ), .B(\b[31] ), .Y(new_n2610_));
  AOI21X1  g02354(.A0(new_n2494_), .A1(new_n2493_), .B0(new_n2610_), .Y(new_n2611_));
  INVX1    g02355(.A(\b[32] ), .Y(new_n2612_));
  XOR2X1   g02356(.A(\b[33] ), .B(new_n2612_), .Y(new_n2613_));
  XOR2X1   g02357(.A(new_n2613_), .B(new_n2611_), .Y(new_n2614_));
  INVX1    g02358(.A(\b[31] ), .Y(new_n2615_));
  AOI22X1  g02359(.A0(new_n267_), .A1(\b[33] ), .B0(new_n266_), .B1(\b[32] ), .Y(new_n2616_));
  OAI21X1  g02360(.A0(new_n350_), .A1(new_n2615_), .B0(new_n2616_), .Y(new_n2617_));
  AOI21X1  g02361(.A0(new_n2614_), .A1(new_n318_), .B0(new_n2617_), .Y(new_n2618_));
  XOR2X1   g02362(.A(new_n2618_), .B(\a[2] ), .Y(new_n2619_));
  XOR2X1   g02363(.A(new_n2619_), .B(new_n2609_), .Y(new_n2620_));
  XOR2X1   g02364(.A(new_n2620_), .B(new_n2515_), .Y(\f[33] ));
  OR2X1    g02365(.A(new_n2619_), .B(new_n2609_), .Y(new_n2622_));
  OAI21X1  g02366(.A0(new_n2514_), .A1(new_n2513_), .B0(new_n2620_), .Y(new_n2623_));
  AND2X1   g02367(.A(new_n2623_), .B(new_n2622_), .Y(new_n2624_));
  AOI21X1  g02368(.A0(new_n2507_), .A1(new_n2384_), .B0(new_n2487_), .Y(new_n2625_));
  XOR2X1   g02369(.A(new_n2596_), .B(new_n2592_), .Y(new_n2626_));
  XOR2X1   g02370(.A(new_n2602_), .B(new_n2626_), .Y(new_n2627_));
  OR2X1    g02371(.A(new_n2607_), .B(new_n2627_), .Y(new_n2628_));
  OAI21X1  g02372(.A0(new_n2608_), .A1(new_n2625_), .B0(new_n2628_), .Y(new_n2629_));
  AND2X1   g02373(.A(new_n2590_), .B(new_n2586_), .Y(new_n2630_));
  OR2X1    g02374(.A(new_n2590_), .B(new_n2586_), .Y(new_n2631_));
  OAI21X1  g02375(.A0(new_n2630_), .A1(new_n2520_), .B0(new_n2631_), .Y(new_n2632_));
  INVX1    g02376(.A(new_n2550_), .Y(new_n2633_));
  NOR2X1   g02377(.A(new_n2554_), .B(new_n2633_), .Y(new_n2634_));
  INVX1    g02378(.A(new_n2555_), .Y(new_n2635_));
  AOI21X1  g02379(.A0(new_n2635_), .A1(new_n2415_), .B0(new_n2634_), .Y(new_n2636_));
  AOI22X1  g02380(.A0(new_n2163_), .A1(\b[7] ), .B0(new_n2162_), .B1(\b[6] ), .Y(new_n2637_));
  OAI21X1  g02381(.A0(new_n2161_), .A1(new_n395_), .B0(new_n2637_), .Y(new_n2638_));
  AOI21X1  g02382(.A0(new_n1907_), .A1(new_n394_), .B0(new_n2638_), .Y(new_n2639_));
  XOR2X1   g02383(.A(new_n2639_), .B(new_n1911_), .Y(new_n2640_));
  OR2X1    g02384(.A(new_n2540_), .B(new_n2538_), .Y(new_n2641_));
  OAI21X1  g02385(.A0(new_n2549_), .A1(new_n2542_), .B0(new_n2641_), .Y(new_n2642_));
  AND2X1   g02386(.A(new_n2260_), .B(new_n323_), .Y(new_n2643_));
  NOR3X1   g02387(.A(new_n2401_), .B(new_n2259_), .C(new_n277_), .Y(new_n2644_));
  OAI22X1  g02388(.A0(new_n2263_), .A1(new_n325_), .B0(new_n2262_), .B1(new_n297_), .Y(new_n2645_));
  NOR3X1   g02389(.A(new_n2645_), .B(new_n2644_), .C(new_n2643_), .Y(new_n2646_));
  XOR2X1   g02390(.A(new_n2646_), .B(new_n2258_), .Y(new_n2647_));
  NAND2X1  g02391(.A(new_n2540_), .B(\a[35] ), .Y(new_n2648_));
  XOR2X1   g02392(.A(\a[33] ), .B(new_n2258_), .Y(new_n2649_));
  INVX1    g02393(.A(\a[35] ), .Y(new_n2650_));
  XOR2X1   g02394(.A(new_n2650_), .B(\a[34] ), .Y(new_n2651_));
  NOR2X1   g02395(.A(new_n2651_), .B(new_n2649_), .Y(new_n2652_));
  XOR2X1   g02396(.A(\a[34] ), .B(\a[33] ), .Y(new_n2653_));
  NAND2X1  g02397(.A(new_n2653_), .B(new_n2649_), .Y(new_n2654_));
  NAND2X1  g02398(.A(new_n2651_), .B(new_n2539_), .Y(new_n2655_));
  OAI22X1  g02399(.A0(new_n2655_), .A1(new_n275_), .B0(new_n2654_), .B1(new_n274_), .Y(new_n2656_));
  AOI21X1  g02400(.A0(new_n2652_), .A1(new_n263_), .B0(new_n2656_), .Y(new_n2657_));
  XOR2X1   g02401(.A(new_n2657_), .B(\a[35] ), .Y(new_n2658_));
  XOR2X1   g02402(.A(new_n2658_), .B(new_n2648_), .Y(new_n2659_));
  XOR2X1   g02403(.A(new_n2659_), .B(new_n2647_), .Y(new_n2660_));
  XOR2X1   g02404(.A(new_n2660_), .B(new_n2642_), .Y(new_n2661_));
  XOR2X1   g02405(.A(new_n2661_), .B(new_n2640_), .Y(new_n2662_));
  XOR2X1   g02406(.A(new_n2662_), .B(new_n2636_), .Y(new_n2663_));
  AOI22X1  g02407(.A0(new_n1814_), .A1(\b[10] ), .B0(new_n1813_), .B1(\b[9] ), .Y(new_n2664_));
  OAI21X1  g02408(.A0(new_n1812_), .A1(new_n489_), .B0(new_n2664_), .Y(new_n2665_));
  AOI21X1  g02409(.A0(new_n1617_), .A1(new_n543_), .B0(new_n2665_), .Y(new_n2666_));
  XOR2X1   g02410(.A(new_n2666_), .B(\a[26] ), .Y(new_n2667_));
  XOR2X1   g02411(.A(new_n2667_), .B(new_n2663_), .Y(new_n2668_));
  OR2X1    g02412(.A(new_n2560_), .B(new_n2556_), .Y(new_n2669_));
  OAI21X1  g02413(.A0(new_n2536_), .A1(new_n2535_), .B0(new_n2561_), .Y(new_n2670_));
  AND2X1   g02414(.A(new_n2670_), .B(new_n2669_), .Y(new_n2671_));
  XOR2X1   g02415(.A(new_n2671_), .B(new_n2668_), .Y(new_n2672_));
  AOI22X1  g02416(.A0(new_n1526_), .A1(\b[13] ), .B0(new_n1525_), .B1(\b[12] ), .Y(new_n2673_));
  OAI21X1  g02417(.A0(new_n1524_), .A1(new_n716_), .B0(new_n2673_), .Y(new_n2674_));
  AOI21X1  g02418(.A0(new_n1347_), .A1(new_n715_), .B0(new_n2674_), .Y(new_n2675_));
  XOR2X1   g02419(.A(new_n2675_), .B(\a[23] ), .Y(new_n2676_));
  NAND2X1  g02420(.A(new_n2676_), .B(new_n2672_), .Y(new_n2677_));
  NOR2X1   g02421(.A(new_n2395_), .B(new_n2394_), .Y(new_n2678_));
  OR2X1    g02422(.A(new_n2430_), .B(new_n2426_), .Y(new_n2679_));
  OAI21X1  g02423(.A0(new_n2433_), .A1(new_n2678_), .B0(new_n2679_), .Y(new_n2680_));
  NOR2X1   g02424(.A(new_n2566_), .B(new_n2562_), .Y(new_n2681_));
  AOI21X1  g02425(.A0(new_n2567_), .A1(new_n2680_), .B0(new_n2681_), .Y(new_n2682_));
  XOR2X1   g02426(.A(new_n2676_), .B(new_n2672_), .Y(new_n2683_));
  NOR2X1   g02427(.A(new_n2683_), .B(new_n2682_), .Y(new_n2684_));
  AND2X1   g02428(.A(new_n2566_), .B(new_n2562_), .Y(new_n2685_));
  OR2X1    g02429(.A(new_n2566_), .B(new_n2562_), .Y(new_n2686_));
  OAI21X1  g02430(.A0(new_n2685_), .A1(new_n2435_), .B0(new_n2686_), .Y(new_n2687_));
  NOR2X1   g02431(.A(new_n2676_), .B(new_n2672_), .Y(new_n2688_));
  AOI21X1  g02432(.A0(new_n2677_), .A1(new_n2687_), .B0(new_n2688_), .Y(new_n2689_));
  AOI21X1  g02433(.A0(new_n2689_), .A1(new_n2677_), .B0(new_n2684_), .Y(new_n2690_));
  AOI22X1  g02434(.A0(new_n1263_), .A1(\b[16] ), .B0(new_n1262_), .B1(\b[15] ), .Y(new_n2691_));
  OAI21X1  g02435(.A0(new_n1261_), .A1(new_n792_), .B0(new_n2691_), .Y(new_n2692_));
  AOI21X1  g02436(.A0(new_n1075_), .A1(new_n842_), .B0(new_n2692_), .Y(new_n2693_));
  XOR2X1   g02437(.A(new_n2693_), .B(\a[20] ), .Y(new_n2694_));
  XOR2X1   g02438(.A(new_n2694_), .B(new_n2690_), .Y(new_n2695_));
  NOR2X1   g02439(.A(new_n2286_), .B(new_n2282_), .Y(new_n2696_));
  NOR2X1   g02440(.A(new_n2181_), .B(new_n2152_), .Y(new_n2697_));
  NAND2X1  g02441(.A(new_n2181_), .B(new_n2152_), .Y(new_n2698_));
  OAI21X1  g02442(.A0(new_n2697_), .A1(new_n2148_), .B0(new_n2698_), .Y(new_n2699_));
  AOI21X1  g02443(.A0(new_n2699_), .A1(new_n2287_), .B0(new_n2696_), .Y(new_n2700_));
  AND2X1   g02444(.A(new_n2440_), .B(new_n2436_), .Y(new_n2701_));
  OR2X1    g02445(.A(new_n2440_), .B(new_n2436_), .Y(new_n2702_));
  OAI21X1  g02446(.A0(new_n2701_), .A1(new_n2700_), .B0(new_n2702_), .Y(new_n2703_));
  NOR2X1   g02447(.A(new_n2572_), .B(new_n2568_), .Y(new_n2704_));
  AOI21X1  g02448(.A0(new_n2573_), .A1(new_n2703_), .B0(new_n2704_), .Y(new_n2705_));
  XOR2X1   g02449(.A(new_n2705_), .B(new_n2695_), .Y(new_n2706_));
  AOI22X1  g02450(.A0(new_n1017_), .A1(\b[19] ), .B0(new_n1016_), .B1(\b[18] ), .Y(new_n2707_));
  OAI21X1  g02451(.A0(new_n1015_), .A1(new_n1118_), .B0(new_n2707_), .Y(new_n2708_));
  AOI21X1  g02452(.A0(new_n1117_), .A1(new_n882_), .B0(new_n2708_), .Y(new_n2709_));
  XOR2X1   g02453(.A(new_n2709_), .B(\a[17] ), .Y(new_n2710_));
  XOR2X1   g02454(.A(new_n2710_), .B(new_n2706_), .Y(new_n2711_));
  NOR2X1   g02455(.A(new_n2578_), .B(new_n2574_), .Y(new_n2712_));
  AOI21X1  g02456(.A0(new_n2579_), .A1(new_n2529_), .B0(new_n2712_), .Y(new_n2713_));
  XOR2X1   g02457(.A(new_n2713_), .B(new_n2711_), .Y(new_n2714_));
  AOI22X1  g02458(.A0(new_n818_), .A1(\b[22] ), .B0(new_n817_), .B1(\b[21] ), .Y(new_n2715_));
  OAI21X1  g02459(.A0(new_n816_), .A1(new_n1297_), .B0(new_n2715_), .Y(new_n2716_));
  AOI21X1  g02460(.A0(new_n1399_), .A1(new_n668_), .B0(new_n2716_), .Y(new_n2717_));
  XOR2X1   g02461(.A(new_n2717_), .B(\a[14] ), .Y(new_n2718_));
  XOR2X1   g02462(.A(new_n2718_), .B(new_n2714_), .Y(new_n2719_));
  INVX1    g02463(.A(new_n2584_), .Y(new_n2720_));
  AND2X1   g02464(.A(new_n2720_), .B(new_n2580_), .Y(new_n2721_));
  XOR2X1   g02465(.A(new_n2720_), .B(new_n2580_), .Y(new_n2722_));
  AOI21X1  g02466(.A0(new_n2722_), .A1(new_n2526_), .B0(new_n2721_), .Y(new_n2723_));
  XOR2X1   g02467(.A(new_n2723_), .B(new_n2719_), .Y(new_n2724_));
  AOI22X1  g02468(.A0(new_n603_), .A1(\b[25] ), .B0(new_n602_), .B1(\b[24] ), .Y(new_n2725_));
  OAI21X1  g02469(.A0(new_n601_), .A1(new_n1591_), .B0(new_n2725_), .Y(new_n2726_));
  AOI21X1  g02470(.A0(new_n1590_), .A1(new_n518_), .B0(new_n2726_), .Y(new_n2727_));
  XOR2X1   g02471(.A(new_n2727_), .B(\a[11] ), .Y(new_n2728_));
  NAND2X1  g02472(.A(new_n2728_), .B(new_n2724_), .Y(new_n2729_));
  NOR2X1   g02473(.A(new_n2728_), .B(new_n2724_), .Y(new_n2730_));
  AND2X1   g02474(.A(new_n2728_), .B(new_n2724_), .Y(new_n2731_));
  OR2X1    g02475(.A(new_n2731_), .B(new_n2730_), .Y(new_n2732_));
  AOI21X1  g02476(.A0(new_n2729_), .A1(new_n2632_), .B0(new_n2730_), .Y(new_n2733_));
  AOI22X1  g02477(.A0(new_n2733_), .A1(new_n2729_), .B0(new_n2732_), .B1(new_n2632_), .Y(new_n2734_));
  AOI22X1  g02478(.A0(new_n469_), .A1(\b[28] ), .B0(new_n468_), .B1(\b[27] ), .Y(new_n2735_));
  OAI21X1  g02479(.A0(new_n467_), .A1(new_n1877_), .B0(new_n2735_), .Y(new_n2736_));
  AOI21X1  g02480(.A0(new_n2004_), .A1(new_n404_), .B0(new_n2736_), .Y(new_n2737_));
  XOR2X1   g02481(.A(new_n2737_), .B(\a[8] ), .Y(new_n2738_));
  XOR2X1   g02482(.A(new_n2738_), .B(new_n2734_), .Y(new_n2739_));
  NOR2X1   g02483(.A(new_n2596_), .B(new_n2592_), .Y(new_n2740_));
  OR2X1    g02484(.A(new_n2470_), .B(new_n2466_), .Y(new_n2741_));
  XOR2X1   g02485(.A(new_n2465_), .B(new_n2518_), .Y(new_n2742_));
  XOR2X1   g02486(.A(new_n2470_), .B(new_n2742_), .Y(new_n2743_));
  OAI21X1  g02487(.A0(new_n2481_), .A1(new_n2743_), .B0(new_n2741_), .Y(new_n2744_));
  AOI21X1  g02488(.A0(new_n2744_), .A1(new_n2626_), .B0(new_n2740_), .Y(new_n2745_));
  XOR2X1   g02489(.A(new_n2745_), .B(new_n2739_), .Y(new_n2746_));
  AOI22X1  g02490(.A0(new_n369_), .A1(\b[31] ), .B0(new_n368_), .B1(\b[30] ), .Y(new_n2747_));
  OAI21X1  g02491(.A0(new_n367_), .A1(new_n2359_), .B0(new_n2747_), .Y(new_n2748_));
  AOI21X1  g02492(.A0(new_n2358_), .A1(new_n308_), .B0(new_n2748_), .Y(new_n2749_));
  XOR2X1   g02493(.A(new_n2749_), .B(\a[5] ), .Y(new_n2750_));
  NOR2X1   g02494(.A(new_n2750_), .B(new_n2746_), .Y(new_n2751_));
  AND2X1   g02495(.A(new_n2750_), .B(new_n2746_), .Y(new_n2752_));
  OR2X1    g02496(.A(new_n2752_), .B(new_n2751_), .Y(new_n2753_));
  AND2X1   g02497(.A(new_n2753_), .B(new_n2629_), .Y(new_n2754_));
  NOR3X1   g02498(.A(new_n2752_), .B(new_n2751_), .C(new_n2629_), .Y(new_n2755_));
  NAND2X1  g02499(.A(\b[33] ), .B(\b[32] ), .Y(new_n2756_));
  OAI21X1  g02500(.A0(new_n2613_), .A1(new_n2611_), .B0(new_n2756_), .Y(new_n2757_));
  XOR2X1   g02501(.A(\b[34] ), .B(\b[33] ), .Y(new_n2758_));
  XOR2X1   g02502(.A(new_n2758_), .B(new_n2757_), .Y(new_n2759_));
  AOI22X1  g02503(.A0(new_n267_), .A1(\b[34] ), .B0(new_n266_), .B1(\b[33] ), .Y(new_n2760_));
  OAI21X1  g02504(.A0(new_n350_), .A1(new_n2612_), .B0(new_n2760_), .Y(new_n2761_));
  AOI21X1  g02505(.A0(new_n2759_), .A1(new_n318_), .B0(new_n2761_), .Y(new_n2762_));
  XOR2X1   g02506(.A(new_n2762_), .B(\a[2] ), .Y(new_n2763_));
  OAI21X1  g02507(.A0(new_n2755_), .A1(new_n2754_), .B0(new_n2763_), .Y(new_n2764_));
  NAND2X1  g02508(.A(new_n2753_), .B(new_n2629_), .Y(new_n2765_));
  NOR2X1   g02509(.A(new_n2607_), .B(new_n2627_), .Y(new_n2766_));
  XOR2X1   g02510(.A(new_n2607_), .B(new_n2627_), .Y(new_n2767_));
  AOI21X1  g02511(.A0(new_n2767_), .A1(new_n2516_), .B0(new_n2766_), .Y(new_n2768_));
  OR2X1    g02512(.A(new_n2750_), .B(new_n2746_), .Y(new_n2769_));
  NAND2X1  g02513(.A(new_n2750_), .B(new_n2746_), .Y(new_n2770_));
  NAND3X1  g02514(.A(new_n2770_), .B(new_n2769_), .C(new_n2768_), .Y(new_n2771_));
  XOR2X1   g02515(.A(new_n2762_), .B(new_n257_), .Y(new_n2772_));
  NAND3X1  g02516(.A(new_n2772_), .B(new_n2771_), .C(new_n2765_), .Y(new_n2773_));
  AND2X1   g02517(.A(new_n2773_), .B(new_n2764_), .Y(new_n2774_));
  XOR2X1   g02518(.A(new_n2774_), .B(new_n2624_), .Y(\f[34] ));
  AOI22X1  g02519(.A0(new_n2773_), .A1(new_n2764_), .B0(new_n2623_), .B1(new_n2622_), .Y(new_n2776_));
  AOI21X1  g02520(.A0(new_n2771_), .A1(new_n2765_), .B0(new_n2763_), .Y(new_n2777_));
  AOI21X1  g02521(.A0(new_n2770_), .A1(new_n2629_), .B0(new_n2751_), .Y(new_n2778_));
  AOI22X1  g02522(.A0(new_n603_), .A1(\b[26] ), .B0(new_n602_), .B1(\b[25] ), .Y(new_n2779_));
  OAI21X1  g02523(.A0(new_n601_), .A1(new_n1588_), .B0(new_n2779_), .Y(new_n2780_));
  AOI21X1  g02524(.A0(new_n1783_), .A1(new_n518_), .B0(new_n2780_), .Y(new_n2781_));
  XOR2X1   g02525(.A(new_n2781_), .B(new_n515_), .Y(new_n2782_));
  OR2X1    g02526(.A(new_n2718_), .B(new_n2714_), .Y(new_n2783_));
  AND2X1   g02527(.A(new_n2676_), .B(new_n2672_), .Y(new_n2784_));
  OR2X1    g02528(.A(new_n2676_), .B(new_n2672_), .Y(new_n2785_));
  OAI21X1  g02529(.A0(new_n2784_), .A1(new_n2682_), .B0(new_n2785_), .Y(new_n2786_));
  OAI22X1  g02530(.A0(new_n2786_), .A1(new_n2784_), .B0(new_n2683_), .B1(new_n2682_), .Y(new_n2787_));
  XOR2X1   g02531(.A(new_n2694_), .B(new_n2787_), .Y(new_n2788_));
  XOR2X1   g02532(.A(new_n2705_), .B(new_n2788_), .Y(new_n2789_));
  XOR2X1   g02533(.A(new_n2710_), .B(new_n2789_), .Y(new_n2790_));
  XOR2X1   g02534(.A(new_n2713_), .B(new_n2790_), .Y(new_n2791_));
  XOR2X1   g02535(.A(new_n2718_), .B(new_n2791_), .Y(new_n2792_));
  OAI21X1  g02536(.A0(new_n2723_), .A1(new_n2792_), .B0(new_n2783_), .Y(new_n2793_));
  OR2X1    g02537(.A(new_n2710_), .B(new_n2706_), .Y(new_n2794_));
  OAI21X1  g02538(.A0(new_n2713_), .A1(new_n2790_), .B0(new_n2794_), .Y(new_n2795_));
  OR2X1    g02539(.A(new_n2667_), .B(new_n2663_), .Y(new_n2796_));
  INVX1    g02540(.A(new_n2668_), .Y(new_n2797_));
  OAI21X1  g02541(.A0(new_n2671_), .A1(new_n2797_), .B0(new_n2796_), .Y(new_n2798_));
  AOI22X1  g02542(.A0(new_n1814_), .A1(\b[11] ), .B0(new_n1813_), .B1(\b[10] ), .Y(new_n2799_));
  OAI21X1  g02543(.A0(new_n1812_), .A1(new_n590_), .B0(new_n2799_), .Y(new_n2800_));
  AOI21X1  g02544(.A0(new_n1617_), .A1(new_n589_), .B0(new_n2800_), .Y(new_n2801_));
  XOR2X1   g02545(.A(new_n2801_), .B(\a[26] ), .Y(new_n2802_));
  NAND2X1  g02546(.A(new_n2661_), .B(new_n2640_), .Y(new_n2803_));
  AND2X1   g02547(.A(new_n2635_), .B(new_n2415_), .Y(new_n2804_));
  OAI21X1  g02548(.A0(new_n2804_), .A1(new_n2634_), .B0(new_n2662_), .Y(new_n2805_));
  AND2X1   g02549(.A(new_n2805_), .B(new_n2803_), .Y(new_n2806_));
  AND2X1   g02550(.A(new_n2659_), .B(new_n2647_), .Y(new_n2807_));
  AOI21X1  g02551(.A0(new_n2660_), .A1(new_n2642_), .B0(new_n2807_), .Y(new_n2808_));
  NAND3X1  g02552(.A(new_n2657_), .B(new_n2540_), .C(\a[35] ), .Y(new_n2809_));
  NAND2X1  g02553(.A(new_n2652_), .B(new_n341_), .Y(new_n2810_));
  OR4X1    g02554(.A(new_n2653_), .B(new_n2651_), .C(new_n2539_), .D(new_n274_), .Y(new_n2811_));
  AND2X1   g02555(.A(new_n2653_), .B(new_n2649_), .Y(new_n2812_));
  AND2X1   g02556(.A(new_n2651_), .B(new_n2539_), .Y(new_n2813_));
  AOI22X1  g02557(.A0(new_n2813_), .A1(\b[2] ), .B0(new_n2812_), .B1(\b[1] ), .Y(new_n2814_));
  NAND3X1  g02558(.A(new_n2814_), .B(new_n2811_), .C(new_n2810_), .Y(new_n2815_));
  XOR2X1   g02559(.A(new_n2815_), .B(new_n2650_), .Y(new_n2816_));
  XOR2X1   g02560(.A(new_n2816_), .B(new_n2809_), .Y(new_n2817_));
  INVX1    g02561(.A(new_n2817_), .Y(new_n2818_));
  AOI22X1  g02562(.A0(new_n2545_), .A1(\b[5] ), .B0(new_n2544_), .B1(\b[4] ), .Y(new_n2819_));
  OAI21X1  g02563(.A0(new_n2543_), .A1(new_n297_), .B0(new_n2819_), .Y(new_n2820_));
  AOI21X1  g02564(.A0(new_n2260_), .A1(new_n349_), .B0(new_n2820_), .Y(new_n2821_));
  XOR2X1   g02565(.A(new_n2821_), .B(\a[32] ), .Y(new_n2822_));
  AND2X1   g02566(.A(new_n2822_), .B(new_n2818_), .Y(new_n2823_));
  XOR2X1   g02567(.A(new_n2822_), .B(new_n2818_), .Y(new_n2824_));
  NOR2X1   g02568(.A(new_n2822_), .B(new_n2818_), .Y(new_n2825_));
  INVX1    g02569(.A(new_n2825_), .Y(new_n2826_));
  OAI21X1  g02570(.A0(new_n2823_), .A1(new_n2808_), .B0(new_n2826_), .Y(new_n2827_));
  OAI22X1  g02571(.A0(new_n2827_), .A1(new_n2823_), .B0(new_n2824_), .B1(new_n2808_), .Y(new_n2828_));
  AOI22X1  g02572(.A0(new_n2163_), .A1(\b[8] ), .B0(new_n2162_), .B1(\b[7] ), .Y(new_n2829_));
  OAI21X1  g02573(.A0(new_n2161_), .A1(new_n392_), .B0(new_n2829_), .Y(new_n2830_));
  AOI21X1  g02574(.A0(new_n1907_), .A1(new_n454_), .B0(new_n2830_), .Y(new_n2831_));
  XOR2X1   g02575(.A(new_n2831_), .B(\a[29] ), .Y(new_n2832_));
  XOR2X1   g02576(.A(new_n2832_), .B(new_n2828_), .Y(new_n2833_));
  XOR2X1   g02577(.A(new_n2833_), .B(new_n2806_), .Y(new_n2834_));
  XOR2X1   g02578(.A(new_n2834_), .B(new_n2802_), .Y(new_n2835_));
  XOR2X1   g02579(.A(new_n2835_), .B(new_n2798_), .Y(new_n2836_));
  AOI22X1  g02580(.A0(new_n1526_), .A1(\b[14] ), .B0(new_n1525_), .B1(\b[13] ), .Y(new_n2837_));
  OAI21X1  g02581(.A0(new_n1524_), .A1(new_n713_), .B0(new_n2837_), .Y(new_n2838_));
  AOI21X1  g02582(.A0(new_n1347_), .A1(new_n734_), .B0(new_n2838_), .Y(new_n2839_));
  XOR2X1   g02583(.A(new_n2839_), .B(\a[23] ), .Y(new_n2840_));
  XOR2X1   g02584(.A(new_n2840_), .B(new_n2836_), .Y(new_n2841_));
  XOR2X1   g02585(.A(new_n2841_), .B(new_n2786_), .Y(new_n2842_));
  AOI22X1  g02586(.A0(new_n1263_), .A1(\b[17] ), .B0(new_n1262_), .B1(\b[16] ), .Y(new_n2843_));
  OAI21X1  g02587(.A0(new_n1261_), .A1(new_n977_), .B0(new_n2843_), .Y(new_n2844_));
  AOI21X1  g02588(.A0(new_n1075_), .A1(new_n976_), .B0(new_n2844_), .Y(new_n2845_));
  XOR2X1   g02589(.A(new_n2845_), .B(\a[20] ), .Y(new_n2846_));
  XOR2X1   g02590(.A(new_n2846_), .B(new_n2842_), .Y(new_n2847_));
  OR2X1    g02591(.A(new_n2694_), .B(new_n2690_), .Y(new_n2848_));
  OAI21X1  g02592(.A0(new_n2705_), .A1(new_n2788_), .B0(new_n2848_), .Y(new_n2849_));
  XOR2X1   g02593(.A(new_n2849_), .B(new_n2847_), .Y(new_n2850_));
  AOI22X1  g02594(.A0(new_n1017_), .A1(\b[20] ), .B0(new_n1016_), .B1(\b[19] ), .Y(new_n2851_));
  OAI21X1  g02595(.A0(new_n1015_), .A1(new_n1115_), .B0(new_n2851_), .Y(new_n2852_));
  AOI21X1  g02596(.A0(new_n1217_), .A1(new_n882_), .B0(new_n2852_), .Y(new_n2853_));
  XOR2X1   g02597(.A(new_n2853_), .B(\a[17] ), .Y(new_n2854_));
  NAND2X1  g02598(.A(new_n2854_), .B(new_n2850_), .Y(new_n2855_));
  OR2X1    g02599(.A(new_n2854_), .B(new_n2850_), .Y(new_n2856_));
  NAND3X1  g02600(.A(new_n2855_), .B(new_n2856_), .C(new_n2795_), .Y(new_n2857_));
  NOR2X1   g02601(.A(new_n2854_), .B(new_n2850_), .Y(new_n2858_));
  AOI21X1  g02602(.A0(new_n2855_), .A1(new_n2795_), .B0(new_n2858_), .Y(new_n2859_));
  AOI22X1  g02603(.A0(new_n2859_), .A1(new_n2855_), .B0(new_n2857_), .B1(new_n2795_), .Y(new_n2860_));
  AOI22X1  g02604(.A0(new_n818_), .A1(\b[23] ), .B0(new_n817_), .B1(\b[22] ), .Y(new_n2861_));
  OAI21X1  g02605(.A0(new_n816_), .A1(new_n1482_), .B0(new_n2861_), .Y(new_n2862_));
  AOI21X1  g02606(.A0(new_n1481_), .A1(new_n668_), .B0(new_n2862_), .Y(new_n2863_));
  XOR2X1   g02607(.A(new_n2863_), .B(\a[14] ), .Y(new_n2864_));
  XOR2X1   g02608(.A(new_n2864_), .B(new_n2860_), .Y(new_n2865_));
  XOR2X1   g02609(.A(new_n2865_), .B(new_n2793_), .Y(new_n2866_));
  XOR2X1   g02610(.A(new_n2866_), .B(new_n2782_), .Y(new_n2867_));
  XOR2X1   g02611(.A(new_n2867_), .B(new_n2733_), .Y(new_n2868_));
  AOI22X1  g02612(.A0(new_n469_), .A1(\b[29] ), .B0(new_n468_), .B1(\b[28] ), .Y(new_n2869_));
  OAI21X1  g02613(.A0(new_n467_), .A1(new_n2126_), .B0(new_n2869_), .Y(new_n2870_));
  AOI21X1  g02614(.A0(new_n2125_), .A1(new_n404_), .B0(new_n2870_), .Y(new_n2871_));
  XOR2X1   g02615(.A(new_n2871_), .B(\a[8] ), .Y(new_n2872_));
  XOR2X1   g02616(.A(new_n2872_), .B(new_n2868_), .Y(new_n2873_));
  NOR2X1   g02617(.A(new_n2738_), .B(new_n2734_), .Y(new_n2874_));
  OR2X1    g02618(.A(new_n2596_), .B(new_n2592_), .Y(new_n2875_));
  OAI21X1  g02619(.A0(new_n2602_), .A1(new_n2598_), .B0(new_n2875_), .Y(new_n2876_));
  AOI21X1  g02620(.A0(new_n2876_), .A1(new_n2739_), .B0(new_n2874_), .Y(new_n2877_));
  XOR2X1   g02621(.A(new_n2877_), .B(new_n2873_), .Y(new_n2878_));
  AOI22X1  g02622(.A0(new_n369_), .A1(\b[32] ), .B0(new_n368_), .B1(\b[31] ), .Y(new_n2879_));
  OAI21X1  g02623(.A0(new_n367_), .A1(new_n2356_), .B0(new_n2879_), .Y(new_n2880_));
  AOI21X1  g02624(.A0(new_n2495_), .A1(new_n308_), .B0(new_n2880_), .Y(new_n2881_));
  XOR2X1   g02625(.A(new_n2881_), .B(\a[5] ), .Y(new_n2882_));
  XOR2X1   g02626(.A(new_n2882_), .B(new_n2878_), .Y(new_n2883_));
  OR2X1    g02627(.A(new_n2883_), .B(new_n2778_), .Y(new_n2884_));
  OR2X1    g02628(.A(new_n2882_), .B(new_n2878_), .Y(new_n2885_));
  NAND2X1  g02629(.A(new_n2882_), .B(new_n2878_), .Y(new_n2886_));
  NAND3X1  g02630(.A(new_n2886_), .B(new_n2885_), .C(new_n2778_), .Y(new_n2887_));
  AND2X1   g02631(.A(\b[34] ), .B(\b[33] ), .Y(new_n2888_));
  AOI21X1  g02632(.A0(new_n2758_), .A1(new_n2757_), .B0(new_n2888_), .Y(new_n2889_));
  INVX1    g02633(.A(\b[34] ), .Y(new_n2890_));
  XOR2X1   g02634(.A(\b[35] ), .B(new_n2890_), .Y(new_n2891_));
  XOR2X1   g02635(.A(new_n2891_), .B(new_n2889_), .Y(new_n2892_));
  INVX1    g02636(.A(\b[33] ), .Y(new_n2893_));
  AOI22X1  g02637(.A0(new_n267_), .A1(\b[35] ), .B0(new_n266_), .B1(\b[34] ), .Y(new_n2894_));
  OAI21X1  g02638(.A0(new_n350_), .A1(new_n2893_), .B0(new_n2894_), .Y(new_n2895_));
  AOI21X1  g02639(.A0(new_n2892_), .A1(new_n318_), .B0(new_n2895_), .Y(new_n2896_));
  XOR2X1   g02640(.A(new_n2896_), .B(new_n257_), .Y(new_n2897_));
  AOI21X1  g02641(.A0(new_n2887_), .A1(new_n2884_), .B0(new_n2897_), .Y(new_n2898_));
  NOR2X1   g02642(.A(new_n2883_), .B(new_n2778_), .Y(new_n2899_));
  OAI21X1  g02643(.A0(new_n2752_), .A1(new_n2768_), .B0(new_n2769_), .Y(new_n2900_));
  NOR2X1   g02644(.A(new_n2882_), .B(new_n2878_), .Y(new_n2901_));
  AND2X1   g02645(.A(new_n2882_), .B(new_n2878_), .Y(new_n2902_));
  NOR3X1   g02646(.A(new_n2902_), .B(new_n2901_), .C(new_n2900_), .Y(new_n2903_));
  XOR2X1   g02647(.A(new_n2896_), .B(\a[2] ), .Y(new_n2904_));
  NOR3X1   g02648(.A(new_n2904_), .B(new_n2903_), .C(new_n2899_), .Y(new_n2905_));
  OAI22X1  g02649(.A0(new_n2905_), .A1(new_n2898_), .B0(new_n2777_), .B1(new_n2776_), .Y(new_n2906_));
  OR4X1    g02650(.A(new_n2905_), .B(new_n2898_), .C(new_n2777_), .D(new_n2776_), .Y(new_n2907_));
  AND2X1   g02651(.A(new_n2907_), .B(new_n2906_), .Y(\f[35] ));
  OAI21X1  g02652(.A0(new_n2902_), .A1(new_n2778_), .B0(new_n2885_), .Y(new_n2909_));
  AOI22X1  g02653(.A0(new_n369_), .A1(\b[33] ), .B0(new_n368_), .B1(\b[32] ), .Y(new_n2910_));
  OAI21X1  g02654(.A0(new_n367_), .A1(new_n2615_), .B0(new_n2910_), .Y(new_n2911_));
  AOI21X1  g02655(.A0(new_n2614_), .A1(new_n308_), .B0(new_n2911_), .Y(new_n2912_));
  XOR2X1   g02656(.A(new_n2912_), .B(new_n305_), .Y(new_n2913_));
  OR2X1    g02657(.A(new_n2872_), .B(new_n2868_), .Y(new_n2914_));
  AND2X1   g02658(.A(new_n2464_), .B(new_n2460_), .Y(new_n2915_));
  OR2X1    g02659(.A(new_n2464_), .B(new_n2460_), .Y(new_n2916_));
  OAI21X1  g02660(.A0(new_n2915_), .A1(new_n2388_), .B0(new_n2916_), .Y(new_n2917_));
  NOR2X1   g02661(.A(new_n2590_), .B(new_n2586_), .Y(new_n2918_));
  AOI21X1  g02662(.A0(new_n2591_), .A1(new_n2917_), .B0(new_n2918_), .Y(new_n2919_));
  OR2X1    g02663(.A(new_n2728_), .B(new_n2724_), .Y(new_n2920_));
  OAI21X1  g02664(.A0(new_n2731_), .A1(new_n2919_), .B0(new_n2920_), .Y(new_n2921_));
  XOR2X1   g02665(.A(new_n2867_), .B(new_n2921_), .Y(new_n2922_));
  XOR2X1   g02666(.A(new_n2872_), .B(new_n2922_), .Y(new_n2923_));
  OAI21X1  g02667(.A0(new_n2877_), .A1(new_n2923_), .B0(new_n2914_), .Y(new_n2924_));
  NAND2X1  g02668(.A(new_n2866_), .B(new_n2782_), .Y(new_n2925_));
  NAND2X1  g02669(.A(new_n2867_), .B(new_n2921_), .Y(new_n2926_));
  NAND2X1  g02670(.A(new_n2926_), .B(new_n2925_), .Y(new_n2927_));
  NOR2X1   g02671(.A(new_n2864_), .B(new_n2860_), .Y(new_n2928_));
  AOI21X1  g02672(.A0(new_n2865_), .A1(new_n2793_), .B0(new_n2928_), .Y(new_n2929_));
  XOR2X1   g02673(.A(new_n2841_), .B(new_n2689_), .Y(new_n2930_));
  NOR2X1   g02674(.A(new_n2846_), .B(new_n2930_), .Y(new_n2931_));
  XOR2X1   g02675(.A(new_n2846_), .B(new_n2930_), .Y(new_n2932_));
  AOI21X1  g02676(.A0(new_n2849_), .A1(new_n2932_), .B0(new_n2931_), .Y(new_n2933_));
  OR2X1    g02677(.A(new_n2840_), .B(new_n2836_), .Y(new_n2934_));
  NAND2X1  g02678(.A(new_n2841_), .B(new_n2786_), .Y(new_n2935_));
  NAND2X1  g02679(.A(new_n2935_), .B(new_n2934_), .Y(new_n2936_));
  XOR2X1   g02680(.A(new_n2831_), .B(new_n1911_), .Y(new_n2937_));
  NAND2X1  g02681(.A(new_n2937_), .B(new_n2828_), .Y(new_n2938_));
  OAI21X1  g02682(.A0(new_n2833_), .A1(new_n2806_), .B0(new_n2938_), .Y(new_n2939_));
  OR2X1    g02683(.A(new_n2816_), .B(new_n2809_), .Y(new_n2940_));
  XOR2X1   g02684(.A(\a[36] ), .B(\a[35] ), .Y(new_n2941_));
  NAND2X1  g02685(.A(new_n2941_), .B(\b[0] ), .Y(new_n2942_));
  INVX1    g02686(.A(new_n2942_), .Y(new_n2943_));
  XOR2X1   g02687(.A(new_n2943_), .B(new_n2940_), .Y(new_n2944_));
  OR2X1    g02688(.A(new_n2653_), .B(new_n2539_), .Y(new_n2945_));
  OR2X1    g02689(.A(new_n2945_), .B(new_n2651_), .Y(new_n2946_));
  AOI22X1  g02690(.A0(new_n2813_), .A1(\b[3] ), .B0(new_n2812_), .B1(\b[2] ), .Y(new_n2947_));
  OAI21X1  g02691(.A0(new_n2946_), .A1(new_n275_), .B0(new_n2947_), .Y(new_n2948_));
  AOI21X1  g02692(.A0(new_n2652_), .A1(new_n366_), .B0(new_n2948_), .Y(new_n2949_));
  XOR2X1   g02693(.A(new_n2949_), .B(\a[35] ), .Y(new_n2950_));
  XOR2X1   g02694(.A(new_n2950_), .B(new_n2944_), .Y(new_n2951_));
  AOI22X1  g02695(.A0(new_n2545_), .A1(\b[6] ), .B0(new_n2544_), .B1(\b[5] ), .Y(new_n2952_));
  OAI21X1  g02696(.A0(new_n2543_), .A1(new_n325_), .B0(new_n2952_), .Y(new_n2953_));
  AOI21X1  g02697(.A0(new_n2260_), .A1(new_n378_), .B0(new_n2953_), .Y(new_n2954_));
  XOR2X1   g02698(.A(new_n2954_), .B(\a[32] ), .Y(new_n2955_));
  XOR2X1   g02699(.A(new_n2955_), .B(new_n2951_), .Y(new_n2956_));
  XOR2X1   g02700(.A(new_n2956_), .B(new_n2827_), .Y(new_n2957_));
  AOI22X1  g02701(.A0(new_n2163_), .A1(\b[9] ), .B0(new_n2162_), .B1(\b[8] ), .Y(new_n2958_));
  OAI21X1  g02702(.A0(new_n2161_), .A1(new_n492_), .B0(new_n2958_), .Y(new_n2959_));
  AOI21X1  g02703(.A0(new_n1907_), .A1(new_n491_), .B0(new_n2959_), .Y(new_n2960_));
  XOR2X1   g02704(.A(new_n2960_), .B(\a[29] ), .Y(new_n2961_));
  XOR2X1   g02705(.A(new_n2961_), .B(new_n2957_), .Y(new_n2962_));
  XOR2X1   g02706(.A(new_n2962_), .B(new_n2939_), .Y(new_n2963_));
  AOI22X1  g02707(.A0(new_n1814_), .A1(\b[12] ), .B0(new_n1813_), .B1(\b[11] ), .Y(new_n2964_));
  OAI21X1  g02708(.A0(new_n1812_), .A1(new_n587_), .B0(new_n2964_), .Y(new_n2965_));
  AOI21X1  g02709(.A0(new_n1617_), .A1(new_n635_), .B0(new_n2965_), .Y(new_n2966_));
  XOR2X1   g02710(.A(new_n2966_), .B(\a[26] ), .Y(new_n2967_));
  XOR2X1   g02711(.A(new_n2967_), .B(new_n2963_), .Y(new_n2968_));
  INVX1    g02712(.A(new_n2802_), .Y(new_n2969_));
  AND2X1   g02713(.A(new_n2834_), .B(new_n2969_), .Y(new_n2970_));
  XOR2X1   g02714(.A(new_n2834_), .B(new_n2969_), .Y(new_n2971_));
  AOI21X1  g02715(.A0(new_n2971_), .A1(new_n2798_), .B0(new_n2970_), .Y(new_n2972_));
  XOR2X1   g02716(.A(new_n2972_), .B(new_n2968_), .Y(new_n2973_));
  AOI22X1  g02717(.A0(new_n1526_), .A1(\b[15] ), .B0(new_n1525_), .B1(\b[14] ), .Y(new_n2974_));
  OAI21X1  g02718(.A0(new_n1524_), .A1(new_n795_), .B0(new_n2974_), .Y(new_n2975_));
  AOI21X1  g02719(.A0(new_n1347_), .A1(new_n794_), .B0(new_n2975_), .Y(new_n2976_));
  XOR2X1   g02720(.A(new_n2976_), .B(\a[23] ), .Y(new_n2977_));
  XOR2X1   g02721(.A(new_n2977_), .B(new_n2973_), .Y(new_n2978_));
  XOR2X1   g02722(.A(new_n2978_), .B(new_n2936_), .Y(new_n2979_));
  AOI22X1  g02723(.A0(new_n1263_), .A1(\b[18] ), .B0(new_n1262_), .B1(\b[17] ), .Y(new_n2980_));
  OAI21X1  g02724(.A0(new_n1261_), .A1(new_n974_), .B0(new_n2980_), .Y(new_n2981_));
  AOI21X1  g02725(.A0(new_n1075_), .A1(new_n1042_), .B0(new_n2981_), .Y(new_n2982_));
  XOR2X1   g02726(.A(new_n2982_), .B(new_n1072_), .Y(new_n2983_));
  XOR2X1   g02727(.A(new_n2983_), .B(new_n2979_), .Y(new_n2984_));
  XOR2X1   g02728(.A(new_n2984_), .B(new_n2933_), .Y(new_n2985_));
  AOI22X1  g02729(.A0(new_n1017_), .A1(\b[21] ), .B0(new_n1016_), .B1(\b[20] ), .Y(new_n2986_));
  OAI21X1  g02730(.A0(new_n1015_), .A1(new_n1300_), .B0(new_n2986_), .Y(new_n2987_));
  AOI21X1  g02731(.A0(new_n1299_), .A1(new_n882_), .B0(new_n2987_), .Y(new_n2988_));
  XOR2X1   g02732(.A(new_n2988_), .B(\a[17] ), .Y(new_n2989_));
  XOR2X1   g02733(.A(new_n2989_), .B(new_n2985_), .Y(new_n2990_));
  XOR2X1   g02734(.A(new_n2990_), .B(new_n2859_), .Y(new_n2991_));
  AOI22X1  g02735(.A0(new_n818_), .A1(\b[24] ), .B0(new_n817_), .B1(\b[23] ), .Y(new_n2992_));
  OAI21X1  g02736(.A0(new_n816_), .A1(new_n1479_), .B0(new_n2992_), .Y(new_n2993_));
  AOI21X1  g02737(.A0(new_n1572_), .A1(new_n668_), .B0(new_n2993_), .Y(new_n2994_));
  XOR2X1   g02738(.A(new_n2994_), .B(\a[14] ), .Y(new_n2995_));
  XOR2X1   g02739(.A(new_n2995_), .B(new_n2991_), .Y(new_n2996_));
  XOR2X1   g02740(.A(new_n2996_), .B(new_n2929_), .Y(new_n2997_));
  AOI22X1  g02741(.A0(new_n603_), .A1(\b[27] ), .B0(new_n602_), .B1(\b[26] ), .Y(new_n2998_));
  OAI21X1  g02742(.A0(new_n601_), .A1(new_n1880_), .B0(new_n2998_), .Y(new_n2999_));
  AOI21X1  g02743(.A0(new_n1879_), .A1(new_n518_), .B0(new_n2999_), .Y(new_n3000_));
  XOR2X1   g02744(.A(new_n3000_), .B(\a[11] ), .Y(new_n3001_));
  XOR2X1   g02745(.A(new_n3001_), .B(new_n2997_), .Y(new_n3002_));
  XOR2X1   g02746(.A(new_n3002_), .B(new_n2927_), .Y(new_n3003_));
  AOI22X1  g02747(.A0(new_n469_), .A1(\b[30] ), .B0(new_n468_), .B1(\b[29] ), .Y(new_n3004_));
  OAI21X1  g02748(.A0(new_n467_), .A1(new_n2231_), .B0(new_n3004_), .Y(new_n3005_));
  AOI21X1  g02749(.A0(new_n2230_), .A1(new_n404_), .B0(new_n3005_), .Y(new_n3006_));
  XOR2X1   g02750(.A(new_n3006_), .B(\a[8] ), .Y(new_n3007_));
  XOR2X1   g02751(.A(new_n3007_), .B(new_n3003_), .Y(new_n3008_));
  XOR2X1   g02752(.A(new_n3008_), .B(new_n2924_), .Y(new_n3009_));
  XOR2X1   g02753(.A(new_n3009_), .B(new_n2913_), .Y(new_n3010_));
  XOR2X1   g02754(.A(new_n3010_), .B(new_n2909_), .Y(new_n3011_));
  NAND2X1  g02755(.A(\b[35] ), .B(\b[34] ), .Y(new_n3012_));
  OAI21X1  g02756(.A0(new_n2891_), .A1(new_n2889_), .B0(new_n3012_), .Y(new_n3013_));
  XOR2X1   g02757(.A(\b[36] ), .B(\b[35] ), .Y(new_n3014_));
  XOR2X1   g02758(.A(new_n3014_), .B(new_n3013_), .Y(new_n3015_));
  AOI22X1  g02759(.A0(new_n267_), .A1(\b[36] ), .B0(new_n266_), .B1(\b[35] ), .Y(new_n3016_));
  OAI21X1  g02760(.A0(new_n350_), .A1(new_n2890_), .B0(new_n3016_), .Y(new_n3017_));
  AOI21X1  g02761(.A0(new_n3015_), .A1(new_n318_), .B0(new_n3017_), .Y(new_n3018_));
  XOR2X1   g02762(.A(new_n3018_), .B(\a[2] ), .Y(new_n3019_));
  XOR2X1   g02763(.A(new_n3019_), .B(new_n3011_), .Y(new_n3020_));
  OAI21X1  g02764(.A0(new_n2903_), .A1(new_n2899_), .B0(new_n2897_), .Y(new_n3021_));
  AND2X1   g02765(.A(new_n3021_), .B(new_n2906_), .Y(new_n3022_));
  XOR2X1   g02766(.A(new_n3022_), .B(new_n3020_), .Y(\f[36] ));
  AOI21X1  g02767(.A0(new_n2886_), .A1(new_n2900_), .B0(new_n2901_), .Y(new_n3024_));
  XOR2X1   g02768(.A(new_n3010_), .B(new_n3024_), .Y(new_n3025_));
  NOR2X1   g02769(.A(new_n3019_), .B(new_n3025_), .Y(new_n3026_));
  AOI21X1  g02770(.A0(new_n3021_), .A1(new_n2906_), .B0(new_n3020_), .Y(new_n3027_));
  OR2X1    g02771(.A(new_n3027_), .B(new_n3026_), .Y(new_n3028_));
  NOR2X1   g02772(.A(new_n3007_), .B(new_n3003_), .Y(new_n3029_));
  AOI21X1  g02773(.A0(new_n3008_), .A1(new_n2924_), .B0(new_n3029_), .Y(new_n3030_));
  AOI22X1  g02774(.A0(new_n469_), .A1(\b[31] ), .B0(new_n468_), .B1(\b[30] ), .Y(new_n3031_));
  OAI21X1  g02775(.A0(new_n467_), .A1(new_n2359_), .B0(new_n3031_), .Y(new_n3032_));
  AOI21X1  g02776(.A0(new_n2358_), .A1(new_n404_), .B0(new_n3032_), .Y(new_n3033_));
  XOR2X1   g02777(.A(new_n3033_), .B(new_n400_), .Y(new_n3034_));
  XOR2X1   g02778(.A(new_n3000_), .B(new_n515_), .Y(new_n3035_));
  AND2X1   g02779(.A(new_n3035_), .B(new_n2997_), .Y(new_n3036_));
  AOI21X1  g02780(.A0(new_n2926_), .A1(new_n2925_), .B0(new_n3002_), .Y(new_n3037_));
  OR2X1    g02781(.A(new_n3037_), .B(new_n3036_), .Y(new_n3038_));
  XOR2X1   g02782(.A(new_n2982_), .B(\a[20] ), .Y(new_n3039_));
  XOR2X1   g02783(.A(new_n3039_), .B(new_n2979_), .Y(new_n3040_));
  XOR2X1   g02784(.A(new_n3040_), .B(new_n2933_), .Y(new_n3041_));
  XOR2X1   g02785(.A(new_n2989_), .B(new_n3041_), .Y(new_n3042_));
  XOR2X1   g02786(.A(new_n3042_), .B(new_n2859_), .Y(new_n3043_));
  OR2X1    g02787(.A(new_n2995_), .B(new_n3043_), .Y(new_n3044_));
  OAI21X1  g02788(.A0(new_n2996_), .A1(new_n2929_), .B0(new_n3044_), .Y(new_n3045_));
  INVX1    g02789(.A(new_n2963_), .Y(new_n3046_));
  OR2X1    g02790(.A(new_n2967_), .B(new_n3046_), .Y(new_n3047_));
  OAI21X1  g02791(.A0(new_n2972_), .A1(new_n2968_), .B0(new_n3047_), .Y(new_n3048_));
  AOI22X1  g02792(.A0(new_n1814_), .A1(\b[13] ), .B0(new_n1813_), .B1(\b[12] ), .Y(new_n3049_));
  OAI21X1  g02793(.A0(new_n1812_), .A1(new_n716_), .B0(new_n3049_), .Y(new_n3050_));
  AOI21X1  g02794(.A0(new_n1617_), .A1(new_n715_), .B0(new_n3050_), .Y(new_n3051_));
  XOR2X1   g02795(.A(new_n3051_), .B(\a[26] ), .Y(new_n3052_));
  INVX1    g02796(.A(new_n3052_), .Y(new_n3053_));
  NOR2X1   g02797(.A(new_n2961_), .B(new_n2957_), .Y(new_n3054_));
  AOI21X1  g02798(.A0(new_n2962_), .A1(new_n2939_), .B0(new_n3054_), .Y(new_n3055_));
  AOI22X1  g02799(.A0(new_n2163_), .A1(\b[10] ), .B0(new_n2162_), .B1(\b[9] ), .Y(new_n3056_));
  OAI21X1  g02800(.A0(new_n2161_), .A1(new_n489_), .B0(new_n3056_), .Y(new_n3057_));
  AOI21X1  g02801(.A0(new_n1907_), .A1(new_n543_), .B0(new_n3057_), .Y(new_n3058_));
  XOR2X1   g02802(.A(new_n3058_), .B(\a[29] ), .Y(new_n3059_));
  INVX1    g02803(.A(new_n3059_), .Y(new_n3060_));
  INVX1    g02804(.A(new_n2827_), .Y(new_n3061_));
  INVX1    g02805(.A(new_n2955_), .Y(new_n3062_));
  NAND2X1  g02806(.A(new_n3062_), .B(new_n2951_), .Y(new_n3063_));
  OAI21X1  g02807(.A0(new_n2956_), .A1(new_n3061_), .B0(new_n3063_), .Y(new_n3064_));
  AOI22X1  g02808(.A0(new_n2545_), .A1(\b[7] ), .B0(new_n2544_), .B1(\b[6] ), .Y(new_n3065_));
  OAI21X1  g02809(.A0(new_n2543_), .A1(new_n395_), .B0(new_n3065_), .Y(new_n3066_));
  AOI21X1  g02810(.A0(new_n2260_), .A1(new_n394_), .B0(new_n3066_), .Y(new_n3067_));
  XOR2X1   g02811(.A(new_n3067_), .B(new_n2258_), .Y(new_n3068_));
  OR4X1    g02812(.A(new_n2942_), .B(new_n2816_), .C(new_n2658_), .D(new_n2648_), .Y(new_n3069_));
  OAI21X1  g02813(.A0(new_n2950_), .A1(new_n2944_), .B0(new_n3069_), .Y(new_n3070_));
  AND2X1   g02814(.A(new_n2652_), .B(new_n323_), .Y(new_n3071_));
  NOR3X1   g02815(.A(new_n2945_), .B(new_n2651_), .C(new_n277_), .Y(new_n3072_));
  OAI22X1  g02816(.A0(new_n2655_), .A1(new_n325_), .B0(new_n2654_), .B1(new_n297_), .Y(new_n3073_));
  NOR3X1   g02817(.A(new_n3073_), .B(new_n3072_), .C(new_n3071_), .Y(new_n3074_));
  XOR2X1   g02818(.A(new_n3074_), .B(new_n2650_), .Y(new_n3075_));
  NAND2X1  g02819(.A(new_n2942_), .B(\a[38] ), .Y(new_n3076_));
  XOR2X1   g02820(.A(\a[36] ), .B(new_n2650_), .Y(new_n3077_));
  INVX1    g02821(.A(\a[38] ), .Y(new_n3078_));
  XOR2X1   g02822(.A(new_n3078_), .B(\a[37] ), .Y(new_n3079_));
  NOR2X1   g02823(.A(new_n3079_), .B(new_n3077_), .Y(new_n3080_));
  XOR2X1   g02824(.A(\a[37] ), .B(\a[36] ), .Y(new_n3081_));
  NAND2X1  g02825(.A(new_n3081_), .B(new_n3077_), .Y(new_n3082_));
  NAND2X1  g02826(.A(new_n3079_), .B(new_n2941_), .Y(new_n3083_));
  OAI22X1  g02827(.A0(new_n3083_), .A1(new_n275_), .B0(new_n3082_), .B1(new_n274_), .Y(new_n3084_));
  AOI21X1  g02828(.A0(new_n3080_), .A1(new_n263_), .B0(new_n3084_), .Y(new_n3085_));
  XOR2X1   g02829(.A(new_n3085_), .B(\a[38] ), .Y(new_n3086_));
  XOR2X1   g02830(.A(new_n3086_), .B(new_n3076_), .Y(new_n3087_));
  XOR2X1   g02831(.A(new_n3087_), .B(new_n3075_), .Y(new_n3088_));
  XOR2X1   g02832(.A(new_n3088_), .B(new_n3070_), .Y(new_n3089_));
  XOR2X1   g02833(.A(new_n3089_), .B(new_n3068_), .Y(new_n3090_));
  XOR2X1   g02834(.A(new_n3090_), .B(new_n3064_), .Y(new_n3091_));
  XOR2X1   g02835(.A(new_n3091_), .B(new_n3060_), .Y(new_n3092_));
  INVX1    g02836(.A(new_n3092_), .Y(new_n3093_));
  XOR2X1   g02837(.A(new_n3093_), .B(new_n3055_), .Y(new_n3094_));
  XOR2X1   g02838(.A(new_n3094_), .B(new_n3053_), .Y(new_n3095_));
  INVX1    g02839(.A(new_n3095_), .Y(new_n3096_));
  XOR2X1   g02840(.A(new_n3096_), .B(new_n3048_), .Y(new_n3097_));
  AOI22X1  g02841(.A0(new_n1526_), .A1(\b[16] ), .B0(new_n1525_), .B1(\b[15] ), .Y(new_n3098_));
  OAI21X1  g02842(.A0(new_n1524_), .A1(new_n792_), .B0(new_n3098_), .Y(new_n3099_));
  AOI21X1  g02843(.A0(new_n1347_), .A1(new_n842_), .B0(new_n3099_), .Y(new_n3100_));
  XOR2X1   g02844(.A(new_n3100_), .B(\a[23] ), .Y(new_n3101_));
  XOR2X1   g02845(.A(new_n3101_), .B(new_n3097_), .Y(new_n3102_));
  XOR2X1   g02846(.A(new_n2976_), .B(new_n1351_), .Y(new_n3103_));
  AND2X1   g02847(.A(new_n3103_), .B(new_n2973_), .Y(new_n3104_));
  AOI21X1  g02848(.A0(new_n2935_), .A1(new_n2934_), .B0(new_n2978_), .Y(new_n3105_));
  NOR2X1   g02849(.A(new_n3105_), .B(new_n3104_), .Y(new_n3106_));
  XOR2X1   g02850(.A(new_n3106_), .B(new_n3102_), .Y(new_n3107_));
  AOI22X1  g02851(.A0(new_n1263_), .A1(\b[19] ), .B0(new_n1262_), .B1(\b[18] ), .Y(new_n3108_));
  OAI21X1  g02852(.A0(new_n1261_), .A1(new_n1118_), .B0(new_n3108_), .Y(new_n3109_));
  AOI21X1  g02853(.A0(new_n1117_), .A1(new_n1075_), .B0(new_n3109_), .Y(new_n3110_));
  XOR2X1   g02854(.A(new_n3110_), .B(new_n1072_), .Y(new_n3111_));
  XOR2X1   g02855(.A(new_n3111_), .B(new_n3107_), .Y(new_n3112_));
  OR2X1    g02856(.A(new_n3039_), .B(new_n2979_), .Y(new_n3113_));
  OAI21X1  g02857(.A0(new_n2984_), .A1(new_n2933_), .B0(new_n3113_), .Y(new_n3114_));
  XOR2X1   g02858(.A(new_n3114_), .B(new_n3112_), .Y(new_n3115_));
  AOI22X1  g02859(.A0(new_n1017_), .A1(\b[22] ), .B0(new_n1016_), .B1(\b[21] ), .Y(new_n3116_));
  OAI21X1  g02860(.A0(new_n1015_), .A1(new_n1297_), .B0(new_n3116_), .Y(new_n3117_));
  AOI21X1  g02861(.A0(new_n1399_), .A1(new_n882_), .B0(new_n3117_), .Y(new_n3118_));
  XOR2X1   g02862(.A(new_n3118_), .B(\a[17] ), .Y(new_n3119_));
  XOR2X1   g02863(.A(new_n3119_), .B(new_n3115_), .Y(new_n3120_));
  OR2X1    g02864(.A(new_n2989_), .B(new_n3041_), .Y(new_n3121_));
  OAI21X1  g02865(.A0(new_n2990_), .A1(new_n2859_), .B0(new_n3121_), .Y(new_n3122_));
  NOR2X1   g02866(.A(new_n3122_), .B(new_n3120_), .Y(new_n3123_));
  AND2X1   g02867(.A(new_n3122_), .B(new_n3120_), .Y(new_n3124_));
  AOI22X1  g02868(.A0(new_n818_), .A1(\b[25] ), .B0(new_n817_), .B1(\b[24] ), .Y(new_n3125_));
  OAI21X1  g02869(.A0(new_n816_), .A1(new_n1591_), .B0(new_n3125_), .Y(new_n3126_));
  AOI21X1  g02870(.A0(new_n1590_), .A1(new_n668_), .B0(new_n3126_), .Y(new_n3127_));
  XOR2X1   g02871(.A(new_n3127_), .B(\a[14] ), .Y(new_n3128_));
  OAI21X1  g02872(.A0(new_n3124_), .A1(new_n3123_), .B0(new_n3128_), .Y(new_n3129_));
  XOR2X1   g02873(.A(new_n3122_), .B(new_n3120_), .Y(new_n3130_));
  XOR2X1   g02874(.A(new_n3128_), .B(new_n3130_), .Y(new_n3131_));
  NOR3X1   g02875(.A(new_n3128_), .B(new_n3124_), .C(new_n3123_), .Y(new_n3132_));
  AOI21X1  g02876(.A0(new_n3129_), .A1(new_n3045_), .B0(new_n3132_), .Y(new_n3133_));
  AOI22X1  g02877(.A0(new_n3133_), .A1(new_n3129_), .B0(new_n3131_), .B1(new_n3045_), .Y(new_n3134_));
  AOI22X1  g02878(.A0(new_n603_), .A1(\b[28] ), .B0(new_n602_), .B1(\b[27] ), .Y(new_n3135_));
  OAI21X1  g02879(.A0(new_n601_), .A1(new_n1877_), .B0(new_n3135_), .Y(new_n3136_));
  AOI21X1  g02880(.A0(new_n2004_), .A1(new_n518_), .B0(new_n3136_), .Y(new_n3137_));
  XOR2X1   g02881(.A(new_n3137_), .B(\a[11] ), .Y(new_n3138_));
  XOR2X1   g02882(.A(new_n3138_), .B(new_n3134_), .Y(new_n3139_));
  XOR2X1   g02883(.A(new_n3139_), .B(new_n3038_), .Y(new_n3140_));
  XOR2X1   g02884(.A(new_n3140_), .B(new_n3034_), .Y(new_n3141_));
  XOR2X1   g02885(.A(new_n3141_), .B(new_n3030_), .Y(new_n3142_));
  AOI22X1  g02886(.A0(new_n369_), .A1(\b[34] ), .B0(new_n368_), .B1(\b[33] ), .Y(new_n3143_));
  OAI21X1  g02887(.A0(new_n367_), .A1(new_n2612_), .B0(new_n3143_), .Y(new_n3144_));
  AOI21X1  g02888(.A0(new_n2759_), .A1(new_n308_), .B0(new_n3144_), .Y(new_n3145_));
  XOR2X1   g02889(.A(new_n3145_), .B(\a[5] ), .Y(new_n3146_));
  XOR2X1   g02890(.A(new_n3146_), .B(new_n3142_), .Y(new_n3147_));
  AND2X1   g02891(.A(new_n3009_), .B(new_n2913_), .Y(new_n3148_));
  AOI21X1  g02892(.A0(new_n3010_), .A1(new_n2909_), .B0(new_n3148_), .Y(new_n3149_));
  XOR2X1   g02893(.A(new_n3149_), .B(new_n3147_), .Y(new_n3150_));
  AND2X1   g02894(.A(\b[36] ), .B(\b[35] ), .Y(new_n3151_));
  AOI21X1  g02895(.A0(new_n3014_), .A1(new_n3013_), .B0(new_n3151_), .Y(new_n3152_));
  XOR2X1   g02896(.A(\b[37] ), .B(\b[36] ), .Y(new_n3153_));
  INVX1    g02897(.A(new_n3153_), .Y(new_n3154_));
  XOR2X1   g02898(.A(new_n3154_), .B(new_n3152_), .Y(new_n3155_));
  INVX1    g02899(.A(\b[35] ), .Y(new_n3156_));
  AOI22X1  g02900(.A0(new_n267_), .A1(\b[37] ), .B0(new_n266_), .B1(\b[36] ), .Y(new_n3157_));
  OAI21X1  g02901(.A0(new_n350_), .A1(new_n3156_), .B0(new_n3157_), .Y(new_n3158_));
  AOI21X1  g02902(.A0(new_n3155_), .A1(new_n318_), .B0(new_n3158_), .Y(new_n3159_));
  XOR2X1   g02903(.A(new_n3159_), .B(\a[2] ), .Y(new_n3160_));
  XOR2X1   g02904(.A(new_n3160_), .B(new_n3150_), .Y(new_n3161_));
  XOR2X1   g02905(.A(new_n3161_), .B(new_n3028_), .Y(\f[37] ));
  OR2X1    g02906(.A(new_n3146_), .B(new_n3142_), .Y(new_n3163_));
  INVX1    g02907(.A(new_n3146_), .Y(new_n3164_));
  XOR2X1   g02908(.A(new_n3164_), .B(new_n3142_), .Y(new_n3165_));
  OAI21X1  g02909(.A0(new_n3149_), .A1(new_n3165_), .B0(new_n3163_), .Y(new_n3166_));
  AOI22X1  g02910(.A0(new_n369_), .A1(\b[35] ), .B0(new_n368_), .B1(\b[34] ), .Y(new_n3167_));
  OAI21X1  g02911(.A0(new_n367_), .A1(new_n2893_), .B0(new_n3167_), .Y(new_n3168_));
  AOI21X1  g02912(.A0(new_n2892_), .A1(new_n308_), .B0(new_n3168_), .Y(new_n3169_));
  XOR2X1   g02913(.A(new_n3169_), .B(new_n305_), .Y(new_n3170_));
  NOR2X1   g02914(.A(new_n3140_), .B(new_n3034_), .Y(new_n3171_));
  NAND2X1  g02915(.A(new_n3140_), .B(new_n3034_), .Y(new_n3172_));
  OAI21X1  g02916(.A0(new_n3171_), .A1(new_n3030_), .B0(new_n3172_), .Y(new_n3173_));
  AOI22X1  g02917(.A0(new_n469_), .A1(\b[32] ), .B0(new_n468_), .B1(\b[31] ), .Y(new_n3174_));
  OAI21X1  g02918(.A0(new_n467_), .A1(new_n2356_), .B0(new_n3174_), .Y(new_n3175_));
  AOI21X1  g02919(.A0(new_n2495_), .A1(new_n404_), .B0(new_n3175_), .Y(new_n3176_));
  XOR2X1   g02920(.A(new_n3176_), .B(new_n400_), .Y(new_n3177_));
  NOR2X1   g02921(.A(new_n3138_), .B(new_n3134_), .Y(new_n3178_));
  AOI21X1  g02922(.A0(new_n3139_), .A1(new_n3038_), .B0(new_n3178_), .Y(new_n3179_));
  AOI22X1  g02923(.A0(new_n603_), .A1(\b[29] ), .B0(new_n602_), .B1(\b[28] ), .Y(new_n3180_));
  OAI21X1  g02924(.A0(new_n601_), .A1(new_n2126_), .B0(new_n3180_), .Y(new_n3181_));
  AOI21X1  g02925(.A0(new_n2125_), .A1(new_n518_), .B0(new_n3181_), .Y(new_n3182_));
  XOR2X1   g02926(.A(new_n3182_), .B(\a[11] ), .Y(new_n3183_));
  NOR2X1   g02927(.A(new_n3119_), .B(new_n3115_), .Y(new_n3184_));
  AOI21X1  g02928(.A0(new_n3122_), .A1(new_n3120_), .B0(new_n3184_), .Y(new_n3185_));
  AND2X1   g02929(.A(new_n3094_), .B(new_n3053_), .Y(new_n3186_));
  AOI21X1  g02930(.A0(new_n3095_), .A1(new_n3048_), .B0(new_n3186_), .Y(new_n3187_));
  AND2X1   g02931(.A(new_n3091_), .B(new_n3060_), .Y(new_n3188_));
  INVX1    g02932(.A(new_n3188_), .Y(new_n3189_));
  OAI21X1  g02933(.A0(new_n3093_), .A1(new_n3055_), .B0(new_n3189_), .Y(new_n3190_));
  AOI22X1  g02934(.A0(new_n2163_), .A1(\b[11] ), .B0(new_n2162_), .B1(\b[10] ), .Y(new_n3191_));
  OAI21X1  g02935(.A0(new_n2161_), .A1(new_n590_), .B0(new_n3191_), .Y(new_n3192_));
  AOI21X1  g02936(.A0(new_n1907_), .A1(new_n589_), .B0(new_n3192_), .Y(new_n3193_));
  XOR2X1   g02937(.A(new_n3193_), .B(\a[29] ), .Y(new_n3194_));
  AND2X1   g02938(.A(new_n3089_), .B(new_n3068_), .Y(new_n3195_));
  AOI21X1  g02939(.A0(new_n3090_), .A1(new_n3064_), .B0(new_n3195_), .Y(new_n3196_));
  AND2X1   g02940(.A(new_n3087_), .B(new_n3075_), .Y(new_n3197_));
  AND2X1   g02941(.A(new_n3088_), .B(new_n3070_), .Y(new_n3198_));
  OR2X1    g02942(.A(new_n3198_), .B(new_n3197_), .Y(new_n3199_));
  NAND3X1  g02943(.A(new_n3085_), .B(new_n2942_), .C(\a[38] ), .Y(new_n3200_));
  NAND2X1  g02944(.A(new_n3080_), .B(new_n341_), .Y(new_n3201_));
  OR4X1    g02945(.A(new_n3081_), .B(new_n3079_), .C(new_n2941_), .D(new_n274_), .Y(new_n3202_));
  AND2X1   g02946(.A(new_n3081_), .B(new_n3077_), .Y(new_n3203_));
  AND2X1   g02947(.A(new_n3079_), .B(new_n2941_), .Y(new_n3204_));
  AOI22X1  g02948(.A0(new_n3204_), .A1(\b[2] ), .B0(new_n3203_), .B1(\b[1] ), .Y(new_n3205_));
  NAND3X1  g02949(.A(new_n3205_), .B(new_n3202_), .C(new_n3201_), .Y(new_n3206_));
  XOR2X1   g02950(.A(new_n3206_), .B(new_n3078_), .Y(new_n3207_));
  XOR2X1   g02951(.A(new_n3207_), .B(new_n3200_), .Y(new_n3208_));
  AOI22X1  g02952(.A0(new_n2813_), .A1(\b[5] ), .B0(new_n2812_), .B1(\b[4] ), .Y(new_n3209_));
  OAI21X1  g02953(.A0(new_n2946_), .A1(new_n297_), .B0(new_n3209_), .Y(new_n3210_));
  AOI21X1  g02954(.A0(new_n2652_), .A1(new_n349_), .B0(new_n3210_), .Y(new_n3211_));
  XOR2X1   g02955(.A(new_n3211_), .B(\a[35] ), .Y(new_n3212_));
  XOR2X1   g02956(.A(new_n3212_), .B(new_n3208_), .Y(new_n3213_));
  XOR2X1   g02957(.A(new_n3213_), .B(new_n3199_), .Y(new_n3214_));
  AOI22X1  g02958(.A0(new_n2545_), .A1(\b[8] ), .B0(new_n2544_), .B1(\b[7] ), .Y(new_n3215_));
  OAI21X1  g02959(.A0(new_n2543_), .A1(new_n392_), .B0(new_n3215_), .Y(new_n3216_));
  AOI21X1  g02960(.A0(new_n2260_), .A1(new_n454_), .B0(new_n3216_), .Y(new_n3217_));
  XOR2X1   g02961(.A(new_n3217_), .B(\a[32] ), .Y(new_n3218_));
  XOR2X1   g02962(.A(new_n3218_), .B(new_n3214_), .Y(new_n3219_));
  INVX1    g02963(.A(new_n3219_), .Y(new_n3220_));
  XOR2X1   g02964(.A(new_n3220_), .B(new_n3196_), .Y(new_n3221_));
  XOR2X1   g02965(.A(new_n3221_), .B(new_n3194_), .Y(new_n3222_));
  XOR2X1   g02966(.A(new_n3222_), .B(new_n3190_), .Y(new_n3223_));
  AOI22X1  g02967(.A0(new_n1814_), .A1(\b[14] ), .B0(new_n1813_), .B1(\b[13] ), .Y(new_n3224_));
  OAI21X1  g02968(.A0(new_n1812_), .A1(new_n713_), .B0(new_n3224_), .Y(new_n3225_));
  AOI21X1  g02969(.A0(new_n1617_), .A1(new_n734_), .B0(new_n3225_), .Y(new_n3226_));
  XOR2X1   g02970(.A(new_n3226_), .B(\a[26] ), .Y(new_n3227_));
  XOR2X1   g02971(.A(new_n3227_), .B(new_n3223_), .Y(new_n3228_));
  INVX1    g02972(.A(new_n3228_), .Y(new_n3229_));
  XOR2X1   g02973(.A(new_n3229_), .B(new_n3187_), .Y(new_n3230_));
  AOI22X1  g02974(.A0(new_n1526_), .A1(\b[17] ), .B0(new_n1525_), .B1(\b[16] ), .Y(new_n3231_));
  OAI21X1  g02975(.A0(new_n1524_), .A1(new_n977_), .B0(new_n3231_), .Y(new_n3232_));
  AOI21X1  g02976(.A0(new_n1347_), .A1(new_n976_), .B0(new_n3232_), .Y(new_n3233_));
  XOR2X1   g02977(.A(new_n3233_), .B(\a[23] ), .Y(new_n3234_));
  XOR2X1   g02978(.A(new_n3234_), .B(new_n3230_), .Y(new_n3235_));
  INVX1    g02979(.A(new_n3235_), .Y(new_n3236_));
  OR2X1    g02980(.A(new_n3101_), .B(new_n3097_), .Y(new_n3237_));
  OAI21X1  g02981(.A0(new_n3105_), .A1(new_n3104_), .B0(new_n3102_), .Y(new_n3238_));
  AND2X1   g02982(.A(new_n3238_), .B(new_n3237_), .Y(new_n3239_));
  XOR2X1   g02983(.A(new_n3239_), .B(new_n3236_), .Y(new_n3240_));
  AOI22X1  g02984(.A0(new_n1263_), .A1(\b[20] ), .B0(new_n1262_), .B1(\b[19] ), .Y(new_n3241_));
  OAI21X1  g02985(.A0(new_n1261_), .A1(new_n1115_), .B0(new_n3241_), .Y(new_n3242_));
  AOI21X1  g02986(.A0(new_n1217_), .A1(new_n1075_), .B0(new_n3242_), .Y(new_n3243_));
  XOR2X1   g02987(.A(new_n3243_), .B(\a[20] ), .Y(new_n3244_));
  XOR2X1   g02988(.A(new_n3244_), .B(new_n3240_), .Y(new_n3245_));
  XOR2X1   g02989(.A(new_n3110_), .B(\a[20] ), .Y(new_n3246_));
  NOR2X1   g02990(.A(new_n3246_), .B(new_n3107_), .Y(new_n3247_));
  XOR2X1   g02991(.A(new_n3246_), .B(new_n3107_), .Y(new_n3248_));
  AOI21X1  g02992(.A0(new_n3114_), .A1(new_n3248_), .B0(new_n3247_), .Y(new_n3249_));
  XOR2X1   g02993(.A(new_n3249_), .B(new_n3245_), .Y(new_n3250_));
  AOI22X1  g02994(.A0(new_n1017_), .A1(\b[23] ), .B0(new_n1016_), .B1(\b[22] ), .Y(new_n3251_));
  OAI21X1  g02995(.A0(new_n1015_), .A1(new_n1482_), .B0(new_n3251_), .Y(new_n3252_));
  AOI21X1  g02996(.A0(new_n1481_), .A1(new_n882_), .B0(new_n3252_), .Y(new_n3253_));
  XOR2X1   g02997(.A(new_n3253_), .B(\a[17] ), .Y(new_n3254_));
  AND2X1   g02998(.A(new_n3254_), .B(new_n3250_), .Y(new_n3255_));
  XOR2X1   g02999(.A(new_n3254_), .B(new_n3250_), .Y(new_n3256_));
  OR2X1    g03000(.A(new_n3254_), .B(new_n3250_), .Y(new_n3257_));
  OAI21X1  g03001(.A0(new_n3255_), .A1(new_n3185_), .B0(new_n3257_), .Y(new_n3258_));
  OAI22X1  g03002(.A0(new_n3258_), .A1(new_n3255_), .B0(new_n3256_), .B1(new_n3185_), .Y(new_n3259_));
  AOI22X1  g03003(.A0(new_n818_), .A1(\b[26] ), .B0(new_n817_), .B1(\b[25] ), .Y(new_n3260_));
  OAI21X1  g03004(.A0(new_n816_), .A1(new_n1588_), .B0(new_n3260_), .Y(new_n3261_));
  AOI21X1  g03005(.A0(new_n1783_), .A1(new_n668_), .B0(new_n3261_), .Y(new_n3262_));
  XOR2X1   g03006(.A(new_n3262_), .B(\a[14] ), .Y(new_n3263_));
  XOR2X1   g03007(.A(new_n3263_), .B(new_n3259_), .Y(new_n3264_));
  XOR2X1   g03008(.A(new_n3264_), .B(new_n3133_), .Y(new_n3265_));
  XOR2X1   g03009(.A(new_n3265_), .B(new_n3183_), .Y(new_n3266_));
  XOR2X1   g03010(.A(new_n3266_), .B(new_n3179_), .Y(new_n3267_));
  XOR2X1   g03011(.A(new_n3267_), .B(new_n3177_), .Y(new_n3268_));
  XOR2X1   g03012(.A(new_n3268_), .B(new_n3173_), .Y(new_n3269_));
  XOR2X1   g03013(.A(new_n3269_), .B(new_n3170_), .Y(new_n3270_));
  XOR2X1   g03014(.A(new_n3270_), .B(new_n3166_), .Y(new_n3271_));
  NAND2X1  g03015(.A(\b[37] ), .B(\b[36] ), .Y(new_n3272_));
  OAI21X1  g03016(.A0(new_n3154_), .A1(new_n3152_), .B0(new_n3272_), .Y(new_n3273_));
  XOR2X1   g03017(.A(\b[38] ), .B(\b[37] ), .Y(new_n3274_));
  XOR2X1   g03018(.A(new_n3274_), .B(new_n3273_), .Y(new_n3275_));
  INVX1    g03019(.A(\b[36] ), .Y(new_n3276_));
  AOI22X1  g03020(.A0(new_n267_), .A1(\b[38] ), .B0(new_n266_), .B1(\b[37] ), .Y(new_n3277_));
  OAI21X1  g03021(.A0(new_n350_), .A1(new_n3276_), .B0(new_n3277_), .Y(new_n3278_));
  AOI21X1  g03022(.A0(new_n3275_), .A1(new_n318_), .B0(new_n3278_), .Y(new_n3279_));
  XOR2X1   g03023(.A(new_n3279_), .B(\a[2] ), .Y(new_n3280_));
  XOR2X1   g03024(.A(new_n3280_), .B(new_n3271_), .Y(new_n3281_));
  OR2X1    g03025(.A(new_n3160_), .B(new_n3150_), .Y(new_n3282_));
  OAI21X1  g03026(.A0(new_n3027_), .A1(new_n3026_), .B0(new_n3161_), .Y(new_n3283_));
  AND2X1   g03027(.A(new_n3283_), .B(new_n3282_), .Y(new_n3284_));
  XOR2X1   g03028(.A(new_n3284_), .B(new_n3281_), .Y(\f[38] ));
  AND2X1   g03029(.A(new_n3269_), .B(new_n3170_), .Y(new_n3286_));
  AOI21X1  g03030(.A0(new_n3270_), .A1(new_n3166_), .B0(new_n3286_), .Y(new_n3287_));
  NOR2X1   g03031(.A(new_n2872_), .B(new_n2868_), .Y(new_n3288_));
  OR2X1    g03032(.A(new_n2738_), .B(new_n2734_), .Y(new_n3289_));
  INVX1    g03033(.A(new_n2738_), .Y(new_n3290_));
  XOR2X1   g03034(.A(new_n3290_), .B(new_n2734_), .Y(new_n3291_));
  OAI21X1  g03035(.A0(new_n2745_), .A1(new_n3291_), .B0(new_n3289_), .Y(new_n3292_));
  AOI21X1  g03036(.A0(new_n3292_), .A1(new_n2873_), .B0(new_n3288_), .Y(new_n3293_));
  AND2X1   g03037(.A(new_n3007_), .B(new_n3003_), .Y(new_n3294_));
  OR2X1    g03038(.A(new_n3007_), .B(new_n3003_), .Y(new_n3295_));
  OAI21X1  g03039(.A0(new_n3294_), .A1(new_n3293_), .B0(new_n3295_), .Y(new_n3296_));
  AND2X1   g03040(.A(new_n3140_), .B(new_n3034_), .Y(new_n3297_));
  AOI21X1  g03041(.A0(new_n3141_), .A1(new_n3296_), .B0(new_n3297_), .Y(new_n3298_));
  NOR2X1   g03042(.A(new_n3267_), .B(new_n3177_), .Y(new_n3299_));
  NAND2X1  g03043(.A(new_n3267_), .B(new_n3177_), .Y(new_n3300_));
  OAI21X1  g03044(.A0(new_n3299_), .A1(new_n3298_), .B0(new_n3300_), .Y(new_n3301_));
  INVX1    g03045(.A(new_n3183_), .Y(new_n3302_));
  NAND2X1  g03046(.A(new_n3265_), .B(new_n3302_), .Y(new_n3303_));
  OAI21X1  g03047(.A0(new_n3266_), .A1(new_n3179_), .B0(new_n3303_), .Y(new_n3304_));
  XOR2X1   g03048(.A(new_n3262_), .B(new_n665_), .Y(new_n3305_));
  AND2X1   g03049(.A(new_n3305_), .B(new_n3259_), .Y(new_n3306_));
  NOR2X1   g03050(.A(new_n3264_), .B(new_n3133_), .Y(new_n3307_));
  NOR2X1   g03051(.A(new_n3307_), .B(new_n3306_), .Y(new_n3308_));
  INVX1    g03052(.A(new_n3230_), .Y(new_n3309_));
  NOR2X1   g03053(.A(new_n3234_), .B(new_n3309_), .Y(new_n3310_));
  AOI21X1  g03054(.A0(new_n3238_), .A1(new_n3237_), .B0(new_n3235_), .Y(new_n3311_));
  NOR2X1   g03055(.A(new_n3311_), .B(new_n3310_), .Y(new_n3312_));
  OR2X1    g03056(.A(new_n3227_), .B(new_n3223_), .Y(new_n3313_));
  OAI21X1  g03057(.A0(new_n3229_), .A1(new_n3187_), .B0(new_n3313_), .Y(new_n3314_));
  OR2X1    g03058(.A(new_n3207_), .B(new_n3200_), .Y(new_n3315_));
  XOR2X1   g03059(.A(\a[39] ), .B(\a[38] ), .Y(new_n3316_));
  NAND2X1  g03060(.A(new_n3316_), .B(\b[0] ), .Y(new_n3317_));
  INVX1    g03061(.A(new_n3317_), .Y(new_n3318_));
  XOR2X1   g03062(.A(new_n3318_), .B(new_n3315_), .Y(new_n3319_));
  OR2X1    g03063(.A(new_n3081_), .B(new_n2941_), .Y(new_n3320_));
  OR2X1    g03064(.A(new_n3320_), .B(new_n3079_), .Y(new_n3321_));
  AOI22X1  g03065(.A0(new_n3204_), .A1(\b[3] ), .B0(new_n3203_), .B1(\b[2] ), .Y(new_n3322_));
  OAI21X1  g03066(.A0(new_n3321_), .A1(new_n275_), .B0(new_n3322_), .Y(new_n3323_));
  AOI21X1  g03067(.A0(new_n3080_), .A1(new_n366_), .B0(new_n3323_), .Y(new_n3324_));
  XOR2X1   g03068(.A(new_n3324_), .B(\a[38] ), .Y(new_n3325_));
  XOR2X1   g03069(.A(new_n3325_), .B(new_n3319_), .Y(new_n3326_));
  AOI22X1  g03070(.A0(new_n2813_), .A1(\b[6] ), .B0(new_n2812_), .B1(\b[5] ), .Y(new_n3327_));
  OAI21X1  g03071(.A0(new_n2946_), .A1(new_n325_), .B0(new_n3327_), .Y(new_n3328_));
  AOI21X1  g03072(.A0(new_n2652_), .A1(new_n378_), .B0(new_n3328_), .Y(new_n3329_));
  XOR2X1   g03073(.A(new_n3329_), .B(\a[35] ), .Y(new_n3330_));
  XOR2X1   g03074(.A(new_n3330_), .B(new_n3326_), .Y(new_n3331_));
  XOR2X1   g03075(.A(new_n3211_), .B(new_n2650_), .Y(new_n3332_));
  AND2X1   g03076(.A(new_n3332_), .B(new_n3208_), .Y(new_n3333_));
  INVX1    g03077(.A(new_n3213_), .Y(new_n3334_));
  AOI21X1  g03078(.A0(new_n3334_), .A1(new_n3199_), .B0(new_n3333_), .Y(new_n3335_));
  XOR2X1   g03079(.A(new_n3335_), .B(new_n3331_), .Y(new_n3336_));
  AOI22X1  g03080(.A0(new_n2545_), .A1(\b[9] ), .B0(new_n2544_), .B1(\b[8] ), .Y(new_n3337_));
  OAI21X1  g03081(.A0(new_n2543_), .A1(new_n492_), .B0(new_n3337_), .Y(new_n3338_));
  AOI21X1  g03082(.A0(new_n2260_), .A1(new_n491_), .B0(new_n3338_), .Y(new_n3339_));
  XOR2X1   g03083(.A(new_n3339_), .B(\a[32] ), .Y(new_n3340_));
  XOR2X1   g03084(.A(new_n3340_), .B(new_n3336_), .Y(new_n3341_));
  INVX1    g03085(.A(new_n3341_), .Y(new_n3342_));
  OR2X1    g03086(.A(new_n3220_), .B(new_n3196_), .Y(new_n3343_));
  OAI21X1  g03087(.A0(new_n3218_), .A1(new_n3214_), .B0(new_n3343_), .Y(new_n3344_));
  XOR2X1   g03088(.A(new_n3344_), .B(new_n3342_), .Y(new_n3345_));
  AOI22X1  g03089(.A0(new_n2163_), .A1(\b[12] ), .B0(new_n2162_), .B1(\b[11] ), .Y(new_n3346_));
  OAI21X1  g03090(.A0(new_n2161_), .A1(new_n587_), .B0(new_n3346_), .Y(new_n3347_));
  AOI21X1  g03091(.A0(new_n1907_), .A1(new_n635_), .B0(new_n3347_), .Y(new_n3348_));
  XOR2X1   g03092(.A(new_n3348_), .B(\a[29] ), .Y(new_n3349_));
  XOR2X1   g03093(.A(new_n3349_), .B(new_n3345_), .Y(new_n3350_));
  INVX1    g03094(.A(new_n3194_), .Y(new_n3351_));
  AND2X1   g03095(.A(new_n3221_), .B(new_n3351_), .Y(new_n3352_));
  INVX1    g03096(.A(new_n3222_), .Y(new_n3353_));
  AOI21X1  g03097(.A0(new_n3353_), .A1(new_n3190_), .B0(new_n3352_), .Y(new_n3354_));
  XOR2X1   g03098(.A(new_n3354_), .B(new_n3350_), .Y(new_n3355_));
  AOI22X1  g03099(.A0(new_n1814_), .A1(\b[15] ), .B0(new_n1813_), .B1(\b[14] ), .Y(new_n3356_));
  OAI21X1  g03100(.A0(new_n1812_), .A1(new_n795_), .B0(new_n3356_), .Y(new_n3357_));
  AOI21X1  g03101(.A0(new_n1617_), .A1(new_n794_), .B0(new_n3357_), .Y(new_n3358_));
  XOR2X1   g03102(.A(new_n3358_), .B(\a[26] ), .Y(new_n3359_));
  XOR2X1   g03103(.A(new_n3359_), .B(new_n3355_), .Y(new_n3360_));
  XOR2X1   g03104(.A(new_n3360_), .B(new_n3314_), .Y(new_n3361_));
  AOI22X1  g03105(.A0(new_n1526_), .A1(\b[18] ), .B0(new_n1525_), .B1(\b[17] ), .Y(new_n3362_));
  OAI21X1  g03106(.A0(new_n1524_), .A1(new_n974_), .B0(new_n3362_), .Y(new_n3363_));
  AOI21X1  g03107(.A0(new_n1347_), .A1(new_n1042_), .B0(new_n3363_), .Y(new_n3364_));
  XOR2X1   g03108(.A(new_n3364_), .B(\a[23] ), .Y(new_n3365_));
  XOR2X1   g03109(.A(new_n3365_), .B(new_n3361_), .Y(new_n3366_));
  XOR2X1   g03110(.A(new_n3366_), .B(new_n3312_), .Y(new_n3367_));
  AOI22X1  g03111(.A0(new_n1263_), .A1(\b[21] ), .B0(new_n1262_), .B1(\b[20] ), .Y(new_n3368_));
  OAI21X1  g03112(.A0(new_n1261_), .A1(new_n1300_), .B0(new_n3368_), .Y(new_n3369_));
  AOI21X1  g03113(.A0(new_n1299_), .A1(new_n1075_), .B0(new_n3369_), .Y(new_n3370_));
  XOR2X1   g03114(.A(new_n3370_), .B(\a[20] ), .Y(new_n3371_));
  XOR2X1   g03115(.A(new_n3371_), .B(new_n3367_), .Y(new_n3372_));
  OR2X1    g03116(.A(new_n3244_), .B(new_n3240_), .Y(new_n3373_));
  XOR2X1   g03117(.A(new_n3239_), .B(new_n3235_), .Y(new_n3374_));
  XOR2X1   g03118(.A(new_n3244_), .B(new_n3374_), .Y(new_n3375_));
  OAI21X1  g03119(.A0(new_n3249_), .A1(new_n3375_), .B0(new_n3373_), .Y(new_n3376_));
  XOR2X1   g03120(.A(new_n3376_), .B(new_n3372_), .Y(new_n3377_));
  AOI22X1  g03121(.A0(new_n1017_), .A1(\b[24] ), .B0(new_n1016_), .B1(\b[23] ), .Y(new_n3378_));
  OAI21X1  g03122(.A0(new_n1015_), .A1(new_n1479_), .B0(new_n3378_), .Y(new_n3379_));
  AOI21X1  g03123(.A0(new_n1572_), .A1(new_n882_), .B0(new_n3379_), .Y(new_n3380_));
  XOR2X1   g03124(.A(new_n3380_), .B(\a[17] ), .Y(new_n3381_));
  XOR2X1   g03125(.A(new_n3381_), .B(new_n3377_), .Y(new_n3382_));
  XOR2X1   g03126(.A(new_n3382_), .B(new_n3258_), .Y(new_n3383_));
  AOI22X1  g03127(.A0(new_n818_), .A1(\b[27] ), .B0(new_n817_), .B1(\b[26] ), .Y(new_n3384_));
  OAI21X1  g03128(.A0(new_n816_), .A1(new_n1880_), .B0(new_n3384_), .Y(new_n3385_));
  AOI21X1  g03129(.A0(new_n1879_), .A1(new_n668_), .B0(new_n3385_), .Y(new_n3386_));
  XOR2X1   g03130(.A(new_n3386_), .B(\a[14] ), .Y(new_n3387_));
  XOR2X1   g03131(.A(new_n3387_), .B(new_n3383_), .Y(new_n3388_));
  XOR2X1   g03132(.A(new_n3388_), .B(new_n3308_), .Y(new_n3389_));
  AOI22X1  g03133(.A0(new_n603_), .A1(\b[30] ), .B0(new_n602_), .B1(\b[29] ), .Y(new_n3390_));
  OAI21X1  g03134(.A0(new_n601_), .A1(new_n2231_), .B0(new_n3390_), .Y(new_n3391_));
  AOI21X1  g03135(.A0(new_n2230_), .A1(new_n518_), .B0(new_n3391_), .Y(new_n3392_));
  XOR2X1   g03136(.A(new_n3392_), .B(\a[11] ), .Y(new_n3393_));
  XOR2X1   g03137(.A(new_n3393_), .B(new_n3389_), .Y(new_n3394_));
  XOR2X1   g03138(.A(new_n3394_), .B(new_n3304_), .Y(new_n3395_));
  AOI22X1  g03139(.A0(new_n469_), .A1(\b[33] ), .B0(new_n468_), .B1(\b[32] ), .Y(new_n3396_));
  OAI21X1  g03140(.A0(new_n467_), .A1(new_n2615_), .B0(new_n3396_), .Y(new_n3397_));
  AOI21X1  g03141(.A0(new_n2614_), .A1(new_n404_), .B0(new_n3397_), .Y(new_n3398_));
  XOR2X1   g03142(.A(new_n3398_), .B(\a[8] ), .Y(new_n3399_));
  XOR2X1   g03143(.A(new_n3399_), .B(new_n3395_), .Y(new_n3400_));
  XOR2X1   g03144(.A(new_n3400_), .B(new_n3301_), .Y(new_n3401_));
  AOI22X1  g03145(.A0(new_n369_), .A1(\b[36] ), .B0(new_n368_), .B1(\b[35] ), .Y(new_n3402_));
  OAI21X1  g03146(.A0(new_n367_), .A1(new_n2890_), .B0(new_n3402_), .Y(new_n3403_));
  AOI21X1  g03147(.A0(new_n3015_), .A1(new_n308_), .B0(new_n3403_), .Y(new_n3404_));
  XOR2X1   g03148(.A(new_n3404_), .B(\a[5] ), .Y(new_n3405_));
  XOR2X1   g03149(.A(new_n3405_), .B(new_n3401_), .Y(new_n3406_));
  XOR2X1   g03150(.A(new_n3406_), .B(new_n3287_), .Y(new_n3407_));
  AND2X1   g03151(.A(\b[38] ), .B(\b[37] ), .Y(new_n3408_));
  AOI21X1  g03152(.A0(new_n3274_), .A1(new_n3273_), .B0(new_n3408_), .Y(new_n3409_));
  XOR2X1   g03153(.A(\b[39] ), .B(\b[38] ), .Y(new_n3410_));
  INVX1    g03154(.A(new_n3410_), .Y(new_n3411_));
  XOR2X1   g03155(.A(new_n3411_), .B(new_n3409_), .Y(new_n3412_));
  INVX1    g03156(.A(\b[37] ), .Y(new_n3413_));
  AOI22X1  g03157(.A0(new_n267_), .A1(\b[39] ), .B0(new_n266_), .B1(\b[38] ), .Y(new_n3414_));
  OAI21X1  g03158(.A0(new_n350_), .A1(new_n3413_), .B0(new_n3414_), .Y(new_n3415_));
  AOI21X1  g03159(.A0(new_n3412_), .A1(new_n318_), .B0(new_n3415_), .Y(new_n3416_));
  XOR2X1   g03160(.A(new_n3416_), .B(\a[2] ), .Y(new_n3417_));
  XOR2X1   g03161(.A(new_n3417_), .B(new_n3407_), .Y(new_n3418_));
  INVX1    g03162(.A(new_n3280_), .Y(new_n3419_));
  AND2X1   g03163(.A(new_n3419_), .B(new_n3271_), .Y(new_n3420_));
  AOI21X1  g03164(.A0(new_n3283_), .A1(new_n3282_), .B0(new_n3281_), .Y(new_n3421_));
  OR2X1    g03165(.A(new_n3421_), .B(new_n3420_), .Y(new_n3422_));
  XOR2X1   g03166(.A(new_n3422_), .B(new_n3418_), .Y(\f[39] ));
  OR2X1    g03167(.A(new_n3417_), .B(new_n3407_), .Y(new_n3424_));
  OAI21X1  g03168(.A0(new_n3421_), .A1(new_n3420_), .B0(new_n3418_), .Y(new_n3425_));
  AND2X1   g03169(.A(new_n3425_), .B(new_n3424_), .Y(new_n3426_));
  NOR2X1   g03170(.A(new_n3146_), .B(new_n3142_), .Y(new_n3427_));
  NAND2X1  g03171(.A(new_n3009_), .B(new_n2913_), .Y(new_n3428_));
  NOR2X1   g03172(.A(new_n3009_), .B(new_n2913_), .Y(new_n3429_));
  OAI21X1  g03173(.A0(new_n3429_), .A1(new_n3024_), .B0(new_n3428_), .Y(new_n3430_));
  AOI21X1  g03174(.A0(new_n3430_), .A1(new_n3147_), .B0(new_n3427_), .Y(new_n3431_));
  NOR2X1   g03175(.A(new_n3269_), .B(new_n3170_), .Y(new_n3432_));
  NAND2X1  g03176(.A(new_n3269_), .B(new_n3170_), .Y(new_n3433_));
  OAI21X1  g03177(.A0(new_n3432_), .A1(new_n3431_), .B0(new_n3433_), .Y(new_n3434_));
  NOR2X1   g03178(.A(new_n3405_), .B(new_n3401_), .Y(new_n3435_));
  AOI21X1  g03179(.A0(new_n3406_), .A1(new_n3434_), .B0(new_n3435_), .Y(new_n3436_));
  AND2X1   g03180(.A(new_n3267_), .B(new_n3177_), .Y(new_n3437_));
  AOI21X1  g03181(.A0(new_n3268_), .A1(new_n3173_), .B0(new_n3437_), .Y(new_n3438_));
  NOR2X1   g03182(.A(new_n3037_), .B(new_n3036_), .Y(new_n3439_));
  AND2X1   g03183(.A(new_n3138_), .B(new_n3134_), .Y(new_n3440_));
  OR2X1    g03184(.A(new_n3138_), .B(new_n3134_), .Y(new_n3441_));
  OAI21X1  g03185(.A0(new_n3440_), .A1(new_n3439_), .B0(new_n3441_), .Y(new_n3442_));
  AND2X1   g03186(.A(new_n3265_), .B(new_n3302_), .Y(new_n3443_));
  XOR2X1   g03187(.A(new_n3265_), .B(new_n3302_), .Y(new_n3444_));
  AOI21X1  g03188(.A0(new_n3444_), .A1(new_n3442_), .B0(new_n3443_), .Y(new_n3445_));
  XOR2X1   g03189(.A(new_n3394_), .B(new_n3445_), .Y(new_n3446_));
  OR2X1    g03190(.A(new_n3399_), .B(new_n3446_), .Y(new_n3447_));
  OAI21X1  g03191(.A0(new_n3400_), .A1(new_n3438_), .B0(new_n3447_), .Y(new_n3448_));
  AOI22X1  g03192(.A0(new_n469_), .A1(\b[34] ), .B0(new_n468_), .B1(\b[33] ), .Y(new_n3449_));
  OAI21X1  g03193(.A0(new_n467_), .A1(new_n2612_), .B0(new_n3449_), .Y(new_n3450_));
  AOI21X1  g03194(.A0(new_n2759_), .A1(new_n404_), .B0(new_n3450_), .Y(new_n3451_));
  XOR2X1   g03195(.A(new_n3451_), .B(new_n400_), .Y(new_n3452_));
  OR2X1    g03196(.A(new_n3393_), .B(new_n3389_), .Y(new_n3453_));
  AND2X1   g03197(.A(new_n3393_), .B(new_n3389_), .Y(new_n3454_));
  OAI21X1  g03198(.A0(new_n3454_), .A1(new_n3445_), .B0(new_n3453_), .Y(new_n3455_));
  OR2X1    g03199(.A(new_n3387_), .B(new_n3383_), .Y(new_n3456_));
  OAI21X1  g03200(.A0(new_n3307_), .A1(new_n3306_), .B0(new_n3388_), .Y(new_n3457_));
  NAND2X1  g03201(.A(new_n3457_), .B(new_n3456_), .Y(new_n3458_));
  AOI22X1  g03202(.A0(new_n818_), .A1(\b[28] ), .B0(new_n817_), .B1(\b[27] ), .Y(new_n3459_));
  OAI21X1  g03203(.A0(new_n816_), .A1(new_n1877_), .B0(new_n3459_), .Y(new_n3460_));
  AOI21X1  g03204(.A0(new_n2004_), .A1(new_n668_), .B0(new_n3460_), .Y(new_n3461_));
  XOR2X1   g03205(.A(new_n3461_), .B(\a[14] ), .Y(new_n3462_));
  XOR2X1   g03206(.A(new_n3348_), .B(new_n1911_), .Y(new_n3463_));
  NAND2X1  g03207(.A(new_n3463_), .B(new_n3345_), .Y(new_n3464_));
  OAI21X1  g03208(.A0(new_n3354_), .A1(new_n3350_), .B0(new_n3464_), .Y(new_n3465_));
  XOR2X1   g03209(.A(new_n3339_), .B(new_n2258_), .Y(new_n3466_));
  AND2X1   g03210(.A(new_n3466_), .B(new_n3336_), .Y(new_n3467_));
  AND2X1   g03211(.A(new_n3344_), .B(new_n3342_), .Y(new_n3468_));
  OR4X1    g03212(.A(new_n3317_), .B(new_n3207_), .C(new_n3086_), .D(new_n3076_), .Y(new_n3469_));
  OAI21X1  g03213(.A0(new_n3325_), .A1(new_n3319_), .B0(new_n3469_), .Y(new_n3470_));
  AND2X1   g03214(.A(new_n3080_), .B(new_n323_), .Y(new_n3471_));
  NOR3X1   g03215(.A(new_n3320_), .B(new_n3079_), .C(new_n277_), .Y(new_n3472_));
  OAI22X1  g03216(.A0(new_n3083_), .A1(new_n325_), .B0(new_n3082_), .B1(new_n297_), .Y(new_n3473_));
  NOR3X1   g03217(.A(new_n3473_), .B(new_n3472_), .C(new_n3471_), .Y(new_n3474_));
  XOR2X1   g03218(.A(new_n3474_), .B(new_n3078_), .Y(new_n3475_));
  NAND2X1  g03219(.A(new_n3317_), .B(\a[41] ), .Y(new_n3476_));
  XOR2X1   g03220(.A(\a[39] ), .B(new_n3078_), .Y(new_n3477_));
  INVX1    g03221(.A(\a[41] ), .Y(new_n3478_));
  XOR2X1   g03222(.A(new_n3478_), .B(\a[40] ), .Y(new_n3479_));
  NOR2X1   g03223(.A(new_n3479_), .B(new_n3477_), .Y(new_n3480_));
  XOR2X1   g03224(.A(\a[40] ), .B(\a[39] ), .Y(new_n3481_));
  NAND2X1  g03225(.A(new_n3481_), .B(new_n3477_), .Y(new_n3482_));
  NAND2X1  g03226(.A(new_n3479_), .B(new_n3316_), .Y(new_n3483_));
  OAI22X1  g03227(.A0(new_n3483_), .A1(new_n275_), .B0(new_n3482_), .B1(new_n274_), .Y(new_n3484_));
  AOI21X1  g03228(.A0(new_n3480_), .A1(new_n263_), .B0(new_n3484_), .Y(new_n3485_));
  XOR2X1   g03229(.A(new_n3485_), .B(\a[41] ), .Y(new_n3486_));
  XOR2X1   g03230(.A(new_n3486_), .B(new_n3476_), .Y(new_n3487_));
  XOR2X1   g03231(.A(new_n3487_), .B(new_n3475_), .Y(new_n3488_));
  XOR2X1   g03232(.A(new_n3488_), .B(new_n3470_), .Y(new_n3489_));
  AOI22X1  g03233(.A0(new_n2813_), .A1(\b[7] ), .B0(new_n2812_), .B1(\b[6] ), .Y(new_n3490_));
  OAI21X1  g03234(.A0(new_n2946_), .A1(new_n395_), .B0(new_n3490_), .Y(new_n3491_));
  AOI21X1  g03235(.A0(new_n2652_), .A1(new_n394_), .B0(new_n3491_), .Y(new_n3492_));
  XOR2X1   g03236(.A(new_n3492_), .B(\a[35] ), .Y(new_n3493_));
  XOR2X1   g03237(.A(new_n3493_), .B(new_n3489_), .Y(new_n3494_));
  INVX1    g03238(.A(new_n3494_), .Y(new_n3495_));
  INVX1    g03239(.A(new_n3330_), .Y(new_n3496_));
  NOR2X1   g03240(.A(new_n3335_), .B(new_n3331_), .Y(new_n3497_));
  AOI21X1  g03241(.A0(new_n3496_), .A1(new_n3326_), .B0(new_n3497_), .Y(new_n3498_));
  XOR2X1   g03242(.A(new_n3498_), .B(new_n3495_), .Y(new_n3499_));
  AOI22X1  g03243(.A0(new_n2545_), .A1(\b[10] ), .B0(new_n2544_), .B1(\b[9] ), .Y(new_n3500_));
  OAI21X1  g03244(.A0(new_n2543_), .A1(new_n489_), .B0(new_n3500_), .Y(new_n3501_));
  AOI21X1  g03245(.A0(new_n2260_), .A1(new_n543_), .B0(new_n3501_), .Y(new_n3502_));
  XOR2X1   g03246(.A(new_n3502_), .B(\a[32] ), .Y(new_n3503_));
  NOR2X1   g03247(.A(new_n3503_), .B(new_n3499_), .Y(new_n3504_));
  AND2X1   g03248(.A(new_n3503_), .B(new_n3499_), .Y(new_n3505_));
  OAI22X1  g03249(.A0(new_n3505_), .A1(new_n3504_), .B0(new_n3468_), .B1(new_n3467_), .Y(new_n3506_));
  OR4X1    g03250(.A(new_n3505_), .B(new_n3504_), .C(new_n3468_), .D(new_n3467_), .Y(new_n3507_));
  AND2X1   g03251(.A(new_n3507_), .B(new_n3506_), .Y(new_n3508_));
  AOI22X1  g03252(.A0(new_n2163_), .A1(\b[13] ), .B0(new_n2162_), .B1(\b[12] ), .Y(new_n3509_));
  OAI21X1  g03253(.A0(new_n2161_), .A1(new_n716_), .B0(new_n3509_), .Y(new_n3510_));
  AOI21X1  g03254(.A0(new_n1907_), .A1(new_n715_), .B0(new_n3510_), .Y(new_n3511_));
  XOR2X1   g03255(.A(new_n3511_), .B(\a[29] ), .Y(new_n3512_));
  XOR2X1   g03256(.A(new_n3512_), .B(new_n3508_), .Y(new_n3513_));
  XOR2X1   g03257(.A(new_n3513_), .B(new_n3465_), .Y(new_n3514_));
  AOI22X1  g03258(.A0(new_n1814_), .A1(\b[16] ), .B0(new_n1813_), .B1(\b[15] ), .Y(new_n3515_));
  OAI21X1  g03259(.A0(new_n1812_), .A1(new_n792_), .B0(new_n3515_), .Y(new_n3516_));
  AOI21X1  g03260(.A0(new_n1617_), .A1(new_n842_), .B0(new_n3516_), .Y(new_n3517_));
  XOR2X1   g03261(.A(new_n3517_), .B(\a[26] ), .Y(new_n3518_));
  XOR2X1   g03262(.A(new_n3518_), .B(new_n3514_), .Y(new_n3519_));
  INVX1    g03263(.A(new_n3355_), .Y(new_n3520_));
  NOR2X1   g03264(.A(new_n3359_), .B(new_n3520_), .Y(new_n3521_));
  INVX1    g03265(.A(new_n3360_), .Y(new_n3522_));
  AOI21X1  g03266(.A0(new_n3522_), .A1(new_n3314_), .B0(new_n3521_), .Y(new_n3523_));
  XOR2X1   g03267(.A(new_n3523_), .B(new_n3519_), .Y(new_n3524_));
  AOI22X1  g03268(.A0(new_n1526_), .A1(\b[19] ), .B0(new_n1525_), .B1(\b[18] ), .Y(new_n3525_));
  OAI21X1  g03269(.A0(new_n1524_), .A1(new_n1118_), .B0(new_n3525_), .Y(new_n3526_));
  AOI21X1  g03270(.A0(new_n1347_), .A1(new_n1117_), .B0(new_n3526_), .Y(new_n3527_));
  XOR2X1   g03271(.A(new_n3527_), .B(\a[23] ), .Y(new_n3528_));
  XOR2X1   g03272(.A(new_n3528_), .B(new_n3524_), .Y(new_n3529_));
  OR2X1    g03273(.A(new_n3365_), .B(new_n3361_), .Y(new_n3530_));
  OAI21X1  g03274(.A0(new_n3311_), .A1(new_n3310_), .B0(new_n3366_), .Y(new_n3531_));
  AND2X1   g03275(.A(new_n3531_), .B(new_n3530_), .Y(new_n3532_));
  XOR2X1   g03276(.A(new_n3532_), .B(new_n3529_), .Y(new_n3533_));
  AOI22X1  g03277(.A0(new_n1263_), .A1(\b[22] ), .B0(new_n1262_), .B1(\b[21] ), .Y(new_n3534_));
  OAI21X1  g03278(.A0(new_n1261_), .A1(new_n1297_), .B0(new_n3534_), .Y(new_n3535_));
  AOI21X1  g03279(.A0(new_n1399_), .A1(new_n1075_), .B0(new_n3535_), .Y(new_n3536_));
  XOR2X1   g03280(.A(new_n3536_), .B(\a[20] ), .Y(new_n3537_));
  XOR2X1   g03281(.A(new_n3537_), .B(new_n3533_), .Y(new_n3538_));
  NOR2X1   g03282(.A(new_n3371_), .B(new_n3367_), .Y(new_n3539_));
  AOI21X1  g03283(.A0(new_n3376_), .A1(new_n3372_), .B0(new_n3539_), .Y(new_n3540_));
  XOR2X1   g03284(.A(new_n3540_), .B(new_n3538_), .Y(new_n3541_));
  AOI22X1  g03285(.A0(new_n1017_), .A1(\b[25] ), .B0(new_n1016_), .B1(\b[24] ), .Y(new_n3542_));
  OAI21X1  g03286(.A0(new_n1015_), .A1(new_n1591_), .B0(new_n3542_), .Y(new_n3543_));
  AOI21X1  g03287(.A0(new_n1590_), .A1(new_n882_), .B0(new_n3543_), .Y(new_n3544_));
  XOR2X1   g03288(.A(new_n3544_), .B(\a[17] ), .Y(new_n3545_));
  XOR2X1   g03289(.A(new_n3545_), .B(new_n3541_), .Y(new_n3546_));
  XOR2X1   g03290(.A(new_n3370_), .B(new_n1072_), .Y(new_n3547_));
  XOR2X1   g03291(.A(new_n3547_), .B(new_n3367_), .Y(new_n3548_));
  XOR2X1   g03292(.A(new_n3376_), .B(new_n3548_), .Y(new_n3549_));
  OR2X1    g03293(.A(new_n3381_), .B(new_n3549_), .Y(new_n3550_));
  XOR2X1   g03294(.A(new_n3381_), .B(new_n3549_), .Y(new_n3551_));
  NAND2X1  g03295(.A(new_n3551_), .B(new_n3258_), .Y(new_n3552_));
  AND2X1   g03296(.A(new_n3552_), .B(new_n3550_), .Y(new_n3553_));
  XOR2X1   g03297(.A(new_n3553_), .B(new_n3546_), .Y(new_n3554_));
  XOR2X1   g03298(.A(new_n3554_), .B(new_n3462_), .Y(new_n3555_));
  XOR2X1   g03299(.A(new_n3555_), .B(new_n3458_), .Y(new_n3556_));
  AOI22X1  g03300(.A0(new_n603_), .A1(\b[31] ), .B0(new_n602_), .B1(\b[30] ), .Y(new_n3557_));
  OAI21X1  g03301(.A0(new_n601_), .A1(new_n2359_), .B0(new_n3557_), .Y(new_n3558_));
  AOI21X1  g03302(.A0(new_n2358_), .A1(new_n518_), .B0(new_n3558_), .Y(new_n3559_));
  XOR2X1   g03303(.A(new_n3559_), .B(\a[11] ), .Y(new_n3560_));
  XOR2X1   g03304(.A(new_n3560_), .B(new_n3556_), .Y(new_n3561_));
  XOR2X1   g03305(.A(new_n3561_), .B(new_n3455_), .Y(new_n3562_));
  XOR2X1   g03306(.A(new_n3562_), .B(new_n3452_), .Y(new_n3563_));
  XOR2X1   g03307(.A(new_n3563_), .B(new_n3448_), .Y(new_n3564_));
  AOI22X1  g03308(.A0(new_n369_), .A1(\b[37] ), .B0(new_n368_), .B1(\b[36] ), .Y(new_n3565_));
  OAI21X1  g03309(.A0(new_n367_), .A1(new_n3156_), .B0(new_n3565_), .Y(new_n3566_));
  AOI21X1  g03310(.A0(new_n3155_), .A1(new_n308_), .B0(new_n3566_), .Y(new_n3567_));
  XOR2X1   g03311(.A(new_n3567_), .B(\a[5] ), .Y(new_n3568_));
  XOR2X1   g03312(.A(new_n3568_), .B(new_n3564_), .Y(new_n3569_));
  XOR2X1   g03313(.A(new_n3569_), .B(new_n3436_), .Y(new_n3570_));
  NAND2X1  g03314(.A(\b[39] ), .B(\b[38] ), .Y(new_n3571_));
  OAI21X1  g03315(.A0(new_n3411_), .A1(new_n3409_), .B0(new_n3571_), .Y(new_n3572_));
  XOR2X1   g03316(.A(\b[40] ), .B(\b[39] ), .Y(new_n3573_));
  XOR2X1   g03317(.A(new_n3573_), .B(new_n3572_), .Y(new_n3574_));
  INVX1    g03318(.A(\b[38] ), .Y(new_n3575_));
  AOI22X1  g03319(.A0(new_n267_), .A1(\b[40] ), .B0(new_n266_), .B1(\b[39] ), .Y(new_n3576_));
  OAI21X1  g03320(.A0(new_n350_), .A1(new_n3575_), .B0(new_n3576_), .Y(new_n3577_));
  AOI21X1  g03321(.A0(new_n3574_), .A1(new_n318_), .B0(new_n3577_), .Y(new_n3578_));
  XOR2X1   g03322(.A(new_n3578_), .B(\a[2] ), .Y(new_n3579_));
  XOR2X1   g03323(.A(new_n3579_), .B(new_n3570_), .Y(new_n3580_));
  XOR2X1   g03324(.A(new_n3580_), .B(new_n3426_), .Y(\f[40] ));
  AND2X1   g03325(.A(new_n3405_), .B(new_n3401_), .Y(new_n3582_));
  OR2X1    g03326(.A(new_n3405_), .B(new_n3401_), .Y(new_n3583_));
  OAI21X1  g03327(.A0(new_n3582_), .A1(new_n3287_), .B0(new_n3583_), .Y(new_n3584_));
  XOR2X1   g03328(.A(new_n3569_), .B(new_n3584_), .Y(new_n3585_));
  NOR2X1   g03329(.A(new_n3579_), .B(new_n3585_), .Y(new_n3586_));
  AOI21X1  g03330(.A0(new_n3425_), .A1(new_n3424_), .B0(new_n3580_), .Y(new_n3587_));
  OR2X1    g03331(.A(new_n3587_), .B(new_n3586_), .Y(new_n3588_));
  NOR2X1   g03332(.A(new_n3399_), .B(new_n3446_), .Y(new_n3589_));
  XOR2X1   g03333(.A(new_n3399_), .B(new_n3446_), .Y(new_n3590_));
  AOI21X1  g03334(.A0(new_n3590_), .A1(new_n3301_), .B0(new_n3589_), .Y(new_n3591_));
  XOR2X1   g03335(.A(new_n3563_), .B(new_n3591_), .Y(new_n3592_));
  NOR2X1   g03336(.A(new_n3568_), .B(new_n3592_), .Y(new_n3593_));
  XOR2X1   g03337(.A(new_n3568_), .B(new_n3592_), .Y(new_n3594_));
  AOI21X1  g03338(.A0(new_n3594_), .A1(new_n3584_), .B0(new_n3593_), .Y(new_n3595_));
  AND2X1   g03339(.A(new_n3562_), .B(new_n3452_), .Y(new_n3596_));
  AOI21X1  g03340(.A0(new_n3563_), .A1(new_n3448_), .B0(new_n3596_), .Y(new_n3597_));
  NOR2X1   g03341(.A(new_n3560_), .B(new_n3556_), .Y(new_n3598_));
  AOI21X1  g03342(.A0(new_n3561_), .A1(new_n3455_), .B0(new_n3598_), .Y(new_n3599_));
  AOI22X1  g03343(.A0(new_n603_), .A1(\b[32] ), .B0(new_n602_), .B1(\b[31] ), .Y(new_n3600_));
  OAI21X1  g03344(.A0(new_n601_), .A1(new_n2356_), .B0(new_n3600_), .Y(new_n3601_));
  AOI21X1  g03345(.A0(new_n2495_), .A1(new_n518_), .B0(new_n3601_), .Y(new_n3602_));
  XOR2X1   g03346(.A(new_n3602_), .B(new_n515_), .Y(new_n3603_));
  INVX1    g03347(.A(new_n3462_), .Y(new_n3604_));
  AND2X1   g03348(.A(new_n3554_), .B(new_n3604_), .Y(new_n3605_));
  AOI21X1  g03349(.A0(new_n3457_), .A1(new_n3456_), .B0(new_n3555_), .Y(new_n3606_));
  OR2X1    g03350(.A(new_n3606_), .B(new_n3605_), .Y(new_n3607_));
  AOI22X1  g03351(.A0(new_n818_), .A1(\b[29] ), .B0(new_n817_), .B1(\b[28] ), .Y(new_n3608_));
  OAI21X1  g03352(.A0(new_n816_), .A1(new_n2126_), .B0(new_n3608_), .Y(new_n3609_));
  AOI21X1  g03353(.A0(new_n2125_), .A1(new_n668_), .B0(new_n3609_), .Y(new_n3610_));
  XOR2X1   g03354(.A(new_n3610_), .B(new_n665_), .Y(new_n3611_));
  XOR2X1   g03355(.A(new_n3544_), .B(new_n879_), .Y(new_n3612_));
  AND2X1   g03356(.A(new_n3612_), .B(new_n3541_), .Y(new_n3613_));
  AOI21X1  g03357(.A0(new_n3552_), .A1(new_n3550_), .B0(new_n3546_), .Y(new_n3614_));
  OR2X1    g03358(.A(new_n3614_), .B(new_n3613_), .Y(new_n3615_));
  INVX1    g03359(.A(new_n3529_), .Y(new_n3616_));
  XOR2X1   g03360(.A(new_n3532_), .B(new_n3616_), .Y(new_n3617_));
  OR2X1    g03361(.A(new_n3537_), .B(new_n3617_), .Y(new_n3618_));
  OAI21X1  g03362(.A0(new_n3540_), .A1(new_n3538_), .B0(new_n3618_), .Y(new_n3619_));
  INVX1    g03363(.A(new_n3512_), .Y(new_n3620_));
  XOR2X1   g03364(.A(new_n3620_), .B(new_n3508_), .Y(new_n3621_));
  XOR2X1   g03365(.A(new_n3621_), .B(new_n3465_), .Y(new_n3622_));
  OR2X1    g03366(.A(new_n3518_), .B(new_n3622_), .Y(new_n3623_));
  OAI21X1  g03367(.A0(new_n3523_), .A1(new_n3519_), .B0(new_n3623_), .Y(new_n3624_));
  AOI22X1  g03368(.A0(new_n1814_), .A1(\b[17] ), .B0(new_n1813_), .B1(\b[16] ), .Y(new_n3625_));
  OAI21X1  g03369(.A0(new_n1812_), .A1(new_n977_), .B0(new_n3625_), .Y(new_n3626_));
  AOI21X1  g03370(.A0(new_n1617_), .A1(new_n976_), .B0(new_n3626_), .Y(new_n3627_));
  XOR2X1   g03371(.A(new_n3627_), .B(\a[26] ), .Y(new_n3628_));
  AOI21X1  g03372(.A0(new_n3507_), .A1(new_n3506_), .B0(new_n3512_), .Y(new_n3629_));
  AOI21X1  g03373(.A0(new_n3513_), .A1(new_n3465_), .B0(new_n3629_), .Y(new_n3630_));
  AOI22X1  g03374(.A0(new_n2163_), .A1(\b[14] ), .B0(new_n2162_), .B1(\b[13] ), .Y(new_n3631_));
  OAI21X1  g03375(.A0(new_n2161_), .A1(new_n713_), .B0(new_n3631_), .Y(new_n3632_));
  AOI21X1  g03376(.A0(new_n1907_), .A1(new_n734_), .B0(new_n3632_), .Y(new_n3633_));
  XOR2X1   g03377(.A(new_n3633_), .B(\a[29] ), .Y(new_n3634_));
  INVX1    g03378(.A(new_n3634_), .Y(new_n3635_));
  AOI21X1  g03379(.A0(new_n3344_), .A1(new_n3342_), .B0(new_n3467_), .Y(new_n3636_));
  OR2X1    g03380(.A(new_n3503_), .B(new_n3499_), .Y(new_n3637_));
  OAI21X1  g03381(.A0(new_n3505_), .A1(new_n3636_), .B0(new_n3637_), .Y(new_n3638_));
  XOR2X1   g03382(.A(new_n3492_), .B(new_n2650_), .Y(new_n3639_));
  NAND2X1  g03383(.A(new_n3639_), .B(new_n3489_), .Y(new_n3640_));
  OAI21X1  g03384(.A0(new_n3498_), .A1(new_n3494_), .B0(new_n3640_), .Y(new_n3641_));
  AOI22X1  g03385(.A0(new_n2813_), .A1(\b[8] ), .B0(new_n2812_), .B1(\b[7] ), .Y(new_n3642_));
  OAI21X1  g03386(.A0(new_n2946_), .A1(new_n392_), .B0(new_n3642_), .Y(new_n3643_));
  AOI21X1  g03387(.A0(new_n2652_), .A1(new_n454_), .B0(new_n3643_), .Y(new_n3644_));
  XOR2X1   g03388(.A(new_n3644_), .B(\a[35] ), .Y(new_n3645_));
  AND2X1   g03389(.A(new_n3487_), .B(new_n3475_), .Y(new_n3646_));
  AOI21X1  g03390(.A0(new_n3488_), .A1(new_n3470_), .B0(new_n3646_), .Y(new_n3647_));
  NAND3X1  g03391(.A(new_n3485_), .B(new_n3317_), .C(\a[41] ), .Y(new_n3648_));
  NAND2X1  g03392(.A(new_n3480_), .B(new_n341_), .Y(new_n3649_));
  OR4X1    g03393(.A(new_n3481_), .B(new_n3479_), .C(new_n3316_), .D(new_n274_), .Y(new_n3650_));
  AND2X1   g03394(.A(new_n3481_), .B(new_n3477_), .Y(new_n3651_));
  AND2X1   g03395(.A(new_n3479_), .B(new_n3316_), .Y(new_n3652_));
  AOI22X1  g03396(.A0(new_n3652_), .A1(\b[2] ), .B0(new_n3651_), .B1(\b[1] ), .Y(new_n3653_));
  NAND3X1  g03397(.A(new_n3653_), .B(new_n3650_), .C(new_n3649_), .Y(new_n3654_));
  XOR2X1   g03398(.A(new_n3654_), .B(new_n3478_), .Y(new_n3655_));
  XOR2X1   g03399(.A(new_n3655_), .B(new_n3648_), .Y(new_n3656_));
  AOI22X1  g03400(.A0(new_n3204_), .A1(\b[5] ), .B0(new_n3203_), .B1(\b[4] ), .Y(new_n3657_));
  OAI21X1  g03401(.A0(new_n3321_), .A1(new_n297_), .B0(new_n3657_), .Y(new_n3658_));
  AOI21X1  g03402(.A0(new_n3080_), .A1(new_n349_), .B0(new_n3658_), .Y(new_n3659_));
  XOR2X1   g03403(.A(new_n3659_), .B(\a[38] ), .Y(new_n3660_));
  XOR2X1   g03404(.A(new_n3660_), .B(new_n3656_), .Y(new_n3661_));
  XOR2X1   g03405(.A(new_n3661_), .B(new_n3647_), .Y(new_n3662_));
  XOR2X1   g03406(.A(new_n3662_), .B(new_n3645_), .Y(new_n3663_));
  XOR2X1   g03407(.A(new_n3663_), .B(new_n3641_), .Y(new_n3664_));
  AOI22X1  g03408(.A0(new_n2545_), .A1(\b[11] ), .B0(new_n2544_), .B1(\b[10] ), .Y(new_n3665_));
  OAI21X1  g03409(.A0(new_n2543_), .A1(new_n590_), .B0(new_n3665_), .Y(new_n3666_));
  AOI21X1  g03410(.A0(new_n2260_), .A1(new_n589_), .B0(new_n3666_), .Y(new_n3667_));
  XOR2X1   g03411(.A(new_n3667_), .B(\a[32] ), .Y(new_n3668_));
  XOR2X1   g03412(.A(new_n3668_), .B(new_n3664_), .Y(new_n3669_));
  XOR2X1   g03413(.A(new_n3669_), .B(new_n3638_), .Y(new_n3670_));
  XOR2X1   g03414(.A(new_n3670_), .B(new_n3635_), .Y(new_n3671_));
  INVX1    g03415(.A(new_n3671_), .Y(new_n3672_));
  XOR2X1   g03416(.A(new_n3672_), .B(new_n3630_), .Y(new_n3673_));
  XOR2X1   g03417(.A(new_n3673_), .B(new_n3628_), .Y(new_n3674_));
  XOR2X1   g03418(.A(new_n3674_), .B(new_n3624_), .Y(new_n3675_));
  AOI22X1  g03419(.A0(new_n1526_), .A1(\b[20] ), .B0(new_n1525_), .B1(\b[19] ), .Y(new_n3676_));
  OAI21X1  g03420(.A0(new_n1524_), .A1(new_n1115_), .B0(new_n3676_), .Y(new_n3677_));
  AOI21X1  g03421(.A0(new_n1347_), .A1(new_n1217_), .B0(new_n3677_), .Y(new_n3678_));
  XOR2X1   g03422(.A(new_n3678_), .B(\a[23] ), .Y(new_n3679_));
  XOR2X1   g03423(.A(new_n3679_), .B(new_n3675_), .Y(new_n3680_));
  INVX1    g03424(.A(new_n3524_), .Y(new_n3681_));
  NOR2X1   g03425(.A(new_n3528_), .B(new_n3681_), .Y(new_n3682_));
  AOI21X1  g03426(.A0(new_n3531_), .A1(new_n3530_), .B0(new_n3529_), .Y(new_n3683_));
  NOR2X1   g03427(.A(new_n3683_), .B(new_n3682_), .Y(new_n3684_));
  XOR2X1   g03428(.A(new_n3684_), .B(new_n3680_), .Y(new_n3685_));
  AOI22X1  g03429(.A0(new_n1263_), .A1(\b[23] ), .B0(new_n1262_), .B1(\b[22] ), .Y(new_n3686_));
  OAI21X1  g03430(.A0(new_n1261_), .A1(new_n1482_), .B0(new_n3686_), .Y(new_n3687_));
  AOI21X1  g03431(.A0(new_n1481_), .A1(new_n1075_), .B0(new_n3687_), .Y(new_n3688_));
  XOR2X1   g03432(.A(new_n3688_), .B(\a[20] ), .Y(new_n3689_));
  NAND2X1  g03433(.A(new_n3689_), .B(new_n3685_), .Y(new_n3690_));
  XOR2X1   g03434(.A(new_n3689_), .B(new_n3685_), .Y(new_n3691_));
  NAND2X1  g03435(.A(new_n3691_), .B(new_n3619_), .Y(new_n3692_));
  NOR2X1   g03436(.A(new_n3689_), .B(new_n3685_), .Y(new_n3693_));
  AOI21X1  g03437(.A0(new_n3690_), .A1(new_n3619_), .B0(new_n3693_), .Y(new_n3694_));
  AOI22X1  g03438(.A0(new_n3694_), .A1(new_n3690_), .B0(new_n3692_), .B1(new_n3619_), .Y(new_n3695_));
  AOI22X1  g03439(.A0(new_n1017_), .A1(\b[26] ), .B0(new_n1016_), .B1(\b[25] ), .Y(new_n3696_));
  OAI21X1  g03440(.A0(new_n1015_), .A1(new_n1588_), .B0(new_n3696_), .Y(new_n3697_));
  AOI21X1  g03441(.A0(new_n1783_), .A1(new_n882_), .B0(new_n3697_), .Y(new_n3698_));
  XOR2X1   g03442(.A(new_n3698_), .B(\a[17] ), .Y(new_n3699_));
  XOR2X1   g03443(.A(new_n3699_), .B(new_n3695_), .Y(new_n3700_));
  XOR2X1   g03444(.A(new_n3700_), .B(new_n3615_), .Y(new_n3701_));
  XOR2X1   g03445(.A(new_n3701_), .B(new_n3611_), .Y(new_n3702_));
  XOR2X1   g03446(.A(new_n3702_), .B(new_n3607_), .Y(new_n3703_));
  XOR2X1   g03447(.A(new_n3703_), .B(new_n3603_), .Y(new_n3704_));
  XOR2X1   g03448(.A(new_n3704_), .B(new_n3599_), .Y(new_n3705_));
  AOI22X1  g03449(.A0(new_n469_), .A1(\b[35] ), .B0(new_n468_), .B1(\b[34] ), .Y(new_n3706_));
  OAI21X1  g03450(.A0(new_n467_), .A1(new_n2893_), .B0(new_n3706_), .Y(new_n3707_));
  AOI21X1  g03451(.A0(new_n2892_), .A1(new_n404_), .B0(new_n3707_), .Y(new_n3708_));
  XOR2X1   g03452(.A(new_n3708_), .B(\a[8] ), .Y(new_n3709_));
  XOR2X1   g03453(.A(new_n3709_), .B(new_n3705_), .Y(new_n3710_));
  XOR2X1   g03454(.A(new_n3710_), .B(new_n3597_), .Y(new_n3711_));
  AOI22X1  g03455(.A0(new_n369_), .A1(\b[38] ), .B0(new_n368_), .B1(\b[37] ), .Y(new_n3712_));
  OAI21X1  g03456(.A0(new_n367_), .A1(new_n3276_), .B0(new_n3712_), .Y(new_n3713_));
  AOI21X1  g03457(.A0(new_n3275_), .A1(new_n308_), .B0(new_n3713_), .Y(new_n3714_));
  XOR2X1   g03458(.A(new_n3714_), .B(\a[5] ), .Y(new_n3715_));
  XOR2X1   g03459(.A(new_n3715_), .B(new_n3711_), .Y(new_n3716_));
  XOR2X1   g03460(.A(new_n3716_), .B(new_n3595_), .Y(new_n3717_));
  AND2X1   g03461(.A(\b[40] ), .B(\b[39] ), .Y(new_n3718_));
  AOI21X1  g03462(.A0(new_n3573_), .A1(new_n3572_), .B0(new_n3718_), .Y(new_n3719_));
  INVX1    g03463(.A(\b[40] ), .Y(new_n3720_));
  XOR2X1   g03464(.A(\b[41] ), .B(new_n3720_), .Y(new_n3721_));
  XOR2X1   g03465(.A(new_n3721_), .B(new_n3719_), .Y(new_n3722_));
  INVX1    g03466(.A(\b[39] ), .Y(new_n3723_));
  AOI22X1  g03467(.A0(new_n267_), .A1(\b[41] ), .B0(new_n266_), .B1(\b[40] ), .Y(new_n3724_));
  OAI21X1  g03468(.A0(new_n350_), .A1(new_n3723_), .B0(new_n3724_), .Y(new_n3725_));
  AOI21X1  g03469(.A0(new_n3722_), .A1(new_n318_), .B0(new_n3725_), .Y(new_n3726_));
  XOR2X1   g03470(.A(new_n3726_), .B(\a[2] ), .Y(new_n3727_));
  XOR2X1   g03471(.A(new_n3727_), .B(new_n3717_), .Y(new_n3728_));
  XOR2X1   g03472(.A(new_n3728_), .B(new_n3588_), .Y(\f[41] ));
  OR2X1    g03473(.A(new_n3568_), .B(new_n3592_), .Y(new_n3730_));
  OAI21X1  g03474(.A0(new_n3569_), .A1(new_n3436_), .B0(new_n3730_), .Y(new_n3731_));
  NOR2X1   g03475(.A(new_n3715_), .B(new_n3711_), .Y(new_n3732_));
  AOI21X1  g03476(.A0(new_n3716_), .A1(new_n3731_), .B0(new_n3732_), .Y(new_n3733_));
  AOI22X1  g03477(.A0(new_n369_), .A1(\b[39] ), .B0(new_n368_), .B1(\b[38] ), .Y(new_n3734_));
  OAI21X1  g03478(.A0(new_n367_), .A1(new_n3413_), .B0(new_n3734_), .Y(new_n3735_));
  AOI21X1  g03479(.A0(new_n3412_), .A1(new_n308_), .B0(new_n3735_), .Y(new_n3736_));
  XOR2X1   g03480(.A(new_n3736_), .B(\a[5] ), .Y(new_n3737_));
  OR2X1    g03481(.A(new_n3709_), .B(new_n3705_), .Y(new_n3738_));
  NOR2X1   g03482(.A(new_n3393_), .B(new_n3389_), .Y(new_n3739_));
  AOI21X1  g03483(.A0(new_n3394_), .A1(new_n3304_), .B0(new_n3739_), .Y(new_n3740_));
  AND2X1   g03484(.A(new_n3560_), .B(new_n3556_), .Y(new_n3741_));
  OR2X1    g03485(.A(new_n3560_), .B(new_n3556_), .Y(new_n3742_));
  OAI21X1  g03486(.A0(new_n3741_), .A1(new_n3740_), .B0(new_n3742_), .Y(new_n3743_));
  XOR2X1   g03487(.A(new_n3704_), .B(new_n3743_), .Y(new_n3744_));
  XOR2X1   g03488(.A(new_n3709_), .B(new_n3744_), .Y(new_n3745_));
  OAI21X1  g03489(.A0(new_n3745_), .A1(new_n3597_), .B0(new_n3738_), .Y(new_n3746_));
  NOR2X1   g03490(.A(new_n3703_), .B(new_n3603_), .Y(new_n3747_));
  NAND2X1  g03491(.A(new_n3703_), .B(new_n3603_), .Y(new_n3748_));
  OAI21X1  g03492(.A0(new_n3747_), .A1(new_n3599_), .B0(new_n3748_), .Y(new_n3749_));
  NAND2X1  g03493(.A(new_n3701_), .B(new_n3611_), .Y(new_n3750_));
  OAI21X1  g03494(.A0(new_n3606_), .A1(new_n3605_), .B0(new_n3702_), .Y(new_n3751_));
  NAND2X1  g03495(.A(new_n3751_), .B(new_n3750_), .Y(new_n3752_));
  NOR2X1   g03496(.A(new_n3699_), .B(new_n3695_), .Y(new_n3753_));
  AOI21X1  g03497(.A0(new_n3700_), .A1(new_n3615_), .B0(new_n3753_), .Y(new_n3754_));
  INVX1    g03498(.A(new_n3628_), .Y(new_n3755_));
  AND2X1   g03499(.A(new_n3673_), .B(new_n3755_), .Y(new_n3756_));
  XOR2X1   g03500(.A(new_n3673_), .B(new_n3755_), .Y(new_n3757_));
  AOI21X1  g03501(.A0(new_n3757_), .A1(new_n3624_), .B0(new_n3756_), .Y(new_n3758_));
  AND2X1   g03502(.A(new_n3670_), .B(new_n3635_), .Y(new_n3759_));
  INVX1    g03503(.A(new_n3759_), .Y(new_n3760_));
  OAI21X1  g03504(.A0(new_n3672_), .A1(new_n3630_), .B0(new_n3760_), .Y(new_n3761_));
  NOR2X1   g03505(.A(new_n3668_), .B(new_n3664_), .Y(new_n3762_));
  AOI21X1  g03506(.A0(new_n3669_), .A1(new_n3638_), .B0(new_n3762_), .Y(new_n3763_));
  AOI22X1  g03507(.A0(new_n2545_), .A1(\b[12] ), .B0(new_n2544_), .B1(\b[11] ), .Y(new_n3764_));
  OAI21X1  g03508(.A0(new_n2543_), .A1(new_n587_), .B0(new_n3764_), .Y(new_n3765_));
  AOI21X1  g03509(.A0(new_n2260_), .A1(new_n635_), .B0(new_n3765_), .Y(new_n3766_));
  XOR2X1   g03510(.A(new_n3766_), .B(\a[32] ), .Y(new_n3767_));
  INVX1    g03511(.A(new_n3645_), .Y(new_n3768_));
  AND2X1   g03512(.A(new_n3662_), .B(new_n3768_), .Y(new_n3769_));
  INVX1    g03513(.A(new_n3663_), .Y(new_n3770_));
  AOI21X1  g03514(.A0(new_n3770_), .A1(new_n3641_), .B0(new_n3769_), .Y(new_n3771_));
  OR2X1    g03515(.A(new_n3655_), .B(new_n3648_), .Y(new_n3772_));
  XOR2X1   g03516(.A(\a[42] ), .B(\a[41] ), .Y(new_n3773_));
  NAND2X1  g03517(.A(new_n3773_), .B(\b[0] ), .Y(new_n3774_));
  INVX1    g03518(.A(new_n3774_), .Y(new_n3775_));
  XOR2X1   g03519(.A(new_n3775_), .B(new_n3772_), .Y(new_n3776_));
  OR2X1    g03520(.A(new_n3481_), .B(new_n3316_), .Y(new_n3777_));
  OR2X1    g03521(.A(new_n3777_), .B(new_n3479_), .Y(new_n3778_));
  AOI22X1  g03522(.A0(new_n3652_), .A1(\b[3] ), .B0(new_n3651_), .B1(\b[2] ), .Y(new_n3779_));
  OAI21X1  g03523(.A0(new_n3778_), .A1(new_n275_), .B0(new_n3779_), .Y(new_n3780_));
  AOI21X1  g03524(.A0(new_n3480_), .A1(new_n366_), .B0(new_n3780_), .Y(new_n3781_));
  XOR2X1   g03525(.A(new_n3781_), .B(\a[41] ), .Y(new_n3782_));
  XOR2X1   g03526(.A(new_n3782_), .B(new_n3776_), .Y(new_n3783_));
  AOI22X1  g03527(.A0(new_n3204_), .A1(\b[6] ), .B0(new_n3203_), .B1(\b[5] ), .Y(new_n3784_));
  OAI21X1  g03528(.A0(new_n3321_), .A1(new_n325_), .B0(new_n3784_), .Y(new_n3785_));
  AOI21X1  g03529(.A0(new_n3080_), .A1(new_n378_), .B0(new_n3785_), .Y(new_n3786_));
  XOR2X1   g03530(.A(new_n3786_), .B(\a[38] ), .Y(new_n3787_));
  XOR2X1   g03531(.A(new_n3787_), .B(new_n3783_), .Y(new_n3788_));
  INVX1    g03532(.A(new_n3660_), .Y(new_n3789_));
  NOR2X1   g03533(.A(new_n3661_), .B(new_n3647_), .Y(new_n3790_));
  AOI21X1  g03534(.A0(new_n3789_), .A1(new_n3656_), .B0(new_n3790_), .Y(new_n3791_));
  XOR2X1   g03535(.A(new_n3791_), .B(new_n3788_), .Y(new_n3792_));
  AOI22X1  g03536(.A0(new_n2813_), .A1(\b[9] ), .B0(new_n2812_), .B1(\b[8] ), .Y(new_n3793_));
  OAI21X1  g03537(.A0(new_n2946_), .A1(new_n492_), .B0(new_n3793_), .Y(new_n3794_));
  AOI21X1  g03538(.A0(new_n2652_), .A1(new_n491_), .B0(new_n3794_), .Y(new_n3795_));
  XOR2X1   g03539(.A(new_n3795_), .B(\a[35] ), .Y(new_n3796_));
  XOR2X1   g03540(.A(new_n3796_), .B(new_n3792_), .Y(new_n3797_));
  XOR2X1   g03541(.A(new_n3797_), .B(new_n3771_), .Y(new_n3798_));
  XOR2X1   g03542(.A(new_n3798_), .B(new_n3767_), .Y(new_n3799_));
  XOR2X1   g03543(.A(new_n3799_), .B(new_n3763_), .Y(new_n3800_));
  AOI22X1  g03544(.A0(new_n2163_), .A1(\b[15] ), .B0(new_n2162_), .B1(\b[14] ), .Y(new_n3801_));
  OAI21X1  g03545(.A0(new_n2161_), .A1(new_n795_), .B0(new_n3801_), .Y(new_n3802_));
  AOI21X1  g03546(.A0(new_n1907_), .A1(new_n794_), .B0(new_n3802_), .Y(new_n3803_));
  XOR2X1   g03547(.A(new_n3803_), .B(\a[29] ), .Y(new_n3804_));
  XOR2X1   g03548(.A(new_n3804_), .B(new_n3800_), .Y(new_n3805_));
  XOR2X1   g03549(.A(new_n3805_), .B(new_n3761_), .Y(new_n3806_));
  AOI22X1  g03550(.A0(new_n1814_), .A1(\b[18] ), .B0(new_n1813_), .B1(\b[17] ), .Y(new_n3807_));
  OAI21X1  g03551(.A0(new_n1812_), .A1(new_n974_), .B0(new_n3807_), .Y(new_n3808_));
  AOI21X1  g03552(.A0(new_n1617_), .A1(new_n1042_), .B0(new_n3808_), .Y(new_n3809_));
  XOR2X1   g03553(.A(new_n3809_), .B(\a[26] ), .Y(new_n3810_));
  XOR2X1   g03554(.A(new_n3810_), .B(new_n3806_), .Y(new_n3811_));
  XOR2X1   g03555(.A(new_n3811_), .B(new_n3758_), .Y(new_n3812_));
  AOI22X1  g03556(.A0(new_n1526_), .A1(\b[21] ), .B0(new_n1525_), .B1(\b[20] ), .Y(new_n3813_));
  OAI21X1  g03557(.A0(new_n1524_), .A1(new_n1300_), .B0(new_n3813_), .Y(new_n3814_));
  AOI21X1  g03558(.A0(new_n1347_), .A1(new_n1299_), .B0(new_n3814_), .Y(new_n3815_));
  XOR2X1   g03559(.A(new_n3815_), .B(\a[23] ), .Y(new_n3816_));
  INVX1    g03560(.A(new_n3816_), .Y(new_n3817_));
  XOR2X1   g03561(.A(new_n3817_), .B(new_n3812_), .Y(new_n3818_));
  OR2X1    g03562(.A(new_n3679_), .B(new_n3675_), .Y(new_n3819_));
  OAI21X1  g03563(.A0(new_n3683_), .A1(new_n3682_), .B0(new_n3680_), .Y(new_n3820_));
  NAND2X1  g03564(.A(new_n3820_), .B(new_n3819_), .Y(new_n3821_));
  XOR2X1   g03565(.A(new_n3821_), .B(new_n3818_), .Y(new_n3822_));
  AOI22X1  g03566(.A0(new_n1263_), .A1(\b[24] ), .B0(new_n1262_), .B1(\b[23] ), .Y(new_n3823_));
  OAI21X1  g03567(.A0(new_n1261_), .A1(new_n1479_), .B0(new_n3823_), .Y(new_n3824_));
  AOI21X1  g03568(.A0(new_n1572_), .A1(new_n1075_), .B0(new_n3824_), .Y(new_n3825_));
  XOR2X1   g03569(.A(new_n3825_), .B(\a[20] ), .Y(new_n3826_));
  XOR2X1   g03570(.A(new_n3826_), .B(new_n3822_), .Y(new_n3827_));
  XOR2X1   g03571(.A(new_n3827_), .B(new_n3694_), .Y(new_n3828_));
  AOI22X1  g03572(.A0(new_n1017_), .A1(\b[27] ), .B0(new_n1016_), .B1(\b[26] ), .Y(new_n3829_));
  OAI21X1  g03573(.A0(new_n1015_), .A1(new_n1880_), .B0(new_n3829_), .Y(new_n3830_));
  AOI21X1  g03574(.A0(new_n1879_), .A1(new_n882_), .B0(new_n3830_), .Y(new_n3831_));
  XOR2X1   g03575(.A(new_n3831_), .B(\a[17] ), .Y(new_n3832_));
  INVX1    g03576(.A(new_n3832_), .Y(new_n3833_));
  XOR2X1   g03577(.A(new_n3833_), .B(new_n3828_), .Y(new_n3834_));
  INVX1    g03578(.A(new_n3834_), .Y(new_n3835_));
  XOR2X1   g03579(.A(new_n3835_), .B(new_n3754_), .Y(new_n3836_));
  AOI22X1  g03580(.A0(new_n818_), .A1(\b[30] ), .B0(new_n817_), .B1(\b[29] ), .Y(new_n3837_));
  OAI21X1  g03581(.A0(new_n816_), .A1(new_n2231_), .B0(new_n3837_), .Y(new_n3838_));
  AOI21X1  g03582(.A0(new_n2230_), .A1(new_n668_), .B0(new_n3838_), .Y(new_n3839_));
  XOR2X1   g03583(.A(new_n3839_), .B(\a[14] ), .Y(new_n3840_));
  XOR2X1   g03584(.A(new_n3840_), .B(new_n3836_), .Y(new_n3841_));
  XOR2X1   g03585(.A(new_n3841_), .B(new_n3752_), .Y(new_n3842_));
  AOI22X1  g03586(.A0(new_n603_), .A1(\b[33] ), .B0(new_n602_), .B1(\b[32] ), .Y(new_n3843_));
  OAI21X1  g03587(.A0(new_n601_), .A1(new_n2615_), .B0(new_n3843_), .Y(new_n3844_));
  AOI21X1  g03588(.A0(new_n2614_), .A1(new_n518_), .B0(new_n3844_), .Y(new_n3845_));
  XOR2X1   g03589(.A(new_n3845_), .B(\a[11] ), .Y(new_n3846_));
  XOR2X1   g03590(.A(new_n3846_), .B(new_n3842_), .Y(new_n3847_));
  XOR2X1   g03591(.A(new_n3847_), .B(new_n3749_), .Y(new_n3848_));
  AOI22X1  g03592(.A0(new_n469_), .A1(\b[36] ), .B0(new_n468_), .B1(\b[35] ), .Y(new_n3849_));
  OAI21X1  g03593(.A0(new_n467_), .A1(new_n2890_), .B0(new_n3849_), .Y(new_n3850_));
  AOI21X1  g03594(.A0(new_n3015_), .A1(new_n404_), .B0(new_n3850_), .Y(new_n3851_));
  XOR2X1   g03595(.A(new_n3851_), .B(\a[8] ), .Y(new_n3852_));
  XOR2X1   g03596(.A(new_n3852_), .B(new_n3848_), .Y(new_n3853_));
  XOR2X1   g03597(.A(new_n3853_), .B(new_n3746_), .Y(new_n3854_));
  XOR2X1   g03598(.A(new_n3854_), .B(new_n3737_), .Y(new_n3855_));
  XOR2X1   g03599(.A(new_n3855_), .B(new_n3733_), .Y(new_n3856_));
  NAND2X1  g03600(.A(\b[41] ), .B(\b[40] ), .Y(new_n3857_));
  OAI21X1  g03601(.A0(new_n3721_), .A1(new_n3719_), .B0(new_n3857_), .Y(new_n3858_));
  XOR2X1   g03602(.A(\b[42] ), .B(\b[41] ), .Y(new_n3859_));
  XOR2X1   g03603(.A(new_n3859_), .B(new_n3858_), .Y(new_n3860_));
  AOI22X1  g03604(.A0(new_n267_), .A1(\b[42] ), .B0(new_n266_), .B1(\b[41] ), .Y(new_n3861_));
  OAI21X1  g03605(.A0(new_n350_), .A1(new_n3720_), .B0(new_n3861_), .Y(new_n3862_));
  AOI21X1  g03606(.A0(new_n3860_), .A1(new_n318_), .B0(new_n3862_), .Y(new_n3863_));
  XOR2X1   g03607(.A(new_n3863_), .B(\a[2] ), .Y(new_n3864_));
  XOR2X1   g03608(.A(new_n3864_), .B(new_n3856_), .Y(new_n3865_));
  OR2X1    g03609(.A(new_n3727_), .B(new_n3717_), .Y(new_n3866_));
  OAI21X1  g03610(.A0(new_n3587_), .A1(new_n3586_), .B0(new_n3728_), .Y(new_n3867_));
  AND2X1   g03611(.A(new_n3867_), .B(new_n3866_), .Y(new_n3868_));
  XOR2X1   g03612(.A(new_n3868_), .B(new_n3865_), .Y(\f[42] ));
  INVX1    g03613(.A(new_n3737_), .Y(new_n3870_));
  NAND2X1  g03614(.A(new_n3854_), .B(new_n3870_), .Y(new_n3871_));
  OAI21X1  g03615(.A0(new_n3855_), .A1(new_n3733_), .B0(new_n3871_), .Y(new_n3872_));
  NOR2X1   g03616(.A(new_n3852_), .B(new_n3848_), .Y(new_n3873_));
  AOI21X1  g03617(.A0(new_n3853_), .A1(new_n3746_), .B0(new_n3873_), .Y(new_n3874_));
  NOR2X1   g03618(.A(new_n3840_), .B(new_n3836_), .Y(new_n3875_));
  AOI21X1  g03619(.A0(new_n3841_), .A1(new_n3752_), .B0(new_n3875_), .Y(new_n3876_));
  OR2X1    g03620(.A(new_n3832_), .B(new_n3828_), .Y(new_n3877_));
  OAI21X1  g03621(.A0(new_n3834_), .A1(new_n3754_), .B0(new_n3877_), .Y(new_n3878_));
  AOI22X1  g03622(.A0(new_n1017_), .A1(\b[28] ), .B0(new_n1016_), .B1(\b[27] ), .Y(new_n3879_));
  OAI21X1  g03623(.A0(new_n1015_), .A1(new_n1877_), .B0(new_n3879_), .Y(new_n3880_));
  AOI21X1  g03624(.A0(new_n2004_), .A1(new_n882_), .B0(new_n3880_), .Y(new_n3881_));
  XOR2X1   g03625(.A(new_n3881_), .B(\a[17] ), .Y(new_n3882_));
  INVX1    g03626(.A(new_n3767_), .Y(new_n3883_));
  AND2X1   g03627(.A(new_n3798_), .B(new_n3883_), .Y(new_n3884_));
  NOR2X1   g03628(.A(new_n3799_), .B(new_n3763_), .Y(new_n3885_));
  OR2X1    g03629(.A(new_n3885_), .B(new_n3884_), .Y(new_n3886_));
  XOR2X1   g03630(.A(new_n3795_), .B(new_n2650_), .Y(new_n3887_));
  NAND2X1  g03631(.A(new_n3887_), .B(new_n3792_), .Y(new_n3888_));
  OAI21X1  g03632(.A0(new_n3797_), .A1(new_n3771_), .B0(new_n3888_), .Y(new_n3889_));
  OR4X1    g03633(.A(new_n3774_), .B(new_n3655_), .C(new_n3486_), .D(new_n3476_), .Y(new_n3890_));
  OAI21X1  g03634(.A0(new_n3782_), .A1(new_n3776_), .B0(new_n3890_), .Y(new_n3891_));
  AND2X1   g03635(.A(new_n3480_), .B(new_n323_), .Y(new_n3892_));
  NOR3X1   g03636(.A(new_n3777_), .B(new_n3479_), .C(new_n277_), .Y(new_n3893_));
  OAI22X1  g03637(.A0(new_n3483_), .A1(new_n325_), .B0(new_n3482_), .B1(new_n297_), .Y(new_n3894_));
  NOR3X1   g03638(.A(new_n3894_), .B(new_n3893_), .C(new_n3892_), .Y(new_n3895_));
  XOR2X1   g03639(.A(new_n3895_), .B(new_n3478_), .Y(new_n3896_));
  NAND2X1  g03640(.A(new_n3774_), .B(\a[44] ), .Y(new_n3897_));
  XOR2X1   g03641(.A(\a[42] ), .B(new_n3478_), .Y(new_n3898_));
  INVX1    g03642(.A(\a[44] ), .Y(new_n3899_));
  XOR2X1   g03643(.A(new_n3899_), .B(\a[43] ), .Y(new_n3900_));
  NOR2X1   g03644(.A(new_n3900_), .B(new_n3898_), .Y(new_n3901_));
  XOR2X1   g03645(.A(\a[43] ), .B(\a[42] ), .Y(new_n3902_));
  NAND2X1  g03646(.A(new_n3902_), .B(new_n3898_), .Y(new_n3903_));
  NAND2X1  g03647(.A(new_n3900_), .B(new_n3773_), .Y(new_n3904_));
  OAI22X1  g03648(.A0(new_n3904_), .A1(new_n275_), .B0(new_n3903_), .B1(new_n274_), .Y(new_n3905_));
  AOI21X1  g03649(.A0(new_n3901_), .A1(new_n263_), .B0(new_n3905_), .Y(new_n3906_));
  XOR2X1   g03650(.A(new_n3906_), .B(\a[44] ), .Y(new_n3907_));
  XOR2X1   g03651(.A(new_n3907_), .B(new_n3897_), .Y(new_n3908_));
  XOR2X1   g03652(.A(new_n3908_), .B(new_n3896_), .Y(new_n3909_));
  XOR2X1   g03653(.A(new_n3909_), .B(new_n3891_), .Y(new_n3910_));
  AOI22X1  g03654(.A0(new_n3204_), .A1(\b[7] ), .B0(new_n3203_), .B1(\b[6] ), .Y(new_n3911_));
  OAI21X1  g03655(.A0(new_n3321_), .A1(new_n395_), .B0(new_n3911_), .Y(new_n3912_));
  AOI21X1  g03656(.A0(new_n3080_), .A1(new_n394_), .B0(new_n3912_), .Y(new_n3913_));
  XOR2X1   g03657(.A(new_n3913_), .B(\a[38] ), .Y(new_n3914_));
  XOR2X1   g03658(.A(new_n3914_), .B(new_n3910_), .Y(new_n3915_));
  INVX1    g03659(.A(new_n3915_), .Y(new_n3916_));
  INVX1    g03660(.A(new_n3787_), .Y(new_n3917_));
  NOR2X1   g03661(.A(new_n3791_), .B(new_n3788_), .Y(new_n3918_));
  AOI21X1  g03662(.A0(new_n3917_), .A1(new_n3783_), .B0(new_n3918_), .Y(new_n3919_));
  XOR2X1   g03663(.A(new_n3919_), .B(new_n3916_), .Y(new_n3920_));
  AOI22X1  g03664(.A0(new_n2813_), .A1(\b[10] ), .B0(new_n2812_), .B1(\b[9] ), .Y(new_n3921_));
  OAI21X1  g03665(.A0(new_n2946_), .A1(new_n489_), .B0(new_n3921_), .Y(new_n3922_));
  AOI21X1  g03666(.A0(new_n2652_), .A1(new_n543_), .B0(new_n3922_), .Y(new_n3923_));
  XOR2X1   g03667(.A(new_n3923_), .B(\a[35] ), .Y(new_n3924_));
  NAND2X1  g03668(.A(new_n3924_), .B(new_n3920_), .Y(new_n3925_));
  XOR2X1   g03669(.A(new_n3924_), .B(new_n3920_), .Y(new_n3926_));
  INVX1    g03670(.A(new_n3926_), .Y(new_n3927_));
  NOR2X1   g03671(.A(new_n3924_), .B(new_n3920_), .Y(new_n3928_));
  AOI21X1  g03672(.A0(new_n3925_), .A1(new_n3889_), .B0(new_n3928_), .Y(new_n3929_));
  AOI22X1  g03673(.A0(new_n3929_), .A1(new_n3925_), .B0(new_n3927_), .B1(new_n3889_), .Y(new_n3930_));
  AOI22X1  g03674(.A0(new_n2545_), .A1(\b[13] ), .B0(new_n2544_), .B1(\b[12] ), .Y(new_n3931_));
  OAI21X1  g03675(.A0(new_n2543_), .A1(new_n716_), .B0(new_n3931_), .Y(new_n3932_));
  AOI21X1  g03676(.A0(new_n2260_), .A1(new_n715_), .B0(new_n3932_), .Y(new_n3933_));
  XOR2X1   g03677(.A(new_n3933_), .B(\a[32] ), .Y(new_n3934_));
  XOR2X1   g03678(.A(new_n3934_), .B(new_n3930_), .Y(new_n3935_));
  XOR2X1   g03679(.A(new_n3935_), .B(new_n3886_), .Y(new_n3936_));
  AOI22X1  g03680(.A0(new_n2163_), .A1(\b[16] ), .B0(new_n2162_), .B1(\b[15] ), .Y(new_n3937_));
  OAI21X1  g03681(.A0(new_n2161_), .A1(new_n792_), .B0(new_n3937_), .Y(new_n3938_));
  AOI21X1  g03682(.A0(new_n1907_), .A1(new_n842_), .B0(new_n3938_), .Y(new_n3939_));
  XOR2X1   g03683(.A(new_n3939_), .B(\a[29] ), .Y(new_n3940_));
  XOR2X1   g03684(.A(new_n3940_), .B(new_n3936_), .Y(new_n3941_));
  XOR2X1   g03685(.A(new_n3803_), .B(new_n1911_), .Y(new_n3942_));
  AND2X1   g03686(.A(new_n3942_), .B(new_n3800_), .Y(new_n3943_));
  INVX1    g03687(.A(new_n3805_), .Y(new_n3944_));
  AOI21X1  g03688(.A0(new_n3944_), .A1(new_n3761_), .B0(new_n3943_), .Y(new_n3945_));
  XOR2X1   g03689(.A(new_n3945_), .B(new_n3941_), .Y(new_n3946_));
  AOI22X1  g03690(.A0(new_n1814_), .A1(\b[19] ), .B0(new_n1813_), .B1(\b[18] ), .Y(new_n3947_));
  OAI21X1  g03691(.A0(new_n1812_), .A1(new_n1118_), .B0(new_n3947_), .Y(new_n3948_));
  AOI21X1  g03692(.A0(new_n1617_), .A1(new_n1117_), .B0(new_n3948_), .Y(new_n3949_));
  XOR2X1   g03693(.A(new_n3949_), .B(\a[26] ), .Y(new_n3950_));
  XOR2X1   g03694(.A(new_n3950_), .B(new_n3946_), .Y(new_n3951_));
  OR2X1    g03695(.A(new_n3810_), .B(new_n3806_), .Y(new_n3952_));
  AND2X1   g03696(.A(new_n3810_), .B(new_n3806_), .Y(new_n3953_));
  OAI21X1  g03697(.A0(new_n3953_), .A1(new_n3758_), .B0(new_n3952_), .Y(new_n3954_));
  XOR2X1   g03698(.A(new_n3954_), .B(new_n3951_), .Y(new_n3955_));
  AOI22X1  g03699(.A0(new_n1526_), .A1(\b[22] ), .B0(new_n1525_), .B1(\b[21] ), .Y(new_n3956_));
  OAI21X1  g03700(.A0(new_n1524_), .A1(new_n1297_), .B0(new_n3956_), .Y(new_n3957_));
  AOI21X1  g03701(.A0(new_n1399_), .A1(new_n1347_), .B0(new_n3957_), .Y(new_n3958_));
  XOR2X1   g03702(.A(new_n3958_), .B(\a[23] ), .Y(new_n3959_));
  XOR2X1   g03703(.A(new_n3959_), .B(new_n3955_), .Y(new_n3960_));
  INVX1    g03704(.A(new_n3960_), .Y(new_n3961_));
  NOR2X1   g03705(.A(new_n3816_), .B(new_n3812_), .Y(new_n3962_));
  AOI21X1  g03706(.A0(new_n3820_), .A1(new_n3819_), .B0(new_n3818_), .Y(new_n3963_));
  NOR2X1   g03707(.A(new_n3963_), .B(new_n3962_), .Y(new_n3964_));
  XOR2X1   g03708(.A(new_n3964_), .B(new_n3961_), .Y(new_n3965_));
  AOI22X1  g03709(.A0(new_n1263_), .A1(\b[25] ), .B0(new_n1262_), .B1(\b[24] ), .Y(new_n3966_));
  OAI21X1  g03710(.A0(new_n1261_), .A1(new_n1591_), .B0(new_n3966_), .Y(new_n3967_));
  AOI21X1  g03711(.A0(new_n1590_), .A1(new_n1075_), .B0(new_n3967_), .Y(new_n3968_));
  XOR2X1   g03712(.A(new_n3968_), .B(\a[20] ), .Y(new_n3969_));
  XOR2X1   g03713(.A(new_n3969_), .B(new_n3965_), .Y(new_n3970_));
  OR2X1    g03714(.A(new_n3826_), .B(new_n3822_), .Y(new_n3971_));
  AND2X1   g03715(.A(new_n3691_), .B(new_n3619_), .Y(new_n3972_));
  OAI21X1  g03716(.A0(new_n3972_), .A1(new_n3693_), .B0(new_n3827_), .Y(new_n3973_));
  AND2X1   g03717(.A(new_n3973_), .B(new_n3971_), .Y(new_n3974_));
  XOR2X1   g03718(.A(new_n3974_), .B(new_n3970_), .Y(new_n3975_));
  XOR2X1   g03719(.A(new_n3975_), .B(new_n3882_), .Y(new_n3976_));
  XOR2X1   g03720(.A(new_n3976_), .B(new_n3878_), .Y(new_n3977_));
  AOI22X1  g03721(.A0(new_n818_), .A1(\b[31] ), .B0(new_n817_), .B1(\b[30] ), .Y(new_n3978_));
  OAI21X1  g03722(.A0(new_n816_), .A1(new_n2359_), .B0(new_n3978_), .Y(new_n3979_));
  AOI21X1  g03723(.A0(new_n2358_), .A1(new_n668_), .B0(new_n3979_), .Y(new_n3980_));
  XOR2X1   g03724(.A(new_n3980_), .B(\a[14] ), .Y(new_n3981_));
  XOR2X1   g03725(.A(new_n3981_), .B(new_n3977_), .Y(new_n3982_));
  XOR2X1   g03726(.A(new_n3982_), .B(new_n3876_), .Y(new_n3983_));
  AOI22X1  g03727(.A0(new_n603_), .A1(\b[34] ), .B0(new_n602_), .B1(\b[33] ), .Y(new_n3984_));
  OAI21X1  g03728(.A0(new_n601_), .A1(new_n2612_), .B0(new_n3984_), .Y(new_n3985_));
  AOI21X1  g03729(.A0(new_n2759_), .A1(new_n518_), .B0(new_n3985_), .Y(new_n3986_));
  XOR2X1   g03730(.A(new_n3986_), .B(\a[11] ), .Y(new_n3987_));
  XOR2X1   g03731(.A(new_n3987_), .B(new_n3983_), .Y(new_n3988_));
  AND2X1   g03732(.A(new_n3751_), .B(new_n3750_), .Y(new_n3989_));
  XOR2X1   g03733(.A(new_n3841_), .B(new_n3989_), .Y(new_n3990_));
  NOR2X1   g03734(.A(new_n3846_), .B(new_n3990_), .Y(new_n3991_));
  XOR2X1   g03735(.A(new_n3846_), .B(new_n3990_), .Y(new_n3992_));
  AOI21X1  g03736(.A0(new_n3992_), .A1(new_n3749_), .B0(new_n3991_), .Y(new_n3993_));
  XOR2X1   g03737(.A(new_n3993_), .B(new_n3988_), .Y(new_n3994_));
  AOI22X1  g03738(.A0(new_n469_), .A1(\b[37] ), .B0(new_n468_), .B1(\b[36] ), .Y(new_n3995_));
  OAI21X1  g03739(.A0(new_n467_), .A1(new_n3156_), .B0(new_n3995_), .Y(new_n3996_));
  AOI21X1  g03740(.A0(new_n3155_), .A1(new_n404_), .B0(new_n3996_), .Y(new_n3997_));
  XOR2X1   g03741(.A(new_n3997_), .B(\a[8] ), .Y(new_n3998_));
  AND2X1   g03742(.A(new_n3998_), .B(new_n3994_), .Y(new_n3999_));
  XOR2X1   g03743(.A(new_n3998_), .B(new_n3994_), .Y(new_n4000_));
  OR2X1    g03744(.A(new_n3998_), .B(new_n3994_), .Y(new_n4001_));
  OAI21X1  g03745(.A0(new_n3999_), .A1(new_n3874_), .B0(new_n4001_), .Y(new_n4002_));
  OAI22X1  g03746(.A0(new_n4002_), .A1(new_n3999_), .B0(new_n4000_), .B1(new_n3874_), .Y(new_n4003_));
  AOI22X1  g03747(.A0(new_n369_), .A1(\b[40] ), .B0(new_n368_), .B1(\b[39] ), .Y(new_n4004_));
  OAI21X1  g03748(.A0(new_n367_), .A1(new_n3575_), .B0(new_n4004_), .Y(new_n4005_));
  AOI21X1  g03749(.A0(new_n3574_), .A1(new_n308_), .B0(new_n4005_), .Y(new_n4006_));
  XOR2X1   g03750(.A(new_n4006_), .B(new_n305_), .Y(new_n4007_));
  XOR2X1   g03751(.A(new_n4007_), .B(new_n4003_), .Y(new_n4008_));
  XOR2X1   g03752(.A(new_n4008_), .B(new_n3872_), .Y(new_n4009_));
  AND2X1   g03753(.A(\b[42] ), .B(\b[41] ), .Y(new_n4010_));
  AOI21X1  g03754(.A0(new_n3859_), .A1(new_n3858_), .B0(new_n4010_), .Y(new_n4011_));
  INVX1    g03755(.A(\b[42] ), .Y(new_n4012_));
  XOR2X1   g03756(.A(\b[43] ), .B(new_n4012_), .Y(new_n4013_));
  XOR2X1   g03757(.A(new_n4013_), .B(new_n4011_), .Y(new_n4014_));
  INVX1    g03758(.A(\b[41] ), .Y(new_n4015_));
  AOI22X1  g03759(.A0(new_n267_), .A1(\b[43] ), .B0(new_n266_), .B1(\b[42] ), .Y(new_n4016_));
  OAI21X1  g03760(.A0(new_n350_), .A1(new_n4015_), .B0(new_n4016_), .Y(new_n4017_));
  AOI21X1  g03761(.A0(new_n4014_), .A1(new_n318_), .B0(new_n4017_), .Y(new_n4018_));
  XOR2X1   g03762(.A(new_n4018_), .B(new_n257_), .Y(new_n4019_));
  XOR2X1   g03763(.A(new_n4019_), .B(new_n4009_), .Y(new_n4020_));
  OR2X1    g03764(.A(new_n3715_), .B(new_n3711_), .Y(new_n4021_));
  AND2X1   g03765(.A(new_n3715_), .B(new_n3711_), .Y(new_n4022_));
  OAI21X1  g03766(.A0(new_n4022_), .A1(new_n3595_), .B0(new_n4021_), .Y(new_n4023_));
  XOR2X1   g03767(.A(new_n3855_), .B(new_n4023_), .Y(new_n4024_));
  NOR2X1   g03768(.A(new_n3864_), .B(new_n4024_), .Y(new_n4025_));
  AOI21X1  g03769(.A0(new_n3867_), .A1(new_n3866_), .B0(new_n3865_), .Y(new_n4026_));
  OR2X1    g03770(.A(new_n4026_), .B(new_n4025_), .Y(new_n4027_));
  XOR2X1   g03771(.A(new_n4027_), .B(new_n4020_), .Y(\f[43] ));
  NAND2X1  g03772(.A(new_n4019_), .B(new_n4009_), .Y(new_n4029_));
  OAI21X1  g03773(.A0(new_n4026_), .A1(new_n4025_), .B0(new_n4020_), .Y(new_n4030_));
  AND2X1   g03774(.A(new_n4030_), .B(new_n4029_), .Y(new_n4031_));
  AND2X1   g03775(.A(new_n4007_), .B(new_n4003_), .Y(new_n4032_));
  AOI21X1  g03776(.A0(new_n4008_), .A1(new_n3872_), .B0(new_n4032_), .Y(new_n4033_));
  AOI22X1  g03777(.A0(new_n369_), .A1(\b[41] ), .B0(new_n368_), .B1(\b[40] ), .Y(new_n4034_));
  OAI21X1  g03778(.A0(new_n367_), .A1(new_n3723_), .B0(new_n4034_), .Y(new_n4035_));
  AOI21X1  g03779(.A0(new_n3722_), .A1(new_n308_), .B0(new_n4035_), .Y(new_n4036_));
  XOR2X1   g03780(.A(new_n4036_), .B(\a[5] ), .Y(new_n4037_));
  NOR2X1   g03781(.A(new_n3562_), .B(new_n3452_), .Y(new_n4038_));
  NAND2X1  g03782(.A(new_n3562_), .B(new_n3452_), .Y(new_n4039_));
  OAI21X1  g03783(.A0(new_n4038_), .A1(new_n3591_), .B0(new_n4039_), .Y(new_n4040_));
  NOR2X1   g03784(.A(new_n3709_), .B(new_n3705_), .Y(new_n4041_));
  AOI21X1  g03785(.A0(new_n3710_), .A1(new_n4040_), .B0(new_n4041_), .Y(new_n4042_));
  AND2X1   g03786(.A(new_n3852_), .B(new_n3848_), .Y(new_n4043_));
  OR2X1    g03787(.A(new_n3852_), .B(new_n3848_), .Y(new_n4044_));
  OAI21X1  g03788(.A0(new_n4043_), .A1(new_n4042_), .B0(new_n4044_), .Y(new_n4045_));
  NOR2X1   g03789(.A(new_n3998_), .B(new_n3994_), .Y(new_n4046_));
  AOI21X1  g03790(.A0(new_n4000_), .A1(new_n4045_), .B0(new_n4046_), .Y(new_n4047_));
  AND2X1   g03791(.A(new_n3981_), .B(new_n3977_), .Y(new_n4048_));
  OR2X1    g03792(.A(new_n3981_), .B(new_n3977_), .Y(new_n4049_));
  OAI21X1  g03793(.A0(new_n4048_), .A1(new_n3876_), .B0(new_n4049_), .Y(new_n4050_));
  AOI22X1  g03794(.A0(new_n818_), .A1(\b[32] ), .B0(new_n817_), .B1(\b[31] ), .Y(new_n4051_));
  OAI21X1  g03795(.A0(new_n816_), .A1(new_n2356_), .B0(new_n4051_), .Y(new_n4052_));
  AOI21X1  g03796(.A0(new_n2495_), .A1(new_n668_), .B0(new_n4052_), .Y(new_n4053_));
  XOR2X1   g03797(.A(new_n4053_), .B(new_n665_), .Y(new_n4054_));
  INVX1    g03798(.A(new_n3882_), .Y(new_n4055_));
  AND2X1   g03799(.A(new_n3975_), .B(new_n4055_), .Y(new_n4056_));
  XOR2X1   g03800(.A(new_n3975_), .B(new_n4055_), .Y(new_n4057_));
  AOI21X1  g03801(.A0(new_n4057_), .A1(new_n3878_), .B0(new_n4056_), .Y(new_n4058_));
  AOI22X1  g03802(.A0(new_n1017_), .A1(\b[29] ), .B0(new_n1016_), .B1(\b[28] ), .Y(new_n4059_));
  OAI21X1  g03803(.A0(new_n1015_), .A1(new_n2126_), .B0(new_n4059_), .Y(new_n4060_));
  AOI21X1  g03804(.A0(new_n2125_), .A1(new_n882_), .B0(new_n4060_), .Y(new_n4061_));
  XOR2X1   g03805(.A(new_n4061_), .B(\a[17] ), .Y(new_n4062_));
  XOR2X1   g03806(.A(new_n3964_), .B(new_n3960_), .Y(new_n4063_));
  OR2X1    g03807(.A(new_n3969_), .B(new_n4063_), .Y(new_n4064_));
  OAI21X1  g03808(.A0(new_n3974_), .A1(new_n3970_), .B0(new_n4064_), .Y(new_n4065_));
  NOR2X1   g03809(.A(new_n3885_), .B(new_n3884_), .Y(new_n4066_));
  XOR2X1   g03810(.A(new_n3935_), .B(new_n4066_), .Y(new_n4067_));
  OR2X1    g03811(.A(new_n3940_), .B(new_n4067_), .Y(new_n4068_));
  OAI21X1  g03812(.A0(new_n3945_), .A1(new_n3941_), .B0(new_n4068_), .Y(new_n4069_));
  AOI22X1  g03813(.A0(new_n2163_), .A1(\b[17] ), .B0(new_n2162_), .B1(\b[16] ), .Y(new_n4070_));
  OAI21X1  g03814(.A0(new_n2161_), .A1(new_n977_), .B0(new_n4070_), .Y(new_n4071_));
  AOI21X1  g03815(.A0(new_n1907_), .A1(new_n976_), .B0(new_n4071_), .Y(new_n4072_));
  XOR2X1   g03816(.A(new_n4072_), .B(\a[29] ), .Y(new_n4073_));
  INVX1    g03817(.A(new_n4073_), .Y(new_n4074_));
  NOR2X1   g03818(.A(new_n3934_), .B(new_n3930_), .Y(new_n4075_));
  AOI21X1  g03819(.A0(new_n3935_), .A1(new_n3886_), .B0(new_n4075_), .Y(new_n4076_));
  AOI22X1  g03820(.A0(new_n2545_), .A1(\b[14] ), .B0(new_n2544_), .B1(\b[13] ), .Y(new_n4077_));
  OAI21X1  g03821(.A0(new_n2543_), .A1(new_n713_), .B0(new_n4077_), .Y(new_n4078_));
  AOI21X1  g03822(.A0(new_n2260_), .A1(new_n734_), .B0(new_n4078_), .Y(new_n4079_));
  XOR2X1   g03823(.A(new_n4079_), .B(\a[32] ), .Y(new_n4080_));
  INVX1    g03824(.A(new_n4080_), .Y(new_n4081_));
  INVX1    g03825(.A(new_n3910_), .Y(new_n4082_));
  OR2X1    g03826(.A(new_n3919_), .B(new_n3915_), .Y(new_n4083_));
  OAI21X1  g03827(.A0(new_n3914_), .A1(new_n4082_), .B0(new_n4083_), .Y(new_n4084_));
  AOI22X1  g03828(.A0(new_n3204_), .A1(\b[8] ), .B0(new_n3203_), .B1(\b[7] ), .Y(new_n4085_));
  OAI21X1  g03829(.A0(new_n3321_), .A1(new_n392_), .B0(new_n4085_), .Y(new_n4086_));
  AOI21X1  g03830(.A0(new_n3080_), .A1(new_n454_), .B0(new_n4086_), .Y(new_n4087_));
  XOR2X1   g03831(.A(new_n4087_), .B(\a[38] ), .Y(new_n4088_));
  AND2X1   g03832(.A(new_n3908_), .B(new_n3896_), .Y(new_n4089_));
  AOI21X1  g03833(.A0(new_n3909_), .A1(new_n3891_), .B0(new_n4089_), .Y(new_n4090_));
  NAND3X1  g03834(.A(new_n3906_), .B(new_n3774_), .C(\a[44] ), .Y(new_n4091_));
  NAND2X1  g03835(.A(new_n3901_), .B(new_n341_), .Y(new_n4092_));
  OR4X1    g03836(.A(new_n3902_), .B(new_n3900_), .C(new_n3773_), .D(new_n274_), .Y(new_n4093_));
  AND2X1   g03837(.A(new_n3902_), .B(new_n3898_), .Y(new_n4094_));
  AND2X1   g03838(.A(new_n3900_), .B(new_n3773_), .Y(new_n4095_));
  AOI22X1  g03839(.A0(new_n4095_), .A1(\b[2] ), .B0(new_n4094_), .B1(\b[1] ), .Y(new_n4096_));
  NAND3X1  g03840(.A(new_n4096_), .B(new_n4093_), .C(new_n4092_), .Y(new_n4097_));
  XOR2X1   g03841(.A(new_n4097_), .B(new_n3899_), .Y(new_n4098_));
  XOR2X1   g03842(.A(new_n4098_), .B(new_n4091_), .Y(new_n4099_));
  AOI22X1  g03843(.A0(new_n3652_), .A1(\b[5] ), .B0(new_n3651_), .B1(\b[4] ), .Y(new_n4100_));
  OAI21X1  g03844(.A0(new_n3778_), .A1(new_n297_), .B0(new_n4100_), .Y(new_n4101_));
  AOI21X1  g03845(.A0(new_n3480_), .A1(new_n349_), .B0(new_n4101_), .Y(new_n4102_));
  XOR2X1   g03846(.A(new_n4102_), .B(\a[41] ), .Y(new_n4103_));
  XOR2X1   g03847(.A(new_n4103_), .B(new_n4099_), .Y(new_n4104_));
  XOR2X1   g03848(.A(new_n4104_), .B(new_n4090_), .Y(new_n4105_));
  XOR2X1   g03849(.A(new_n4105_), .B(new_n4088_), .Y(new_n4106_));
  INVX1    g03850(.A(new_n4106_), .Y(new_n4107_));
  XOR2X1   g03851(.A(new_n4107_), .B(new_n4084_), .Y(new_n4108_));
  AOI22X1  g03852(.A0(new_n2813_), .A1(\b[11] ), .B0(new_n2812_), .B1(\b[10] ), .Y(new_n4109_));
  OAI21X1  g03853(.A0(new_n2946_), .A1(new_n590_), .B0(new_n4109_), .Y(new_n4110_));
  AOI21X1  g03854(.A0(new_n2652_), .A1(new_n589_), .B0(new_n4110_), .Y(new_n4111_));
  XOR2X1   g03855(.A(new_n4111_), .B(\a[35] ), .Y(new_n4112_));
  XOR2X1   g03856(.A(new_n4112_), .B(new_n4108_), .Y(new_n4113_));
  XOR2X1   g03857(.A(new_n4113_), .B(new_n3929_), .Y(new_n4114_));
  XOR2X1   g03858(.A(new_n4114_), .B(new_n4081_), .Y(new_n4115_));
  INVX1    g03859(.A(new_n4115_), .Y(new_n4116_));
  XOR2X1   g03860(.A(new_n4116_), .B(new_n4076_), .Y(new_n4117_));
  XOR2X1   g03861(.A(new_n4117_), .B(new_n4074_), .Y(new_n4118_));
  XOR2X1   g03862(.A(new_n4118_), .B(new_n4069_), .Y(new_n4119_));
  AOI22X1  g03863(.A0(new_n1814_), .A1(\b[20] ), .B0(new_n1813_), .B1(\b[19] ), .Y(new_n4120_));
  OAI21X1  g03864(.A0(new_n1812_), .A1(new_n1115_), .B0(new_n4120_), .Y(new_n4121_));
  AOI21X1  g03865(.A0(new_n1617_), .A1(new_n1217_), .B0(new_n4121_), .Y(new_n4122_));
  XOR2X1   g03866(.A(new_n4122_), .B(\a[26] ), .Y(new_n4123_));
  XOR2X1   g03867(.A(new_n4123_), .B(new_n4119_), .Y(new_n4124_));
  INVX1    g03868(.A(new_n4124_), .Y(new_n4125_));
  XOR2X1   g03869(.A(new_n3940_), .B(new_n4067_), .Y(new_n4126_));
  XOR2X1   g03870(.A(new_n3945_), .B(new_n4126_), .Y(new_n4127_));
  NOR2X1   g03871(.A(new_n3950_), .B(new_n4127_), .Y(new_n4128_));
  XOR2X1   g03872(.A(new_n3950_), .B(new_n4127_), .Y(new_n4129_));
  AOI21X1  g03873(.A0(new_n3954_), .A1(new_n4129_), .B0(new_n4128_), .Y(new_n4130_));
  XOR2X1   g03874(.A(new_n4130_), .B(new_n4125_), .Y(new_n4131_));
  AOI22X1  g03875(.A0(new_n1526_), .A1(\b[23] ), .B0(new_n1525_), .B1(\b[22] ), .Y(new_n4132_));
  OAI21X1  g03876(.A0(new_n1524_), .A1(new_n1482_), .B0(new_n4132_), .Y(new_n4133_));
  AOI21X1  g03877(.A0(new_n1481_), .A1(new_n1347_), .B0(new_n4133_), .Y(new_n4134_));
  XOR2X1   g03878(.A(new_n4134_), .B(\a[23] ), .Y(new_n4135_));
  NAND2X1  g03879(.A(new_n4135_), .B(new_n4131_), .Y(new_n4136_));
  OR2X1    g03880(.A(new_n3959_), .B(new_n3955_), .Y(new_n4137_));
  OAI21X1  g03881(.A0(new_n3963_), .A1(new_n3962_), .B0(new_n3960_), .Y(new_n4138_));
  OR2X1    g03882(.A(new_n4135_), .B(new_n4131_), .Y(new_n4139_));
  AOI22X1  g03883(.A0(new_n4136_), .A1(new_n4139_), .B0(new_n4138_), .B1(new_n4137_), .Y(new_n4140_));
  NAND2X1  g03884(.A(new_n4138_), .B(new_n4137_), .Y(new_n4141_));
  NOR2X1   g03885(.A(new_n4135_), .B(new_n4131_), .Y(new_n4142_));
  AOI21X1  g03886(.A0(new_n4136_), .A1(new_n4141_), .B0(new_n4142_), .Y(new_n4143_));
  AOI21X1  g03887(.A0(new_n4143_), .A1(new_n4136_), .B0(new_n4140_), .Y(new_n4144_));
  AOI22X1  g03888(.A0(new_n1263_), .A1(\b[26] ), .B0(new_n1262_), .B1(\b[25] ), .Y(new_n4145_));
  OAI21X1  g03889(.A0(new_n1261_), .A1(new_n1588_), .B0(new_n4145_), .Y(new_n4146_));
  AOI21X1  g03890(.A0(new_n1783_), .A1(new_n1075_), .B0(new_n4146_), .Y(new_n4147_));
  XOR2X1   g03891(.A(new_n4147_), .B(\a[20] ), .Y(new_n4148_));
  XOR2X1   g03892(.A(new_n4148_), .B(new_n4144_), .Y(new_n4149_));
  XOR2X1   g03893(.A(new_n4149_), .B(new_n4065_), .Y(new_n4150_));
  XOR2X1   g03894(.A(new_n4150_), .B(new_n4062_), .Y(new_n4151_));
  XOR2X1   g03895(.A(new_n4151_), .B(new_n4058_), .Y(new_n4152_));
  XOR2X1   g03896(.A(new_n4152_), .B(new_n4054_), .Y(new_n4153_));
  XOR2X1   g03897(.A(new_n4153_), .B(new_n4050_), .Y(new_n4154_));
  AOI22X1  g03898(.A0(new_n603_), .A1(\b[35] ), .B0(new_n602_), .B1(\b[34] ), .Y(new_n4155_));
  OAI21X1  g03899(.A0(new_n601_), .A1(new_n2893_), .B0(new_n4155_), .Y(new_n4156_));
  AOI21X1  g03900(.A0(new_n2892_), .A1(new_n518_), .B0(new_n4156_), .Y(new_n4157_));
  XOR2X1   g03901(.A(new_n4157_), .B(\a[11] ), .Y(new_n4158_));
  XOR2X1   g03902(.A(new_n4158_), .B(new_n4154_), .Y(new_n4159_));
  NOR2X1   g03903(.A(new_n3987_), .B(new_n3983_), .Y(new_n4160_));
  AND2X1   g03904(.A(new_n3703_), .B(new_n3603_), .Y(new_n4161_));
  AOI21X1  g03905(.A0(new_n3704_), .A1(new_n3743_), .B0(new_n4161_), .Y(new_n4162_));
  OR2X1    g03906(.A(new_n3846_), .B(new_n3990_), .Y(new_n4163_));
  OAI21X1  g03907(.A0(new_n3847_), .A1(new_n4162_), .B0(new_n4163_), .Y(new_n4164_));
  AOI21X1  g03908(.A0(new_n4164_), .A1(new_n3988_), .B0(new_n4160_), .Y(new_n4165_));
  XOR2X1   g03909(.A(new_n4165_), .B(new_n4159_), .Y(new_n4166_));
  AOI22X1  g03910(.A0(new_n469_), .A1(\b[38] ), .B0(new_n468_), .B1(\b[37] ), .Y(new_n4167_));
  OAI21X1  g03911(.A0(new_n467_), .A1(new_n3276_), .B0(new_n4167_), .Y(new_n4168_));
  AOI21X1  g03912(.A0(new_n3275_), .A1(new_n404_), .B0(new_n4168_), .Y(new_n4169_));
  XOR2X1   g03913(.A(new_n4169_), .B(\a[8] ), .Y(new_n4170_));
  XOR2X1   g03914(.A(new_n4170_), .B(new_n4166_), .Y(new_n4171_));
  XOR2X1   g03915(.A(new_n4171_), .B(new_n4047_), .Y(new_n4172_));
  XOR2X1   g03916(.A(new_n4172_), .B(new_n4037_), .Y(new_n4173_));
  XOR2X1   g03917(.A(new_n4173_), .B(new_n4033_), .Y(new_n4174_));
  NAND2X1  g03918(.A(\b[43] ), .B(\b[42] ), .Y(new_n4175_));
  OAI21X1  g03919(.A0(new_n4013_), .A1(new_n4011_), .B0(new_n4175_), .Y(new_n4176_));
  XOR2X1   g03920(.A(\b[44] ), .B(\b[43] ), .Y(new_n4177_));
  XOR2X1   g03921(.A(new_n4177_), .B(new_n4176_), .Y(new_n4178_));
  AOI22X1  g03922(.A0(new_n267_), .A1(\b[44] ), .B0(new_n266_), .B1(\b[43] ), .Y(new_n4179_));
  OAI21X1  g03923(.A0(new_n350_), .A1(new_n4012_), .B0(new_n4179_), .Y(new_n4180_));
  AOI21X1  g03924(.A0(new_n4178_), .A1(new_n318_), .B0(new_n4180_), .Y(new_n4181_));
  XOR2X1   g03925(.A(new_n4181_), .B(\a[2] ), .Y(new_n4182_));
  XOR2X1   g03926(.A(new_n4182_), .B(new_n4174_), .Y(new_n4183_));
  XOR2X1   g03927(.A(new_n4183_), .B(new_n4031_), .Y(\f[44] ));
  AOI21X1  g03928(.A0(new_n4030_), .A1(new_n4029_), .B0(new_n4183_), .Y(new_n4185_));
  INVX1    g03929(.A(new_n4037_), .Y(new_n4186_));
  XOR2X1   g03930(.A(new_n4172_), .B(new_n4186_), .Y(new_n4187_));
  XOR2X1   g03931(.A(new_n4187_), .B(new_n4033_), .Y(new_n4188_));
  NOR2X1   g03932(.A(new_n4182_), .B(new_n4188_), .Y(new_n4189_));
  OR2X1    g03933(.A(new_n4189_), .B(new_n4185_), .Y(new_n4190_));
  OR2X1    g03934(.A(new_n3840_), .B(new_n3836_), .Y(new_n4191_));
  AND2X1   g03935(.A(new_n3840_), .B(new_n3836_), .Y(new_n4192_));
  OAI21X1  g03936(.A0(new_n4192_), .A1(new_n3989_), .B0(new_n4191_), .Y(new_n4193_));
  NOR2X1   g03937(.A(new_n3981_), .B(new_n3977_), .Y(new_n4194_));
  AOI21X1  g03938(.A0(new_n3982_), .A1(new_n4193_), .B0(new_n4194_), .Y(new_n4195_));
  XOR2X1   g03939(.A(new_n4153_), .B(new_n4195_), .Y(new_n4196_));
  NOR2X1   g03940(.A(new_n4158_), .B(new_n4196_), .Y(new_n4197_));
  XOR2X1   g03941(.A(new_n4158_), .B(new_n4196_), .Y(new_n4198_));
  OR2X1    g03942(.A(new_n3987_), .B(new_n3983_), .Y(new_n4199_));
  XOR2X1   g03943(.A(new_n3982_), .B(new_n4193_), .Y(new_n4200_));
  XOR2X1   g03944(.A(new_n3987_), .B(new_n4200_), .Y(new_n4201_));
  OAI21X1  g03945(.A0(new_n3993_), .A1(new_n4201_), .B0(new_n4199_), .Y(new_n4202_));
  AOI21X1  g03946(.A0(new_n4202_), .A1(new_n4198_), .B0(new_n4197_), .Y(new_n4203_));
  NOR2X1   g03947(.A(new_n4152_), .B(new_n4054_), .Y(new_n4204_));
  NAND2X1  g03948(.A(new_n4152_), .B(new_n4054_), .Y(new_n4205_));
  OAI21X1  g03949(.A0(new_n4204_), .A1(new_n4195_), .B0(new_n4205_), .Y(new_n4206_));
  INVX1    g03950(.A(new_n4062_), .Y(new_n4207_));
  NAND2X1  g03951(.A(new_n4150_), .B(new_n4207_), .Y(new_n4208_));
  OAI21X1  g03952(.A0(new_n4151_), .A1(new_n4058_), .B0(new_n4208_), .Y(new_n4209_));
  NOR2X1   g03953(.A(new_n4148_), .B(new_n4144_), .Y(new_n4210_));
  AOI21X1  g03954(.A0(new_n4149_), .A1(new_n4065_), .B0(new_n4210_), .Y(new_n4211_));
  AND2X1   g03955(.A(new_n4117_), .B(new_n4074_), .Y(new_n4212_));
  AOI21X1  g03956(.A0(new_n4118_), .A1(new_n4069_), .B0(new_n4212_), .Y(new_n4213_));
  AND2X1   g03957(.A(new_n4114_), .B(new_n4081_), .Y(new_n4214_));
  INVX1    g03958(.A(new_n4214_), .Y(new_n4215_));
  OAI21X1  g03959(.A0(new_n4116_), .A1(new_n4076_), .B0(new_n4215_), .Y(new_n4216_));
  XOR2X1   g03960(.A(new_n4106_), .B(new_n4084_), .Y(new_n4217_));
  OR2X1    g03961(.A(new_n4112_), .B(new_n4217_), .Y(new_n4218_));
  OAI21X1  g03962(.A0(new_n4113_), .A1(new_n3929_), .B0(new_n4218_), .Y(new_n4219_));
  AOI22X1  g03963(.A0(new_n2813_), .A1(\b[12] ), .B0(new_n2812_), .B1(\b[11] ), .Y(new_n4220_));
  OAI21X1  g03964(.A0(new_n2946_), .A1(new_n587_), .B0(new_n4220_), .Y(new_n4221_));
  AOI21X1  g03965(.A0(new_n2652_), .A1(new_n635_), .B0(new_n4221_), .Y(new_n4222_));
  XOR2X1   g03966(.A(new_n4222_), .B(\a[35] ), .Y(new_n4223_));
  INVX1    g03967(.A(new_n4088_), .Y(new_n4224_));
  AND2X1   g03968(.A(new_n4105_), .B(new_n4224_), .Y(new_n4225_));
  AOI21X1  g03969(.A0(new_n4107_), .A1(new_n4084_), .B0(new_n4225_), .Y(new_n4226_));
  OR2X1    g03970(.A(new_n4098_), .B(new_n4091_), .Y(new_n4227_));
  XOR2X1   g03971(.A(\a[45] ), .B(\a[44] ), .Y(new_n4228_));
  NAND2X1  g03972(.A(new_n4228_), .B(\b[0] ), .Y(new_n4229_));
  INVX1    g03973(.A(new_n4229_), .Y(new_n4230_));
  XOR2X1   g03974(.A(new_n4230_), .B(new_n4227_), .Y(new_n4231_));
  OR2X1    g03975(.A(new_n3902_), .B(new_n3773_), .Y(new_n4232_));
  OR2X1    g03976(.A(new_n4232_), .B(new_n3900_), .Y(new_n4233_));
  AOI22X1  g03977(.A0(new_n4095_), .A1(\b[3] ), .B0(new_n4094_), .B1(\b[2] ), .Y(new_n4234_));
  OAI21X1  g03978(.A0(new_n4233_), .A1(new_n275_), .B0(new_n4234_), .Y(new_n4235_));
  AOI21X1  g03979(.A0(new_n3901_), .A1(new_n366_), .B0(new_n4235_), .Y(new_n4236_));
  XOR2X1   g03980(.A(new_n4236_), .B(\a[44] ), .Y(new_n4237_));
  XOR2X1   g03981(.A(new_n4237_), .B(new_n4231_), .Y(new_n4238_));
  AOI22X1  g03982(.A0(new_n3652_), .A1(\b[6] ), .B0(new_n3651_), .B1(\b[5] ), .Y(new_n4239_));
  OAI21X1  g03983(.A0(new_n3778_), .A1(new_n325_), .B0(new_n4239_), .Y(new_n4240_));
  AOI21X1  g03984(.A0(new_n3480_), .A1(new_n378_), .B0(new_n4240_), .Y(new_n4241_));
  XOR2X1   g03985(.A(new_n4241_), .B(\a[41] ), .Y(new_n4242_));
  XOR2X1   g03986(.A(new_n4242_), .B(new_n4238_), .Y(new_n4243_));
  INVX1    g03987(.A(new_n4103_), .Y(new_n4244_));
  NOR2X1   g03988(.A(new_n4104_), .B(new_n4090_), .Y(new_n4245_));
  AOI21X1  g03989(.A0(new_n4244_), .A1(new_n4099_), .B0(new_n4245_), .Y(new_n4246_));
  XOR2X1   g03990(.A(new_n4246_), .B(new_n4243_), .Y(new_n4247_));
  AOI22X1  g03991(.A0(new_n3204_), .A1(\b[9] ), .B0(new_n3203_), .B1(\b[8] ), .Y(new_n4248_));
  OAI21X1  g03992(.A0(new_n3321_), .A1(new_n492_), .B0(new_n4248_), .Y(new_n4249_));
  AOI21X1  g03993(.A0(new_n3080_), .A1(new_n491_), .B0(new_n4249_), .Y(new_n4250_));
  XOR2X1   g03994(.A(new_n4250_), .B(\a[38] ), .Y(new_n4251_));
  XOR2X1   g03995(.A(new_n4251_), .B(new_n4247_), .Y(new_n4252_));
  XOR2X1   g03996(.A(new_n4252_), .B(new_n4226_), .Y(new_n4253_));
  XOR2X1   g03997(.A(new_n4253_), .B(new_n4223_), .Y(new_n4254_));
  XOR2X1   g03998(.A(new_n4254_), .B(new_n4219_), .Y(new_n4255_));
  AOI22X1  g03999(.A0(new_n2545_), .A1(\b[15] ), .B0(new_n2544_), .B1(\b[14] ), .Y(new_n4256_));
  OAI21X1  g04000(.A0(new_n2543_), .A1(new_n795_), .B0(new_n4256_), .Y(new_n4257_));
  AOI21X1  g04001(.A0(new_n2260_), .A1(new_n794_), .B0(new_n4257_), .Y(new_n4258_));
  XOR2X1   g04002(.A(new_n4258_), .B(\a[32] ), .Y(new_n4259_));
  XOR2X1   g04003(.A(new_n4259_), .B(new_n4255_), .Y(new_n4260_));
  INVX1    g04004(.A(new_n4260_), .Y(new_n4261_));
  XOR2X1   g04005(.A(new_n4261_), .B(new_n4216_), .Y(new_n4262_));
  AOI22X1  g04006(.A0(new_n2163_), .A1(\b[18] ), .B0(new_n2162_), .B1(\b[17] ), .Y(new_n4263_));
  OAI21X1  g04007(.A0(new_n2161_), .A1(new_n974_), .B0(new_n4263_), .Y(new_n4264_));
  AOI21X1  g04008(.A0(new_n1907_), .A1(new_n1042_), .B0(new_n4264_), .Y(new_n4265_));
  XOR2X1   g04009(.A(new_n4265_), .B(\a[29] ), .Y(new_n4266_));
  XOR2X1   g04010(.A(new_n4266_), .B(new_n4262_), .Y(new_n4267_));
  XOR2X1   g04011(.A(new_n4267_), .B(new_n4213_), .Y(new_n4268_));
  AOI22X1  g04012(.A0(new_n1814_), .A1(\b[21] ), .B0(new_n1813_), .B1(\b[20] ), .Y(new_n4269_));
  OAI21X1  g04013(.A0(new_n1812_), .A1(new_n1300_), .B0(new_n4269_), .Y(new_n4270_));
  AOI21X1  g04014(.A0(new_n1617_), .A1(new_n1299_), .B0(new_n4270_), .Y(new_n4271_));
  XOR2X1   g04015(.A(new_n4271_), .B(\a[26] ), .Y(new_n4272_));
  XOR2X1   g04016(.A(new_n4272_), .B(new_n4268_), .Y(new_n4273_));
  INVX1    g04017(.A(new_n4273_), .Y(new_n4274_));
  XOR2X1   g04018(.A(new_n4117_), .B(new_n4073_), .Y(new_n4275_));
  XOR2X1   g04019(.A(new_n4275_), .B(new_n4069_), .Y(new_n4276_));
  OR2X1    g04020(.A(new_n4123_), .B(new_n4276_), .Y(new_n4277_));
  OAI21X1  g04021(.A0(new_n4130_), .A1(new_n4124_), .B0(new_n4277_), .Y(new_n4278_));
  XOR2X1   g04022(.A(new_n4278_), .B(new_n4274_), .Y(new_n4279_));
  AOI22X1  g04023(.A0(new_n1526_), .A1(\b[24] ), .B0(new_n1525_), .B1(\b[23] ), .Y(new_n4280_));
  OAI21X1  g04024(.A0(new_n1524_), .A1(new_n1479_), .B0(new_n4280_), .Y(new_n4281_));
  AOI21X1  g04025(.A0(new_n1572_), .A1(new_n1347_), .B0(new_n4281_), .Y(new_n4282_));
  XOR2X1   g04026(.A(new_n4282_), .B(\a[23] ), .Y(new_n4283_));
  XOR2X1   g04027(.A(new_n4283_), .B(new_n4279_), .Y(new_n4284_));
  XOR2X1   g04028(.A(new_n4284_), .B(new_n4143_), .Y(new_n4285_));
  AOI22X1  g04029(.A0(new_n1263_), .A1(\b[27] ), .B0(new_n1262_), .B1(\b[26] ), .Y(new_n4286_));
  OAI21X1  g04030(.A0(new_n1261_), .A1(new_n1880_), .B0(new_n4286_), .Y(new_n4287_));
  AOI21X1  g04031(.A0(new_n1879_), .A1(new_n1075_), .B0(new_n4287_), .Y(new_n4288_));
  XOR2X1   g04032(.A(new_n4288_), .B(\a[20] ), .Y(new_n4289_));
  XOR2X1   g04033(.A(new_n4289_), .B(new_n4285_), .Y(new_n4290_));
  XOR2X1   g04034(.A(new_n4290_), .B(new_n4211_), .Y(new_n4291_));
  AOI22X1  g04035(.A0(new_n1017_), .A1(\b[30] ), .B0(new_n1016_), .B1(\b[29] ), .Y(new_n4292_));
  OAI21X1  g04036(.A0(new_n1015_), .A1(new_n2231_), .B0(new_n4292_), .Y(new_n4293_));
  AOI21X1  g04037(.A0(new_n2230_), .A1(new_n882_), .B0(new_n4293_), .Y(new_n4294_));
  XOR2X1   g04038(.A(new_n4294_), .B(\a[17] ), .Y(new_n4295_));
  XOR2X1   g04039(.A(new_n4295_), .B(new_n4291_), .Y(new_n4296_));
  XOR2X1   g04040(.A(new_n4296_), .B(new_n4209_), .Y(new_n4297_));
  AOI22X1  g04041(.A0(new_n818_), .A1(\b[33] ), .B0(new_n817_), .B1(\b[32] ), .Y(new_n4298_));
  OAI21X1  g04042(.A0(new_n816_), .A1(new_n2615_), .B0(new_n4298_), .Y(new_n4299_));
  AOI21X1  g04043(.A0(new_n2614_), .A1(new_n668_), .B0(new_n4299_), .Y(new_n4300_));
  XOR2X1   g04044(.A(new_n4300_), .B(\a[14] ), .Y(new_n4301_));
  XOR2X1   g04045(.A(new_n4301_), .B(new_n4297_), .Y(new_n4302_));
  XOR2X1   g04046(.A(new_n4302_), .B(new_n4206_), .Y(new_n4303_));
  AOI22X1  g04047(.A0(new_n603_), .A1(\b[36] ), .B0(new_n602_), .B1(\b[35] ), .Y(new_n4304_));
  OAI21X1  g04048(.A0(new_n601_), .A1(new_n2890_), .B0(new_n4304_), .Y(new_n4305_));
  AOI21X1  g04049(.A0(new_n3015_), .A1(new_n518_), .B0(new_n4305_), .Y(new_n4306_));
  XOR2X1   g04050(.A(new_n4306_), .B(\a[11] ), .Y(new_n4307_));
  XOR2X1   g04051(.A(new_n4307_), .B(new_n4303_), .Y(new_n4308_));
  XOR2X1   g04052(.A(new_n4308_), .B(new_n4203_), .Y(new_n4309_));
  AOI22X1  g04053(.A0(new_n469_), .A1(\b[39] ), .B0(new_n468_), .B1(\b[38] ), .Y(new_n4310_));
  OAI21X1  g04054(.A0(new_n467_), .A1(new_n3413_), .B0(new_n4310_), .Y(new_n4311_));
  AOI21X1  g04055(.A0(new_n3412_), .A1(new_n404_), .B0(new_n4311_), .Y(new_n4312_));
  XOR2X1   g04056(.A(new_n4312_), .B(\a[8] ), .Y(new_n4313_));
  XOR2X1   g04057(.A(new_n4313_), .B(new_n4309_), .Y(new_n4314_));
  XOR2X1   g04058(.A(new_n4165_), .B(new_n4198_), .Y(new_n4315_));
  NOR2X1   g04059(.A(new_n4170_), .B(new_n4315_), .Y(new_n4316_));
  XOR2X1   g04060(.A(new_n4170_), .B(new_n4315_), .Y(new_n4317_));
  AOI21X1  g04061(.A0(new_n4317_), .A1(new_n4002_), .B0(new_n4316_), .Y(new_n4318_));
  XOR2X1   g04062(.A(new_n4318_), .B(new_n4314_), .Y(new_n4319_));
  AOI22X1  g04063(.A0(new_n369_), .A1(\b[42] ), .B0(new_n368_), .B1(\b[41] ), .Y(new_n4320_));
  OAI21X1  g04064(.A0(new_n367_), .A1(new_n3720_), .B0(new_n4320_), .Y(new_n4321_));
  AOI21X1  g04065(.A0(new_n3860_), .A1(new_n308_), .B0(new_n4321_), .Y(new_n4322_));
  XOR2X1   g04066(.A(new_n4322_), .B(\a[5] ), .Y(new_n4323_));
  XOR2X1   g04067(.A(new_n4323_), .B(new_n4319_), .Y(new_n4324_));
  AND2X1   g04068(.A(new_n3854_), .B(new_n3870_), .Y(new_n4325_));
  XOR2X1   g04069(.A(new_n3854_), .B(new_n3870_), .Y(new_n4326_));
  AOI21X1  g04070(.A0(new_n4326_), .A1(new_n4023_), .B0(new_n4325_), .Y(new_n4327_));
  NOR2X1   g04071(.A(new_n4007_), .B(new_n4003_), .Y(new_n4328_));
  NAND2X1  g04072(.A(new_n4007_), .B(new_n4003_), .Y(new_n4329_));
  OAI21X1  g04073(.A0(new_n4328_), .A1(new_n4327_), .B0(new_n4329_), .Y(new_n4330_));
  AND2X1   g04074(.A(new_n4172_), .B(new_n4186_), .Y(new_n4331_));
  AOI21X1  g04075(.A0(new_n4187_), .A1(new_n4330_), .B0(new_n4331_), .Y(new_n4332_));
  XOR2X1   g04076(.A(new_n4332_), .B(new_n4324_), .Y(new_n4333_));
  AND2X1   g04077(.A(\b[44] ), .B(\b[43] ), .Y(new_n4334_));
  AOI21X1  g04078(.A0(new_n4177_), .A1(new_n4176_), .B0(new_n4334_), .Y(new_n4335_));
  INVX1    g04079(.A(\b[44] ), .Y(new_n4336_));
  XOR2X1   g04080(.A(\b[45] ), .B(new_n4336_), .Y(new_n4337_));
  XOR2X1   g04081(.A(new_n4337_), .B(new_n4335_), .Y(new_n4338_));
  INVX1    g04082(.A(\b[43] ), .Y(new_n4339_));
  AOI22X1  g04083(.A0(new_n267_), .A1(\b[45] ), .B0(new_n266_), .B1(\b[44] ), .Y(new_n4340_));
  OAI21X1  g04084(.A0(new_n350_), .A1(new_n4339_), .B0(new_n4340_), .Y(new_n4341_));
  AOI21X1  g04085(.A0(new_n4338_), .A1(new_n318_), .B0(new_n4341_), .Y(new_n4342_));
  XOR2X1   g04086(.A(new_n4342_), .B(\a[2] ), .Y(new_n4343_));
  XOR2X1   g04087(.A(new_n4343_), .B(new_n4333_), .Y(new_n4344_));
  XOR2X1   g04088(.A(new_n4344_), .B(new_n4190_), .Y(\f[45] ));
  NOR2X1   g04089(.A(new_n4295_), .B(new_n4291_), .Y(new_n4346_));
  AOI21X1  g04090(.A0(new_n4296_), .A1(new_n4209_), .B0(new_n4346_), .Y(new_n4347_));
  OR2X1    g04091(.A(new_n4289_), .B(new_n4285_), .Y(new_n4348_));
  AND2X1   g04092(.A(new_n4138_), .B(new_n4137_), .Y(new_n4349_));
  AND2X1   g04093(.A(new_n4135_), .B(new_n4131_), .Y(new_n4350_));
  OAI21X1  g04094(.A0(new_n4350_), .A1(new_n4349_), .B0(new_n4139_), .Y(new_n4351_));
  XOR2X1   g04095(.A(new_n4284_), .B(new_n4351_), .Y(new_n4352_));
  XOR2X1   g04096(.A(new_n4289_), .B(new_n4352_), .Y(new_n4353_));
  OAI21X1  g04097(.A0(new_n4353_), .A1(new_n4211_), .B0(new_n4348_), .Y(new_n4354_));
  AOI22X1  g04098(.A0(new_n1263_), .A1(\b[28] ), .B0(new_n1262_), .B1(\b[27] ), .Y(new_n4355_));
  OAI21X1  g04099(.A0(new_n1261_), .A1(new_n1877_), .B0(new_n4355_), .Y(new_n4356_));
  AOI21X1  g04100(.A0(new_n2004_), .A1(new_n1075_), .B0(new_n4356_), .Y(new_n4357_));
  XOR2X1   g04101(.A(new_n4357_), .B(\a[20] ), .Y(new_n4358_));
  INVX1    g04102(.A(new_n4223_), .Y(new_n4359_));
  AND2X1   g04103(.A(new_n4253_), .B(new_n4359_), .Y(new_n4360_));
  XOR2X1   g04104(.A(new_n4253_), .B(new_n4359_), .Y(new_n4361_));
  AOI21X1  g04105(.A0(new_n4361_), .A1(new_n4219_), .B0(new_n4360_), .Y(new_n4362_));
  XOR2X1   g04106(.A(new_n4250_), .B(new_n3078_), .Y(new_n4363_));
  NAND2X1  g04107(.A(new_n4363_), .B(new_n4247_), .Y(new_n4364_));
  OAI21X1  g04108(.A0(new_n4252_), .A1(new_n4226_), .B0(new_n4364_), .Y(new_n4365_));
  OR4X1    g04109(.A(new_n4229_), .B(new_n4098_), .C(new_n3907_), .D(new_n3897_), .Y(new_n4366_));
  OAI21X1  g04110(.A0(new_n4237_), .A1(new_n4231_), .B0(new_n4366_), .Y(new_n4367_));
  AND2X1   g04111(.A(new_n3901_), .B(new_n323_), .Y(new_n4368_));
  NOR3X1   g04112(.A(new_n4232_), .B(new_n3900_), .C(new_n277_), .Y(new_n4369_));
  OAI22X1  g04113(.A0(new_n3904_), .A1(new_n325_), .B0(new_n3903_), .B1(new_n297_), .Y(new_n4370_));
  NOR3X1   g04114(.A(new_n4370_), .B(new_n4369_), .C(new_n4368_), .Y(new_n4371_));
  XOR2X1   g04115(.A(new_n4371_), .B(new_n3899_), .Y(new_n4372_));
  NAND2X1  g04116(.A(new_n4229_), .B(\a[47] ), .Y(new_n4373_));
  XOR2X1   g04117(.A(\a[47] ), .B(\a[46] ), .Y(new_n4374_));
  AND2X1   g04118(.A(new_n4374_), .B(new_n4228_), .Y(new_n4375_));
  INVX1    g04119(.A(new_n4228_), .Y(new_n4376_));
  XOR2X1   g04120(.A(\a[46] ), .B(\a[45] ), .Y(new_n4377_));
  NAND2X1  g04121(.A(new_n4377_), .B(new_n4376_), .Y(new_n4378_));
  INVX1    g04122(.A(new_n4374_), .Y(new_n4379_));
  NAND2X1  g04123(.A(new_n4379_), .B(new_n4228_), .Y(new_n4380_));
  OAI22X1  g04124(.A0(new_n4380_), .A1(new_n275_), .B0(new_n4378_), .B1(new_n274_), .Y(new_n4381_));
  AOI21X1  g04125(.A0(new_n4375_), .A1(new_n263_), .B0(new_n4381_), .Y(new_n4382_));
  XOR2X1   g04126(.A(new_n4382_), .B(\a[47] ), .Y(new_n4383_));
  XOR2X1   g04127(.A(new_n4383_), .B(new_n4373_), .Y(new_n4384_));
  XOR2X1   g04128(.A(new_n4384_), .B(new_n4372_), .Y(new_n4385_));
  XOR2X1   g04129(.A(new_n4385_), .B(new_n4367_), .Y(new_n4386_));
  AOI22X1  g04130(.A0(new_n3652_), .A1(\b[7] ), .B0(new_n3651_), .B1(\b[6] ), .Y(new_n4387_));
  OAI21X1  g04131(.A0(new_n3778_), .A1(new_n395_), .B0(new_n4387_), .Y(new_n4388_));
  AOI21X1  g04132(.A0(new_n3480_), .A1(new_n394_), .B0(new_n4388_), .Y(new_n4389_));
  XOR2X1   g04133(.A(new_n4389_), .B(\a[41] ), .Y(new_n4390_));
  XOR2X1   g04134(.A(new_n4390_), .B(new_n4386_), .Y(new_n4391_));
  INVX1    g04135(.A(new_n4391_), .Y(new_n4392_));
  INVX1    g04136(.A(new_n4242_), .Y(new_n4393_));
  NOR2X1   g04137(.A(new_n4246_), .B(new_n4243_), .Y(new_n4394_));
  AOI21X1  g04138(.A0(new_n4393_), .A1(new_n4238_), .B0(new_n4394_), .Y(new_n4395_));
  XOR2X1   g04139(.A(new_n4395_), .B(new_n4392_), .Y(new_n4396_));
  AOI22X1  g04140(.A0(new_n3204_), .A1(\b[10] ), .B0(new_n3203_), .B1(\b[9] ), .Y(new_n4397_));
  OAI21X1  g04141(.A0(new_n3321_), .A1(new_n489_), .B0(new_n4397_), .Y(new_n4398_));
  AOI21X1  g04142(.A0(new_n3080_), .A1(new_n543_), .B0(new_n4398_), .Y(new_n4399_));
  XOR2X1   g04143(.A(new_n4399_), .B(\a[38] ), .Y(new_n4400_));
  NAND2X1  g04144(.A(new_n4400_), .B(new_n4396_), .Y(new_n4401_));
  XOR2X1   g04145(.A(new_n4400_), .B(new_n4396_), .Y(new_n4402_));
  INVX1    g04146(.A(new_n4402_), .Y(new_n4403_));
  NOR2X1   g04147(.A(new_n4400_), .B(new_n4396_), .Y(new_n4404_));
  AOI21X1  g04148(.A0(new_n4401_), .A1(new_n4365_), .B0(new_n4404_), .Y(new_n4405_));
  AOI22X1  g04149(.A0(new_n4405_), .A1(new_n4401_), .B0(new_n4403_), .B1(new_n4365_), .Y(new_n4406_));
  AOI22X1  g04150(.A0(new_n2813_), .A1(\b[13] ), .B0(new_n2812_), .B1(\b[12] ), .Y(new_n4407_));
  OAI21X1  g04151(.A0(new_n2946_), .A1(new_n716_), .B0(new_n4407_), .Y(new_n4408_));
  AOI21X1  g04152(.A0(new_n2652_), .A1(new_n715_), .B0(new_n4408_), .Y(new_n4409_));
  XOR2X1   g04153(.A(new_n4409_), .B(\a[35] ), .Y(new_n4410_));
  XOR2X1   g04154(.A(new_n4410_), .B(new_n4406_), .Y(new_n4411_));
  XOR2X1   g04155(.A(new_n4411_), .B(new_n4362_), .Y(new_n4412_));
  AOI22X1  g04156(.A0(new_n2545_), .A1(\b[16] ), .B0(new_n2544_), .B1(\b[15] ), .Y(new_n4413_));
  OAI21X1  g04157(.A0(new_n2543_), .A1(new_n792_), .B0(new_n4413_), .Y(new_n4414_));
  AOI21X1  g04158(.A0(new_n2260_), .A1(new_n842_), .B0(new_n4414_), .Y(new_n4415_));
  XOR2X1   g04159(.A(new_n4415_), .B(\a[32] ), .Y(new_n4416_));
  XOR2X1   g04160(.A(new_n4416_), .B(new_n4412_), .Y(new_n4417_));
  NOR2X1   g04161(.A(new_n4259_), .B(new_n4255_), .Y(new_n4418_));
  AOI21X1  g04162(.A0(new_n4260_), .A1(new_n4216_), .B0(new_n4418_), .Y(new_n4419_));
  XOR2X1   g04163(.A(new_n4419_), .B(new_n4417_), .Y(new_n4420_));
  AOI22X1  g04164(.A0(new_n2163_), .A1(\b[19] ), .B0(new_n2162_), .B1(\b[18] ), .Y(new_n4421_));
  OAI21X1  g04165(.A0(new_n2161_), .A1(new_n1118_), .B0(new_n4421_), .Y(new_n4422_));
  AOI21X1  g04166(.A0(new_n1907_), .A1(new_n1117_), .B0(new_n4422_), .Y(new_n4423_));
  XOR2X1   g04167(.A(new_n4423_), .B(\a[29] ), .Y(new_n4424_));
  XOR2X1   g04168(.A(new_n4424_), .B(new_n4420_), .Y(new_n4425_));
  OR2X1    g04169(.A(new_n4266_), .B(new_n4262_), .Y(new_n4426_));
  AND2X1   g04170(.A(new_n4266_), .B(new_n4262_), .Y(new_n4427_));
  OAI21X1  g04171(.A0(new_n4427_), .A1(new_n4213_), .B0(new_n4426_), .Y(new_n4428_));
  XOR2X1   g04172(.A(new_n4428_), .B(new_n4425_), .Y(new_n4429_));
  AOI22X1  g04173(.A0(new_n1814_), .A1(\b[22] ), .B0(new_n1813_), .B1(\b[21] ), .Y(new_n4430_));
  OAI21X1  g04174(.A0(new_n1812_), .A1(new_n1297_), .B0(new_n4430_), .Y(new_n4431_));
  AOI21X1  g04175(.A0(new_n1617_), .A1(new_n1399_), .B0(new_n4431_), .Y(new_n4432_));
  XOR2X1   g04176(.A(new_n4432_), .B(\a[26] ), .Y(new_n4433_));
  XOR2X1   g04177(.A(new_n4433_), .B(new_n4429_), .Y(new_n4434_));
  NOR2X1   g04178(.A(new_n4272_), .B(new_n4268_), .Y(new_n4435_));
  AOI21X1  g04179(.A0(new_n4278_), .A1(new_n4273_), .B0(new_n4435_), .Y(new_n4436_));
  XOR2X1   g04180(.A(new_n4436_), .B(new_n4434_), .Y(new_n4437_));
  AOI22X1  g04181(.A0(new_n1526_), .A1(\b[25] ), .B0(new_n1525_), .B1(\b[24] ), .Y(new_n4438_));
  OAI21X1  g04182(.A0(new_n1524_), .A1(new_n1591_), .B0(new_n4438_), .Y(new_n4439_));
  AOI21X1  g04183(.A0(new_n1590_), .A1(new_n1347_), .B0(new_n4439_), .Y(new_n4440_));
  XOR2X1   g04184(.A(new_n4440_), .B(\a[23] ), .Y(new_n4441_));
  XOR2X1   g04185(.A(new_n4441_), .B(new_n4437_), .Y(new_n4442_));
  OR2X1    g04186(.A(new_n4283_), .B(new_n4279_), .Y(new_n4443_));
  NAND2X1  g04187(.A(new_n4284_), .B(new_n4351_), .Y(new_n4444_));
  AND2X1   g04188(.A(new_n4444_), .B(new_n4443_), .Y(new_n4445_));
  XOR2X1   g04189(.A(new_n4445_), .B(new_n4442_), .Y(new_n4446_));
  XOR2X1   g04190(.A(new_n4446_), .B(new_n4358_), .Y(new_n4447_));
  XOR2X1   g04191(.A(new_n4447_), .B(new_n4354_), .Y(new_n4448_));
  AOI22X1  g04192(.A0(new_n1017_), .A1(\b[31] ), .B0(new_n1016_), .B1(\b[30] ), .Y(new_n4449_));
  OAI21X1  g04193(.A0(new_n1015_), .A1(new_n2359_), .B0(new_n4449_), .Y(new_n4450_));
  AOI21X1  g04194(.A0(new_n2358_), .A1(new_n882_), .B0(new_n4450_), .Y(new_n4451_));
  XOR2X1   g04195(.A(new_n4451_), .B(\a[17] ), .Y(new_n4452_));
  XOR2X1   g04196(.A(new_n4452_), .B(new_n4448_), .Y(new_n4453_));
  XOR2X1   g04197(.A(new_n4453_), .B(new_n4347_), .Y(new_n4454_));
  AOI22X1  g04198(.A0(new_n818_), .A1(\b[34] ), .B0(new_n817_), .B1(\b[33] ), .Y(new_n4455_));
  OAI21X1  g04199(.A0(new_n816_), .A1(new_n2612_), .B0(new_n4455_), .Y(new_n4456_));
  AOI21X1  g04200(.A0(new_n2759_), .A1(new_n668_), .B0(new_n4456_), .Y(new_n4457_));
  XOR2X1   g04201(.A(new_n4457_), .B(\a[14] ), .Y(new_n4458_));
  XOR2X1   g04202(.A(new_n4458_), .B(new_n4454_), .Y(new_n4459_));
  XOR2X1   g04203(.A(new_n4353_), .B(new_n4211_), .Y(new_n4460_));
  XOR2X1   g04204(.A(new_n4295_), .B(new_n4460_), .Y(new_n4461_));
  XOR2X1   g04205(.A(new_n4461_), .B(new_n4209_), .Y(new_n4462_));
  NOR2X1   g04206(.A(new_n4301_), .B(new_n4462_), .Y(new_n4463_));
  XOR2X1   g04207(.A(new_n4301_), .B(new_n4462_), .Y(new_n4464_));
  AOI21X1  g04208(.A0(new_n4464_), .A1(new_n4206_), .B0(new_n4463_), .Y(new_n4465_));
  XOR2X1   g04209(.A(new_n4465_), .B(new_n4459_), .Y(new_n4466_));
  AOI22X1  g04210(.A0(new_n603_), .A1(\b[37] ), .B0(new_n602_), .B1(\b[36] ), .Y(new_n4467_));
  OAI21X1  g04211(.A0(new_n601_), .A1(new_n3156_), .B0(new_n4467_), .Y(new_n4468_));
  AOI21X1  g04212(.A0(new_n3155_), .A1(new_n518_), .B0(new_n4468_), .Y(new_n4469_));
  XOR2X1   g04213(.A(new_n4469_), .B(\a[11] ), .Y(new_n4470_));
  XOR2X1   g04214(.A(new_n4470_), .B(new_n4466_), .Y(new_n4471_));
  OR2X1    g04215(.A(new_n4158_), .B(new_n4196_), .Y(new_n4472_));
  OAI21X1  g04216(.A0(new_n4165_), .A1(new_n4159_), .B0(new_n4472_), .Y(new_n4473_));
  NOR2X1   g04217(.A(new_n4307_), .B(new_n4303_), .Y(new_n4474_));
  AOI21X1  g04218(.A0(new_n4308_), .A1(new_n4473_), .B0(new_n4474_), .Y(new_n4475_));
  XOR2X1   g04219(.A(new_n4475_), .B(new_n4471_), .Y(new_n4476_));
  AOI22X1  g04220(.A0(new_n469_), .A1(\b[40] ), .B0(new_n468_), .B1(\b[39] ), .Y(new_n4477_));
  OAI21X1  g04221(.A0(new_n467_), .A1(new_n3575_), .B0(new_n4477_), .Y(new_n4478_));
  AOI21X1  g04222(.A0(new_n3574_), .A1(new_n404_), .B0(new_n4478_), .Y(new_n4479_));
  XOR2X1   g04223(.A(new_n4479_), .B(\a[8] ), .Y(new_n4480_));
  NAND2X1  g04224(.A(new_n4480_), .B(new_n4476_), .Y(new_n4481_));
  NOR2X1   g04225(.A(new_n4313_), .B(new_n4309_), .Y(new_n4482_));
  OR2X1    g04226(.A(new_n4170_), .B(new_n4315_), .Y(new_n4483_));
  OAI21X1  g04227(.A0(new_n4171_), .A1(new_n4047_), .B0(new_n4483_), .Y(new_n4484_));
  AOI21X1  g04228(.A0(new_n4484_), .A1(new_n4314_), .B0(new_n4482_), .Y(new_n4485_));
  OR2X1    g04229(.A(new_n4480_), .B(new_n4476_), .Y(new_n4486_));
  AOI21X1  g04230(.A0(new_n4481_), .A1(new_n4486_), .B0(new_n4485_), .Y(new_n4487_));
  OR2X1    g04231(.A(new_n4313_), .B(new_n4309_), .Y(new_n4488_));
  XOR2X1   g04232(.A(new_n4308_), .B(new_n4473_), .Y(new_n4489_));
  XOR2X1   g04233(.A(new_n4313_), .B(new_n4489_), .Y(new_n4490_));
  OAI21X1  g04234(.A0(new_n4318_), .A1(new_n4490_), .B0(new_n4488_), .Y(new_n4491_));
  NOR2X1   g04235(.A(new_n4480_), .B(new_n4476_), .Y(new_n4492_));
  AOI21X1  g04236(.A0(new_n4481_), .A1(new_n4491_), .B0(new_n4492_), .Y(new_n4493_));
  AOI21X1  g04237(.A0(new_n4493_), .A1(new_n4481_), .B0(new_n4487_), .Y(new_n4494_));
  AOI22X1  g04238(.A0(new_n369_), .A1(\b[43] ), .B0(new_n368_), .B1(\b[42] ), .Y(new_n4495_));
  OAI21X1  g04239(.A0(new_n367_), .A1(new_n4015_), .B0(new_n4495_), .Y(new_n4496_));
  AOI21X1  g04240(.A0(new_n4014_), .A1(new_n308_), .B0(new_n4496_), .Y(new_n4497_));
  XOR2X1   g04241(.A(new_n4497_), .B(\a[5] ), .Y(new_n4498_));
  INVX1    g04242(.A(new_n4498_), .Y(new_n4499_));
  XOR2X1   g04243(.A(new_n4499_), .B(new_n4494_), .Y(new_n4500_));
  NOR2X1   g04244(.A(new_n4323_), .B(new_n4319_), .Y(new_n4501_));
  NAND2X1  g04245(.A(new_n4172_), .B(new_n4186_), .Y(new_n4502_));
  OAI21X1  g04246(.A0(new_n4173_), .A1(new_n4033_), .B0(new_n4502_), .Y(new_n4503_));
  AOI21X1  g04247(.A0(new_n4503_), .A1(new_n4324_), .B0(new_n4501_), .Y(new_n4504_));
  XOR2X1   g04248(.A(new_n4504_), .B(new_n4500_), .Y(new_n4505_));
  NAND2X1  g04249(.A(\b[45] ), .B(\b[44] ), .Y(new_n4506_));
  OAI21X1  g04250(.A0(new_n4337_), .A1(new_n4335_), .B0(new_n4506_), .Y(new_n4507_));
  XOR2X1   g04251(.A(\b[46] ), .B(\b[45] ), .Y(new_n4508_));
  XOR2X1   g04252(.A(new_n4508_), .B(new_n4507_), .Y(new_n4509_));
  AOI22X1  g04253(.A0(new_n267_), .A1(\b[46] ), .B0(new_n266_), .B1(\b[45] ), .Y(new_n4510_));
  OAI21X1  g04254(.A0(new_n350_), .A1(new_n4336_), .B0(new_n4510_), .Y(new_n4511_));
  AOI21X1  g04255(.A0(new_n4509_), .A1(new_n318_), .B0(new_n4511_), .Y(new_n4512_));
  XOR2X1   g04256(.A(new_n4512_), .B(\a[2] ), .Y(new_n4513_));
  XOR2X1   g04257(.A(new_n4513_), .B(new_n4505_), .Y(new_n4514_));
  OR2X1    g04258(.A(new_n4343_), .B(new_n4333_), .Y(new_n4515_));
  OAI21X1  g04259(.A0(new_n4189_), .A1(new_n4185_), .B0(new_n4344_), .Y(new_n4516_));
  AND2X1   g04260(.A(new_n4516_), .B(new_n4515_), .Y(new_n4517_));
  XOR2X1   g04261(.A(new_n4517_), .B(new_n4514_), .Y(\f[46] ));
  OR2X1    g04262(.A(new_n4498_), .B(new_n4494_), .Y(new_n4519_));
  OAI21X1  g04263(.A0(new_n4504_), .A1(new_n4500_), .B0(new_n4519_), .Y(new_n4520_));
  OR2X1    g04264(.A(new_n4452_), .B(new_n4448_), .Y(new_n4521_));
  INVX1    g04265(.A(new_n4452_), .Y(new_n4522_));
  XOR2X1   g04266(.A(new_n4522_), .B(new_n4448_), .Y(new_n4523_));
  OAI21X1  g04267(.A0(new_n4523_), .A1(new_n4347_), .B0(new_n4521_), .Y(new_n4524_));
  AOI22X1  g04268(.A0(new_n1017_), .A1(\b[32] ), .B0(new_n1016_), .B1(\b[31] ), .Y(new_n4525_));
  OAI21X1  g04269(.A0(new_n1015_), .A1(new_n2356_), .B0(new_n4525_), .Y(new_n4526_));
  AOI21X1  g04270(.A0(new_n2495_), .A1(new_n882_), .B0(new_n4526_), .Y(new_n4527_));
  XOR2X1   g04271(.A(new_n4527_), .B(\a[17] ), .Y(new_n4528_));
  INVX1    g04272(.A(new_n4358_), .Y(new_n4529_));
  AND2X1   g04273(.A(new_n4446_), .B(new_n4529_), .Y(new_n4530_));
  XOR2X1   g04274(.A(new_n4446_), .B(new_n4529_), .Y(new_n4531_));
  AOI21X1  g04275(.A0(new_n4531_), .A1(new_n4354_), .B0(new_n4530_), .Y(new_n4532_));
  AOI22X1  g04276(.A0(new_n1263_), .A1(\b[29] ), .B0(new_n1262_), .B1(\b[28] ), .Y(new_n4533_));
  OAI21X1  g04277(.A0(new_n1261_), .A1(new_n2126_), .B0(new_n4533_), .Y(new_n4534_));
  AOI21X1  g04278(.A0(new_n2125_), .A1(new_n1075_), .B0(new_n4534_), .Y(new_n4535_));
  XOR2X1   g04279(.A(new_n4535_), .B(\a[20] ), .Y(new_n4536_));
  XOR2X1   g04280(.A(new_n4440_), .B(new_n1351_), .Y(new_n4537_));
  AND2X1   g04281(.A(new_n4537_), .B(new_n4437_), .Y(new_n4538_));
  AOI21X1  g04282(.A0(new_n4444_), .A1(new_n4443_), .B0(new_n4442_), .Y(new_n4539_));
  OR2X1    g04283(.A(new_n4539_), .B(new_n4538_), .Y(new_n4540_));
  AND2X1   g04284(.A(new_n4361_), .B(new_n4219_), .Y(new_n4541_));
  OR2X1    g04285(.A(new_n4541_), .B(new_n4360_), .Y(new_n4542_));
  XOR2X1   g04286(.A(new_n4411_), .B(new_n4542_), .Y(new_n4543_));
  XOR2X1   g04287(.A(new_n4416_), .B(new_n4543_), .Y(new_n4544_));
  XOR2X1   g04288(.A(new_n4419_), .B(new_n4544_), .Y(new_n4545_));
  XOR2X1   g04289(.A(new_n4424_), .B(new_n4545_), .Y(new_n4546_));
  XOR2X1   g04290(.A(new_n4428_), .B(new_n4546_), .Y(new_n4547_));
  OR2X1    g04291(.A(new_n4433_), .B(new_n4547_), .Y(new_n4548_));
  OAI21X1  g04292(.A0(new_n4436_), .A1(new_n4434_), .B0(new_n4548_), .Y(new_n4549_));
  OR2X1    g04293(.A(new_n4416_), .B(new_n4412_), .Y(new_n4550_));
  OAI21X1  g04294(.A0(new_n4419_), .A1(new_n4544_), .B0(new_n4550_), .Y(new_n4551_));
  AOI22X1  g04295(.A0(new_n2545_), .A1(\b[17] ), .B0(new_n2544_), .B1(\b[16] ), .Y(new_n4552_));
  OAI21X1  g04296(.A0(new_n2543_), .A1(new_n977_), .B0(new_n4552_), .Y(new_n4553_));
  AOI21X1  g04297(.A0(new_n2260_), .A1(new_n976_), .B0(new_n4553_), .Y(new_n4554_));
  XOR2X1   g04298(.A(new_n4554_), .B(\a[32] ), .Y(new_n4555_));
  NOR2X1   g04299(.A(new_n4410_), .B(new_n4406_), .Y(new_n4556_));
  AOI21X1  g04300(.A0(new_n4411_), .A1(new_n4542_), .B0(new_n4556_), .Y(new_n4557_));
  INVX1    g04301(.A(new_n4386_), .Y(new_n4558_));
  OR2X1    g04302(.A(new_n4395_), .B(new_n4391_), .Y(new_n4559_));
  OAI21X1  g04303(.A0(new_n4390_), .A1(new_n4558_), .B0(new_n4559_), .Y(new_n4560_));
  AOI22X1  g04304(.A0(new_n3652_), .A1(\b[8] ), .B0(new_n3651_), .B1(\b[7] ), .Y(new_n4561_));
  OAI21X1  g04305(.A0(new_n3778_), .A1(new_n392_), .B0(new_n4561_), .Y(new_n4562_));
  AOI21X1  g04306(.A0(new_n3480_), .A1(new_n454_), .B0(new_n4562_), .Y(new_n4563_));
  XOR2X1   g04307(.A(new_n4563_), .B(\a[41] ), .Y(new_n4564_));
  AND2X1   g04308(.A(new_n4384_), .B(new_n4372_), .Y(new_n4565_));
  AOI21X1  g04309(.A0(new_n4385_), .A1(new_n4367_), .B0(new_n4565_), .Y(new_n4566_));
  NAND3X1  g04310(.A(new_n4382_), .B(new_n4229_), .C(\a[47] ), .Y(new_n4567_));
  INVX1    g04311(.A(\a[47] ), .Y(new_n4568_));
  NAND2X1  g04312(.A(new_n4375_), .B(new_n341_), .Y(new_n4569_));
  OR4X1    g04313(.A(new_n4377_), .B(new_n4379_), .C(new_n4228_), .D(new_n274_), .Y(new_n4570_));
  AND2X1   g04314(.A(new_n4377_), .B(new_n4376_), .Y(new_n4571_));
  AND2X1   g04315(.A(new_n4379_), .B(new_n4228_), .Y(new_n4572_));
  AOI22X1  g04316(.A0(new_n4572_), .A1(\b[2] ), .B0(new_n4571_), .B1(\b[1] ), .Y(new_n4573_));
  NAND3X1  g04317(.A(new_n4573_), .B(new_n4570_), .C(new_n4569_), .Y(new_n4574_));
  XOR2X1   g04318(.A(new_n4574_), .B(new_n4568_), .Y(new_n4575_));
  XOR2X1   g04319(.A(new_n4575_), .B(new_n4567_), .Y(new_n4576_));
  AOI22X1  g04320(.A0(new_n4095_), .A1(\b[5] ), .B0(new_n4094_), .B1(\b[4] ), .Y(new_n4577_));
  OAI21X1  g04321(.A0(new_n4233_), .A1(new_n297_), .B0(new_n4577_), .Y(new_n4578_));
  AOI21X1  g04322(.A0(new_n3901_), .A1(new_n349_), .B0(new_n4578_), .Y(new_n4579_));
  XOR2X1   g04323(.A(new_n4579_), .B(\a[44] ), .Y(new_n4580_));
  XOR2X1   g04324(.A(new_n4580_), .B(new_n4576_), .Y(new_n4581_));
  XOR2X1   g04325(.A(new_n4581_), .B(new_n4566_), .Y(new_n4582_));
  XOR2X1   g04326(.A(new_n4582_), .B(new_n4564_), .Y(new_n4583_));
  XOR2X1   g04327(.A(new_n4583_), .B(new_n4560_), .Y(new_n4584_));
  AOI22X1  g04328(.A0(new_n3204_), .A1(\b[11] ), .B0(new_n3203_), .B1(\b[10] ), .Y(new_n4585_));
  OAI21X1  g04329(.A0(new_n3321_), .A1(new_n590_), .B0(new_n4585_), .Y(new_n4586_));
  AOI21X1  g04330(.A0(new_n3080_), .A1(new_n589_), .B0(new_n4586_), .Y(new_n4587_));
  XOR2X1   g04331(.A(new_n4587_), .B(\a[38] ), .Y(new_n4588_));
  XOR2X1   g04332(.A(new_n4588_), .B(new_n4584_), .Y(new_n4589_));
  XOR2X1   g04333(.A(new_n4589_), .B(new_n4405_), .Y(new_n4590_));
  AOI22X1  g04334(.A0(new_n2813_), .A1(\b[14] ), .B0(new_n2812_), .B1(\b[13] ), .Y(new_n4591_));
  OAI21X1  g04335(.A0(new_n2946_), .A1(new_n713_), .B0(new_n4591_), .Y(new_n4592_));
  AOI21X1  g04336(.A0(new_n2652_), .A1(new_n734_), .B0(new_n4592_), .Y(new_n4593_));
  XOR2X1   g04337(.A(new_n4593_), .B(\a[35] ), .Y(new_n4594_));
  INVX1    g04338(.A(new_n4594_), .Y(new_n4595_));
  XOR2X1   g04339(.A(new_n4595_), .B(new_n4590_), .Y(new_n4596_));
  XOR2X1   g04340(.A(new_n4596_), .B(new_n4557_), .Y(new_n4597_));
  XOR2X1   g04341(.A(new_n4597_), .B(new_n4555_), .Y(new_n4598_));
  XOR2X1   g04342(.A(new_n4598_), .B(new_n4551_), .Y(new_n4599_));
  AOI22X1  g04343(.A0(new_n2163_), .A1(\b[20] ), .B0(new_n2162_), .B1(\b[19] ), .Y(new_n4600_));
  OAI21X1  g04344(.A0(new_n2161_), .A1(new_n1115_), .B0(new_n4600_), .Y(new_n4601_));
  AOI21X1  g04345(.A0(new_n1907_), .A1(new_n1217_), .B0(new_n4601_), .Y(new_n4602_));
  XOR2X1   g04346(.A(new_n4602_), .B(\a[29] ), .Y(new_n4603_));
  XOR2X1   g04347(.A(new_n4603_), .B(new_n4599_), .Y(new_n4604_));
  NOR2X1   g04348(.A(new_n4424_), .B(new_n4420_), .Y(new_n4605_));
  AOI21X1  g04349(.A0(new_n4428_), .A1(new_n4425_), .B0(new_n4605_), .Y(new_n4606_));
  XOR2X1   g04350(.A(new_n4606_), .B(new_n4604_), .Y(new_n4607_));
  AOI22X1  g04351(.A0(new_n1814_), .A1(\b[23] ), .B0(new_n1813_), .B1(\b[22] ), .Y(new_n4608_));
  OAI21X1  g04352(.A0(new_n1812_), .A1(new_n1482_), .B0(new_n4608_), .Y(new_n4609_));
  AOI21X1  g04353(.A0(new_n1617_), .A1(new_n1481_), .B0(new_n4609_), .Y(new_n4610_));
  XOR2X1   g04354(.A(new_n4610_), .B(\a[26] ), .Y(new_n4611_));
  NAND2X1  g04355(.A(new_n4611_), .B(new_n4607_), .Y(new_n4612_));
  XOR2X1   g04356(.A(new_n4610_), .B(new_n1621_), .Y(new_n4613_));
  XOR2X1   g04357(.A(new_n4613_), .B(new_n4607_), .Y(new_n4614_));
  NOR2X1   g04358(.A(new_n4611_), .B(new_n4607_), .Y(new_n4615_));
  AOI21X1  g04359(.A0(new_n4612_), .A1(new_n4549_), .B0(new_n4615_), .Y(new_n4616_));
  AOI22X1  g04360(.A0(new_n4616_), .A1(new_n4612_), .B0(new_n4614_), .B1(new_n4549_), .Y(new_n4617_));
  AOI22X1  g04361(.A0(new_n1526_), .A1(\b[26] ), .B0(new_n1525_), .B1(\b[25] ), .Y(new_n4618_));
  OAI21X1  g04362(.A0(new_n1524_), .A1(new_n1588_), .B0(new_n4618_), .Y(new_n4619_));
  AOI21X1  g04363(.A0(new_n1783_), .A1(new_n1347_), .B0(new_n4619_), .Y(new_n4620_));
  XOR2X1   g04364(.A(new_n4620_), .B(\a[23] ), .Y(new_n4621_));
  XOR2X1   g04365(.A(new_n4621_), .B(new_n4617_), .Y(new_n4622_));
  XOR2X1   g04366(.A(new_n4622_), .B(new_n4540_), .Y(new_n4623_));
  XOR2X1   g04367(.A(new_n4623_), .B(new_n4536_), .Y(new_n4624_));
  XOR2X1   g04368(.A(new_n4624_), .B(new_n4532_), .Y(new_n4625_));
  XOR2X1   g04369(.A(new_n4625_), .B(new_n4528_), .Y(new_n4626_));
  XOR2X1   g04370(.A(new_n4626_), .B(new_n4524_), .Y(new_n4627_));
  AOI22X1  g04371(.A0(new_n818_), .A1(\b[35] ), .B0(new_n817_), .B1(\b[34] ), .Y(new_n4628_));
  OAI21X1  g04372(.A0(new_n816_), .A1(new_n2893_), .B0(new_n4628_), .Y(new_n4629_));
  AOI21X1  g04373(.A0(new_n2892_), .A1(new_n668_), .B0(new_n4629_), .Y(new_n4630_));
  XOR2X1   g04374(.A(new_n4630_), .B(\a[14] ), .Y(new_n4631_));
  XOR2X1   g04375(.A(new_n4631_), .B(new_n4627_), .Y(new_n4632_));
  NOR2X1   g04376(.A(new_n4458_), .B(new_n4454_), .Y(new_n4633_));
  AND2X1   g04377(.A(new_n4152_), .B(new_n4054_), .Y(new_n4634_));
  AOI21X1  g04378(.A0(new_n4153_), .A1(new_n4050_), .B0(new_n4634_), .Y(new_n4635_));
  OR2X1    g04379(.A(new_n4301_), .B(new_n4462_), .Y(new_n4636_));
  OAI21X1  g04380(.A0(new_n4302_), .A1(new_n4635_), .B0(new_n4636_), .Y(new_n4637_));
  AOI21X1  g04381(.A0(new_n4637_), .A1(new_n4459_), .B0(new_n4633_), .Y(new_n4638_));
  XOR2X1   g04382(.A(new_n4638_), .B(new_n4632_), .Y(new_n4639_));
  AOI22X1  g04383(.A0(new_n603_), .A1(\b[38] ), .B0(new_n602_), .B1(\b[37] ), .Y(new_n4640_));
  OAI21X1  g04384(.A0(new_n601_), .A1(new_n3276_), .B0(new_n4640_), .Y(new_n4641_));
  AOI21X1  g04385(.A0(new_n3275_), .A1(new_n518_), .B0(new_n4641_), .Y(new_n4642_));
  XOR2X1   g04386(.A(new_n4642_), .B(\a[11] ), .Y(new_n4643_));
  XOR2X1   g04387(.A(new_n4643_), .B(new_n4639_), .Y(new_n4644_));
  NOR2X1   g04388(.A(new_n4470_), .B(new_n4466_), .Y(new_n4645_));
  OR2X1    g04389(.A(new_n4307_), .B(new_n4303_), .Y(new_n4646_));
  AND2X1   g04390(.A(new_n4307_), .B(new_n4303_), .Y(new_n4647_));
  OAI21X1  g04391(.A0(new_n4647_), .A1(new_n4203_), .B0(new_n4646_), .Y(new_n4648_));
  AOI21X1  g04392(.A0(new_n4648_), .A1(new_n4471_), .B0(new_n4645_), .Y(new_n4649_));
  XOR2X1   g04393(.A(new_n4649_), .B(new_n4644_), .Y(new_n4650_));
  AOI22X1  g04394(.A0(new_n469_), .A1(\b[41] ), .B0(new_n468_), .B1(\b[40] ), .Y(new_n4651_));
  OAI21X1  g04395(.A0(new_n467_), .A1(new_n3723_), .B0(new_n4651_), .Y(new_n4652_));
  AOI21X1  g04396(.A0(new_n3722_), .A1(new_n404_), .B0(new_n4652_), .Y(new_n4653_));
  XOR2X1   g04397(.A(new_n4653_), .B(\a[8] ), .Y(new_n4654_));
  NAND2X1  g04398(.A(new_n4654_), .B(new_n4650_), .Y(new_n4655_));
  OR2X1    g04399(.A(new_n4654_), .B(new_n4650_), .Y(new_n4656_));
  AOI21X1  g04400(.A0(new_n4655_), .A1(new_n4656_), .B0(new_n4493_), .Y(new_n4657_));
  AND2X1   g04401(.A(new_n4480_), .B(new_n4476_), .Y(new_n4658_));
  OAI21X1  g04402(.A0(new_n4658_), .A1(new_n4485_), .B0(new_n4486_), .Y(new_n4659_));
  NOR2X1   g04403(.A(new_n4654_), .B(new_n4650_), .Y(new_n4660_));
  AOI21X1  g04404(.A0(new_n4655_), .A1(new_n4659_), .B0(new_n4660_), .Y(new_n4661_));
  AOI21X1  g04405(.A0(new_n4661_), .A1(new_n4655_), .B0(new_n4657_), .Y(new_n4662_));
  AOI22X1  g04406(.A0(new_n369_), .A1(\b[44] ), .B0(new_n368_), .B1(\b[43] ), .Y(new_n4663_));
  OAI21X1  g04407(.A0(new_n367_), .A1(new_n4012_), .B0(new_n4663_), .Y(new_n4664_));
  AOI21X1  g04408(.A0(new_n4178_), .A1(new_n308_), .B0(new_n4664_), .Y(new_n4665_));
  XOR2X1   g04409(.A(new_n4665_), .B(\a[5] ), .Y(new_n4666_));
  XOR2X1   g04410(.A(new_n4666_), .B(new_n4662_), .Y(new_n4667_));
  XOR2X1   g04411(.A(new_n4667_), .B(new_n4520_), .Y(new_n4668_));
  AND2X1   g04412(.A(\b[46] ), .B(\b[45] ), .Y(new_n4669_));
  AOI21X1  g04413(.A0(new_n4508_), .A1(new_n4507_), .B0(new_n4669_), .Y(new_n4670_));
  XOR2X1   g04414(.A(\b[47] ), .B(\b[46] ), .Y(new_n4671_));
  INVX1    g04415(.A(new_n4671_), .Y(new_n4672_));
  XOR2X1   g04416(.A(new_n4672_), .B(new_n4670_), .Y(new_n4673_));
  INVX1    g04417(.A(\b[45] ), .Y(new_n4674_));
  AOI22X1  g04418(.A0(new_n267_), .A1(\b[47] ), .B0(new_n266_), .B1(\b[46] ), .Y(new_n4675_));
  OAI21X1  g04419(.A0(new_n350_), .A1(new_n4674_), .B0(new_n4675_), .Y(new_n4676_));
  AOI21X1  g04420(.A0(new_n4673_), .A1(new_n318_), .B0(new_n4676_), .Y(new_n4677_));
  XOR2X1   g04421(.A(new_n4677_), .B(new_n257_), .Y(new_n4678_));
  XOR2X1   g04422(.A(new_n4678_), .B(new_n4668_), .Y(new_n4679_));
  XOR2X1   g04423(.A(new_n4498_), .B(new_n4494_), .Y(new_n4680_));
  XOR2X1   g04424(.A(new_n4504_), .B(new_n4680_), .Y(new_n4681_));
  NOR2X1   g04425(.A(new_n4513_), .B(new_n4681_), .Y(new_n4682_));
  AOI21X1  g04426(.A0(new_n4516_), .A1(new_n4515_), .B0(new_n4514_), .Y(new_n4683_));
  OR2X1    g04427(.A(new_n4683_), .B(new_n4682_), .Y(new_n4684_));
  XOR2X1   g04428(.A(new_n4684_), .B(new_n4679_), .Y(\f[47] ));
  NAND2X1  g04429(.A(new_n4678_), .B(new_n4668_), .Y(new_n4686_));
  OAI21X1  g04430(.A0(new_n4683_), .A1(new_n4682_), .B0(new_n4679_), .Y(new_n4687_));
  AND2X1   g04431(.A(new_n4687_), .B(new_n4686_), .Y(new_n4688_));
  NAND2X1  g04432(.A(\b[47] ), .B(\b[46] ), .Y(new_n4689_));
  OAI21X1  g04433(.A0(new_n4672_), .A1(new_n4670_), .B0(new_n4689_), .Y(new_n4690_));
  XOR2X1   g04434(.A(\b[48] ), .B(\b[47] ), .Y(new_n4691_));
  XOR2X1   g04435(.A(new_n4691_), .B(new_n4690_), .Y(new_n4692_));
  INVX1    g04436(.A(\b[46] ), .Y(new_n4693_));
  AOI22X1  g04437(.A0(new_n267_), .A1(\b[48] ), .B0(new_n266_), .B1(\b[47] ), .Y(new_n4694_));
  OAI21X1  g04438(.A0(new_n350_), .A1(new_n4693_), .B0(new_n4694_), .Y(new_n4695_));
  AOI21X1  g04439(.A0(new_n4692_), .A1(new_n318_), .B0(new_n4695_), .Y(new_n4696_));
  XOR2X1   g04440(.A(new_n4696_), .B(\a[2] ), .Y(new_n4697_));
  NOR2X1   g04441(.A(new_n4666_), .B(new_n4662_), .Y(new_n4698_));
  AOI21X1  g04442(.A0(new_n4667_), .A1(new_n4520_), .B0(new_n4698_), .Y(new_n4699_));
  OR2X1    g04443(.A(new_n4631_), .B(new_n4627_), .Y(new_n4700_));
  INVX1    g04444(.A(new_n4528_), .Y(new_n4701_));
  XOR2X1   g04445(.A(new_n4625_), .B(new_n4701_), .Y(new_n4702_));
  XOR2X1   g04446(.A(new_n4702_), .B(new_n4524_), .Y(new_n4703_));
  XOR2X1   g04447(.A(new_n4631_), .B(new_n4703_), .Y(new_n4704_));
  OAI21X1  g04448(.A0(new_n4638_), .A1(new_n4704_), .B0(new_n4700_), .Y(new_n4705_));
  AND2X1   g04449(.A(new_n4625_), .B(new_n4701_), .Y(new_n4706_));
  AOI21X1  g04450(.A0(new_n4702_), .A1(new_n4524_), .B0(new_n4706_), .Y(new_n4707_));
  INVX1    g04451(.A(new_n4536_), .Y(new_n4708_));
  NAND2X1  g04452(.A(new_n4623_), .B(new_n4708_), .Y(new_n4709_));
  OAI21X1  g04453(.A0(new_n4624_), .A1(new_n4532_), .B0(new_n4709_), .Y(new_n4710_));
  OR2X1    g04454(.A(new_n4621_), .B(new_n4617_), .Y(new_n4711_));
  OAI21X1  g04455(.A0(new_n4539_), .A1(new_n4538_), .B0(new_n4622_), .Y(new_n4712_));
  AND2X1   g04456(.A(new_n4712_), .B(new_n4711_), .Y(new_n4713_));
  OR2X1    g04457(.A(new_n4594_), .B(new_n4590_), .Y(new_n4714_));
  OAI21X1  g04458(.A0(new_n4596_), .A1(new_n4557_), .B0(new_n4714_), .Y(new_n4715_));
  AOI22X1  g04459(.A0(new_n2813_), .A1(\b[15] ), .B0(new_n2812_), .B1(\b[14] ), .Y(new_n4716_));
  OAI21X1  g04460(.A0(new_n2946_), .A1(new_n795_), .B0(new_n4716_), .Y(new_n4717_));
  AOI21X1  g04461(.A0(new_n2652_), .A1(new_n794_), .B0(new_n4717_), .Y(new_n4718_));
  XOR2X1   g04462(.A(new_n4718_), .B(\a[35] ), .Y(new_n4719_));
  INVX1    g04463(.A(new_n4719_), .Y(new_n4720_));
  NOR2X1   g04464(.A(new_n4588_), .B(new_n4584_), .Y(new_n4721_));
  INVX1    g04465(.A(new_n4721_), .Y(new_n4722_));
  AND2X1   g04466(.A(new_n4402_), .B(new_n4365_), .Y(new_n4723_));
  OAI21X1  g04467(.A0(new_n4723_), .A1(new_n4404_), .B0(new_n4589_), .Y(new_n4724_));
  AND2X1   g04468(.A(new_n4724_), .B(new_n4722_), .Y(new_n4725_));
  AOI22X1  g04469(.A0(new_n3204_), .A1(\b[12] ), .B0(new_n3203_), .B1(\b[11] ), .Y(new_n4726_));
  OAI21X1  g04470(.A0(new_n3321_), .A1(new_n587_), .B0(new_n4726_), .Y(new_n4727_));
  AOI21X1  g04471(.A0(new_n3080_), .A1(new_n635_), .B0(new_n4727_), .Y(new_n4728_));
  XOR2X1   g04472(.A(new_n4728_), .B(\a[38] ), .Y(new_n4729_));
  INVX1    g04473(.A(new_n4564_), .Y(new_n4730_));
  AND2X1   g04474(.A(new_n4582_), .B(new_n4730_), .Y(new_n4731_));
  INVX1    g04475(.A(new_n4583_), .Y(new_n4732_));
  AOI21X1  g04476(.A0(new_n4732_), .A1(new_n4560_), .B0(new_n4731_), .Y(new_n4733_));
  OR2X1    g04477(.A(new_n4575_), .B(new_n4567_), .Y(new_n4734_));
  XOR2X1   g04478(.A(\a[48] ), .B(new_n4568_), .Y(new_n4735_));
  OR2X1    g04479(.A(new_n4735_), .B(new_n274_), .Y(new_n4736_));
  INVX1    g04480(.A(new_n4736_), .Y(new_n4737_));
  XOR2X1   g04481(.A(new_n4737_), .B(new_n4734_), .Y(new_n4738_));
  OR2X1    g04482(.A(new_n4377_), .B(new_n4228_), .Y(new_n4739_));
  OR2X1    g04483(.A(new_n4739_), .B(new_n4379_), .Y(new_n4740_));
  AOI22X1  g04484(.A0(new_n4572_), .A1(\b[3] ), .B0(new_n4571_), .B1(\b[2] ), .Y(new_n4741_));
  OAI21X1  g04485(.A0(new_n4740_), .A1(new_n275_), .B0(new_n4741_), .Y(new_n4742_));
  AOI21X1  g04486(.A0(new_n4375_), .A1(new_n366_), .B0(new_n4742_), .Y(new_n4743_));
  XOR2X1   g04487(.A(new_n4743_), .B(\a[47] ), .Y(new_n4744_));
  XOR2X1   g04488(.A(new_n4744_), .B(new_n4738_), .Y(new_n4745_));
  AOI22X1  g04489(.A0(new_n4095_), .A1(\b[6] ), .B0(new_n4094_), .B1(\b[5] ), .Y(new_n4746_));
  OAI21X1  g04490(.A0(new_n4233_), .A1(new_n325_), .B0(new_n4746_), .Y(new_n4747_));
  AOI21X1  g04491(.A0(new_n3901_), .A1(new_n378_), .B0(new_n4747_), .Y(new_n4748_));
  XOR2X1   g04492(.A(new_n4748_), .B(\a[44] ), .Y(new_n4749_));
  XOR2X1   g04493(.A(new_n4749_), .B(new_n4745_), .Y(new_n4750_));
  INVX1    g04494(.A(new_n4580_), .Y(new_n4751_));
  NOR2X1   g04495(.A(new_n4581_), .B(new_n4566_), .Y(new_n4752_));
  AOI21X1  g04496(.A0(new_n4751_), .A1(new_n4576_), .B0(new_n4752_), .Y(new_n4753_));
  XOR2X1   g04497(.A(new_n4753_), .B(new_n4750_), .Y(new_n4754_));
  INVX1    g04498(.A(new_n4754_), .Y(new_n4755_));
  AOI22X1  g04499(.A0(new_n3652_), .A1(\b[9] ), .B0(new_n3651_), .B1(\b[8] ), .Y(new_n4756_));
  OAI21X1  g04500(.A0(new_n3778_), .A1(new_n492_), .B0(new_n4756_), .Y(new_n4757_));
  AOI21X1  g04501(.A0(new_n3480_), .A1(new_n491_), .B0(new_n4757_), .Y(new_n4758_));
  XOR2X1   g04502(.A(new_n4758_), .B(\a[41] ), .Y(new_n4759_));
  XOR2X1   g04503(.A(new_n4759_), .B(new_n4755_), .Y(new_n4760_));
  INVX1    g04504(.A(new_n4760_), .Y(new_n4761_));
  XOR2X1   g04505(.A(new_n4761_), .B(new_n4733_), .Y(new_n4762_));
  XOR2X1   g04506(.A(new_n4762_), .B(new_n4729_), .Y(new_n4763_));
  XOR2X1   g04507(.A(new_n4763_), .B(new_n4725_), .Y(new_n4764_));
  XOR2X1   g04508(.A(new_n4764_), .B(new_n4720_), .Y(new_n4765_));
  XOR2X1   g04509(.A(new_n4765_), .B(new_n4715_), .Y(new_n4766_));
  AOI22X1  g04510(.A0(new_n2545_), .A1(\b[18] ), .B0(new_n2544_), .B1(\b[17] ), .Y(new_n4767_));
  OAI21X1  g04511(.A0(new_n2543_), .A1(new_n974_), .B0(new_n4767_), .Y(new_n4768_));
  AOI21X1  g04512(.A0(new_n2260_), .A1(new_n1042_), .B0(new_n4768_), .Y(new_n4769_));
  XOR2X1   g04513(.A(new_n4769_), .B(\a[32] ), .Y(new_n4770_));
  XOR2X1   g04514(.A(new_n4770_), .B(new_n4766_), .Y(new_n4771_));
  INVX1    g04515(.A(new_n4555_), .Y(new_n4772_));
  AND2X1   g04516(.A(new_n4597_), .B(new_n4772_), .Y(new_n4773_));
  XOR2X1   g04517(.A(new_n4597_), .B(new_n4772_), .Y(new_n4774_));
  AOI21X1  g04518(.A0(new_n4774_), .A1(new_n4551_), .B0(new_n4773_), .Y(new_n4775_));
  XOR2X1   g04519(.A(new_n4775_), .B(new_n4771_), .Y(new_n4776_));
  AOI22X1  g04520(.A0(new_n2163_), .A1(\b[21] ), .B0(new_n2162_), .B1(\b[20] ), .Y(new_n4777_));
  OAI21X1  g04521(.A0(new_n2161_), .A1(new_n1300_), .B0(new_n4777_), .Y(new_n4778_));
  AOI21X1  g04522(.A0(new_n1907_), .A1(new_n1299_), .B0(new_n4778_), .Y(new_n4779_));
  XOR2X1   g04523(.A(new_n4779_), .B(\a[29] ), .Y(new_n4780_));
  XOR2X1   g04524(.A(new_n4780_), .B(new_n4776_), .Y(new_n4781_));
  OR2X1    g04525(.A(new_n4603_), .B(new_n4599_), .Y(new_n4782_));
  XOR2X1   g04526(.A(new_n4774_), .B(new_n4551_), .Y(new_n4783_));
  XOR2X1   g04527(.A(new_n4603_), .B(new_n4783_), .Y(new_n4784_));
  OAI21X1  g04528(.A0(new_n4606_), .A1(new_n4784_), .B0(new_n4782_), .Y(new_n4785_));
  XOR2X1   g04529(.A(new_n4785_), .B(new_n4781_), .Y(new_n4786_));
  AOI22X1  g04530(.A0(new_n1814_), .A1(\b[24] ), .B0(new_n1813_), .B1(\b[23] ), .Y(new_n4787_));
  OAI21X1  g04531(.A0(new_n1812_), .A1(new_n1479_), .B0(new_n4787_), .Y(new_n4788_));
  AOI21X1  g04532(.A0(new_n1617_), .A1(new_n1572_), .B0(new_n4788_), .Y(new_n4789_));
  XOR2X1   g04533(.A(new_n4789_), .B(\a[26] ), .Y(new_n4790_));
  XOR2X1   g04534(.A(new_n4790_), .B(new_n4786_), .Y(new_n4791_));
  XOR2X1   g04535(.A(new_n4791_), .B(new_n4616_), .Y(new_n4792_));
  AOI22X1  g04536(.A0(new_n1526_), .A1(\b[27] ), .B0(new_n1525_), .B1(\b[26] ), .Y(new_n4793_));
  OAI21X1  g04537(.A0(new_n1524_), .A1(new_n1880_), .B0(new_n4793_), .Y(new_n4794_));
  AOI21X1  g04538(.A0(new_n1879_), .A1(new_n1347_), .B0(new_n4794_), .Y(new_n4795_));
  XOR2X1   g04539(.A(new_n4795_), .B(\a[23] ), .Y(new_n4796_));
  XOR2X1   g04540(.A(new_n4796_), .B(new_n4792_), .Y(new_n4797_));
  INVX1    g04541(.A(new_n4797_), .Y(new_n4798_));
  XOR2X1   g04542(.A(new_n4798_), .B(new_n4713_), .Y(new_n4799_));
  AOI22X1  g04543(.A0(new_n1263_), .A1(\b[30] ), .B0(new_n1262_), .B1(\b[29] ), .Y(new_n4800_));
  OAI21X1  g04544(.A0(new_n1261_), .A1(new_n2231_), .B0(new_n4800_), .Y(new_n4801_));
  AOI21X1  g04545(.A0(new_n2230_), .A1(new_n1075_), .B0(new_n4801_), .Y(new_n4802_));
  XOR2X1   g04546(.A(new_n4802_), .B(\a[20] ), .Y(new_n4803_));
  XOR2X1   g04547(.A(new_n4803_), .B(new_n4799_), .Y(new_n4804_));
  XOR2X1   g04548(.A(new_n4804_), .B(new_n4710_), .Y(new_n4805_));
  AOI22X1  g04549(.A0(new_n1017_), .A1(\b[33] ), .B0(new_n1016_), .B1(\b[32] ), .Y(new_n4806_));
  OAI21X1  g04550(.A0(new_n1015_), .A1(new_n2615_), .B0(new_n4806_), .Y(new_n4807_));
  AOI21X1  g04551(.A0(new_n2614_), .A1(new_n882_), .B0(new_n4807_), .Y(new_n4808_));
  XOR2X1   g04552(.A(new_n4808_), .B(\a[17] ), .Y(new_n4809_));
  XOR2X1   g04553(.A(new_n4809_), .B(new_n4805_), .Y(new_n4810_));
  XOR2X1   g04554(.A(new_n4810_), .B(new_n4707_), .Y(new_n4811_));
  AOI22X1  g04555(.A0(new_n818_), .A1(\b[36] ), .B0(new_n817_), .B1(\b[35] ), .Y(new_n4812_));
  OAI21X1  g04556(.A0(new_n816_), .A1(new_n2890_), .B0(new_n4812_), .Y(new_n4813_));
  AOI21X1  g04557(.A0(new_n3015_), .A1(new_n668_), .B0(new_n4813_), .Y(new_n4814_));
  XOR2X1   g04558(.A(new_n4814_), .B(\a[14] ), .Y(new_n4815_));
  XOR2X1   g04559(.A(new_n4815_), .B(new_n4811_), .Y(new_n4816_));
  XOR2X1   g04560(.A(new_n4816_), .B(new_n4705_), .Y(new_n4817_));
  AOI22X1  g04561(.A0(new_n603_), .A1(\b[39] ), .B0(new_n602_), .B1(\b[38] ), .Y(new_n4818_));
  OAI21X1  g04562(.A0(new_n601_), .A1(new_n3413_), .B0(new_n4818_), .Y(new_n4819_));
  AOI21X1  g04563(.A0(new_n3412_), .A1(new_n518_), .B0(new_n4819_), .Y(new_n4820_));
  XOR2X1   g04564(.A(new_n4820_), .B(\a[11] ), .Y(new_n4821_));
  XOR2X1   g04565(.A(new_n4821_), .B(new_n4817_), .Y(new_n4822_));
  NOR2X1   g04566(.A(new_n4643_), .B(new_n4639_), .Y(new_n4823_));
  OR2X1    g04567(.A(new_n4470_), .B(new_n4466_), .Y(new_n4824_));
  XOR2X1   g04568(.A(new_n4523_), .B(new_n4347_), .Y(new_n4825_));
  XOR2X1   g04569(.A(new_n4458_), .B(new_n4825_), .Y(new_n4826_));
  XOR2X1   g04570(.A(new_n4465_), .B(new_n4826_), .Y(new_n4827_));
  XOR2X1   g04571(.A(new_n4470_), .B(new_n4827_), .Y(new_n4828_));
  OAI21X1  g04572(.A0(new_n4475_), .A1(new_n4828_), .B0(new_n4824_), .Y(new_n4829_));
  AOI21X1  g04573(.A0(new_n4829_), .A1(new_n4644_), .B0(new_n4823_), .Y(new_n4830_));
  XOR2X1   g04574(.A(new_n4830_), .B(new_n4822_), .Y(new_n4831_));
  AOI22X1  g04575(.A0(new_n469_), .A1(\b[42] ), .B0(new_n468_), .B1(\b[41] ), .Y(new_n4832_));
  OAI21X1  g04576(.A0(new_n467_), .A1(new_n3720_), .B0(new_n4832_), .Y(new_n4833_));
  AOI21X1  g04577(.A0(new_n3860_), .A1(new_n404_), .B0(new_n4833_), .Y(new_n4834_));
  XOR2X1   g04578(.A(new_n4834_), .B(\a[8] ), .Y(new_n4835_));
  XOR2X1   g04579(.A(new_n4835_), .B(new_n4831_), .Y(new_n4836_));
  XOR2X1   g04580(.A(new_n4836_), .B(new_n4661_), .Y(new_n4837_));
  AOI22X1  g04581(.A0(new_n369_), .A1(\b[45] ), .B0(new_n368_), .B1(\b[44] ), .Y(new_n4838_));
  OAI21X1  g04582(.A0(new_n367_), .A1(new_n4339_), .B0(new_n4838_), .Y(new_n4839_));
  AOI21X1  g04583(.A0(new_n4338_), .A1(new_n308_), .B0(new_n4839_), .Y(new_n4840_));
  XOR2X1   g04584(.A(new_n4840_), .B(\a[5] ), .Y(new_n4841_));
  XOR2X1   g04585(.A(new_n4841_), .B(new_n4837_), .Y(new_n4842_));
  XOR2X1   g04586(.A(new_n4842_), .B(new_n4699_), .Y(new_n4843_));
  XOR2X1   g04587(.A(new_n4843_), .B(new_n4697_), .Y(new_n4844_));
  XOR2X1   g04588(.A(new_n4844_), .B(new_n4688_), .Y(\f[48] ));
  INVX1    g04589(.A(new_n4697_), .Y(new_n4846_));
  AND2X1   g04590(.A(new_n4843_), .B(new_n4846_), .Y(new_n4847_));
  AOI21X1  g04591(.A0(new_n4687_), .A1(new_n4686_), .B0(new_n4844_), .Y(new_n4848_));
  OR2X1    g04592(.A(new_n4848_), .B(new_n4847_), .Y(new_n4849_));
  NOR2X1   g04593(.A(new_n4796_), .B(new_n4792_), .Y(new_n4850_));
  AOI21X1  g04594(.A0(new_n4712_), .A1(new_n4711_), .B0(new_n4798_), .Y(new_n4851_));
  NOR2X1   g04595(.A(new_n4851_), .B(new_n4850_), .Y(new_n4852_));
  AOI22X1  g04596(.A0(new_n1526_), .A1(\b[28] ), .B0(new_n1525_), .B1(\b[27] ), .Y(new_n4853_));
  OAI21X1  g04597(.A0(new_n1524_), .A1(new_n1877_), .B0(new_n4853_), .Y(new_n4854_));
  AOI21X1  g04598(.A0(new_n2004_), .A1(new_n1347_), .B0(new_n4854_), .Y(new_n4855_));
  XOR2X1   g04599(.A(new_n4855_), .B(\a[23] ), .Y(new_n4856_));
  INVX1    g04600(.A(new_n4856_), .Y(new_n4857_));
  INVX1    g04601(.A(new_n4729_), .Y(new_n4858_));
  AND2X1   g04602(.A(new_n4762_), .B(new_n4858_), .Y(new_n4859_));
  AOI21X1  g04603(.A0(new_n4724_), .A1(new_n4722_), .B0(new_n4763_), .Y(new_n4860_));
  NOR2X1   g04604(.A(new_n4860_), .B(new_n4859_), .Y(new_n4861_));
  NOR2X1   g04605(.A(new_n4759_), .B(new_n4755_), .Y(new_n4862_));
  INVX1    g04606(.A(new_n4862_), .Y(new_n4863_));
  OAI21X1  g04607(.A0(new_n4761_), .A1(new_n4733_), .B0(new_n4863_), .Y(new_n4864_));
  OR4X1    g04608(.A(new_n4736_), .B(new_n4575_), .C(new_n4383_), .D(new_n4373_), .Y(new_n4865_));
  OAI21X1  g04609(.A0(new_n4744_), .A1(new_n4738_), .B0(new_n4865_), .Y(new_n4866_));
  AND2X1   g04610(.A(new_n4375_), .B(new_n323_), .Y(new_n4867_));
  NOR3X1   g04611(.A(new_n4739_), .B(new_n4379_), .C(new_n277_), .Y(new_n4868_));
  OAI22X1  g04612(.A0(new_n4380_), .A1(new_n325_), .B0(new_n4378_), .B1(new_n297_), .Y(new_n4869_));
  NOR3X1   g04613(.A(new_n4869_), .B(new_n4868_), .C(new_n4867_), .Y(new_n4870_));
  XOR2X1   g04614(.A(new_n4870_), .B(new_n4568_), .Y(new_n4871_));
  OAI21X1  g04615(.A0(new_n4735_), .A1(new_n274_), .B0(\a[50] ), .Y(new_n4872_));
  INVX1    g04616(.A(\a[50] ), .Y(new_n4873_));
  XOR2X1   g04617(.A(new_n4873_), .B(\a[49] ), .Y(new_n4874_));
  NOR2X1   g04618(.A(new_n4874_), .B(new_n4735_), .Y(new_n4875_));
  XOR2X1   g04619(.A(\a[49] ), .B(\a[48] ), .Y(new_n4876_));
  AND2X1   g04620(.A(new_n4876_), .B(new_n4735_), .Y(new_n4877_));
  INVX1    g04621(.A(new_n4877_), .Y(new_n4878_));
  INVX1    g04622(.A(new_n4735_), .Y(new_n4879_));
  AND2X1   g04623(.A(new_n4874_), .B(new_n4879_), .Y(new_n4880_));
  INVX1    g04624(.A(new_n4880_), .Y(new_n4881_));
  OAI22X1  g04625(.A0(new_n4881_), .A1(new_n275_), .B0(new_n4878_), .B1(new_n274_), .Y(new_n4882_));
  AOI21X1  g04626(.A0(new_n4875_), .A1(new_n263_), .B0(new_n4882_), .Y(new_n4883_));
  XOR2X1   g04627(.A(new_n4883_), .B(\a[50] ), .Y(new_n4884_));
  XOR2X1   g04628(.A(new_n4884_), .B(new_n4872_), .Y(new_n4885_));
  XOR2X1   g04629(.A(new_n4885_), .B(new_n4871_), .Y(new_n4886_));
  XOR2X1   g04630(.A(new_n4886_), .B(new_n4866_), .Y(new_n4887_));
  AOI22X1  g04631(.A0(new_n4095_), .A1(\b[7] ), .B0(new_n4094_), .B1(\b[6] ), .Y(new_n4888_));
  OAI21X1  g04632(.A0(new_n4233_), .A1(new_n395_), .B0(new_n4888_), .Y(new_n4889_));
  AOI21X1  g04633(.A0(new_n3901_), .A1(new_n394_), .B0(new_n4889_), .Y(new_n4890_));
  XOR2X1   g04634(.A(new_n4890_), .B(\a[44] ), .Y(new_n4891_));
  XOR2X1   g04635(.A(new_n4891_), .B(new_n4887_), .Y(new_n4892_));
  INVX1    g04636(.A(new_n4749_), .Y(new_n4893_));
  NOR2X1   g04637(.A(new_n4753_), .B(new_n4750_), .Y(new_n4894_));
  AOI21X1  g04638(.A0(new_n4893_), .A1(new_n4745_), .B0(new_n4894_), .Y(new_n4895_));
  XOR2X1   g04639(.A(new_n4895_), .B(new_n4892_), .Y(new_n4896_));
  INVX1    g04640(.A(new_n4896_), .Y(new_n4897_));
  AOI22X1  g04641(.A0(new_n3652_), .A1(\b[10] ), .B0(new_n3651_), .B1(\b[9] ), .Y(new_n4898_));
  OAI21X1  g04642(.A0(new_n3778_), .A1(new_n489_), .B0(new_n4898_), .Y(new_n4899_));
  AOI21X1  g04643(.A0(new_n3480_), .A1(new_n543_), .B0(new_n4899_), .Y(new_n4900_));
  XOR2X1   g04644(.A(new_n4900_), .B(\a[41] ), .Y(new_n4901_));
  NAND2X1  g04645(.A(new_n4901_), .B(new_n4897_), .Y(new_n4902_));
  XOR2X1   g04646(.A(new_n4901_), .B(new_n4897_), .Y(new_n4903_));
  INVX1    g04647(.A(new_n4903_), .Y(new_n4904_));
  NOR2X1   g04648(.A(new_n4901_), .B(new_n4897_), .Y(new_n4905_));
  AOI21X1  g04649(.A0(new_n4902_), .A1(new_n4864_), .B0(new_n4905_), .Y(new_n4906_));
  AOI22X1  g04650(.A0(new_n4906_), .A1(new_n4902_), .B0(new_n4904_), .B1(new_n4864_), .Y(new_n4907_));
  AOI22X1  g04651(.A0(new_n3204_), .A1(\b[13] ), .B0(new_n3203_), .B1(\b[12] ), .Y(new_n4908_));
  OAI21X1  g04652(.A0(new_n3321_), .A1(new_n716_), .B0(new_n4908_), .Y(new_n4909_));
  AOI21X1  g04653(.A0(new_n3080_), .A1(new_n715_), .B0(new_n4909_), .Y(new_n4910_));
  XOR2X1   g04654(.A(new_n4910_), .B(\a[38] ), .Y(new_n4911_));
  XOR2X1   g04655(.A(new_n4911_), .B(new_n4907_), .Y(new_n4912_));
  XOR2X1   g04656(.A(new_n4912_), .B(new_n4861_), .Y(new_n4913_));
  AOI22X1  g04657(.A0(new_n2813_), .A1(\b[16] ), .B0(new_n2812_), .B1(\b[15] ), .Y(new_n4914_));
  OAI21X1  g04658(.A0(new_n2946_), .A1(new_n792_), .B0(new_n4914_), .Y(new_n4915_));
  AOI21X1  g04659(.A0(new_n2652_), .A1(new_n842_), .B0(new_n4915_), .Y(new_n4916_));
  XOR2X1   g04660(.A(new_n4916_), .B(\a[35] ), .Y(new_n4917_));
  XOR2X1   g04661(.A(new_n4917_), .B(new_n4913_), .Y(new_n4918_));
  AND2X1   g04662(.A(new_n4764_), .B(new_n4720_), .Y(new_n4919_));
  AOI21X1  g04663(.A0(new_n4765_), .A1(new_n4715_), .B0(new_n4919_), .Y(new_n4920_));
  XOR2X1   g04664(.A(new_n4920_), .B(new_n4918_), .Y(new_n4921_));
  AOI22X1  g04665(.A0(new_n2545_), .A1(\b[19] ), .B0(new_n2544_), .B1(\b[18] ), .Y(new_n4922_));
  OAI21X1  g04666(.A0(new_n2543_), .A1(new_n1118_), .B0(new_n4922_), .Y(new_n4923_));
  AOI21X1  g04667(.A0(new_n2260_), .A1(new_n1117_), .B0(new_n4923_), .Y(new_n4924_));
  XOR2X1   g04668(.A(new_n4924_), .B(\a[32] ), .Y(new_n4925_));
  XOR2X1   g04669(.A(new_n4925_), .B(new_n4921_), .Y(new_n4926_));
  INVX1    g04670(.A(new_n4770_), .Y(new_n4927_));
  NAND2X1  g04671(.A(new_n4927_), .B(new_n4766_), .Y(new_n4928_));
  OAI21X1  g04672(.A0(new_n4775_), .A1(new_n4771_), .B0(new_n4928_), .Y(new_n4929_));
  XOR2X1   g04673(.A(new_n4929_), .B(new_n4926_), .Y(new_n4930_));
  AOI22X1  g04674(.A0(new_n2163_), .A1(\b[22] ), .B0(new_n2162_), .B1(\b[21] ), .Y(new_n4931_));
  OAI21X1  g04675(.A0(new_n2161_), .A1(new_n1297_), .B0(new_n4931_), .Y(new_n4932_));
  AOI21X1  g04676(.A0(new_n1907_), .A1(new_n1399_), .B0(new_n4932_), .Y(new_n4933_));
  XOR2X1   g04677(.A(new_n4933_), .B(\a[29] ), .Y(new_n4934_));
  XOR2X1   g04678(.A(new_n4934_), .B(new_n4930_), .Y(new_n4935_));
  XOR2X1   g04679(.A(new_n4927_), .B(new_n4766_), .Y(new_n4936_));
  XOR2X1   g04680(.A(new_n4775_), .B(new_n4936_), .Y(new_n4937_));
  NOR2X1   g04681(.A(new_n4780_), .B(new_n4937_), .Y(new_n4938_));
  XOR2X1   g04682(.A(new_n4780_), .B(new_n4937_), .Y(new_n4939_));
  AOI21X1  g04683(.A0(new_n4785_), .A1(new_n4939_), .B0(new_n4938_), .Y(new_n4940_));
  XOR2X1   g04684(.A(new_n4940_), .B(new_n4935_), .Y(new_n4941_));
  AOI22X1  g04685(.A0(new_n1814_), .A1(\b[25] ), .B0(new_n1813_), .B1(\b[24] ), .Y(new_n4942_));
  OAI21X1  g04686(.A0(new_n1812_), .A1(new_n1591_), .B0(new_n4942_), .Y(new_n4943_));
  AOI21X1  g04687(.A0(new_n1617_), .A1(new_n1590_), .B0(new_n4943_), .Y(new_n4944_));
  XOR2X1   g04688(.A(new_n4944_), .B(\a[26] ), .Y(new_n4945_));
  XOR2X1   g04689(.A(new_n4945_), .B(new_n4941_), .Y(new_n4946_));
  NOR2X1   g04690(.A(new_n4790_), .B(new_n4786_), .Y(new_n4947_));
  INVX1    g04691(.A(new_n4947_), .Y(new_n4948_));
  OR2X1    g04692(.A(new_n4436_), .B(new_n4434_), .Y(new_n4949_));
  AOI21X1  g04693(.A0(new_n4949_), .A1(new_n4548_), .B0(new_n4614_), .Y(new_n4950_));
  OAI21X1  g04694(.A0(new_n4950_), .A1(new_n4615_), .B0(new_n4791_), .Y(new_n4951_));
  AND2X1   g04695(.A(new_n4951_), .B(new_n4948_), .Y(new_n4952_));
  XOR2X1   g04696(.A(new_n4952_), .B(new_n4946_), .Y(new_n4953_));
  XOR2X1   g04697(.A(new_n4953_), .B(new_n4857_), .Y(new_n4954_));
  XOR2X1   g04698(.A(new_n4954_), .B(new_n4852_), .Y(new_n4955_));
  AOI22X1  g04699(.A0(new_n1263_), .A1(\b[31] ), .B0(new_n1262_), .B1(\b[30] ), .Y(new_n4956_));
  OAI21X1  g04700(.A0(new_n1261_), .A1(new_n2359_), .B0(new_n4956_), .Y(new_n4957_));
  AOI21X1  g04701(.A0(new_n2358_), .A1(new_n1075_), .B0(new_n4957_), .Y(new_n4958_));
  XOR2X1   g04702(.A(new_n4958_), .B(\a[20] ), .Y(new_n4959_));
  INVX1    g04703(.A(new_n4959_), .Y(new_n4960_));
  XOR2X1   g04704(.A(new_n4960_), .B(new_n4955_), .Y(new_n4961_));
  XOR2X1   g04705(.A(new_n4797_), .B(new_n4713_), .Y(new_n4962_));
  NOR2X1   g04706(.A(new_n4803_), .B(new_n4962_), .Y(new_n4963_));
  XOR2X1   g04707(.A(new_n4803_), .B(new_n4962_), .Y(new_n4964_));
  AOI21X1  g04708(.A0(new_n4964_), .A1(new_n4710_), .B0(new_n4963_), .Y(new_n4965_));
  XOR2X1   g04709(.A(new_n4965_), .B(new_n4961_), .Y(new_n4966_));
  AOI22X1  g04710(.A0(new_n1017_), .A1(\b[34] ), .B0(new_n1016_), .B1(\b[33] ), .Y(new_n4967_));
  OAI21X1  g04711(.A0(new_n1015_), .A1(new_n2612_), .B0(new_n4967_), .Y(new_n4968_));
  AOI21X1  g04712(.A0(new_n2759_), .A1(new_n882_), .B0(new_n4968_), .Y(new_n4969_));
  XOR2X1   g04713(.A(new_n4969_), .B(\a[17] ), .Y(new_n4970_));
  XOR2X1   g04714(.A(new_n4970_), .B(new_n4966_), .Y(new_n4971_));
  OR2X1    g04715(.A(new_n4809_), .B(new_n4805_), .Y(new_n4972_));
  XOR2X1   g04716(.A(new_n4964_), .B(new_n4710_), .Y(new_n4973_));
  XOR2X1   g04717(.A(new_n4809_), .B(new_n4973_), .Y(new_n4974_));
  OAI21X1  g04718(.A0(new_n4974_), .A1(new_n4707_), .B0(new_n4972_), .Y(new_n4975_));
  XOR2X1   g04719(.A(new_n4975_), .B(new_n4971_), .Y(new_n4976_));
  AOI22X1  g04720(.A0(new_n818_), .A1(\b[37] ), .B0(new_n817_), .B1(\b[36] ), .Y(new_n4977_));
  OAI21X1  g04721(.A0(new_n816_), .A1(new_n3156_), .B0(new_n4977_), .Y(new_n4978_));
  AOI21X1  g04722(.A0(new_n3155_), .A1(new_n668_), .B0(new_n4978_), .Y(new_n4979_));
  XOR2X1   g04723(.A(new_n4979_), .B(\a[14] ), .Y(new_n4980_));
  XOR2X1   g04724(.A(new_n4980_), .B(new_n4976_), .Y(new_n4981_));
  NOR2X1   g04725(.A(new_n4815_), .B(new_n4811_), .Y(new_n4982_));
  AOI21X1  g04726(.A0(new_n4816_), .A1(new_n4705_), .B0(new_n4982_), .Y(new_n4983_));
  XOR2X1   g04727(.A(new_n4983_), .B(new_n4981_), .Y(new_n4984_));
  AOI22X1  g04728(.A0(new_n603_), .A1(\b[40] ), .B0(new_n602_), .B1(\b[39] ), .Y(new_n4985_));
  OAI21X1  g04729(.A0(new_n601_), .A1(new_n3575_), .B0(new_n4985_), .Y(new_n4986_));
  AOI21X1  g04730(.A0(new_n3574_), .A1(new_n518_), .B0(new_n4986_), .Y(new_n4987_));
  XOR2X1   g04731(.A(new_n4987_), .B(\a[11] ), .Y(new_n4988_));
  XOR2X1   g04732(.A(new_n4988_), .B(new_n4984_), .Y(new_n4989_));
  NOR2X1   g04733(.A(new_n4631_), .B(new_n4627_), .Y(new_n4990_));
  OR2X1    g04734(.A(new_n4458_), .B(new_n4454_), .Y(new_n4991_));
  OAI21X1  g04735(.A0(new_n4465_), .A1(new_n4826_), .B0(new_n4991_), .Y(new_n4992_));
  AOI21X1  g04736(.A0(new_n4992_), .A1(new_n4632_), .B0(new_n4990_), .Y(new_n4993_));
  XOR2X1   g04737(.A(new_n4816_), .B(new_n4993_), .Y(new_n4994_));
  NOR2X1   g04738(.A(new_n4821_), .B(new_n4994_), .Y(new_n4995_));
  XOR2X1   g04739(.A(new_n4821_), .B(new_n4994_), .Y(new_n4996_));
  OR2X1    g04740(.A(new_n4643_), .B(new_n4639_), .Y(new_n4997_));
  XOR2X1   g04741(.A(new_n4638_), .B(new_n4704_), .Y(new_n4998_));
  XOR2X1   g04742(.A(new_n4643_), .B(new_n4998_), .Y(new_n4999_));
  OAI21X1  g04743(.A0(new_n4649_), .A1(new_n4999_), .B0(new_n4997_), .Y(new_n5000_));
  AOI21X1  g04744(.A0(new_n5000_), .A1(new_n4996_), .B0(new_n4995_), .Y(new_n5001_));
  XOR2X1   g04745(.A(new_n5001_), .B(new_n4989_), .Y(new_n5002_));
  AOI22X1  g04746(.A0(new_n469_), .A1(\b[43] ), .B0(new_n468_), .B1(\b[42] ), .Y(new_n5003_));
  OAI21X1  g04747(.A0(new_n467_), .A1(new_n4015_), .B0(new_n5003_), .Y(new_n5004_));
  AOI21X1  g04748(.A0(new_n4014_), .A1(new_n404_), .B0(new_n5004_), .Y(new_n5005_));
  XOR2X1   g04749(.A(new_n5005_), .B(\a[8] ), .Y(new_n5006_));
  XOR2X1   g04750(.A(new_n5006_), .B(new_n5002_), .Y(new_n5007_));
  AND2X1   g04751(.A(new_n4654_), .B(new_n4650_), .Y(new_n5008_));
  OAI21X1  g04752(.A0(new_n5008_), .A1(new_n4493_), .B0(new_n4656_), .Y(new_n5009_));
  XOR2X1   g04753(.A(new_n4830_), .B(new_n4996_), .Y(new_n5010_));
  NOR2X1   g04754(.A(new_n4835_), .B(new_n5010_), .Y(new_n5011_));
  XOR2X1   g04755(.A(new_n4835_), .B(new_n5010_), .Y(new_n5012_));
  AOI21X1  g04756(.A0(new_n5012_), .A1(new_n5009_), .B0(new_n5011_), .Y(new_n5013_));
  XOR2X1   g04757(.A(new_n5013_), .B(new_n5007_), .Y(new_n5014_));
  AOI22X1  g04758(.A0(new_n369_), .A1(\b[46] ), .B0(new_n368_), .B1(\b[45] ), .Y(new_n5015_));
  OAI21X1  g04759(.A0(new_n367_), .A1(new_n4336_), .B0(new_n5015_), .Y(new_n5016_));
  AOI21X1  g04760(.A0(new_n4509_), .A1(new_n308_), .B0(new_n5016_), .Y(new_n5017_));
  XOR2X1   g04761(.A(new_n5017_), .B(\a[5] ), .Y(new_n5018_));
  XOR2X1   g04762(.A(new_n5018_), .B(new_n5014_), .Y(new_n5019_));
  NOR2X1   g04763(.A(new_n4498_), .B(new_n4494_), .Y(new_n5020_));
  OR2X1    g04764(.A(new_n4323_), .B(new_n4319_), .Y(new_n5021_));
  XOR2X1   g04765(.A(new_n4318_), .B(new_n4490_), .Y(new_n5022_));
  XOR2X1   g04766(.A(new_n4323_), .B(new_n5022_), .Y(new_n5023_));
  OAI21X1  g04767(.A0(new_n4332_), .A1(new_n5023_), .B0(new_n5021_), .Y(new_n5024_));
  AOI21X1  g04768(.A0(new_n5024_), .A1(new_n4680_), .B0(new_n5020_), .Y(new_n5025_));
  AND2X1   g04769(.A(new_n4666_), .B(new_n4662_), .Y(new_n5026_));
  OR2X1    g04770(.A(new_n4666_), .B(new_n4662_), .Y(new_n5027_));
  OAI21X1  g04771(.A0(new_n5026_), .A1(new_n5025_), .B0(new_n5027_), .Y(new_n5028_));
  XOR2X1   g04772(.A(new_n4836_), .B(new_n5009_), .Y(new_n5029_));
  NOR2X1   g04773(.A(new_n4841_), .B(new_n5029_), .Y(new_n5030_));
  XOR2X1   g04774(.A(new_n4841_), .B(new_n5029_), .Y(new_n5031_));
  AOI21X1  g04775(.A0(new_n5031_), .A1(new_n5028_), .B0(new_n5030_), .Y(new_n5032_));
  XOR2X1   g04776(.A(new_n5032_), .B(new_n5019_), .Y(new_n5033_));
  AND2X1   g04777(.A(\b[48] ), .B(\b[47] ), .Y(new_n5034_));
  AOI21X1  g04778(.A0(new_n4691_), .A1(new_n4690_), .B0(new_n5034_), .Y(new_n5035_));
  INVX1    g04779(.A(\b[48] ), .Y(new_n5036_));
  XOR2X1   g04780(.A(\b[49] ), .B(new_n5036_), .Y(new_n5037_));
  XOR2X1   g04781(.A(new_n5037_), .B(new_n5035_), .Y(new_n5038_));
  INVX1    g04782(.A(\b[47] ), .Y(new_n5039_));
  AOI22X1  g04783(.A0(new_n267_), .A1(\b[49] ), .B0(new_n266_), .B1(\b[48] ), .Y(new_n5040_));
  OAI21X1  g04784(.A0(new_n350_), .A1(new_n5039_), .B0(new_n5040_), .Y(new_n5041_));
  AOI21X1  g04785(.A0(new_n5038_), .A1(new_n318_), .B0(new_n5041_), .Y(new_n5042_));
  XOR2X1   g04786(.A(new_n5042_), .B(\a[2] ), .Y(new_n5043_));
  XOR2X1   g04787(.A(new_n5043_), .B(new_n5033_), .Y(new_n5044_));
  XOR2X1   g04788(.A(new_n5044_), .B(new_n4849_), .Y(\f[49] ));
  NOR2X1   g04789(.A(new_n5006_), .B(new_n5002_), .Y(new_n5046_));
  OR2X1    g04790(.A(new_n4835_), .B(new_n5010_), .Y(new_n5047_));
  OAI21X1  g04791(.A0(new_n4836_), .A1(new_n4661_), .B0(new_n5047_), .Y(new_n5048_));
  AOI21X1  g04792(.A0(new_n5048_), .A1(new_n5007_), .B0(new_n5046_), .Y(new_n5049_));
  OR2X1    g04793(.A(new_n4959_), .B(new_n4955_), .Y(new_n5050_));
  OAI21X1  g04794(.A0(new_n4965_), .A1(new_n4961_), .B0(new_n5050_), .Y(new_n5051_));
  AOI22X1  g04795(.A0(new_n1263_), .A1(\b[32] ), .B0(new_n1262_), .B1(\b[31] ), .Y(new_n5052_));
  OAI21X1  g04796(.A0(new_n1261_), .A1(new_n2356_), .B0(new_n5052_), .Y(new_n5053_));
  AOI21X1  g04797(.A0(new_n2495_), .A1(new_n1075_), .B0(new_n5053_), .Y(new_n5054_));
  XOR2X1   g04798(.A(new_n5054_), .B(\a[20] ), .Y(new_n5055_));
  INVX1    g04799(.A(new_n5055_), .Y(new_n5056_));
  NAND2X1  g04800(.A(new_n4953_), .B(new_n4857_), .Y(new_n5057_));
  OAI21X1  g04801(.A0(new_n4851_), .A1(new_n4850_), .B0(new_n4954_), .Y(new_n5058_));
  AND2X1   g04802(.A(new_n5058_), .B(new_n5057_), .Y(new_n5059_));
  AOI22X1  g04803(.A0(new_n1526_), .A1(\b[29] ), .B0(new_n1525_), .B1(\b[28] ), .Y(new_n5060_));
  OAI21X1  g04804(.A0(new_n1524_), .A1(new_n2126_), .B0(new_n5060_), .Y(new_n5061_));
  AOI21X1  g04805(.A0(new_n2125_), .A1(new_n1347_), .B0(new_n5061_), .Y(new_n5062_));
  XOR2X1   g04806(.A(new_n5062_), .B(\a[23] ), .Y(new_n5063_));
  XOR2X1   g04807(.A(new_n4944_), .B(new_n1621_), .Y(new_n5064_));
  AND2X1   g04808(.A(new_n5064_), .B(new_n4941_), .Y(new_n5065_));
  AOI21X1  g04809(.A0(new_n4951_), .A1(new_n4948_), .B0(new_n4946_), .Y(new_n5066_));
  OR2X1    g04810(.A(new_n5066_), .B(new_n5065_), .Y(new_n5067_));
  XOR2X1   g04811(.A(new_n4933_), .B(new_n1911_), .Y(new_n5068_));
  NAND2X1  g04812(.A(new_n5068_), .B(new_n4930_), .Y(new_n5069_));
  OAI21X1  g04813(.A0(new_n4940_), .A1(new_n4935_), .B0(new_n5069_), .Y(new_n5070_));
  OR2X1    g04814(.A(new_n4917_), .B(new_n4913_), .Y(new_n5071_));
  XOR2X1   g04815(.A(new_n4916_), .B(new_n2650_), .Y(new_n5072_));
  XOR2X1   g04816(.A(new_n5072_), .B(new_n4913_), .Y(new_n5073_));
  OAI21X1  g04817(.A0(new_n4920_), .A1(new_n5073_), .B0(new_n5071_), .Y(new_n5074_));
  AOI22X1  g04818(.A0(new_n2813_), .A1(\b[17] ), .B0(new_n2812_), .B1(\b[16] ), .Y(new_n5075_));
  OAI21X1  g04819(.A0(new_n2946_), .A1(new_n977_), .B0(new_n5075_), .Y(new_n5076_));
  AOI21X1  g04820(.A0(new_n2652_), .A1(new_n976_), .B0(new_n5076_), .Y(new_n5077_));
  XOR2X1   g04821(.A(new_n5077_), .B(\a[35] ), .Y(new_n5078_));
  OR2X1    g04822(.A(new_n4911_), .B(new_n4907_), .Y(new_n5079_));
  OAI21X1  g04823(.A0(new_n4860_), .A1(new_n4859_), .B0(new_n4912_), .Y(new_n5080_));
  AND2X1   g04824(.A(new_n5080_), .B(new_n5079_), .Y(new_n5081_));
  INVX1    g04825(.A(new_n4887_), .Y(new_n5082_));
  OR2X1    g04826(.A(new_n4895_), .B(new_n4892_), .Y(new_n5083_));
  OAI21X1  g04827(.A0(new_n4891_), .A1(new_n5082_), .B0(new_n5083_), .Y(new_n5084_));
  AOI22X1  g04828(.A0(new_n4095_), .A1(\b[8] ), .B0(new_n4094_), .B1(\b[7] ), .Y(new_n5085_));
  OAI21X1  g04829(.A0(new_n4233_), .A1(new_n392_), .B0(new_n5085_), .Y(new_n5086_));
  AOI21X1  g04830(.A0(new_n3901_), .A1(new_n454_), .B0(new_n5086_), .Y(new_n5087_));
  XOR2X1   g04831(.A(new_n5087_), .B(\a[44] ), .Y(new_n5088_));
  AND2X1   g04832(.A(new_n4885_), .B(new_n4871_), .Y(new_n5089_));
  AOI21X1  g04833(.A0(new_n4886_), .A1(new_n4866_), .B0(new_n5089_), .Y(new_n5090_));
  NAND3X1  g04834(.A(new_n4883_), .B(new_n4736_), .C(\a[50] ), .Y(new_n5091_));
  NAND2X1  g04835(.A(new_n4875_), .B(new_n341_), .Y(new_n5092_));
  OR4X1    g04836(.A(new_n4876_), .B(new_n4874_), .C(new_n4879_), .D(new_n274_), .Y(new_n5093_));
  AOI22X1  g04837(.A0(new_n4880_), .A1(\b[2] ), .B0(new_n4877_), .B1(\b[1] ), .Y(new_n5094_));
  NAND3X1  g04838(.A(new_n5094_), .B(new_n5093_), .C(new_n5092_), .Y(new_n5095_));
  XOR2X1   g04839(.A(new_n5095_), .B(new_n4873_), .Y(new_n5096_));
  XOR2X1   g04840(.A(new_n5096_), .B(new_n5091_), .Y(new_n5097_));
  AOI22X1  g04841(.A0(new_n4572_), .A1(\b[5] ), .B0(new_n4571_), .B1(\b[4] ), .Y(new_n5098_));
  OAI21X1  g04842(.A0(new_n4740_), .A1(new_n297_), .B0(new_n5098_), .Y(new_n5099_));
  AOI21X1  g04843(.A0(new_n4375_), .A1(new_n349_), .B0(new_n5099_), .Y(new_n5100_));
  XOR2X1   g04844(.A(new_n5100_), .B(\a[47] ), .Y(new_n5101_));
  XOR2X1   g04845(.A(new_n5101_), .B(new_n5097_), .Y(new_n5102_));
  XOR2X1   g04846(.A(new_n5102_), .B(new_n5090_), .Y(new_n5103_));
  XOR2X1   g04847(.A(new_n5103_), .B(new_n5088_), .Y(new_n5104_));
  XOR2X1   g04848(.A(new_n5104_), .B(new_n5084_), .Y(new_n5105_));
  AOI22X1  g04849(.A0(new_n3652_), .A1(\b[11] ), .B0(new_n3651_), .B1(\b[10] ), .Y(new_n5106_));
  OAI21X1  g04850(.A0(new_n3778_), .A1(new_n590_), .B0(new_n5106_), .Y(new_n5107_));
  AOI21X1  g04851(.A0(new_n3480_), .A1(new_n589_), .B0(new_n5107_), .Y(new_n5108_));
  XOR2X1   g04852(.A(new_n5108_), .B(\a[41] ), .Y(new_n5109_));
  XOR2X1   g04853(.A(new_n5109_), .B(new_n5105_), .Y(new_n5110_));
  XOR2X1   g04854(.A(new_n5110_), .B(new_n4906_), .Y(new_n5111_));
  AOI22X1  g04855(.A0(new_n3204_), .A1(\b[14] ), .B0(new_n3203_), .B1(\b[13] ), .Y(new_n5112_));
  OAI21X1  g04856(.A0(new_n3321_), .A1(new_n713_), .B0(new_n5112_), .Y(new_n5113_));
  AOI21X1  g04857(.A0(new_n3080_), .A1(new_n734_), .B0(new_n5113_), .Y(new_n5114_));
  XOR2X1   g04858(.A(new_n5114_), .B(\a[38] ), .Y(new_n5115_));
  XOR2X1   g04859(.A(new_n5115_), .B(new_n5111_), .Y(new_n5116_));
  INVX1    g04860(.A(new_n5116_), .Y(new_n5117_));
  XOR2X1   g04861(.A(new_n5117_), .B(new_n5081_), .Y(new_n5118_));
  XOR2X1   g04862(.A(new_n5118_), .B(new_n5078_), .Y(new_n5119_));
  XOR2X1   g04863(.A(new_n5119_), .B(new_n5074_), .Y(new_n5120_));
  AOI22X1  g04864(.A0(new_n2545_), .A1(\b[20] ), .B0(new_n2544_), .B1(\b[19] ), .Y(new_n5121_));
  OAI21X1  g04865(.A0(new_n2543_), .A1(new_n1115_), .B0(new_n5121_), .Y(new_n5122_));
  AOI21X1  g04866(.A0(new_n2260_), .A1(new_n1217_), .B0(new_n5122_), .Y(new_n5123_));
  XOR2X1   g04867(.A(new_n5123_), .B(\a[32] ), .Y(new_n5124_));
  XOR2X1   g04868(.A(new_n5124_), .B(new_n5120_), .Y(new_n5125_));
  NOR2X1   g04869(.A(new_n4925_), .B(new_n4921_), .Y(new_n5126_));
  AOI21X1  g04870(.A0(new_n4929_), .A1(new_n4926_), .B0(new_n5126_), .Y(new_n5127_));
  XOR2X1   g04871(.A(new_n5127_), .B(new_n5125_), .Y(new_n5128_));
  AOI22X1  g04872(.A0(new_n2163_), .A1(\b[23] ), .B0(new_n2162_), .B1(\b[22] ), .Y(new_n5129_));
  OAI21X1  g04873(.A0(new_n2161_), .A1(new_n1482_), .B0(new_n5129_), .Y(new_n5130_));
  AOI21X1  g04874(.A0(new_n1907_), .A1(new_n1481_), .B0(new_n5130_), .Y(new_n5131_));
  XOR2X1   g04875(.A(new_n5131_), .B(\a[29] ), .Y(new_n5132_));
  NAND2X1  g04876(.A(new_n5132_), .B(new_n5128_), .Y(new_n5133_));
  XOR2X1   g04877(.A(new_n5132_), .B(new_n5128_), .Y(new_n5134_));
  INVX1    g04878(.A(new_n5134_), .Y(new_n5135_));
  NOR2X1   g04879(.A(new_n5132_), .B(new_n5128_), .Y(new_n5136_));
  AOI21X1  g04880(.A0(new_n5133_), .A1(new_n5070_), .B0(new_n5136_), .Y(new_n5137_));
  AOI22X1  g04881(.A0(new_n5137_), .A1(new_n5133_), .B0(new_n5135_), .B1(new_n5070_), .Y(new_n5138_));
  AOI22X1  g04882(.A0(new_n1814_), .A1(\b[26] ), .B0(new_n1813_), .B1(\b[25] ), .Y(new_n5139_));
  OAI21X1  g04883(.A0(new_n1812_), .A1(new_n1588_), .B0(new_n5139_), .Y(new_n5140_));
  AOI21X1  g04884(.A0(new_n1783_), .A1(new_n1617_), .B0(new_n5140_), .Y(new_n5141_));
  XOR2X1   g04885(.A(new_n5141_), .B(\a[26] ), .Y(new_n5142_));
  XOR2X1   g04886(.A(new_n5142_), .B(new_n5138_), .Y(new_n5143_));
  XOR2X1   g04887(.A(new_n5143_), .B(new_n5067_), .Y(new_n5144_));
  XOR2X1   g04888(.A(new_n5144_), .B(new_n5063_), .Y(new_n5145_));
  XOR2X1   g04889(.A(new_n5145_), .B(new_n5059_), .Y(new_n5146_));
  XOR2X1   g04890(.A(new_n5146_), .B(new_n5056_), .Y(new_n5147_));
  XOR2X1   g04891(.A(new_n5147_), .B(new_n5051_), .Y(new_n5148_));
  AOI22X1  g04892(.A0(new_n1017_), .A1(\b[35] ), .B0(new_n1016_), .B1(\b[34] ), .Y(new_n5149_));
  OAI21X1  g04893(.A0(new_n1015_), .A1(new_n2893_), .B0(new_n5149_), .Y(new_n5150_));
  AOI21X1  g04894(.A0(new_n2892_), .A1(new_n882_), .B0(new_n5150_), .Y(new_n5151_));
  XOR2X1   g04895(.A(new_n5151_), .B(\a[17] ), .Y(new_n5152_));
  INVX1    g04896(.A(new_n5152_), .Y(new_n5153_));
  XOR2X1   g04897(.A(new_n5153_), .B(new_n5148_), .Y(new_n5154_));
  XOR2X1   g04898(.A(new_n4959_), .B(new_n4955_), .Y(new_n5155_));
  XOR2X1   g04899(.A(new_n4965_), .B(new_n5155_), .Y(new_n5156_));
  NOR2X1   g04900(.A(new_n4970_), .B(new_n5156_), .Y(new_n5157_));
  XOR2X1   g04901(.A(new_n4970_), .B(new_n5156_), .Y(new_n5158_));
  AOI21X1  g04902(.A0(new_n4975_), .A1(new_n5158_), .B0(new_n5157_), .Y(new_n5159_));
  XOR2X1   g04903(.A(new_n5159_), .B(new_n5154_), .Y(new_n5160_));
  AOI22X1  g04904(.A0(new_n818_), .A1(\b[38] ), .B0(new_n817_), .B1(\b[37] ), .Y(new_n5161_));
  OAI21X1  g04905(.A0(new_n816_), .A1(new_n3276_), .B0(new_n5161_), .Y(new_n5162_));
  AOI21X1  g04906(.A0(new_n3275_), .A1(new_n668_), .B0(new_n5162_), .Y(new_n5163_));
  XOR2X1   g04907(.A(new_n5163_), .B(\a[14] ), .Y(new_n5164_));
  XOR2X1   g04908(.A(new_n5164_), .B(new_n5160_), .Y(new_n5165_));
  NOR2X1   g04909(.A(new_n4980_), .B(new_n4976_), .Y(new_n5166_));
  OR2X1    g04910(.A(new_n4815_), .B(new_n4811_), .Y(new_n5167_));
  AND2X1   g04911(.A(new_n4815_), .B(new_n4811_), .Y(new_n5168_));
  OAI21X1  g04912(.A0(new_n5168_), .A1(new_n4993_), .B0(new_n5167_), .Y(new_n5169_));
  AOI21X1  g04913(.A0(new_n5169_), .A1(new_n4981_), .B0(new_n5166_), .Y(new_n5170_));
  XOR2X1   g04914(.A(new_n5170_), .B(new_n5165_), .Y(new_n5171_));
  AOI22X1  g04915(.A0(new_n603_), .A1(\b[41] ), .B0(new_n602_), .B1(\b[40] ), .Y(new_n5172_));
  OAI21X1  g04916(.A0(new_n601_), .A1(new_n3723_), .B0(new_n5172_), .Y(new_n5173_));
  AOI21X1  g04917(.A0(new_n3722_), .A1(new_n518_), .B0(new_n5173_), .Y(new_n5174_));
  XOR2X1   g04918(.A(new_n5174_), .B(\a[11] ), .Y(new_n5175_));
  XOR2X1   g04919(.A(new_n5175_), .B(new_n5171_), .Y(new_n5176_));
  NOR2X1   g04920(.A(new_n4988_), .B(new_n4984_), .Y(new_n5177_));
  OR2X1    g04921(.A(new_n4821_), .B(new_n4994_), .Y(new_n5178_));
  OAI21X1  g04922(.A0(new_n4830_), .A1(new_n4822_), .B0(new_n5178_), .Y(new_n5179_));
  AOI21X1  g04923(.A0(new_n5179_), .A1(new_n4989_), .B0(new_n5177_), .Y(new_n5180_));
  XOR2X1   g04924(.A(new_n5180_), .B(new_n5176_), .Y(new_n5181_));
  AOI22X1  g04925(.A0(new_n469_), .A1(\b[44] ), .B0(new_n468_), .B1(\b[43] ), .Y(new_n5182_));
  OAI21X1  g04926(.A0(new_n467_), .A1(new_n4012_), .B0(new_n5182_), .Y(new_n5183_));
  AOI21X1  g04927(.A0(new_n4178_), .A1(new_n404_), .B0(new_n5183_), .Y(new_n5184_));
  XOR2X1   g04928(.A(new_n5184_), .B(\a[8] ), .Y(new_n5185_));
  AND2X1   g04929(.A(new_n5185_), .B(new_n5181_), .Y(new_n5186_));
  XOR2X1   g04930(.A(new_n5185_), .B(new_n5181_), .Y(new_n5187_));
  OR2X1    g04931(.A(new_n5185_), .B(new_n5181_), .Y(new_n5188_));
  OAI21X1  g04932(.A0(new_n5186_), .A1(new_n5049_), .B0(new_n5188_), .Y(new_n5189_));
  OAI22X1  g04933(.A0(new_n5189_), .A1(new_n5186_), .B0(new_n5187_), .B1(new_n5049_), .Y(new_n5190_));
  AOI22X1  g04934(.A0(new_n369_), .A1(\b[47] ), .B0(new_n368_), .B1(\b[46] ), .Y(new_n5191_));
  OAI21X1  g04935(.A0(new_n367_), .A1(new_n4674_), .B0(new_n5191_), .Y(new_n5192_));
  AOI21X1  g04936(.A0(new_n4673_), .A1(new_n308_), .B0(new_n5192_), .Y(new_n5193_));
  XOR2X1   g04937(.A(new_n5193_), .B(\a[5] ), .Y(new_n5194_));
  XOR2X1   g04938(.A(new_n5194_), .B(new_n5190_), .Y(new_n5195_));
  NOR2X1   g04939(.A(new_n5018_), .B(new_n5014_), .Y(new_n5196_));
  OR2X1    g04940(.A(new_n4841_), .B(new_n5029_), .Y(new_n5197_));
  OAI21X1  g04941(.A0(new_n4842_), .A1(new_n4699_), .B0(new_n5197_), .Y(new_n5198_));
  AOI21X1  g04942(.A0(new_n5198_), .A1(new_n5019_), .B0(new_n5196_), .Y(new_n5199_));
  XOR2X1   g04943(.A(new_n5199_), .B(new_n5195_), .Y(new_n5200_));
  NAND2X1  g04944(.A(\b[49] ), .B(\b[48] ), .Y(new_n5201_));
  OAI21X1  g04945(.A0(new_n5037_), .A1(new_n5035_), .B0(new_n5201_), .Y(new_n5202_));
  XOR2X1   g04946(.A(\b[50] ), .B(\b[49] ), .Y(new_n5203_));
  XOR2X1   g04947(.A(new_n5203_), .B(new_n5202_), .Y(new_n5204_));
  AOI22X1  g04948(.A0(new_n267_), .A1(\b[50] ), .B0(new_n266_), .B1(\b[49] ), .Y(new_n5205_));
  OAI21X1  g04949(.A0(new_n350_), .A1(new_n5036_), .B0(new_n5205_), .Y(new_n5206_));
  AOI21X1  g04950(.A0(new_n5204_), .A1(new_n318_), .B0(new_n5206_), .Y(new_n5207_));
  XOR2X1   g04951(.A(new_n5207_), .B(\a[2] ), .Y(new_n5208_));
  XOR2X1   g04952(.A(new_n5208_), .B(new_n5200_), .Y(new_n5209_));
  OR2X1    g04953(.A(new_n5043_), .B(new_n5033_), .Y(new_n5210_));
  OAI21X1  g04954(.A0(new_n4848_), .A1(new_n4847_), .B0(new_n5044_), .Y(new_n5211_));
  AND2X1   g04955(.A(new_n5211_), .B(new_n5210_), .Y(new_n5212_));
  XOR2X1   g04956(.A(new_n5212_), .B(new_n5209_), .Y(\f[50] ));
  NAND2X1  g04957(.A(new_n5185_), .B(new_n5181_), .Y(new_n5214_));
  NOR2X1   g04958(.A(new_n5187_), .B(new_n5049_), .Y(new_n5215_));
  OR2X1    g04959(.A(new_n5006_), .B(new_n5002_), .Y(new_n5216_));
  XOR2X1   g04960(.A(new_n4975_), .B(new_n5158_), .Y(new_n5217_));
  XOR2X1   g04961(.A(new_n4980_), .B(new_n5217_), .Y(new_n5218_));
  XOR2X1   g04962(.A(new_n4983_), .B(new_n5218_), .Y(new_n5219_));
  XOR2X1   g04963(.A(new_n4988_), .B(new_n5219_), .Y(new_n5220_));
  XOR2X1   g04964(.A(new_n5001_), .B(new_n5220_), .Y(new_n5221_));
  XOR2X1   g04965(.A(new_n5006_), .B(new_n5221_), .Y(new_n5222_));
  OAI21X1  g04966(.A0(new_n5013_), .A1(new_n5222_), .B0(new_n5216_), .Y(new_n5223_));
  NOR2X1   g04967(.A(new_n5185_), .B(new_n5181_), .Y(new_n5224_));
  AOI21X1  g04968(.A0(new_n5214_), .A1(new_n5223_), .B0(new_n5224_), .Y(new_n5225_));
  AOI21X1  g04969(.A0(new_n5225_), .A1(new_n5214_), .B0(new_n5215_), .Y(new_n5226_));
  XOR2X1   g04970(.A(new_n5194_), .B(new_n5226_), .Y(new_n5227_));
  XOR2X1   g04971(.A(new_n5199_), .B(new_n5227_), .Y(new_n5228_));
  NOR2X1   g04972(.A(new_n5208_), .B(new_n5228_), .Y(new_n5229_));
  AOI21X1  g04973(.A0(new_n5211_), .A1(new_n5210_), .B0(new_n5209_), .Y(new_n5230_));
  OR2X1    g04974(.A(new_n5230_), .B(new_n5229_), .Y(new_n5231_));
  AND2X1   g04975(.A(\b[50] ), .B(\b[49] ), .Y(new_n5232_));
  AOI21X1  g04976(.A0(new_n5203_), .A1(new_n5202_), .B0(new_n5232_), .Y(new_n5233_));
  INVX1    g04977(.A(\b[50] ), .Y(new_n5234_));
  XOR2X1   g04978(.A(\b[51] ), .B(new_n5234_), .Y(new_n5235_));
  XOR2X1   g04979(.A(new_n5235_), .B(new_n5233_), .Y(new_n5236_));
  INVX1    g04980(.A(\b[49] ), .Y(new_n5237_));
  AOI22X1  g04981(.A0(new_n267_), .A1(\b[51] ), .B0(new_n266_), .B1(\b[50] ), .Y(new_n5238_));
  OAI21X1  g04982(.A0(new_n350_), .A1(new_n5237_), .B0(new_n5238_), .Y(new_n5239_));
  AOI21X1  g04983(.A0(new_n5236_), .A1(new_n318_), .B0(new_n5239_), .Y(new_n5240_));
  XOR2X1   g04984(.A(new_n5240_), .B(new_n257_), .Y(new_n5241_));
  OR2X1    g04985(.A(new_n5194_), .B(new_n5226_), .Y(new_n5242_));
  OAI21X1  g04986(.A0(new_n5199_), .A1(new_n5195_), .B0(new_n5242_), .Y(new_n5243_));
  NAND2X1  g04987(.A(new_n5153_), .B(new_n5148_), .Y(new_n5244_));
  XOR2X1   g04988(.A(new_n5152_), .B(new_n5148_), .Y(new_n5245_));
  OAI21X1  g04989(.A0(new_n5159_), .A1(new_n5245_), .B0(new_n5244_), .Y(new_n5246_));
  AND2X1   g04990(.A(new_n5146_), .B(new_n5056_), .Y(new_n5247_));
  AOI21X1  g04991(.A0(new_n5147_), .A1(new_n5051_), .B0(new_n5247_), .Y(new_n5248_));
  INVX1    g04992(.A(new_n5063_), .Y(new_n5249_));
  AND2X1   g04993(.A(new_n5144_), .B(new_n5249_), .Y(new_n5250_));
  AOI21X1  g04994(.A0(new_n5058_), .A1(new_n5057_), .B0(new_n5145_), .Y(new_n5251_));
  NOR2X1   g04995(.A(new_n5251_), .B(new_n5250_), .Y(new_n5252_));
  OR2X1    g04996(.A(new_n5142_), .B(new_n5138_), .Y(new_n5253_));
  NAND2X1  g04997(.A(new_n5143_), .B(new_n5067_), .Y(new_n5254_));
  AND2X1   g04998(.A(new_n5254_), .B(new_n5253_), .Y(new_n5255_));
  INVX1    g04999(.A(new_n5078_), .Y(new_n5256_));
  AND2X1   g05000(.A(new_n5118_), .B(new_n5256_), .Y(new_n5257_));
  XOR2X1   g05001(.A(new_n5118_), .B(new_n5256_), .Y(new_n5258_));
  AOI21X1  g05002(.A0(new_n5258_), .A1(new_n5074_), .B0(new_n5257_), .Y(new_n5259_));
  AOI22X1  g05003(.A0(new_n2813_), .A1(\b[18] ), .B0(new_n2812_), .B1(\b[17] ), .Y(new_n5260_));
  OAI21X1  g05004(.A0(new_n2946_), .A1(new_n974_), .B0(new_n5260_), .Y(new_n5261_));
  AOI21X1  g05005(.A0(new_n2652_), .A1(new_n1042_), .B0(new_n5261_), .Y(new_n5262_));
  XOR2X1   g05006(.A(new_n5262_), .B(\a[35] ), .Y(new_n5263_));
  NOR2X1   g05007(.A(new_n5115_), .B(new_n5111_), .Y(new_n5264_));
  AOI21X1  g05008(.A0(new_n5080_), .A1(new_n5079_), .B0(new_n5117_), .Y(new_n5265_));
  OR2X1    g05009(.A(new_n5265_), .B(new_n5264_), .Y(new_n5266_));
  AOI22X1  g05010(.A0(new_n3204_), .A1(\b[15] ), .B0(new_n3203_), .B1(\b[14] ), .Y(new_n5267_));
  OAI21X1  g05011(.A0(new_n3321_), .A1(new_n795_), .B0(new_n5267_), .Y(new_n5268_));
  AOI21X1  g05012(.A0(new_n3080_), .A1(new_n794_), .B0(new_n5268_), .Y(new_n5269_));
  XOR2X1   g05013(.A(new_n5269_), .B(\a[38] ), .Y(new_n5270_));
  INVX1    g05014(.A(new_n5270_), .Y(new_n5271_));
  NOR2X1   g05015(.A(new_n5109_), .B(new_n5105_), .Y(new_n5272_));
  INVX1    g05016(.A(new_n5272_), .Y(new_n5273_));
  AND2X1   g05017(.A(new_n4903_), .B(new_n4864_), .Y(new_n5274_));
  OAI21X1  g05018(.A0(new_n5274_), .A1(new_n4905_), .B0(new_n5110_), .Y(new_n5275_));
  AND2X1   g05019(.A(new_n5275_), .B(new_n5273_), .Y(new_n5276_));
  AOI22X1  g05020(.A0(new_n3652_), .A1(\b[12] ), .B0(new_n3651_), .B1(\b[11] ), .Y(new_n5277_));
  OAI21X1  g05021(.A0(new_n3778_), .A1(new_n587_), .B0(new_n5277_), .Y(new_n5278_));
  AOI21X1  g05022(.A0(new_n3480_), .A1(new_n635_), .B0(new_n5278_), .Y(new_n5279_));
  XOR2X1   g05023(.A(new_n5279_), .B(\a[41] ), .Y(new_n5280_));
  INVX1    g05024(.A(new_n5088_), .Y(new_n5281_));
  AND2X1   g05025(.A(new_n5103_), .B(new_n5281_), .Y(new_n5282_));
  INVX1    g05026(.A(new_n5104_), .Y(new_n5283_));
  AND2X1   g05027(.A(new_n5283_), .B(new_n5084_), .Y(new_n5284_));
  OR2X1    g05028(.A(new_n5284_), .B(new_n5282_), .Y(new_n5285_));
  OR2X1    g05029(.A(new_n5096_), .B(new_n5091_), .Y(new_n5286_));
  XOR2X1   g05030(.A(\a[51] ), .B(new_n4873_), .Y(new_n5287_));
  NOR2X1   g05031(.A(new_n5287_), .B(new_n274_), .Y(new_n5288_));
  XOR2X1   g05032(.A(new_n5288_), .B(new_n5286_), .Y(new_n5289_));
  OR2X1    g05033(.A(new_n4876_), .B(new_n4879_), .Y(new_n5290_));
  OR2X1    g05034(.A(new_n5290_), .B(new_n4874_), .Y(new_n5291_));
  AOI22X1  g05035(.A0(new_n4880_), .A1(\b[3] ), .B0(new_n4877_), .B1(\b[2] ), .Y(new_n5292_));
  OAI21X1  g05036(.A0(new_n5291_), .A1(new_n275_), .B0(new_n5292_), .Y(new_n5293_));
  AOI21X1  g05037(.A0(new_n4875_), .A1(new_n366_), .B0(new_n5293_), .Y(new_n5294_));
  XOR2X1   g05038(.A(new_n5294_), .B(\a[50] ), .Y(new_n5295_));
  XOR2X1   g05039(.A(new_n5295_), .B(new_n5289_), .Y(new_n5296_));
  AOI22X1  g05040(.A0(new_n4572_), .A1(\b[6] ), .B0(new_n4571_), .B1(\b[5] ), .Y(new_n5297_));
  OAI21X1  g05041(.A0(new_n4740_), .A1(new_n325_), .B0(new_n5297_), .Y(new_n5298_));
  AOI21X1  g05042(.A0(new_n4375_), .A1(new_n378_), .B0(new_n5298_), .Y(new_n5299_));
  XOR2X1   g05043(.A(new_n5299_), .B(\a[47] ), .Y(new_n5300_));
  XOR2X1   g05044(.A(new_n5300_), .B(new_n5296_), .Y(new_n5301_));
  INVX1    g05045(.A(new_n5301_), .Y(new_n5302_));
  INVX1    g05046(.A(new_n5101_), .Y(new_n5303_));
  NOR2X1   g05047(.A(new_n5102_), .B(new_n5090_), .Y(new_n5304_));
  AOI21X1  g05048(.A0(new_n5303_), .A1(new_n5097_), .B0(new_n5304_), .Y(new_n5305_));
  XOR2X1   g05049(.A(new_n5305_), .B(new_n5302_), .Y(new_n5306_));
  AOI22X1  g05050(.A0(new_n4095_), .A1(\b[9] ), .B0(new_n4094_), .B1(\b[8] ), .Y(new_n5307_));
  OAI21X1  g05051(.A0(new_n4233_), .A1(new_n492_), .B0(new_n5307_), .Y(new_n5308_));
  AOI21X1  g05052(.A0(new_n3901_), .A1(new_n491_), .B0(new_n5308_), .Y(new_n5309_));
  XOR2X1   g05053(.A(new_n5309_), .B(\a[44] ), .Y(new_n5310_));
  XOR2X1   g05054(.A(new_n5310_), .B(new_n5306_), .Y(new_n5311_));
  XOR2X1   g05055(.A(new_n5311_), .B(new_n5285_), .Y(new_n5312_));
  XOR2X1   g05056(.A(new_n5312_), .B(new_n5280_), .Y(new_n5313_));
  XOR2X1   g05057(.A(new_n5313_), .B(new_n5276_), .Y(new_n5314_));
  XOR2X1   g05058(.A(new_n5314_), .B(new_n5271_), .Y(new_n5315_));
  XOR2X1   g05059(.A(new_n5315_), .B(new_n5266_), .Y(new_n5316_));
  XOR2X1   g05060(.A(new_n5316_), .B(new_n5263_), .Y(new_n5317_));
  XOR2X1   g05061(.A(new_n5317_), .B(new_n5259_), .Y(new_n5318_));
  AOI22X1  g05062(.A0(new_n2545_), .A1(\b[21] ), .B0(new_n2544_), .B1(\b[20] ), .Y(new_n5319_));
  OAI21X1  g05063(.A0(new_n2543_), .A1(new_n1300_), .B0(new_n5319_), .Y(new_n5320_));
  AOI21X1  g05064(.A0(new_n2260_), .A1(new_n1299_), .B0(new_n5320_), .Y(new_n5321_));
  XOR2X1   g05065(.A(new_n5321_), .B(\a[32] ), .Y(new_n5322_));
  XOR2X1   g05066(.A(new_n5322_), .B(new_n5318_), .Y(new_n5323_));
  OR2X1    g05067(.A(new_n5124_), .B(new_n5120_), .Y(new_n5324_));
  INVX1    g05068(.A(new_n5124_), .Y(new_n5325_));
  XOR2X1   g05069(.A(new_n5325_), .B(new_n5120_), .Y(new_n5326_));
  OAI21X1  g05070(.A0(new_n5127_), .A1(new_n5326_), .B0(new_n5324_), .Y(new_n5327_));
  XOR2X1   g05071(.A(new_n5327_), .B(new_n5323_), .Y(new_n5328_));
  AOI22X1  g05072(.A0(new_n2163_), .A1(\b[24] ), .B0(new_n2162_), .B1(\b[23] ), .Y(new_n5329_));
  OAI21X1  g05073(.A0(new_n2161_), .A1(new_n1479_), .B0(new_n5329_), .Y(new_n5330_));
  AOI21X1  g05074(.A0(new_n1907_), .A1(new_n1572_), .B0(new_n5330_), .Y(new_n5331_));
  XOR2X1   g05075(.A(new_n5331_), .B(\a[29] ), .Y(new_n5332_));
  XOR2X1   g05076(.A(new_n5332_), .B(new_n5328_), .Y(new_n5333_));
  XOR2X1   g05077(.A(new_n5333_), .B(new_n5137_), .Y(new_n5334_));
  AOI22X1  g05078(.A0(new_n1814_), .A1(\b[27] ), .B0(new_n1813_), .B1(\b[26] ), .Y(new_n5335_));
  OAI21X1  g05079(.A0(new_n1812_), .A1(new_n1880_), .B0(new_n5335_), .Y(new_n5336_));
  AOI21X1  g05080(.A0(new_n1879_), .A1(new_n1617_), .B0(new_n5336_), .Y(new_n5337_));
  XOR2X1   g05081(.A(new_n5337_), .B(\a[26] ), .Y(new_n5338_));
  XOR2X1   g05082(.A(new_n5338_), .B(new_n5334_), .Y(new_n5339_));
  XOR2X1   g05083(.A(new_n5339_), .B(new_n5255_), .Y(new_n5340_));
  AOI22X1  g05084(.A0(new_n1526_), .A1(\b[30] ), .B0(new_n1525_), .B1(\b[29] ), .Y(new_n5341_));
  OAI21X1  g05085(.A0(new_n1524_), .A1(new_n2231_), .B0(new_n5341_), .Y(new_n5342_));
  AOI21X1  g05086(.A0(new_n2230_), .A1(new_n1347_), .B0(new_n5342_), .Y(new_n5343_));
  XOR2X1   g05087(.A(new_n5343_), .B(\a[23] ), .Y(new_n5344_));
  XOR2X1   g05088(.A(new_n5344_), .B(new_n5340_), .Y(new_n5345_));
  XOR2X1   g05089(.A(new_n5345_), .B(new_n5252_), .Y(new_n5346_));
  AOI22X1  g05090(.A0(new_n1263_), .A1(\b[33] ), .B0(new_n1262_), .B1(\b[32] ), .Y(new_n5347_));
  OAI21X1  g05091(.A0(new_n1261_), .A1(new_n2615_), .B0(new_n5347_), .Y(new_n5348_));
  AOI21X1  g05092(.A0(new_n2614_), .A1(new_n1075_), .B0(new_n5348_), .Y(new_n5349_));
  XOR2X1   g05093(.A(new_n5349_), .B(\a[20] ), .Y(new_n5350_));
  XOR2X1   g05094(.A(new_n5350_), .B(new_n5346_), .Y(new_n5351_));
  XOR2X1   g05095(.A(new_n5351_), .B(new_n5248_), .Y(new_n5352_));
  AOI22X1  g05096(.A0(new_n1017_), .A1(\b[36] ), .B0(new_n1016_), .B1(\b[35] ), .Y(new_n5353_));
  OAI21X1  g05097(.A0(new_n1015_), .A1(new_n2890_), .B0(new_n5353_), .Y(new_n5354_));
  AOI21X1  g05098(.A0(new_n3015_), .A1(new_n882_), .B0(new_n5354_), .Y(new_n5355_));
  XOR2X1   g05099(.A(new_n5355_), .B(\a[17] ), .Y(new_n5356_));
  XOR2X1   g05100(.A(new_n5356_), .B(new_n5352_), .Y(new_n5357_));
  XOR2X1   g05101(.A(new_n5357_), .B(new_n5246_), .Y(new_n5358_));
  AOI22X1  g05102(.A0(new_n818_), .A1(\b[39] ), .B0(new_n817_), .B1(\b[38] ), .Y(new_n5359_));
  OAI21X1  g05103(.A0(new_n816_), .A1(new_n3413_), .B0(new_n5359_), .Y(new_n5360_));
  AOI21X1  g05104(.A0(new_n3412_), .A1(new_n668_), .B0(new_n5360_), .Y(new_n5361_));
  XOR2X1   g05105(.A(new_n5361_), .B(\a[14] ), .Y(new_n5362_));
  XOR2X1   g05106(.A(new_n5362_), .B(new_n5358_), .Y(new_n5363_));
  NOR2X1   g05107(.A(new_n5164_), .B(new_n5160_), .Y(new_n5364_));
  OR2X1    g05108(.A(new_n4980_), .B(new_n4976_), .Y(new_n5365_));
  OAI21X1  g05109(.A0(new_n4983_), .A1(new_n5218_), .B0(new_n5365_), .Y(new_n5366_));
  AOI21X1  g05110(.A0(new_n5366_), .A1(new_n5165_), .B0(new_n5364_), .Y(new_n5367_));
  XOR2X1   g05111(.A(new_n5367_), .B(new_n5363_), .Y(new_n5368_));
  AOI22X1  g05112(.A0(new_n603_), .A1(\b[42] ), .B0(new_n602_), .B1(\b[41] ), .Y(new_n5369_));
  OAI21X1  g05113(.A0(new_n601_), .A1(new_n3720_), .B0(new_n5369_), .Y(new_n5370_));
  AOI21X1  g05114(.A0(new_n3860_), .A1(new_n518_), .B0(new_n5370_), .Y(new_n5371_));
  XOR2X1   g05115(.A(new_n5371_), .B(\a[11] ), .Y(new_n5372_));
  XOR2X1   g05116(.A(new_n5372_), .B(new_n5368_), .Y(new_n5373_));
  NOR2X1   g05117(.A(new_n5175_), .B(new_n5171_), .Y(new_n5374_));
  OR2X1    g05118(.A(new_n4988_), .B(new_n4984_), .Y(new_n5375_));
  OAI21X1  g05119(.A0(new_n5001_), .A1(new_n5220_), .B0(new_n5375_), .Y(new_n5376_));
  AOI21X1  g05120(.A0(new_n5376_), .A1(new_n5176_), .B0(new_n5374_), .Y(new_n5377_));
  XOR2X1   g05121(.A(new_n5377_), .B(new_n5373_), .Y(new_n5378_));
  AOI22X1  g05122(.A0(new_n469_), .A1(\b[45] ), .B0(new_n468_), .B1(\b[44] ), .Y(new_n5379_));
  OAI21X1  g05123(.A0(new_n467_), .A1(new_n4339_), .B0(new_n5379_), .Y(new_n5380_));
  AOI21X1  g05124(.A0(new_n4338_), .A1(new_n404_), .B0(new_n5380_), .Y(new_n5381_));
  XOR2X1   g05125(.A(new_n5381_), .B(\a[8] ), .Y(new_n5382_));
  XOR2X1   g05126(.A(new_n5382_), .B(new_n5378_), .Y(new_n5383_));
  XOR2X1   g05127(.A(new_n5383_), .B(new_n5189_), .Y(new_n5384_));
  AOI22X1  g05128(.A0(new_n369_), .A1(\b[48] ), .B0(new_n368_), .B1(\b[47] ), .Y(new_n5385_));
  OAI21X1  g05129(.A0(new_n367_), .A1(new_n4693_), .B0(new_n5385_), .Y(new_n5386_));
  AOI21X1  g05130(.A0(new_n4692_), .A1(new_n308_), .B0(new_n5386_), .Y(new_n5387_));
  XOR2X1   g05131(.A(new_n5387_), .B(\a[5] ), .Y(new_n5388_));
  XOR2X1   g05132(.A(new_n5388_), .B(new_n5384_), .Y(new_n5389_));
  XOR2X1   g05133(.A(new_n5389_), .B(new_n5243_), .Y(new_n5390_));
  XOR2X1   g05134(.A(new_n5390_), .B(new_n5241_), .Y(new_n5391_));
  XOR2X1   g05135(.A(new_n5391_), .B(new_n5231_), .Y(\f[51] ));
  NAND2X1  g05136(.A(new_n5390_), .B(new_n5241_), .Y(new_n5393_));
  OAI21X1  g05137(.A0(new_n5230_), .A1(new_n5229_), .B0(new_n5391_), .Y(new_n5394_));
  AND2X1   g05138(.A(new_n5394_), .B(new_n5393_), .Y(new_n5395_));
  NOR2X1   g05139(.A(new_n5388_), .B(new_n5384_), .Y(new_n5396_));
  AOI21X1  g05140(.A0(new_n5389_), .A1(new_n5243_), .B0(new_n5396_), .Y(new_n5397_));
  NOR2X1   g05141(.A(new_n5338_), .B(new_n5334_), .Y(new_n5398_));
  INVX1    g05142(.A(new_n5339_), .Y(new_n5399_));
  AOI21X1  g05143(.A0(new_n5254_), .A1(new_n5253_), .B0(new_n5399_), .Y(new_n5400_));
  OR2X1    g05144(.A(new_n5400_), .B(new_n5398_), .Y(new_n5401_));
  NOR2X1   g05145(.A(new_n5332_), .B(new_n5328_), .Y(new_n5402_));
  INVX1    g05146(.A(new_n5402_), .Y(new_n5403_));
  AND2X1   g05147(.A(new_n5134_), .B(new_n5070_), .Y(new_n5404_));
  OAI21X1  g05148(.A0(new_n5404_), .A1(new_n5136_), .B0(new_n5333_), .Y(new_n5405_));
  NAND2X1  g05149(.A(new_n5405_), .B(new_n5403_), .Y(new_n5406_));
  INVX1    g05150(.A(new_n5263_), .Y(new_n5407_));
  NAND2X1  g05151(.A(new_n5316_), .B(new_n5407_), .Y(new_n5408_));
  OAI21X1  g05152(.A0(new_n5317_), .A1(new_n5259_), .B0(new_n5408_), .Y(new_n5409_));
  INVX1    g05153(.A(new_n5280_), .Y(new_n5410_));
  AND2X1   g05154(.A(new_n5312_), .B(new_n5410_), .Y(new_n5411_));
  AOI21X1  g05155(.A0(new_n5275_), .A1(new_n5273_), .B0(new_n5313_), .Y(new_n5412_));
  NOR2X1   g05156(.A(new_n5412_), .B(new_n5411_), .Y(new_n5413_));
  INVX1    g05157(.A(new_n5288_), .Y(new_n5414_));
  OR4X1    g05158(.A(new_n5414_), .B(new_n5096_), .C(new_n4884_), .D(new_n4872_), .Y(new_n5415_));
  OAI21X1  g05159(.A0(new_n5295_), .A1(new_n5289_), .B0(new_n5415_), .Y(new_n5416_));
  AND2X1   g05160(.A(new_n4875_), .B(new_n323_), .Y(new_n5417_));
  NOR4X1   g05161(.A(new_n4876_), .B(new_n4874_), .C(new_n4879_), .D(new_n277_), .Y(new_n5418_));
  OAI22X1  g05162(.A0(new_n4881_), .A1(new_n325_), .B0(new_n4878_), .B1(new_n297_), .Y(new_n5419_));
  NOR3X1   g05163(.A(new_n5419_), .B(new_n5418_), .C(new_n5417_), .Y(new_n5420_));
  XOR2X1   g05164(.A(new_n5420_), .B(new_n4873_), .Y(new_n5421_));
  OAI21X1  g05165(.A0(new_n5287_), .A1(new_n274_), .B0(\a[53] ), .Y(new_n5422_));
  INVX1    g05166(.A(\a[53] ), .Y(new_n5423_));
  XOR2X1   g05167(.A(new_n5423_), .B(\a[52] ), .Y(new_n5424_));
  NOR2X1   g05168(.A(new_n5424_), .B(new_n5287_), .Y(new_n5425_));
  XOR2X1   g05169(.A(\a[52] ), .B(\a[51] ), .Y(new_n5426_));
  AND2X1   g05170(.A(new_n5426_), .B(new_n5287_), .Y(new_n5427_));
  INVX1    g05171(.A(new_n5427_), .Y(new_n5428_));
  INVX1    g05172(.A(new_n5287_), .Y(new_n5429_));
  AND2X1   g05173(.A(new_n5424_), .B(new_n5429_), .Y(new_n5430_));
  INVX1    g05174(.A(new_n5430_), .Y(new_n5431_));
  OAI22X1  g05175(.A0(new_n5431_), .A1(new_n275_), .B0(new_n5428_), .B1(new_n274_), .Y(new_n5432_));
  AOI21X1  g05176(.A0(new_n5425_), .A1(new_n263_), .B0(new_n5432_), .Y(new_n5433_));
  XOR2X1   g05177(.A(new_n5433_), .B(\a[53] ), .Y(new_n5434_));
  XOR2X1   g05178(.A(new_n5434_), .B(new_n5422_), .Y(new_n5435_));
  XOR2X1   g05179(.A(new_n5435_), .B(new_n5421_), .Y(new_n5436_));
  XOR2X1   g05180(.A(new_n5436_), .B(new_n5416_), .Y(new_n5437_));
  AOI22X1  g05181(.A0(new_n4572_), .A1(\b[7] ), .B0(new_n4571_), .B1(\b[6] ), .Y(new_n5438_));
  OAI21X1  g05182(.A0(new_n4740_), .A1(new_n395_), .B0(new_n5438_), .Y(new_n5439_));
  AOI21X1  g05183(.A0(new_n4375_), .A1(new_n394_), .B0(new_n5439_), .Y(new_n5440_));
  XOR2X1   g05184(.A(new_n5440_), .B(\a[47] ), .Y(new_n5441_));
  XOR2X1   g05185(.A(new_n5441_), .B(new_n5437_), .Y(new_n5442_));
  INVX1    g05186(.A(new_n5300_), .Y(new_n5443_));
  NOR2X1   g05187(.A(new_n5305_), .B(new_n5301_), .Y(new_n5444_));
  AOI21X1  g05188(.A0(new_n5443_), .A1(new_n5296_), .B0(new_n5444_), .Y(new_n5445_));
  XOR2X1   g05189(.A(new_n5445_), .B(new_n5442_), .Y(new_n5446_));
  INVX1    g05190(.A(new_n5446_), .Y(new_n5447_));
  AOI22X1  g05191(.A0(new_n4095_), .A1(\b[10] ), .B0(new_n4094_), .B1(\b[9] ), .Y(new_n5448_));
  OAI21X1  g05192(.A0(new_n4233_), .A1(new_n489_), .B0(new_n5448_), .Y(new_n5449_));
  AOI21X1  g05193(.A0(new_n3901_), .A1(new_n543_), .B0(new_n5449_), .Y(new_n5450_));
  XOR2X1   g05194(.A(new_n5450_), .B(\a[44] ), .Y(new_n5451_));
  AND2X1   g05195(.A(new_n5451_), .B(new_n5447_), .Y(new_n5452_));
  INVX1    g05196(.A(new_n5452_), .Y(new_n5453_));
  NOR2X1   g05197(.A(new_n5310_), .B(new_n5306_), .Y(new_n5454_));
  INVX1    g05198(.A(new_n5454_), .Y(new_n5455_));
  OAI21X1  g05199(.A0(new_n5284_), .A1(new_n5282_), .B0(new_n5311_), .Y(new_n5456_));
  NOR2X1   g05200(.A(new_n5451_), .B(new_n5447_), .Y(new_n5457_));
  INVX1    g05201(.A(new_n5457_), .Y(new_n5458_));
  AOI22X1  g05202(.A0(new_n5453_), .A1(new_n5458_), .B0(new_n5456_), .B1(new_n5455_), .Y(new_n5459_));
  NAND2X1  g05203(.A(new_n5456_), .B(new_n5455_), .Y(new_n5460_));
  AOI21X1  g05204(.A0(new_n5453_), .A1(new_n5460_), .B0(new_n5457_), .Y(new_n5461_));
  AOI21X1  g05205(.A0(new_n5461_), .A1(new_n5453_), .B0(new_n5459_), .Y(new_n5462_));
  AOI22X1  g05206(.A0(new_n3652_), .A1(\b[13] ), .B0(new_n3651_), .B1(\b[12] ), .Y(new_n5463_));
  OAI21X1  g05207(.A0(new_n3778_), .A1(new_n716_), .B0(new_n5463_), .Y(new_n5464_));
  AOI21X1  g05208(.A0(new_n3480_), .A1(new_n715_), .B0(new_n5464_), .Y(new_n5465_));
  XOR2X1   g05209(.A(new_n5465_), .B(\a[41] ), .Y(new_n5466_));
  XOR2X1   g05210(.A(new_n5466_), .B(new_n5462_), .Y(new_n5467_));
  XOR2X1   g05211(.A(new_n5467_), .B(new_n5413_), .Y(new_n5468_));
  AOI22X1  g05212(.A0(new_n3204_), .A1(\b[16] ), .B0(new_n3203_), .B1(\b[15] ), .Y(new_n5469_));
  OAI21X1  g05213(.A0(new_n3321_), .A1(new_n792_), .B0(new_n5469_), .Y(new_n5470_));
  AOI21X1  g05214(.A0(new_n3080_), .A1(new_n842_), .B0(new_n5470_), .Y(new_n5471_));
  XOR2X1   g05215(.A(new_n5471_), .B(\a[38] ), .Y(new_n5472_));
  XOR2X1   g05216(.A(new_n5472_), .B(new_n5468_), .Y(new_n5473_));
  AND2X1   g05217(.A(new_n5314_), .B(new_n5271_), .Y(new_n5474_));
  AOI21X1  g05218(.A0(new_n5315_), .A1(new_n5266_), .B0(new_n5474_), .Y(new_n5475_));
  XOR2X1   g05219(.A(new_n5475_), .B(new_n5473_), .Y(new_n5476_));
  AOI22X1  g05220(.A0(new_n2813_), .A1(\b[19] ), .B0(new_n2812_), .B1(\b[18] ), .Y(new_n5477_));
  OAI21X1  g05221(.A0(new_n2946_), .A1(new_n1118_), .B0(new_n5477_), .Y(new_n5478_));
  AOI21X1  g05222(.A0(new_n2652_), .A1(new_n1117_), .B0(new_n5478_), .Y(new_n5479_));
  XOR2X1   g05223(.A(new_n5479_), .B(\a[35] ), .Y(new_n5480_));
  NOR2X1   g05224(.A(new_n5480_), .B(new_n5476_), .Y(new_n5481_));
  AND2X1   g05225(.A(new_n5480_), .B(new_n5476_), .Y(new_n5482_));
  OAI21X1  g05226(.A0(new_n5482_), .A1(new_n5481_), .B0(new_n5409_), .Y(new_n5483_));
  NAND2X1  g05227(.A(new_n5480_), .B(new_n5476_), .Y(new_n5484_));
  AOI21X1  g05228(.A0(new_n5484_), .A1(new_n5409_), .B0(new_n5481_), .Y(new_n5485_));
  NAND2X1  g05229(.A(new_n5485_), .B(new_n5484_), .Y(new_n5486_));
  NAND2X1  g05230(.A(new_n5486_), .B(new_n5483_), .Y(new_n5487_));
  AOI22X1  g05231(.A0(new_n2545_), .A1(\b[22] ), .B0(new_n2544_), .B1(\b[21] ), .Y(new_n5488_));
  OAI21X1  g05232(.A0(new_n2543_), .A1(new_n1297_), .B0(new_n5488_), .Y(new_n5489_));
  AOI21X1  g05233(.A0(new_n2260_), .A1(new_n1399_), .B0(new_n5489_), .Y(new_n5490_));
  XOR2X1   g05234(.A(new_n5490_), .B(\a[32] ), .Y(new_n5491_));
  XOR2X1   g05235(.A(new_n5491_), .B(new_n5487_), .Y(new_n5492_));
  INVX1    g05236(.A(new_n5318_), .Y(new_n5493_));
  NOR2X1   g05237(.A(new_n5322_), .B(new_n5493_), .Y(new_n5494_));
  INVX1    g05238(.A(new_n5323_), .Y(new_n5495_));
  AOI21X1  g05239(.A0(new_n5327_), .A1(new_n5495_), .B0(new_n5494_), .Y(new_n5496_));
  XOR2X1   g05240(.A(new_n5496_), .B(new_n5492_), .Y(new_n5497_));
  AOI22X1  g05241(.A0(new_n2163_), .A1(\b[25] ), .B0(new_n2162_), .B1(\b[24] ), .Y(new_n5498_));
  OAI21X1  g05242(.A0(new_n2161_), .A1(new_n1591_), .B0(new_n5498_), .Y(new_n5499_));
  AOI21X1  g05243(.A0(new_n1907_), .A1(new_n1590_), .B0(new_n5499_), .Y(new_n5500_));
  XOR2X1   g05244(.A(new_n5500_), .B(\a[29] ), .Y(new_n5501_));
  XOR2X1   g05245(.A(new_n5501_), .B(new_n5497_), .Y(new_n5502_));
  XOR2X1   g05246(.A(new_n5502_), .B(new_n5406_), .Y(new_n5503_));
  AOI22X1  g05247(.A0(new_n1814_), .A1(\b[28] ), .B0(new_n1813_), .B1(\b[27] ), .Y(new_n5504_));
  OAI21X1  g05248(.A0(new_n1812_), .A1(new_n1877_), .B0(new_n5504_), .Y(new_n5505_));
  AOI21X1  g05249(.A0(new_n2004_), .A1(new_n1617_), .B0(new_n5505_), .Y(new_n5506_));
  XOR2X1   g05250(.A(new_n5506_), .B(\a[26] ), .Y(new_n5507_));
  XOR2X1   g05251(.A(new_n5507_), .B(new_n5503_), .Y(new_n5508_));
  XOR2X1   g05252(.A(new_n5508_), .B(new_n5401_), .Y(new_n5509_));
  AOI22X1  g05253(.A0(new_n1526_), .A1(\b[31] ), .B0(new_n1525_), .B1(\b[30] ), .Y(new_n5510_));
  OAI21X1  g05254(.A0(new_n1524_), .A1(new_n2359_), .B0(new_n5510_), .Y(new_n5511_));
  AOI21X1  g05255(.A0(new_n2358_), .A1(new_n1347_), .B0(new_n5511_), .Y(new_n5512_));
  XOR2X1   g05256(.A(new_n5512_), .B(\a[23] ), .Y(new_n5513_));
  INVX1    g05257(.A(new_n5513_), .Y(new_n5514_));
  XOR2X1   g05258(.A(new_n5514_), .B(new_n5509_), .Y(new_n5515_));
  OR2X1    g05259(.A(new_n5344_), .B(new_n5340_), .Y(new_n5516_));
  OAI21X1  g05260(.A0(new_n5251_), .A1(new_n5250_), .B0(new_n5345_), .Y(new_n5517_));
  AND2X1   g05261(.A(new_n5517_), .B(new_n5516_), .Y(new_n5518_));
  XOR2X1   g05262(.A(new_n5518_), .B(new_n5515_), .Y(new_n5519_));
  AOI22X1  g05263(.A0(new_n1263_), .A1(\b[34] ), .B0(new_n1262_), .B1(\b[33] ), .Y(new_n5520_));
  OAI21X1  g05264(.A0(new_n1261_), .A1(new_n2612_), .B0(new_n5520_), .Y(new_n5521_));
  AOI21X1  g05265(.A0(new_n2759_), .A1(new_n1075_), .B0(new_n5521_), .Y(new_n5522_));
  XOR2X1   g05266(.A(new_n5522_), .B(\a[20] ), .Y(new_n5523_));
  XOR2X1   g05267(.A(new_n5523_), .B(new_n5519_), .Y(new_n5524_));
  OR2X1    g05268(.A(new_n5350_), .B(new_n5346_), .Y(new_n5525_));
  XOR2X1   g05269(.A(new_n5349_), .B(new_n1072_), .Y(new_n5526_));
  XOR2X1   g05270(.A(new_n5526_), .B(new_n5346_), .Y(new_n5527_));
  OAI21X1  g05271(.A0(new_n5527_), .A1(new_n5248_), .B0(new_n5525_), .Y(new_n5528_));
  XOR2X1   g05272(.A(new_n5528_), .B(new_n5524_), .Y(new_n5529_));
  AOI22X1  g05273(.A0(new_n1017_), .A1(\b[37] ), .B0(new_n1016_), .B1(\b[36] ), .Y(new_n5530_));
  OAI21X1  g05274(.A0(new_n1015_), .A1(new_n3156_), .B0(new_n5530_), .Y(new_n5531_));
  AOI21X1  g05275(.A0(new_n3155_), .A1(new_n882_), .B0(new_n5531_), .Y(new_n5532_));
  XOR2X1   g05276(.A(new_n5532_), .B(\a[17] ), .Y(new_n5533_));
  XOR2X1   g05277(.A(new_n5533_), .B(new_n5529_), .Y(new_n5534_));
  NOR2X1   g05278(.A(new_n5356_), .B(new_n5352_), .Y(new_n5535_));
  AOI21X1  g05279(.A0(new_n5357_), .A1(new_n5246_), .B0(new_n5535_), .Y(new_n5536_));
  XOR2X1   g05280(.A(new_n5536_), .B(new_n5534_), .Y(new_n5537_));
  AOI22X1  g05281(.A0(new_n818_), .A1(\b[40] ), .B0(new_n817_), .B1(\b[39] ), .Y(new_n5538_));
  OAI21X1  g05282(.A0(new_n816_), .A1(new_n3575_), .B0(new_n5538_), .Y(new_n5539_));
  AOI21X1  g05283(.A0(new_n3574_), .A1(new_n668_), .B0(new_n5539_), .Y(new_n5540_));
  XOR2X1   g05284(.A(new_n5540_), .B(\a[14] ), .Y(new_n5541_));
  XOR2X1   g05285(.A(new_n5541_), .B(new_n5537_), .Y(new_n5542_));
  INVX1    g05286(.A(new_n5362_), .Y(new_n5543_));
  NAND2X1  g05287(.A(new_n5543_), .B(new_n5358_), .Y(new_n5544_));
  OAI21X1  g05288(.A0(new_n5367_), .A1(new_n5363_), .B0(new_n5544_), .Y(new_n5545_));
  XOR2X1   g05289(.A(new_n5545_), .B(new_n5542_), .Y(new_n5546_));
  AOI22X1  g05290(.A0(new_n603_), .A1(\b[43] ), .B0(new_n602_), .B1(\b[42] ), .Y(new_n5547_));
  OAI21X1  g05291(.A0(new_n601_), .A1(new_n4015_), .B0(new_n5547_), .Y(new_n5548_));
  AOI21X1  g05292(.A0(new_n4014_), .A1(new_n518_), .B0(new_n5548_), .Y(new_n5549_));
  XOR2X1   g05293(.A(new_n5549_), .B(\a[11] ), .Y(new_n5550_));
  NAND2X1  g05294(.A(new_n5550_), .B(new_n5546_), .Y(new_n5551_));
  XOR2X1   g05295(.A(new_n5543_), .B(new_n5358_), .Y(new_n5552_));
  XOR2X1   g05296(.A(new_n5367_), .B(new_n5552_), .Y(new_n5553_));
  NOR2X1   g05297(.A(new_n5372_), .B(new_n5553_), .Y(new_n5554_));
  XOR2X1   g05298(.A(new_n5372_), .B(new_n5553_), .Y(new_n5555_));
  OR2X1    g05299(.A(new_n5175_), .B(new_n5171_), .Y(new_n5556_));
  XOR2X1   g05300(.A(new_n5159_), .B(new_n5245_), .Y(new_n5557_));
  XOR2X1   g05301(.A(new_n5164_), .B(new_n5557_), .Y(new_n5558_));
  XOR2X1   g05302(.A(new_n5170_), .B(new_n5558_), .Y(new_n5559_));
  XOR2X1   g05303(.A(new_n5175_), .B(new_n5559_), .Y(new_n5560_));
  OAI21X1  g05304(.A0(new_n5180_), .A1(new_n5560_), .B0(new_n5556_), .Y(new_n5561_));
  AOI21X1  g05305(.A0(new_n5561_), .A1(new_n5555_), .B0(new_n5554_), .Y(new_n5562_));
  OR2X1    g05306(.A(new_n5550_), .B(new_n5546_), .Y(new_n5563_));
  AOI21X1  g05307(.A0(new_n5551_), .A1(new_n5563_), .B0(new_n5562_), .Y(new_n5564_));
  OR2X1    g05308(.A(new_n5372_), .B(new_n5553_), .Y(new_n5565_));
  OAI21X1  g05309(.A0(new_n5377_), .A1(new_n5373_), .B0(new_n5565_), .Y(new_n5566_));
  NOR2X1   g05310(.A(new_n5550_), .B(new_n5546_), .Y(new_n5567_));
  AOI21X1  g05311(.A0(new_n5551_), .A1(new_n5566_), .B0(new_n5567_), .Y(new_n5568_));
  AOI21X1  g05312(.A0(new_n5568_), .A1(new_n5551_), .B0(new_n5564_), .Y(new_n5569_));
  AOI22X1  g05313(.A0(new_n469_), .A1(\b[46] ), .B0(new_n468_), .B1(\b[45] ), .Y(new_n5570_));
  OAI21X1  g05314(.A0(new_n467_), .A1(new_n4336_), .B0(new_n5570_), .Y(new_n5571_));
  AOI21X1  g05315(.A0(new_n4509_), .A1(new_n404_), .B0(new_n5571_), .Y(new_n5572_));
  XOR2X1   g05316(.A(new_n5572_), .B(\a[8] ), .Y(new_n5573_));
  INVX1    g05317(.A(new_n5573_), .Y(new_n5574_));
  XOR2X1   g05318(.A(new_n5574_), .B(new_n5569_), .Y(new_n5575_));
  XOR2X1   g05319(.A(new_n5377_), .B(new_n5555_), .Y(new_n5576_));
  OR2X1    g05320(.A(new_n5382_), .B(new_n5576_), .Y(new_n5577_));
  OR2X1    g05321(.A(new_n5383_), .B(new_n5225_), .Y(new_n5578_));
  AND2X1   g05322(.A(new_n5578_), .B(new_n5577_), .Y(new_n5579_));
  XOR2X1   g05323(.A(new_n5579_), .B(new_n5575_), .Y(new_n5580_));
  AOI22X1  g05324(.A0(new_n369_), .A1(\b[49] ), .B0(new_n368_), .B1(\b[48] ), .Y(new_n5581_));
  OAI21X1  g05325(.A0(new_n367_), .A1(new_n5039_), .B0(new_n5581_), .Y(new_n5582_));
  AOI21X1  g05326(.A0(new_n5038_), .A1(new_n308_), .B0(new_n5582_), .Y(new_n5583_));
  XOR2X1   g05327(.A(new_n5583_), .B(\a[5] ), .Y(new_n5584_));
  XOR2X1   g05328(.A(new_n5584_), .B(new_n5580_), .Y(new_n5585_));
  XOR2X1   g05329(.A(new_n5585_), .B(new_n5397_), .Y(new_n5586_));
  NAND2X1  g05330(.A(\b[51] ), .B(\b[50] ), .Y(new_n5587_));
  OAI21X1  g05331(.A0(new_n5235_), .A1(new_n5233_), .B0(new_n5587_), .Y(new_n5588_));
  XOR2X1   g05332(.A(\b[52] ), .B(\b[51] ), .Y(new_n5589_));
  XOR2X1   g05333(.A(new_n5589_), .B(new_n5588_), .Y(new_n5590_));
  AOI22X1  g05334(.A0(new_n267_), .A1(\b[52] ), .B0(new_n266_), .B1(\b[51] ), .Y(new_n5591_));
  OAI21X1  g05335(.A0(new_n350_), .A1(new_n5234_), .B0(new_n5591_), .Y(new_n5592_));
  AOI21X1  g05336(.A0(new_n5590_), .A1(new_n318_), .B0(new_n5592_), .Y(new_n5593_));
  XOR2X1   g05337(.A(new_n5593_), .B(\a[2] ), .Y(new_n5594_));
  XOR2X1   g05338(.A(new_n5594_), .B(new_n5586_), .Y(new_n5595_));
  XOR2X1   g05339(.A(new_n5595_), .B(new_n5395_), .Y(\f[52] ));
  NOR2X1   g05340(.A(new_n5194_), .B(new_n5226_), .Y(new_n5597_));
  OR2X1    g05341(.A(new_n5018_), .B(new_n5014_), .Y(new_n5598_));
  XOR2X1   g05342(.A(new_n5013_), .B(new_n5222_), .Y(new_n5599_));
  XOR2X1   g05343(.A(new_n5018_), .B(new_n5599_), .Y(new_n5600_));
  OAI21X1  g05344(.A0(new_n5032_), .A1(new_n5600_), .B0(new_n5598_), .Y(new_n5601_));
  AOI21X1  g05345(.A0(new_n5601_), .A1(new_n5227_), .B0(new_n5597_), .Y(new_n5602_));
  AND2X1   g05346(.A(new_n5388_), .B(new_n5384_), .Y(new_n5603_));
  OR2X1    g05347(.A(new_n5388_), .B(new_n5384_), .Y(new_n5604_));
  OAI21X1  g05348(.A0(new_n5603_), .A1(new_n5602_), .B0(new_n5604_), .Y(new_n5605_));
  XOR2X1   g05349(.A(new_n5585_), .B(new_n5605_), .Y(new_n5606_));
  NOR2X1   g05350(.A(new_n5594_), .B(new_n5606_), .Y(new_n5607_));
  AOI21X1  g05351(.A0(new_n5394_), .A1(new_n5393_), .B0(new_n5595_), .Y(new_n5608_));
  XOR2X1   g05352(.A(new_n5573_), .B(new_n5569_), .Y(new_n5609_));
  XOR2X1   g05353(.A(new_n5579_), .B(new_n5609_), .Y(new_n5610_));
  OR2X1    g05354(.A(new_n5584_), .B(new_n5610_), .Y(new_n5611_));
  OAI21X1  g05355(.A0(new_n5585_), .A1(new_n5397_), .B0(new_n5611_), .Y(new_n5612_));
  NAND2X1  g05356(.A(new_n5514_), .B(new_n5509_), .Y(new_n5613_));
  XOR2X1   g05357(.A(new_n5513_), .B(new_n5509_), .Y(new_n5614_));
  OAI21X1  g05358(.A0(new_n5518_), .A1(new_n5614_), .B0(new_n5613_), .Y(new_n5615_));
  AOI22X1  g05359(.A0(new_n1526_), .A1(\b[32] ), .B0(new_n1525_), .B1(\b[31] ), .Y(new_n5616_));
  OAI21X1  g05360(.A0(new_n1524_), .A1(new_n2356_), .B0(new_n5616_), .Y(new_n5617_));
  AOI21X1  g05361(.A0(new_n2495_), .A1(new_n1347_), .B0(new_n5617_), .Y(new_n5618_));
  XOR2X1   g05362(.A(new_n5618_), .B(\a[23] ), .Y(new_n5619_));
  INVX1    g05363(.A(new_n5619_), .Y(new_n5620_));
  OAI21X1  g05364(.A0(new_n5400_), .A1(new_n5398_), .B0(new_n5508_), .Y(new_n5621_));
  OAI21X1  g05365(.A0(new_n5507_), .A1(new_n5503_), .B0(new_n5621_), .Y(new_n5622_));
  AOI22X1  g05366(.A0(new_n1814_), .A1(\b[29] ), .B0(new_n1813_), .B1(\b[28] ), .Y(new_n5623_));
  OAI21X1  g05367(.A0(new_n1812_), .A1(new_n2126_), .B0(new_n5623_), .Y(new_n5624_));
  AOI21X1  g05368(.A0(new_n2125_), .A1(new_n1617_), .B0(new_n5624_), .Y(new_n5625_));
  XOR2X1   g05369(.A(new_n5625_), .B(\a[26] ), .Y(new_n5626_));
  INVX1    g05370(.A(new_n5626_), .Y(new_n5627_));
  AND2X1   g05371(.A(new_n5405_), .B(new_n5403_), .Y(new_n5628_));
  XOR2X1   g05372(.A(new_n5500_), .B(new_n1911_), .Y(new_n5629_));
  NAND2X1  g05373(.A(new_n5629_), .B(new_n5497_), .Y(new_n5630_));
  OAI21X1  g05374(.A0(new_n5502_), .A1(new_n5628_), .B0(new_n5630_), .Y(new_n5631_));
  AND2X1   g05375(.A(new_n5486_), .B(new_n5483_), .Y(new_n5632_));
  OR2X1    g05376(.A(new_n5491_), .B(new_n5632_), .Y(new_n5633_));
  OAI21X1  g05377(.A0(new_n5496_), .A1(new_n5492_), .B0(new_n5633_), .Y(new_n5634_));
  AOI22X1  g05378(.A0(new_n2545_), .A1(\b[23] ), .B0(new_n2544_), .B1(\b[22] ), .Y(new_n5635_));
  OAI21X1  g05379(.A0(new_n2543_), .A1(new_n1482_), .B0(new_n5635_), .Y(new_n5636_));
  AOI21X1  g05380(.A0(new_n2260_), .A1(new_n1481_), .B0(new_n5636_), .Y(new_n5637_));
  XOR2X1   g05381(.A(new_n5637_), .B(\a[32] ), .Y(new_n5638_));
  OR2X1    g05382(.A(new_n5472_), .B(new_n5468_), .Y(new_n5639_));
  INVX1    g05383(.A(new_n5473_), .Y(new_n5640_));
  OAI21X1  g05384(.A0(new_n5475_), .A1(new_n5640_), .B0(new_n5639_), .Y(new_n5641_));
  AOI22X1  g05385(.A0(new_n3204_), .A1(\b[17] ), .B0(new_n3203_), .B1(\b[16] ), .Y(new_n5642_));
  OAI21X1  g05386(.A0(new_n3321_), .A1(new_n977_), .B0(new_n5642_), .Y(new_n5643_));
  AOI21X1  g05387(.A0(new_n3080_), .A1(new_n976_), .B0(new_n5643_), .Y(new_n5644_));
  XOR2X1   g05388(.A(new_n5644_), .B(\a[38] ), .Y(new_n5645_));
  INVX1    g05389(.A(new_n5645_), .Y(new_n5646_));
  INVX1    g05390(.A(new_n5413_), .Y(new_n5647_));
  NOR2X1   g05391(.A(new_n5466_), .B(new_n5462_), .Y(new_n5648_));
  AOI21X1  g05392(.A0(new_n5467_), .A1(new_n5647_), .B0(new_n5648_), .Y(new_n5649_));
  INVX1    g05393(.A(new_n5461_), .Y(new_n5650_));
  AOI22X1  g05394(.A0(new_n4095_), .A1(\b[11] ), .B0(new_n4094_), .B1(\b[10] ), .Y(new_n5651_));
  OAI21X1  g05395(.A0(new_n4233_), .A1(new_n590_), .B0(new_n5651_), .Y(new_n5652_));
  AOI21X1  g05396(.A0(new_n3901_), .A1(new_n589_), .B0(new_n5652_), .Y(new_n5653_));
  XOR2X1   g05397(.A(new_n5653_), .B(new_n3899_), .Y(new_n5654_));
  XOR2X1   g05398(.A(new_n5440_), .B(new_n4568_), .Y(new_n5655_));
  NAND2X1  g05399(.A(new_n5655_), .B(new_n5437_), .Y(new_n5656_));
  OAI21X1  g05400(.A0(new_n5445_), .A1(new_n5442_), .B0(new_n5656_), .Y(new_n5657_));
  AND2X1   g05401(.A(new_n5435_), .B(new_n5421_), .Y(new_n5658_));
  AND2X1   g05402(.A(new_n5436_), .B(new_n5416_), .Y(new_n5659_));
  OR2X1    g05403(.A(new_n5659_), .B(new_n5658_), .Y(new_n5660_));
  NAND3X1  g05404(.A(new_n5433_), .B(new_n5414_), .C(\a[53] ), .Y(new_n5661_));
  NAND2X1  g05405(.A(new_n5425_), .B(new_n341_), .Y(new_n5662_));
  OR4X1    g05406(.A(new_n5426_), .B(new_n5424_), .C(new_n5429_), .D(new_n274_), .Y(new_n5663_));
  AOI22X1  g05407(.A0(new_n5430_), .A1(\b[2] ), .B0(new_n5427_), .B1(\b[1] ), .Y(new_n5664_));
  NAND3X1  g05408(.A(new_n5664_), .B(new_n5663_), .C(new_n5662_), .Y(new_n5665_));
  XOR2X1   g05409(.A(new_n5665_), .B(new_n5423_), .Y(new_n5666_));
  XOR2X1   g05410(.A(new_n5666_), .B(new_n5661_), .Y(new_n5667_));
  INVX1    g05411(.A(new_n5667_), .Y(new_n5668_));
  AOI22X1  g05412(.A0(new_n4880_), .A1(\b[5] ), .B0(new_n4877_), .B1(\b[4] ), .Y(new_n5669_));
  OAI21X1  g05413(.A0(new_n5291_), .A1(new_n297_), .B0(new_n5669_), .Y(new_n5670_));
  AOI21X1  g05414(.A0(new_n4875_), .A1(new_n349_), .B0(new_n5670_), .Y(new_n5671_));
  XOR2X1   g05415(.A(new_n5671_), .B(\a[50] ), .Y(new_n5672_));
  NAND2X1  g05416(.A(new_n5672_), .B(new_n5668_), .Y(new_n5673_));
  XOR2X1   g05417(.A(new_n5672_), .B(new_n5668_), .Y(new_n5674_));
  INVX1    g05418(.A(new_n5674_), .Y(new_n5675_));
  NOR2X1   g05419(.A(new_n5672_), .B(new_n5668_), .Y(new_n5676_));
  AOI21X1  g05420(.A0(new_n5673_), .A1(new_n5660_), .B0(new_n5676_), .Y(new_n5677_));
  AOI22X1  g05421(.A0(new_n5677_), .A1(new_n5673_), .B0(new_n5675_), .B1(new_n5660_), .Y(new_n5678_));
  AOI22X1  g05422(.A0(new_n4572_), .A1(\b[8] ), .B0(new_n4571_), .B1(\b[7] ), .Y(new_n5679_));
  OAI21X1  g05423(.A0(new_n4740_), .A1(new_n392_), .B0(new_n5679_), .Y(new_n5680_));
  AOI21X1  g05424(.A0(new_n4375_), .A1(new_n454_), .B0(new_n5680_), .Y(new_n5681_));
  XOR2X1   g05425(.A(new_n5681_), .B(\a[47] ), .Y(new_n5682_));
  XOR2X1   g05426(.A(new_n5682_), .B(new_n5678_), .Y(new_n5683_));
  XOR2X1   g05427(.A(new_n5683_), .B(new_n5657_), .Y(new_n5684_));
  XOR2X1   g05428(.A(new_n5684_), .B(new_n5654_), .Y(new_n5685_));
  XOR2X1   g05429(.A(new_n5685_), .B(new_n5650_), .Y(new_n5686_));
  AOI22X1  g05430(.A0(new_n3652_), .A1(\b[14] ), .B0(new_n3651_), .B1(\b[13] ), .Y(new_n5687_));
  OAI21X1  g05431(.A0(new_n3778_), .A1(new_n713_), .B0(new_n5687_), .Y(new_n5688_));
  AOI21X1  g05432(.A0(new_n3480_), .A1(new_n734_), .B0(new_n5688_), .Y(new_n5689_));
  XOR2X1   g05433(.A(new_n5689_), .B(\a[41] ), .Y(new_n5690_));
  XOR2X1   g05434(.A(new_n5690_), .B(new_n5686_), .Y(new_n5691_));
  XOR2X1   g05435(.A(new_n5691_), .B(new_n5649_), .Y(new_n5692_));
  XOR2X1   g05436(.A(new_n5692_), .B(new_n5646_), .Y(new_n5693_));
  XOR2X1   g05437(.A(new_n5693_), .B(new_n5641_), .Y(new_n5694_));
  AOI22X1  g05438(.A0(new_n2813_), .A1(\b[20] ), .B0(new_n2812_), .B1(\b[19] ), .Y(new_n5695_));
  OAI21X1  g05439(.A0(new_n2946_), .A1(new_n1115_), .B0(new_n5695_), .Y(new_n5696_));
  AOI21X1  g05440(.A0(new_n2652_), .A1(new_n1217_), .B0(new_n5696_), .Y(new_n5697_));
  XOR2X1   g05441(.A(new_n5697_), .B(\a[35] ), .Y(new_n5698_));
  XOR2X1   g05442(.A(new_n5698_), .B(new_n5694_), .Y(new_n5699_));
  XOR2X1   g05443(.A(new_n5699_), .B(new_n5485_), .Y(new_n5700_));
  XOR2X1   g05444(.A(new_n5700_), .B(new_n5638_), .Y(new_n5701_));
  XOR2X1   g05445(.A(new_n5701_), .B(new_n5634_), .Y(new_n5702_));
  AOI22X1  g05446(.A0(new_n2163_), .A1(\b[26] ), .B0(new_n2162_), .B1(\b[25] ), .Y(new_n5703_));
  OAI21X1  g05447(.A0(new_n2161_), .A1(new_n1588_), .B0(new_n5703_), .Y(new_n5704_));
  AOI21X1  g05448(.A0(new_n1907_), .A1(new_n1783_), .B0(new_n5704_), .Y(new_n5705_));
  XOR2X1   g05449(.A(new_n5705_), .B(\a[29] ), .Y(new_n5706_));
  XOR2X1   g05450(.A(new_n5706_), .B(new_n5702_), .Y(new_n5707_));
  XOR2X1   g05451(.A(new_n5707_), .B(new_n5631_), .Y(new_n5708_));
  XOR2X1   g05452(.A(new_n5708_), .B(new_n5627_), .Y(new_n5709_));
  XOR2X1   g05453(.A(new_n5709_), .B(new_n5622_), .Y(new_n5710_));
  XOR2X1   g05454(.A(new_n5710_), .B(new_n5620_), .Y(new_n5711_));
  XOR2X1   g05455(.A(new_n5711_), .B(new_n5615_), .Y(new_n5712_));
  AOI22X1  g05456(.A0(new_n1263_), .A1(\b[35] ), .B0(new_n1262_), .B1(\b[34] ), .Y(new_n5713_));
  OAI21X1  g05457(.A0(new_n1261_), .A1(new_n2893_), .B0(new_n5713_), .Y(new_n5714_));
  AOI21X1  g05458(.A0(new_n2892_), .A1(new_n1075_), .B0(new_n5714_), .Y(new_n5715_));
  XOR2X1   g05459(.A(new_n5715_), .B(\a[20] ), .Y(new_n5716_));
  XOR2X1   g05460(.A(new_n5716_), .B(new_n5712_), .Y(new_n5717_));
  NOR2X1   g05461(.A(new_n5523_), .B(new_n5519_), .Y(new_n5718_));
  AOI21X1  g05462(.A0(new_n5528_), .A1(new_n5524_), .B0(new_n5718_), .Y(new_n5719_));
  XOR2X1   g05463(.A(new_n5719_), .B(new_n5717_), .Y(new_n5720_));
  AOI22X1  g05464(.A0(new_n1017_), .A1(\b[38] ), .B0(new_n1016_), .B1(\b[37] ), .Y(new_n5721_));
  OAI21X1  g05465(.A0(new_n1015_), .A1(new_n3276_), .B0(new_n5721_), .Y(new_n5722_));
  AOI21X1  g05466(.A0(new_n3275_), .A1(new_n882_), .B0(new_n5722_), .Y(new_n5723_));
  XOR2X1   g05467(.A(new_n5723_), .B(\a[17] ), .Y(new_n5724_));
  XOR2X1   g05468(.A(new_n5724_), .B(new_n5720_), .Y(new_n5725_));
  XOR2X1   g05469(.A(new_n5518_), .B(new_n5614_), .Y(new_n5726_));
  XOR2X1   g05470(.A(new_n5523_), .B(new_n5726_), .Y(new_n5727_));
  XOR2X1   g05471(.A(new_n5528_), .B(new_n5727_), .Y(new_n5728_));
  OR2X1    g05472(.A(new_n5533_), .B(new_n5728_), .Y(new_n5729_));
  OAI21X1  g05473(.A0(new_n5536_), .A1(new_n5534_), .B0(new_n5729_), .Y(new_n5730_));
  XOR2X1   g05474(.A(new_n5730_), .B(new_n5725_), .Y(new_n5731_));
  AOI22X1  g05475(.A0(new_n818_), .A1(\b[41] ), .B0(new_n817_), .B1(\b[40] ), .Y(new_n5732_));
  OAI21X1  g05476(.A0(new_n816_), .A1(new_n3723_), .B0(new_n5732_), .Y(new_n5733_));
  AOI21X1  g05477(.A0(new_n3722_), .A1(new_n668_), .B0(new_n5733_), .Y(new_n5734_));
  XOR2X1   g05478(.A(new_n5734_), .B(\a[14] ), .Y(new_n5735_));
  XOR2X1   g05479(.A(new_n5735_), .B(new_n5731_), .Y(new_n5736_));
  XOR2X1   g05480(.A(new_n5533_), .B(new_n5728_), .Y(new_n5737_));
  XOR2X1   g05481(.A(new_n5536_), .B(new_n5737_), .Y(new_n5738_));
  NOR2X1   g05482(.A(new_n5541_), .B(new_n5738_), .Y(new_n5739_));
  XOR2X1   g05483(.A(new_n5541_), .B(new_n5738_), .Y(new_n5740_));
  AOI21X1  g05484(.A0(new_n5545_), .A1(new_n5740_), .B0(new_n5739_), .Y(new_n5741_));
  XOR2X1   g05485(.A(new_n5741_), .B(new_n5736_), .Y(new_n5742_));
  AOI22X1  g05486(.A0(new_n603_), .A1(\b[44] ), .B0(new_n602_), .B1(\b[43] ), .Y(new_n5743_));
  OAI21X1  g05487(.A0(new_n601_), .A1(new_n4012_), .B0(new_n5743_), .Y(new_n5744_));
  AOI21X1  g05488(.A0(new_n4178_), .A1(new_n518_), .B0(new_n5744_), .Y(new_n5745_));
  XOR2X1   g05489(.A(new_n5745_), .B(\a[11] ), .Y(new_n5746_));
  AND2X1   g05490(.A(new_n5746_), .B(new_n5742_), .Y(new_n5747_));
  XOR2X1   g05491(.A(new_n5746_), .B(new_n5742_), .Y(new_n5748_));
  OR2X1    g05492(.A(new_n5746_), .B(new_n5742_), .Y(new_n5749_));
  OAI21X1  g05493(.A0(new_n5747_), .A1(new_n5568_), .B0(new_n5749_), .Y(new_n5750_));
  OAI22X1  g05494(.A0(new_n5750_), .A1(new_n5747_), .B0(new_n5748_), .B1(new_n5568_), .Y(new_n5751_));
  AOI22X1  g05495(.A0(new_n469_), .A1(\b[47] ), .B0(new_n468_), .B1(\b[46] ), .Y(new_n5752_));
  OAI21X1  g05496(.A0(new_n467_), .A1(new_n4674_), .B0(new_n5752_), .Y(new_n5753_));
  AOI21X1  g05497(.A0(new_n4673_), .A1(new_n404_), .B0(new_n5753_), .Y(new_n5754_));
  XOR2X1   g05498(.A(new_n5754_), .B(\a[8] ), .Y(new_n5755_));
  XOR2X1   g05499(.A(new_n5755_), .B(new_n5751_), .Y(new_n5756_));
  NOR2X1   g05500(.A(new_n5573_), .B(new_n5569_), .Y(new_n5757_));
  OAI21X1  g05501(.A0(new_n5383_), .A1(new_n5225_), .B0(new_n5577_), .Y(new_n5758_));
  AOI21X1  g05502(.A0(new_n5758_), .A1(new_n5609_), .B0(new_n5757_), .Y(new_n5759_));
  XOR2X1   g05503(.A(new_n5759_), .B(new_n5756_), .Y(new_n5760_));
  AOI22X1  g05504(.A0(new_n369_), .A1(\b[50] ), .B0(new_n368_), .B1(\b[49] ), .Y(new_n5761_));
  OAI21X1  g05505(.A0(new_n367_), .A1(new_n5036_), .B0(new_n5761_), .Y(new_n5762_));
  AOI21X1  g05506(.A0(new_n5204_), .A1(new_n308_), .B0(new_n5762_), .Y(new_n5763_));
  XOR2X1   g05507(.A(new_n5763_), .B(\a[5] ), .Y(new_n5764_));
  XOR2X1   g05508(.A(new_n5764_), .B(new_n5760_), .Y(new_n5765_));
  NAND2X1  g05509(.A(new_n5765_), .B(new_n5612_), .Y(new_n5766_));
  NOR2X1   g05510(.A(new_n5584_), .B(new_n5610_), .Y(new_n5767_));
  XOR2X1   g05511(.A(new_n5584_), .B(new_n5610_), .Y(new_n5768_));
  AOI21X1  g05512(.A0(new_n5768_), .A1(new_n5605_), .B0(new_n5767_), .Y(new_n5769_));
  NAND2X1  g05513(.A(new_n5746_), .B(new_n5742_), .Y(new_n5770_));
  NOR2X1   g05514(.A(new_n5748_), .B(new_n5568_), .Y(new_n5771_));
  AND2X1   g05515(.A(new_n5550_), .B(new_n5546_), .Y(new_n5772_));
  OAI21X1  g05516(.A0(new_n5772_), .A1(new_n5562_), .B0(new_n5563_), .Y(new_n5773_));
  NOR2X1   g05517(.A(new_n5746_), .B(new_n5742_), .Y(new_n5774_));
  AOI21X1  g05518(.A0(new_n5770_), .A1(new_n5773_), .B0(new_n5774_), .Y(new_n5775_));
  AOI21X1  g05519(.A0(new_n5775_), .A1(new_n5770_), .B0(new_n5771_), .Y(new_n5776_));
  XOR2X1   g05520(.A(new_n5755_), .B(new_n5776_), .Y(new_n5777_));
  XOR2X1   g05521(.A(new_n5759_), .B(new_n5777_), .Y(new_n5778_));
  OR2X1    g05522(.A(new_n5764_), .B(new_n5778_), .Y(new_n5779_));
  NAND2X1  g05523(.A(new_n5764_), .B(new_n5778_), .Y(new_n5780_));
  NAND3X1  g05524(.A(new_n5780_), .B(new_n5779_), .C(new_n5769_), .Y(new_n5781_));
  AND2X1   g05525(.A(\b[52] ), .B(\b[51] ), .Y(new_n5782_));
  AOI21X1  g05526(.A0(new_n5589_), .A1(new_n5588_), .B0(new_n5782_), .Y(new_n5783_));
  XOR2X1   g05527(.A(\b[53] ), .B(\b[52] ), .Y(new_n5784_));
  INVX1    g05528(.A(new_n5784_), .Y(new_n5785_));
  XOR2X1   g05529(.A(new_n5785_), .B(new_n5783_), .Y(new_n5786_));
  INVX1    g05530(.A(\b[51] ), .Y(new_n5787_));
  AOI22X1  g05531(.A0(new_n267_), .A1(\b[53] ), .B0(new_n266_), .B1(\b[52] ), .Y(new_n5788_));
  OAI21X1  g05532(.A0(new_n350_), .A1(new_n5787_), .B0(new_n5788_), .Y(new_n5789_));
  AOI21X1  g05533(.A0(new_n5786_), .A1(new_n318_), .B0(new_n5789_), .Y(new_n5790_));
  XOR2X1   g05534(.A(new_n5790_), .B(new_n257_), .Y(new_n5791_));
  AOI21X1  g05535(.A0(new_n5781_), .A1(new_n5766_), .B0(new_n5791_), .Y(new_n5792_));
  AND2X1   g05536(.A(new_n5765_), .B(new_n5612_), .Y(new_n5793_));
  NOR2X1   g05537(.A(new_n5764_), .B(new_n5778_), .Y(new_n5794_));
  AND2X1   g05538(.A(new_n5764_), .B(new_n5778_), .Y(new_n5795_));
  NOR3X1   g05539(.A(new_n5795_), .B(new_n5794_), .C(new_n5612_), .Y(new_n5796_));
  XOR2X1   g05540(.A(new_n5790_), .B(\a[2] ), .Y(new_n5797_));
  NOR3X1   g05541(.A(new_n5797_), .B(new_n5796_), .C(new_n5793_), .Y(new_n5798_));
  OAI22X1  g05542(.A0(new_n5798_), .A1(new_n5792_), .B0(new_n5608_), .B1(new_n5607_), .Y(new_n5799_));
  OR4X1    g05543(.A(new_n5798_), .B(new_n5792_), .C(new_n5608_), .D(new_n5607_), .Y(new_n5800_));
  AND2X1   g05544(.A(new_n5800_), .B(new_n5799_), .Y(\f[53] ));
  OAI21X1  g05545(.A0(new_n5796_), .A1(new_n5793_), .B0(new_n5791_), .Y(new_n5802_));
  AND2X1   g05546(.A(new_n5802_), .B(new_n5799_), .Y(new_n5803_));
  NAND2X1  g05547(.A(\b[53] ), .B(\b[52] ), .Y(new_n5804_));
  OAI21X1  g05548(.A0(new_n5785_), .A1(new_n5783_), .B0(new_n5804_), .Y(new_n5805_));
  XOR2X1   g05549(.A(\b[54] ), .B(\b[53] ), .Y(new_n5806_));
  XOR2X1   g05550(.A(new_n5806_), .B(new_n5805_), .Y(new_n5807_));
  INVX1    g05551(.A(\b[52] ), .Y(new_n5808_));
  AOI22X1  g05552(.A0(new_n267_), .A1(\b[54] ), .B0(new_n266_), .B1(\b[53] ), .Y(new_n5809_));
  OAI21X1  g05553(.A0(new_n350_), .A1(new_n5808_), .B0(new_n5809_), .Y(new_n5810_));
  AOI21X1  g05554(.A0(new_n5807_), .A1(new_n318_), .B0(new_n5810_), .Y(new_n5811_));
  XOR2X1   g05555(.A(new_n5811_), .B(\a[2] ), .Y(new_n5812_));
  OAI21X1  g05556(.A0(new_n5795_), .A1(new_n5769_), .B0(new_n5779_), .Y(new_n5813_));
  AOI22X1  g05557(.A0(new_n603_), .A1(\b[45] ), .B0(new_n602_), .B1(\b[44] ), .Y(new_n5814_));
  OAI21X1  g05558(.A0(new_n601_), .A1(new_n4339_), .B0(new_n5814_), .Y(new_n5815_));
  AOI21X1  g05559(.A0(new_n4338_), .A1(new_n518_), .B0(new_n5815_), .Y(new_n5816_));
  XOR2X1   g05560(.A(new_n5816_), .B(\a[11] ), .Y(new_n5817_));
  OR2X1    g05561(.A(new_n5735_), .B(new_n5731_), .Y(new_n5818_));
  INVX1    g05562(.A(new_n5716_), .Y(new_n5819_));
  XOR2X1   g05563(.A(new_n5819_), .B(new_n5712_), .Y(new_n5820_));
  XOR2X1   g05564(.A(new_n5719_), .B(new_n5820_), .Y(new_n5821_));
  XOR2X1   g05565(.A(new_n5724_), .B(new_n5821_), .Y(new_n5822_));
  XOR2X1   g05566(.A(new_n5730_), .B(new_n5822_), .Y(new_n5823_));
  XOR2X1   g05567(.A(new_n5735_), .B(new_n5823_), .Y(new_n5824_));
  OAI21X1  g05568(.A0(new_n5741_), .A1(new_n5824_), .B0(new_n5818_), .Y(new_n5825_));
  NAND2X1  g05569(.A(new_n5819_), .B(new_n5712_), .Y(new_n5826_));
  OAI21X1  g05570(.A0(new_n5719_), .A1(new_n5717_), .B0(new_n5826_), .Y(new_n5827_));
  AND2X1   g05571(.A(new_n5710_), .B(new_n5620_), .Y(new_n5828_));
  AOI21X1  g05572(.A0(new_n5711_), .A1(new_n5615_), .B0(new_n5828_), .Y(new_n5829_));
  NAND2X1  g05573(.A(new_n5708_), .B(new_n5627_), .Y(new_n5830_));
  NAND2X1  g05574(.A(new_n5709_), .B(new_n5622_), .Y(new_n5831_));
  NAND2X1  g05575(.A(new_n5831_), .B(new_n5830_), .Y(new_n5832_));
  AOI22X1  g05576(.A0(new_n1814_), .A1(\b[30] ), .B0(new_n1813_), .B1(\b[29] ), .Y(new_n5833_));
  OAI21X1  g05577(.A0(new_n1812_), .A1(new_n2231_), .B0(new_n5833_), .Y(new_n5834_));
  AOI21X1  g05578(.A0(new_n2230_), .A1(new_n1617_), .B0(new_n5834_), .Y(new_n5835_));
  XOR2X1   g05579(.A(new_n5835_), .B(\a[26] ), .Y(new_n5836_));
  NOR2X1   g05580(.A(new_n5706_), .B(new_n5702_), .Y(new_n5837_));
  AOI21X1  g05581(.A0(new_n5707_), .A1(new_n5631_), .B0(new_n5837_), .Y(new_n5838_));
  AOI22X1  g05582(.A0(new_n2163_), .A1(\b[27] ), .B0(new_n2162_), .B1(\b[26] ), .Y(new_n5839_));
  OAI21X1  g05583(.A0(new_n2161_), .A1(new_n1880_), .B0(new_n5839_), .Y(new_n5840_));
  AOI21X1  g05584(.A0(new_n1907_), .A1(new_n1879_), .B0(new_n5840_), .Y(new_n5841_));
  XOR2X1   g05585(.A(new_n5841_), .B(\a[29] ), .Y(new_n5842_));
  INVX1    g05586(.A(new_n5638_), .Y(new_n5843_));
  AND2X1   g05587(.A(new_n5700_), .B(new_n5843_), .Y(new_n5844_));
  INVX1    g05588(.A(new_n5701_), .Y(new_n5845_));
  AOI21X1  g05589(.A0(new_n5845_), .A1(new_n5634_), .B0(new_n5844_), .Y(new_n5846_));
  AOI22X1  g05590(.A0(new_n2545_), .A1(\b[24] ), .B0(new_n2544_), .B1(\b[23] ), .Y(new_n5847_));
  OAI21X1  g05591(.A0(new_n2543_), .A1(new_n1479_), .B0(new_n5847_), .Y(new_n5848_));
  AOI21X1  g05592(.A0(new_n2260_), .A1(new_n1572_), .B0(new_n5848_), .Y(new_n5849_));
  XOR2X1   g05593(.A(new_n5849_), .B(\a[32] ), .Y(new_n5850_));
  INVX1    g05594(.A(new_n5693_), .Y(new_n5851_));
  XOR2X1   g05595(.A(new_n5851_), .B(new_n5641_), .Y(new_n5852_));
  OR2X1    g05596(.A(new_n5698_), .B(new_n5852_), .Y(new_n5853_));
  OAI21X1  g05597(.A0(new_n5699_), .A1(new_n5485_), .B0(new_n5853_), .Y(new_n5854_));
  AOI22X1  g05598(.A0(new_n2813_), .A1(\b[21] ), .B0(new_n2812_), .B1(\b[20] ), .Y(new_n5855_));
  OAI21X1  g05599(.A0(new_n2946_), .A1(new_n1300_), .B0(new_n5855_), .Y(new_n5856_));
  AOI21X1  g05600(.A0(new_n2652_), .A1(new_n1299_), .B0(new_n5856_), .Y(new_n5857_));
  XOR2X1   g05601(.A(new_n5857_), .B(\a[35] ), .Y(new_n5858_));
  INVX1    g05602(.A(new_n5858_), .Y(new_n5859_));
  AND2X1   g05603(.A(new_n5692_), .B(new_n5646_), .Y(new_n5860_));
  AOI21X1  g05604(.A0(new_n5693_), .A1(new_n5641_), .B0(new_n5860_), .Y(new_n5861_));
  AOI22X1  g05605(.A0(new_n3204_), .A1(\b[18] ), .B0(new_n3203_), .B1(\b[17] ), .Y(new_n5862_));
  OAI21X1  g05606(.A0(new_n3321_), .A1(new_n974_), .B0(new_n5862_), .Y(new_n5863_));
  AOI21X1  g05607(.A0(new_n3080_), .A1(new_n1042_), .B0(new_n5863_), .Y(new_n5864_));
  XOR2X1   g05608(.A(new_n5864_), .B(\a[38] ), .Y(new_n5865_));
  XOR2X1   g05609(.A(new_n5689_), .B(new_n3478_), .Y(new_n5866_));
  NAND2X1  g05610(.A(new_n5866_), .B(new_n5686_), .Y(new_n5867_));
  OAI21X1  g05611(.A0(new_n5691_), .A1(new_n5649_), .B0(new_n5867_), .Y(new_n5868_));
  AOI22X1  g05612(.A0(new_n3652_), .A1(\b[15] ), .B0(new_n3651_), .B1(\b[14] ), .Y(new_n5869_));
  OAI21X1  g05613(.A0(new_n3778_), .A1(new_n795_), .B0(new_n5869_), .Y(new_n5870_));
  AOI21X1  g05614(.A0(new_n3480_), .A1(new_n794_), .B0(new_n5870_), .Y(new_n5871_));
  XOR2X1   g05615(.A(new_n5871_), .B(\a[41] ), .Y(new_n5872_));
  INVX1    g05616(.A(new_n5872_), .Y(new_n5873_));
  AND2X1   g05617(.A(new_n5684_), .B(new_n5654_), .Y(new_n5874_));
  AOI21X1  g05618(.A0(new_n5685_), .A1(new_n5650_), .B0(new_n5874_), .Y(new_n5875_));
  AOI22X1  g05619(.A0(new_n4095_), .A1(\b[12] ), .B0(new_n4094_), .B1(\b[11] ), .Y(new_n5876_));
  OAI21X1  g05620(.A0(new_n4233_), .A1(new_n587_), .B0(new_n5876_), .Y(new_n5877_));
  AOI21X1  g05621(.A0(new_n3901_), .A1(new_n635_), .B0(new_n5877_), .Y(new_n5878_));
  XOR2X1   g05622(.A(new_n5878_), .B(\a[44] ), .Y(new_n5879_));
  NOR2X1   g05623(.A(new_n5682_), .B(new_n5678_), .Y(new_n5880_));
  AOI21X1  g05624(.A0(new_n5683_), .A1(new_n5657_), .B0(new_n5880_), .Y(new_n5881_));
  AOI22X1  g05625(.A0(new_n4572_), .A1(\b[9] ), .B0(new_n4571_), .B1(\b[8] ), .Y(new_n5882_));
  OAI21X1  g05626(.A0(new_n4740_), .A1(new_n492_), .B0(new_n5882_), .Y(new_n5883_));
  AOI21X1  g05627(.A0(new_n4375_), .A1(new_n491_), .B0(new_n5883_), .Y(new_n5884_));
  XOR2X1   g05628(.A(new_n5884_), .B(\a[47] ), .Y(new_n5885_));
  OR2X1    g05629(.A(new_n5666_), .B(new_n5661_), .Y(new_n5886_));
  XOR2X1   g05630(.A(\a[54] ), .B(\a[53] ), .Y(new_n5887_));
  AND2X1   g05631(.A(new_n5887_), .B(\b[0] ), .Y(new_n5888_));
  XOR2X1   g05632(.A(new_n5888_), .B(new_n5886_), .Y(new_n5889_));
  NOR3X1   g05633(.A(new_n5426_), .B(new_n5424_), .C(new_n5429_), .Y(new_n5890_));
  INVX1    g05634(.A(new_n5890_), .Y(new_n5891_));
  AOI22X1  g05635(.A0(new_n5430_), .A1(\b[3] ), .B0(new_n5427_), .B1(\b[2] ), .Y(new_n5892_));
  OAI21X1  g05636(.A0(new_n5891_), .A1(new_n275_), .B0(new_n5892_), .Y(new_n5893_));
  AOI21X1  g05637(.A0(new_n5425_), .A1(new_n366_), .B0(new_n5893_), .Y(new_n5894_));
  XOR2X1   g05638(.A(new_n5894_), .B(\a[53] ), .Y(new_n5895_));
  XOR2X1   g05639(.A(new_n5895_), .B(new_n5889_), .Y(new_n5896_));
  AOI22X1  g05640(.A0(new_n4880_), .A1(\b[6] ), .B0(new_n4877_), .B1(\b[5] ), .Y(new_n5897_));
  OAI21X1  g05641(.A0(new_n5291_), .A1(new_n325_), .B0(new_n5897_), .Y(new_n5898_));
  AOI21X1  g05642(.A0(new_n4875_), .A1(new_n378_), .B0(new_n5898_), .Y(new_n5899_));
  XOR2X1   g05643(.A(new_n5899_), .B(\a[50] ), .Y(new_n5900_));
  XOR2X1   g05644(.A(new_n5900_), .B(new_n5896_), .Y(new_n5901_));
  XOR2X1   g05645(.A(new_n5901_), .B(new_n5677_), .Y(new_n5902_));
  XOR2X1   g05646(.A(new_n5902_), .B(new_n5885_), .Y(new_n5903_));
  XOR2X1   g05647(.A(new_n5903_), .B(new_n5881_), .Y(new_n5904_));
  XOR2X1   g05648(.A(new_n5904_), .B(new_n5879_), .Y(new_n5905_));
  XOR2X1   g05649(.A(new_n5905_), .B(new_n5875_), .Y(new_n5906_));
  XOR2X1   g05650(.A(new_n5906_), .B(new_n5873_), .Y(new_n5907_));
  XOR2X1   g05651(.A(new_n5907_), .B(new_n5868_), .Y(new_n5908_));
  XOR2X1   g05652(.A(new_n5908_), .B(new_n5865_), .Y(new_n5909_));
  XOR2X1   g05653(.A(new_n5909_), .B(new_n5861_), .Y(new_n5910_));
  XOR2X1   g05654(.A(new_n5910_), .B(new_n5859_), .Y(new_n5911_));
  XOR2X1   g05655(.A(new_n5911_), .B(new_n5854_), .Y(new_n5912_));
  XOR2X1   g05656(.A(new_n5912_), .B(new_n5850_), .Y(new_n5913_));
  XOR2X1   g05657(.A(new_n5913_), .B(new_n5846_), .Y(new_n5914_));
  XOR2X1   g05658(.A(new_n5914_), .B(new_n5842_), .Y(new_n5915_));
  XOR2X1   g05659(.A(new_n5915_), .B(new_n5838_), .Y(new_n5916_));
  XOR2X1   g05660(.A(new_n5916_), .B(new_n5836_), .Y(new_n5917_));
  XOR2X1   g05661(.A(new_n5917_), .B(new_n5832_), .Y(new_n5918_));
  AOI22X1  g05662(.A0(new_n1526_), .A1(\b[33] ), .B0(new_n1525_), .B1(\b[32] ), .Y(new_n5919_));
  OAI21X1  g05663(.A0(new_n1524_), .A1(new_n2615_), .B0(new_n5919_), .Y(new_n5920_));
  AOI21X1  g05664(.A0(new_n2614_), .A1(new_n1347_), .B0(new_n5920_), .Y(new_n5921_));
  XOR2X1   g05665(.A(new_n5921_), .B(\a[23] ), .Y(new_n5922_));
  XOR2X1   g05666(.A(new_n5922_), .B(new_n5918_), .Y(new_n5923_));
  XOR2X1   g05667(.A(new_n5923_), .B(new_n5829_), .Y(new_n5924_));
  AOI22X1  g05668(.A0(new_n1263_), .A1(\b[36] ), .B0(new_n1262_), .B1(\b[35] ), .Y(new_n5925_));
  OAI21X1  g05669(.A0(new_n1261_), .A1(new_n2890_), .B0(new_n5925_), .Y(new_n5926_));
  AOI21X1  g05670(.A0(new_n3015_), .A1(new_n1075_), .B0(new_n5926_), .Y(new_n5927_));
  XOR2X1   g05671(.A(new_n5927_), .B(\a[20] ), .Y(new_n5928_));
  XOR2X1   g05672(.A(new_n5928_), .B(new_n5924_), .Y(new_n5929_));
  XOR2X1   g05673(.A(new_n5929_), .B(new_n5827_), .Y(new_n5930_));
  AOI22X1  g05674(.A0(new_n1017_), .A1(\b[39] ), .B0(new_n1016_), .B1(\b[38] ), .Y(new_n5931_));
  OAI21X1  g05675(.A0(new_n1015_), .A1(new_n3413_), .B0(new_n5931_), .Y(new_n5932_));
  AOI21X1  g05676(.A0(new_n3412_), .A1(new_n882_), .B0(new_n5932_), .Y(new_n5933_));
  XOR2X1   g05677(.A(new_n5933_), .B(\a[17] ), .Y(new_n5934_));
  INVX1    g05678(.A(new_n5934_), .Y(new_n5935_));
  XOR2X1   g05679(.A(new_n5935_), .B(new_n5930_), .Y(new_n5936_));
  NOR2X1   g05680(.A(new_n5724_), .B(new_n5821_), .Y(new_n5937_));
  AOI21X1  g05681(.A0(new_n5730_), .A1(new_n5822_), .B0(new_n5937_), .Y(new_n5938_));
  XOR2X1   g05682(.A(new_n5938_), .B(new_n5936_), .Y(new_n5939_));
  AOI22X1  g05683(.A0(new_n818_), .A1(\b[42] ), .B0(new_n817_), .B1(\b[41] ), .Y(new_n5940_));
  OAI21X1  g05684(.A0(new_n816_), .A1(new_n3720_), .B0(new_n5940_), .Y(new_n5941_));
  AOI21X1  g05685(.A0(new_n3860_), .A1(new_n668_), .B0(new_n5941_), .Y(new_n5942_));
  XOR2X1   g05686(.A(new_n5942_), .B(\a[14] ), .Y(new_n5943_));
  XOR2X1   g05687(.A(new_n5943_), .B(new_n5939_), .Y(new_n5944_));
  XOR2X1   g05688(.A(new_n5944_), .B(new_n5825_), .Y(new_n5945_));
  XOR2X1   g05689(.A(new_n5945_), .B(new_n5817_), .Y(new_n5946_));
  XOR2X1   g05690(.A(new_n5946_), .B(new_n5750_), .Y(new_n5947_));
  AOI22X1  g05691(.A0(new_n469_), .A1(\b[48] ), .B0(new_n468_), .B1(\b[47] ), .Y(new_n5948_));
  OAI21X1  g05692(.A0(new_n467_), .A1(new_n4693_), .B0(new_n5948_), .Y(new_n5949_));
  AOI21X1  g05693(.A0(new_n4692_), .A1(new_n404_), .B0(new_n5949_), .Y(new_n5950_));
  XOR2X1   g05694(.A(new_n5950_), .B(\a[8] ), .Y(new_n5951_));
  XOR2X1   g05695(.A(new_n5951_), .B(new_n5947_), .Y(new_n5952_));
  NOR2X1   g05696(.A(new_n5755_), .B(new_n5776_), .Y(new_n5953_));
  OR2X1    g05697(.A(new_n5573_), .B(new_n5569_), .Y(new_n5954_));
  OAI21X1  g05698(.A0(new_n5579_), .A1(new_n5575_), .B0(new_n5954_), .Y(new_n5955_));
  AOI21X1  g05699(.A0(new_n5955_), .A1(new_n5777_), .B0(new_n5953_), .Y(new_n5956_));
  XOR2X1   g05700(.A(new_n5956_), .B(new_n5952_), .Y(new_n5957_));
  AOI22X1  g05701(.A0(new_n369_), .A1(\b[51] ), .B0(new_n368_), .B1(\b[50] ), .Y(new_n5958_));
  OAI21X1  g05702(.A0(new_n367_), .A1(new_n5237_), .B0(new_n5958_), .Y(new_n5959_));
  AOI21X1  g05703(.A0(new_n5236_), .A1(new_n308_), .B0(new_n5959_), .Y(new_n5960_));
  XOR2X1   g05704(.A(new_n5960_), .B(\a[5] ), .Y(new_n5961_));
  XOR2X1   g05705(.A(new_n5961_), .B(new_n5957_), .Y(new_n5962_));
  XOR2X1   g05706(.A(new_n5962_), .B(new_n5813_), .Y(new_n5963_));
  XOR2X1   g05707(.A(new_n5963_), .B(new_n5812_), .Y(new_n5964_));
  XOR2X1   g05708(.A(new_n5964_), .B(new_n5803_), .Y(\f[54] ));
  INVX1    g05709(.A(new_n5812_), .Y(new_n5966_));
  AND2X1   g05710(.A(new_n5963_), .B(new_n5966_), .Y(new_n5967_));
  AOI21X1  g05711(.A0(new_n5802_), .A1(new_n5799_), .B0(new_n5964_), .Y(new_n5968_));
  OR2X1    g05712(.A(new_n5968_), .B(new_n5967_), .Y(new_n5969_));
  NOR2X1   g05713(.A(new_n5961_), .B(new_n5957_), .Y(new_n5970_));
  AOI21X1  g05714(.A0(new_n5962_), .A1(new_n5813_), .B0(new_n5970_), .Y(new_n5971_));
  OR2X1    g05715(.A(new_n5951_), .B(new_n5947_), .Y(new_n5972_));
  XOR2X1   g05716(.A(new_n5946_), .B(new_n5775_), .Y(new_n5973_));
  XOR2X1   g05717(.A(new_n5951_), .B(new_n5973_), .Y(new_n5974_));
  OAI21X1  g05718(.A0(new_n5956_), .A1(new_n5974_), .B0(new_n5972_), .Y(new_n5975_));
  AOI22X1  g05719(.A0(new_n469_), .A1(\b[49] ), .B0(new_n468_), .B1(\b[48] ), .Y(new_n5976_));
  OAI21X1  g05720(.A0(new_n467_), .A1(new_n5039_), .B0(new_n5976_), .Y(new_n5977_));
  AOI21X1  g05721(.A0(new_n5038_), .A1(new_n404_), .B0(new_n5977_), .Y(new_n5978_));
  XOR2X1   g05722(.A(new_n5978_), .B(new_n400_), .Y(new_n5979_));
  INVX1    g05723(.A(new_n5817_), .Y(new_n5980_));
  NAND2X1  g05724(.A(new_n5945_), .B(new_n5980_), .Y(new_n5981_));
  OAI21X1  g05725(.A0(new_n5946_), .A1(new_n5775_), .B0(new_n5981_), .Y(new_n5982_));
  NOR2X1   g05726(.A(new_n5943_), .B(new_n5939_), .Y(new_n5983_));
  AOI21X1  g05727(.A0(new_n5944_), .A1(new_n5825_), .B0(new_n5983_), .Y(new_n5984_));
  INVX1    g05728(.A(new_n5865_), .Y(new_n5985_));
  NAND2X1  g05729(.A(new_n5908_), .B(new_n5985_), .Y(new_n5986_));
  OAI21X1  g05730(.A0(new_n5909_), .A1(new_n5861_), .B0(new_n5986_), .Y(new_n5987_));
  INVX1    g05731(.A(new_n5879_), .Y(new_n5988_));
  AND2X1   g05732(.A(new_n5904_), .B(new_n5988_), .Y(new_n5989_));
  INVX1    g05733(.A(new_n5989_), .Y(new_n5990_));
  OAI21X1  g05734(.A0(new_n5905_), .A1(new_n5875_), .B0(new_n5990_), .Y(new_n5991_));
  AOI22X1  g05735(.A0(new_n4095_), .A1(\b[13] ), .B0(new_n4094_), .B1(\b[12] ), .Y(new_n5992_));
  OAI21X1  g05736(.A0(new_n4233_), .A1(new_n716_), .B0(new_n5992_), .Y(new_n5993_));
  AOI21X1  g05737(.A0(new_n3901_), .A1(new_n715_), .B0(new_n5993_), .Y(new_n5994_));
  XOR2X1   g05738(.A(new_n5994_), .B(\a[44] ), .Y(new_n5995_));
  INVX1    g05739(.A(new_n5995_), .Y(new_n5996_));
  INVX1    g05740(.A(new_n5885_), .Y(new_n5997_));
  NAND2X1  g05741(.A(new_n5902_), .B(new_n5997_), .Y(new_n5998_));
  OAI21X1  g05742(.A0(new_n5903_), .A1(new_n5881_), .B0(new_n5998_), .Y(new_n5999_));
  AOI22X1  g05743(.A0(new_n4572_), .A1(\b[10] ), .B0(new_n4571_), .B1(\b[9] ), .Y(new_n6000_));
  OAI21X1  g05744(.A0(new_n4740_), .A1(new_n489_), .B0(new_n6000_), .Y(new_n6001_));
  AOI21X1  g05745(.A0(new_n4375_), .A1(new_n543_), .B0(new_n6001_), .Y(new_n6002_));
  XOR2X1   g05746(.A(new_n6002_), .B(new_n4568_), .Y(new_n6003_));
  XOR2X1   g05747(.A(new_n5899_), .B(new_n4873_), .Y(new_n6004_));
  NAND2X1  g05748(.A(new_n6004_), .B(new_n5896_), .Y(new_n6005_));
  OAI21X1  g05749(.A0(new_n5901_), .A1(new_n5677_), .B0(new_n6005_), .Y(new_n6006_));
  AOI22X1  g05750(.A0(new_n4880_), .A1(\b[7] ), .B0(new_n4877_), .B1(\b[6] ), .Y(new_n6007_));
  OAI21X1  g05751(.A0(new_n5291_), .A1(new_n395_), .B0(new_n6007_), .Y(new_n6008_));
  AOI21X1  g05752(.A0(new_n4875_), .A1(new_n394_), .B0(new_n6008_), .Y(new_n6009_));
  XOR2X1   g05753(.A(new_n6009_), .B(new_n4873_), .Y(new_n6010_));
  INVX1    g05754(.A(new_n5888_), .Y(new_n6011_));
  OR4X1    g05755(.A(new_n6011_), .B(new_n5666_), .C(new_n5434_), .D(new_n5422_), .Y(new_n6012_));
  OAI21X1  g05756(.A0(new_n5895_), .A1(new_n5889_), .B0(new_n6012_), .Y(new_n6013_));
  AND2X1   g05757(.A(new_n5425_), .B(new_n323_), .Y(new_n6014_));
  NOR4X1   g05758(.A(new_n5426_), .B(new_n5424_), .C(new_n5429_), .D(new_n277_), .Y(new_n6015_));
  OAI22X1  g05759(.A0(new_n5431_), .A1(new_n325_), .B0(new_n5428_), .B1(new_n297_), .Y(new_n6016_));
  NOR3X1   g05760(.A(new_n6016_), .B(new_n6015_), .C(new_n6014_), .Y(new_n6017_));
  XOR2X1   g05761(.A(new_n6017_), .B(new_n5423_), .Y(new_n6018_));
  INVX1    g05762(.A(\a[56] ), .Y(new_n6019_));
  OR2X1    g05763(.A(new_n5888_), .B(new_n6019_), .Y(new_n6020_));
  INVX1    g05764(.A(new_n5887_), .Y(new_n6021_));
  XOR2X1   g05765(.A(new_n6019_), .B(\a[55] ), .Y(new_n6022_));
  NOR2X1   g05766(.A(new_n6022_), .B(new_n6021_), .Y(new_n6023_));
  XOR2X1   g05767(.A(\a[55] ), .B(\a[54] ), .Y(new_n6024_));
  NAND2X1  g05768(.A(new_n6024_), .B(new_n6021_), .Y(new_n6025_));
  NAND2X1  g05769(.A(new_n6022_), .B(new_n5887_), .Y(new_n6026_));
  OAI22X1  g05770(.A0(new_n6026_), .A1(new_n275_), .B0(new_n6025_), .B1(new_n274_), .Y(new_n6027_));
  AOI21X1  g05771(.A0(new_n6023_), .A1(new_n263_), .B0(new_n6027_), .Y(new_n6028_));
  XOR2X1   g05772(.A(new_n6028_), .B(\a[56] ), .Y(new_n6029_));
  XOR2X1   g05773(.A(new_n6029_), .B(new_n6020_), .Y(new_n6030_));
  XOR2X1   g05774(.A(new_n6030_), .B(new_n6018_), .Y(new_n6031_));
  XOR2X1   g05775(.A(new_n6031_), .B(new_n6013_), .Y(new_n6032_));
  XOR2X1   g05776(.A(new_n6032_), .B(new_n6010_), .Y(new_n6033_));
  XOR2X1   g05777(.A(new_n6033_), .B(new_n6006_), .Y(new_n6034_));
  XOR2X1   g05778(.A(new_n6034_), .B(new_n6003_), .Y(new_n6035_));
  XOR2X1   g05779(.A(new_n6035_), .B(new_n5999_), .Y(new_n6036_));
  XOR2X1   g05780(.A(new_n6036_), .B(new_n5996_), .Y(new_n6037_));
  XOR2X1   g05781(.A(new_n6037_), .B(new_n5991_), .Y(new_n6038_));
  AOI22X1  g05782(.A0(new_n3652_), .A1(\b[16] ), .B0(new_n3651_), .B1(\b[15] ), .Y(new_n6039_));
  OAI21X1  g05783(.A0(new_n3778_), .A1(new_n792_), .B0(new_n6039_), .Y(new_n6040_));
  AOI21X1  g05784(.A0(new_n3480_), .A1(new_n842_), .B0(new_n6040_), .Y(new_n6041_));
  XOR2X1   g05785(.A(new_n6041_), .B(\a[41] ), .Y(new_n6042_));
  XOR2X1   g05786(.A(new_n6042_), .B(new_n6038_), .Y(new_n6043_));
  INVX1    g05787(.A(new_n6043_), .Y(new_n6044_));
  AND2X1   g05788(.A(new_n5906_), .B(new_n5873_), .Y(new_n6045_));
  AOI21X1  g05789(.A0(new_n5907_), .A1(new_n5868_), .B0(new_n6045_), .Y(new_n6046_));
  XOR2X1   g05790(.A(new_n6046_), .B(new_n6044_), .Y(new_n6047_));
  AOI22X1  g05791(.A0(new_n3204_), .A1(\b[19] ), .B0(new_n3203_), .B1(\b[18] ), .Y(new_n6048_));
  OAI21X1  g05792(.A0(new_n3321_), .A1(new_n1118_), .B0(new_n6048_), .Y(new_n6049_));
  AOI21X1  g05793(.A0(new_n3080_), .A1(new_n1117_), .B0(new_n6049_), .Y(new_n6050_));
  XOR2X1   g05794(.A(new_n6050_), .B(\a[38] ), .Y(new_n6051_));
  NAND2X1  g05795(.A(new_n6051_), .B(new_n6047_), .Y(new_n6052_));
  XOR2X1   g05796(.A(new_n6051_), .B(new_n6047_), .Y(new_n6053_));
  INVX1    g05797(.A(new_n6053_), .Y(new_n6054_));
  NOR2X1   g05798(.A(new_n6051_), .B(new_n6047_), .Y(new_n6055_));
  AOI21X1  g05799(.A0(new_n6052_), .A1(new_n5987_), .B0(new_n6055_), .Y(new_n6056_));
  AOI22X1  g05800(.A0(new_n6056_), .A1(new_n6052_), .B0(new_n6054_), .B1(new_n5987_), .Y(new_n6057_));
  AOI22X1  g05801(.A0(new_n2813_), .A1(\b[22] ), .B0(new_n2812_), .B1(\b[21] ), .Y(new_n6058_));
  OAI21X1  g05802(.A0(new_n2946_), .A1(new_n1297_), .B0(new_n6058_), .Y(new_n6059_));
  AOI21X1  g05803(.A0(new_n2652_), .A1(new_n1399_), .B0(new_n6059_), .Y(new_n6060_));
  XOR2X1   g05804(.A(new_n6060_), .B(\a[35] ), .Y(new_n6061_));
  XOR2X1   g05805(.A(new_n6061_), .B(new_n6057_), .Y(new_n6062_));
  AND2X1   g05806(.A(new_n5910_), .B(new_n5859_), .Y(new_n6063_));
  AOI21X1  g05807(.A0(new_n5911_), .A1(new_n5854_), .B0(new_n6063_), .Y(new_n6064_));
  XOR2X1   g05808(.A(new_n6064_), .B(new_n6062_), .Y(new_n6065_));
  AOI22X1  g05809(.A0(new_n2545_), .A1(\b[25] ), .B0(new_n2544_), .B1(\b[24] ), .Y(new_n6066_));
  OAI21X1  g05810(.A0(new_n2543_), .A1(new_n1591_), .B0(new_n6066_), .Y(new_n6067_));
  AOI21X1  g05811(.A0(new_n2260_), .A1(new_n1590_), .B0(new_n6067_), .Y(new_n6068_));
  XOR2X1   g05812(.A(new_n6068_), .B(\a[32] ), .Y(new_n6069_));
  XOR2X1   g05813(.A(new_n6069_), .B(new_n6065_), .Y(new_n6070_));
  INVX1    g05814(.A(new_n6070_), .Y(new_n6071_));
  INVX1    g05815(.A(new_n5850_), .Y(new_n6072_));
  NAND2X1  g05816(.A(new_n5912_), .B(new_n6072_), .Y(new_n6073_));
  OAI21X1  g05817(.A0(new_n5913_), .A1(new_n5846_), .B0(new_n6073_), .Y(new_n6074_));
  XOR2X1   g05818(.A(new_n6074_), .B(new_n6071_), .Y(new_n6075_));
  AOI22X1  g05819(.A0(new_n2163_), .A1(\b[28] ), .B0(new_n2162_), .B1(\b[27] ), .Y(new_n6076_));
  OAI21X1  g05820(.A0(new_n2161_), .A1(new_n1877_), .B0(new_n6076_), .Y(new_n6077_));
  AOI21X1  g05821(.A0(new_n2004_), .A1(new_n1907_), .B0(new_n6077_), .Y(new_n6078_));
  XOR2X1   g05822(.A(new_n6078_), .B(\a[29] ), .Y(new_n6079_));
  XOR2X1   g05823(.A(new_n6079_), .B(new_n6075_), .Y(new_n6080_));
  INVX1    g05824(.A(new_n5842_), .Y(new_n6081_));
  NAND2X1  g05825(.A(new_n5914_), .B(new_n6081_), .Y(new_n6082_));
  OAI21X1  g05826(.A0(new_n5915_), .A1(new_n5838_), .B0(new_n6082_), .Y(new_n6083_));
  XOR2X1   g05827(.A(new_n6083_), .B(new_n6080_), .Y(new_n6084_));
  AOI22X1  g05828(.A0(new_n1814_), .A1(\b[31] ), .B0(new_n1813_), .B1(\b[30] ), .Y(new_n6085_));
  OAI21X1  g05829(.A0(new_n1812_), .A1(new_n2359_), .B0(new_n6085_), .Y(new_n6086_));
  AOI21X1  g05830(.A0(new_n2358_), .A1(new_n1617_), .B0(new_n6086_), .Y(new_n6087_));
  XOR2X1   g05831(.A(new_n6087_), .B(\a[26] ), .Y(new_n6088_));
  XOR2X1   g05832(.A(new_n6088_), .B(new_n6084_), .Y(new_n6089_));
  INVX1    g05833(.A(new_n6089_), .Y(new_n6090_));
  INVX1    g05834(.A(new_n5836_), .Y(new_n6091_));
  AOI21X1  g05835(.A0(new_n5831_), .A1(new_n5830_), .B0(new_n5917_), .Y(new_n6092_));
  AOI21X1  g05836(.A0(new_n5916_), .A1(new_n6091_), .B0(new_n6092_), .Y(new_n6093_));
  XOR2X1   g05837(.A(new_n6093_), .B(new_n6090_), .Y(new_n6094_));
  AOI22X1  g05838(.A0(new_n1526_), .A1(\b[34] ), .B0(new_n1525_), .B1(\b[33] ), .Y(new_n6095_));
  OAI21X1  g05839(.A0(new_n1524_), .A1(new_n2612_), .B0(new_n6095_), .Y(new_n6096_));
  AOI21X1  g05840(.A0(new_n2759_), .A1(new_n1347_), .B0(new_n6096_), .Y(new_n6097_));
  XOR2X1   g05841(.A(new_n6097_), .B(\a[23] ), .Y(new_n6098_));
  XOR2X1   g05842(.A(new_n6098_), .B(new_n6094_), .Y(new_n6099_));
  OR2X1    g05843(.A(new_n5922_), .B(new_n5918_), .Y(new_n6100_));
  XOR2X1   g05844(.A(new_n5921_), .B(new_n1351_), .Y(new_n6101_));
  XOR2X1   g05845(.A(new_n6101_), .B(new_n5918_), .Y(new_n6102_));
  OAI21X1  g05846(.A0(new_n6102_), .A1(new_n5829_), .B0(new_n6100_), .Y(new_n6103_));
  XOR2X1   g05847(.A(new_n6103_), .B(new_n6099_), .Y(new_n6104_));
  AOI22X1  g05848(.A0(new_n1263_), .A1(\b[37] ), .B0(new_n1262_), .B1(\b[36] ), .Y(new_n6105_));
  OAI21X1  g05849(.A0(new_n1261_), .A1(new_n3156_), .B0(new_n6105_), .Y(new_n6106_));
  AOI21X1  g05850(.A0(new_n3155_), .A1(new_n1075_), .B0(new_n6106_), .Y(new_n6107_));
  XOR2X1   g05851(.A(new_n6107_), .B(\a[20] ), .Y(new_n6108_));
  XOR2X1   g05852(.A(new_n6108_), .B(new_n6104_), .Y(new_n6109_));
  NOR2X1   g05853(.A(new_n5928_), .B(new_n5924_), .Y(new_n6110_));
  AOI21X1  g05854(.A0(new_n5929_), .A1(new_n5827_), .B0(new_n6110_), .Y(new_n6111_));
  XOR2X1   g05855(.A(new_n6111_), .B(new_n6109_), .Y(new_n6112_));
  AOI22X1  g05856(.A0(new_n1017_), .A1(\b[40] ), .B0(new_n1016_), .B1(\b[39] ), .Y(new_n6113_));
  OAI21X1  g05857(.A0(new_n1015_), .A1(new_n3575_), .B0(new_n6113_), .Y(new_n6114_));
  AOI21X1  g05858(.A0(new_n3574_), .A1(new_n882_), .B0(new_n6114_), .Y(new_n6115_));
  XOR2X1   g05859(.A(new_n6115_), .B(\a[17] ), .Y(new_n6116_));
  XOR2X1   g05860(.A(new_n6116_), .B(new_n6112_), .Y(new_n6117_));
  NAND2X1  g05861(.A(new_n5935_), .B(new_n5930_), .Y(new_n6118_));
  XOR2X1   g05862(.A(new_n5934_), .B(new_n5930_), .Y(new_n6119_));
  OAI21X1  g05863(.A0(new_n5938_), .A1(new_n6119_), .B0(new_n6118_), .Y(new_n6120_));
  XOR2X1   g05864(.A(new_n6120_), .B(new_n6117_), .Y(new_n6121_));
  AOI22X1  g05865(.A0(new_n818_), .A1(\b[43] ), .B0(new_n817_), .B1(\b[42] ), .Y(new_n6122_));
  OAI21X1  g05866(.A0(new_n816_), .A1(new_n4015_), .B0(new_n6122_), .Y(new_n6123_));
  AOI21X1  g05867(.A0(new_n4014_), .A1(new_n668_), .B0(new_n6123_), .Y(new_n6124_));
  XOR2X1   g05868(.A(new_n6124_), .B(\a[14] ), .Y(new_n6125_));
  AND2X1   g05869(.A(new_n6125_), .B(new_n6121_), .Y(new_n6126_));
  XOR2X1   g05870(.A(new_n6125_), .B(new_n6121_), .Y(new_n6127_));
  OR2X1    g05871(.A(new_n6125_), .B(new_n6121_), .Y(new_n6128_));
  OAI21X1  g05872(.A0(new_n6126_), .A1(new_n5984_), .B0(new_n6128_), .Y(new_n6129_));
  OAI22X1  g05873(.A0(new_n6129_), .A1(new_n6126_), .B0(new_n6127_), .B1(new_n5984_), .Y(new_n6130_));
  AOI22X1  g05874(.A0(new_n603_), .A1(\b[46] ), .B0(new_n602_), .B1(\b[45] ), .Y(new_n6131_));
  OAI21X1  g05875(.A0(new_n601_), .A1(new_n4336_), .B0(new_n6131_), .Y(new_n6132_));
  AOI21X1  g05876(.A0(new_n4509_), .A1(new_n518_), .B0(new_n6132_), .Y(new_n6133_));
  XOR2X1   g05877(.A(new_n6133_), .B(new_n515_), .Y(new_n6134_));
  XOR2X1   g05878(.A(new_n6134_), .B(new_n6130_), .Y(new_n6135_));
  XOR2X1   g05879(.A(new_n6135_), .B(new_n5982_), .Y(new_n6136_));
  XOR2X1   g05880(.A(new_n6136_), .B(new_n5979_), .Y(new_n6137_));
  XOR2X1   g05881(.A(new_n6137_), .B(new_n5975_), .Y(new_n6138_));
  AOI22X1  g05882(.A0(new_n369_), .A1(\b[52] ), .B0(new_n368_), .B1(\b[51] ), .Y(new_n6139_));
  OAI21X1  g05883(.A0(new_n367_), .A1(new_n5234_), .B0(new_n6139_), .Y(new_n6140_));
  AOI21X1  g05884(.A0(new_n5590_), .A1(new_n308_), .B0(new_n6140_), .Y(new_n6141_));
  XOR2X1   g05885(.A(new_n6141_), .B(\a[5] ), .Y(new_n6142_));
  INVX1    g05886(.A(new_n6142_), .Y(new_n6143_));
  XOR2X1   g05887(.A(new_n6143_), .B(new_n6138_), .Y(new_n6144_));
  XOR2X1   g05888(.A(new_n6144_), .B(new_n5971_), .Y(new_n6145_));
  AND2X1   g05889(.A(\b[54] ), .B(\b[53] ), .Y(new_n6146_));
  AOI21X1  g05890(.A0(new_n5806_), .A1(new_n5805_), .B0(new_n6146_), .Y(new_n6147_));
  INVX1    g05891(.A(\b[54] ), .Y(new_n6148_));
  XOR2X1   g05892(.A(\b[55] ), .B(new_n6148_), .Y(new_n6149_));
  XOR2X1   g05893(.A(new_n6149_), .B(new_n6147_), .Y(new_n6150_));
  INVX1    g05894(.A(\b[53] ), .Y(new_n6151_));
  AOI22X1  g05895(.A0(new_n267_), .A1(\b[55] ), .B0(new_n266_), .B1(\b[54] ), .Y(new_n6152_));
  OAI21X1  g05896(.A0(new_n350_), .A1(new_n6151_), .B0(new_n6152_), .Y(new_n6153_));
  AOI21X1  g05897(.A0(new_n6150_), .A1(new_n318_), .B0(new_n6153_), .Y(new_n6154_));
  XOR2X1   g05898(.A(new_n6154_), .B(\a[2] ), .Y(new_n6155_));
  XOR2X1   g05899(.A(new_n6155_), .B(new_n6145_), .Y(new_n6156_));
  XOR2X1   g05900(.A(new_n6156_), .B(new_n5969_), .Y(\f[55] ));
  NAND2X1  g05901(.A(new_n6143_), .B(new_n6138_), .Y(new_n6158_));
  XOR2X1   g05902(.A(new_n6142_), .B(new_n6138_), .Y(new_n6159_));
  OAI21X1  g05903(.A0(new_n6159_), .A1(new_n5971_), .B0(new_n6158_), .Y(new_n6160_));
  NOR2X1   g05904(.A(new_n5951_), .B(new_n5947_), .Y(new_n6161_));
  OR2X1    g05905(.A(new_n5755_), .B(new_n5776_), .Y(new_n6162_));
  OAI21X1  g05906(.A0(new_n5759_), .A1(new_n5756_), .B0(new_n6162_), .Y(new_n6163_));
  AOI21X1  g05907(.A0(new_n6163_), .A1(new_n5952_), .B0(new_n6161_), .Y(new_n6164_));
  NOR2X1   g05908(.A(new_n6136_), .B(new_n5979_), .Y(new_n6165_));
  NAND2X1  g05909(.A(new_n6136_), .B(new_n5979_), .Y(new_n6166_));
  OAI21X1  g05910(.A0(new_n6165_), .A1(new_n6164_), .B0(new_n6166_), .Y(new_n6167_));
  AOI22X1  g05911(.A0(new_n469_), .A1(\b[50] ), .B0(new_n468_), .B1(\b[49] ), .Y(new_n6168_));
  OAI21X1  g05912(.A0(new_n467_), .A1(new_n5036_), .B0(new_n6168_), .Y(new_n6169_));
  AOI21X1  g05913(.A0(new_n5204_), .A1(new_n404_), .B0(new_n6169_), .Y(new_n6170_));
  XOR2X1   g05914(.A(new_n6170_), .B(\a[8] ), .Y(new_n6171_));
  INVX1    g05915(.A(new_n6171_), .Y(new_n6172_));
  AND2X1   g05916(.A(new_n6134_), .B(new_n6130_), .Y(new_n6173_));
  AOI21X1  g05917(.A0(new_n6135_), .A1(new_n5982_), .B0(new_n6173_), .Y(new_n6174_));
  INVX1    g05918(.A(new_n6084_), .Y(new_n6175_));
  OR2X1    g05919(.A(new_n6088_), .B(new_n6175_), .Y(new_n6176_));
  OAI21X1  g05920(.A0(new_n6093_), .A1(new_n6089_), .B0(new_n6176_), .Y(new_n6177_));
  AOI22X1  g05921(.A0(new_n1814_), .A1(\b[32] ), .B0(new_n1813_), .B1(\b[31] ), .Y(new_n6178_));
  OAI21X1  g05922(.A0(new_n1812_), .A1(new_n2356_), .B0(new_n6178_), .Y(new_n6179_));
  AOI21X1  g05923(.A0(new_n2495_), .A1(new_n1617_), .B0(new_n6179_), .Y(new_n6180_));
  XOR2X1   g05924(.A(new_n6180_), .B(\a[26] ), .Y(new_n6181_));
  INVX1    g05925(.A(new_n6181_), .Y(new_n6182_));
  NAND2X1  g05926(.A(new_n6083_), .B(new_n6080_), .Y(new_n6183_));
  OAI21X1  g05927(.A0(new_n6079_), .A1(new_n6075_), .B0(new_n6183_), .Y(new_n6184_));
  OR2X1    g05928(.A(new_n6061_), .B(new_n6057_), .Y(new_n6185_));
  INVX1    g05929(.A(new_n6061_), .Y(new_n6186_));
  XOR2X1   g05930(.A(new_n6186_), .B(new_n6057_), .Y(new_n6187_));
  OAI21X1  g05931(.A0(new_n6064_), .A1(new_n6187_), .B0(new_n6185_), .Y(new_n6188_));
  XOR2X1   g05932(.A(new_n6041_), .B(new_n3478_), .Y(new_n6189_));
  NAND2X1  g05933(.A(new_n6189_), .B(new_n6038_), .Y(new_n6190_));
  OAI21X1  g05934(.A0(new_n6046_), .A1(new_n6043_), .B0(new_n6190_), .Y(new_n6191_));
  AOI22X1  g05935(.A0(new_n3652_), .A1(\b[17] ), .B0(new_n3651_), .B1(\b[16] ), .Y(new_n6192_));
  OAI21X1  g05936(.A0(new_n3778_), .A1(new_n977_), .B0(new_n6192_), .Y(new_n6193_));
  AOI21X1  g05937(.A0(new_n3480_), .A1(new_n976_), .B0(new_n6193_), .Y(new_n6194_));
  XOR2X1   g05938(.A(new_n6194_), .B(\a[41] ), .Y(new_n6195_));
  AND2X1   g05939(.A(new_n6036_), .B(new_n5996_), .Y(new_n6196_));
  AOI21X1  g05940(.A0(new_n6037_), .A1(new_n5991_), .B0(new_n6196_), .Y(new_n6197_));
  AND2X1   g05941(.A(new_n6034_), .B(new_n6003_), .Y(new_n6198_));
  AOI21X1  g05942(.A0(new_n6035_), .A1(new_n5999_), .B0(new_n6198_), .Y(new_n6199_));
  AOI22X1  g05943(.A0(new_n4572_), .A1(\b[11] ), .B0(new_n4571_), .B1(\b[10] ), .Y(new_n6200_));
  OAI21X1  g05944(.A0(new_n4740_), .A1(new_n590_), .B0(new_n6200_), .Y(new_n6201_));
  AOI21X1  g05945(.A0(new_n4375_), .A1(new_n589_), .B0(new_n6201_), .Y(new_n6202_));
  XOR2X1   g05946(.A(new_n6202_), .B(\a[47] ), .Y(new_n6203_));
  INVX1    g05947(.A(new_n6203_), .Y(new_n6204_));
  AND2X1   g05948(.A(new_n6032_), .B(new_n6010_), .Y(new_n6205_));
  AND2X1   g05949(.A(new_n6033_), .B(new_n6006_), .Y(new_n6206_));
  OR2X1    g05950(.A(new_n6206_), .B(new_n6205_), .Y(new_n6207_));
  AND2X1   g05951(.A(new_n6030_), .B(new_n6018_), .Y(new_n6208_));
  AND2X1   g05952(.A(new_n6031_), .B(new_n6013_), .Y(new_n6209_));
  OR2X1    g05953(.A(new_n6209_), .B(new_n6208_), .Y(new_n6210_));
  NAND3X1  g05954(.A(new_n6028_), .B(new_n6011_), .C(\a[56] ), .Y(new_n6211_));
  NAND2X1  g05955(.A(new_n6023_), .B(new_n341_), .Y(new_n6212_));
  OR2X1    g05956(.A(new_n6024_), .B(new_n5887_), .Y(new_n6213_));
  NOR2X1   g05957(.A(new_n6213_), .B(new_n6022_), .Y(new_n6214_));
  OAI22X1  g05958(.A0(new_n6026_), .A1(new_n277_), .B0(new_n6025_), .B1(new_n275_), .Y(new_n6215_));
  AOI21X1  g05959(.A0(new_n6214_), .A1(\b[0] ), .B0(new_n6215_), .Y(new_n6216_));
  NAND2X1  g05960(.A(new_n6216_), .B(new_n6212_), .Y(new_n6217_));
  XOR2X1   g05961(.A(new_n6217_), .B(new_n6019_), .Y(new_n6218_));
  XOR2X1   g05962(.A(new_n6218_), .B(new_n6211_), .Y(new_n6219_));
  INVX1    g05963(.A(new_n6219_), .Y(new_n6220_));
  AOI22X1  g05964(.A0(new_n5430_), .A1(\b[5] ), .B0(new_n5427_), .B1(\b[4] ), .Y(new_n6221_));
  OAI21X1  g05965(.A0(new_n5891_), .A1(new_n297_), .B0(new_n6221_), .Y(new_n6222_));
  AOI21X1  g05966(.A0(new_n5425_), .A1(new_n349_), .B0(new_n6222_), .Y(new_n6223_));
  XOR2X1   g05967(.A(new_n6223_), .B(\a[53] ), .Y(new_n6224_));
  NAND2X1  g05968(.A(new_n6224_), .B(new_n6220_), .Y(new_n6225_));
  NOR2X1   g05969(.A(new_n6224_), .B(new_n6220_), .Y(new_n6226_));
  INVX1    g05970(.A(new_n6226_), .Y(new_n6227_));
  NAND3X1  g05971(.A(new_n6225_), .B(new_n6227_), .C(new_n6210_), .Y(new_n6228_));
  AOI21X1  g05972(.A0(new_n6225_), .A1(new_n6210_), .B0(new_n6226_), .Y(new_n6229_));
  AOI22X1  g05973(.A0(new_n6229_), .A1(new_n6225_), .B0(new_n6228_), .B1(new_n6210_), .Y(new_n6230_));
  AOI22X1  g05974(.A0(new_n4880_), .A1(\b[8] ), .B0(new_n4877_), .B1(\b[7] ), .Y(new_n6231_));
  OAI21X1  g05975(.A0(new_n5291_), .A1(new_n392_), .B0(new_n6231_), .Y(new_n6232_));
  AOI21X1  g05976(.A0(new_n4875_), .A1(new_n454_), .B0(new_n6232_), .Y(new_n6233_));
  XOR2X1   g05977(.A(new_n6233_), .B(\a[50] ), .Y(new_n6234_));
  XOR2X1   g05978(.A(new_n6234_), .B(new_n6230_), .Y(new_n6235_));
  XOR2X1   g05979(.A(new_n6235_), .B(new_n6207_), .Y(new_n6236_));
  XOR2X1   g05980(.A(new_n6236_), .B(new_n6204_), .Y(new_n6237_));
  INVX1    g05981(.A(new_n6237_), .Y(new_n6238_));
  XOR2X1   g05982(.A(new_n6238_), .B(new_n6199_), .Y(new_n6239_));
  AOI22X1  g05983(.A0(new_n4095_), .A1(\b[14] ), .B0(new_n4094_), .B1(\b[13] ), .Y(new_n6240_));
  OAI21X1  g05984(.A0(new_n4233_), .A1(new_n713_), .B0(new_n6240_), .Y(new_n6241_));
  AOI21X1  g05985(.A0(new_n3901_), .A1(new_n734_), .B0(new_n6241_), .Y(new_n6242_));
  XOR2X1   g05986(.A(new_n6242_), .B(\a[44] ), .Y(new_n6243_));
  XOR2X1   g05987(.A(new_n6243_), .B(new_n6239_), .Y(new_n6244_));
  XOR2X1   g05988(.A(new_n6244_), .B(new_n6197_), .Y(new_n6245_));
  XOR2X1   g05989(.A(new_n6245_), .B(new_n6195_), .Y(new_n6246_));
  XOR2X1   g05990(.A(new_n6246_), .B(new_n6191_), .Y(new_n6247_));
  AOI22X1  g05991(.A0(new_n3204_), .A1(\b[20] ), .B0(new_n3203_), .B1(\b[19] ), .Y(new_n6248_));
  OAI21X1  g05992(.A0(new_n3321_), .A1(new_n1115_), .B0(new_n6248_), .Y(new_n6249_));
  AOI21X1  g05993(.A0(new_n3080_), .A1(new_n1217_), .B0(new_n6249_), .Y(new_n6250_));
  XOR2X1   g05994(.A(new_n6250_), .B(\a[38] ), .Y(new_n6251_));
  INVX1    g05995(.A(new_n6251_), .Y(new_n6252_));
  XOR2X1   g05996(.A(new_n6252_), .B(new_n6247_), .Y(new_n6253_));
  INVX1    g05997(.A(new_n6253_), .Y(new_n6254_));
  XOR2X1   g05998(.A(new_n6254_), .B(new_n6056_), .Y(new_n6255_));
  AOI22X1  g05999(.A0(new_n2813_), .A1(\b[23] ), .B0(new_n2812_), .B1(\b[22] ), .Y(new_n6256_));
  OAI21X1  g06000(.A0(new_n2946_), .A1(new_n1482_), .B0(new_n6256_), .Y(new_n6257_));
  AOI21X1  g06001(.A0(new_n2652_), .A1(new_n1481_), .B0(new_n6257_), .Y(new_n6258_));
  XOR2X1   g06002(.A(new_n6258_), .B(\a[35] ), .Y(new_n6259_));
  XOR2X1   g06003(.A(new_n6259_), .B(new_n6255_), .Y(new_n6260_));
  XOR2X1   g06004(.A(new_n6260_), .B(new_n6188_), .Y(new_n6261_));
  AOI22X1  g06005(.A0(new_n2545_), .A1(\b[26] ), .B0(new_n2544_), .B1(\b[25] ), .Y(new_n6262_));
  OAI21X1  g06006(.A0(new_n2543_), .A1(new_n1588_), .B0(new_n6262_), .Y(new_n6263_));
  AOI21X1  g06007(.A0(new_n2260_), .A1(new_n1783_), .B0(new_n6263_), .Y(new_n6264_));
  XOR2X1   g06008(.A(new_n6264_), .B(\a[32] ), .Y(new_n6265_));
  INVX1    g06009(.A(new_n6265_), .Y(new_n6266_));
  OR2X1    g06010(.A(new_n6266_), .B(new_n6261_), .Y(new_n6267_));
  NOR2X1   g06011(.A(new_n6069_), .B(new_n6065_), .Y(new_n6268_));
  AOI21X1  g06012(.A0(new_n6074_), .A1(new_n6070_), .B0(new_n6268_), .Y(new_n6269_));
  NAND2X1  g06013(.A(new_n6266_), .B(new_n6261_), .Y(new_n6270_));
  AOI21X1  g06014(.A0(new_n6267_), .A1(new_n6270_), .B0(new_n6269_), .Y(new_n6271_));
  XOR2X1   g06015(.A(new_n6265_), .B(new_n6261_), .Y(new_n6272_));
  OR2X1    g06016(.A(new_n6272_), .B(new_n6269_), .Y(new_n6273_));
  AND2X1   g06017(.A(new_n6273_), .B(new_n6270_), .Y(new_n6274_));
  AOI21X1  g06018(.A0(new_n6274_), .A1(new_n6267_), .B0(new_n6271_), .Y(new_n6275_));
  AOI22X1  g06019(.A0(new_n2163_), .A1(\b[29] ), .B0(new_n2162_), .B1(\b[28] ), .Y(new_n6276_));
  OAI21X1  g06020(.A0(new_n2161_), .A1(new_n2126_), .B0(new_n6276_), .Y(new_n6277_));
  AOI21X1  g06021(.A0(new_n2125_), .A1(new_n1907_), .B0(new_n6277_), .Y(new_n6278_));
  XOR2X1   g06022(.A(new_n6278_), .B(\a[29] ), .Y(new_n6279_));
  XOR2X1   g06023(.A(new_n6279_), .B(new_n6275_), .Y(new_n6280_));
  XOR2X1   g06024(.A(new_n6280_), .B(new_n6184_), .Y(new_n6281_));
  XOR2X1   g06025(.A(new_n6281_), .B(new_n6182_), .Y(new_n6282_));
  XOR2X1   g06026(.A(new_n6282_), .B(new_n6177_), .Y(new_n6283_));
  AOI22X1  g06027(.A0(new_n1526_), .A1(\b[35] ), .B0(new_n1525_), .B1(\b[34] ), .Y(new_n6284_));
  OAI21X1  g06028(.A0(new_n1524_), .A1(new_n2893_), .B0(new_n6284_), .Y(new_n6285_));
  AOI21X1  g06029(.A0(new_n2892_), .A1(new_n1347_), .B0(new_n6285_), .Y(new_n6286_));
  XOR2X1   g06030(.A(new_n6286_), .B(\a[23] ), .Y(new_n6287_));
  XOR2X1   g06031(.A(new_n6287_), .B(new_n6283_), .Y(new_n6288_));
  NOR2X1   g06032(.A(new_n6098_), .B(new_n6094_), .Y(new_n6289_));
  AOI21X1  g06033(.A0(new_n6103_), .A1(new_n6099_), .B0(new_n6289_), .Y(new_n6290_));
  XOR2X1   g06034(.A(new_n6290_), .B(new_n6288_), .Y(new_n6291_));
  AOI22X1  g06035(.A0(new_n1263_), .A1(\b[38] ), .B0(new_n1262_), .B1(\b[37] ), .Y(new_n6292_));
  OAI21X1  g06036(.A0(new_n1261_), .A1(new_n3276_), .B0(new_n6292_), .Y(new_n6293_));
  AOI21X1  g06037(.A0(new_n3275_), .A1(new_n1075_), .B0(new_n6293_), .Y(new_n6294_));
  XOR2X1   g06038(.A(new_n6294_), .B(\a[20] ), .Y(new_n6295_));
  XOR2X1   g06039(.A(new_n6295_), .B(new_n6291_), .Y(new_n6296_));
  XOR2X1   g06040(.A(new_n6093_), .B(new_n6089_), .Y(new_n6297_));
  XOR2X1   g06041(.A(new_n6098_), .B(new_n6297_), .Y(new_n6298_));
  XOR2X1   g06042(.A(new_n6103_), .B(new_n6298_), .Y(new_n6299_));
  OR2X1    g06043(.A(new_n6108_), .B(new_n6299_), .Y(new_n6300_));
  OAI21X1  g06044(.A0(new_n6111_), .A1(new_n6109_), .B0(new_n6300_), .Y(new_n6301_));
  XOR2X1   g06045(.A(new_n6301_), .B(new_n6296_), .Y(new_n6302_));
  AOI22X1  g06046(.A0(new_n1017_), .A1(\b[41] ), .B0(new_n1016_), .B1(\b[40] ), .Y(new_n6303_));
  OAI21X1  g06047(.A0(new_n1015_), .A1(new_n3723_), .B0(new_n6303_), .Y(new_n6304_));
  AOI21X1  g06048(.A0(new_n3722_), .A1(new_n882_), .B0(new_n6304_), .Y(new_n6305_));
  XOR2X1   g06049(.A(new_n6305_), .B(\a[17] ), .Y(new_n6306_));
  XOR2X1   g06050(.A(new_n6306_), .B(new_n6302_), .Y(new_n6307_));
  XOR2X1   g06051(.A(new_n6108_), .B(new_n6299_), .Y(new_n6308_));
  XOR2X1   g06052(.A(new_n6111_), .B(new_n6308_), .Y(new_n6309_));
  NOR2X1   g06053(.A(new_n6116_), .B(new_n6309_), .Y(new_n6310_));
  XOR2X1   g06054(.A(new_n6116_), .B(new_n6309_), .Y(new_n6311_));
  AOI21X1  g06055(.A0(new_n6120_), .A1(new_n6311_), .B0(new_n6310_), .Y(new_n6312_));
  XOR2X1   g06056(.A(new_n6312_), .B(new_n6307_), .Y(new_n6313_));
  AOI22X1  g06057(.A0(new_n818_), .A1(\b[44] ), .B0(new_n817_), .B1(\b[43] ), .Y(new_n6314_));
  OAI21X1  g06058(.A0(new_n816_), .A1(new_n4012_), .B0(new_n6314_), .Y(new_n6315_));
  AOI21X1  g06059(.A0(new_n4178_), .A1(new_n668_), .B0(new_n6315_), .Y(new_n6316_));
  XOR2X1   g06060(.A(new_n6316_), .B(\a[14] ), .Y(new_n6317_));
  NOR2X1   g06061(.A(new_n6317_), .B(new_n6313_), .Y(new_n6318_));
  AND2X1   g06062(.A(new_n6317_), .B(new_n6313_), .Y(new_n6319_));
  OR2X1    g06063(.A(new_n6319_), .B(new_n6318_), .Y(new_n6320_));
  AND2X1   g06064(.A(new_n6320_), .B(new_n6129_), .Y(new_n6321_));
  NOR3X1   g06065(.A(new_n6319_), .B(new_n6318_), .C(new_n6129_), .Y(new_n6322_));
  OR2X1    g06066(.A(new_n6322_), .B(new_n6321_), .Y(new_n6323_));
  AOI22X1  g06067(.A0(new_n603_), .A1(\b[47] ), .B0(new_n602_), .B1(\b[46] ), .Y(new_n6324_));
  OAI21X1  g06068(.A0(new_n601_), .A1(new_n4674_), .B0(new_n6324_), .Y(new_n6325_));
  AOI21X1  g06069(.A0(new_n4673_), .A1(new_n518_), .B0(new_n6325_), .Y(new_n6326_));
  XOR2X1   g06070(.A(new_n6326_), .B(\a[11] ), .Y(new_n6327_));
  XOR2X1   g06071(.A(new_n6327_), .B(new_n6323_), .Y(new_n6328_));
  XOR2X1   g06072(.A(new_n6328_), .B(new_n6174_), .Y(new_n6329_));
  XOR2X1   g06073(.A(new_n6329_), .B(new_n6172_), .Y(new_n6330_));
  XOR2X1   g06074(.A(new_n6330_), .B(new_n6167_), .Y(new_n6331_));
  AOI22X1  g06075(.A0(new_n369_), .A1(\b[53] ), .B0(new_n368_), .B1(\b[52] ), .Y(new_n6332_));
  OAI21X1  g06076(.A0(new_n367_), .A1(new_n5787_), .B0(new_n6332_), .Y(new_n6333_));
  AOI21X1  g06077(.A0(new_n5786_), .A1(new_n308_), .B0(new_n6333_), .Y(new_n6334_));
  XOR2X1   g06078(.A(new_n6334_), .B(\a[5] ), .Y(new_n6335_));
  INVX1    g06079(.A(new_n6335_), .Y(new_n6336_));
  XOR2X1   g06080(.A(new_n6336_), .B(new_n6331_), .Y(new_n6337_));
  XOR2X1   g06081(.A(new_n6337_), .B(new_n6160_), .Y(new_n6338_));
  NAND2X1  g06082(.A(\b[55] ), .B(\b[54] ), .Y(new_n6339_));
  OAI21X1  g06083(.A0(new_n6149_), .A1(new_n6147_), .B0(new_n6339_), .Y(new_n6340_));
  XOR2X1   g06084(.A(\b[56] ), .B(\b[55] ), .Y(new_n6341_));
  XOR2X1   g06085(.A(new_n6341_), .B(new_n6340_), .Y(new_n6342_));
  AOI22X1  g06086(.A0(new_n267_), .A1(\b[56] ), .B0(new_n266_), .B1(\b[55] ), .Y(new_n6343_));
  OAI21X1  g06087(.A0(new_n350_), .A1(new_n6148_), .B0(new_n6343_), .Y(new_n6344_));
  AOI21X1  g06088(.A0(new_n6342_), .A1(new_n318_), .B0(new_n6344_), .Y(new_n6345_));
  XOR2X1   g06089(.A(new_n6345_), .B(\a[2] ), .Y(new_n6346_));
  XOR2X1   g06090(.A(new_n6346_), .B(new_n6338_), .Y(new_n6347_));
  OR2X1    g06091(.A(new_n6155_), .B(new_n6145_), .Y(new_n6348_));
  OAI21X1  g06092(.A0(new_n5968_), .A1(new_n5967_), .B0(new_n6156_), .Y(new_n6349_));
  AND2X1   g06093(.A(new_n6349_), .B(new_n6348_), .Y(new_n6350_));
  XOR2X1   g06094(.A(new_n6350_), .B(new_n6347_), .Y(\f[56] ));
  AND2X1   g06095(.A(new_n6336_), .B(new_n6331_), .Y(new_n6352_));
  AOI21X1  g06096(.A0(new_n6337_), .A1(new_n6160_), .B0(new_n6352_), .Y(new_n6353_));
  AOI22X1  g06097(.A0(new_n369_), .A1(\b[54] ), .B0(new_n368_), .B1(\b[53] ), .Y(new_n6354_));
  OAI21X1  g06098(.A0(new_n367_), .A1(new_n5808_), .B0(new_n6354_), .Y(new_n6355_));
  AOI21X1  g06099(.A0(new_n5807_), .A1(new_n308_), .B0(new_n6355_), .Y(new_n6356_));
  XOR2X1   g06100(.A(new_n6356_), .B(\a[5] ), .Y(new_n6357_));
  AND2X1   g06101(.A(new_n6329_), .B(new_n6172_), .Y(new_n6358_));
  AOI21X1  g06102(.A0(new_n6330_), .A1(new_n6167_), .B0(new_n6358_), .Y(new_n6359_));
  AOI22X1  g06103(.A0(new_n469_), .A1(\b[51] ), .B0(new_n468_), .B1(\b[50] ), .Y(new_n6360_));
  OAI21X1  g06104(.A0(new_n467_), .A1(new_n5237_), .B0(new_n6360_), .Y(new_n6361_));
  AOI21X1  g06105(.A0(new_n5236_), .A1(new_n404_), .B0(new_n6361_), .Y(new_n6362_));
  XOR2X1   g06106(.A(new_n6362_), .B(\a[8] ), .Y(new_n6363_));
  NOR2X1   g06107(.A(new_n6322_), .B(new_n6321_), .Y(new_n6364_));
  OR2X1    g06108(.A(new_n6327_), .B(new_n6364_), .Y(new_n6365_));
  OAI21X1  g06109(.A0(new_n6328_), .A1(new_n6174_), .B0(new_n6365_), .Y(new_n6366_));
  AOI22X1  g06110(.A0(new_n603_), .A1(\b[48] ), .B0(new_n602_), .B1(\b[47] ), .Y(new_n6367_));
  OAI21X1  g06111(.A0(new_n601_), .A1(new_n4693_), .B0(new_n6367_), .Y(new_n6368_));
  AOI21X1  g06112(.A0(new_n4692_), .A1(new_n518_), .B0(new_n6368_), .Y(new_n6369_));
  XOR2X1   g06113(.A(new_n6369_), .B(\a[11] ), .Y(new_n6370_));
  INVX1    g06114(.A(new_n6370_), .Y(new_n6371_));
  NAND2X1  g06115(.A(new_n6317_), .B(new_n6313_), .Y(new_n6372_));
  AOI21X1  g06116(.A0(new_n6372_), .A1(new_n6129_), .B0(new_n6318_), .Y(new_n6373_));
  AOI22X1  g06117(.A0(new_n818_), .A1(\b[45] ), .B0(new_n817_), .B1(\b[44] ), .Y(new_n6374_));
  OAI21X1  g06118(.A0(new_n816_), .A1(new_n4339_), .B0(new_n6374_), .Y(new_n6375_));
  AOI21X1  g06119(.A0(new_n4338_), .A1(new_n668_), .B0(new_n6375_), .Y(new_n6376_));
  XOR2X1   g06120(.A(new_n6376_), .B(\a[14] ), .Y(new_n6377_));
  OR2X1    g06121(.A(new_n6306_), .B(new_n6302_), .Y(new_n6378_));
  INVX1    g06122(.A(new_n6287_), .Y(new_n6379_));
  XOR2X1   g06123(.A(new_n6379_), .B(new_n6283_), .Y(new_n6380_));
  XOR2X1   g06124(.A(new_n6290_), .B(new_n6380_), .Y(new_n6381_));
  XOR2X1   g06125(.A(new_n6295_), .B(new_n6381_), .Y(new_n6382_));
  XOR2X1   g06126(.A(new_n6301_), .B(new_n6382_), .Y(new_n6383_));
  XOR2X1   g06127(.A(new_n6306_), .B(new_n6383_), .Y(new_n6384_));
  OAI21X1  g06128(.A0(new_n6312_), .A1(new_n6384_), .B0(new_n6378_), .Y(new_n6385_));
  NAND2X1  g06129(.A(new_n6379_), .B(new_n6283_), .Y(new_n6386_));
  OAI21X1  g06130(.A0(new_n6290_), .A1(new_n6288_), .B0(new_n6386_), .Y(new_n6387_));
  AND2X1   g06131(.A(new_n6281_), .B(new_n6182_), .Y(new_n6388_));
  AOI21X1  g06132(.A0(new_n6282_), .A1(new_n6177_), .B0(new_n6388_), .Y(new_n6389_));
  NOR2X1   g06133(.A(new_n6279_), .B(new_n6275_), .Y(new_n6390_));
  AOI21X1  g06134(.A0(new_n6280_), .A1(new_n6184_), .B0(new_n6390_), .Y(new_n6391_));
  AOI22X1  g06135(.A0(new_n2163_), .A1(\b[30] ), .B0(new_n2162_), .B1(\b[29] ), .Y(new_n6392_));
  OAI21X1  g06136(.A0(new_n2161_), .A1(new_n2231_), .B0(new_n6392_), .Y(new_n6393_));
  AOI21X1  g06137(.A0(new_n2230_), .A1(new_n1907_), .B0(new_n6393_), .Y(new_n6394_));
  XOR2X1   g06138(.A(new_n6394_), .B(\a[29] ), .Y(new_n6395_));
  INVX1    g06139(.A(new_n6395_), .Y(new_n6396_));
  OAI21X1  g06140(.A0(new_n6272_), .A1(new_n6269_), .B0(new_n6270_), .Y(new_n6397_));
  OR2X1    g06141(.A(new_n6251_), .B(new_n6247_), .Y(new_n6398_));
  OAI21X1  g06142(.A0(new_n6253_), .A1(new_n6056_), .B0(new_n6398_), .Y(new_n6399_));
  AOI22X1  g06143(.A0(new_n3204_), .A1(\b[21] ), .B0(new_n3203_), .B1(\b[20] ), .Y(new_n6400_));
  OAI21X1  g06144(.A0(new_n3321_), .A1(new_n1300_), .B0(new_n6400_), .Y(new_n6401_));
  AOI21X1  g06145(.A0(new_n3080_), .A1(new_n1299_), .B0(new_n6401_), .Y(new_n6402_));
  XOR2X1   g06146(.A(new_n6402_), .B(new_n3078_), .Y(new_n6403_));
  INVX1    g06147(.A(new_n6195_), .Y(new_n6404_));
  AND2X1   g06148(.A(new_n6245_), .B(new_n6404_), .Y(new_n6405_));
  INVX1    g06149(.A(new_n6246_), .Y(new_n6406_));
  AOI21X1  g06150(.A0(new_n6406_), .A1(new_n6191_), .B0(new_n6405_), .Y(new_n6407_));
  AOI22X1  g06151(.A0(new_n3652_), .A1(\b[18] ), .B0(new_n3651_), .B1(\b[17] ), .Y(new_n6408_));
  OAI21X1  g06152(.A0(new_n3778_), .A1(new_n974_), .B0(new_n6408_), .Y(new_n6409_));
  AOI21X1  g06153(.A0(new_n3480_), .A1(new_n1042_), .B0(new_n6409_), .Y(new_n6410_));
  XOR2X1   g06154(.A(new_n6410_), .B(\a[41] ), .Y(new_n6411_));
  INVX1    g06155(.A(new_n6239_), .Y(new_n6412_));
  OR2X1    g06156(.A(new_n6244_), .B(new_n6197_), .Y(new_n6413_));
  OAI21X1  g06157(.A0(new_n6243_), .A1(new_n6412_), .B0(new_n6413_), .Y(new_n6414_));
  AOI22X1  g06158(.A0(new_n4095_), .A1(\b[15] ), .B0(new_n4094_), .B1(\b[14] ), .Y(new_n6415_));
  OAI21X1  g06159(.A0(new_n4233_), .A1(new_n795_), .B0(new_n6415_), .Y(new_n6416_));
  AOI21X1  g06160(.A0(new_n3901_), .A1(new_n794_), .B0(new_n6416_), .Y(new_n6417_));
  XOR2X1   g06161(.A(new_n6417_), .B(\a[44] ), .Y(new_n6418_));
  INVX1    g06162(.A(new_n6418_), .Y(new_n6419_));
  AND2X1   g06163(.A(new_n6236_), .B(new_n6204_), .Y(new_n6420_));
  INVX1    g06164(.A(new_n6420_), .Y(new_n6421_));
  OR2X1    g06165(.A(new_n6238_), .B(new_n6199_), .Y(new_n6422_));
  AND2X1   g06166(.A(new_n6422_), .B(new_n6421_), .Y(new_n6423_));
  AOI22X1  g06167(.A0(new_n4572_), .A1(\b[12] ), .B0(new_n4571_), .B1(\b[11] ), .Y(new_n6424_));
  OAI21X1  g06168(.A0(new_n4740_), .A1(new_n587_), .B0(new_n6424_), .Y(new_n6425_));
  AOI21X1  g06169(.A0(new_n4375_), .A1(new_n635_), .B0(new_n6425_), .Y(new_n6426_));
  XOR2X1   g06170(.A(new_n6426_), .B(\a[47] ), .Y(new_n6427_));
  INVX1    g06171(.A(new_n6427_), .Y(new_n6428_));
  OAI21X1  g06172(.A0(new_n6206_), .A1(new_n6205_), .B0(new_n6235_), .Y(new_n6429_));
  OAI21X1  g06173(.A0(new_n6234_), .A1(new_n6230_), .B0(new_n6429_), .Y(new_n6430_));
  NOR4X1   g06174(.A(new_n6217_), .B(new_n6029_), .C(new_n5888_), .D(new_n6019_), .Y(new_n6431_));
  XOR2X1   g06175(.A(\a[57] ), .B(new_n6019_), .Y(new_n6432_));
  NOR2X1   g06176(.A(new_n6432_), .B(new_n274_), .Y(new_n6433_));
  INVX1    g06177(.A(new_n6433_), .Y(new_n6434_));
  XOR2X1   g06178(.A(new_n6434_), .B(new_n6431_), .Y(new_n6435_));
  INVX1    g06179(.A(new_n6214_), .Y(new_n6436_));
  INVX1    g06180(.A(new_n6025_), .Y(new_n6437_));
  INVX1    g06181(.A(new_n6026_), .Y(new_n6438_));
  AOI22X1  g06182(.A0(new_n6438_), .A1(\b[3] ), .B0(new_n6437_), .B1(\b[2] ), .Y(new_n6439_));
  OAI21X1  g06183(.A0(new_n6436_), .A1(new_n275_), .B0(new_n6439_), .Y(new_n6440_));
  AOI21X1  g06184(.A0(new_n6023_), .A1(new_n366_), .B0(new_n6440_), .Y(new_n6441_));
  XOR2X1   g06185(.A(new_n6441_), .B(\a[56] ), .Y(new_n6442_));
  XOR2X1   g06186(.A(new_n6442_), .B(new_n6435_), .Y(new_n6443_));
  AOI22X1  g06187(.A0(new_n5430_), .A1(\b[6] ), .B0(new_n5427_), .B1(\b[5] ), .Y(new_n6444_));
  OAI21X1  g06188(.A0(new_n5891_), .A1(new_n325_), .B0(new_n6444_), .Y(new_n6445_));
  AOI21X1  g06189(.A0(new_n5425_), .A1(new_n378_), .B0(new_n6445_), .Y(new_n6446_));
  XOR2X1   g06190(.A(new_n6446_), .B(\a[53] ), .Y(new_n6447_));
  XOR2X1   g06191(.A(new_n6447_), .B(new_n6443_), .Y(new_n6448_));
  INVX1    g06192(.A(new_n6448_), .Y(new_n6449_));
  XOR2X1   g06193(.A(new_n6449_), .B(new_n6229_), .Y(new_n6450_));
  AOI22X1  g06194(.A0(new_n4880_), .A1(\b[9] ), .B0(new_n4877_), .B1(\b[8] ), .Y(new_n6451_));
  OAI21X1  g06195(.A0(new_n5291_), .A1(new_n492_), .B0(new_n6451_), .Y(new_n6452_));
  AOI21X1  g06196(.A0(new_n4875_), .A1(new_n491_), .B0(new_n6452_), .Y(new_n6453_));
  XOR2X1   g06197(.A(new_n6453_), .B(\a[50] ), .Y(new_n6454_));
  XOR2X1   g06198(.A(new_n6454_), .B(new_n6450_), .Y(new_n6455_));
  XOR2X1   g06199(.A(new_n6455_), .B(new_n6430_), .Y(new_n6456_));
  XOR2X1   g06200(.A(new_n6456_), .B(new_n6428_), .Y(new_n6457_));
  INVX1    g06201(.A(new_n6457_), .Y(new_n6458_));
  XOR2X1   g06202(.A(new_n6458_), .B(new_n6423_), .Y(new_n6459_));
  XOR2X1   g06203(.A(new_n6459_), .B(new_n6419_), .Y(new_n6460_));
  XOR2X1   g06204(.A(new_n6460_), .B(new_n6414_), .Y(new_n6461_));
  XOR2X1   g06205(.A(new_n6461_), .B(new_n6411_), .Y(new_n6462_));
  XOR2X1   g06206(.A(new_n6462_), .B(new_n6407_), .Y(new_n6463_));
  XOR2X1   g06207(.A(new_n6463_), .B(new_n6403_), .Y(new_n6464_));
  XOR2X1   g06208(.A(new_n6464_), .B(new_n6399_), .Y(new_n6465_));
  AOI22X1  g06209(.A0(new_n2813_), .A1(\b[24] ), .B0(new_n2812_), .B1(\b[23] ), .Y(new_n6466_));
  OAI21X1  g06210(.A0(new_n2946_), .A1(new_n1479_), .B0(new_n6466_), .Y(new_n6467_));
  AOI21X1  g06211(.A0(new_n2652_), .A1(new_n1572_), .B0(new_n6467_), .Y(new_n6468_));
  XOR2X1   g06212(.A(new_n6468_), .B(\a[35] ), .Y(new_n6469_));
  XOR2X1   g06213(.A(new_n6469_), .B(new_n6465_), .Y(new_n6470_));
  INVX1    g06214(.A(new_n6470_), .Y(new_n6471_));
  NOR2X1   g06215(.A(new_n6259_), .B(new_n6255_), .Y(new_n6472_));
  AOI21X1  g06216(.A0(new_n6260_), .A1(new_n6188_), .B0(new_n6472_), .Y(new_n6473_));
  XOR2X1   g06217(.A(new_n6473_), .B(new_n6471_), .Y(new_n6474_));
  AOI22X1  g06218(.A0(new_n2545_), .A1(\b[27] ), .B0(new_n2544_), .B1(\b[26] ), .Y(new_n6475_));
  OAI21X1  g06219(.A0(new_n2543_), .A1(new_n1880_), .B0(new_n6475_), .Y(new_n6476_));
  AOI21X1  g06220(.A0(new_n2260_), .A1(new_n1879_), .B0(new_n6476_), .Y(new_n6477_));
  XOR2X1   g06221(.A(new_n6477_), .B(\a[32] ), .Y(new_n6478_));
  XOR2X1   g06222(.A(new_n6478_), .B(new_n6474_), .Y(new_n6479_));
  XOR2X1   g06223(.A(new_n6479_), .B(new_n6397_), .Y(new_n6480_));
  XOR2X1   g06224(.A(new_n6480_), .B(new_n6396_), .Y(new_n6481_));
  XOR2X1   g06225(.A(new_n6481_), .B(new_n6391_), .Y(new_n6482_));
  AOI22X1  g06226(.A0(new_n1814_), .A1(\b[33] ), .B0(new_n1813_), .B1(\b[32] ), .Y(new_n6483_));
  OAI21X1  g06227(.A0(new_n1812_), .A1(new_n2615_), .B0(new_n6483_), .Y(new_n6484_));
  AOI21X1  g06228(.A0(new_n2614_), .A1(new_n1617_), .B0(new_n6484_), .Y(new_n6485_));
  XOR2X1   g06229(.A(new_n6485_), .B(\a[26] ), .Y(new_n6486_));
  XOR2X1   g06230(.A(new_n6486_), .B(new_n6482_), .Y(new_n6487_));
  XOR2X1   g06231(.A(new_n6487_), .B(new_n6389_), .Y(new_n6488_));
  AOI22X1  g06232(.A0(new_n1526_), .A1(\b[36] ), .B0(new_n1525_), .B1(\b[35] ), .Y(new_n6489_));
  OAI21X1  g06233(.A0(new_n1524_), .A1(new_n2890_), .B0(new_n6489_), .Y(new_n6490_));
  AOI21X1  g06234(.A0(new_n3015_), .A1(new_n1347_), .B0(new_n6490_), .Y(new_n6491_));
  XOR2X1   g06235(.A(new_n6491_), .B(\a[23] ), .Y(new_n6492_));
  XOR2X1   g06236(.A(new_n6492_), .B(new_n6488_), .Y(new_n6493_));
  XOR2X1   g06237(.A(new_n6493_), .B(new_n6387_), .Y(new_n6494_));
  AOI22X1  g06238(.A0(new_n1263_), .A1(\b[39] ), .B0(new_n1262_), .B1(\b[38] ), .Y(new_n6495_));
  OAI21X1  g06239(.A0(new_n1261_), .A1(new_n3413_), .B0(new_n6495_), .Y(new_n6496_));
  AOI21X1  g06240(.A0(new_n3412_), .A1(new_n1075_), .B0(new_n6496_), .Y(new_n6497_));
  XOR2X1   g06241(.A(new_n6497_), .B(\a[20] ), .Y(new_n6498_));
  INVX1    g06242(.A(new_n6498_), .Y(new_n6499_));
  XOR2X1   g06243(.A(new_n6499_), .B(new_n6494_), .Y(new_n6500_));
  NOR2X1   g06244(.A(new_n6295_), .B(new_n6381_), .Y(new_n6501_));
  AOI21X1  g06245(.A0(new_n6301_), .A1(new_n6382_), .B0(new_n6501_), .Y(new_n6502_));
  XOR2X1   g06246(.A(new_n6502_), .B(new_n6500_), .Y(new_n6503_));
  AOI22X1  g06247(.A0(new_n1017_), .A1(\b[42] ), .B0(new_n1016_), .B1(\b[41] ), .Y(new_n6504_));
  OAI21X1  g06248(.A0(new_n1015_), .A1(new_n3720_), .B0(new_n6504_), .Y(new_n6505_));
  AOI21X1  g06249(.A0(new_n3860_), .A1(new_n882_), .B0(new_n6505_), .Y(new_n6506_));
  XOR2X1   g06250(.A(new_n6506_), .B(\a[17] ), .Y(new_n6507_));
  XOR2X1   g06251(.A(new_n6507_), .B(new_n6503_), .Y(new_n6508_));
  XOR2X1   g06252(.A(new_n6508_), .B(new_n6385_), .Y(new_n6509_));
  XOR2X1   g06253(.A(new_n6509_), .B(new_n6377_), .Y(new_n6510_));
  XOR2X1   g06254(.A(new_n6510_), .B(new_n6373_), .Y(new_n6511_));
  XOR2X1   g06255(.A(new_n6511_), .B(new_n6371_), .Y(new_n6512_));
  XOR2X1   g06256(.A(new_n6512_), .B(new_n6366_), .Y(new_n6513_));
  XOR2X1   g06257(.A(new_n6513_), .B(new_n6363_), .Y(new_n6514_));
  XOR2X1   g06258(.A(new_n6514_), .B(new_n6359_), .Y(new_n6515_));
  XOR2X1   g06259(.A(new_n6515_), .B(new_n6357_), .Y(new_n6516_));
  XOR2X1   g06260(.A(new_n6516_), .B(new_n6353_), .Y(new_n6517_));
  AND2X1   g06261(.A(\b[56] ), .B(\b[55] ), .Y(new_n6518_));
  AOI21X1  g06262(.A0(new_n6341_), .A1(new_n6340_), .B0(new_n6518_), .Y(new_n6519_));
  INVX1    g06263(.A(\b[56] ), .Y(new_n6520_));
  XOR2X1   g06264(.A(\b[57] ), .B(new_n6520_), .Y(new_n6521_));
  XOR2X1   g06265(.A(new_n6521_), .B(new_n6519_), .Y(new_n6522_));
  INVX1    g06266(.A(\b[55] ), .Y(new_n6523_));
  AOI22X1  g06267(.A0(new_n267_), .A1(\b[57] ), .B0(new_n266_), .B1(\b[56] ), .Y(new_n6524_));
  OAI21X1  g06268(.A0(new_n350_), .A1(new_n6523_), .B0(new_n6524_), .Y(new_n6525_));
  AOI21X1  g06269(.A0(new_n6522_), .A1(new_n318_), .B0(new_n6525_), .Y(new_n6526_));
  XOR2X1   g06270(.A(new_n6526_), .B(new_n257_), .Y(new_n6527_));
  XOR2X1   g06271(.A(new_n6527_), .B(new_n6517_), .Y(new_n6528_));
  XOR2X1   g06272(.A(new_n6345_), .B(new_n257_), .Y(new_n6529_));
  AND2X1   g06273(.A(new_n6529_), .B(new_n6338_), .Y(new_n6530_));
  AOI21X1  g06274(.A0(new_n6349_), .A1(new_n6348_), .B0(new_n6347_), .Y(new_n6531_));
  OR2X1    g06275(.A(new_n6531_), .B(new_n6530_), .Y(new_n6532_));
  XOR2X1   g06276(.A(new_n6532_), .B(new_n6528_), .Y(\f[57] ));
  INVX1    g06277(.A(new_n6357_), .Y(new_n6534_));
  NAND2X1  g06278(.A(new_n6515_), .B(new_n6534_), .Y(new_n6535_));
  OAI21X1  g06279(.A0(new_n6516_), .A1(new_n6353_), .B0(new_n6535_), .Y(new_n6536_));
  AOI22X1  g06280(.A0(new_n369_), .A1(\b[55] ), .B0(new_n368_), .B1(\b[54] ), .Y(new_n6537_));
  OAI21X1  g06281(.A0(new_n367_), .A1(new_n6151_), .B0(new_n6537_), .Y(new_n6538_));
  AOI21X1  g06282(.A0(new_n6150_), .A1(new_n308_), .B0(new_n6538_), .Y(new_n6539_));
  XOR2X1   g06283(.A(new_n6539_), .B(new_n305_), .Y(new_n6540_));
  INVX1    g06284(.A(new_n6363_), .Y(new_n6541_));
  NAND2X1  g06285(.A(new_n6513_), .B(new_n6541_), .Y(new_n6542_));
  OAI21X1  g06286(.A0(new_n6514_), .A1(new_n6359_), .B0(new_n6542_), .Y(new_n6543_));
  AOI22X1  g06287(.A0(new_n469_), .A1(\b[52] ), .B0(new_n468_), .B1(\b[51] ), .Y(new_n6544_));
  OAI21X1  g06288(.A0(new_n467_), .A1(new_n5234_), .B0(new_n6544_), .Y(new_n6545_));
  AOI21X1  g06289(.A0(new_n5590_), .A1(new_n404_), .B0(new_n6545_), .Y(new_n6546_));
  XOR2X1   g06290(.A(new_n6546_), .B(new_n400_), .Y(new_n6547_));
  OR2X1    g06291(.A(new_n5946_), .B(new_n5775_), .Y(new_n6548_));
  AND2X1   g06292(.A(new_n6548_), .B(new_n5981_), .Y(new_n6549_));
  NOR2X1   g06293(.A(new_n6134_), .B(new_n6130_), .Y(new_n6550_));
  NAND2X1  g06294(.A(new_n6134_), .B(new_n6130_), .Y(new_n6551_));
  OAI21X1  g06295(.A0(new_n6550_), .A1(new_n6549_), .B0(new_n6551_), .Y(new_n6552_));
  NOR2X1   g06296(.A(new_n6327_), .B(new_n6364_), .Y(new_n6553_));
  XOR2X1   g06297(.A(new_n6327_), .B(new_n6364_), .Y(new_n6554_));
  AOI21X1  g06298(.A0(new_n6554_), .A1(new_n6552_), .B0(new_n6553_), .Y(new_n6555_));
  NAND2X1  g06299(.A(new_n6511_), .B(new_n6371_), .Y(new_n6556_));
  XOR2X1   g06300(.A(new_n6511_), .B(new_n6370_), .Y(new_n6557_));
  OAI21X1  g06301(.A0(new_n6557_), .A1(new_n6555_), .B0(new_n6556_), .Y(new_n6558_));
  AOI22X1  g06302(.A0(new_n603_), .A1(\b[49] ), .B0(new_n602_), .B1(\b[48] ), .Y(new_n6559_));
  OAI21X1  g06303(.A0(new_n601_), .A1(new_n5039_), .B0(new_n6559_), .Y(new_n6560_));
  AOI21X1  g06304(.A0(new_n5038_), .A1(new_n518_), .B0(new_n6560_), .Y(new_n6561_));
  XOR2X1   g06305(.A(new_n6561_), .B(new_n515_), .Y(new_n6562_));
  INVX1    g06306(.A(new_n6377_), .Y(new_n6563_));
  NAND2X1  g06307(.A(new_n6509_), .B(new_n6563_), .Y(new_n6564_));
  OAI21X1  g06308(.A0(new_n6510_), .A1(new_n6373_), .B0(new_n6564_), .Y(new_n6565_));
  NOR2X1   g06309(.A(new_n6507_), .B(new_n6503_), .Y(new_n6566_));
  AOI21X1  g06310(.A0(new_n6508_), .A1(new_n6385_), .B0(new_n6566_), .Y(new_n6567_));
  NAND2X1  g06311(.A(new_n6480_), .B(new_n6396_), .Y(new_n6568_));
  INVX1    g06312(.A(new_n6481_), .Y(new_n6569_));
  OAI21X1  g06313(.A0(new_n6569_), .A1(new_n6391_), .B0(new_n6568_), .Y(new_n6570_));
  NOR2X1   g06314(.A(new_n6478_), .B(new_n6474_), .Y(new_n6571_));
  AOI21X1  g06315(.A0(new_n6479_), .A1(new_n6397_), .B0(new_n6571_), .Y(new_n6572_));
  INVX1    g06316(.A(new_n6411_), .Y(new_n6573_));
  AND2X1   g06317(.A(new_n6461_), .B(new_n6573_), .Y(new_n6574_));
  NOR2X1   g06318(.A(new_n6462_), .B(new_n6407_), .Y(new_n6575_));
  OR2X1    g06319(.A(new_n6575_), .B(new_n6574_), .Y(new_n6576_));
  AOI21X1  g06320(.A0(new_n6422_), .A1(new_n6421_), .B0(new_n6458_), .Y(new_n6577_));
  AOI21X1  g06321(.A0(new_n6456_), .A1(new_n6428_), .B0(new_n6577_), .Y(new_n6578_));
  XOR2X1   g06322(.A(new_n6446_), .B(new_n5423_), .Y(new_n6579_));
  AND2X1   g06323(.A(new_n6579_), .B(new_n6443_), .Y(new_n6580_));
  NOR2X1   g06324(.A(new_n6448_), .B(new_n6229_), .Y(new_n6581_));
  NOR2X1   g06325(.A(new_n6581_), .B(new_n6580_), .Y(new_n6582_));
  INVX1    g06326(.A(new_n6582_), .Y(new_n6583_));
  AOI22X1  g06327(.A0(new_n5430_), .A1(\b[7] ), .B0(new_n5427_), .B1(\b[6] ), .Y(new_n6584_));
  OAI21X1  g06328(.A0(new_n5891_), .A1(new_n395_), .B0(new_n6584_), .Y(new_n6585_));
  AOI21X1  g06329(.A0(new_n5425_), .A1(new_n394_), .B0(new_n6585_), .Y(new_n6586_));
  XOR2X1   g06330(.A(new_n6586_), .B(new_n5423_), .Y(new_n6587_));
  NAND2X1  g06331(.A(new_n6433_), .B(new_n6431_), .Y(new_n6588_));
  OAI21X1  g06332(.A0(new_n6442_), .A1(new_n6435_), .B0(new_n6588_), .Y(new_n6589_));
  AND2X1   g06333(.A(new_n6023_), .B(new_n323_), .Y(new_n6590_));
  NOR3X1   g06334(.A(new_n6213_), .B(new_n6022_), .C(new_n277_), .Y(new_n6591_));
  OAI22X1  g06335(.A0(new_n6026_), .A1(new_n325_), .B0(new_n6025_), .B1(new_n297_), .Y(new_n6592_));
  NOR3X1   g06336(.A(new_n6592_), .B(new_n6591_), .C(new_n6590_), .Y(new_n6593_));
  XOR2X1   g06337(.A(new_n6593_), .B(new_n6019_), .Y(new_n6594_));
  OAI21X1  g06338(.A0(new_n6432_), .A1(new_n274_), .B0(\a[59] ), .Y(new_n6595_));
  INVX1    g06339(.A(\a[59] ), .Y(new_n6596_));
  XOR2X1   g06340(.A(new_n6596_), .B(\a[58] ), .Y(new_n6597_));
  NOR2X1   g06341(.A(new_n6597_), .B(new_n6432_), .Y(new_n6598_));
  XOR2X1   g06342(.A(\a[58] ), .B(\a[57] ), .Y(new_n6599_));
  AND2X1   g06343(.A(new_n6599_), .B(new_n6432_), .Y(new_n6600_));
  INVX1    g06344(.A(new_n6600_), .Y(new_n6601_));
  INVX1    g06345(.A(new_n6432_), .Y(new_n6602_));
  AND2X1   g06346(.A(new_n6597_), .B(new_n6602_), .Y(new_n6603_));
  INVX1    g06347(.A(new_n6603_), .Y(new_n6604_));
  OAI22X1  g06348(.A0(new_n6604_), .A1(new_n275_), .B0(new_n6601_), .B1(new_n274_), .Y(new_n6605_));
  AOI21X1  g06349(.A0(new_n6598_), .A1(new_n263_), .B0(new_n6605_), .Y(new_n6606_));
  XOR2X1   g06350(.A(new_n6606_), .B(\a[59] ), .Y(new_n6607_));
  XOR2X1   g06351(.A(new_n6607_), .B(new_n6595_), .Y(new_n6608_));
  XOR2X1   g06352(.A(new_n6608_), .B(new_n6594_), .Y(new_n6609_));
  XOR2X1   g06353(.A(new_n6609_), .B(new_n6589_), .Y(new_n6610_));
  XOR2X1   g06354(.A(new_n6610_), .B(new_n6587_), .Y(new_n6611_));
  XOR2X1   g06355(.A(new_n6611_), .B(new_n6583_), .Y(new_n6612_));
  AOI22X1  g06356(.A0(new_n4880_), .A1(\b[10] ), .B0(new_n4877_), .B1(\b[9] ), .Y(new_n6613_));
  OAI21X1  g06357(.A0(new_n5291_), .A1(new_n489_), .B0(new_n6613_), .Y(new_n6614_));
  AOI21X1  g06358(.A0(new_n4875_), .A1(new_n543_), .B0(new_n6614_), .Y(new_n6615_));
  XOR2X1   g06359(.A(new_n6615_), .B(\a[50] ), .Y(new_n6616_));
  XOR2X1   g06360(.A(new_n6616_), .B(new_n6612_), .Y(new_n6617_));
  NOR2X1   g06361(.A(new_n6454_), .B(new_n6450_), .Y(new_n6618_));
  AOI21X1  g06362(.A0(new_n6455_), .A1(new_n6430_), .B0(new_n6618_), .Y(new_n6619_));
  XOR2X1   g06363(.A(new_n6619_), .B(new_n6617_), .Y(new_n6620_));
  INVX1    g06364(.A(new_n6620_), .Y(new_n6621_));
  AOI22X1  g06365(.A0(new_n4572_), .A1(\b[13] ), .B0(new_n4571_), .B1(\b[12] ), .Y(new_n6622_));
  OAI21X1  g06366(.A0(new_n4740_), .A1(new_n716_), .B0(new_n6622_), .Y(new_n6623_));
  AOI21X1  g06367(.A0(new_n4375_), .A1(new_n715_), .B0(new_n6623_), .Y(new_n6624_));
  XOR2X1   g06368(.A(new_n6624_), .B(\a[47] ), .Y(new_n6625_));
  AND2X1   g06369(.A(new_n6625_), .B(new_n6621_), .Y(new_n6626_));
  XOR2X1   g06370(.A(new_n6625_), .B(new_n6621_), .Y(new_n6627_));
  NOR2X1   g06371(.A(new_n6625_), .B(new_n6621_), .Y(new_n6628_));
  INVX1    g06372(.A(new_n6628_), .Y(new_n6629_));
  OAI21X1  g06373(.A0(new_n6626_), .A1(new_n6578_), .B0(new_n6629_), .Y(new_n6630_));
  OAI22X1  g06374(.A0(new_n6630_), .A1(new_n6626_), .B0(new_n6627_), .B1(new_n6578_), .Y(new_n6631_));
  AOI22X1  g06375(.A0(new_n4095_), .A1(\b[16] ), .B0(new_n4094_), .B1(\b[15] ), .Y(new_n6632_));
  OAI21X1  g06376(.A0(new_n4233_), .A1(new_n792_), .B0(new_n6632_), .Y(new_n6633_));
  AOI21X1  g06377(.A0(new_n3901_), .A1(new_n842_), .B0(new_n6633_), .Y(new_n6634_));
  XOR2X1   g06378(.A(new_n6634_), .B(\a[44] ), .Y(new_n6635_));
  XOR2X1   g06379(.A(new_n6635_), .B(new_n6631_), .Y(new_n6636_));
  AND2X1   g06380(.A(new_n6459_), .B(new_n6419_), .Y(new_n6637_));
  AOI21X1  g06381(.A0(new_n6460_), .A1(new_n6414_), .B0(new_n6637_), .Y(new_n6638_));
  XOR2X1   g06382(.A(new_n6638_), .B(new_n6636_), .Y(new_n6639_));
  INVX1    g06383(.A(new_n6639_), .Y(new_n6640_));
  AOI22X1  g06384(.A0(new_n3652_), .A1(\b[19] ), .B0(new_n3651_), .B1(\b[18] ), .Y(new_n6641_));
  OAI21X1  g06385(.A0(new_n3778_), .A1(new_n1118_), .B0(new_n6641_), .Y(new_n6642_));
  AOI21X1  g06386(.A0(new_n3480_), .A1(new_n1117_), .B0(new_n6642_), .Y(new_n6643_));
  XOR2X1   g06387(.A(new_n6643_), .B(\a[41] ), .Y(new_n6644_));
  NAND2X1  g06388(.A(new_n6644_), .B(new_n6640_), .Y(new_n6645_));
  XOR2X1   g06389(.A(new_n6644_), .B(new_n6640_), .Y(new_n6646_));
  INVX1    g06390(.A(new_n6646_), .Y(new_n6647_));
  NOR2X1   g06391(.A(new_n6644_), .B(new_n6640_), .Y(new_n6648_));
  AOI21X1  g06392(.A0(new_n6645_), .A1(new_n6576_), .B0(new_n6648_), .Y(new_n6649_));
  AOI22X1  g06393(.A0(new_n6649_), .A1(new_n6645_), .B0(new_n6647_), .B1(new_n6576_), .Y(new_n6650_));
  AOI22X1  g06394(.A0(new_n3204_), .A1(\b[22] ), .B0(new_n3203_), .B1(\b[21] ), .Y(new_n6651_));
  OAI21X1  g06395(.A0(new_n3321_), .A1(new_n1297_), .B0(new_n6651_), .Y(new_n6652_));
  AOI21X1  g06396(.A0(new_n3080_), .A1(new_n1399_), .B0(new_n6652_), .Y(new_n6653_));
  XOR2X1   g06397(.A(new_n6653_), .B(\a[38] ), .Y(new_n6654_));
  XOR2X1   g06398(.A(new_n6654_), .B(new_n6650_), .Y(new_n6655_));
  AND2X1   g06399(.A(new_n6463_), .B(new_n6403_), .Y(new_n6656_));
  AOI21X1  g06400(.A0(new_n6464_), .A1(new_n6399_), .B0(new_n6656_), .Y(new_n6657_));
  XOR2X1   g06401(.A(new_n6657_), .B(new_n6655_), .Y(new_n6658_));
  AOI22X1  g06402(.A0(new_n2813_), .A1(\b[25] ), .B0(new_n2812_), .B1(\b[24] ), .Y(new_n6659_));
  OAI21X1  g06403(.A0(new_n2946_), .A1(new_n1591_), .B0(new_n6659_), .Y(new_n6660_));
  AOI21X1  g06404(.A0(new_n2652_), .A1(new_n1590_), .B0(new_n6660_), .Y(new_n6661_));
  XOR2X1   g06405(.A(new_n6661_), .B(\a[35] ), .Y(new_n6662_));
  XOR2X1   g06406(.A(new_n6662_), .B(new_n6658_), .Y(new_n6663_));
  INVX1    g06407(.A(new_n6465_), .Y(new_n6664_));
  OR2X1    g06408(.A(new_n6469_), .B(new_n6664_), .Y(new_n6665_));
  OAI21X1  g06409(.A0(new_n6473_), .A1(new_n6470_), .B0(new_n6665_), .Y(new_n6666_));
  XOR2X1   g06410(.A(new_n6666_), .B(new_n6663_), .Y(new_n6667_));
  AOI22X1  g06411(.A0(new_n2545_), .A1(\b[28] ), .B0(new_n2544_), .B1(\b[27] ), .Y(new_n6668_));
  OAI21X1  g06412(.A0(new_n2543_), .A1(new_n1877_), .B0(new_n6668_), .Y(new_n6669_));
  AOI21X1  g06413(.A0(new_n2260_), .A1(new_n2004_), .B0(new_n6669_), .Y(new_n6670_));
  XOR2X1   g06414(.A(new_n6670_), .B(\a[32] ), .Y(new_n6671_));
  XOR2X1   g06415(.A(new_n6671_), .B(new_n6667_), .Y(new_n6672_));
  XOR2X1   g06416(.A(new_n6672_), .B(new_n6572_), .Y(new_n6673_));
  AOI22X1  g06417(.A0(new_n2163_), .A1(\b[31] ), .B0(new_n2162_), .B1(\b[30] ), .Y(new_n6674_));
  OAI21X1  g06418(.A0(new_n2161_), .A1(new_n2359_), .B0(new_n6674_), .Y(new_n6675_));
  AOI21X1  g06419(.A0(new_n2358_), .A1(new_n1907_), .B0(new_n6675_), .Y(new_n6676_));
  XOR2X1   g06420(.A(new_n6676_), .B(\a[29] ), .Y(new_n6677_));
  XOR2X1   g06421(.A(new_n6677_), .B(new_n6673_), .Y(new_n6678_));
  XOR2X1   g06422(.A(new_n6678_), .B(new_n6570_), .Y(new_n6679_));
  AOI22X1  g06423(.A0(new_n1814_), .A1(\b[34] ), .B0(new_n1813_), .B1(\b[33] ), .Y(new_n6680_));
  OAI21X1  g06424(.A0(new_n1812_), .A1(new_n2612_), .B0(new_n6680_), .Y(new_n6681_));
  AOI21X1  g06425(.A0(new_n2759_), .A1(new_n1617_), .B0(new_n6681_), .Y(new_n6682_));
  XOR2X1   g06426(.A(new_n6682_), .B(\a[26] ), .Y(new_n6683_));
  XOR2X1   g06427(.A(new_n6683_), .B(new_n6679_), .Y(new_n6684_));
  OR2X1    g06428(.A(new_n6486_), .B(new_n6482_), .Y(new_n6685_));
  INVX1    g06429(.A(new_n6486_), .Y(new_n6686_));
  XOR2X1   g06430(.A(new_n6686_), .B(new_n6482_), .Y(new_n6687_));
  OAI21X1  g06431(.A0(new_n6687_), .A1(new_n6389_), .B0(new_n6685_), .Y(new_n6688_));
  XOR2X1   g06432(.A(new_n6688_), .B(new_n6684_), .Y(new_n6689_));
  AOI22X1  g06433(.A0(new_n1526_), .A1(\b[37] ), .B0(new_n1525_), .B1(\b[36] ), .Y(new_n6690_));
  OAI21X1  g06434(.A0(new_n1524_), .A1(new_n3156_), .B0(new_n6690_), .Y(new_n6691_));
  AOI21X1  g06435(.A0(new_n3155_), .A1(new_n1347_), .B0(new_n6691_), .Y(new_n6692_));
  XOR2X1   g06436(.A(new_n6692_), .B(\a[23] ), .Y(new_n6693_));
  XOR2X1   g06437(.A(new_n6693_), .B(new_n6689_), .Y(new_n6694_));
  NOR2X1   g06438(.A(new_n6492_), .B(new_n6488_), .Y(new_n6695_));
  AOI21X1  g06439(.A0(new_n6493_), .A1(new_n6387_), .B0(new_n6695_), .Y(new_n6696_));
  XOR2X1   g06440(.A(new_n6696_), .B(new_n6694_), .Y(new_n6697_));
  AOI22X1  g06441(.A0(new_n1263_), .A1(\b[40] ), .B0(new_n1262_), .B1(\b[39] ), .Y(new_n6698_));
  OAI21X1  g06442(.A0(new_n1261_), .A1(new_n3575_), .B0(new_n6698_), .Y(new_n6699_));
  AOI21X1  g06443(.A0(new_n3574_), .A1(new_n1075_), .B0(new_n6699_), .Y(new_n6700_));
  XOR2X1   g06444(.A(new_n6700_), .B(\a[20] ), .Y(new_n6701_));
  XOR2X1   g06445(.A(new_n6701_), .B(new_n6697_), .Y(new_n6702_));
  NAND2X1  g06446(.A(new_n6499_), .B(new_n6494_), .Y(new_n6703_));
  XOR2X1   g06447(.A(new_n6498_), .B(new_n6494_), .Y(new_n6704_));
  OAI21X1  g06448(.A0(new_n6502_), .A1(new_n6704_), .B0(new_n6703_), .Y(new_n6705_));
  XOR2X1   g06449(.A(new_n6705_), .B(new_n6702_), .Y(new_n6706_));
  AOI22X1  g06450(.A0(new_n1017_), .A1(\b[43] ), .B0(new_n1016_), .B1(\b[42] ), .Y(new_n6707_));
  OAI21X1  g06451(.A0(new_n1015_), .A1(new_n4015_), .B0(new_n6707_), .Y(new_n6708_));
  AOI21X1  g06452(.A0(new_n4014_), .A1(new_n882_), .B0(new_n6708_), .Y(new_n6709_));
  XOR2X1   g06453(.A(new_n6709_), .B(\a[17] ), .Y(new_n6710_));
  AND2X1   g06454(.A(new_n6710_), .B(new_n6706_), .Y(new_n6711_));
  XOR2X1   g06455(.A(new_n6710_), .B(new_n6706_), .Y(new_n6712_));
  OR2X1    g06456(.A(new_n6710_), .B(new_n6706_), .Y(new_n6713_));
  OAI21X1  g06457(.A0(new_n6711_), .A1(new_n6567_), .B0(new_n6713_), .Y(new_n6714_));
  OAI22X1  g06458(.A0(new_n6714_), .A1(new_n6711_), .B0(new_n6712_), .B1(new_n6567_), .Y(new_n6715_));
  AOI22X1  g06459(.A0(new_n818_), .A1(\b[46] ), .B0(new_n817_), .B1(\b[45] ), .Y(new_n6716_));
  OAI21X1  g06460(.A0(new_n816_), .A1(new_n4336_), .B0(new_n6716_), .Y(new_n6717_));
  AOI21X1  g06461(.A0(new_n4509_), .A1(new_n668_), .B0(new_n6717_), .Y(new_n6718_));
  XOR2X1   g06462(.A(new_n6718_), .B(\a[14] ), .Y(new_n6719_));
  INVX1    g06463(.A(new_n6719_), .Y(new_n6720_));
  XOR2X1   g06464(.A(new_n6720_), .B(new_n6715_), .Y(new_n6721_));
  XOR2X1   g06465(.A(new_n6721_), .B(new_n6565_), .Y(new_n6722_));
  XOR2X1   g06466(.A(new_n6722_), .B(new_n6562_), .Y(new_n6723_));
  XOR2X1   g06467(.A(new_n6723_), .B(new_n6558_), .Y(new_n6724_));
  XOR2X1   g06468(.A(new_n6724_), .B(new_n6547_), .Y(new_n6725_));
  XOR2X1   g06469(.A(new_n6725_), .B(new_n6543_), .Y(new_n6726_));
  XOR2X1   g06470(.A(new_n6726_), .B(new_n6540_), .Y(new_n6727_));
  XOR2X1   g06471(.A(new_n6727_), .B(new_n6536_), .Y(new_n6728_));
  NAND2X1  g06472(.A(\b[57] ), .B(\b[56] ), .Y(new_n6729_));
  OAI21X1  g06473(.A0(new_n6521_), .A1(new_n6519_), .B0(new_n6729_), .Y(new_n6730_));
  XOR2X1   g06474(.A(\b[58] ), .B(\b[57] ), .Y(new_n6731_));
  XOR2X1   g06475(.A(new_n6731_), .B(new_n6730_), .Y(new_n6732_));
  AOI22X1  g06476(.A0(new_n267_), .A1(\b[58] ), .B0(new_n266_), .B1(\b[57] ), .Y(new_n6733_));
  OAI21X1  g06477(.A0(new_n350_), .A1(new_n6520_), .B0(new_n6733_), .Y(new_n6734_));
  AOI21X1  g06478(.A0(new_n6732_), .A1(new_n318_), .B0(new_n6734_), .Y(new_n6735_));
  XOR2X1   g06479(.A(new_n6735_), .B(\a[2] ), .Y(new_n6736_));
  XOR2X1   g06480(.A(new_n6736_), .B(new_n6728_), .Y(new_n6737_));
  NAND2X1  g06481(.A(new_n6527_), .B(new_n6517_), .Y(new_n6738_));
  OAI21X1  g06482(.A0(new_n6531_), .A1(new_n6530_), .B0(new_n6528_), .Y(new_n6739_));
  AND2X1   g06483(.A(new_n6739_), .B(new_n6738_), .Y(new_n6740_));
  XOR2X1   g06484(.A(new_n6740_), .B(new_n6737_), .Y(\f[58] ));
  AND2X1   g06485(.A(new_n6727_), .B(new_n6536_), .Y(new_n6742_));
  NOR2X1   g06486(.A(new_n6727_), .B(new_n6536_), .Y(new_n6743_));
  NOR3X1   g06487(.A(new_n6736_), .B(new_n6743_), .C(new_n6742_), .Y(new_n6744_));
  AOI21X1  g06488(.A0(new_n6739_), .A1(new_n6738_), .B0(new_n6737_), .Y(new_n6745_));
  OR2X1    g06489(.A(new_n6745_), .B(new_n6744_), .Y(new_n6746_));
  AND2X1   g06490(.A(new_n6726_), .B(new_n6540_), .Y(new_n6747_));
  OR2X1    g06491(.A(new_n6742_), .B(new_n6747_), .Y(new_n6748_));
  AND2X1   g06492(.A(new_n6724_), .B(new_n6547_), .Y(new_n6749_));
  AOI21X1  g06493(.A0(new_n6725_), .A1(new_n6543_), .B0(new_n6749_), .Y(new_n6750_));
  AOI22X1  g06494(.A0(new_n469_), .A1(\b[53] ), .B0(new_n468_), .B1(\b[52] ), .Y(new_n6751_));
  OAI21X1  g06495(.A0(new_n467_), .A1(new_n5787_), .B0(new_n6751_), .Y(new_n6752_));
  AOI21X1  g06496(.A0(new_n5786_), .A1(new_n404_), .B0(new_n6752_), .Y(new_n6753_));
  XOR2X1   g06497(.A(new_n6753_), .B(\a[8] ), .Y(new_n6754_));
  AND2X1   g06498(.A(new_n6722_), .B(new_n6562_), .Y(new_n6755_));
  AOI21X1  g06499(.A0(new_n6723_), .A1(new_n6558_), .B0(new_n6755_), .Y(new_n6756_));
  AND2X1   g06500(.A(new_n6720_), .B(new_n6715_), .Y(new_n6757_));
  AOI21X1  g06501(.A0(new_n6721_), .A1(new_n6565_), .B0(new_n6757_), .Y(new_n6758_));
  INVX1    g06502(.A(new_n6678_), .Y(new_n6759_));
  XOR2X1   g06503(.A(new_n6759_), .B(new_n6570_), .Y(new_n6760_));
  XOR2X1   g06504(.A(new_n6683_), .B(new_n6760_), .Y(new_n6761_));
  XOR2X1   g06505(.A(new_n6688_), .B(new_n6761_), .Y(new_n6762_));
  XOR2X1   g06506(.A(new_n6693_), .B(new_n6762_), .Y(new_n6763_));
  XOR2X1   g06507(.A(new_n6696_), .B(new_n6763_), .Y(new_n6764_));
  NOR2X1   g06508(.A(new_n6701_), .B(new_n6764_), .Y(new_n6765_));
  XOR2X1   g06509(.A(new_n6701_), .B(new_n6764_), .Y(new_n6766_));
  AOI21X1  g06510(.A0(new_n6705_), .A1(new_n6766_), .B0(new_n6765_), .Y(new_n6767_));
  INVX1    g06511(.A(new_n6673_), .Y(new_n6768_));
  NOR2X1   g06512(.A(new_n6677_), .B(new_n6768_), .Y(new_n6769_));
  AOI21X1  g06513(.A0(new_n6759_), .A1(new_n6570_), .B0(new_n6769_), .Y(new_n6770_));
  INVX1    g06514(.A(new_n6654_), .Y(new_n6771_));
  XOR2X1   g06515(.A(new_n6771_), .B(new_n6650_), .Y(new_n6772_));
  XOR2X1   g06516(.A(new_n6657_), .B(new_n6772_), .Y(new_n6773_));
  XOR2X1   g06517(.A(new_n6662_), .B(new_n6773_), .Y(new_n6774_));
  XOR2X1   g06518(.A(new_n6666_), .B(new_n6774_), .Y(new_n6775_));
  OR2X1    g06519(.A(new_n6671_), .B(new_n6775_), .Y(new_n6776_));
  OAI21X1  g06520(.A0(new_n6672_), .A1(new_n6572_), .B0(new_n6776_), .Y(new_n6777_));
  OR2X1    g06521(.A(new_n6654_), .B(new_n6650_), .Y(new_n6778_));
  OAI21X1  g06522(.A0(new_n6657_), .A1(new_n6772_), .B0(new_n6778_), .Y(new_n6779_));
  INVX1    g06523(.A(new_n6631_), .Y(new_n6780_));
  OR2X1    g06524(.A(new_n6635_), .B(new_n6780_), .Y(new_n6781_));
  OAI21X1  g06525(.A0(new_n6638_), .A1(new_n6636_), .B0(new_n6781_), .Y(new_n6782_));
  AOI22X1  g06526(.A0(new_n4095_), .A1(\b[17] ), .B0(new_n4094_), .B1(\b[16] ), .Y(new_n6783_));
  OAI21X1  g06527(.A0(new_n4233_), .A1(new_n977_), .B0(new_n6783_), .Y(new_n6784_));
  AOI21X1  g06528(.A0(new_n3901_), .A1(new_n976_), .B0(new_n6784_), .Y(new_n6785_));
  XOR2X1   g06529(.A(new_n6785_), .B(\a[44] ), .Y(new_n6786_));
  INVX1    g06530(.A(new_n6630_), .Y(new_n6787_));
  XOR2X1   g06531(.A(new_n6615_), .B(new_n4873_), .Y(new_n6788_));
  AND2X1   g06532(.A(new_n6788_), .B(new_n6612_), .Y(new_n6789_));
  NOR2X1   g06533(.A(new_n6619_), .B(new_n6617_), .Y(new_n6790_));
  OR2X1    g06534(.A(new_n6790_), .B(new_n6789_), .Y(new_n6791_));
  AOI22X1  g06535(.A0(new_n4880_), .A1(\b[11] ), .B0(new_n4877_), .B1(\b[10] ), .Y(new_n6792_));
  OAI21X1  g06536(.A0(new_n5291_), .A1(new_n590_), .B0(new_n6792_), .Y(new_n6793_));
  AOI21X1  g06537(.A0(new_n4875_), .A1(new_n589_), .B0(new_n6793_), .Y(new_n6794_));
  XOR2X1   g06538(.A(new_n6794_), .B(new_n4873_), .Y(new_n6795_));
  NAND2X1  g06539(.A(new_n6610_), .B(new_n6587_), .Y(new_n6796_));
  OAI21X1  g06540(.A0(new_n6581_), .A1(new_n6580_), .B0(new_n6611_), .Y(new_n6797_));
  NAND2X1  g06541(.A(new_n6797_), .B(new_n6796_), .Y(new_n6798_));
  AND2X1   g06542(.A(new_n6608_), .B(new_n6594_), .Y(new_n6799_));
  AND2X1   g06543(.A(new_n6609_), .B(new_n6589_), .Y(new_n6800_));
  OR2X1    g06544(.A(new_n6800_), .B(new_n6799_), .Y(new_n6801_));
  NOR2X1   g06545(.A(new_n6607_), .B(new_n6595_), .Y(new_n6802_));
  NOR3X1   g06546(.A(new_n6599_), .B(new_n6597_), .C(new_n6602_), .Y(new_n6803_));
  INVX1    g06547(.A(new_n6803_), .Y(new_n6804_));
  AOI22X1  g06548(.A0(new_n6603_), .A1(\b[2] ), .B0(new_n6600_), .B1(\b[1] ), .Y(new_n6805_));
  OAI21X1  g06549(.A0(new_n6804_), .A1(new_n274_), .B0(new_n6805_), .Y(new_n6806_));
  AOI21X1  g06550(.A0(new_n6598_), .A1(new_n341_), .B0(new_n6806_), .Y(new_n6807_));
  XOR2X1   g06551(.A(new_n6807_), .B(\a[59] ), .Y(new_n6808_));
  XOR2X1   g06552(.A(new_n6808_), .B(new_n6802_), .Y(new_n6809_));
  AOI22X1  g06553(.A0(new_n6438_), .A1(\b[5] ), .B0(new_n6437_), .B1(\b[4] ), .Y(new_n6810_));
  OAI21X1  g06554(.A0(new_n6436_), .A1(new_n297_), .B0(new_n6810_), .Y(new_n6811_));
  AOI21X1  g06555(.A0(new_n6023_), .A1(new_n349_), .B0(new_n6811_), .Y(new_n6812_));
  XOR2X1   g06556(.A(new_n6812_), .B(\a[56] ), .Y(new_n6813_));
  NAND2X1  g06557(.A(new_n6813_), .B(new_n6809_), .Y(new_n6814_));
  XOR2X1   g06558(.A(new_n6813_), .B(new_n6809_), .Y(new_n6815_));
  INVX1    g06559(.A(new_n6815_), .Y(new_n6816_));
  NOR2X1   g06560(.A(new_n6813_), .B(new_n6809_), .Y(new_n6817_));
  AOI21X1  g06561(.A0(new_n6814_), .A1(new_n6801_), .B0(new_n6817_), .Y(new_n6818_));
  AOI22X1  g06562(.A0(new_n6818_), .A1(new_n6814_), .B0(new_n6816_), .B1(new_n6801_), .Y(new_n6819_));
  AOI22X1  g06563(.A0(new_n5430_), .A1(\b[8] ), .B0(new_n5427_), .B1(\b[7] ), .Y(new_n6820_));
  OAI21X1  g06564(.A0(new_n5891_), .A1(new_n392_), .B0(new_n6820_), .Y(new_n6821_));
  AOI21X1  g06565(.A0(new_n5425_), .A1(new_n454_), .B0(new_n6821_), .Y(new_n6822_));
  XOR2X1   g06566(.A(new_n6822_), .B(\a[53] ), .Y(new_n6823_));
  XOR2X1   g06567(.A(new_n6823_), .B(new_n6819_), .Y(new_n6824_));
  XOR2X1   g06568(.A(new_n6824_), .B(new_n6798_), .Y(new_n6825_));
  XOR2X1   g06569(.A(new_n6825_), .B(new_n6795_), .Y(new_n6826_));
  XOR2X1   g06570(.A(new_n6826_), .B(new_n6791_), .Y(new_n6827_));
  AOI22X1  g06571(.A0(new_n4572_), .A1(\b[14] ), .B0(new_n4571_), .B1(\b[13] ), .Y(new_n6828_));
  OAI21X1  g06572(.A0(new_n4740_), .A1(new_n713_), .B0(new_n6828_), .Y(new_n6829_));
  AOI21X1  g06573(.A0(new_n4375_), .A1(new_n734_), .B0(new_n6829_), .Y(new_n6830_));
  XOR2X1   g06574(.A(new_n6830_), .B(\a[47] ), .Y(new_n6831_));
  XOR2X1   g06575(.A(new_n6831_), .B(new_n6827_), .Y(new_n6832_));
  XOR2X1   g06576(.A(new_n6832_), .B(new_n6787_), .Y(new_n6833_));
  XOR2X1   g06577(.A(new_n6833_), .B(new_n6786_), .Y(new_n6834_));
  XOR2X1   g06578(.A(new_n6834_), .B(new_n6782_), .Y(new_n6835_));
  AOI22X1  g06579(.A0(new_n3652_), .A1(\b[20] ), .B0(new_n3651_), .B1(\b[19] ), .Y(new_n6836_));
  OAI21X1  g06580(.A0(new_n3778_), .A1(new_n1115_), .B0(new_n6836_), .Y(new_n6837_));
  AOI21X1  g06581(.A0(new_n3480_), .A1(new_n1217_), .B0(new_n6837_), .Y(new_n6838_));
  XOR2X1   g06582(.A(new_n6838_), .B(\a[41] ), .Y(new_n6839_));
  INVX1    g06583(.A(new_n6839_), .Y(new_n6840_));
  XOR2X1   g06584(.A(new_n6840_), .B(new_n6835_), .Y(new_n6841_));
  XOR2X1   g06585(.A(new_n6841_), .B(new_n6649_), .Y(new_n6842_));
  AOI22X1  g06586(.A0(new_n3204_), .A1(\b[23] ), .B0(new_n3203_), .B1(\b[22] ), .Y(new_n6843_));
  OAI21X1  g06587(.A0(new_n3321_), .A1(new_n1482_), .B0(new_n6843_), .Y(new_n6844_));
  AOI21X1  g06588(.A0(new_n3080_), .A1(new_n1481_), .B0(new_n6844_), .Y(new_n6845_));
  XOR2X1   g06589(.A(new_n6845_), .B(\a[38] ), .Y(new_n6846_));
  XOR2X1   g06590(.A(new_n6846_), .B(new_n6842_), .Y(new_n6847_));
  XOR2X1   g06591(.A(new_n6847_), .B(new_n6779_), .Y(new_n6848_));
  AOI22X1  g06592(.A0(new_n2813_), .A1(\b[26] ), .B0(new_n2812_), .B1(\b[25] ), .Y(new_n6849_));
  OAI21X1  g06593(.A0(new_n2946_), .A1(new_n1588_), .B0(new_n6849_), .Y(new_n6850_));
  AOI21X1  g06594(.A0(new_n2652_), .A1(new_n1783_), .B0(new_n6850_), .Y(new_n6851_));
  XOR2X1   g06595(.A(new_n6851_), .B(\a[35] ), .Y(new_n6852_));
  XOR2X1   g06596(.A(new_n6852_), .B(new_n6848_), .Y(new_n6853_));
  NOR2X1   g06597(.A(new_n6662_), .B(new_n6658_), .Y(new_n6854_));
  AOI21X1  g06598(.A0(new_n6666_), .A1(new_n6663_), .B0(new_n6854_), .Y(new_n6855_));
  XOR2X1   g06599(.A(new_n6855_), .B(new_n6853_), .Y(new_n6856_));
  AOI22X1  g06600(.A0(new_n2545_), .A1(\b[29] ), .B0(new_n2544_), .B1(\b[28] ), .Y(new_n6857_));
  OAI21X1  g06601(.A0(new_n2543_), .A1(new_n2126_), .B0(new_n6857_), .Y(new_n6858_));
  AOI21X1  g06602(.A0(new_n2260_), .A1(new_n2125_), .B0(new_n6858_), .Y(new_n6859_));
  XOR2X1   g06603(.A(new_n6859_), .B(\a[32] ), .Y(new_n6860_));
  NAND2X1  g06604(.A(new_n6860_), .B(new_n6856_), .Y(new_n6861_));
  INVX1    g06605(.A(new_n6847_), .Y(new_n6862_));
  XOR2X1   g06606(.A(new_n6862_), .B(new_n6779_), .Y(new_n6863_));
  XOR2X1   g06607(.A(new_n6852_), .B(new_n6863_), .Y(new_n6864_));
  XOR2X1   g06608(.A(new_n6855_), .B(new_n6864_), .Y(new_n6865_));
  XOR2X1   g06609(.A(new_n6860_), .B(new_n6865_), .Y(new_n6866_));
  NOR2X1   g06610(.A(new_n6860_), .B(new_n6856_), .Y(new_n6867_));
  AOI21X1  g06611(.A0(new_n6861_), .A1(new_n6777_), .B0(new_n6867_), .Y(new_n6868_));
  AOI22X1  g06612(.A0(new_n6868_), .A1(new_n6861_), .B0(new_n6866_), .B1(new_n6777_), .Y(new_n6869_));
  AOI22X1  g06613(.A0(new_n2163_), .A1(\b[32] ), .B0(new_n2162_), .B1(\b[31] ), .Y(new_n6870_));
  OAI21X1  g06614(.A0(new_n2161_), .A1(new_n2356_), .B0(new_n6870_), .Y(new_n6871_));
  AOI21X1  g06615(.A0(new_n2495_), .A1(new_n1907_), .B0(new_n6871_), .Y(new_n6872_));
  XOR2X1   g06616(.A(new_n6872_), .B(\a[29] ), .Y(new_n6873_));
  INVX1    g06617(.A(new_n6873_), .Y(new_n6874_));
  XOR2X1   g06618(.A(new_n6874_), .B(new_n6869_), .Y(new_n6875_));
  XOR2X1   g06619(.A(new_n6875_), .B(new_n6770_), .Y(new_n6876_));
  AOI22X1  g06620(.A0(new_n1814_), .A1(\b[35] ), .B0(new_n1813_), .B1(\b[34] ), .Y(new_n6877_));
  OAI21X1  g06621(.A0(new_n1812_), .A1(new_n2893_), .B0(new_n6877_), .Y(new_n6878_));
  AOI21X1  g06622(.A0(new_n2892_), .A1(new_n1617_), .B0(new_n6878_), .Y(new_n6879_));
  XOR2X1   g06623(.A(new_n6879_), .B(\a[26] ), .Y(new_n6880_));
  XOR2X1   g06624(.A(new_n6880_), .B(new_n6876_), .Y(new_n6881_));
  NOR2X1   g06625(.A(new_n6683_), .B(new_n6679_), .Y(new_n6882_));
  AOI21X1  g06626(.A0(new_n6688_), .A1(new_n6684_), .B0(new_n6882_), .Y(new_n6883_));
  XOR2X1   g06627(.A(new_n6883_), .B(new_n6881_), .Y(new_n6884_));
  AOI22X1  g06628(.A0(new_n1526_), .A1(\b[38] ), .B0(new_n1525_), .B1(\b[37] ), .Y(new_n6885_));
  OAI21X1  g06629(.A0(new_n1524_), .A1(new_n3276_), .B0(new_n6885_), .Y(new_n6886_));
  AOI21X1  g06630(.A0(new_n3275_), .A1(new_n1347_), .B0(new_n6886_), .Y(new_n6887_));
  XOR2X1   g06631(.A(new_n6887_), .B(\a[23] ), .Y(new_n6888_));
  XOR2X1   g06632(.A(new_n6888_), .B(new_n6884_), .Y(new_n6889_));
  OR2X1    g06633(.A(new_n6693_), .B(new_n6762_), .Y(new_n6890_));
  OAI21X1  g06634(.A0(new_n6696_), .A1(new_n6694_), .B0(new_n6890_), .Y(new_n6891_));
  XOR2X1   g06635(.A(new_n6891_), .B(new_n6889_), .Y(new_n6892_));
  AOI22X1  g06636(.A0(new_n1263_), .A1(\b[41] ), .B0(new_n1262_), .B1(\b[40] ), .Y(new_n6893_));
  OAI21X1  g06637(.A0(new_n1261_), .A1(new_n3723_), .B0(new_n6893_), .Y(new_n6894_));
  AOI21X1  g06638(.A0(new_n3722_), .A1(new_n1075_), .B0(new_n6894_), .Y(new_n6895_));
  XOR2X1   g06639(.A(new_n6895_), .B(\a[20] ), .Y(new_n6896_));
  AND2X1   g06640(.A(new_n6896_), .B(new_n6892_), .Y(new_n6897_));
  XOR2X1   g06641(.A(new_n6896_), .B(new_n6892_), .Y(new_n6898_));
  OR2X1    g06642(.A(new_n6896_), .B(new_n6892_), .Y(new_n6899_));
  OAI21X1  g06643(.A0(new_n6897_), .A1(new_n6767_), .B0(new_n6899_), .Y(new_n6900_));
  OAI22X1  g06644(.A0(new_n6900_), .A1(new_n6897_), .B0(new_n6898_), .B1(new_n6767_), .Y(new_n6901_));
  AOI22X1  g06645(.A0(new_n1017_), .A1(\b[44] ), .B0(new_n1016_), .B1(\b[43] ), .Y(new_n6902_));
  OAI21X1  g06646(.A0(new_n1015_), .A1(new_n4012_), .B0(new_n6902_), .Y(new_n6903_));
  AOI21X1  g06647(.A0(new_n4178_), .A1(new_n882_), .B0(new_n6903_), .Y(new_n6904_));
  XOR2X1   g06648(.A(new_n6904_), .B(\a[17] ), .Y(new_n6905_));
  XOR2X1   g06649(.A(new_n6905_), .B(new_n6901_), .Y(new_n6906_));
  XOR2X1   g06650(.A(new_n6906_), .B(new_n6714_), .Y(new_n6907_));
  AOI22X1  g06651(.A0(new_n818_), .A1(\b[47] ), .B0(new_n817_), .B1(\b[46] ), .Y(new_n6908_));
  OAI21X1  g06652(.A0(new_n816_), .A1(new_n4674_), .B0(new_n6908_), .Y(new_n6909_));
  AOI21X1  g06653(.A0(new_n4673_), .A1(new_n668_), .B0(new_n6909_), .Y(new_n6910_));
  XOR2X1   g06654(.A(new_n6910_), .B(\a[14] ), .Y(new_n6911_));
  XOR2X1   g06655(.A(new_n6911_), .B(new_n6907_), .Y(new_n6912_));
  XOR2X1   g06656(.A(new_n6912_), .B(new_n6758_), .Y(new_n6913_));
  AOI22X1  g06657(.A0(new_n603_), .A1(\b[50] ), .B0(new_n602_), .B1(\b[49] ), .Y(new_n6914_));
  OAI21X1  g06658(.A0(new_n601_), .A1(new_n5036_), .B0(new_n6914_), .Y(new_n6915_));
  AOI21X1  g06659(.A0(new_n5204_), .A1(new_n518_), .B0(new_n6915_), .Y(new_n6916_));
  XOR2X1   g06660(.A(new_n6916_), .B(\a[11] ), .Y(new_n6917_));
  INVX1    g06661(.A(new_n6917_), .Y(new_n6918_));
  XOR2X1   g06662(.A(new_n6918_), .B(new_n6913_), .Y(new_n6919_));
  XOR2X1   g06663(.A(new_n6919_), .B(new_n6756_), .Y(new_n6920_));
  XOR2X1   g06664(.A(new_n6920_), .B(new_n6754_), .Y(new_n6921_));
  XOR2X1   g06665(.A(new_n6921_), .B(new_n6750_), .Y(new_n6922_));
  AOI22X1  g06666(.A0(new_n369_), .A1(\b[56] ), .B0(new_n368_), .B1(\b[55] ), .Y(new_n6923_));
  OAI21X1  g06667(.A0(new_n367_), .A1(new_n6148_), .B0(new_n6923_), .Y(new_n6924_));
  AOI21X1  g06668(.A0(new_n6342_), .A1(new_n308_), .B0(new_n6924_), .Y(new_n6925_));
  XOR2X1   g06669(.A(new_n6925_), .B(\a[5] ), .Y(new_n6926_));
  XOR2X1   g06670(.A(new_n6926_), .B(new_n6922_), .Y(new_n6927_));
  AND2X1   g06671(.A(\b[58] ), .B(\b[57] ), .Y(new_n6928_));
  AOI21X1  g06672(.A0(new_n6731_), .A1(new_n6730_), .B0(new_n6928_), .Y(new_n6929_));
  INVX1    g06673(.A(\b[58] ), .Y(new_n6930_));
  XOR2X1   g06674(.A(\b[59] ), .B(new_n6930_), .Y(new_n6931_));
  XOR2X1   g06675(.A(new_n6931_), .B(new_n6929_), .Y(new_n6932_));
  INVX1    g06676(.A(\b[57] ), .Y(new_n6933_));
  AOI22X1  g06677(.A0(new_n267_), .A1(\b[59] ), .B0(new_n266_), .B1(\b[58] ), .Y(new_n6934_));
  OAI21X1  g06678(.A0(new_n350_), .A1(new_n6933_), .B0(new_n6934_), .Y(new_n6935_));
  AOI21X1  g06679(.A0(new_n6932_), .A1(new_n318_), .B0(new_n6935_), .Y(new_n6936_));
  XOR2X1   g06680(.A(new_n6936_), .B(\a[2] ), .Y(new_n6937_));
  XOR2X1   g06681(.A(new_n6937_), .B(new_n6927_), .Y(new_n6938_));
  XOR2X1   g06682(.A(new_n6938_), .B(new_n6748_), .Y(new_n6939_));
  XOR2X1   g06683(.A(new_n6939_), .B(new_n6746_), .Y(\f[59] ));
  NAND2X1  g06684(.A(new_n6938_), .B(new_n6748_), .Y(new_n6941_));
  OAI21X1  g06685(.A0(new_n6745_), .A1(new_n6744_), .B0(new_n6939_), .Y(new_n6942_));
  AND2X1   g06686(.A(new_n6942_), .B(new_n6941_), .Y(new_n6943_));
  XOR2X1   g06687(.A(new_n6925_), .B(new_n305_), .Y(new_n6944_));
  NAND2X1  g06688(.A(new_n6944_), .B(new_n6922_), .Y(new_n6945_));
  OR2X1    g06689(.A(new_n6937_), .B(new_n6927_), .Y(new_n6946_));
  AND2X1   g06690(.A(new_n6946_), .B(new_n6945_), .Y(new_n6947_));
  NAND2X1  g06691(.A(\b[59] ), .B(\b[58] ), .Y(new_n6948_));
  OAI21X1  g06692(.A0(new_n6931_), .A1(new_n6929_), .B0(new_n6948_), .Y(new_n6949_));
  XOR2X1   g06693(.A(\b[60] ), .B(\b[59] ), .Y(new_n6950_));
  XOR2X1   g06694(.A(new_n6950_), .B(new_n6949_), .Y(new_n6951_));
  AOI22X1  g06695(.A0(new_n267_), .A1(\b[60] ), .B0(new_n266_), .B1(\b[59] ), .Y(new_n6952_));
  OAI21X1  g06696(.A0(new_n350_), .A1(new_n6930_), .B0(new_n6952_), .Y(new_n6953_));
  AOI21X1  g06697(.A0(new_n6951_), .A1(new_n318_), .B0(new_n6953_), .Y(new_n6954_));
  XOR2X1   g06698(.A(new_n6954_), .B(new_n257_), .Y(new_n6955_));
  AOI22X1  g06699(.A0(new_n369_), .A1(\b[57] ), .B0(new_n368_), .B1(\b[56] ), .Y(new_n6956_));
  OAI21X1  g06700(.A0(new_n367_), .A1(new_n6523_), .B0(new_n6956_), .Y(new_n6957_));
  AOI21X1  g06701(.A0(new_n6522_), .A1(new_n308_), .B0(new_n6957_), .Y(new_n6958_));
  XOR2X1   g06702(.A(new_n6958_), .B(new_n305_), .Y(new_n6959_));
  INVX1    g06703(.A(new_n6754_), .Y(new_n6960_));
  NAND2X1  g06704(.A(new_n6920_), .B(new_n6960_), .Y(new_n6961_));
  OAI21X1  g06705(.A0(new_n6921_), .A1(new_n6750_), .B0(new_n6961_), .Y(new_n6962_));
  AOI22X1  g06706(.A0(new_n469_), .A1(\b[54] ), .B0(new_n468_), .B1(\b[53] ), .Y(new_n6963_));
  OAI21X1  g06707(.A0(new_n467_), .A1(new_n5808_), .B0(new_n6963_), .Y(new_n6964_));
  AOI21X1  g06708(.A0(new_n5807_), .A1(new_n404_), .B0(new_n6964_), .Y(new_n6965_));
  XOR2X1   g06709(.A(new_n6965_), .B(new_n400_), .Y(new_n6966_));
  AND2X1   g06710(.A(new_n6511_), .B(new_n6371_), .Y(new_n6967_));
  AOI21X1  g06711(.A0(new_n6512_), .A1(new_n6366_), .B0(new_n6967_), .Y(new_n6968_));
  NOR2X1   g06712(.A(new_n6722_), .B(new_n6562_), .Y(new_n6969_));
  NAND2X1  g06713(.A(new_n6722_), .B(new_n6562_), .Y(new_n6970_));
  OAI21X1  g06714(.A0(new_n6969_), .A1(new_n6968_), .B0(new_n6970_), .Y(new_n6971_));
  NOR2X1   g06715(.A(new_n6917_), .B(new_n6913_), .Y(new_n6972_));
  XOR2X1   g06716(.A(new_n6917_), .B(new_n6913_), .Y(new_n6973_));
  AOI21X1  g06717(.A0(new_n6973_), .A1(new_n6971_), .B0(new_n6972_), .Y(new_n6974_));
  AOI22X1  g06718(.A0(new_n603_), .A1(\b[51] ), .B0(new_n602_), .B1(\b[50] ), .Y(new_n6975_));
  OAI21X1  g06719(.A0(new_n601_), .A1(new_n5237_), .B0(new_n6975_), .Y(new_n6976_));
  AOI21X1  g06720(.A0(new_n5236_), .A1(new_n518_), .B0(new_n6976_), .Y(new_n6977_));
  XOR2X1   g06721(.A(new_n6977_), .B(\a[11] ), .Y(new_n6978_));
  OR2X1    g06722(.A(new_n6911_), .B(new_n6907_), .Y(new_n6979_));
  AND2X1   g06723(.A(new_n6721_), .B(new_n6565_), .Y(new_n6980_));
  OAI21X1  g06724(.A0(new_n6980_), .A1(new_n6757_), .B0(new_n6912_), .Y(new_n6981_));
  AND2X1   g06725(.A(new_n6981_), .B(new_n6979_), .Y(new_n6982_));
  AOI22X1  g06726(.A0(new_n818_), .A1(\b[48] ), .B0(new_n817_), .B1(\b[47] ), .Y(new_n6983_));
  OAI21X1  g06727(.A0(new_n816_), .A1(new_n4693_), .B0(new_n6983_), .Y(new_n6984_));
  AOI21X1  g06728(.A0(new_n4692_), .A1(new_n668_), .B0(new_n6984_), .Y(new_n6985_));
  XOR2X1   g06729(.A(new_n6985_), .B(\a[14] ), .Y(new_n6986_));
  XOR2X1   g06730(.A(new_n6904_), .B(new_n879_), .Y(new_n6987_));
  AND2X1   g06731(.A(new_n6987_), .B(new_n6901_), .Y(new_n6988_));
  XOR2X1   g06732(.A(new_n6987_), .B(new_n6901_), .Y(new_n6989_));
  AOI21X1  g06733(.A0(new_n6989_), .A1(new_n6714_), .B0(new_n6988_), .Y(new_n6990_));
  AOI22X1  g06734(.A0(new_n1017_), .A1(\b[45] ), .B0(new_n1016_), .B1(\b[44] ), .Y(new_n6991_));
  OAI21X1  g06735(.A0(new_n1015_), .A1(new_n4339_), .B0(new_n6991_), .Y(new_n6992_));
  AOI21X1  g06736(.A0(new_n4338_), .A1(new_n882_), .B0(new_n6992_), .Y(new_n6993_));
  XOR2X1   g06737(.A(new_n6993_), .B(\a[17] ), .Y(new_n6994_));
  INVX1    g06738(.A(new_n6994_), .Y(new_n6995_));
  XOR2X1   g06739(.A(new_n6873_), .B(new_n6869_), .Y(new_n6996_));
  XOR2X1   g06740(.A(new_n6996_), .B(new_n6770_), .Y(new_n6997_));
  OR2X1    g06741(.A(new_n6880_), .B(new_n6997_), .Y(new_n6998_));
  OAI21X1  g06742(.A0(new_n6883_), .A1(new_n6881_), .B0(new_n6998_), .Y(new_n6999_));
  OR2X1    g06743(.A(new_n6873_), .B(new_n6869_), .Y(new_n7000_));
  OAI21X1  g06744(.A0(new_n6875_), .A1(new_n6770_), .B0(new_n7000_), .Y(new_n7001_));
  OR2X1    g06745(.A(new_n6839_), .B(new_n6835_), .Y(new_n7002_));
  OAI21X1  g06746(.A0(new_n6841_), .A1(new_n6649_), .B0(new_n7002_), .Y(new_n7003_));
  AOI22X1  g06747(.A0(new_n3652_), .A1(\b[21] ), .B0(new_n3651_), .B1(\b[20] ), .Y(new_n7004_));
  OAI21X1  g06748(.A0(new_n3778_), .A1(new_n1300_), .B0(new_n7004_), .Y(new_n7005_));
  AOI21X1  g06749(.A0(new_n3480_), .A1(new_n1299_), .B0(new_n7005_), .Y(new_n7006_));
  XOR2X1   g06750(.A(new_n7006_), .B(new_n3478_), .Y(new_n7007_));
  XOR2X1   g06751(.A(new_n6832_), .B(new_n6630_), .Y(new_n7008_));
  NOR2X1   g06752(.A(new_n7008_), .B(new_n6786_), .Y(new_n7009_));
  INVX1    g06753(.A(new_n6834_), .Y(new_n7010_));
  AOI21X1  g06754(.A0(new_n7010_), .A1(new_n6782_), .B0(new_n7009_), .Y(new_n7011_));
  AOI22X1  g06755(.A0(new_n4095_), .A1(\b[18] ), .B0(new_n4094_), .B1(\b[17] ), .Y(new_n7012_));
  OAI21X1  g06756(.A0(new_n4233_), .A1(new_n974_), .B0(new_n7012_), .Y(new_n7013_));
  AOI21X1  g06757(.A0(new_n3901_), .A1(new_n1042_), .B0(new_n7013_), .Y(new_n7014_));
  XOR2X1   g06758(.A(new_n7014_), .B(\a[44] ), .Y(new_n7015_));
  XOR2X1   g06759(.A(new_n6830_), .B(new_n4568_), .Y(new_n7016_));
  NAND2X1  g06760(.A(new_n7016_), .B(new_n6827_), .Y(new_n7017_));
  OAI21X1  g06761(.A0(new_n6832_), .A1(new_n6787_), .B0(new_n7017_), .Y(new_n7018_));
  AOI22X1  g06762(.A0(new_n4572_), .A1(\b[15] ), .B0(new_n4571_), .B1(\b[14] ), .Y(new_n7019_));
  OAI21X1  g06763(.A0(new_n4740_), .A1(new_n795_), .B0(new_n7019_), .Y(new_n7020_));
  AOI21X1  g06764(.A0(new_n4375_), .A1(new_n794_), .B0(new_n7020_), .Y(new_n7021_));
  XOR2X1   g06765(.A(new_n7021_), .B(new_n4568_), .Y(new_n7022_));
  AND2X1   g06766(.A(new_n6825_), .B(new_n6795_), .Y(new_n7023_));
  AOI21X1  g06767(.A0(new_n6826_), .A1(new_n6791_), .B0(new_n7023_), .Y(new_n7024_));
  AOI22X1  g06768(.A0(new_n4880_), .A1(\b[12] ), .B0(new_n4877_), .B1(\b[11] ), .Y(new_n7025_));
  OAI21X1  g06769(.A0(new_n5291_), .A1(new_n587_), .B0(new_n7025_), .Y(new_n7026_));
  AOI21X1  g06770(.A0(new_n4875_), .A1(new_n635_), .B0(new_n7026_), .Y(new_n7027_));
  XOR2X1   g06771(.A(new_n7027_), .B(\a[50] ), .Y(new_n7028_));
  INVX1    g06772(.A(new_n7028_), .Y(new_n7029_));
  NAND2X1  g06773(.A(new_n6824_), .B(new_n6798_), .Y(new_n7030_));
  OAI21X1  g06774(.A0(new_n6823_), .A1(new_n6819_), .B0(new_n7030_), .Y(new_n7031_));
  NOR3X1   g06775(.A(new_n6808_), .B(new_n6607_), .C(new_n6595_), .Y(new_n7032_));
  XOR2X1   g06776(.A(\a[60] ), .B(new_n6596_), .Y(new_n7033_));
  NOR2X1   g06777(.A(new_n7033_), .B(new_n274_), .Y(new_n7034_));
  INVX1    g06778(.A(new_n7034_), .Y(new_n7035_));
  XOR2X1   g06779(.A(new_n7035_), .B(new_n7032_), .Y(new_n7036_));
  AOI22X1  g06780(.A0(new_n6603_), .A1(\b[3] ), .B0(new_n6600_), .B1(\b[2] ), .Y(new_n7037_));
  OAI21X1  g06781(.A0(new_n6804_), .A1(new_n275_), .B0(new_n7037_), .Y(new_n7038_));
  AOI21X1  g06782(.A0(new_n6598_), .A1(new_n366_), .B0(new_n7038_), .Y(new_n7039_));
  XOR2X1   g06783(.A(new_n7039_), .B(\a[59] ), .Y(new_n7040_));
  XOR2X1   g06784(.A(new_n7040_), .B(new_n7036_), .Y(new_n7041_));
  AOI22X1  g06785(.A0(new_n6438_), .A1(\b[6] ), .B0(new_n6437_), .B1(\b[5] ), .Y(new_n7042_));
  OAI21X1  g06786(.A0(new_n6436_), .A1(new_n325_), .B0(new_n7042_), .Y(new_n7043_));
  AOI21X1  g06787(.A0(new_n6023_), .A1(new_n378_), .B0(new_n7043_), .Y(new_n7044_));
  XOR2X1   g06788(.A(new_n7044_), .B(\a[56] ), .Y(new_n7045_));
  XOR2X1   g06789(.A(new_n7045_), .B(new_n7041_), .Y(new_n7046_));
  INVX1    g06790(.A(new_n7046_), .Y(new_n7047_));
  XOR2X1   g06791(.A(new_n7047_), .B(new_n6818_), .Y(new_n7048_));
  AOI22X1  g06792(.A0(new_n5430_), .A1(\b[9] ), .B0(new_n5427_), .B1(\b[8] ), .Y(new_n7049_));
  OAI21X1  g06793(.A0(new_n5891_), .A1(new_n492_), .B0(new_n7049_), .Y(new_n7050_));
  AOI21X1  g06794(.A0(new_n5425_), .A1(new_n491_), .B0(new_n7050_), .Y(new_n7051_));
  XOR2X1   g06795(.A(new_n7051_), .B(\a[53] ), .Y(new_n7052_));
  XOR2X1   g06796(.A(new_n7052_), .B(new_n7048_), .Y(new_n7053_));
  XOR2X1   g06797(.A(new_n7053_), .B(new_n7031_), .Y(new_n7054_));
  XOR2X1   g06798(.A(new_n7054_), .B(new_n7029_), .Y(new_n7055_));
  INVX1    g06799(.A(new_n7055_), .Y(new_n7056_));
  XOR2X1   g06800(.A(new_n7056_), .B(new_n7024_), .Y(new_n7057_));
  XOR2X1   g06801(.A(new_n7057_), .B(new_n7022_), .Y(new_n7058_));
  XOR2X1   g06802(.A(new_n7058_), .B(new_n7018_), .Y(new_n7059_));
  XOR2X1   g06803(.A(new_n7059_), .B(new_n7015_), .Y(new_n7060_));
  XOR2X1   g06804(.A(new_n7060_), .B(new_n7011_), .Y(new_n7061_));
  XOR2X1   g06805(.A(new_n7061_), .B(new_n7007_), .Y(new_n7062_));
  XOR2X1   g06806(.A(new_n7062_), .B(new_n7003_), .Y(new_n7063_));
  AOI22X1  g06807(.A0(new_n3204_), .A1(\b[24] ), .B0(new_n3203_), .B1(\b[23] ), .Y(new_n7064_));
  OAI21X1  g06808(.A0(new_n3321_), .A1(new_n1479_), .B0(new_n7064_), .Y(new_n7065_));
  AOI21X1  g06809(.A0(new_n3080_), .A1(new_n1572_), .B0(new_n7065_), .Y(new_n7066_));
  XOR2X1   g06810(.A(new_n7066_), .B(\a[38] ), .Y(new_n7067_));
  XOR2X1   g06811(.A(new_n7067_), .B(new_n7063_), .Y(new_n7068_));
  INVX1    g06812(.A(new_n7068_), .Y(new_n7069_));
  XOR2X1   g06813(.A(new_n6845_), .B(new_n3078_), .Y(new_n7070_));
  AND2X1   g06814(.A(new_n7070_), .B(new_n6842_), .Y(new_n7071_));
  AOI21X1  g06815(.A0(new_n6862_), .A1(new_n6779_), .B0(new_n7071_), .Y(new_n7072_));
  XOR2X1   g06816(.A(new_n7072_), .B(new_n7069_), .Y(new_n7073_));
  AOI22X1  g06817(.A0(new_n2813_), .A1(\b[27] ), .B0(new_n2812_), .B1(\b[26] ), .Y(new_n7074_));
  OAI21X1  g06818(.A0(new_n2946_), .A1(new_n1880_), .B0(new_n7074_), .Y(new_n7075_));
  AOI21X1  g06819(.A0(new_n2652_), .A1(new_n1879_), .B0(new_n7075_), .Y(new_n7076_));
  XOR2X1   g06820(.A(new_n7076_), .B(\a[35] ), .Y(new_n7077_));
  XOR2X1   g06821(.A(new_n7077_), .B(new_n7073_), .Y(new_n7078_));
  OR2X1    g06822(.A(new_n6852_), .B(new_n6848_), .Y(new_n7079_));
  OAI21X1  g06823(.A0(new_n6855_), .A1(new_n6864_), .B0(new_n7079_), .Y(new_n7080_));
  XOR2X1   g06824(.A(new_n7080_), .B(new_n7078_), .Y(new_n7081_));
  AOI22X1  g06825(.A0(new_n2545_), .A1(\b[30] ), .B0(new_n2544_), .B1(\b[29] ), .Y(new_n7082_));
  OAI21X1  g06826(.A0(new_n2543_), .A1(new_n2231_), .B0(new_n7082_), .Y(new_n7083_));
  AOI21X1  g06827(.A0(new_n2260_), .A1(new_n2230_), .B0(new_n7083_), .Y(new_n7084_));
  XOR2X1   g06828(.A(new_n7084_), .B(\a[32] ), .Y(new_n7085_));
  XOR2X1   g06829(.A(new_n7085_), .B(new_n7081_), .Y(new_n7086_));
  XOR2X1   g06830(.A(new_n7086_), .B(new_n6868_), .Y(new_n7087_));
  AOI22X1  g06831(.A0(new_n2163_), .A1(\b[33] ), .B0(new_n2162_), .B1(\b[32] ), .Y(new_n7088_));
  OAI21X1  g06832(.A0(new_n2161_), .A1(new_n2615_), .B0(new_n7088_), .Y(new_n7089_));
  AOI21X1  g06833(.A0(new_n2614_), .A1(new_n1907_), .B0(new_n7089_), .Y(new_n7090_));
  XOR2X1   g06834(.A(new_n7090_), .B(\a[29] ), .Y(new_n7091_));
  XOR2X1   g06835(.A(new_n7091_), .B(new_n7087_), .Y(new_n7092_));
  XOR2X1   g06836(.A(new_n7092_), .B(new_n7001_), .Y(new_n7093_));
  AOI22X1  g06837(.A0(new_n1814_), .A1(\b[36] ), .B0(new_n1813_), .B1(\b[35] ), .Y(new_n7094_));
  OAI21X1  g06838(.A0(new_n1812_), .A1(new_n2890_), .B0(new_n7094_), .Y(new_n7095_));
  AOI21X1  g06839(.A0(new_n3015_), .A1(new_n1617_), .B0(new_n7095_), .Y(new_n7096_));
  XOR2X1   g06840(.A(new_n7096_), .B(\a[26] ), .Y(new_n7097_));
  XOR2X1   g06841(.A(new_n7097_), .B(new_n7093_), .Y(new_n7098_));
  XOR2X1   g06842(.A(new_n7098_), .B(new_n6999_), .Y(new_n7099_));
  AOI22X1  g06843(.A0(new_n1526_), .A1(\b[39] ), .B0(new_n1525_), .B1(\b[38] ), .Y(new_n7100_));
  OAI21X1  g06844(.A0(new_n1524_), .A1(new_n3413_), .B0(new_n7100_), .Y(new_n7101_));
  AOI21X1  g06845(.A0(new_n3412_), .A1(new_n1347_), .B0(new_n7101_), .Y(new_n7102_));
  XOR2X1   g06846(.A(new_n7102_), .B(\a[23] ), .Y(new_n7103_));
  INVX1    g06847(.A(new_n7103_), .Y(new_n7104_));
  XOR2X1   g06848(.A(new_n7104_), .B(new_n7099_), .Y(new_n7105_));
  XOR2X1   g06849(.A(new_n6880_), .B(new_n6997_), .Y(new_n7106_));
  XOR2X1   g06850(.A(new_n6883_), .B(new_n7106_), .Y(new_n7107_));
  NOR2X1   g06851(.A(new_n6888_), .B(new_n7107_), .Y(new_n7108_));
  XOR2X1   g06852(.A(new_n6888_), .B(new_n7107_), .Y(new_n7109_));
  AOI21X1  g06853(.A0(new_n6891_), .A1(new_n7109_), .B0(new_n7108_), .Y(new_n7110_));
  XOR2X1   g06854(.A(new_n7110_), .B(new_n7105_), .Y(new_n7111_));
  AOI22X1  g06855(.A0(new_n1263_), .A1(\b[42] ), .B0(new_n1262_), .B1(\b[41] ), .Y(new_n7112_));
  OAI21X1  g06856(.A0(new_n1261_), .A1(new_n3720_), .B0(new_n7112_), .Y(new_n7113_));
  AOI21X1  g06857(.A0(new_n3860_), .A1(new_n1075_), .B0(new_n7113_), .Y(new_n7114_));
  XOR2X1   g06858(.A(new_n7114_), .B(\a[20] ), .Y(new_n7115_));
  XOR2X1   g06859(.A(new_n7115_), .B(new_n7111_), .Y(new_n7116_));
  XOR2X1   g06860(.A(new_n7116_), .B(new_n6900_), .Y(new_n7117_));
  XOR2X1   g06861(.A(new_n7117_), .B(new_n6995_), .Y(new_n7118_));
  INVX1    g06862(.A(new_n7118_), .Y(new_n7119_));
  XOR2X1   g06863(.A(new_n7119_), .B(new_n6990_), .Y(new_n7120_));
  XOR2X1   g06864(.A(new_n7120_), .B(new_n6986_), .Y(new_n7121_));
  XOR2X1   g06865(.A(new_n7121_), .B(new_n6982_), .Y(new_n7122_));
  XOR2X1   g06866(.A(new_n7122_), .B(new_n6978_), .Y(new_n7123_));
  XOR2X1   g06867(.A(new_n7123_), .B(new_n6974_), .Y(new_n7124_));
  XOR2X1   g06868(.A(new_n7124_), .B(new_n6966_), .Y(new_n7125_));
  XOR2X1   g06869(.A(new_n7125_), .B(new_n6962_), .Y(new_n7126_));
  XOR2X1   g06870(.A(new_n7126_), .B(new_n6959_), .Y(new_n7127_));
  XOR2X1   g06871(.A(new_n7127_), .B(new_n6955_), .Y(new_n7128_));
  XOR2X1   g06872(.A(new_n7128_), .B(new_n6947_), .Y(new_n7129_));
  XOR2X1   g06873(.A(new_n7129_), .B(new_n6943_), .Y(\f[60] ));
  OR2X1    g06874(.A(new_n6917_), .B(new_n6913_), .Y(new_n7131_));
  OAI21X1  g06875(.A0(new_n6919_), .A1(new_n6756_), .B0(new_n7131_), .Y(new_n7132_));
  INVX1    g06876(.A(new_n6978_), .Y(new_n7133_));
  AND2X1   g06877(.A(new_n7122_), .B(new_n7133_), .Y(new_n7134_));
  XOR2X1   g06878(.A(new_n7122_), .B(new_n7133_), .Y(new_n7135_));
  AOI21X1  g06879(.A0(new_n7135_), .A1(new_n7132_), .B0(new_n7134_), .Y(new_n7136_));
  AOI22X1  g06880(.A0(new_n603_), .A1(\b[52] ), .B0(new_n602_), .B1(\b[51] ), .Y(new_n7137_));
  OAI21X1  g06881(.A0(new_n601_), .A1(new_n5234_), .B0(new_n7137_), .Y(new_n7138_));
  AOI21X1  g06882(.A0(new_n5590_), .A1(new_n518_), .B0(new_n7138_), .Y(new_n7139_));
  XOR2X1   g06883(.A(new_n7139_), .B(new_n515_), .Y(new_n7140_));
  INVX1    g06884(.A(new_n6986_), .Y(new_n7141_));
  AND2X1   g06885(.A(new_n7120_), .B(new_n7141_), .Y(new_n7142_));
  AOI21X1  g06886(.A0(new_n6981_), .A1(new_n6979_), .B0(new_n7121_), .Y(new_n7143_));
  OR2X1    g06887(.A(new_n7143_), .B(new_n7142_), .Y(new_n7144_));
  AOI22X1  g06888(.A0(new_n818_), .A1(\b[49] ), .B0(new_n817_), .B1(\b[48] ), .Y(new_n7145_));
  OAI21X1  g06889(.A0(new_n816_), .A1(new_n5039_), .B0(new_n7145_), .Y(new_n7146_));
  AOI21X1  g06890(.A0(new_n5038_), .A1(new_n668_), .B0(new_n7146_), .Y(new_n7147_));
  XOR2X1   g06891(.A(new_n7147_), .B(\a[14] ), .Y(new_n7148_));
  INVX1    g06892(.A(new_n7148_), .Y(new_n7149_));
  NAND2X1  g06893(.A(new_n7117_), .B(new_n6995_), .Y(new_n7150_));
  OR2X1    g06894(.A(new_n7119_), .B(new_n6990_), .Y(new_n7151_));
  AND2X1   g06895(.A(new_n7151_), .B(new_n7150_), .Y(new_n7152_));
  NOR2X1   g06896(.A(new_n7115_), .B(new_n7111_), .Y(new_n7153_));
  AOI21X1  g06897(.A0(new_n7116_), .A1(new_n6900_), .B0(new_n7153_), .Y(new_n7154_));
  INVX1    g06898(.A(new_n7087_), .Y(new_n7155_));
  NOR2X1   g06899(.A(new_n7091_), .B(new_n7155_), .Y(new_n7156_));
  INVX1    g06900(.A(new_n7092_), .Y(new_n7157_));
  AOI21X1  g06901(.A0(new_n7157_), .A1(new_n7001_), .B0(new_n7156_), .Y(new_n7158_));
  XOR2X1   g06902(.A(new_n7072_), .B(new_n7068_), .Y(new_n7159_));
  XOR2X1   g06903(.A(new_n7077_), .B(new_n7159_), .Y(new_n7160_));
  XOR2X1   g06904(.A(new_n7080_), .B(new_n7160_), .Y(new_n7161_));
  OR2X1    g06905(.A(new_n7085_), .B(new_n7161_), .Y(new_n7162_));
  OAI21X1  g06906(.A0(new_n7086_), .A1(new_n6868_), .B0(new_n7162_), .Y(new_n7163_));
  INVX1    g06907(.A(new_n7015_), .Y(new_n7164_));
  AND2X1   g06908(.A(new_n7059_), .B(new_n7164_), .Y(new_n7165_));
  INVX1    g06909(.A(new_n7165_), .Y(new_n7166_));
  OAI21X1  g06910(.A0(new_n7060_), .A1(new_n7011_), .B0(new_n7166_), .Y(new_n7167_));
  XOR2X1   g06911(.A(new_n7044_), .B(new_n6019_), .Y(new_n7168_));
  AND2X1   g06912(.A(new_n7168_), .B(new_n7041_), .Y(new_n7169_));
  NOR2X1   g06913(.A(new_n7046_), .B(new_n6818_), .Y(new_n7170_));
  NOR2X1   g06914(.A(new_n7170_), .B(new_n7169_), .Y(new_n7171_));
  INVX1    g06915(.A(new_n7171_), .Y(new_n7172_));
  AOI22X1  g06916(.A0(new_n6438_), .A1(\b[7] ), .B0(new_n6437_), .B1(\b[6] ), .Y(new_n7173_));
  OAI21X1  g06917(.A0(new_n6436_), .A1(new_n395_), .B0(new_n7173_), .Y(new_n7174_));
  AOI21X1  g06918(.A0(new_n6023_), .A1(new_n394_), .B0(new_n7174_), .Y(new_n7175_));
  XOR2X1   g06919(.A(new_n7175_), .B(new_n6019_), .Y(new_n7176_));
  OR4X1    g06920(.A(new_n7035_), .B(new_n6808_), .C(new_n6607_), .D(new_n6595_), .Y(new_n7177_));
  OAI21X1  g06921(.A0(new_n7040_), .A1(new_n7036_), .B0(new_n7177_), .Y(new_n7178_));
  AND2X1   g06922(.A(new_n6598_), .B(new_n323_), .Y(new_n7179_));
  NOR4X1   g06923(.A(new_n6599_), .B(new_n6597_), .C(new_n6602_), .D(new_n277_), .Y(new_n7180_));
  OAI22X1  g06924(.A0(new_n6604_), .A1(new_n325_), .B0(new_n6601_), .B1(new_n297_), .Y(new_n7181_));
  NOR3X1   g06925(.A(new_n7181_), .B(new_n7180_), .C(new_n7179_), .Y(new_n7182_));
  XOR2X1   g06926(.A(new_n7182_), .B(new_n6596_), .Y(new_n7183_));
  OAI21X1  g06927(.A0(new_n7033_), .A1(new_n274_), .B0(\a[62] ), .Y(new_n7184_));
  INVX1    g06928(.A(\a[62] ), .Y(new_n7185_));
  XOR2X1   g06929(.A(new_n7185_), .B(\a[61] ), .Y(new_n7186_));
  NOR2X1   g06930(.A(new_n7186_), .B(new_n7033_), .Y(new_n7187_));
  XOR2X1   g06931(.A(\a[61] ), .B(\a[60] ), .Y(new_n7188_));
  AND2X1   g06932(.A(new_n7188_), .B(new_n7033_), .Y(new_n7189_));
  INVX1    g06933(.A(new_n7189_), .Y(new_n7190_));
  INVX1    g06934(.A(new_n7033_), .Y(new_n7191_));
  AND2X1   g06935(.A(new_n7186_), .B(new_n7191_), .Y(new_n7192_));
  INVX1    g06936(.A(new_n7192_), .Y(new_n7193_));
  OAI22X1  g06937(.A0(new_n7193_), .A1(new_n275_), .B0(new_n7190_), .B1(new_n274_), .Y(new_n7194_));
  AOI21X1  g06938(.A0(new_n7187_), .A1(new_n263_), .B0(new_n7194_), .Y(new_n7195_));
  XOR2X1   g06939(.A(new_n7195_), .B(\a[62] ), .Y(new_n7196_));
  XOR2X1   g06940(.A(new_n7196_), .B(new_n7184_), .Y(new_n7197_));
  XOR2X1   g06941(.A(new_n7197_), .B(new_n7183_), .Y(new_n7198_));
  XOR2X1   g06942(.A(new_n7198_), .B(new_n7178_), .Y(new_n7199_));
  XOR2X1   g06943(.A(new_n7199_), .B(new_n7176_), .Y(new_n7200_));
  XOR2X1   g06944(.A(new_n7200_), .B(new_n7172_), .Y(new_n7201_));
  AOI22X1  g06945(.A0(new_n5430_), .A1(\b[10] ), .B0(new_n5427_), .B1(\b[9] ), .Y(new_n7202_));
  OAI21X1  g06946(.A0(new_n5891_), .A1(new_n489_), .B0(new_n7202_), .Y(new_n7203_));
  AOI21X1  g06947(.A0(new_n5425_), .A1(new_n543_), .B0(new_n7203_), .Y(new_n7204_));
  XOR2X1   g06948(.A(new_n7204_), .B(\a[53] ), .Y(new_n7205_));
  XOR2X1   g06949(.A(new_n7205_), .B(new_n7201_), .Y(new_n7206_));
  NOR2X1   g06950(.A(new_n7052_), .B(new_n7048_), .Y(new_n7207_));
  AOI21X1  g06951(.A0(new_n7053_), .A1(new_n7031_), .B0(new_n7207_), .Y(new_n7208_));
  XOR2X1   g06952(.A(new_n7208_), .B(new_n7206_), .Y(new_n7209_));
  INVX1    g06953(.A(new_n7209_), .Y(new_n7210_));
  AOI22X1  g06954(.A0(new_n4880_), .A1(\b[13] ), .B0(new_n4877_), .B1(\b[12] ), .Y(new_n7211_));
  OAI21X1  g06955(.A0(new_n5291_), .A1(new_n716_), .B0(new_n7211_), .Y(new_n7212_));
  AOI21X1  g06956(.A0(new_n4875_), .A1(new_n715_), .B0(new_n7212_), .Y(new_n7213_));
  XOR2X1   g06957(.A(new_n7213_), .B(\a[50] ), .Y(new_n7214_));
  AND2X1   g06958(.A(new_n7214_), .B(new_n7210_), .Y(new_n7215_));
  INVX1    g06959(.A(new_n7215_), .Y(new_n7216_));
  AND2X1   g06960(.A(new_n7054_), .B(new_n7029_), .Y(new_n7217_));
  INVX1    g06961(.A(new_n7217_), .Y(new_n7218_));
  OR2X1    g06962(.A(new_n7056_), .B(new_n7024_), .Y(new_n7219_));
  XOR2X1   g06963(.A(new_n7214_), .B(new_n7210_), .Y(new_n7220_));
  AOI21X1  g06964(.A0(new_n7219_), .A1(new_n7218_), .B0(new_n7220_), .Y(new_n7221_));
  AND2X1   g06965(.A(new_n7219_), .B(new_n7218_), .Y(new_n7222_));
  INVX1    g06966(.A(new_n7222_), .Y(new_n7223_));
  NOR2X1   g06967(.A(new_n7214_), .B(new_n7210_), .Y(new_n7224_));
  AOI21X1  g06968(.A0(new_n7216_), .A1(new_n7223_), .B0(new_n7224_), .Y(new_n7225_));
  AOI21X1  g06969(.A0(new_n7225_), .A1(new_n7216_), .B0(new_n7221_), .Y(new_n7226_));
  AOI22X1  g06970(.A0(new_n4572_), .A1(\b[16] ), .B0(new_n4571_), .B1(\b[15] ), .Y(new_n7227_));
  OAI21X1  g06971(.A0(new_n4740_), .A1(new_n792_), .B0(new_n7227_), .Y(new_n7228_));
  AOI21X1  g06972(.A0(new_n4375_), .A1(new_n842_), .B0(new_n7228_), .Y(new_n7229_));
  XOR2X1   g06973(.A(new_n7229_), .B(\a[47] ), .Y(new_n7230_));
  XOR2X1   g06974(.A(new_n7230_), .B(new_n7226_), .Y(new_n7231_));
  AND2X1   g06975(.A(new_n7057_), .B(new_n7022_), .Y(new_n7232_));
  AOI21X1  g06976(.A0(new_n7058_), .A1(new_n7018_), .B0(new_n7232_), .Y(new_n7233_));
  XOR2X1   g06977(.A(new_n7233_), .B(new_n7231_), .Y(new_n7234_));
  AOI22X1  g06978(.A0(new_n4095_), .A1(\b[19] ), .B0(new_n4094_), .B1(\b[18] ), .Y(new_n7235_));
  OAI21X1  g06979(.A0(new_n4233_), .A1(new_n1118_), .B0(new_n7235_), .Y(new_n7236_));
  AOI21X1  g06980(.A0(new_n3901_), .A1(new_n1117_), .B0(new_n7236_), .Y(new_n7237_));
  XOR2X1   g06981(.A(new_n7237_), .B(\a[44] ), .Y(new_n7238_));
  XOR2X1   g06982(.A(new_n7238_), .B(new_n7234_), .Y(new_n7239_));
  NAND2X1  g06983(.A(new_n7239_), .B(new_n7167_), .Y(new_n7240_));
  NOR2X1   g06984(.A(new_n7238_), .B(new_n7234_), .Y(new_n7241_));
  AND2X1   g06985(.A(new_n7238_), .B(new_n7234_), .Y(new_n7242_));
  NOR3X1   g06986(.A(new_n7242_), .B(new_n7241_), .C(new_n7167_), .Y(new_n7243_));
  AOI21X1  g06987(.A0(new_n7240_), .A1(new_n7167_), .B0(new_n7243_), .Y(new_n7244_));
  AOI22X1  g06988(.A0(new_n3652_), .A1(\b[22] ), .B0(new_n3651_), .B1(\b[21] ), .Y(new_n7245_));
  OAI21X1  g06989(.A0(new_n3778_), .A1(new_n1297_), .B0(new_n7245_), .Y(new_n7246_));
  AOI21X1  g06990(.A0(new_n3480_), .A1(new_n1399_), .B0(new_n7246_), .Y(new_n7247_));
  XOR2X1   g06991(.A(new_n7247_), .B(\a[41] ), .Y(new_n7248_));
  XOR2X1   g06992(.A(new_n7248_), .B(new_n7244_), .Y(new_n7249_));
  AND2X1   g06993(.A(new_n7061_), .B(new_n7007_), .Y(new_n7250_));
  AOI21X1  g06994(.A0(new_n7062_), .A1(new_n7003_), .B0(new_n7250_), .Y(new_n7251_));
  XOR2X1   g06995(.A(new_n7251_), .B(new_n7249_), .Y(new_n7252_));
  AOI22X1  g06996(.A0(new_n3204_), .A1(\b[25] ), .B0(new_n3203_), .B1(\b[24] ), .Y(new_n7253_));
  OAI21X1  g06997(.A0(new_n3321_), .A1(new_n1591_), .B0(new_n7253_), .Y(new_n7254_));
  AOI21X1  g06998(.A0(new_n3080_), .A1(new_n1590_), .B0(new_n7254_), .Y(new_n7255_));
  XOR2X1   g06999(.A(new_n7255_), .B(\a[38] ), .Y(new_n7256_));
  XOR2X1   g07000(.A(new_n7256_), .B(new_n7252_), .Y(new_n7257_));
  INVX1    g07001(.A(new_n7257_), .Y(new_n7258_));
  XOR2X1   g07002(.A(new_n7066_), .B(new_n3078_), .Y(new_n7259_));
  NAND2X1  g07003(.A(new_n7259_), .B(new_n7063_), .Y(new_n7260_));
  OAI21X1  g07004(.A0(new_n7072_), .A1(new_n7068_), .B0(new_n7260_), .Y(new_n7261_));
  XOR2X1   g07005(.A(new_n7261_), .B(new_n7258_), .Y(new_n7262_));
  AOI22X1  g07006(.A0(new_n2813_), .A1(\b[28] ), .B0(new_n2812_), .B1(\b[27] ), .Y(new_n7263_));
  OAI21X1  g07007(.A0(new_n2946_), .A1(new_n1877_), .B0(new_n7263_), .Y(new_n7264_));
  AOI21X1  g07008(.A0(new_n2652_), .A1(new_n2004_), .B0(new_n7264_), .Y(new_n7265_));
  XOR2X1   g07009(.A(new_n7265_), .B(\a[35] ), .Y(new_n7266_));
  XOR2X1   g07010(.A(new_n7266_), .B(new_n7262_), .Y(new_n7267_));
  NOR2X1   g07011(.A(new_n7077_), .B(new_n7073_), .Y(new_n7268_));
  AOI21X1  g07012(.A0(new_n7080_), .A1(new_n7078_), .B0(new_n7268_), .Y(new_n7269_));
  XOR2X1   g07013(.A(new_n7269_), .B(new_n7267_), .Y(new_n7270_));
  AOI22X1  g07014(.A0(new_n2545_), .A1(\b[31] ), .B0(new_n2544_), .B1(\b[30] ), .Y(new_n7271_));
  OAI21X1  g07015(.A0(new_n2543_), .A1(new_n2359_), .B0(new_n7271_), .Y(new_n7272_));
  AOI21X1  g07016(.A0(new_n2358_), .A1(new_n2260_), .B0(new_n7272_), .Y(new_n7273_));
  XOR2X1   g07017(.A(new_n7273_), .B(\a[32] ), .Y(new_n7274_));
  XOR2X1   g07018(.A(new_n7274_), .B(new_n7270_), .Y(new_n7275_));
  INVX1    g07019(.A(new_n7275_), .Y(new_n7276_));
  XOR2X1   g07020(.A(new_n7276_), .B(new_n7163_), .Y(new_n7277_));
  AOI22X1  g07021(.A0(new_n2163_), .A1(\b[34] ), .B0(new_n2162_), .B1(\b[33] ), .Y(new_n7278_));
  OAI21X1  g07022(.A0(new_n2161_), .A1(new_n2612_), .B0(new_n7278_), .Y(new_n7279_));
  AOI21X1  g07023(.A0(new_n2759_), .A1(new_n1907_), .B0(new_n7279_), .Y(new_n7280_));
  XOR2X1   g07024(.A(new_n7280_), .B(\a[29] ), .Y(new_n7281_));
  XOR2X1   g07025(.A(new_n7281_), .B(new_n7277_), .Y(new_n7282_));
  XOR2X1   g07026(.A(new_n7282_), .B(new_n7158_), .Y(new_n7283_));
  AOI22X1  g07027(.A0(new_n1814_), .A1(\b[37] ), .B0(new_n1813_), .B1(\b[36] ), .Y(new_n7284_));
  OAI21X1  g07028(.A0(new_n1812_), .A1(new_n3156_), .B0(new_n7284_), .Y(new_n7285_));
  AOI21X1  g07029(.A0(new_n3155_), .A1(new_n1617_), .B0(new_n7285_), .Y(new_n7286_));
  XOR2X1   g07030(.A(new_n7286_), .B(\a[26] ), .Y(new_n7287_));
  INVX1    g07031(.A(new_n7287_), .Y(new_n7288_));
  XOR2X1   g07032(.A(new_n7288_), .B(new_n7283_), .Y(new_n7289_));
  NOR2X1   g07033(.A(new_n7097_), .B(new_n7093_), .Y(new_n7290_));
  AOI21X1  g07034(.A0(new_n7098_), .A1(new_n6999_), .B0(new_n7290_), .Y(new_n7291_));
  XOR2X1   g07035(.A(new_n7291_), .B(new_n7289_), .Y(new_n7292_));
  AOI22X1  g07036(.A0(new_n1526_), .A1(\b[40] ), .B0(new_n1525_), .B1(\b[39] ), .Y(new_n7293_));
  OAI21X1  g07037(.A0(new_n1524_), .A1(new_n3575_), .B0(new_n7293_), .Y(new_n7294_));
  AOI21X1  g07038(.A0(new_n3574_), .A1(new_n1347_), .B0(new_n7294_), .Y(new_n7295_));
  XOR2X1   g07039(.A(new_n7295_), .B(\a[23] ), .Y(new_n7296_));
  XOR2X1   g07040(.A(new_n7296_), .B(new_n7292_), .Y(new_n7297_));
  NAND2X1  g07041(.A(new_n7104_), .B(new_n7099_), .Y(new_n7298_));
  XOR2X1   g07042(.A(new_n7103_), .B(new_n7099_), .Y(new_n7299_));
  OAI21X1  g07043(.A0(new_n7110_), .A1(new_n7299_), .B0(new_n7298_), .Y(new_n7300_));
  XOR2X1   g07044(.A(new_n7300_), .B(new_n7297_), .Y(new_n7301_));
  AOI22X1  g07045(.A0(new_n1263_), .A1(\b[43] ), .B0(new_n1262_), .B1(\b[42] ), .Y(new_n7302_));
  OAI21X1  g07046(.A0(new_n1261_), .A1(new_n4015_), .B0(new_n7302_), .Y(new_n7303_));
  AOI21X1  g07047(.A0(new_n4014_), .A1(new_n1075_), .B0(new_n7303_), .Y(new_n7304_));
  XOR2X1   g07048(.A(new_n7304_), .B(\a[20] ), .Y(new_n7305_));
  AND2X1   g07049(.A(new_n7305_), .B(new_n7301_), .Y(new_n7306_));
  XOR2X1   g07050(.A(new_n7305_), .B(new_n7301_), .Y(new_n7307_));
  OR2X1    g07051(.A(new_n7305_), .B(new_n7301_), .Y(new_n7308_));
  OAI21X1  g07052(.A0(new_n7306_), .A1(new_n7154_), .B0(new_n7308_), .Y(new_n7309_));
  OAI22X1  g07053(.A0(new_n7309_), .A1(new_n7306_), .B0(new_n7307_), .B1(new_n7154_), .Y(new_n7310_));
  AOI22X1  g07054(.A0(new_n1017_), .A1(\b[46] ), .B0(new_n1016_), .B1(\b[45] ), .Y(new_n7311_));
  OAI21X1  g07055(.A0(new_n1015_), .A1(new_n4336_), .B0(new_n7311_), .Y(new_n7312_));
  AOI21X1  g07056(.A0(new_n4509_), .A1(new_n882_), .B0(new_n7312_), .Y(new_n7313_));
  XOR2X1   g07057(.A(new_n7313_), .B(\a[17] ), .Y(new_n7314_));
  XOR2X1   g07058(.A(new_n7314_), .B(new_n7310_), .Y(new_n7315_));
  XOR2X1   g07059(.A(new_n7315_), .B(new_n7152_), .Y(new_n7316_));
  XOR2X1   g07060(.A(new_n7316_), .B(new_n7149_), .Y(new_n7317_));
  XOR2X1   g07061(.A(new_n7317_), .B(new_n7144_), .Y(new_n7318_));
  XOR2X1   g07062(.A(new_n7318_), .B(new_n7140_), .Y(new_n7319_));
  XOR2X1   g07063(.A(new_n7319_), .B(new_n7136_), .Y(new_n7320_));
  AOI22X1  g07064(.A0(new_n469_), .A1(\b[55] ), .B0(new_n468_), .B1(\b[54] ), .Y(new_n7321_));
  OAI21X1  g07065(.A0(new_n467_), .A1(new_n6151_), .B0(new_n7321_), .Y(new_n7322_));
  AOI21X1  g07066(.A0(new_n6150_), .A1(new_n404_), .B0(new_n7322_), .Y(new_n7323_));
  XOR2X1   g07067(.A(new_n7323_), .B(\a[8] ), .Y(new_n7324_));
  XOR2X1   g07068(.A(new_n7324_), .B(new_n7320_), .Y(new_n7325_));
  AND2X1   g07069(.A(new_n7124_), .B(new_n6966_), .Y(new_n7326_));
  AOI21X1  g07070(.A0(new_n7125_), .A1(new_n6962_), .B0(new_n7326_), .Y(new_n7327_));
  XOR2X1   g07071(.A(new_n7327_), .B(new_n7325_), .Y(new_n7328_));
  AOI22X1  g07072(.A0(new_n369_), .A1(\b[58] ), .B0(new_n368_), .B1(\b[57] ), .Y(new_n7329_));
  OAI21X1  g07073(.A0(new_n367_), .A1(new_n6520_), .B0(new_n7329_), .Y(new_n7330_));
  AOI21X1  g07074(.A0(new_n6732_), .A1(new_n308_), .B0(new_n7330_), .Y(new_n7331_));
  XOR2X1   g07075(.A(new_n7331_), .B(\a[5] ), .Y(new_n7332_));
  XOR2X1   g07076(.A(new_n7332_), .B(new_n7328_), .Y(new_n7333_));
  AND2X1   g07077(.A(\b[60] ), .B(\b[59] ), .Y(new_n7334_));
  AOI21X1  g07078(.A0(new_n6950_), .A1(new_n6949_), .B0(new_n7334_), .Y(new_n7335_));
  XOR2X1   g07079(.A(\b[61] ), .B(\b[60] ), .Y(new_n7336_));
  INVX1    g07080(.A(new_n7336_), .Y(new_n7337_));
  XOR2X1   g07081(.A(new_n7337_), .B(new_n7335_), .Y(new_n7338_));
  INVX1    g07082(.A(\b[59] ), .Y(new_n7339_));
  AOI22X1  g07083(.A0(new_n267_), .A1(\b[61] ), .B0(new_n266_), .B1(\b[60] ), .Y(new_n7340_));
  OAI21X1  g07084(.A0(new_n350_), .A1(new_n7339_), .B0(new_n7340_), .Y(new_n7341_));
  AOI21X1  g07085(.A0(new_n7338_), .A1(new_n318_), .B0(new_n7341_), .Y(new_n7342_));
  XOR2X1   g07086(.A(new_n7342_), .B(\a[2] ), .Y(new_n7343_));
  XOR2X1   g07087(.A(new_n7343_), .B(new_n7333_), .Y(new_n7344_));
  AND2X1   g07088(.A(new_n7126_), .B(new_n6959_), .Y(new_n7345_));
  AOI21X1  g07089(.A0(new_n7127_), .A1(new_n6955_), .B0(new_n7345_), .Y(new_n7346_));
  XOR2X1   g07090(.A(new_n7346_), .B(new_n7344_), .Y(new_n7347_));
  OAI21X1  g07091(.A0(new_n6937_), .A1(new_n6927_), .B0(new_n6945_), .Y(new_n7348_));
  AND2X1   g07092(.A(new_n7128_), .B(new_n7348_), .Y(new_n7349_));
  AOI21X1  g07093(.A0(new_n6942_), .A1(new_n6941_), .B0(new_n7129_), .Y(new_n7350_));
  OR2X1    g07094(.A(new_n7350_), .B(new_n7349_), .Y(new_n7351_));
  XOR2X1   g07095(.A(new_n7351_), .B(new_n7347_), .Y(\f[61] ));
  OR2X1    g07096(.A(new_n7346_), .B(new_n7344_), .Y(new_n7353_));
  OAI21X1  g07097(.A0(new_n7350_), .A1(new_n7349_), .B0(new_n7347_), .Y(new_n7354_));
  AND2X1   g07098(.A(new_n7354_), .B(new_n7353_), .Y(new_n7355_));
  OR2X1    g07099(.A(new_n7332_), .B(new_n7328_), .Y(new_n7356_));
  XOR2X1   g07100(.A(new_n7323_), .B(new_n400_), .Y(new_n7357_));
  XOR2X1   g07101(.A(new_n7357_), .B(new_n7320_), .Y(new_n7358_));
  XOR2X1   g07102(.A(new_n7327_), .B(new_n7358_), .Y(new_n7359_));
  XOR2X1   g07103(.A(new_n7332_), .B(new_n7359_), .Y(new_n7360_));
  OR2X1    g07104(.A(new_n7343_), .B(new_n7360_), .Y(new_n7361_));
  AND2X1   g07105(.A(new_n7361_), .B(new_n7356_), .Y(new_n7362_));
  NOR2X1   g07106(.A(new_n7318_), .B(new_n7140_), .Y(new_n7363_));
  NAND2X1  g07107(.A(new_n7318_), .B(new_n7140_), .Y(new_n7364_));
  OAI21X1  g07108(.A0(new_n7363_), .A1(new_n7136_), .B0(new_n7364_), .Y(new_n7365_));
  AND2X1   g07109(.A(new_n7316_), .B(new_n7149_), .Y(new_n7366_));
  AOI21X1  g07110(.A0(new_n7317_), .A1(new_n7144_), .B0(new_n7366_), .Y(new_n7367_));
  NAND2X1  g07111(.A(new_n7305_), .B(new_n7301_), .Y(new_n7368_));
  NOR2X1   g07112(.A(new_n7307_), .B(new_n7154_), .Y(new_n7369_));
  AND2X1   g07113(.A(new_n7116_), .B(new_n6900_), .Y(new_n7370_));
  OAI21X1  g07114(.A0(new_n7370_), .A1(new_n7153_), .B0(new_n7307_), .Y(new_n7371_));
  AND2X1   g07115(.A(new_n7371_), .B(new_n7308_), .Y(new_n7372_));
  AOI21X1  g07116(.A0(new_n7372_), .A1(new_n7368_), .B0(new_n7369_), .Y(new_n7373_));
  NOR2X1   g07117(.A(new_n7314_), .B(new_n7373_), .Y(new_n7374_));
  AOI21X1  g07118(.A0(new_n7151_), .A1(new_n7150_), .B0(new_n7315_), .Y(new_n7375_));
  NOR2X1   g07119(.A(new_n7375_), .B(new_n7374_), .Y(new_n7376_));
  XOR2X1   g07120(.A(new_n7287_), .B(new_n7283_), .Y(new_n7377_));
  XOR2X1   g07121(.A(new_n7291_), .B(new_n7377_), .Y(new_n7378_));
  NOR2X1   g07122(.A(new_n7296_), .B(new_n7378_), .Y(new_n7379_));
  XOR2X1   g07123(.A(new_n7296_), .B(new_n7378_), .Y(new_n7380_));
  AND2X1   g07124(.A(new_n7300_), .B(new_n7380_), .Y(new_n7381_));
  OR2X1    g07125(.A(new_n7381_), .B(new_n7379_), .Y(new_n7382_));
  OR2X1    g07126(.A(new_n7248_), .B(new_n7244_), .Y(new_n7383_));
  INVX1    g07127(.A(new_n7249_), .Y(new_n7384_));
  OAI21X1  g07128(.A0(new_n7251_), .A1(new_n7384_), .B0(new_n7383_), .Y(new_n7385_));
  AOI21X1  g07129(.A0(new_n7239_), .A1(new_n7167_), .B0(new_n7241_), .Y(new_n7386_));
  NOR2X1   g07130(.A(new_n7230_), .B(new_n7226_), .Y(new_n7387_));
  INVX1    g07131(.A(new_n7387_), .Y(new_n7388_));
  INVX1    g07132(.A(new_n7231_), .Y(new_n7389_));
  OAI21X1  g07133(.A0(new_n7233_), .A1(new_n7389_), .B0(new_n7388_), .Y(new_n7390_));
  AOI22X1  g07134(.A0(new_n4572_), .A1(\b[17] ), .B0(new_n4571_), .B1(\b[16] ), .Y(new_n7391_));
  OAI21X1  g07135(.A0(new_n4740_), .A1(new_n977_), .B0(new_n7391_), .Y(new_n7392_));
  AOI21X1  g07136(.A0(new_n4375_), .A1(new_n976_), .B0(new_n7392_), .Y(new_n7393_));
  XOR2X1   g07137(.A(new_n7393_), .B(\a[47] ), .Y(new_n7394_));
  XOR2X1   g07138(.A(new_n7204_), .B(new_n5423_), .Y(new_n7395_));
  NOR2X1   g07139(.A(new_n7208_), .B(new_n7206_), .Y(new_n7396_));
  AOI21X1  g07140(.A0(new_n7395_), .A1(new_n7201_), .B0(new_n7396_), .Y(new_n7397_));
  INVX1    g07141(.A(new_n7397_), .Y(new_n7398_));
  AOI22X1  g07142(.A0(new_n5430_), .A1(\b[11] ), .B0(new_n5427_), .B1(\b[10] ), .Y(new_n7399_));
  OAI21X1  g07143(.A0(new_n5891_), .A1(new_n590_), .B0(new_n7399_), .Y(new_n7400_));
  AOI21X1  g07144(.A0(new_n5425_), .A1(new_n589_), .B0(new_n7400_), .Y(new_n7401_));
  XOR2X1   g07145(.A(new_n7401_), .B(new_n5423_), .Y(new_n7402_));
  NAND2X1  g07146(.A(new_n7199_), .B(new_n7176_), .Y(new_n7403_));
  OAI21X1  g07147(.A0(new_n7170_), .A1(new_n7169_), .B0(new_n7200_), .Y(new_n7404_));
  NAND2X1  g07148(.A(new_n7404_), .B(new_n7403_), .Y(new_n7405_));
  AND2X1   g07149(.A(new_n7197_), .B(new_n7183_), .Y(new_n7406_));
  AND2X1   g07150(.A(new_n7198_), .B(new_n7178_), .Y(new_n7407_));
  OR2X1    g07151(.A(new_n7407_), .B(new_n7406_), .Y(new_n7408_));
  NOR2X1   g07152(.A(new_n7196_), .B(new_n7184_), .Y(new_n7409_));
  INVX1    g07153(.A(new_n7187_), .Y(new_n7410_));
  NOR3X1   g07154(.A(new_n7188_), .B(new_n7186_), .C(new_n7191_), .Y(new_n7411_));
  OAI22X1  g07155(.A0(new_n7193_), .A1(new_n277_), .B0(new_n7190_), .B1(new_n275_), .Y(new_n7412_));
  AOI21X1  g07156(.A0(new_n7411_), .A1(\b[0] ), .B0(new_n7412_), .Y(new_n7413_));
  OAI21X1  g07157(.A0(new_n7410_), .A1(new_n281_), .B0(new_n7413_), .Y(new_n7414_));
  XOR2X1   g07158(.A(new_n7414_), .B(new_n7185_), .Y(new_n7415_));
  XOR2X1   g07159(.A(new_n7415_), .B(new_n7409_), .Y(new_n7416_));
  AOI22X1  g07160(.A0(new_n6603_), .A1(\b[5] ), .B0(new_n6600_), .B1(\b[4] ), .Y(new_n7417_));
  OAI21X1  g07161(.A0(new_n6804_), .A1(new_n297_), .B0(new_n7417_), .Y(new_n7418_));
  AOI21X1  g07162(.A0(new_n6598_), .A1(new_n349_), .B0(new_n7418_), .Y(new_n7419_));
  XOR2X1   g07163(.A(new_n7419_), .B(\a[59] ), .Y(new_n7420_));
  NAND2X1  g07164(.A(new_n7420_), .B(new_n7416_), .Y(new_n7421_));
  XOR2X1   g07165(.A(new_n7420_), .B(new_n7416_), .Y(new_n7422_));
  INVX1    g07166(.A(new_n7422_), .Y(new_n7423_));
  NOR2X1   g07167(.A(new_n7420_), .B(new_n7416_), .Y(new_n7424_));
  AOI21X1  g07168(.A0(new_n7421_), .A1(new_n7408_), .B0(new_n7424_), .Y(new_n7425_));
  AOI22X1  g07169(.A0(new_n7425_), .A1(new_n7421_), .B0(new_n7423_), .B1(new_n7408_), .Y(new_n7426_));
  AOI22X1  g07170(.A0(new_n6438_), .A1(\b[8] ), .B0(new_n6437_), .B1(\b[7] ), .Y(new_n7427_));
  OAI21X1  g07171(.A0(new_n6436_), .A1(new_n392_), .B0(new_n7427_), .Y(new_n7428_));
  AOI21X1  g07172(.A0(new_n6023_), .A1(new_n454_), .B0(new_n7428_), .Y(new_n7429_));
  XOR2X1   g07173(.A(new_n7429_), .B(\a[56] ), .Y(new_n7430_));
  XOR2X1   g07174(.A(new_n7430_), .B(new_n7426_), .Y(new_n7431_));
  XOR2X1   g07175(.A(new_n7431_), .B(new_n7405_), .Y(new_n7432_));
  XOR2X1   g07176(.A(new_n7432_), .B(new_n7402_), .Y(new_n7433_));
  XOR2X1   g07177(.A(new_n7433_), .B(new_n7398_), .Y(new_n7434_));
  AOI22X1  g07178(.A0(new_n4880_), .A1(\b[14] ), .B0(new_n4877_), .B1(\b[13] ), .Y(new_n7435_));
  OAI21X1  g07179(.A0(new_n5291_), .A1(new_n713_), .B0(new_n7435_), .Y(new_n7436_));
  AOI21X1  g07180(.A0(new_n4875_), .A1(new_n734_), .B0(new_n7436_), .Y(new_n7437_));
  XOR2X1   g07181(.A(new_n7437_), .B(\a[50] ), .Y(new_n7438_));
  XOR2X1   g07182(.A(new_n7438_), .B(new_n7434_), .Y(new_n7439_));
  XOR2X1   g07183(.A(new_n7439_), .B(new_n7225_), .Y(new_n7440_));
  XOR2X1   g07184(.A(new_n7440_), .B(new_n7394_), .Y(new_n7441_));
  XOR2X1   g07185(.A(new_n7441_), .B(new_n7390_), .Y(new_n7442_));
  AOI22X1  g07186(.A0(new_n4095_), .A1(\b[20] ), .B0(new_n4094_), .B1(\b[19] ), .Y(new_n7443_));
  OAI21X1  g07187(.A0(new_n4233_), .A1(new_n1115_), .B0(new_n7443_), .Y(new_n7444_));
  AOI21X1  g07188(.A0(new_n3901_), .A1(new_n1217_), .B0(new_n7444_), .Y(new_n7445_));
  XOR2X1   g07189(.A(new_n7445_), .B(\a[44] ), .Y(new_n7446_));
  XOR2X1   g07190(.A(new_n7446_), .B(new_n7442_), .Y(new_n7447_));
  XOR2X1   g07191(.A(new_n7447_), .B(new_n7386_), .Y(new_n7448_));
  AOI22X1  g07192(.A0(new_n3652_), .A1(\b[23] ), .B0(new_n3651_), .B1(\b[22] ), .Y(new_n7449_));
  OAI21X1  g07193(.A0(new_n3778_), .A1(new_n1482_), .B0(new_n7449_), .Y(new_n7450_));
  AOI21X1  g07194(.A0(new_n3480_), .A1(new_n1481_), .B0(new_n7450_), .Y(new_n7451_));
  XOR2X1   g07195(.A(new_n7451_), .B(\a[41] ), .Y(new_n7452_));
  XOR2X1   g07196(.A(new_n7452_), .B(new_n7448_), .Y(new_n7453_));
  XOR2X1   g07197(.A(new_n7453_), .B(new_n7385_), .Y(new_n7454_));
  AOI22X1  g07198(.A0(new_n3204_), .A1(\b[26] ), .B0(new_n3203_), .B1(\b[25] ), .Y(new_n7455_));
  OAI21X1  g07199(.A0(new_n3321_), .A1(new_n1588_), .B0(new_n7455_), .Y(new_n7456_));
  AOI21X1  g07200(.A0(new_n3080_), .A1(new_n1783_), .B0(new_n7456_), .Y(new_n7457_));
  XOR2X1   g07201(.A(new_n7457_), .B(\a[38] ), .Y(new_n7458_));
  XOR2X1   g07202(.A(new_n7458_), .B(new_n7454_), .Y(new_n7459_));
  NOR2X1   g07203(.A(new_n7256_), .B(new_n7252_), .Y(new_n7460_));
  AOI21X1  g07204(.A0(new_n7261_), .A1(new_n7257_), .B0(new_n7460_), .Y(new_n7461_));
  XOR2X1   g07205(.A(new_n7461_), .B(new_n7459_), .Y(new_n7462_));
  AOI22X1  g07206(.A0(new_n2813_), .A1(\b[29] ), .B0(new_n2812_), .B1(\b[28] ), .Y(new_n7463_));
  OAI21X1  g07207(.A0(new_n2946_), .A1(new_n2126_), .B0(new_n7463_), .Y(new_n7464_));
  AOI21X1  g07208(.A0(new_n2652_), .A1(new_n2125_), .B0(new_n7464_), .Y(new_n7465_));
  XOR2X1   g07209(.A(new_n7465_), .B(\a[35] ), .Y(new_n7466_));
  INVX1    g07210(.A(new_n7466_), .Y(new_n7467_));
  XOR2X1   g07211(.A(new_n7467_), .B(new_n7462_), .Y(new_n7468_));
  INVX1    g07212(.A(new_n7468_), .Y(new_n7469_));
  OR2X1    g07213(.A(new_n7266_), .B(new_n7262_), .Y(new_n7470_));
  INVX1    g07214(.A(new_n7267_), .Y(new_n7471_));
  OAI21X1  g07215(.A0(new_n7269_), .A1(new_n7471_), .B0(new_n7470_), .Y(new_n7472_));
  XOR2X1   g07216(.A(new_n7472_), .B(new_n7469_), .Y(new_n7473_));
  AOI22X1  g07217(.A0(new_n2545_), .A1(\b[32] ), .B0(new_n2544_), .B1(\b[31] ), .Y(new_n7474_));
  OAI21X1  g07218(.A0(new_n2543_), .A1(new_n2356_), .B0(new_n7474_), .Y(new_n7475_));
  AOI21X1  g07219(.A0(new_n2495_), .A1(new_n2260_), .B0(new_n7475_), .Y(new_n7476_));
  XOR2X1   g07220(.A(new_n7476_), .B(\a[32] ), .Y(new_n7477_));
  NAND2X1  g07221(.A(new_n7477_), .B(new_n7473_), .Y(new_n7478_));
  NOR2X1   g07222(.A(new_n7274_), .B(new_n7270_), .Y(new_n7479_));
  AOI21X1  g07223(.A0(new_n7275_), .A1(new_n7163_), .B0(new_n7479_), .Y(new_n7480_));
  XOR2X1   g07224(.A(new_n7477_), .B(new_n7473_), .Y(new_n7481_));
  NOR2X1   g07225(.A(new_n7481_), .B(new_n7480_), .Y(new_n7482_));
  INVX1    g07226(.A(new_n7480_), .Y(new_n7483_));
  NOR2X1   g07227(.A(new_n7477_), .B(new_n7473_), .Y(new_n7484_));
  AOI21X1  g07228(.A0(new_n7478_), .A1(new_n7483_), .B0(new_n7484_), .Y(new_n7485_));
  AOI21X1  g07229(.A0(new_n7485_), .A1(new_n7478_), .B0(new_n7482_), .Y(new_n7486_));
  AOI22X1  g07230(.A0(new_n2163_), .A1(\b[35] ), .B0(new_n2162_), .B1(\b[34] ), .Y(new_n7487_));
  OAI21X1  g07231(.A0(new_n2161_), .A1(new_n2893_), .B0(new_n7487_), .Y(new_n7488_));
  AOI21X1  g07232(.A0(new_n2892_), .A1(new_n1907_), .B0(new_n7488_), .Y(new_n7489_));
  XOR2X1   g07233(.A(new_n7489_), .B(\a[29] ), .Y(new_n7490_));
  XOR2X1   g07234(.A(new_n7490_), .B(new_n7486_), .Y(new_n7491_));
  OR2X1    g07235(.A(new_n7281_), .B(new_n7277_), .Y(new_n7492_));
  AND2X1   g07236(.A(new_n7157_), .B(new_n7001_), .Y(new_n7493_));
  OAI21X1  g07237(.A0(new_n7493_), .A1(new_n7156_), .B0(new_n7282_), .Y(new_n7494_));
  AND2X1   g07238(.A(new_n7494_), .B(new_n7492_), .Y(new_n7495_));
  XOR2X1   g07239(.A(new_n7495_), .B(new_n7491_), .Y(new_n7496_));
  AOI22X1  g07240(.A0(new_n1814_), .A1(\b[38] ), .B0(new_n1813_), .B1(\b[37] ), .Y(new_n7497_));
  OAI21X1  g07241(.A0(new_n1812_), .A1(new_n3276_), .B0(new_n7497_), .Y(new_n7498_));
  AOI21X1  g07242(.A0(new_n3275_), .A1(new_n1617_), .B0(new_n7498_), .Y(new_n7499_));
  XOR2X1   g07243(.A(new_n7499_), .B(\a[26] ), .Y(new_n7500_));
  XOR2X1   g07244(.A(new_n7500_), .B(new_n7496_), .Y(new_n7501_));
  OR2X1    g07245(.A(new_n7287_), .B(new_n7283_), .Y(new_n7502_));
  OR2X1    g07246(.A(new_n7291_), .B(new_n7289_), .Y(new_n7503_));
  AND2X1   g07247(.A(new_n7503_), .B(new_n7502_), .Y(new_n7504_));
  XOR2X1   g07248(.A(new_n7504_), .B(new_n7501_), .Y(new_n7505_));
  AOI22X1  g07249(.A0(new_n1526_), .A1(\b[41] ), .B0(new_n1525_), .B1(\b[40] ), .Y(new_n7506_));
  OAI21X1  g07250(.A0(new_n1524_), .A1(new_n3723_), .B0(new_n7506_), .Y(new_n7507_));
  AOI21X1  g07251(.A0(new_n3722_), .A1(new_n1347_), .B0(new_n7507_), .Y(new_n7508_));
  XOR2X1   g07252(.A(new_n7508_), .B(\a[23] ), .Y(new_n7509_));
  NAND2X1  g07253(.A(new_n7509_), .B(new_n7505_), .Y(new_n7510_));
  OR2X1    g07254(.A(new_n7509_), .B(new_n7505_), .Y(new_n7511_));
  NAND3X1  g07255(.A(new_n7510_), .B(new_n7511_), .C(new_n7382_), .Y(new_n7512_));
  NOR2X1   g07256(.A(new_n7509_), .B(new_n7505_), .Y(new_n7513_));
  AOI21X1  g07257(.A0(new_n7510_), .A1(new_n7382_), .B0(new_n7513_), .Y(new_n7514_));
  AOI22X1  g07258(.A0(new_n7514_), .A1(new_n7510_), .B0(new_n7512_), .B1(new_n7382_), .Y(new_n7515_));
  AOI22X1  g07259(.A0(new_n1263_), .A1(\b[44] ), .B0(new_n1262_), .B1(\b[43] ), .Y(new_n7516_));
  OAI21X1  g07260(.A0(new_n1261_), .A1(new_n4012_), .B0(new_n7516_), .Y(new_n7517_));
  AOI21X1  g07261(.A0(new_n4178_), .A1(new_n1075_), .B0(new_n7517_), .Y(new_n7518_));
  XOR2X1   g07262(.A(new_n7518_), .B(\a[20] ), .Y(new_n7519_));
  INVX1    g07263(.A(new_n7519_), .Y(new_n7520_));
  XOR2X1   g07264(.A(new_n7520_), .B(new_n7515_), .Y(new_n7521_));
  XOR2X1   g07265(.A(new_n7521_), .B(new_n7309_), .Y(new_n7522_));
  AOI22X1  g07266(.A0(new_n1017_), .A1(\b[47] ), .B0(new_n1016_), .B1(\b[46] ), .Y(new_n7523_));
  OAI21X1  g07267(.A0(new_n1015_), .A1(new_n4674_), .B0(new_n7523_), .Y(new_n7524_));
  AOI21X1  g07268(.A0(new_n4673_), .A1(new_n882_), .B0(new_n7524_), .Y(new_n7525_));
  XOR2X1   g07269(.A(new_n7525_), .B(\a[17] ), .Y(new_n7526_));
  XOR2X1   g07270(.A(new_n7526_), .B(new_n7522_), .Y(new_n7527_));
  XOR2X1   g07271(.A(new_n7527_), .B(new_n7376_), .Y(new_n7528_));
  AOI22X1  g07272(.A0(new_n818_), .A1(\b[50] ), .B0(new_n817_), .B1(\b[49] ), .Y(new_n7529_));
  OAI21X1  g07273(.A0(new_n816_), .A1(new_n5036_), .B0(new_n7529_), .Y(new_n7530_));
  AOI21X1  g07274(.A0(new_n5204_), .A1(new_n668_), .B0(new_n7530_), .Y(new_n7531_));
  XOR2X1   g07275(.A(new_n7531_), .B(\a[14] ), .Y(new_n7532_));
  XOR2X1   g07276(.A(new_n7532_), .B(new_n7528_), .Y(new_n7533_));
  XOR2X1   g07277(.A(new_n7533_), .B(new_n7367_), .Y(new_n7534_));
  AOI22X1  g07278(.A0(new_n603_), .A1(\b[53] ), .B0(new_n602_), .B1(\b[52] ), .Y(new_n7535_));
  OAI21X1  g07279(.A0(new_n601_), .A1(new_n5787_), .B0(new_n7535_), .Y(new_n7536_));
  AOI21X1  g07280(.A0(new_n5786_), .A1(new_n518_), .B0(new_n7536_), .Y(new_n7537_));
  XOR2X1   g07281(.A(new_n7537_), .B(\a[11] ), .Y(new_n7538_));
  XOR2X1   g07282(.A(new_n7538_), .B(new_n7534_), .Y(new_n7539_));
  XOR2X1   g07283(.A(new_n7539_), .B(new_n7365_), .Y(new_n7540_));
  AOI22X1  g07284(.A0(new_n469_), .A1(\b[56] ), .B0(new_n468_), .B1(\b[55] ), .Y(new_n7541_));
  OAI21X1  g07285(.A0(new_n467_), .A1(new_n6148_), .B0(new_n7541_), .Y(new_n7542_));
  AOI21X1  g07286(.A0(new_n6342_), .A1(new_n404_), .B0(new_n7542_), .Y(new_n7543_));
  XOR2X1   g07287(.A(new_n7543_), .B(\a[8] ), .Y(new_n7544_));
  XOR2X1   g07288(.A(new_n7544_), .B(new_n7540_), .Y(new_n7545_));
  AOI22X1  g07289(.A0(new_n369_), .A1(\b[59] ), .B0(new_n368_), .B1(\b[58] ), .Y(new_n7546_));
  OAI21X1  g07290(.A0(new_n367_), .A1(new_n6933_), .B0(new_n7546_), .Y(new_n7547_));
  AOI21X1  g07291(.A0(new_n6932_), .A1(new_n308_), .B0(new_n7547_), .Y(new_n7548_));
  XOR2X1   g07292(.A(new_n7548_), .B(\a[5] ), .Y(new_n7549_));
  XOR2X1   g07293(.A(new_n7549_), .B(new_n7545_), .Y(new_n7550_));
  OR2X1    g07294(.A(new_n7324_), .B(new_n7320_), .Y(new_n7551_));
  OR2X1    g07295(.A(new_n7327_), .B(new_n7358_), .Y(new_n7552_));
  AND2X1   g07296(.A(new_n7552_), .B(new_n7551_), .Y(new_n7553_));
  XOR2X1   g07297(.A(new_n7553_), .B(new_n7550_), .Y(new_n7554_));
  NAND2X1  g07298(.A(\b[61] ), .B(\b[60] ), .Y(new_n7555_));
  OAI21X1  g07299(.A0(new_n7337_), .A1(new_n7335_), .B0(new_n7555_), .Y(new_n7556_));
  XOR2X1   g07300(.A(\b[62] ), .B(\b[61] ), .Y(new_n7557_));
  XOR2X1   g07301(.A(new_n7557_), .B(new_n7556_), .Y(new_n7558_));
  INVX1    g07302(.A(\b[60] ), .Y(new_n7559_));
  AOI22X1  g07303(.A0(new_n267_), .A1(\b[62] ), .B0(new_n266_), .B1(\b[61] ), .Y(new_n7560_));
  OAI21X1  g07304(.A0(new_n350_), .A1(new_n7559_), .B0(new_n7560_), .Y(new_n7561_));
  AOI21X1  g07305(.A0(new_n7558_), .A1(new_n318_), .B0(new_n7561_), .Y(new_n7562_));
  XOR2X1   g07306(.A(new_n7562_), .B(\a[2] ), .Y(new_n7563_));
  XOR2X1   g07307(.A(new_n7563_), .B(new_n7554_), .Y(new_n7564_));
  XOR2X1   g07308(.A(new_n7564_), .B(new_n7362_), .Y(new_n7565_));
  XOR2X1   g07309(.A(new_n7565_), .B(new_n7355_), .Y(\f[62] ));
  NOR2X1   g07310(.A(new_n7143_), .B(new_n7142_), .Y(new_n7567_));
  NAND2X1  g07311(.A(new_n7316_), .B(new_n7149_), .Y(new_n7568_));
  XOR2X1   g07312(.A(new_n7316_), .B(new_n7148_), .Y(new_n7569_));
  OAI21X1  g07313(.A0(new_n7569_), .A1(new_n7567_), .B0(new_n7568_), .Y(new_n7570_));
  NOR2X1   g07314(.A(new_n7532_), .B(new_n7528_), .Y(new_n7571_));
  AOI21X1  g07315(.A0(new_n7533_), .A1(new_n7570_), .B0(new_n7571_), .Y(new_n7572_));
  AOI22X1  g07316(.A0(new_n818_), .A1(\b[51] ), .B0(new_n817_), .B1(\b[50] ), .Y(new_n7573_));
  OAI21X1  g07317(.A0(new_n816_), .A1(new_n5237_), .B0(new_n7573_), .Y(new_n7574_));
  AOI21X1  g07318(.A0(new_n5236_), .A1(new_n668_), .B0(new_n7574_), .Y(new_n7575_));
  XOR2X1   g07319(.A(new_n7575_), .B(\a[14] ), .Y(new_n7576_));
  INVX1    g07320(.A(new_n7576_), .Y(new_n7577_));
  OR2X1    g07321(.A(new_n7375_), .B(new_n7374_), .Y(new_n7578_));
  NOR2X1   g07322(.A(new_n7526_), .B(new_n7522_), .Y(new_n7579_));
  AOI21X1  g07323(.A0(new_n7527_), .A1(new_n7578_), .B0(new_n7579_), .Y(new_n7580_));
  AOI22X1  g07324(.A0(new_n1017_), .A1(\b[48] ), .B0(new_n1016_), .B1(\b[47] ), .Y(new_n7581_));
  OAI21X1  g07325(.A0(new_n1015_), .A1(new_n4693_), .B0(new_n7581_), .Y(new_n7582_));
  AOI21X1  g07326(.A0(new_n4692_), .A1(new_n882_), .B0(new_n7582_), .Y(new_n7583_));
  XOR2X1   g07327(.A(new_n7583_), .B(\a[17] ), .Y(new_n7584_));
  OR2X1    g07328(.A(new_n7519_), .B(new_n7515_), .Y(new_n7585_));
  OAI21X1  g07329(.A0(new_n7521_), .A1(new_n7372_), .B0(new_n7585_), .Y(new_n7586_));
  AOI22X1  g07330(.A0(new_n1263_), .A1(\b[45] ), .B0(new_n1262_), .B1(\b[44] ), .Y(new_n7587_));
  OAI21X1  g07331(.A0(new_n1261_), .A1(new_n4339_), .B0(new_n7587_), .Y(new_n7588_));
  AOI21X1  g07332(.A0(new_n4338_), .A1(new_n1075_), .B0(new_n7588_), .Y(new_n7589_));
  XOR2X1   g07333(.A(new_n7589_), .B(\a[20] ), .Y(new_n7590_));
  INVX1    g07334(.A(new_n7590_), .Y(new_n7591_));
  AOI22X1  g07335(.A0(new_n1526_), .A1(\b[42] ), .B0(new_n1525_), .B1(\b[41] ), .Y(new_n7592_));
  OAI21X1  g07336(.A0(new_n1524_), .A1(new_n3720_), .B0(new_n7592_), .Y(new_n7593_));
  AOI21X1  g07337(.A0(new_n3860_), .A1(new_n1347_), .B0(new_n7593_), .Y(new_n7594_));
  XOR2X1   g07338(.A(new_n7594_), .B(\a[23] ), .Y(new_n7595_));
  NOR2X1   g07339(.A(new_n7500_), .B(new_n7496_), .Y(new_n7596_));
  OAI21X1  g07340(.A0(new_n7291_), .A1(new_n7289_), .B0(new_n7502_), .Y(new_n7597_));
  AOI21X1  g07341(.A0(new_n7597_), .A1(new_n7501_), .B0(new_n7596_), .Y(new_n7598_));
  OR2X1    g07342(.A(new_n7490_), .B(new_n7486_), .Y(new_n7599_));
  AND2X1   g07343(.A(new_n7477_), .B(new_n7473_), .Y(new_n7600_));
  OR2X1    g07344(.A(new_n7477_), .B(new_n7473_), .Y(new_n7601_));
  OAI21X1  g07345(.A0(new_n7600_), .A1(new_n7480_), .B0(new_n7601_), .Y(new_n7602_));
  OAI22X1  g07346(.A0(new_n7602_), .A1(new_n7600_), .B0(new_n7481_), .B1(new_n7480_), .Y(new_n7603_));
  XOR2X1   g07347(.A(new_n7490_), .B(new_n7603_), .Y(new_n7604_));
  OAI21X1  g07348(.A0(new_n7495_), .A1(new_n7604_), .B0(new_n7599_), .Y(new_n7605_));
  AND2X1   g07349(.A(new_n7239_), .B(new_n7167_), .Y(new_n7606_));
  OAI21X1  g07350(.A0(new_n7606_), .A1(new_n7241_), .B0(new_n7447_), .Y(new_n7607_));
  OAI21X1  g07351(.A0(new_n7446_), .A1(new_n7442_), .B0(new_n7607_), .Y(new_n7608_));
  AOI22X1  g07352(.A0(new_n4095_), .A1(\b[21] ), .B0(new_n4094_), .B1(\b[20] ), .Y(new_n7609_));
  OAI21X1  g07353(.A0(new_n4233_), .A1(new_n1300_), .B0(new_n7609_), .Y(new_n7610_));
  AOI21X1  g07354(.A0(new_n3901_), .A1(new_n1299_), .B0(new_n7610_), .Y(new_n7611_));
  XOR2X1   g07355(.A(new_n7611_), .B(new_n3899_), .Y(new_n7612_));
  INVX1    g07356(.A(new_n7390_), .Y(new_n7613_));
  INVX1    g07357(.A(new_n7394_), .Y(new_n7614_));
  NAND2X1  g07358(.A(new_n7440_), .B(new_n7614_), .Y(new_n7615_));
  OAI21X1  g07359(.A0(new_n7441_), .A1(new_n7613_), .B0(new_n7615_), .Y(new_n7616_));
  AND2X1   g07360(.A(new_n7432_), .B(new_n7402_), .Y(new_n7617_));
  AOI21X1  g07361(.A0(new_n7433_), .A1(new_n7398_), .B0(new_n7617_), .Y(new_n7618_));
  INVX1    g07362(.A(new_n7618_), .Y(new_n7619_));
  NAND2X1  g07363(.A(new_n7431_), .B(new_n7405_), .Y(new_n7620_));
  OAI21X1  g07364(.A0(new_n7430_), .A1(new_n7426_), .B0(new_n7620_), .Y(new_n7621_));
  INVX1    g07365(.A(new_n7425_), .Y(new_n7622_));
  NOR4X1   g07366(.A(new_n7414_), .B(new_n7196_), .C(new_n7034_), .D(new_n7185_), .Y(new_n7623_));
  XOR2X1   g07367(.A(\a[63] ), .B(new_n7185_), .Y(new_n7624_));
  NOR2X1   g07368(.A(new_n7624_), .B(new_n274_), .Y(new_n7625_));
  XOR2X1   g07369(.A(new_n7625_), .B(new_n7623_), .Y(new_n7626_));
  INVX1    g07370(.A(new_n7411_), .Y(new_n7627_));
  AOI22X1  g07371(.A0(new_n7192_), .A1(\b[3] ), .B0(new_n7189_), .B1(\b[2] ), .Y(new_n7628_));
  OAI21X1  g07372(.A0(new_n7627_), .A1(new_n275_), .B0(new_n7628_), .Y(new_n7629_));
  AOI21X1  g07373(.A0(new_n7187_), .A1(new_n366_), .B0(new_n7629_), .Y(new_n7630_));
  XOR2X1   g07374(.A(new_n7630_), .B(\a[62] ), .Y(new_n7631_));
  XOR2X1   g07375(.A(new_n7631_), .B(new_n7626_), .Y(new_n7632_));
  AOI22X1  g07376(.A0(new_n6603_), .A1(\b[6] ), .B0(new_n6600_), .B1(\b[5] ), .Y(new_n7633_));
  OAI21X1  g07377(.A0(new_n6804_), .A1(new_n325_), .B0(new_n7633_), .Y(new_n7634_));
  AOI21X1  g07378(.A0(new_n6598_), .A1(new_n378_), .B0(new_n7634_), .Y(new_n7635_));
  XOR2X1   g07379(.A(new_n7635_), .B(\a[59] ), .Y(new_n7636_));
  XOR2X1   g07380(.A(new_n7636_), .B(new_n7632_), .Y(new_n7637_));
  XOR2X1   g07381(.A(new_n7637_), .B(new_n7622_), .Y(new_n7638_));
  AOI22X1  g07382(.A0(new_n6438_), .A1(\b[9] ), .B0(new_n6437_), .B1(\b[8] ), .Y(new_n7639_));
  OAI21X1  g07383(.A0(new_n6436_), .A1(new_n492_), .B0(new_n7639_), .Y(new_n7640_));
  AOI21X1  g07384(.A0(new_n6023_), .A1(new_n491_), .B0(new_n7640_), .Y(new_n7641_));
  XOR2X1   g07385(.A(new_n7641_), .B(\a[56] ), .Y(new_n7642_));
  XOR2X1   g07386(.A(new_n7642_), .B(new_n7638_), .Y(new_n7643_));
  XOR2X1   g07387(.A(new_n7643_), .B(new_n7621_), .Y(new_n7644_));
  AOI22X1  g07388(.A0(new_n5430_), .A1(\b[12] ), .B0(new_n5427_), .B1(\b[11] ), .Y(new_n7645_));
  OAI21X1  g07389(.A0(new_n5891_), .A1(new_n587_), .B0(new_n7645_), .Y(new_n7646_));
  AOI21X1  g07390(.A0(new_n5425_), .A1(new_n635_), .B0(new_n7646_), .Y(new_n7647_));
  XOR2X1   g07391(.A(new_n7647_), .B(\a[53] ), .Y(new_n7648_));
  XOR2X1   g07392(.A(new_n7648_), .B(new_n7644_), .Y(new_n7649_));
  XOR2X1   g07393(.A(new_n7649_), .B(new_n7619_), .Y(new_n7650_));
  AOI22X1  g07394(.A0(new_n4880_), .A1(\b[15] ), .B0(new_n4877_), .B1(\b[14] ), .Y(new_n7651_));
  OAI21X1  g07395(.A0(new_n5291_), .A1(new_n795_), .B0(new_n7651_), .Y(new_n7652_));
  AOI21X1  g07396(.A0(new_n4875_), .A1(new_n794_), .B0(new_n7652_), .Y(new_n7653_));
  XOR2X1   g07397(.A(new_n7653_), .B(\a[50] ), .Y(new_n7654_));
  XOR2X1   g07398(.A(new_n7654_), .B(new_n7650_), .Y(new_n7655_));
  INVX1    g07399(.A(new_n7655_), .Y(new_n7656_));
  INVX1    g07400(.A(new_n7438_), .Y(new_n7657_));
  NOR2X1   g07401(.A(new_n7439_), .B(new_n7225_), .Y(new_n7658_));
  AOI21X1  g07402(.A0(new_n7657_), .A1(new_n7434_), .B0(new_n7658_), .Y(new_n7659_));
  XOR2X1   g07403(.A(new_n7659_), .B(new_n7656_), .Y(new_n7660_));
  AOI22X1  g07404(.A0(new_n4572_), .A1(\b[18] ), .B0(new_n4571_), .B1(\b[17] ), .Y(new_n7661_));
  OAI21X1  g07405(.A0(new_n4740_), .A1(new_n974_), .B0(new_n7661_), .Y(new_n7662_));
  AOI21X1  g07406(.A0(new_n4375_), .A1(new_n1042_), .B0(new_n7662_), .Y(new_n7663_));
  XOR2X1   g07407(.A(new_n7663_), .B(\a[47] ), .Y(new_n7664_));
  XOR2X1   g07408(.A(new_n7664_), .B(new_n7660_), .Y(new_n7665_));
  XOR2X1   g07409(.A(new_n7665_), .B(new_n7616_), .Y(new_n7666_));
  XOR2X1   g07410(.A(new_n7666_), .B(new_n7612_), .Y(new_n7667_));
  XOR2X1   g07411(.A(new_n7667_), .B(new_n7608_), .Y(new_n7668_));
  AOI22X1  g07412(.A0(new_n3652_), .A1(\b[24] ), .B0(new_n3651_), .B1(\b[23] ), .Y(new_n7669_));
  OAI21X1  g07413(.A0(new_n3778_), .A1(new_n1479_), .B0(new_n7669_), .Y(new_n7670_));
  AOI21X1  g07414(.A0(new_n3480_), .A1(new_n1572_), .B0(new_n7670_), .Y(new_n7671_));
  XOR2X1   g07415(.A(new_n7671_), .B(\a[41] ), .Y(new_n7672_));
  XOR2X1   g07416(.A(new_n7672_), .B(new_n7668_), .Y(new_n7673_));
  NOR2X1   g07417(.A(new_n7452_), .B(new_n7448_), .Y(new_n7674_));
  AOI21X1  g07418(.A0(new_n7453_), .A1(new_n7385_), .B0(new_n7674_), .Y(new_n7675_));
  XOR2X1   g07419(.A(new_n7675_), .B(new_n7673_), .Y(new_n7676_));
  AOI22X1  g07420(.A0(new_n3204_), .A1(\b[27] ), .B0(new_n3203_), .B1(\b[26] ), .Y(new_n7677_));
  OAI21X1  g07421(.A0(new_n3321_), .A1(new_n1880_), .B0(new_n7677_), .Y(new_n7678_));
  AOI21X1  g07422(.A0(new_n3080_), .A1(new_n1879_), .B0(new_n7678_), .Y(new_n7679_));
  XOR2X1   g07423(.A(new_n7679_), .B(\a[38] ), .Y(new_n7680_));
  XOR2X1   g07424(.A(new_n7680_), .B(new_n7676_), .Y(new_n7681_));
  INVX1    g07425(.A(new_n7681_), .Y(new_n7682_));
  XOR2X1   g07426(.A(new_n7457_), .B(new_n3078_), .Y(new_n7683_));
  NOR2X1   g07427(.A(new_n7461_), .B(new_n7459_), .Y(new_n7684_));
  AOI21X1  g07428(.A0(new_n7683_), .A1(new_n7454_), .B0(new_n7684_), .Y(new_n7685_));
  XOR2X1   g07429(.A(new_n7685_), .B(new_n7682_), .Y(new_n7686_));
  AOI22X1  g07430(.A0(new_n2813_), .A1(\b[30] ), .B0(new_n2812_), .B1(\b[29] ), .Y(new_n7687_));
  OAI21X1  g07431(.A0(new_n2946_), .A1(new_n2231_), .B0(new_n7687_), .Y(new_n7688_));
  AOI21X1  g07432(.A0(new_n2652_), .A1(new_n2230_), .B0(new_n7688_), .Y(new_n7689_));
  XOR2X1   g07433(.A(new_n7689_), .B(\a[35] ), .Y(new_n7690_));
  XOR2X1   g07434(.A(new_n7690_), .B(new_n7686_), .Y(new_n7691_));
  AND2X1   g07435(.A(new_n7472_), .B(new_n7468_), .Y(new_n7692_));
  AOI21X1  g07436(.A0(new_n7467_), .A1(new_n7462_), .B0(new_n7692_), .Y(new_n7693_));
  XOR2X1   g07437(.A(new_n7693_), .B(new_n7691_), .Y(new_n7694_));
  AOI22X1  g07438(.A0(new_n2545_), .A1(\b[33] ), .B0(new_n2544_), .B1(\b[32] ), .Y(new_n7695_));
  OAI21X1  g07439(.A0(new_n2543_), .A1(new_n2615_), .B0(new_n7695_), .Y(new_n7696_));
  AOI21X1  g07440(.A0(new_n2614_), .A1(new_n2260_), .B0(new_n7696_), .Y(new_n7697_));
  XOR2X1   g07441(.A(new_n7697_), .B(\a[32] ), .Y(new_n7698_));
  XOR2X1   g07442(.A(new_n7698_), .B(new_n7694_), .Y(new_n7699_));
  XOR2X1   g07443(.A(new_n7699_), .B(new_n7485_), .Y(new_n7700_));
  AOI22X1  g07444(.A0(new_n2163_), .A1(\b[36] ), .B0(new_n2162_), .B1(\b[35] ), .Y(new_n7701_));
  OAI21X1  g07445(.A0(new_n2161_), .A1(new_n2890_), .B0(new_n7701_), .Y(new_n7702_));
  AOI21X1  g07446(.A0(new_n3015_), .A1(new_n1907_), .B0(new_n7702_), .Y(new_n7703_));
  XOR2X1   g07447(.A(new_n7703_), .B(\a[29] ), .Y(new_n7704_));
  XOR2X1   g07448(.A(new_n7704_), .B(new_n7700_), .Y(new_n7705_));
  XOR2X1   g07449(.A(new_n7705_), .B(new_n7605_), .Y(new_n7706_));
  AOI22X1  g07450(.A0(new_n1814_), .A1(\b[39] ), .B0(new_n1813_), .B1(\b[38] ), .Y(new_n7707_));
  OAI21X1  g07451(.A0(new_n1812_), .A1(new_n3413_), .B0(new_n7707_), .Y(new_n7708_));
  AOI21X1  g07452(.A0(new_n3412_), .A1(new_n1617_), .B0(new_n7708_), .Y(new_n7709_));
  XOR2X1   g07453(.A(new_n7709_), .B(\a[26] ), .Y(new_n7710_));
  XOR2X1   g07454(.A(new_n7710_), .B(new_n7706_), .Y(new_n7711_));
  XOR2X1   g07455(.A(new_n7711_), .B(new_n7598_), .Y(new_n7712_));
  XOR2X1   g07456(.A(new_n7712_), .B(new_n7595_), .Y(new_n7713_));
  XOR2X1   g07457(.A(new_n7713_), .B(new_n7514_), .Y(new_n7714_));
  XOR2X1   g07458(.A(new_n7714_), .B(new_n7591_), .Y(new_n7715_));
  XOR2X1   g07459(.A(new_n7715_), .B(new_n7586_), .Y(new_n7716_));
  XOR2X1   g07460(.A(new_n7716_), .B(new_n7584_), .Y(new_n7717_));
  XOR2X1   g07461(.A(new_n7717_), .B(new_n7580_), .Y(new_n7718_));
  XOR2X1   g07462(.A(new_n7718_), .B(new_n7577_), .Y(new_n7719_));
  XOR2X1   g07463(.A(new_n7719_), .B(new_n7572_), .Y(new_n7720_));
  AOI22X1  g07464(.A0(new_n603_), .A1(\b[54] ), .B0(new_n602_), .B1(\b[53] ), .Y(new_n7721_));
  OAI21X1  g07465(.A0(new_n601_), .A1(new_n5808_), .B0(new_n7721_), .Y(new_n7722_));
  AOI21X1  g07466(.A0(new_n5807_), .A1(new_n518_), .B0(new_n7722_), .Y(new_n7723_));
  XOR2X1   g07467(.A(new_n7723_), .B(\a[11] ), .Y(new_n7724_));
  XOR2X1   g07468(.A(new_n7724_), .B(new_n7720_), .Y(new_n7725_));
  NOR2X1   g07469(.A(new_n7538_), .B(new_n7534_), .Y(new_n7726_));
  AOI21X1  g07470(.A0(new_n7539_), .A1(new_n7365_), .B0(new_n7726_), .Y(new_n7727_));
  XOR2X1   g07471(.A(new_n7727_), .B(new_n7725_), .Y(new_n7728_));
  AOI22X1  g07472(.A0(new_n469_), .A1(\b[57] ), .B0(new_n468_), .B1(\b[56] ), .Y(new_n7729_));
  OAI21X1  g07473(.A0(new_n467_), .A1(new_n6523_), .B0(new_n7729_), .Y(new_n7730_));
  AOI21X1  g07474(.A0(new_n6522_), .A1(new_n404_), .B0(new_n7730_), .Y(new_n7731_));
  XOR2X1   g07475(.A(new_n7731_), .B(\a[8] ), .Y(new_n7732_));
  XOR2X1   g07476(.A(new_n7732_), .B(new_n7728_), .Y(new_n7733_));
  AOI22X1  g07477(.A0(new_n369_), .A1(\b[60] ), .B0(new_n368_), .B1(\b[59] ), .Y(new_n7734_));
  OAI21X1  g07478(.A0(new_n367_), .A1(new_n6930_), .B0(new_n7734_), .Y(new_n7735_));
  AOI21X1  g07479(.A0(new_n6951_), .A1(new_n308_), .B0(new_n7735_), .Y(new_n7736_));
  XOR2X1   g07480(.A(new_n7736_), .B(\a[5] ), .Y(new_n7737_));
  XOR2X1   g07481(.A(new_n7737_), .B(new_n7733_), .Y(new_n7738_));
  INVX1    g07482(.A(new_n7544_), .Y(new_n7739_));
  NOR2X1   g07483(.A(new_n7549_), .B(new_n7545_), .Y(new_n7740_));
  AOI21X1  g07484(.A0(new_n7739_), .A1(new_n7540_), .B0(new_n7740_), .Y(new_n7741_));
  XOR2X1   g07485(.A(new_n7741_), .B(new_n7738_), .Y(new_n7742_));
  AND2X1   g07486(.A(\b[62] ), .B(\b[61] ), .Y(new_n7743_));
  AOI21X1  g07487(.A0(new_n7557_), .A1(new_n7556_), .B0(new_n7743_), .Y(new_n7744_));
  INVX1    g07488(.A(\b[62] ), .Y(new_n7745_));
  XOR2X1   g07489(.A(\b[63] ), .B(new_n7745_), .Y(new_n7746_));
  XOR2X1   g07490(.A(new_n7746_), .B(new_n7744_), .Y(new_n7747_));
  INVX1    g07491(.A(\b[61] ), .Y(new_n7748_));
  AOI22X1  g07492(.A0(new_n267_), .A1(\b[63] ), .B0(new_n266_), .B1(\b[62] ), .Y(new_n7749_));
  OAI21X1  g07493(.A0(new_n350_), .A1(new_n7748_), .B0(new_n7749_), .Y(new_n7750_));
  AOI21X1  g07494(.A0(new_n7747_), .A1(new_n318_), .B0(new_n7750_), .Y(new_n7751_));
  XOR2X1   g07495(.A(new_n7751_), .B(\a[2] ), .Y(new_n7752_));
  XOR2X1   g07496(.A(new_n7752_), .B(new_n7742_), .Y(new_n7753_));
  INVX1    g07497(.A(new_n7553_), .Y(new_n7754_));
  NOR2X1   g07498(.A(new_n7563_), .B(new_n7554_), .Y(new_n7755_));
  AOI21X1  g07499(.A0(new_n7754_), .A1(new_n7550_), .B0(new_n7755_), .Y(new_n7756_));
  XOR2X1   g07500(.A(new_n7756_), .B(new_n7753_), .Y(new_n7757_));
  OAI21X1  g07501(.A0(new_n7343_), .A1(new_n7360_), .B0(new_n7356_), .Y(new_n7758_));
  AND2X1   g07502(.A(new_n7564_), .B(new_n7758_), .Y(new_n7759_));
  AOI21X1  g07503(.A0(new_n7354_), .A1(new_n7353_), .B0(new_n7565_), .Y(new_n7760_));
  OR2X1    g07504(.A(new_n7760_), .B(new_n7759_), .Y(new_n7761_));
  XOR2X1   g07505(.A(new_n7761_), .B(new_n7757_), .Y(\f[63] ));
  OR2X1    g07506(.A(new_n7756_), .B(new_n7753_), .Y(new_n7763_));
  OAI21X1  g07507(.A0(new_n7760_), .A1(new_n7759_), .B0(new_n7757_), .Y(new_n7764_));
  AND2X1   g07508(.A(new_n7764_), .B(new_n7763_), .Y(new_n7765_));
  OR2X1    g07509(.A(new_n7741_), .B(new_n7738_), .Y(new_n7766_));
  XOR2X1   g07510(.A(new_n7736_), .B(new_n305_), .Y(new_n7767_));
  XOR2X1   g07511(.A(new_n7767_), .B(new_n7733_), .Y(new_n7768_));
  XOR2X1   g07512(.A(new_n7741_), .B(new_n7768_), .Y(new_n7769_));
  OR2X1    g07513(.A(new_n7752_), .B(new_n7769_), .Y(new_n7770_));
  AND2X1   g07514(.A(new_n7770_), .B(new_n7766_), .Y(new_n7771_));
  INVX1    g07515(.A(\b[63] ), .Y(new_n7772_));
  OR2X1    g07516(.A(\b[63] ), .B(new_n7745_), .Y(new_n7773_));
  AOI21X1  g07517(.A0(new_n7744_), .A1(new_n7745_), .B0(new_n7772_), .Y(new_n7774_));
  OAI22X1  g07518(.A0(new_n7774_), .A1(new_n7772_), .B0(new_n7773_), .B1(new_n7744_), .Y(new_n7775_));
  OAI22X1  g07519(.A0(new_n350_), .A1(new_n7745_), .B0(new_n284_), .B1(new_n7772_), .Y(new_n7776_));
  AOI21X1  g07520(.A0(new_n7775_), .A1(new_n318_), .B0(new_n7776_), .Y(new_n7777_));
  XOR2X1   g07521(.A(new_n7777_), .B(new_n257_), .Y(new_n7778_));
  NOR2X1   g07522(.A(new_n7732_), .B(new_n7728_), .Y(new_n7779_));
  AOI21X1  g07523(.A0(new_n7767_), .A1(new_n7733_), .B0(new_n7779_), .Y(new_n7780_));
  OR2X1    g07524(.A(new_n7724_), .B(new_n7720_), .Y(new_n7781_));
  XOR2X1   g07525(.A(new_n7718_), .B(new_n7576_), .Y(new_n7782_));
  XOR2X1   g07526(.A(new_n7782_), .B(new_n7572_), .Y(new_n7783_));
  XOR2X1   g07527(.A(new_n7724_), .B(new_n7783_), .Y(new_n7784_));
  OAI21X1  g07528(.A0(new_n7727_), .A1(new_n7784_), .B0(new_n7781_), .Y(new_n7785_));
  AOI22X1  g07529(.A0(new_n603_), .A1(\b[55] ), .B0(new_n602_), .B1(\b[54] ), .Y(new_n7786_));
  OAI21X1  g07530(.A0(new_n601_), .A1(new_n6151_), .B0(new_n7786_), .Y(new_n7787_));
  AOI21X1  g07531(.A0(new_n6150_), .A1(new_n518_), .B0(new_n7787_), .Y(new_n7788_));
  XOR2X1   g07532(.A(new_n7788_), .B(\a[11] ), .Y(new_n7789_));
  NAND2X1  g07533(.A(new_n7718_), .B(new_n7577_), .Y(new_n7790_));
  OAI21X1  g07534(.A0(new_n7782_), .A1(new_n7572_), .B0(new_n7790_), .Y(new_n7791_));
  AOI22X1  g07535(.A0(new_n818_), .A1(\b[52] ), .B0(new_n817_), .B1(\b[51] ), .Y(new_n7792_));
  OAI21X1  g07536(.A0(new_n816_), .A1(new_n5234_), .B0(new_n7792_), .Y(new_n7793_));
  AOI21X1  g07537(.A0(new_n5590_), .A1(new_n668_), .B0(new_n7793_), .Y(new_n7794_));
  XOR2X1   g07538(.A(new_n7794_), .B(\a[14] ), .Y(new_n7795_));
  INVX1    g07539(.A(new_n7795_), .Y(new_n7796_));
  INVX1    g07540(.A(new_n7584_), .Y(new_n7797_));
  NAND2X1  g07541(.A(new_n7716_), .B(new_n7797_), .Y(new_n7798_));
  OAI21X1  g07542(.A0(new_n7717_), .A1(new_n7580_), .B0(new_n7798_), .Y(new_n7799_));
  AOI22X1  g07543(.A0(new_n1017_), .A1(\b[49] ), .B0(new_n1016_), .B1(\b[48] ), .Y(new_n7800_));
  OAI21X1  g07544(.A0(new_n1015_), .A1(new_n5039_), .B0(new_n7800_), .Y(new_n7801_));
  AOI21X1  g07545(.A0(new_n5038_), .A1(new_n882_), .B0(new_n7801_), .Y(new_n7802_));
  XOR2X1   g07546(.A(new_n7802_), .B(\a[17] ), .Y(new_n7803_));
  INVX1    g07547(.A(new_n7803_), .Y(new_n7804_));
  AND2X1   g07548(.A(new_n7714_), .B(new_n7591_), .Y(new_n7805_));
  AOI21X1  g07549(.A0(new_n7715_), .A1(new_n7586_), .B0(new_n7805_), .Y(new_n7806_));
  AOI22X1  g07550(.A0(new_n1263_), .A1(\b[46] ), .B0(new_n1262_), .B1(\b[45] ), .Y(new_n7807_));
  OAI21X1  g07551(.A0(new_n1261_), .A1(new_n4336_), .B0(new_n7807_), .Y(new_n7808_));
  AOI21X1  g07552(.A0(new_n4509_), .A1(new_n1075_), .B0(new_n7808_), .Y(new_n7809_));
  XOR2X1   g07553(.A(new_n7809_), .B(\a[20] ), .Y(new_n7810_));
  INVX1    g07554(.A(new_n7595_), .Y(new_n7811_));
  NAND2X1  g07555(.A(new_n7712_), .B(new_n7811_), .Y(new_n7812_));
  OAI21X1  g07556(.A0(new_n7713_), .A1(new_n7514_), .B0(new_n7812_), .Y(new_n7813_));
  NOR2X1   g07557(.A(new_n7636_), .B(new_n7632_), .Y(new_n7814_));
  AOI21X1  g07558(.A0(new_n7637_), .A1(new_n7622_), .B0(new_n7814_), .Y(new_n7815_));
  INVX1    g07559(.A(new_n7815_), .Y(new_n7816_));
  INVX1    g07560(.A(new_n7624_), .Y(new_n7817_));
  AND2X1   g07561(.A(\a[63] ), .B(\a[62] ), .Y(new_n7818_));
  AOI22X1  g07562(.A0(new_n7818_), .A1(\b[0] ), .B0(new_n7817_), .B1(\b[1] ), .Y(new_n7819_));
  AND2X1   g07563(.A(new_n7187_), .B(new_n323_), .Y(new_n7820_));
  NOR4X1   g07564(.A(new_n7188_), .B(new_n7186_), .C(new_n7191_), .D(new_n277_), .Y(new_n7821_));
  OAI22X1  g07565(.A0(new_n7193_), .A1(new_n325_), .B0(new_n7190_), .B1(new_n297_), .Y(new_n7822_));
  NOR3X1   g07566(.A(new_n7822_), .B(new_n7821_), .C(new_n7820_), .Y(new_n7823_));
  XOR2X1   g07567(.A(new_n7823_), .B(\a[62] ), .Y(new_n7824_));
  XOR2X1   g07568(.A(new_n7824_), .B(new_n7819_), .Y(new_n7825_));
  AND2X1   g07569(.A(new_n7625_), .B(new_n7623_), .Y(new_n7826_));
  INVX1    g07570(.A(new_n7631_), .Y(new_n7827_));
  AOI21X1  g07571(.A0(new_n7827_), .A1(new_n7626_), .B0(new_n7826_), .Y(new_n7828_));
  XOR2X1   g07572(.A(new_n7828_), .B(new_n7825_), .Y(new_n7829_));
  AOI22X1  g07573(.A0(new_n6603_), .A1(\b[7] ), .B0(new_n6600_), .B1(\b[6] ), .Y(new_n7830_));
  OAI21X1  g07574(.A0(new_n6804_), .A1(new_n395_), .B0(new_n7830_), .Y(new_n7831_));
  AOI21X1  g07575(.A0(new_n6598_), .A1(new_n394_), .B0(new_n7831_), .Y(new_n7832_));
  XOR2X1   g07576(.A(new_n7832_), .B(\a[59] ), .Y(new_n7833_));
  XOR2X1   g07577(.A(new_n7833_), .B(new_n7829_), .Y(new_n7834_));
  XOR2X1   g07578(.A(new_n7834_), .B(new_n7816_), .Y(new_n7835_));
  AOI22X1  g07579(.A0(new_n6438_), .A1(\b[10] ), .B0(new_n6437_), .B1(\b[9] ), .Y(new_n7836_));
  OAI21X1  g07580(.A0(new_n6436_), .A1(new_n489_), .B0(new_n7836_), .Y(new_n7837_));
  AOI21X1  g07581(.A0(new_n6023_), .A1(new_n543_), .B0(new_n7837_), .Y(new_n7838_));
  XOR2X1   g07582(.A(new_n7838_), .B(\a[56] ), .Y(new_n7839_));
  XOR2X1   g07583(.A(new_n7839_), .B(new_n7835_), .Y(new_n7840_));
  XOR2X1   g07584(.A(new_n7641_), .B(new_n6019_), .Y(new_n7841_));
  AND2X1   g07585(.A(new_n7841_), .B(new_n7638_), .Y(new_n7842_));
  INVX1    g07586(.A(new_n7643_), .Y(new_n7843_));
  AOI21X1  g07587(.A0(new_n7843_), .A1(new_n7621_), .B0(new_n7842_), .Y(new_n7844_));
  XOR2X1   g07588(.A(new_n7844_), .B(new_n7840_), .Y(new_n7845_));
  INVX1    g07589(.A(new_n7845_), .Y(new_n7846_));
  AOI22X1  g07590(.A0(new_n5430_), .A1(\b[13] ), .B0(new_n5427_), .B1(\b[12] ), .Y(new_n7847_));
  OAI21X1  g07591(.A0(new_n5891_), .A1(new_n716_), .B0(new_n7847_), .Y(new_n7848_));
  AOI21X1  g07592(.A0(new_n5425_), .A1(new_n715_), .B0(new_n7848_), .Y(new_n7849_));
  XOR2X1   g07593(.A(new_n7849_), .B(\a[53] ), .Y(new_n7850_));
  XOR2X1   g07594(.A(new_n7850_), .B(new_n7846_), .Y(new_n7851_));
  INVX1    g07595(.A(new_n7851_), .Y(new_n7852_));
  NOR2X1   g07596(.A(new_n7648_), .B(new_n7644_), .Y(new_n7853_));
  AOI21X1  g07597(.A0(new_n7649_), .A1(new_n7619_), .B0(new_n7853_), .Y(new_n7854_));
  XOR2X1   g07598(.A(new_n7854_), .B(new_n7852_), .Y(new_n7855_));
  AOI22X1  g07599(.A0(new_n4880_), .A1(\b[16] ), .B0(new_n4877_), .B1(\b[15] ), .Y(new_n7856_));
  OAI21X1  g07600(.A0(new_n5291_), .A1(new_n792_), .B0(new_n7856_), .Y(new_n7857_));
  AOI21X1  g07601(.A0(new_n4875_), .A1(new_n842_), .B0(new_n7857_), .Y(new_n7858_));
  XOR2X1   g07602(.A(new_n7858_), .B(\a[50] ), .Y(new_n7859_));
  XOR2X1   g07603(.A(new_n7859_), .B(new_n7855_), .Y(new_n7860_));
  INVX1    g07604(.A(new_n7654_), .Y(new_n7861_));
  NOR2X1   g07605(.A(new_n7659_), .B(new_n7655_), .Y(new_n7862_));
  AOI21X1  g07606(.A0(new_n7861_), .A1(new_n7650_), .B0(new_n7862_), .Y(new_n7863_));
  XOR2X1   g07607(.A(new_n7863_), .B(new_n7860_), .Y(new_n7864_));
  INVX1    g07608(.A(new_n7864_), .Y(new_n7865_));
  AOI22X1  g07609(.A0(new_n4572_), .A1(\b[19] ), .B0(new_n4571_), .B1(\b[18] ), .Y(new_n7866_));
  OAI21X1  g07610(.A0(new_n4740_), .A1(new_n1118_), .B0(new_n7866_), .Y(new_n7867_));
  AOI21X1  g07611(.A0(new_n4375_), .A1(new_n1117_), .B0(new_n7867_), .Y(new_n7868_));
  XOR2X1   g07612(.A(new_n7868_), .B(\a[47] ), .Y(new_n7869_));
  XOR2X1   g07613(.A(new_n7869_), .B(new_n7865_), .Y(new_n7870_));
  NOR2X1   g07614(.A(new_n7664_), .B(new_n7660_), .Y(new_n7871_));
  AOI21X1  g07615(.A0(new_n7665_), .A1(new_n7616_), .B0(new_n7871_), .Y(new_n7872_));
  XOR2X1   g07616(.A(new_n7872_), .B(new_n7870_), .Y(new_n7873_));
  AOI22X1  g07617(.A0(new_n4095_), .A1(\b[22] ), .B0(new_n4094_), .B1(\b[21] ), .Y(new_n7874_));
  OAI21X1  g07618(.A0(new_n4233_), .A1(new_n1297_), .B0(new_n7874_), .Y(new_n7875_));
  AOI21X1  g07619(.A0(new_n3901_), .A1(new_n1399_), .B0(new_n7875_), .Y(new_n7876_));
  XOR2X1   g07620(.A(new_n7876_), .B(\a[44] ), .Y(new_n7877_));
  XOR2X1   g07621(.A(new_n7877_), .B(new_n7873_), .Y(new_n7878_));
  AND2X1   g07622(.A(new_n7666_), .B(new_n7612_), .Y(new_n7879_));
  AOI21X1  g07623(.A0(new_n7667_), .A1(new_n7608_), .B0(new_n7879_), .Y(new_n7880_));
  XOR2X1   g07624(.A(new_n7880_), .B(new_n7878_), .Y(new_n7881_));
  AOI22X1  g07625(.A0(new_n3652_), .A1(\b[25] ), .B0(new_n3651_), .B1(\b[24] ), .Y(new_n7882_));
  OAI21X1  g07626(.A0(new_n3778_), .A1(new_n1591_), .B0(new_n7882_), .Y(new_n7883_));
  AOI21X1  g07627(.A0(new_n3480_), .A1(new_n1590_), .B0(new_n7883_), .Y(new_n7884_));
  XOR2X1   g07628(.A(new_n7884_), .B(\a[41] ), .Y(new_n7885_));
  XOR2X1   g07629(.A(new_n7885_), .B(new_n7881_), .Y(new_n7886_));
  XOR2X1   g07630(.A(new_n7671_), .B(new_n3478_), .Y(new_n7887_));
  AND2X1   g07631(.A(new_n7887_), .B(new_n7668_), .Y(new_n7888_));
  NOR2X1   g07632(.A(new_n7675_), .B(new_n7673_), .Y(new_n7889_));
  OR2X1    g07633(.A(new_n7889_), .B(new_n7888_), .Y(new_n7890_));
  XOR2X1   g07634(.A(new_n7890_), .B(new_n7886_), .Y(new_n7891_));
  AOI22X1  g07635(.A0(new_n3204_), .A1(\b[28] ), .B0(new_n3203_), .B1(\b[27] ), .Y(new_n7892_));
  OAI21X1  g07636(.A0(new_n3321_), .A1(new_n1877_), .B0(new_n7892_), .Y(new_n7893_));
  AOI21X1  g07637(.A0(new_n3080_), .A1(new_n2004_), .B0(new_n7893_), .Y(new_n7894_));
  XOR2X1   g07638(.A(new_n7894_), .B(\a[38] ), .Y(new_n7895_));
  XOR2X1   g07639(.A(new_n7895_), .B(new_n7891_), .Y(new_n7896_));
  XOR2X1   g07640(.A(new_n7679_), .B(new_n3078_), .Y(new_n7897_));
  NAND2X1  g07641(.A(new_n7897_), .B(new_n7676_), .Y(new_n7898_));
  OAI21X1  g07642(.A0(new_n7685_), .A1(new_n7681_), .B0(new_n7898_), .Y(new_n7899_));
  XOR2X1   g07643(.A(new_n7899_), .B(new_n7896_), .Y(new_n7900_));
  AOI22X1  g07644(.A0(new_n2813_), .A1(\b[31] ), .B0(new_n2812_), .B1(\b[30] ), .Y(new_n7901_));
  OAI21X1  g07645(.A0(new_n2946_), .A1(new_n2359_), .B0(new_n7901_), .Y(new_n7902_));
  AOI21X1  g07646(.A0(new_n2652_), .A1(new_n2358_), .B0(new_n7902_), .Y(new_n7903_));
  XOR2X1   g07647(.A(new_n7903_), .B(\a[35] ), .Y(new_n7904_));
  XOR2X1   g07648(.A(new_n7904_), .B(new_n7900_), .Y(new_n7905_));
  AND2X1   g07649(.A(new_n7690_), .B(new_n7686_), .Y(new_n7906_));
  OR2X1    g07650(.A(new_n7690_), .B(new_n7686_), .Y(new_n7907_));
  OAI21X1  g07651(.A0(new_n7693_), .A1(new_n7906_), .B0(new_n7907_), .Y(new_n7908_));
  XOR2X1   g07652(.A(new_n7908_), .B(new_n7905_), .Y(new_n7909_));
  AOI22X1  g07653(.A0(new_n2545_), .A1(\b[34] ), .B0(new_n2544_), .B1(\b[33] ), .Y(new_n7910_));
  OAI21X1  g07654(.A0(new_n2543_), .A1(new_n2612_), .B0(new_n7910_), .Y(new_n7911_));
  AOI21X1  g07655(.A0(new_n2759_), .A1(new_n2260_), .B0(new_n7911_), .Y(new_n7912_));
  XOR2X1   g07656(.A(new_n7912_), .B(\a[32] ), .Y(new_n7913_));
  XOR2X1   g07657(.A(new_n7913_), .B(new_n7909_), .Y(new_n7914_));
  NOR2X1   g07658(.A(new_n7698_), .B(new_n7694_), .Y(new_n7915_));
  AOI21X1  g07659(.A0(new_n7699_), .A1(new_n7602_), .B0(new_n7915_), .Y(new_n7916_));
  XOR2X1   g07660(.A(new_n7916_), .B(new_n7914_), .Y(new_n7917_));
  AOI22X1  g07661(.A0(new_n2163_), .A1(\b[37] ), .B0(new_n2162_), .B1(\b[36] ), .Y(new_n7918_));
  OAI21X1  g07662(.A0(new_n2161_), .A1(new_n3156_), .B0(new_n7918_), .Y(new_n7919_));
  AOI21X1  g07663(.A0(new_n3155_), .A1(new_n1907_), .B0(new_n7919_), .Y(new_n7920_));
  XOR2X1   g07664(.A(new_n7920_), .B(\a[29] ), .Y(new_n7921_));
  XOR2X1   g07665(.A(new_n7921_), .B(new_n7917_), .Y(new_n7922_));
  NOR2X1   g07666(.A(new_n7704_), .B(new_n7700_), .Y(new_n7923_));
  AOI21X1  g07667(.A0(new_n7705_), .A1(new_n7605_), .B0(new_n7923_), .Y(new_n7924_));
  XOR2X1   g07668(.A(new_n7924_), .B(new_n7922_), .Y(new_n7925_));
  AOI22X1  g07669(.A0(new_n1814_), .A1(\b[40] ), .B0(new_n1813_), .B1(\b[39] ), .Y(new_n7926_));
  OAI21X1  g07670(.A0(new_n1812_), .A1(new_n3575_), .B0(new_n7926_), .Y(new_n7927_));
  AOI21X1  g07671(.A0(new_n3574_), .A1(new_n1617_), .B0(new_n7927_), .Y(new_n7928_));
  XOR2X1   g07672(.A(new_n7928_), .B(\a[26] ), .Y(new_n7929_));
  XOR2X1   g07673(.A(new_n7929_), .B(new_n7925_), .Y(new_n7930_));
  XOR2X1   g07674(.A(new_n7709_), .B(new_n1621_), .Y(new_n7931_));
  NAND2X1  g07675(.A(new_n7931_), .B(new_n7706_), .Y(new_n7932_));
  OAI21X1  g07676(.A0(new_n7711_), .A1(new_n7598_), .B0(new_n7932_), .Y(new_n7933_));
  XOR2X1   g07677(.A(new_n7933_), .B(new_n7930_), .Y(new_n7934_));
  AOI22X1  g07678(.A0(new_n1526_), .A1(\b[43] ), .B0(new_n1525_), .B1(\b[42] ), .Y(new_n7935_));
  OAI21X1  g07679(.A0(new_n1524_), .A1(new_n4015_), .B0(new_n7935_), .Y(new_n7936_));
  AOI21X1  g07680(.A0(new_n4014_), .A1(new_n1347_), .B0(new_n7936_), .Y(new_n7937_));
  XOR2X1   g07681(.A(new_n7937_), .B(\a[23] ), .Y(new_n7938_));
  XOR2X1   g07682(.A(new_n7938_), .B(new_n7934_), .Y(new_n7939_));
  XOR2X1   g07683(.A(new_n7939_), .B(new_n7813_), .Y(new_n7940_));
  XOR2X1   g07684(.A(new_n7940_), .B(new_n7810_), .Y(new_n7941_));
  XOR2X1   g07685(.A(new_n7941_), .B(new_n7806_), .Y(new_n7942_));
  XOR2X1   g07686(.A(new_n7942_), .B(new_n7804_), .Y(new_n7943_));
  XOR2X1   g07687(.A(new_n7943_), .B(new_n7799_), .Y(new_n7944_));
  XOR2X1   g07688(.A(new_n7944_), .B(new_n7796_), .Y(new_n7945_));
  XOR2X1   g07689(.A(new_n7945_), .B(new_n7791_), .Y(new_n7946_));
  XOR2X1   g07690(.A(new_n7946_), .B(new_n7789_), .Y(new_n7947_));
  XOR2X1   g07691(.A(new_n7947_), .B(new_n7785_), .Y(new_n7948_));
  AOI22X1  g07692(.A0(new_n469_), .A1(\b[58] ), .B0(new_n468_), .B1(\b[57] ), .Y(new_n7949_));
  OAI21X1  g07693(.A0(new_n467_), .A1(new_n6520_), .B0(new_n7949_), .Y(new_n7950_));
  AOI21X1  g07694(.A0(new_n6732_), .A1(new_n404_), .B0(new_n7950_), .Y(new_n7951_));
  XOR2X1   g07695(.A(new_n7951_), .B(\a[8] ), .Y(new_n7952_));
  XOR2X1   g07696(.A(new_n7952_), .B(new_n7948_), .Y(new_n7953_));
  AOI22X1  g07697(.A0(new_n369_), .A1(\b[61] ), .B0(new_n368_), .B1(\b[60] ), .Y(new_n7954_));
  OAI21X1  g07698(.A0(new_n367_), .A1(new_n7339_), .B0(new_n7954_), .Y(new_n7955_));
  AOI21X1  g07699(.A0(new_n7338_), .A1(new_n308_), .B0(new_n7955_), .Y(new_n7956_));
  XOR2X1   g07700(.A(new_n7956_), .B(\a[5] ), .Y(new_n7957_));
  XOR2X1   g07701(.A(new_n7957_), .B(new_n7953_), .Y(new_n7958_));
  XOR2X1   g07702(.A(new_n7958_), .B(new_n7780_), .Y(new_n7959_));
  XOR2X1   g07703(.A(new_n7959_), .B(new_n7778_), .Y(new_n7960_));
  XOR2X1   g07704(.A(new_n7960_), .B(new_n7771_), .Y(new_n7961_));
  XOR2X1   g07705(.A(new_n7961_), .B(new_n7765_), .Y(\f[64] ));
  AND2X1   g07706(.A(new_n7942_), .B(new_n7804_), .Y(new_n7963_));
  AOI21X1  g07707(.A0(new_n7943_), .A1(new_n7799_), .B0(new_n7963_), .Y(new_n7964_));
  INVX1    g07708(.A(new_n7810_), .Y(new_n7965_));
  NOR2X1   g07709(.A(new_n7941_), .B(new_n7806_), .Y(new_n7966_));
  AOI21X1  g07710(.A0(new_n7940_), .A1(new_n7965_), .B0(new_n7966_), .Y(new_n7967_));
  AOI22X1  g07711(.A0(new_n1263_), .A1(\b[47] ), .B0(new_n1262_), .B1(\b[46] ), .Y(new_n7968_));
  OAI21X1  g07712(.A0(new_n1261_), .A1(new_n4674_), .B0(new_n7968_), .Y(new_n7969_));
  AOI21X1  g07713(.A0(new_n4673_), .A1(new_n1075_), .B0(new_n7969_), .Y(new_n7970_));
  XOR2X1   g07714(.A(new_n7970_), .B(\a[20] ), .Y(new_n7971_));
  NOR2X1   g07715(.A(new_n7904_), .B(new_n7900_), .Y(new_n7972_));
  AOI21X1  g07716(.A0(new_n7908_), .A1(new_n7905_), .B0(new_n7972_), .Y(new_n7973_));
  OR2X1    g07717(.A(new_n7877_), .B(new_n7873_), .Y(new_n7974_));
  INVX1    g07718(.A(new_n7878_), .Y(new_n7975_));
  OAI21X1  g07719(.A0(new_n7880_), .A1(new_n7975_), .B0(new_n7974_), .Y(new_n7976_));
  AND2X1   g07720(.A(new_n7869_), .B(new_n7865_), .Y(new_n7977_));
  OR2X1    g07721(.A(new_n7869_), .B(new_n7865_), .Y(new_n7978_));
  OAI21X1  g07722(.A0(new_n7872_), .A1(new_n7977_), .B0(new_n7978_), .Y(new_n7979_));
  XOR2X1   g07723(.A(new_n7858_), .B(new_n4873_), .Y(new_n7980_));
  AND2X1   g07724(.A(new_n7980_), .B(new_n7855_), .Y(new_n7981_));
  INVX1    g07725(.A(new_n7981_), .Y(new_n7982_));
  OAI21X1  g07726(.A0(new_n7863_), .A1(new_n7860_), .B0(new_n7982_), .Y(new_n7983_));
  OR2X1    g07727(.A(new_n7850_), .B(new_n7846_), .Y(new_n7984_));
  OAI21X1  g07728(.A0(new_n7854_), .A1(new_n7852_), .B0(new_n7984_), .Y(new_n7985_));
  XOR2X1   g07729(.A(new_n7838_), .B(new_n6019_), .Y(new_n7986_));
  NOR2X1   g07730(.A(new_n7844_), .B(new_n7840_), .Y(new_n7987_));
  AOI21X1  g07731(.A0(new_n7986_), .A1(new_n7835_), .B0(new_n7987_), .Y(new_n7988_));
  INVX1    g07732(.A(new_n7988_), .Y(new_n7989_));
  NOR2X1   g07733(.A(new_n7833_), .B(new_n7829_), .Y(new_n7990_));
  AOI21X1  g07734(.A0(new_n7834_), .A1(new_n7816_), .B0(new_n7990_), .Y(new_n7991_));
  INVX1    g07735(.A(new_n7991_), .Y(new_n7992_));
  AOI22X1  g07736(.A0(new_n7818_), .A1(\b[1] ), .B0(new_n7817_), .B1(\b[2] ), .Y(new_n7993_));
  AOI22X1  g07737(.A0(new_n7192_), .A1(\b[5] ), .B0(new_n7189_), .B1(\b[4] ), .Y(new_n7994_));
  OAI21X1  g07738(.A0(new_n7627_), .A1(new_n297_), .B0(new_n7994_), .Y(new_n7995_));
  AOI21X1  g07739(.A0(new_n7187_), .A1(new_n349_), .B0(new_n7995_), .Y(new_n7996_));
  XOR2X1   g07740(.A(new_n7996_), .B(\a[62] ), .Y(new_n7997_));
  XOR2X1   g07741(.A(new_n7997_), .B(new_n7993_), .Y(new_n7998_));
  INVX1    g07742(.A(new_n7998_), .Y(new_n7999_));
  OR2X1    g07743(.A(new_n7824_), .B(new_n7819_), .Y(new_n8000_));
  INVX1    g07744(.A(new_n7825_), .Y(new_n8001_));
  OR2X1    g07745(.A(new_n7828_), .B(new_n8001_), .Y(new_n8002_));
  AND2X1   g07746(.A(new_n8002_), .B(new_n8000_), .Y(new_n8003_));
  XOR2X1   g07747(.A(new_n8003_), .B(new_n7999_), .Y(new_n8004_));
  INVX1    g07748(.A(new_n8004_), .Y(new_n8005_));
  AOI22X1  g07749(.A0(new_n6603_), .A1(\b[8] ), .B0(new_n6600_), .B1(\b[7] ), .Y(new_n8006_));
  OAI21X1  g07750(.A0(new_n6804_), .A1(new_n392_), .B0(new_n8006_), .Y(new_n8007_));
  AOI21X1  g07751(.A0(new_n6598_), .A1(new_n454_), .B0(new_n8007_), .Y(new_n8008_));
  XOR2X1   g07752(.A(new_n8008_), .B(\a[59] ), .Y(new_n8009_));
  AND2X1   g07753(.A(new_n8009_), .B(new_n8005_), .Y(new_n8010_));
  INVX1    g07754(.A(new_n8010_), .Y(new_n8011_));
  XOR2X1   g07755(.A(new_n8009_), .B(new_n8004_), .Y(new_n8012_));
  NOR2X1   g07756(.A(new_n8009_), .B(new_n8005_), .Y(new_n8013_));
  AOI21X1  g07757(.A0(new_n8011_), .A1(new_n7992_), .B0(new_n8013_), .Y(new_n8014_));
  AOI22X1  g07758(.A0(new_n8014_), .A1(new_n8011_), .B0(new_n8012_), .B1(new_n7992_), .Y(new_n8015_));
  AOI22X1  g07759(.A0(new_n6438_), .A1(\b[11] ), .B0(new_n6437_), .B1(\b[10] ), .Y(new_n8016_));
  OAI21X1  g07760(.A0(new_n6436_), .A1(new_n590_), .B0(new_n8016_), .Y(new_n8017_));
  AOI21X1  g07761(.A0(new_n6023_), .A1(new_n589_), .B0(new_n8017_), .Y(new_n8018_));
  XOR2X1   g07762(.A(new_n8018_), .B(\a[56] ), .Y(new_n8019_));
  XOR2X1   g07763(.A(new_n8019_), .B(new_n8015_), .Y(new_n8020_));
  XOR2X1   g07764(.A(new_n8020_), .B(new_n7989_), .Y(new_n8021_));
  AOI22X1  g07765(.A0(new_n5430_), .A1(\b[14] ), .B0(new_n5427_), .B1(\b[13] ), .Y(new_n8022_));
  OAI21X1  g07766(.A0(new_n5891_), .A1(new_n713_), .B0(new_n8022_), .Y(new_n8023_));
  AOI21X1  g07767(.A0(new_n5425_), .A1(new_n734_), .B0(new_n8023_), .Y(new_n8024_));
  XOR2X1   g07768(.A(new_n8024_), .B(\a[53] ), .Y(new_n8025_));
  XOR2X1   g07769(.A(new_n8025_), .B(new_n8021_), .Y(new_n8026_));
  XOR2X1   g07770(.A(new_n8026_), .B(new_n7985_), .Y(new_n8027_));
  AOI22X1  g07771(.A0(new_n4880_), .A1(\b[17] ), .B0(new_n4877_), .B1(\b[16] ), .Y(new_n8028_));
  OAI21X1  g07772(.A0(new_n5291_), .A1(new_n977_), .B0(new_n8028_), .Y(new_n8029_));
  AOI21X1  g07773(.A0(new_n4875_), .A1(new_n976_), .B0(new_n8029_), .Y(new_n8030_));
  XOR2X1   g07774(.A(new_n8030_), .B(\a[50] ), .Y(new_n8031_));
  XOR2X1   g07775(.A(new_n8031_), .B(new_n8027_), .Y(new_n8032_));
  XOR2X1   g07776(.A(new_n8032_), .B(new_n7983_), .Y(new_n8033_));
  AOI22X1  g07777(.A0(new_n4572_), .A1(\b[20] ), .B0(new_n4571_), .B1(\b[19] ), .Y(new_n8034_));
  OAI21X1  g07778(.A0(new_n4740_), .A1(new_n1115_), .B0(new_n8034_), .Y(new_n8035_));
  AOI21X1  g07779(.A0(new_n4375_), .A1(new_n1217_), .B0(new_n8035_), .Y(new_n8036_));
  XOR2X1   g07780(.A(new_n8036_), .B(\a[47] ), .Y(new_n8037_));
  XOR2X1   g07781(.A(new_n8037_), .B(new_n8033_), .Y(new_n8038_));
  XOR2X1   g07782(.A(new_n8038_), .B(new_n7979_), .Y(new_n8039_));
  AOI22X1  g07783(.A0(new_n4095_), .A1(\b[23] ), .B0(new_n4094_), .B1(\b[22] ), .Y(new_n8040_));
  OAI21X1  g07784(.A0(new_n4233_), .A1(new_n1482_), .B0(new_n8040_), .Y(new_n8041_));
  AOI21X1  g07785(.A0(new_n3901_), .A1(new_n1481_), .B0(new_n8041_), .Y(new_n8042_));
  XOR2X1   g07786(.A(new_n8042_), .B(\a[44] ), .Y(new_n8043_));
  XOR2X1   g07787(.A(new_n8043_), .B(new_n8039_), .Y(new_n8044_));
  XOR2X1   g07788(.A(new_n8044_), .B(new_n7976_), .Y(new_n8045_));
  AOI22X1  g07789(.A0(new_n3652_), .A1(\b[26] ), .B0(new_n3651_), .B1(\b[25] ), .Y(new_n8046_));
  OAI21X1  g07790(.A0(new_n3778_), .A1(new_n1588_), .B0(new_n8046_), .Y(new_n8047_));
  AOI21X1  g07791(.A0(new_n3480_), .A1(new_n1783_), .B0(new_n8047_), .Y(new_n8048_));
  XOR2X1   g07792(.A(new_n8048_), .B(\a[41] ), .Y(new_n8049_));
  INVX1    g07793(.A(new_n8049_), .Y(new_n8050_));
  XOR2X1   g07794(.A(new_n8050_), .B(new_n8045_), .Y(new_n8051_));
  NOR2X1   g07795(.A(new_n7885_), .B(new_n7881_), .Y(new_n8052_));
  AOI21X1  g07796(.A0(new_n7890_), .A1(new_n7886_), .B0(new_n8052_), .Y(new_n8053_));
  XOR2X1   g07797(.A(new_n8053_), .B(new_n8051_), .Y(new_n8054_));
  AOI22X1  g07798(.A0(new_n3204_), .A1(\b[29] ), .B0(new_n3203_), .B1(\b[28] ), .Y(new_n8055_));
  OAI21X1  g07799(.A0(new_n3321_), .A1(new_n2126_), .B0(new_n8055_), .Y(new_n8056_));
  AOI21X1  g07800(.A0(new_n3080_), .A1(new_n2125_), .B0(new_n8056_), .Y(new_n8057_));
  XOR2X1   g07801(.A(new_n8057_), .B(\a[38] ), .Y(new_n8058_));
  XOR2X1   g07802(.A(new_n8058_), .B(new_n8054_), .Y(new_n8059_));
  NOR2X1   g07803(.A(new_n7889_), .B(new_n7888_), .Y(new_n8060_));
  XOR2X1   g07804(.A(new_n8060_), .B(new_n7886_), .Y(new_n8061_));
  NOR2X1   g07805(.A(new_n7895_), .B(new_n8061_), .Y(new_n8062_));
  XOR2X1   g07806(.A(new_n7895_), .B(new_n8061_), .Y(new_n8063_));
  AOI21X1  g07807(.A0(new_n7899_), .A1(new_n8063_), .B0(new_n8062_), .Y(new_n8064_));
  XOR2X1   g07808(.A(new_n8064_), .B(new_n8059_), .Y(new_n8065_));
  AOI22X1  g07809(.A0(new_n2813_), .A1(\b[32] ), .B0(new_n2812_), .B1(\b[31] ), .Y(new_n8066_));
  OAI21X1  g07810(.A0(new_n2946_), .A1(new_n2356_), .B0(new_n8066_), .Y(new_n8067_));
  AOI21X1  g07811(.A0(new_n2652_), .A1(new_n2495_), .B0(new_n8067_), .Y(new_n8068_));
  XOR2X1   g07812(.A(new_n8068_), .B(\a[35] ), .Y(new_n8069_));
  AND2X1   g07813(.A(new_n8069_), .B(new_n8065_), .Y(new_n8070_));
  XOR2X1   g07814(.A(new_n8069_), .B(new_n8065_), .Y(new_n8071_));
  OR2X1    g07815(.A(new_n8069_), .B(new_n8065_), .Y(new_n8072_));
  OAI21X1  g07816(.A0(new_n8070_), .A1(new_n7973_), .B0(new_n8072_), .Y(new_n8073_));
  OAI22X1  g07817(.A0(new_n8073_), .A1(new_n8070_), .B0(new_n8071_), .B1(new_n7973_), .Y(new_n8074_));
  AOI22X1  g07818(.A0(new_n2545_), .A1(\b[35] ), .B0(new_n2544_), .B1(\b[34] ), .Y(new_n8075_));
  OAI21X1  g07819(.A0(new_n2543_), .A1(new_n2893_), .B0(new_n8075_), .Y(new_n8076_));
  AOI21X1  g07820(.A0(new_n2892_), .A1(new_n2260_), .B0(new_n8076_), .Y(new_n8077_));
  XOR2X1   g07821(.A(new_n8077_), .B(\a[32] ), .Y(new_n8078_));
  XOR2X1   g07822(.A(new_n8078_), .B(new_n8074_), .Y(new_n8079_));
  INVX1    g07823(.A(new_n7913_), .Y(new_n8080_));
  NOR2X1   g07824(.A(new_n7916_), .B(new_n7914_), .Y(new_n8081_));
  AOI21X1  g07825(.A0(new_n8080_), .A1(new_n7909_), .B0(new_n8081_), .Y(new_n8082_));
  XOR2X1   g07826(.A(new_n8082_), .B(new_n8079_), .Y(new_n8083_));
  AOI22X1  g07827(.A0(new_n2163_), .A1(\b[38] ), .B0(new_n2162_), .B1(\b[37] ), .Y(new_n8084_));
  OAI21X1  g07828(.A0(new_n2161_), .A1(new_n3276_), .B0(new_n8084_), .Y(new_n8085_));
  AOI21X1  g07829(.A0(new_n3275_), .A1(new_n1907_), .B0(new_n8085_), .Y(new_n8086_));
  XOR2X1   g07830(.A(new_n8086_), .B(\a[29] ), .Y(new_n8087_));
  XOR2X1   g07831(.A(new_n8087_), .B(new_n8083_), .Y(new_n8088_));
  INVX1    g07832(.A(new_n7914_), .Y(new_n8089_));
  XOR2X1   g07833(.A(new_n7916_), .B(new_n8089_), .Y(new_n8090_));
  OR2X1    g07834(.A(new_n7921_), .B(new_n8090_), .Y(new_n8091_));
  OAI21X1  g07835(.A0(new_n7924_), .A1(new_n7922_), .B0(new_n8091_), .Y(new_n8092_));
  XOR2X1   g07836(.A(new_n8092_), .B(new_n8088_), .Y(new_n8093_));
  AOI22X1  g07837(.A0(new_n1814_), .A1(\b[41] ), .B0(new_n1813_), .B1(\b[40] ), .Y(new_n8094_));
  OAI21X1  g07838(.A0(new_n1812_), .A1(new_n3723_), .B0(new_n8094_), .Y(new_n8095_));
  AOI21X1  g07839(.A0(new_n3722_), .A1(new_n1617_), .B0(new_n8095_), .Y(new_n8096_));
  XOR2X1   g07840(.A(new_n8096_), .B(\a[26] ), .Y(new_n8097_));
  NAND2X1  g07841(.A(new_n8097_), .B(new_n8093_), .Y(new_n8098_));
  XOR2X1   g07842(.A(new_n7921_), .B(new_n8090_), .Y(new_n8099_));
  XOR2X1   g07843(.A(new_n7924_), .B(new_n8099_), .Y(new_n8100_));
  NOR2X1   g07844(.A(new_n7929_), .B(new_n8100_), .Y(new_n8101_));
  XOR2X1   g07845(.A(new_n7929_), .B(new_n8100_), .Y(new_n8102_));
  AOI21X1  g07846(.A0(new_n7933_), .A1(new_n8102_), .B0(new_n8101_), .Y(new_n8103_));
  OR2X1    g07847(.A(new_n8097_), .B(new_n8093_), .Y(new_n8104_));
  AOI21X1  g07848(.A0(new_n8098_), .A1(new_n8104_), .B0(new_n8103_), .Y(new_n8105_));
  NOR2X1   g07849(.A(new_n8097_), .B(new_n8093_), .Y(new_n8106_));
  AND2X1   g07850(.A(new_n8097_), .B(new_n8093_), .Y(new_n8107_));
  NOR3X1   g07851(.A(new_n8107_), .B(new_n8106_), .C(new_n8103_), .Y(new_n8108_));
  NOR2X1   g07852(.A(new_n8108_), .B(new_n8106_), .Y(new_n8109_));
  AOI21X1  g07853(.A0(new_n8109_), .A1(new_n8098_), .B0(new_n8105_), .Y(new_n8110_));
  AOI22X1  g07854(.A0(new_n1526_), .A1(\b[44] ), .B0(new_n1525_), .B1(\b[43] ), .Y(new_n8111_));
  OAI21X1  g07855(.A0(new_n1524_), .A1(new_n4012_), .B0(new_n8111_), .Y(new_n8112_));
  AOI21X1  g07856(.A0(new_n4178_), .A1(new_n1347_), .B0(new_n8112_), .Y(new_n8113_));
  XOR2X1   g07857(.A(new_n8113_), .B(\a[23] ), .Y(new_n8114_));
  INVX1    g07858(.A(new_n8114_), .Y(new_n8115_));
  XOR2X1   g07859(.A(new_n8115_), .B(new_n8110_), .Y(new_n8116_));
  NOR2X1   g07860(.A(new_n7938_), .B(new_n7934_), .Y(new_n8117_));
  AOI21X1  g07861(.A0(new_n7939_), .A1(new_n7813_), .B0(new_n8117_), .Y(new_n8118_));
  XOR2X1   g07862(.A(new_n8118_), .B(new_n8116_), .Y(new_n8119_));
  XOR2X1   g07863(.A(new_n8119_), .B(new_n7971_), .Y(new_n8120_));
  XOR2X1   g07864(.A(new_n8120_), .B(new_n7967_), .Y(new_n8121_));
  AOI22X1  g07865(.A0(new_n1017_), .A1(\b[50] ), .B0(new_n1016_), .B1(\b[49] ), .Y(new_n8122_));
  OAI21X1  g07866(.A0(new_n1015_), .A1(new_n5036_), .B0(new_n8122_), .Y(new_n8123_));
  AOI21X1  g07867(.A0(new_n5204_), .A1(new_n882_), .B0(new_n8123_), .Y(new_n8124_));
  XOR2X1   g07868(.A(new_n8124_), .B(\a[17] ), .Y(new_n8125_));
  INVX1    g07869(.A(new_n8125_), .Y(new_n8126_));
  XOR2X1   g07870(.A(new_n8126_), .B(new_n8121_), .Y(new_n8127_));
  XOR2X1   g07871(.A(new_n8127_), .B(new_n7964_), .Y(new_n8128_));
  AOI22X1  g07872(.A0(new_n818_), .A1(\b[53] ), .B0(new_n817_), .B1(\b[52] ), .Y(new_n8129_));
  OAI21X1  g07873(.A0(new_n816_), .A1(new_n5787_), .B0(new_n8129_), .Y(new_n8130_));
  AOI21X1  g07874(.A0(new_n5786_), .A1(new_n668_), .B0(new_n8130_), .Y(new_n8131_));
  XOR2X1   g07875(.A(new_n8131_), .B(\a[14] ), .Y(new_n8132_));
  XOR2X1   g07876(.A(new_n8132_), .B(new_n8128_), .Y(new_n8133_));
  AND2X1   g07877(.A(new_n7944_), .B(new_n7796_), .Y(new_n8134_));
  AOI21X1  g07878(.A0(new_n7945_), .A1(new_n7791_), .B0(new_n8134_), .Y(new_n8135_));
  XOR2X1   g07879(.A(new_n8135_), .B(new_n8133_), .Y(new_n8136_));
  AOI22X1  g07880(.A0(new_n603_), .A1(\b[56] ), .B0(new_n602_), .B1(\b[55] ), .Y(new_n8137_));
  OAI21X1  g07881(.A0(new_n601_), .A1(new_n6148_), .B0(new_n8137_), .Y(new_n8138_));
  AOI21X1  g07882(.A0(new_n6342_), .A1(new_n518_), .B0(new_n8138_), .Y(new_n8139_));
  XOR2X1   g07883(.A(new_n8139_), .B(\a[11] ), .Y(new_n8140_));
  XOR2X1   g07884(.A(new_n8140_), .B(new_n8136_), .Y(new_n8141_));
  AOI22X1  g07885(.A0(new_n469_), .A1(\b[59] ), .B0(new_n468_), .B1(\b[58] ), .Y(new_n8142_));
  OAI21X1  g07886(.A0(new_n467_), .A1(new_n6933_), .B0(new_n8142_), .Y(new_n8143_));
  AOI21X1  g07887(.A0(new_n6932_), .A1(new_n404_), .B0(new_n8143_), .Y(new_n8144_));
  XOR2X1   g07888(.A(new_n8144_), .B(\a[8] ), .Y(new_n8145_));
  XOR2X1   g07889(.A(new_n8145_), .B(new_n8141_), .Y(new_n8146_));
  INVX1    g07890(.A(new_n7789_), .Y(new_n8147_));
  AND2X1   g07891(.A(new_n7946_), .B(new_n8147_), .Y(new_n8148_));
  XOR2X1   g07892(.A(new_n7946_), .B(new_n8147_), .Y(new_n8149_));
  AOI21X1  g07893(.A0(new_n8149_), .A1(new_n7785_), .B0(new_n8148_), .Y(new_n8150_));
  XOR2X1   g07894(.A(new_n8150_), .B(new_n8146_), .Y(new_n8151_));
  AOI22X1  g07895(.A0(new_n369_), .A1(\b[62] ), .B0(new_n368_), .B1(\b[61] ), .Y(new_n8152_));
  OAI21X1  g07896(.A0(new_n367_), .A1(new_n7559_), .B0(new_n8152_), .Y(new_n8153_));
  AOI21X1  g07897(.A0(new_n7558_), .A1(new_n308_), .B0(new_n8153_), .Y(new_n8154_));
  XOR2X1   g07898(.A(new_n8154_), .B(\a[5] ), .Y(new_n8155_));
  XOR2X1   g07899(.A(new_n8155_), .B(new_n8151_), .Y(new_n8156_));
  OR2X1    g07900(.A(new_n7952_), .B(new_n7948_), .Y(new_n8157_));
  XOR2X1   g07901(.A(new_n8149_), .B(new_n7785_), .Y(new_n8158_));
  XOR2X1   g07902(.A(new_n7952_), .B(new_n8158_), .Y(new_n8159_));
  OAI21X1  g07903(.A0(new_n7957_), .A1(new_n8159_), .B0(new_n8157_), .Y(new_n8160_));
  AND2X1   g07904(.A(new_n7774_), .B(new_n318_), .Y(new_n8161_));
  AOI22X1  g07905(.A0(new_n7774_), .A1(new_n318_), .B0(new_n282_), .B1(\b[63] ), .Y(new_n8162_));
  MX2X1    g07906(.A(new_n8162_), .B(new_n8161_), .S0(new_n257_), .Y(new_n8163_));
  XOR2X1   g07907(.A(new_n8163_), .B(new_n8160_), .Y(new_n8164_));
  XOR2X1   g07908(.A(new_n8164_), .B(new_n8156_), .Y(new_n8165_));
  NOR2X1   g07909(.A(new_n7958_), .B(new_n7780_), .Y(new_n8166_));
  AOI21X1  g07910(.A0(new_n7959_), .A1(new_n7778_), .B0(new_n8166_), .Y(new_n8167_));
  XOR2X1   g07911(.A(new_n8167_), .B(new_n8165_), .Y(new_n8168_));
  OAI21X1  g07912(.A0(new_n7752_), .A1(new_n7769_), .B0(new_n7766_), .Y(new_n8169_));
  AND2X1   g07913(.A(new_n7960_), .B(new_n8169_), .Y(new_n8170_));
  AOI21X1  g07914(.A0(new_n7764_), .A1(new_n7763_), .B0(new_n7961_), .Y(new_n8171_));
  OR2X1    g07915(.A(new_n8171_), .B(new_n8170_), .Y(new_n8172_));
  XOR2X1   g07916(.A(new_n8172_), .B(new_n8168_), .Y(\f[65] ));
  OR2X1    g07917(.A(new_n8150_), .B(new_n8146_), .Y(new_n8174_));
  INVX1    g07918(.A(new_n8145_), .Y(new_n8175_));
  XOR2X1   g07919(.A(new_n8175_), .B(new_n8141_), .Y(new_n8176_));
  XOR2X1   g07920(.A(new_n8150_), .B(new_n8176_), .Y(new_n8177_));
  OAI21X1  g07921(.A0(new_n8155_), .A1(new_n8177_), .B0(new_n8174_), .Y(new_n8178_));
  AOI22X1  g07922(.A0(new_n369_), .A1(\b[63] ), .B0(new_n368_), .B1(\b[62] ), .Y(new_n8179_));
  OAI21X1  g07923(.A0(new_n367_), .A1(new_n7748_), .B0(new_n8179_), .Y(new_n8180_));
  AOI21X1  g07924(.A0(new_n7747_), .A1(new_n308_), .B0(new_n8180_), .Y(new_n8181_));
  XOR2X1   g07925(.A(new_n8181_), .B(\a[5] ), .Y(new_n8182_));
  XOR2X1   g07926(.A(new_n8182_), .B(new_n8178_), .Y(new_n8183_));
  AOI22X1  g07927(.A0(new_n603_), .A1(\b[57] ), .B0(new_n602_), .B1(\b[56] ), .Y(new_n8184_));
  OAI21X1  g07928(.A0(new_n601_), .A1(new_n6523_), .B0(new_n8184_), .Y(new_n8185_));
  AOI21X1  g07929(.A0(new_n6522_), .A1(new_n518_), .B0(new_n8185_), .Y(new_n8186_));
  XOR2X1   g07930(.A(new_n8186_), .B(\a[11] ), .Y(new_n8187_));
  INVX1    g07931(.A(new_n8187_), .Y(new_n8188_));
  NOR2X1   g07932(.A(new_n8132_), .B(new_n8128_), .Y(new_n8189_));
  AND2X1   g07933(.A(new_n7945_), .B(new_n7791_), .Y(new_n8190_));
  OR2X1    g07934(.A(new_n8190_), .B(new_n8134_), .Y(new_n8191_));
  AOI21X1  g07935(.A0(new_n8191_), .A1(new_n8133_), .B0(new_n8189_), .Y(new_n8192_));
  XOR2X1   g07936(.A(new_n8192_), .B(new_n8188_), .Y(new_n8193_));
  AOI22X1  g07937(.A0(new_n1017_), .A1(\b[51] ), .B0(new_n1016_), .B1(\b[50] ), .Y(new_n8194_));
  OAI21X1  g07938(.A0(new_n1015_), .A1(new_n5237_), .B0(new_n8194_), .Y(new_n8195_));
  AOI21X1  g07939(.A0(new_n5236_), .A1(new_n882_), .B0(new_n8195_), .Y(new_n8196_));
  XOR2X1   g07940(.A(new_n8196_), .B(\a[17] ), .Y(new_n8197_));
  INVX1    g07941(.A(new_n8197_), .Y(new_n8198_));
  INVX1    g07942(.A(new_n7971_), .Y(new_n8199_));
  NOR2X1   g07943(.A(new_n8120_), .B(new_n7967_), .Y(new_n8200_));
  AOI21X1  g07944(.A0(new_n8119_), .A1(new_n8199_), .B0(new_n8200_), .Y(new_n8201_));
  XOR2X1   g07945(.A(new_n8201_), .B(new_n8198_), .Y(new_n8202_));
  AOI22X1  g07946(.A0(new_n1263_), .A1(\b[48] ), .B0(new_n1262_), .B1(\b[47] ), .Y(new_n8203_));
  OAI21X1  g07947(.A0(new_n1261_), .A1(new_n4693_), .B0(new_n8203_), .Y(new_n8204_));
  AOI21X1  g07948(.A0(new_n4692_), .A1(new_n1075_), .B0(new_n8204_), .Y(new_n8205_));
  XOR2X1   g07949(.A(new_n8205_), .B(\a[20] ), .Y(new_n8206_));
  OR2X1    g07950(.A(new_n8114_), .B(new_n8110_), .Y(new_n8207_));
  OAI21X1  g07951(.A0(new_n8118_), .A1(new_n8116_), .B0(new_n8207_), .Y(new_n8208_));
  XOR2X1   g07952(.A(new_n8208_), .B(new_n8206_), .Y(new_n8209_));
  AOI22X1  g07953(.A0(new_n1526_), .A1(\b[45] ), .B0(new_n1525_), .B1(\b[44] ), .Y(new_n8210_));
  OAI21X1  g07954(.A0(new_n1524_), .A1(new_n4339_), .B0(new_n8210_), .Y(new_n8211_));
  AOI21X1  g07955(.A0(new_n4338_), .A1(new_n1347_), .B0(new_n8211_), .Y(new_n8212_));
  XOR2X1   g07956(.A(new_n8212_), .B(\a[23] ), .Y(new_n8213_));
  XOR2X1   g07957(.A(new_n8213_), .B(new_n8109_), .Y(new_n8214_));
  INVX1    g07958(.A(new_n8214_), .Y(new_n8215_));
  AOI22X1  g07959(.A0(new_n1814_), .A1(\b[42] ), .B0(new_n1813_), .B1(\b[41] ), .Y(new_n8216_));
  OAI21X1  g07960(.A0(new_n1812_), .A1(new_n3720_), .B0(new_n8216_), .Y(new_n8217_));
  AOI21X1  g07961(.A0(new_n3860_), .A1(new_n1617_), .B0(new_n8217_), .Y(new_n8218_));
  XOR2X1   g07962(.A(new_n8218_), .B(\a[26] ), .Y(new_n8219_));
  INVX1    g07963(.A(new_n8219_), .Y(new_n8220_));
  INVX1    g07964(.A(new_n8087_), .Y(new_n8221_));
  AND2X1   g07965(.A(new_n8221_), .B(new_n8083_), .Y(new_n8222_));
  XOR2X1   g07966(.A(new_n8221_), .B(new_n8083_), .Y(new_n8223_));
  AOI21X1  g07967(.A0(new_n8092_), .A1(new_n8223_), .B0(new_n8222_), .Y(new_n8224_));
  XOR2X1   g07968(.A(new_n8224_), .B(new_n8220_), .Y(new_n8225_));
  XOR2X1   g07969(.A(new_n8077_), .B(new_n2258_), .Y(new_n8226_));
  AND2X1   g07970(.A(new_n8226_), .B(new_n8074_), .Y(new_n8227_));
  INVX1    g07971(.A(new_n8227_), .Y(new_n8228_));
  OR2X1    g07972(.A(new_n8082_), .B(new_n8079_), .Y(new_n8229_));
  NAND2X1  g07973(.A(new_n8229_), .B(new_n8228_), .Y(new_n8230_));
  AOI22X1  g07974(.A0(new_n2163_), .A1(\b[39] ), .B0(new_n2162_), .B1(\b[38] ), .Y(new_n8231_));
  OAI21X1  g07975(.A0(new_n2161_), .A1(new_n3413_), .B0(new_n8231_), .Y(new_n8232_));
  AOI21X1  g07976(.A0(new_n3412_), .A1(new_n1907_), .B0(new_n8232_), .Y(new_n8233_));
  XOR2X1   g07977(.A(new_n8233_), .B(\a[29] ), .Y(new_n8234_));
  XOR2X1   g07978(.A(new_n8234_), .B(new_n8230_), .Y(new_n8235_));
  NOR2X1   g07979(.A(new_n8019_), .B(new_n8015_), .Y(new_n8236_));
  AOI21X1  g07980(.A0(new_n8020_), .A1(new_n7989_), .B0(new_n8236_), .Y(new_n8237_));
  INVX1    g07981(.A(new_n8237_), .Y(new_n8238_));
  NOR2X1   g07982(.A(new_n7997_), .B(new_n7993_), .Y(new_n8239_));
  AOI21X1  g07983(.A0(new_n8002_), .A1(new_n8000_), .B0(new_n7999_), .Y(new_n8240_));
  NOR2X1   g07984(.A(new_n8240_), .B(new_n8239_), .Y(new_n8241_));
  AOI22X1  g07985(.A0(new_n7818_), .A1(\b[2] ), .B0(new_n7817_), .B1(\b[3] ), .Y(new_n8242_));
  XOR2X1   g07986(.A(new_n8242_), .B(\a[2] ), .Y(new_n8243_));
  AOI22X1  g07987(.A0(new_n7192_), .A1(\b[6] ), .B0(new_n7189_), .B1(\b[5] ), .Y(new_n8244_));
  OAI21X1  g07988(.A0(new_n7627_), .A1(new_n325_), .B0(new_n8244_), .Y(new_n8245_));
  AOI21X1  g07989(.A0(new_n7187_), .A1(new_n378_), .B0(new_n8245_), .Y(new_n8246_));
  XOR2X1   g07990(.A(new_n8246_), .B(\a[62] ), .Y(new_n8247_));
  XOR2X1   g07991(.A(new_n8247_), .B(new_n8243_), .Y(new_n8248_));
  XOR2X1   g07992(.A(new_n8248_), .B(new_n8241_), .Y(new_n8249_));
  AOI22X1  g07993(.A0(new_n6603_), .A1(\b[9] ), .B0(new_n6600_), .B1(\b[8] ), .Y(new_n8250_));
  OAI21X1  g07994(.A0(new_n6804_), .A1(new_n492_), .B0(new_n8250_), .Y(new_n8251_));
  AOI21X1  g07995(.A0(new_n6598_), .A1(new_n491_), .B0(new_n8251_), .Y(new_n8252_));
  XOR2X1   g07996(.A(new_n8252_), .B(\a[59] ), .Y(new_n8253_));
  XOR2X1   g07997(.A(new_n8253_), .B(new_n8249_), .Y(new_n8254_));
  XOR2X1   g07998(.A(new_n8254_), .B(new_n8014_), .Y(new_n8255_));
  AOI22X1  g07999(.A0(new_n6438_), .A1(\b[12] ), .B0(new_n6437_), .B1(\b[11] ), .Y(new_n8256_));
  OAI21X1  g08000(.A0(new_n6436_), .A1(new_n587_), .B0(new_n8256_), .Y(new_n8257_));
  AOI21X1  g08001(.A0(new_n6023_), .A1(new_n635_), .B0(new_n8257_), .Y(new_n8258_));
  XOR2X1   g08002(.A(new_n8258_), .B(\a[56] ), .Y(new_n8259_));
  XOR2X1   g08003(.A(new_n8259_), .B(new_n8255_), .Y(new_n8260_));
  XOR2X1   g08004(.A(new_n8260_), .B(new_n8238_), .Y(new_n8261_));
  AOI22X1  g08005(.A0(new_n5430_), .A1(\b[15] ), .B0(new_n5427_), .B1(\b[14] ), .Y(new_n8262_));
  OAI21X1  g08006(.A0(new_n5891_), .A1(new_n795_), .B0(new_n8262_), .Y(new_n8263_));
  AOI21X1  g08007(.A0(new_n5425_), .A1(new_n794_), .B0(new_n8263_), .Y(new_n8264_));
  XOR2X1   g08008(.A(new_n8264_), .B(\a[53] ), .Y(new_n8265_));
  XOR2X1   g08009(.A(new_n8265_), .B(new_n8261_), .Y(new_n8266_));
  XOR2X1   g08010(.A(new_n8024_), .B(new_n5423_), .Y(new_n8267_));
  AND2X1   g08011(.A(new_n8267_), .B(new_n8021_), .Y(new_n8268_));
  INVX1    g08012(.A(new_n8026_), .Y(new_n8269_));
  AOI21X1  g08013(.A0(new_n8269_), .A1(new_n7985_), .B0(new_n8268_), .Y(new_n8270_));
  XOR2X1   g08014(.A(new_n8270_), .B(new_n8266_), .Y(new_n8271_));
  AOI22X1  g08015(.A0(new_n4880_), .A1(\b[18] ), .B0(new_n4877_), .B1(\b[17] ), .Y(new_n8272_));
  OAI21X1  g08016(.A0(new_n5291_), .A1(new_n974_), .B0(new_n8272_), .Y(new_n8273_));
  AOI21X1  g08017(.A0(new_n4875_), .A1(new_n1042_), .B0(new_n8273_), .Y(new_n8274_));
  XOR2X1   g08018(.A(new_n8274_), .B(\a[50] ), .Y(new_n8275_));
  XOR2X1   g08019(.A(new_n8275_), .B(new_n8271_), .Y(new_n8276_));
  NOR2X1   g08020(.A(new_n8031_), .B(new_n8027_), .Y(new_n8277_));
  AOI21X1  g08021(.A0(new_n8032_), .A1(new_n7983_), .B0(new_n8277_), .Y(new_n8278_));
  XOR2X1   g08022(.A(new_n8278_), .B(new_n8276_), .Y(new_n8279_));
  AOI22X1  g08023(.A0(new_n4572_), .A1(\b[21] ), .B0(new_n4571_), .B1(\b[20] ), .Y(new_n8280_));
  OAI21X1  g08024(.A0(new_n4740_), .A1(new_n1300_), .B0(new_n8280_), .Y(new_n8281_));
  AOI21X1  g08025(.A0(new_n4375_), .A1(new_n1299_), .B0(new_n8281_), .Y(new_n8282_));
  XOR2X1   g08026(.A(new_n8282_), .B(\a[47] ), .Y(new_n8283_));
  INVX1    g08027(.A(new_n8283_), .Y(new_n8284_));
  XOR2X1   g08028(.A(new_n8284_), .B(new_n8279_), .Y(new_n8285_));
  INVX1    g08029(.A(new_n8285_), .Y(new_n8286_));
  XOR2X1   g08030(.A(new_n8036_), .B(new_n4568_), .Y(new_n8287_));
  AND2X1   g08031(.A(new_n8287_), .B(new_n8033_), .Y(new_n8288_));
  INVX1    g08032(.A(new_n8038_), .Y(new_n8289_));
  AOI21X1  g08033(.A0(new_n8289_), .A1(new_n7979_), .B0(new_n8288_), .Y(new_n8290_));
  XOR2X1   g08034(.A(new_n8290_), .B(new_n8286_), .Y(new_n8291_));
  AOI22X1  g08035(.A0(new_n4095_), .A1(\b[24] ), .B0(new_n4094_), .B1(\b[23] ), .Y(new_n8292_));
  OAI21X1  g08036(.A0(new_n4233_), .A1(new_n1479_), .B0(new_n8292_), .Y(new_n8293_));
  AOI21X1  g08037(.A0(new_n3901_), .A1(new_n1572_), .B0(new_n8293_), .Y(new_n8294_));
  XOR2X1   g08038(.A(new_n8294_), .B(\a[44] ), .Y(new_n8295_));
  XOR2X1   g08039(.A(new_n8295_), .B(new_n8291_), .Y(new_n8296_));
  NOR2X1   g08040(.A(new_n8043_), .B(new_n8039_), .Y(new_n8297_));
  AOI21X1  g08041(.A0(new_n8044_), .A1(new_n7976_), .B0(new_n8297_), .Y(new_n8298_));
  XOR2X1   g08042(.A(new_n8298_), .B(new_n8296_), .Y(new_n8299_));
  AOI22X1  g08043(.A0(new_n3652_), .A1(\b[27] ), .B0(new_n3651_), .B1(\b[26] ), .Y(new_n8300_));
  OAI21X1  g08044(.A0(new_n3778_), .A1(new_n1880_), .B0(new_n8300_), .Y(new_n8301_));
  AOI21X1  g08045(.A0(new_n3480_), .A1(new_n1879_), .B0(new_n8301_), .Y(new_n8302_));
  XOR2X1   g08046(.A(new_n8302_), .B(\a[41] ), .Y(new_n8303_));
  XOR2X1   g08047(.A(new_n8303_), .B(new_n8299_), .Y(new_n8304_));
  INVX1    g08048(.A(new_n8304_), .Y(new_n8305_));
  INVX1    g08049(.A(new_n8051_), .Y(new_n8306_));
  NOR2X1   g08050(.A(new_n8053_), .B(new_n8306_), .Y(new_n8307_));
  AOI21X1  g08051(.A0(new_n8050_), .A1(new_n8045_), .B0(new_n8307_), .Y(new_n8308_));
  XOR2X1   g08052(.A(new_n8308_), .B(new_n8305_), .Y(new_n8309_));
  AOI22X1  g08053(.A0(new_n3204_), .A1(\b[30] ), .B0(new_n3203_), .B1(\b[29] ), .Y(new_n8310_));
  OAI21X1  g08054(.A0(new_n3321_), .A1(new_n2231_), .B0(new_n8310_), .Y(new_n8311_));
  AOI21X1  g08055(.A0(new_n3080_), .A1(new_n2230_), .B0(new_n8311_), .Y(new_n8312_));
  XOR2X1   g08056(.A(new_n8312_), .B(\a[38] ), .Y(new_n8313_));
  XOR2X1   g08057(.A(new_n8313_), .B(new_n8309_), .Y(new_n8314_));
  NOR2X1   g08058(.A(new_n8058_), .B(new_n8054_), .Y(new_n8315_));
  INVX1    g08059(.A(new_n8064_), .Y(new_n8316_));
  AOI21X1  g08060(.A0(new_n8316_), .A1(new_n8059_), .B0(new_n8315_), .Y(new_n8317_));
  XOR2X1   g08061(.A(new_n8317_), .B(new_n8314_), .Y(new_n8318_));
  AOI22X1  g08062(.A0(new_n2813_), .A1(\b[33] ), .B0(new_n2812_), .B1(\b[32] ), .Y(new_n8319_));
  OAI21X1  g08063(.A0(new_n2946_), .A1(new_n2615_), .B0(new_n8319_), .Y(new_n8320_));
  AOI21X1  g08064(.A0(new_n2652_), .A1(new_n2614_), .B0(new_n8320_), .Y(new_n8321_));
  XOR2X1   g08065(.A(new_n8321_), .B(\a[35] ), .Y(new_n8322_));
  XOR2X1   g08066(.A(new_n8322_), .B(new_n8318_), .Y(new_n8323_));
  INVX1    g08067(.A(new_n8323_), .Y(new_n8324_));
  AOI22X1  g08068(.A0(new_n2545_), .A1(\b[36] ), .B0(new_n2544_), .B1(\b[35] ), .Y(new_n8325_));
  OAI21X1  g08069(.A0(new_n2543_), .A1(new_n2890_), .B0(new_n8325_), .Y(new_n8326_));
  AOI21X1  g08070(.A0(new_n3015_), .A1(new_n2260_), .B0(new_n8326_), .Y(new_n8327_));
  XOR2X1   g08071(.A(new_n8327_), .B(\a[32] ), .Y(new_n8328_));
  XOR2X1   g08072(.A(new_n8328_), .B(new_n8073_), .Y(new_n8329_));
  XOR2X1   g08073(.A(new_n8329_), .B(new_n8324_), .Y(new_n8330_));
  XOR2X1   g08074(.A(new_n8330_), .B(new_n8235_), .Y(new_n8331_));
  XOR2X1   g08075(.A(new_n8331_), .B(new_n8225_), .Y(new_n8332_));
  XOR2X1   g08076(.A(new_n8332_), .B(new_n8215_), .Y(new_n8333_));
  XOR2X1   g08077(.A(new_n8333_), .B(new_n8209_), .Y(new_n8334_));
  XOR2X1   g08078(.A(new_n8334_), .B(new_n8202_), .Y(new_n8335_));
  NAND2X1  g08079(.A(new_n8126_), .B(new_n8121_), .Y(new_n8336_));
  XOR2X1   g08080(.A(new_n8125_), .B(new_n8121_), .Y(new_n8337_));
  OAI21X1  g08081(.A0(new_n8337_), .A1(new_n7964_), .B0(new_n8336_), .Y(new_n8338_));
  AOI22X1  g08082(.A0(new_n818_), .A1(\b[54] ), .B0(new_n817_), .B1(\b[53] ), .Y(new_n8339_));
  OAI21X1  g08083(.A0(new_n816_), .A1(new_n5808_), .B0(new_n8339_), .Y(new_n8340_));
  AOI21X1  g08084(.A0(new_n5807_), .A1(new_n668_), .B0(new_n8340_), .Y(new_n8341_));
  XOR2X1   g08085(.A(new_n8341_), .B(new_n665_), .Y(new_n8342_));
  XOR2X1   g08086(.A(new_n8342_), .B(new_n8338_), .Y(new_n8343_));
  XOR2X1   g08087(.A(new_n8343_), .B(new_n8335_), .Y(new_n8344_));
  XOR2X1   g08088(.A(new_n8344_), .B(new_n8193_), .Y(new_n8345_));
  AOI22X1  g08089(.A0(new_n469_), .A1(\b[60] ), .B0(new_n468_), .B1(\b[59] ), .Y(new_n8346_));
  OAI21X1  g08090(.A0(new_n467_), .A1(new_n6930_), .B0(new_n8346_), .Y(new_n8347_));
  AOI21X1  g08091(.A0(new_n6951_), .A1(new_n404_), .B0(new_n8347_), .Y(new_n8348_));
  XOR2X1   g08092(.A(new_n8348_), .B(\a[8] ), .Y(new_n8349_));
  INVX1    g08093(.A(new_n8349_), .Y(new_n8350_));
  NOR2X1   g08094(.A(new_n8140_), .B(new_n8136_), .Y(new_n8351_));
  AOI21X1  g08095(.A0(new_n8175_), .A1(new_n8141_), .B0(new_n8351_), .Y(new_n8352_));
  XOR2X1   g08096(.A(new_n8352_), .B(new_n8350_), .Y(new_n8353_));
  XOR2X1   g08097(.A(new_n8353_), .B(new_n8345_), .Y(new_n8354_));
  XOR2X1   g08098(.A(new_n8354_), .B(new_n8183_), .Y(new_n8355_));
  XOR2X1   g08099(.A(new_n8155_), .B(new_n8177_), .Y(new_n8356_));
  AND2X1   g08100(.A(new_n8163_), .B(new_n8160_), .Y(new_n8357_));
  AOI21X1  g08101(.A0(new_n8164_), .A1(new_n8356_), .B0(new_n8357_), .Y(new_n8358_));
  XOR2X1   g08102(.A(new_n8358_), .B(new_n8355_), .Y(new_n8359_));
  OR2X1    g08103(.A(new_n8167_), .B(new_n8165_), .Y(new_n8360_));
  OAI21X1  g08104(.A0(new_n8171_), .A1(new_n8170_), .B0(new_n8168_), .Y(new_n8361_));
  AND2X1   g08105(.A(new_n8361_), .B(new_n8360_), .Y(new_n8362_));
  XOR2X1   g08106(.A(new_n8362_), .B(new_n8359_), .Y(\f[66] ));
  INVX1    g08107(.A(new_n8354_), .Y(new_n8364_));
  XOR2X1   g08108(.A(new_n8364_), .B(new_n8183_), .Y(new_n8365_));
  NOR2X1   g08109(.A(new_n8358_), .B(new_n8365_), .Y(new_n8366_));
  AOI21X1  g08110(.A0(new_n8361_), .A1(new_n8360_), .B0(new_n8359_), .Y(new_n8367_));
  OR2X1    g08111(.A(new_n8367_), .B(new_n8366_), .Y(new_n8368_));
  OR2X1    g08112(.A(new_n8155_), .B(new_n8177_), .Y(new_n8369_));
  AOI21X1  g08113(.A0(new_n8369_), .A1(new_n8174_), .B0(new_n8182_), .Y(new_n8370_));
  NOR2X1   g08114(.A(new_n8354_), .B(new_n8183_), .Y(new_n8371_));
  OR2X1    g08115(.A(new_n8371_), .B(new_n8370_), .Y(new_n8372_));
  AOI22X1  g08116(.A0(new_n818_), .A1(\b[55] ), .B0(new_n817_), .B1(\b[54] ), .Y(new_n8373_));
  OAI21X1  g08117(.A0(new_n816_), .A1(new_n6151_), .B0(new_n8373_), .Y(new_n8374_));
  AOI21X1  g08118(.A0(new_n6150_), .A1(new_n668_), .B0(new_n8374_), .Y(new_n8375_));
  XOR2X1   g08119(.A(new_n8375_), .B(\a[14] ), .Y(new_n8376_));
  INVX1    g08120(.A(new_n8376_), .Y(new_n8377_));
  NAND2X1  g08121(.A(new_n8201_), .B(new_n8197_), .Y(new_n8378_));
  NOR2X1   g08122(.A(new_n8201_), .B(new_n8197_), .Y(new_n8379_));
  AOI21X1  g08123(.A0(new_n8334_), .A1(new_n8378_), .B0(new_n8379_), .Y(new_n8380_));
  XOR2X1   g08124(.A(new_n8380_), .B(new_n8377_), .Y(new_n8381_));
  AOI22X1  g08125(.A0(new_n1263_), .A1(\b[49] ), .B0(new_n1262_), .B1(\b[48] ), .Y(new_n8382_));
  OAI21X1  g08126(.A0(new_n1261_), .A1(new_n5039_), .B0(new_n8382_), .Y(new_n8383_));
  AOI21X1  g08127(.A0(new_n5038_), .A1(new_n1075_), .B0(new_n8383_), .Y(new_n8384_));
  XOR2X1   g08128(.A(new_n8384_), .B(\a[20] ), .Y(new_n8385_));
  INVX1    g08129(.A(new_n8385_), .Y(new_n8386_));
  NOR2X1   g08130(.A(new_n8213_), .B(new_n8109_), .Y(new_n8387_));
  AOI21X1  g08131(.A0(new_n8332_), .A1(new_n8214_), .B0(new_n8387_), .Y(new_n8388_));
  XOR2X1   g08132(.A(new_n8388_), .B(new_n8386_), .Y(new_n8389_));
  AOI22X1  g08133(.A0(new_n1814_), .A1(\b[43] ), .B0(new_n1813_), .B1(\b[42] ), .Y(new_n8390_));
  OAI21X1  g08134(.A0(new_n1812_), .A1(new_n4015_), .B0(new_n8390_), .Y(new_n8391_));
  AOI21X1  g08135(.A0(new_n4014_), .A1(new_n1617_), .B0(new_n8391_), .Y(new_n8392_));
  XOR2X1   g08136(.A(new_n8392_), .B(\a[26] ), .Y(new_n8393_));
  INVX1    g08137(.A(new_n8393_), .Y(new_n8394_));
  AOI21X1  g08138(.A0(new_n8229_), .A1(new_n8228_), .B0(new_n8234_), .Y(new_n8395_));
  NAND3X1  g08139(.A(new_n8234_), .B(new_n8229_), .C(new_n8228_), .Y(new_n8396_));
  AOI21X1  g08140(.A0(new_n8330_), .A1(new_n8396_), .B0(new_n8395_), .Y(new_n8397_));
  XOR2X1   g08141(.A(new_n8397_), .B(new_n8394_), .Y(new_n8398_));
  AND2X1   g08142(.A(new_n8313_), .B(new_n8309_), .Y(new_n8399_));
  NOR2X1   g08143(.A(new_n8313_), .B(new_n8309_), .Y(new_n8400_));
  NOR3X1   g08144(.A(new_n8317_), .B(new_n8400_), .C(new_n8399_), .Y(new_n8401_));
  NOR2X1   g08145(.A(new_n8322_), .B(new_n8318_), .Y(new_n8402_));
  OR2X1    g08146(.A(new_n8402_), .B(new_n8401_), .Y(new_n8403_));
  AOI22X1  g08147(.A0(new_n2545_), .A1(\b[37] ), .B0(new_n2544_), .B1(\b[36] ), .Y(new_n8404_));
  OAI21X1  g08148(.A0(new_n2543_), .A1(new_n3156_), .B0(new_n8404_), .Y(new_n8405_));
  AOI21X1  g08149(.A0(new_n3155_), .A1(new_n2260_), .B0(new_n8405_), .Y(new_n8406_));
  XOR2X1   g08150(.A(new_n8406_), .B(\a[32] ), .Y(new_n8407_));
  XOR2X1   g08151(.A(new_n8407_), .B(new_n8403_), .Y(new_n8408_));
  AOI22X1  g08152(.A0(new_n2813_), .A1(\b[34] ), .B0(new_n2812_), .B1(\b[33] ), .Y(new_n8409_));
  OAI21X1  g08153(.A0(new_n2946_), .A1(new_n2612_), .B0(new_n8409_), .Y(new_n8410_));
  AOI21X1  g08154(.A0(new_n2759_), .A1(new_n2652_), .B0(new_n8410_), .Y(new_n8411_));
  XOR2X1   g08155(.A(new_n8411_), .B(\a[35] ), .Y(new_n8412_));
  INVX1    g08156(.A(new_n8412_), .Y(new_n8413_));
  NOR2X1   g08157(.A(new_n8308_), .B(new_n8304_), .Y(new_n8414_));
  NOR2X1   g08158(.A(new_n8400_), .B(new_n8414_), .Y(new_n8415_));
  AOI22X1  g08159(.A0(new_n7192_), .A1(\b[7] ), .B0(new_n7189_), .B1(\b[6] ), .Y(new_n8416_));
  OAI21X1  g08160(.A0(new_n7627_), .A1(new_n395_), .B0(new_n8416_), .Y(new_n8417_));
  AOI21X1  g08161(.A0(new_n7187_), .A1(new_n394_), .B0(new_n8417_), .Y(new_n8418_));
  XOR2X1   g08162(.A(new_n8418_), .B(new_n7185_), .Y(new_n8419_));
  AOI22X1  g08163(.A0(new_n7818_), .A1(\b[3] ), .B0(new_n7817_), .B1(\b[4] ), .Y(new_n8420_));
  XOR2X1   g08164(.A(new_n8420_), .B(\a[2] ), .Y(new_n8421_));
  XOR2X1   g08165(.A(new_n8421_), .B(new_n8419_), .Y(new_n8422_));
  OR2X1    g08166(.A(new_n8242_), .B(new_n257_), .Y(new_n8423_));
  OR2X1    g08167(.A(new_n8247_), .B(new_n8243_), .Y(new_n8424_));
  AND2X1   g08168(.A(new_n8424_), .B(new_n8423_), .Y(new_n8425_));
  XOR2X1   g08169(.A(new_n8425_), .B(new_n8422_), .Y(new_n8426_));
  AOI22X1  g08170(.A0(new_n6603_), .A1(\b[10] ), .B0(new_n6600_), .B1(\b[9] ), .Y(new_n8427_));
  OAI21X1  g08171(.A0(new_n6804_), .A1(new_n489_), .B0(new_n8427_), .Y(new_n8428_));
  AOI21X1  g08172(.A0(new_n6598_), .A1(new_n543_), .B0(new_n8428_), .Y(new_n8429_));
  XOR2X1   g08173(.A(new_n8429_), .B(\a[59] ), .Y(new_n8430_));
  XOR2X1   g08174(.A(new_n8430_), .B(new_n8426_), .Y(new_n8431_));
  OAI21X1  g08175(.A0(new_n8240_), .A1(new_n8239_), .B0(new_n8248_), .Y(new_n8432_));
  OR2X1    g08176(.A(new_n8253_), .B(new_n8249_), .Y(new_n8433_));
  AND2X1   g08177(.A(new_n8433_), .B(new_n8432_), .Y(new_n8434_));
  XOR2X1   g08178(.A(new_n8434_), .B(new_n8431_), .Y(new_n8435_));
  AOI22X1  g08179(.A0(new_n6438_), .A1(\b[13] ), .B0(new_n6437_), .B1(\b[12] ), .Y(new_n8436_));
  OAI21X1  g08180(.A0(new_n6436_), .A1(new_n716_), .B0(new_n8436_), .Y(new_n8437_));
  AOI21X1  g08181(.A0(new_n6023_), .A1(new_n715_), .B0(new_n8437_), .Y(new_n8438_));
  XOR2X1   g08182(.A(new_n8438_), .B(\a[56] ), .Y(new_n8439_));
  INVX1    g08183(.A(new_n8439_), .Y(new_n8440_));
  XOR2X1   g08184(.A(new_n8440_), .B(new_n8435_), .Y(new_n8441_));
  INVX1    g08185(.A(new_n8441_), .Y(new_n8442_));
  INVX1    g08186(.A(new_n8014_), .Y(new_n8443_));
  NOR2X1   g08187(.A(new_n8259_), .B(new_n8255_), .Y(new_n8444_));
  AOI21X1  g08188(.A0(new_n8254_), .A1(new_n8443_), .B0(new_n8444_), .Y(new_n8445_));
  XOR2X1   g08189(.A(new_n8445_), .B(new_n8442_), .Y(new_n8446_));
  AOI22X1  g08190(.A0(new_n5430_), .A1(\b[16] ), .B0(new_n5427_), .B1(\b[15] ), .Y(new_n8447_));
  OAI21X1  g08191(.A0(new_n5891_), .A1(new_n792_), .B0(new_n8447_), .Y(new_n8448_));
  AOI21X1  g08192(.A0(new_n5425_), .A1(new_n842_), .B0(new_n8448_), .Y(new_n8449_));
  XOR2X1   g08193(.A(new_n8449_), .B(\a[53] ), .Y(new_n8450_));
  XOR2X1   g08194(.A(new_n8450_), .B(new_n8446_), .Y(new_n8451_));
  AND2X1   g08195(.A(new_n8260_), .B(new_n8238_), .Y(new_n8452_));
  INVX1    g08196(.A(new_n8265_), .Y(new_n8453_));
  AOI21X1  g08197(.A0(new_n8453_), .A1(new_n8261_), .B0(new_n8452_), .Y(new_n8454_));
  XOR2X1   g08198(.A(new_n8454_), .B(new_n8451_), .Y(new_n8455_));
  AOI22X1  g08199(.A0(new_n4880_), .A1(\b[19] ), .B0(new_n4877_), .B1(\b[18] ), .Y(new_n8456_));
  OAI21X1  g08200(.A0(new_n5291_), .A1(new_n1118_), .B0(new_n8456_), .Y(new_n8457_));
  AOI21X1  g08201(.A0(new_n4875_), .A1(new_n1117_), .B0(new_n8457_), .Y(new_n8458_));
  XOR2X1   g08202(.A(new_n8458_), .B(\a[50] ), .Y(new_n8459_));
  XOR2X1   g08203(.A(new_n8459_), .B(new_n8455_), .Y(new_n8460_));
  NOR2X1   g08204(.A(new_n8270_), .B(new_n8266_), .Y(new_n8461_));
  INVX1    g08205(.A(new_n8275_), .Y(new_n8462_));
  AOI21X1  g08206(.A0(new_n8462_), .A1(new_n8271_), .B0(new_n8461_), .Y(new_n8463_));
  XOR2X1   g08207(.A(new_n8463_), .B(new_n8460_), .Y(new_n8464_));
  AOI22X1  g08208(.A0(new_n4572_), .A1(\b[22] ), .B0(new_n4571_), .B1(\b[21] ), .Y(new_n8465_));
  OAI21X1  g08209(.A0(new_n4740_), .A1(new_n1297_), .B0(new_n8465_), .Y(new_n8466_));
  AOI21X1  g08210(.A0(new_n4375_), .A1(new_n1399_), .B0(new_n8466_), .Y(new_n8467_));
  XOR2X1   g08211(.A(new_n8467_), .B(\a[47] ), .Y(new_n8468_));
  XOR2X1   g08212(.A(new_n8468_), .B(new_n8464_), .Y(new_n8469_));
  NOR2X1   g08213(.A(new_n8278_), .B(new_n8276_), .Y(new_n8470_));
  AOI21X1  g08214(.A0(new_n8284_), .A1(new_n8279_), .B0(new_n8470_), .Y(new_n8471_));
  XOR2X1   g08215(.A(new_n8471_), .B(new_n8469_), .Y(new_n8472_));
  AOI22X1  g08216(.A0(new_n4095_), .A1(\b[25] ), .B0(new_n4094_), .B1(\b[24] ), .Y(new_n8473_));
  OAI21X1  g08217(.A0(new_n4233_), .A1(new_n1591_), .B0(new_n8473_), .Y(new_n8474_));
  AOI21X1  g08218(.A0(new_n3901_), .A1(new_n1590_), .B0(new_n8474_), .Y(new_n8475_));
  XOR2X1   g08219(.A(new_n8475_), .B(\a[44] ), .Y(new_n8476_));
  XOR2X1   g08220(.A(new_n8476_), .B(new_n8472_), .Y(new_n8477_));
  NOR2X1   g08221(.A(new_n8290_), .B(new_n8286_), .Y(new_n8478_));
  INVX1    g08222(.A(new_n8295_), .Y(new_n8479_));
  AOI21X1  g08223(.A0(new_n8479_), .A1(new_n8291_), .B0(new_n8478_), .Y(new_n8480_));
  XOR2X1   g08224(.A(new_n8480_), .B(new_n8477_), .Y(new_n8481_));
  AOI22X1  g08225(.A0(new_n3652_), .A1(\b[28] ), .B0(new_n3651_), .B1(\b[27] ), .Y(new_n8482_));
  OAI21X1  g08226(.A0(new_n3778_), .A1(new_n1877_), .B0(new_n8482_), .Y(new_n8483_));
  AOI21X1  g08227(.A0(new_n3480_), .A1(new_n2004_), .B0(new_n8483_), .Y(new_n8484_));
  XOR2X1   g08228(.A(new_n8484_), .B(\a[41] ), .Y(new_n8485_));
  XOR2X1   g08229(.A(new_n8485_), .B(new_n8481_), .Y(new_n8486_));
  INVX1    g08230(.A(new_n8486_), .Y(new_n8487_));
  NOR2X1   g08231(.A(new_n8298_), .B(new_n8296_), .Y(new_n8488_));
  INVX1    g08232(.A(new_n8303_), .Y(new_n8489_));
  AOI21X1  g08233(.A0(new_n8489_), .A1(new_n8299_), .B0(new_n8488_), .Y(new_n8490_));
  XOR2X1   g08234(.A(new_n8490_), .B(new_n8487_), .Y(new_n8491_));
  AOI22X1  g08235(.A0(new_n3204_), .A1(\b[31] ), .B0(new_n3203_), .B1(\b[30] ), .Y(new_n8492_));
  OAI21X1  g08236(.A0(new_n3321_), .A1(new_n2359_), .B0(new_n8492_), .Y(new_n8493_));
  AOI21X1  g08237(.A0(new_n3080_), .A1(new_n2358_), .B0(new_n8493_), .Y(new_n8494_));
  XOR2X1   g08238(.A(new_n8494_), .B(\a[38] ), .Y(new_n8495_));
  XOR2X1   g08239(.A(new_n8495_), .B(new_n8491_), .Y(new_n8496_));
  XOR2X1   g08240(.A(new_n8496_), .B(new_n8415_), .Y(new_n8497_));
  XOR2X1   g08241(.A(new_n8497_), .B(new_n8413_), .Y(new_n8498_));
  XOR2X1   g08242(.A(new_n8498_), .B(new_n8408_), .Y(new_n8499_));
  INVX1    g08243(.A(new_n8499_), .Y(new_n8500_));
  AND2X1   g08244(.A(new_n7908_), .B(new_n7905_), .Y(new_n8501_));
  OAI21X1  g08245(.A0(new_n8501_), .A1(new_n7972_), .B0(new_n8071_), .Y(new_n8502_));
  AOI21X1  g08246(.A0(new_n8502_), .A1(new_n8072_), .B0(new_n8328_), .Y(new_n8503_));
  INVX1    g08247(.A(new_n8503_), .Y(new_n8504_));
  OAI21X1  g08248(.A0(new_n8329_), .A1(new_n8324_), .B0(new_n8504_), .Y(new_n8505_));
  AOI22X1  g08249(.A0(new_n2163_), .A1(\b[40] ), .B0(new_n2162_), .B1(\b[39] ), .Y(new_n8506_));
  OAI21X1  g08250(.A0(new_n2161_), .A1(new_n3575_), .B0(new_n8506_), .Y(new_n8507_));
  AOI21X1  g08251(.A0(new_n3574_), .A1(new_n1907_), .B0(new_n8507_), .Y(new_n8508_));
  XOR2X1   g08252(.A(new_n8508_), .B(new_n1911_), .Y(new_n8509_));
  XOR2X1   g08253(.A(new_n8509_), .B(new_n8505_), .Y(new_n8510_));
  XOR2X1   g08254(.A(new_n8510_), .B(new_n8500_), .Y(new_n8511_));
  XOR2X1   g08255(.A(new_n8511_), .B(new_n8398_), .Y(new_n8512_));
  AOI22X1  g08256(.A0(new_n1526_), .A1(\b[46] ), .B0(new_n1525_), .B1(\b[45] ), .Y(new_n8513_));
  OAI21X1  g08257(.A0(new_n1524_), .A1(new_n4336_), .B0(new_n8513_), .Y(new_n8514_));
  AOI21X1  g08258(.A0(new_n4509_), .A1(new_n1347_), .B0(new_n8514_), .Y(new_n8515_));
  XOR2X1   g08259(.A(new_n8515_), .B(\a[23] ), .Y(new_n8516_));
  OR2X1    g08260(.A(new_n8224_), .B(new_n8219_), .Y(new_n8517_));
  OR2X1    g08261(.A(new_n8331_), .B(new_n8225_), .Y(new_n8518_));
  AND2X1   g08262(.A(new_n8518_), .B(new_n8517_), .Y(new_n8519_));
  XOR2X1   g08263(.A(new_n8519_), .B(new_n8516_), .Y(new_n8520_));
  INVX1    g08264(.A(new_n8520_), .Y(new_n8521_));
  XOR2X1   g08265(.A(new_n8521_), .B(new_n8512_), .Y(new_n8522_));
  XOR2X1   g08266(.A(new_n8522_), .B(new_n8389_), .Y(new_n8523_));
  INVX1    g08267(.A(new_n8523_), .Y(new_n8524_));
  AOI22X1  g08268(.A0(new_n1017_), .A1(\b[52] ), .B0(new_n1016_), .B1(\b[51] ), .Y(new_n8525_));
  OAI21X1  g08269(.A0(new_n1015_), .A1(new_n5234_), .B0(new_n8525_), .Y(new_n8526_));
  AOI21X1  g08270(.A0(new_n5590_), .A1(new_n882_), .B0(new_n8526_), .Y(new_n8527_));
  XOR2X1   g08271(.A(new_n8527_), .B(\a[17] ), .Y(new_n8528_));
  INVX1    g08272(.A(new_n8206_), .Y(new_n8529_));
  NOR2X1   g08273(.A(new_n8333_), .B(new_n8209_), .Y(new_n8530_));
  AOI21X1  g08274(.A0(new_n8208_), .A1(new_n8529_), .B0(new_n8530_), .Y(new_n8531_));
  XOR2X1   g08275(.A(new_n8531_), .B(new_n8528_), .Y(new_n8532_));
  XOR2X1   g08276(.A(new_n8532_), .B(new_n8524_), .Y(new_n8533_));
  XOR2X1   g08277(.A(new_n8533_), .B(new_n8381_), .Y(new_n8534_));
  NAND2X1  g08278(.A(new_n8342_), .B(new_n8338_), .Y(new_n8535_));
  XOR2X1   g08279(.A(new_n8341_), .B(\a[14] ), .Y(new_n8536_));
  XOR2X1   g08280(.A(new_n8536_), .B(new_n8338_), .Y(new_n8537_));
  OR2X1    g08281(.A(new_n8537_), .B(new_n8335_), .Y(new_n8538_));
  AND2X1   g08282(.A(new_n8538_), .B(new_n8535_), .Y(new_n8539_));
  INVX1    g08283(.A(new_n6732_), .Y(new_n8540_));
  INVX1    g08284(.A(new_n601_), .Y(new_n8541_));
  OAI22X1  g08285(.A0(new_n661_), .A1(new_n6930_), .B0(new_n660_), .B1(new_n6933_), .Y(new_n8542_));
  AOI21X1  g08286(.A0(new_n8541_), .A1(\b[56] ), .B0(new_n8542_), .Y(new_n8543_));
  OAI21X1  g08287(.A0(new_n8540_), .A1(new_n567_), .B0(new_n8543_), .Y(new_n8544_));
  XOR2X1   g08288(.A(new_n8544_), .B(new_n515_), .Y(new_n8545_));
  XOR2X1   g08289(.A(new_n8545_), .B(new_n8539_), .Y(new_n8546_));
  XOR2X1   g08290(.A(new_n8546_), .B(new_n8534_), .Y(new_n8547_));
  OR2X1    g08291(.A(new_n8192_), .B(new_n8187_), .Y(new_n8548_));
  OAI21X1  g08292(.A0(new_n8344_), .A1(new_n8193_), .B0(new_n8548_), .Y(new_n8549_));
  INVX1    g08293(.A(new_n7338_), .Y(new_n8550_));
  INVX1    g08294(.A(new_n467_), .Y(new_n8551_));
  OAI22X1  g08295(.A0(new_n511_), .A1(new_n7748_), .B0(new_n510_), .B1(new_n7559_), .Y(new_n8552_));
  AOI21X1  g08296(.A0(new_n8551_), .A1(\b[59] ), .B0(new_n8552_), .Y(new_n8553_));
  OAI21X1  g08297(.A0(new_n8550_), .A1(new_n429_), .B0(new_n8553_), .Y(new_n8554_));
  XOR2X1   g08298(.A(new_n8554_), .B(new_n400_), .Y(new_n8555_));
  INVX1    g08299(.A(new_n8555_), .Y(new_n8556_));
  XOR2X1   g08300(.A(new_n8556_), .B(new_n8549_), .Y(new_n8557_));
  XOR2X1   g08301(.A(new_n8557_), .B(new_n8547_), .Y(new_n8558_));
  INVX1    g08302(.A(new_n8345_), .Y(new_n8559_));
  OR2X1    g08303(.A(new_n8352_), .B(new_n8349_), .Y(new_n8560_));
  OAI21X1  g08304(.A0(new_n8353_), .A1(new_n8559_), .B0(new_n8560_), .Y(new_n8561_));
  OAI22X1  g08305(.A0(new_n367_), .A1(new_n7745_), .B0(new_n416_), .B1(new_n7772_), .Y(new_n8562_));
  AOI21X1  g08306(.A0(new_n7775_), .A1(new_n308_), .B0(new_n8562_), .Y(new_n8563_));
  XOR2X1   g08307(.A(new_n8563_), .B(\a[5] ), .Y(new_n8564_));
  OR2X1    g08308(.A(new_n8564_), .B(new_n8561_), .Y(new_n8565_));
  INVX1    g08309(.A(new_n8564_), .Y(new_n8566_));
  XOR2X1   g08310(.A(new_n8566_), .B(new_n8561_), .Y(new_n8567_));
  AOI21X1  g08311(.A0(new_n8564_), .A1(new_n8561_), .B0(new_n8558_), .Y(new_n8568_));
  AOI22X1  g08312(.A0(new_n8568_), .A1(new_n8565_), .B0(new_n8567_), .B1(new_n8558_), .Y(new_n8569_));
  XOR2X1   g08313(.A(new_n8569_), .B(new_n8372_), .Y(new_n8570_));
  XOR2X1   g08314(.A(new_n8570_), .B(new_n8368_), .Y(\f[67] ));
  OAI21X1  g08315(.A0(new_n8371_), .A1(new_n8370_), .B0(new_n8569_), .Y(new_n8572_));
  OAI21X1  g08316(.A0(new_n8367_), .A1(new_n8366_), .B0(new_n8570_), .Y(new_n8573_));
  AND2X1   g08317(.A(new_n8573_), .B(new_n8572_), .Y(new_n8574_));
  AND2X1   g08318(.A(new_n8566_), .B(new_n8561_), .Y(new_n8575_));
  AOI21X1  g08319(.A0(new_n8567_), .A1(new_n8558_), .B0(new_n8575_), .Y(new_n8576_));
  AND2X1   g08320(.A(new_n8556_), .B(new_n8549_), .Y(new_n8577_));
  AOI21X1  g08321(.A0(new_n8557_), .A1(new_n8547_), .B0(new_n8577_), .Y(new_n8578_));
  NOR4X1   g08322(.A(new_n336_), .B(new_n335_), .C(new_n301_), .D(new_n7772_), .Y(new_n8579_));
  AOI21X1  g08323(.A0(new_n7774_), .A1(new_n308_), .B0(new_n8579_), .Y(new_n8580_));
  XOR2X1   g08324(.A(new_n8580_), .B(\a[5] ), .Y(new_n8581_));
  XOR2X1   g08325(.A(new_n8581_), .B(new_n8578_), .Y(new_n8582_));
  AOI22X1  g08326(.A0(new_n603_), .A1(\b[59] ), .B0(new_n602_), .B1(\b[58] ), .Y(new_n8583_));
  OAI21X1  g08327(.A0(new_n601_), .A1(new_n6933_), .B0(new_n8583_), .Y(new_n8584_));
  AOI21X1  g08328(.A0(new_n6932_), .A1(new_n518_), .B0(new_n8584_), .Y(new_n8585_));
  XOR2X1   g08329(.A(new_n8585_), .B(\a[11] ), .Y(new_n8586_));
  OR2X1    g08330(.A(new_n8380_), .B(new_n8376_), .Y(new_n8587_));
  OAI21X1  g08331(.A0(new_n8533_), .A1(new_n8381_), .B0(new_n8587_), .Y(new_n8588_));
  XOR2X1   g08332(.A(new_n8588_), .B(new_n8586_), .Y(new_n8589_));
  AOI22X1  g08333(.A0(new_n818_), .A1(\b[56] ), .B0(new_n817_), .B1(\b[55] ), .Y(new_n8590_));
  OAI21X1  g08334(.A0(new_n816_), .A1(new_n6148_), .B0(new_n8590_), .Y(new_n8591_));
  AOI21X1  g08335(.A0(new_n6342_), .A1(new_n668_), .B0(new_n8591_), .Y(new_n8592_));
  XOR2X1   g08336(.A(new_n8592_), .B(\a[14] ), .Y(new_n8593_));
  NOR2X1   g08337(.A(new_n8531_), .B(new_n8528_), .Y(new_n8594_));
  AOI21X1  g08338(.A0(new_n8532_), .A1(new_n8523_), .B0(new_n8594_), .Y(new_n8595_));
  XOR2X1   g08339(.A(new_n8595_), .B(new_n8593_), .Y(new_n8596_));
  OR2X1    g08340(.A(new_n8388_), .B(new_n8385_), .Y(new_n8597_));
  OAI21X1  g08341(.A0(new_n8522_), .A1(new_n8389_), .B0(new_n8597_), .Y(new_n8598_));
  INVX1    g08342(.A(new_n5786_), .Y(new_n8599_));
  INVX1    g08343(.A(new_n1015_), .Y(new_n8600_));
  OAI22X1  g08344(.A0(new_n1068_), .A1(new_n6151_), .B0(new_n1067_), .B1(new_n5808_), .Y(new_n8601_));
  AOI21X1  g08345(.A0(new_n8600_), .A1(\b[51] ), .B0(new_n8601_), .Y(new_n8602_));
  OAI21X1  g08346(.A0(new_n8599_), .A1(new_n934_), .B0(new_n8602_), .Y(new_n8603_));
  XOR2X1   g08347(.A(new_n8603_), .B(new_n879_), .Y(new_n8604_));
  XOR2X1   g08348(.A(new_n8604_), .B(new_n8598_), .Y(new_n8605_));
  AOI22X1  g08349(.A0(new_n1263_), .A1(\b[50] ), .B0(new_n1262_), .B1(\b[49] ), .Y(new_n8606_));
  OAI21X1  g08350(.A0(new_n1261_), .A1(new_n5036_), .B0(new_n8606_), .Y(new_n8607_));
  AOI21X1  g08351(.A0(new_n5204_), .A1(new_n1075_), .B0(new_n8607_), .Y(new_n8608_));
  XOR2X1   g08352(.A(new_n8608_), .B(\a[20] ), .Y(new_n8609_));
  AOI21X1  g08353(.A0(new_n8518_), .A1(new_n8517_), .B0(new_n8516_), .Y(new_n8610_));
  AOI21X1  g08354(.A0(new_n8520_), .A1(new_n8512_), .B0(new_n8610_), .Y(new_n8611_));
  XOR2X1   g08355(.A(new_n8611_), .B(new_n8609_), .Y(new_n8612_));
  AOI22X1  g08356(.A0(new_n1526_), .A1(\b[47] ), .B0(new_n1525_), .B1(\b[46] ), .Y(new_n8613_));
  OAI21X1  g08357(.A0(new_n1524_), .A1(new_n4674_), .B0(new_n8613_), .Y(new_n8614_));
  AOI21X1  g08358(.A0(new_n4673_), .A1(new_n1347_), .B0(new_n8614_), .Y(new_n8615_));
  XOR2X1   g08359(.A(new_n8615_), .B(\a[23] ), .Y(new_n8616_));
  OR2X1    g08360(.A(new_n8397_), .B(new_n8393_), .Y(new_n8617_));
  OR2X1    g08361(.A(new_n8511_), .B(new_n8398_), .Y(new_n8618_));
  AND2X1   g08362(.A(new_n8618_), .B(new_n8617_), .Y(new_n8619_));
  XOR2X1   g08363(.A(new_n8619_), .B(new_n8616_), .Y(new_n8620_));
  AOI22X1  g08364(.A0(new_n2163_), .A1(\b[41] ), .B0(new_n2162_), .B1(\b[40] ), .Y(new_n8621_));
  OAI21X1  g08365(.A0(new_n2161_), .A1(new_n3723_), .B0(new_n8621_), .Y(new_n8622_));
  AOI21X1  g08366(.A0(new_n3722_), .A1(new_n1907_), .B0(new_n8622_), .Y(new_n8623_));
  XOR2X1   g08367(.A(new_n8623_), .B(\a[29] ), .Y(new_n8624_));
  INVX1    g08368(.A(new_n8624_), .Y(new_n8625_));
  XOR2X1   g08369(.A(new_n8406_), .B(new_n2258_), .Y(new_n8626_));
  NOR2X1   g08370(.A(new_n8498_), .B(new_n8408_), .Y(new_n8627_));
  AOI21X1  g08371(.A0(new_n8626_), .A1(new_n8403_), .B0(new_n8627_), .Y(new_n8628_));
  XOR2X1   g08372(.A(new_n8628_), .B(new_n8625_), .Y(new_n8629_));
  AOI22X1  g08373(.A0(new_n7192_), .A1(\b[8] ), .B0(new_n7189_), .B1(\b[7] ), .Y(new_n8630_));
  OAI21X1  g08374(.A0(new_n7627_), .A1(new_n392_), .B0(new_n8630_), .Y(new_n8631_));
  AOI21X1  g08375(.A0(new_n7187_), .A1(new_n454_), .B0(new_n8631_), .Y(new_n8632_));
  XOR2X1   g08376(.A(new_n8632_), .B(\a[62] ), .Y(new_n8633_));
  AOI22X1  g08377(.A0(new_n7818_), .A1(\b[4] ), .B0(new_n7817_), .B1(\b[5] ), .Y(new_n8634_));
  XOR2X1   g08378(.A(new_n8634_), .B(\a[2] ), .Y(new_n8635_));
  XOR2X1   g08379(.A(new_n8635_), .B(new_n8633_), .Y(new_n8636_));
  INVX1    g08380(.A(new_n8636_), .Y(new_n8637_));
  NOR2X1   g08381(.A(new_n8420_), .B(new_n257_), .Y(new_n8638_));
  INVX1    g08382(.A(new_n8421_), .Y(new_n8639_));
  AOI21X1  g08383(.A0(new_n8639_), .A1(new_n8419_), .B0(new_n8638_), .Y(new_n8640_));
  XOR2X1   g08384(.A(new_n8640_), .B(new_n8637_), .Y(new_n8641_));
  INVX1    g08385(.A(new_n8641_), .Y(new_n8642_));
  AOI22X1  g08386(.A0(new_n6603_), .A1(\b[11] ), .B0(new_n6600_), .B1(\b[10] ), .Y(new_n8643_));
  OAI21X1  g08387(.A0(new_n6804_), .A1(new_n590_), .B0(new_n8643_), .Y(new_n8644_));
  AOI21X1  g08388(.A0(new_n6598_), .A1(new_n589_), .B0(new_n8644_), .Y(new_n8645_));
  XOR2X1   g08389(.A(new_n8645_), .B(\a[59] ), .Y(new_n8646_));
  XOR2X1   g08390(.A(new_n8646_), .B(new_n8642_), .Y(new_n8647_));
  INVX1    g08391(.A(new_n8647_), .Y(new_n8648_));
  AOI21X1  g08392(.A0(new_n8424_), .A1(new_n8423_), .B0(new_n8422_), .Y(new_n8649_));
  INVX1    g08393(.A(new_n8430_), .Y(new_n8650_));
  AOI21X1  g08394(.A0(new_n8650_), .A1(new_n8426_), .B0(new_n8649_), .Y(new_n8651_));
  XOR2X1   g08395(.A(new_n8651_), .B(new_n8648_), .Y(new_n8652_));
  AOI22X1  g08396(.A0(new_n6438_), .A1(\b[14] ), .B0(new_n6437_), .B1(\b[13] ), .Y(new_n8653_));
  OAI21X1  g08397(.A0(new_n6436_), .A1(new_n713_), .B0(new_n8653_), .Y(new_n8654_));
  AOI21X1  g08398(.A0(new_n6023_), .A1(new_n734_), .B0(new_n8654_), .Y(new_n8655_));
  XOR2X1   g08399(.A(new_n8655_), .B(\a[56] ), .Y(new_n8656_));
  XOR2X1   g08400(.A(new_n8656_), .B(new_n8652_), .Y(new_n8657_));
  AOI21X1  g08401(.A0(new_n8433_), .A1(new_n8432_), .B0(new_n8431_), .Y(new_n8658_));
  AOI21X1  g08402(.A0(new_n8440_), .A1(new_n8435_), .B0(new_n8658_), .Y(new_n8659_));
  XOR2X1   g08403(.A(new_n8659_), .B(new_n8657_), .Y(new_n8660_));
  AOI22X1  g08404(.A0(new_n5430_), .A1(\b[17] ), .B0(new_n5427_), .B1(\b[16] ), .Y(new_n8661_));
  OAI21X1  g08405(.A0(new_n5891_), .A1(new_n977_), .B0(new_n8661_), .Y(new_n8662_));
  AOI21X1  g08406(.A0(new_n5425_), .A1(new_n976_), .B0(new_n8662_), .Y(new_n8663_));
  XOR2X1   g08407(.A(new_n8663_), .B(\a[53] ), .Y(new_n8664_));
  XOR2X1   g08408(.A(new_n8664_), .B(new_n8660_), .Y(new_n8665_));
  NOR2X1   g08409(.A(new_n8445_), .B(new_n8442_), .Y(new_n8666_));
  INVX1    g08410(.A(new_n8450_), .Y(new_n8667_));
  AOI21X1  g08411(.A0(new_n8667_), .A1(new_n8446_), .B0(new_n8666_), .Y(new_n8668_));
  XOR2X1   g08412(.A(new_n8668_), .B(new_n8665_), .Y(new_n8669_));
  INVX1    g08413(.A(new_n8669_), .Y(new_n8670_));
  AOI22X1  g08414(.A0(new_n4880_), .A1(\b[20] ), .B0(new_n4877_), .B1(\b[19] ), .Y(new_n8671_));
  OAI21X1  g08415(.A0(new_n5291_), .A1(new_n1115_), .B0(new_n8671_), .Y(new_n8672_));
  AOI21X1  g08416(.A0(new_n4875_), .A1(new_n1217_), .B0(new_n8672_), .Y(new_n8673_));
  XOR2X1   g08417(.A(new_n8673_), .B(\a[50] ), .Y(new_n8674_));
  XOR2X1   g08418(.A(new_n8674_), .B(new_n8670_), .Y(new_n8675_));
  INVX1    g08419(.A(new_n8675_), .Y(new_n8676_));
  NOR2X1   g08420(.A(new_n8454_), .B(new_n8451_), .Y(new_n8677_));
  INVX1    g08421(.A(new_n8459_), .Y(new_n8678_));
  AOI21X1  g08422(.A0(new_n8678_), .A1(new_n8455_), .B0(new_n8677_), .Y(new_n8679_));
  XOR2X1   g08423(.A(new_n8679_), .B(new_n8676_), .Y(new_n8680_));
  AOI22X1  g08424(.A0(new_n4572_), .A1(\b[23] ), .B0(new_n4571_), .B1(\b[22] ), .Y(new_n8681_));
  OAI21X1  g08425(.A0(new_n4740_), .A1(new_n1482_), .B0(new_n8681_), .Y(new_n8682_));
  AOI21X1  g08426(.A0(new_n4375_), .A1(new_n1481_), .B0(new_n8682_), .Y(new_n8683_));
  XOR2X1   g08427(.A(new_n8683_), .B(\a[47] ), .Y(new_n8684_));
  XOR2X1   g08428(.A(new_n8684_), .B(new_n8680_), .Y(new_n8685_));
  NOR2X1   g08429(.A(new_n8463_), .B(new_n8460_), .Y(new_n8686_));
  INVX1    g08430(.A(new_n8468_), .Y(new_n8687_));
  AOI21X1  g08431(.A0(new_n8687_), .A1(new_n8464_), .B0(new_n8686_), .Y(new_n8688_));
  XOR2X1   g08432(.A(new_n8688_), .B(new_n8685_), .Y(new_n8689_));
  AOI22X1  g08433(.A0(new_n4095_), .A1(\b[26] ), .B0(new_n4094_), .B1(\b[25] ), .Y(new_n8690_));
  OAI21X1  g08434(.A0(new_n4233_), .A1(new_n1588_), .B0(new_n8690_), .Y(new_n8691_));
  AOI21X1  g08435(.A0(new_n3901_), .A1(new_n1783_), .B0(new_n8691_), .Y(new_n8692_));
  XOR2X1   g08436(.A(new_n8692_), .B(\a[44] ), .Y(new_n8693_));
  XOR2X1   g08437(.A(new_n8693_), .B(new_n8689_), .Y(new_n8694_));
  NOR2X1   g08438(.A(new_n8471_), .B(new_n8469_), .Y(new_n8695_));
  INVX1    g08439(.A(new_n8476_), .Y(new_n8696_));
  AOI21X1  g08440(.A0(new_n8696_), .A1(new_n8472_), .B0(new_n8695_), .Y(new_n8697_));
  XOR2X1   g08441(.A(new_n8697_), .B(new_n8694_), .Y(new_n8698_));
  AOI22X1  g08442(.A0(new_n3652_), .A1(\b[29] ), .B0(new_n3651_), .B1(\b[28] ), .Y(new_n8699_));
  OAI21X1  g08443(.A0(new_n3778_), .A1(new_n2126_), .B0(new_n8699_), .Y(new_n8700_));
  AOI21X1  g08444(.A0(new_n3480_), .A1(new_n2125_), .B0(new_n8700_), .Y(new_n8701_));
  XOR2X1   g08445(.A(new_n8701_), .B(\a[41] ), .Y(new_n8702_));
  XOR2X1   g08446(.A(new_n8702_), .B(new_n8698_), .Y(new_n8703_));
  NOR2X1   g08447(.A(new_n8480_), .B(new_n8477_), .Y(new_n8704_));
  INVX1    g08448(.A(new_n8485_), .Y(new_n8705_));
  AOI21X1  g08449(.A0(new_n8705_), .A1(new_n8481_), .B0(new_n8704_), .Y(new_n8706_));
  XOR2X1   g08450(.A(new_n8706_), .B(new_n8703_), .Y(new_n8707_));
  INVX1    g08451(.A(new_n8707_), .Y(new_n8708_));
  AOI22X1  g08452(.A0(new_n3204_), .A1(\b[32] ), .B0(new_n3203_), .B1(\b[31] ), .Y(new_n8709_));
  OAI21X1  g08453(.A0(new_n3321_), .A1(new_n2356_), .B0(new_n8709_), .Y(new_n8710_));
  AOI21X1  g08454(.A0(new_n3080_), .A1(new_n2495_), .B0(new_n8710_), .Y(new_n8711_));
  XOR2X1   g08455(.A(new_n8711_), .B(\a[38] ), .Y(new_n8712_));
  XOR2X1   g08456(.A(new_n8712_), .B(new_n8708_), .Y(new_n8713_));
  INVX1    g08457(.A(new_n8713_), .Y(new_n8714_));
  OR2X1    g08458(.A(new_n8490_), .B(new_n8486_), .Y(new_n8715_));
  OR2X1    g08459(.A(new_n8495_), .B(new_n8491_), .Y(new_n8716_));
  AND2X1   g08460(.A(new_n8716_), .B(new_n8715_), .Y(new_n8717_));
  XOR2X1   g08461(.A(new_n8717_), .B(new_n8714_), .Y(new_n8718_));
  AOI22X1  g08462(.A0(new_n2813_), .A1(\b[35] ), .B0(new_n2812_), .B1(\b[34] ), .Y(new_n8719_));
  OAI21X1  g08463(.A0(new_n2946_), .A1(new_n2893_), .B0(new_n8719_), .Y(new_n8720_));
  AOI21X1  g08464(.A0(new_n2892_), .A1(new_n2652_), .B0(new_n8720_), .Y(new_n8721_));
  XOR2X1   g08465(.A(new_n8721_), .B(\a[35] ), .Y(new_n8722_));
  XOR2X1   g08466(.A(new_n8722_), .B(new_n8718_), .Y(new_n8723_));
  OAI21X1  g08467(.A0(new_n8400_), .A1(new_n8414_), .B0(new_n8496_), .Y(new_n8724_));
  OR2X1    g08468(.A(new_n8497_), .B(new_n8412_), .Y(new_n8725_));
  AND2X1   g08469(.A(new_n8725_), .B(new_n8724_), .Y(new_n8726_));
  AOI22X1  g08470(.A0(new_n2545_), .A1(\b[38] ), .B0(new_n2544_), .B1(\b[37] ), .Y(new_n8727_));
  OAI21X1  g08471(.A0(new_n2543_), .A1(new_n3276_), .B0(new_n8727_), .Y(new_n8728_));
  AOI21X1  g08472(.A0(new_n3275_), .A1(new_n2260_), .B0(new_n8728_), .Y(new_n8729_));
  XOR2X1   g08473(.A(new_n8729_), .B(\a[32] ), .Y(new_n8730_));
  XOR2X1   g08474(.A(new_n8730_), .B(new_n8726_), .Y(new_n8731_));
  XOR2X1   g08475(.A(new_n8731_), .B(new_n8723_), .Y(new_n8732_));
  XOR2X1   g08476(.A(new_n8732_), .B(new_n8629_), .Y(new_n8733_));
  AND2X1   g08477(.A(new_n8509_), .B(new_n8505_), .Y(new_n8734_));
  AOI21X1  g08478(.A0(new_n8510_), .A1(new_n8499_), .B0(new_n8734_), .Y(new_n8735_));
  INVX1    g08479(.A(new_n4178_), .Y(new_n8736_));
  OAI22X1  g08480(.A0(new_n1623_), .A1(new_n4336_), .B0(new_n1620_), .B1(new_n4339_), .Y(new_n8737_));
  AOI21X1  g08481(.A0(new_n1725_), .A1(\b[42] ), .B0(new_n8737_), .Y(new_n8738_));
  OAI21X1  g08482(.A0(new_n8736_), .A1(new_n1723_), .B0(new_n8738_), .Y(new_n8739_));
  XOR2X1   g08483(.A(new_n8739_), .B(new_n1621_), .Y(new_n8740_));
  INVX1    g08484(.A(new_n8740_), .Y(new_n8741_));
  XOR2X1   g08485(.A(new_n8741_), .B(new_n8735_), .Y(new_n8742_));
  XOR2X1   g08486(.A(new_n8742_), .B(new_n8733_), .Y(new_n8743_));
  XOR2X1   g08487(.A(new_n8743_), .B(new_n8620_), .Y(new_n8744_));
  XOR2X1   g08488(.A(new_n8744_), .B(new_n8612_), .Y(new_n8745_));
  XOR2X1   g08489(.A(new_n8745_), .B(new_n8605_), .Y(new_n8746_));
  INVX1    g08490(.A(new_n8746_), .Y(new_n8747_));
  XOR2X1   g08491(.A(new_n8747_), .B(new_n8596_), .Y(new_n8748_));
  XOR2X1   g08492(.A(new_n8748_), .B(new_n8589_), .Y(new_n8749_));
  AOI21X1  g08493(.A0(new_n8538_), .A1(new_n8535_), .B0(new_n8545_), .Y(new_n8750_));
  AOI21X1  g08494(.A0(new_n8546_), .A1(new_n8534_), .B0(new_n8750_), .Y(new_n8751_));
  INVX1    g08495(.A(new_n8751_), .Y(new_n8752_));
  INVX1    g08496(.A(new_n7558_), .Y(new_n8753_));
  OAI22X1  g08497(.A0(new_n511_), .A1(new_n7745_), .B0(new_n510_), .B1(new_n7748_), .Y(new_n8754_));
  AOI21X1  g08498(.A0(new_n8551_), .A1(\b[60] ), .B0(new_n8754_), .Y(new_n8755_));
  OAI21X1  g08499(.A0(new_n8753_), .A1(new_n429_), .B0(new_n8755_), .Y(new_n8756_));
  XOR2X1   g08500(.A(new_n8756_), .B(new_n400_), .Y(new_n8757_));
  OR2X1    g08501(.A(new_n8757_), .B(new_n8752_), .Y(new_n8758_));
  XOR2X1   g08502(.A(new_n8757_), .B(new_n8751_), .Y(new_n8759_));
  AOI21X1  g08503(.A0(new_n8757_), .A1(new_n8752_), .B0(new_n8749_), .Y(new_n8760_));
  AOI22X1  g08504(.A0(new_n8760_), .A1(new_n8758_), .B0(new_n8759_), .B1(new_n8749_), .Y(new_n8761_));
  XOR2X1   g08505(.A(new_n8761_), .B(new_n8582_), .Y(new_n8762_));
  XOR2X1   g08506(.A(new_n8762_), .B(new_n8576_), .Y(new_n8763_));
  XOR2X1   g08507(.A(new_n8763_), .B(new_n8574_), .Y(\f[68] ));
  AND2X1   g08508(.A(new_n8567_), .B(new_n8558_), .Y(new_n8765_));
  OR2X1    g08509(.A(new_n8765_), .B(new_n8575_), .Y(new_n8766_));
  AND2X1   g08510(.A(new_n8762_), .B(new_n8766_), .Y(new_n8767_));
  AOI21X1  g08511(.A0(new_n8573_), .A1(new_n8572_), .B0(new_n8763_), .Y(new_n8768_));
  OR2X1    g08512(.A(new_n8768_), .B(new_n8767_), .Y(new_n8769_));
  NOR2X1   g08513(.A(new_n8581_), .B(new_n8578_), .Y(new_n8770_));
  AOI21X1  g08514(.A0(new_n8761_), .A1(new_n8582_), .B0(new_n8770_), .Y(new_n8771_));
  NOR2X1   g08515(.A(new_n8757_), .B(new_n8751_), .Y(new_n8772_));
  AOI21X1  g08516(.A0(new_n8759_), .A1(new_n8749_), .B0(new_n8772_), .Y(new_n8773_));
  AOI22X1  g08517(.A0(new_n469_), .A1(\b[63] ), .B0(new_n468_), .B1(\b[62] ), .Y(new_n8774_));
  OAI21X1  g08518(.A0(new_n467_), .A1(new_n7748_), .B0(new_n8774_), .Y(new_n8775_));
  AOI21X1  g08519(.A0(new_n7747_), .A1(new_n404_), .B0(new_n8775_), .Y(new_n8776_));
  XOR2X1   g08520(.A(new_n8776_), .B(\a[8] ), .Y(new_n8777_));
  XOR2X1   g08521(.A(new_n8777_), .B(new_n8773_), .Y(new_n8778_));
  AOI22X1  g08522(.A0(new_n603_), .A1(\b[60] ), .B0(new_n602_), .B1(\b[59] ), .Y(new_n8779_));
  OAI21X1  g08523(.A0(new_n601_), .A1(new_n6930_), .B0(new_n8779_), .Y(new_n8780_));
  AOI21X1  g08524(.A0(new_n6951_), .A1(new_n518_), .B0(new_n8780_), .Y(new_n8781_));
  XOR2X1   g08525(.A(new_n8781_), .B(\a[11] ), .Y(new_n8782_));
  INVX1    g08526(.A(new_n8586_), .Y(new_n8783_));
  NOR2X1   g08527(.A(new_n8748_), .B(new_n8589_), .Y(new_n8784_));
  AOI21X1  g08528(.A0(new_n8588_), .A1(new_n8783_), .B0(new_n8784_), .Y(new_n8785_));
  XOR2X1   g08529(.A(new_n8785_), .B(new_n8782_), .Y(new_n8786_));
  OR2X1    g08530(.A(new_n8522_), .B(new_n8389_), .Y(new_n8787_));
  AOI21X1  g08531(.A0(new_n8787_), .A1(new_n8597_), .B0(new_n8604_), .Y(new_n8788_));
  INVX1    g08532(.A(new_n8788_), .Y(new_n8789_));
  OR2X1    g08533(.A(new_n8745_), .B(new_n8605_), .Y(new_n8790_));
  NAND2X1  g08534(.A(new_n8790_), .B(new_n8789_), .Y(new_n8791_));
  AOI22X1  g08535(.A0(new_n1017_), .A1(\b[54] ), .B0(new_n1016_), .B1(\b[53] ), .Y(new_n8792_));
  OAI21X1  g08536(.A0(new_n1015_), .A1(new_n5808_), .B0(new_n8792_), .Y(new_n8793_));
  AOI21X1  g08537(.A0(new_n5807_), .A1(new_n882_), .B0(new_n8793_), .Y(new_n8794_));
  XOR2X1   g08538(.A(new_n8794_), .B(\a[17] ), .Y(new_n8795_));
  XOR2X1   g08539(.A(new_n8795_), .B(new_n8791_), .Y(new_n8796_));
  AOI22X1  g08540(.A0(new_n1526_), .A1(\b[48] ), .B0(new_n1525_), .B1(\b[47] ), .Y(new_n8797_));
  OAI21X1  g08541(.A0(new_n1524_), .A1(new_n4693_), .B0(new_n8797_), .Y(new_n8798_));
  AOI21X1  g08542(.A0(new_n4692_), .A1(new_n1347_), .B0(new_n8798_), .Y(new_n8799_));
  XOR2X1   g08543(.A(new_n8799_), .B(\a[23] ), .Y(new_n8800_));
  AOI21X1  g08544(.A0(new_n8618_), .A1(new_n8617_), .B0(new_n8616_), .Y(new_n8801_));
  INVX1    g08545(.A(new_n8743_), .Y(new_n8802_));
  AOI21X1  g08546(.A0(new_n8802_), .A1(new_n8620_), .B0(new_n8801_), .Y(new_n8803_));
  XOR2X1   g08547(.A(new_n8803_), .B(new_n8800_), .Y(new_n8804_));
  NOR2X1   g08548(.A(new_n8740_), .B(new_n8735_), .Y(new_n8805_));
  XOR2X1   g08549(.A(new_n8740_), .B(new_n8735_), .Y(new_n8806_));
  AOI21X1  g08550(.A0(new_n8806_), .A1(new_n8733_), .B0(new_n8805_), .Y(new_n8807_));
  AOI22X1  g08551(.A0(new_n1814_), .A1(\b[45] ), .B0(new_n1813_), .B1(\b[44] ), .Y(new_n8808_));
  OAI21X1  g08552(.A0(new_n1812_), .A1(new_n4339_), .B0(new_n8808_), .Y(new_n8809_));
  AOI21X1  g08553(.A0(new_n4338_), .A1(new_n1617_), .B0(new_n8809_), .Y(new_n8810_));
  XOR2X1   g08554(.A(new_n8810_), .B(\a[26] ), .Y(new_n8811_));
  XOR2X1   g08555(.A(new_n8811_), .B(new_n8807_), .Y(new_n8812_));
  AOI22X1  g08556(.A0(new_n2163_), .A1(\b[42] ), .B0(new_n2162_), .B1(\b[41] ), .Y(new_n8813_));
  OAI21X1  g08557(.A0(new_n2161_), .A1(new_n3720_), .B0(new_n8813_), .Y(new_n8814_));
  AOI21X1  g08558(.A0(new_n3860_), .A1(new_n1907_), .B0(new_n8814_), .Y(new_n8815_));
  XOR2X1   g08559(.A(new_n8815_), .B(\a[29] ), .Y(new_n8816_));
  OR2X1    g08560(.A(new_n8628_), .B(new_n8624_), .Y(new_n8817_));
  OR2X1    g08561(.A(new_n8732_), .B(new_n8629_), .Y(new_n8818_));
  AND2X1   g08562(.A(new_n8818_), .B(new_n8817_), .Y(new_n8819_));
  XOR2X1   g08563(.A(new_n8819_), .B(new_n8816_), .Y(new_n8820_));
  OR2X1    g08564(.A(new_n8717_), .B(new_n8714_), .Y(new_n8821_));
  AND2X1   g08565(.A(new_n8717_), .B(new_n8714_), .Y(new_n8822_));
  OAI21X1  g08566(.A0(new_n8722_), .A1(new_n8822_), .B0(new_n8821_), .Y(new_n8823_));
  NOR2X1   g08567(.A(new_n8706_), .B(new_n8703_), .Y(new_n8824_));
  INVX1    g08568(.A(new_n8824_), .Y(new_n8825_));
  OAI21X1  g08569(.A0(new_n8712_), .A1(new_n8708_), .B0(new_n8825_), .Y(new_n8826_));
  NOR2X1   g08570(.A(new_n8697_), .B(new_n8694_), .Y(new_n8827_));
  INVX1    g08571(.A(new_n8827_), .Y(new_n8828_));
  INVX1    g08572(.A(new_n8698_), .Y(new_n8829_));
  OAI21X1  g08573(.A0(new_n8702_), .A1(new_n8829_), .B0(new_n8828_), .Y(new_n8830_));
  INVX1    g08574(.A(new_n8830_), .Y(new_n8831_));
  NOR2X1   g08575(.A(new_n8679_), .B(new_n8676_), .Y(new_n8832_));
  INVX1    g08576(.A(new_n8832_), .Y(new_n8833_));
  INVX1    g08577(.A(new_n8680_), .Y(new_n8834_));
  OAI21X1  g08578(.A0(new_n8684_), .A1(new_n8834_), .B0(new_n8833_), .Y(new_n8835_));
  OR2X1    g08579(.A(new_n8668_), .B(new_n8665_), .Y(new_n8836_));
  OAI21X1  g08580(.A0(new_n8674_), .A1(new_n8670_), .B0(new_n8836_), .Y(new_n8837_));
  OR2X1    g08581(.A(new_n8640_), .B(new_n8637_), .Y(new_n8838_));
  OAI21X1  g08582(.A0(new_n8646_), .A1(new_n8642_), .B0(new_n8838_), .Y(new_n8839_));
  AOI22X1  g08583(.A0(new_n6603_), .A1(\b[12] ), .B0(new_n6600_), .B1(\b[11] ), .Y(new_n8840_));
  OAI21X1  g08584(.A0(new_n6804_), .A1(new_n587_), .B0(new_n8840_), .Y(new_n8841_));
  AOI21X1  g08585(.A0(new_n6598_), .A1(new_n635_), .B0(new_n8841_), .Y(new_n8842_));
  XOR2X1   g08586(.A(new_n8842_), .B(\a[59] ), .Y(new_n8843_));
  OR2X1    g08587(.A(new_n8634_), .B(new_n257_), .Y(new_n8844_));
  OAI21X1  g08588(.A0(new_n8635_), .A1(new_n8633_), .B0(new_n8844_), .Y(new_n8845_));
  INVX1    g08589(.A(new_n8845_), .Y(new_n8846_));
  AOI22X1  g08590(.A0(new_n7818_), .A1(\b[5] ), .B0(new_n7817_), .B1(\b[6] ), .Y(new_n8847_));
  XOR2X1   g08591(.A(\a[5] ), .B(new_n257_), .Y(new_n8848_));
  XOR2X1   g08592(.A(new_n8848_), .B(new_n8847_), .Y(new_n8849_));
  XOR2X1   g08593(.A(new_n8849_), .B(new_n8846_), .Y(new_n8850_));
  AOI22X1  g08594(.A0(new_n7192_), .A1(\b[9] ), .B0(new_n7189_), .B1(\b[8] ), .Y(new_n8851_));
  OAI21X1  g08595(.A0(new_n7627_), .A1(new_n492_), .B0(new_n8851_), .Y(new_n8852_));
  AOI21X1  g08596(.A0(new_n7187_), .A1(new_n491_), .B0(new_n8852_), .Y(new_n8853_));
  XOR2X1   g08597(.A(new_n8853_), .B(\a[62] ), .Y(new_n8854_));
  XOR2X1   g08598(.A(new_n8854_), .B(new_n8850_), .Y(new_n8855_));
  XOR2X1   g08599(.A(new_n8855_), .B(new_n8843_), .Y(new_n8856_));
  XOR2X1   g08600(.A(new_n8856_), .B(new_n8839_), .Y(new_n8857_));
  AOI22X1  g08601(.A0(new_n6438_), .A1(\b[15] ), .B0(new_n6437_), .B1(\b[14] ), .Y(new_n8858_));
  OAI21X1  g08602(.A0(new_n6436_), .A1(new_n795_), .B0(new_n8858_), .Y(new_n8859_));
  AOI21X1  g08603(.A0(new_n6023_), .A1(new_n794_), .B0(new_n8859_), .Y(new_n8860_));
  XOR2X1   g08604(.A(new_n8860_), .B(\a[56] ), .Y(new_n8861_));
  XOR2X1   g08605(.A(new_n8861_), .B(new_n8857_), .Y(new_n8862_));
  INVX1    g08606(.A(new_n8862_), .Y(new_n8863_));
  NOR2X1   g08607(.A(new_n8651_), .B(new_n8648_), .Y(new_n8864_));
  INVX1    g08608(.A(new_n8656_), .Y(new_n8865_));
  AOI21X1  g08609(.A0(new_n8865_), .A1(new_n8652_), .B0(new_n8864_), .Y(new_n8866_));
  XOR2X1   g08610(.A(new_n8866_), .B(new_n8863_), .Y(new_n8867_));
  AOI22X1  g08611(.A0(new_n5430_), .A1(\b[18] ), .B0(new_n5427_), .B1(\b[17] ), .Y(new_n8868_));
  OAI21X1  g08612(.A0(new_n5891_), .A1(new_n974_), .B0(new_n8868_), .Y(new_n8869_));
  AOI21X1  g08613(.A0(new_n5425_), .A1(new_n1042_), .B0(new_n8869_), .Y(new_n8870_));
  XOR2X1   g08614(.A(new_n8870_), .B(\a[53] ), .Y(new_n8871_));
  XOR2X1   g08615(.A(new_n8871_), .B(new_n8867_), .Y(new_n8872_));
  NOR2X1   g08616(.A(new_n8659_), .B(new_n8657_), .Y(new_n8873_));
  INVX1    g08617(.A(new_n8664_), .Y(new_n8874_));
  AOI21X1  g08618(.A0(new_n8874_), .A1(new_n8660_), .B0(new_n8873_), .Y(new_n8875_));
  XOR2X1   g08619(.A(new_n8875_), .B(new_n8872_), .Y(new_n8876_));
  AOI22X1  g08620(.A0(new_n4880_), .A1(\b[21] ), .B0(new_n4877_), .B1(\b[20] ), .Y(new_n8877_));
  OAI21X1  g08621(.A0(new_n5291_), .A1(new_n1300_), .B0(new_n8877_), .Y(new_n8878_));
  AOI21X1  g08622(.A0(new_n4875_), .A1(new_n1299_), .B0(new_n8878_), .Y(new_n8879_));
  XOR2X1   g08623(.A(new_n8879_), .B(\a[50] ), .Y(new_n8880_));
  XOR2X1   g08624(.A(new_n8880_), .B(new_n8876_), .Y(new_n8881_));
  XOR2X1   g08625(.A(new_n8881_), .B(new_n8837_), .Y(new_n8882_));
  AOI22X1  g08626(.A0(new_n4572_), .A1(\b[24] ), .B0(new_n4571_), .B1(\b[23] ), .Y(new_n8883_));
  OAI21X1  g08627(.A0(new_n4740_), .A1(new_n1479_), .B0(new_n8883_), .Y(new_n8884_));
  AOI21X1  g08628(.A0(new_n4375_), .A1(new_n1572_), .B0(new_n8884_), .Y(new_n8885_));
  XOR2X1   g08629(.A(new_n8885_), .B(\a[47] ), .Y(new_n8886_));
  XOR2X1   g08630(.A(new_n8886_), .B(new_n8882_), .Y(new_n8887_));
  XOR2X1   g08631(.A(new_n8887_), .B(new_n8835_), .Y(new_n8888_));
  AOI22X1  g08632(.A0(new_n4095_), .A1(\b[27] ), .B0(new_n4094_), .B1(\b[26] ), .Y(new_n8889_));
  OAI21X1  g08633(.A0(new_n4233_), .A1(new_n1880_), .B0(new_n8889_), .Y(new_n8890_));
  AOI21X1  g08634(.A0(new_n3901_), .A1(new_n1879_), .B0(new_n8890_), .Y(new_n8891_));
  XOR2X1   g08635(.A(new_n8891_), .B(\a[44] ), .Y(new_n8892_));
  XOR2X1   g08636(.A(new_n8892_), .B(new_n8888_), .Y(new_n8893_));
  NOR2X1   g08637(.A(new_n8688_), .B(new_n8685_), .Y(new_n8894_));
  INVX1    g08638(.A(new_n8693_), .Y(new_n8895_));
  AOI21X1  g08639(.A0(new_n8895_), .A1(new_n8689_), .B0(new_n8894_), .Y(new_n8896_));
  XOR2X1   g08640(.A(new_n8896_), .B(new_n8893_), .Y(new_n8897_));
  AOI22X1  g08641(.A0(new_n3652_), .A1(\b[30] ), .B0(new_n3651_), .B1(\b[29] ), .Y(new_n8898_));
  OAI21X1  g08642(.A0(new_n3778_), .A1(new_n2231_), .B0(new_n8898_), .Y(new_n8899_));
  AOI21X1  g08643(.A0(new_n3480_), .A1(new_n2230_), .B0(new_n8899_), .Y(new_n8900_));
  XOR2X1   g08644(.A(new_n8900_), .B(\a[41] ), .Y(new_n8901_));
  INVX1    g08645(.A(new_n8901_), .Y(new_n8902_));
  NOR2X1   g08646(.A(new_n8902_), .B(new_n8897_), .Y(new_n8903_));
  AND2X1   g08647(.A(new_n8902_), .B(new_n8897_), .Y(new_n8904_));
  NOR3X1   g08648(.A(new_n8904_), .B(new_n8903_), .C(new_n8831_), .Y(new_n8905_));
  NOR2X1   g08649(.A(new_n8905_), .B(new_n8904_), .Y(new_n8906_));
  INVX1    g08650(.A(new_n8906_), .Y(new_n8907_));
  OAI22X1  g08651(.A0(new_n8907_), .A1(new_n8903_), .B0(new_n8905_), .B1(new_n8831_), .Y(new_n8908_));
  AOI22X1  g08652(.A0(new_n3204_), .A1(\b[33] ), .B0(new_n3203_), .B1(\b[32] ), .Y(new_n8909_));
  OAI21X1  g08653(.A0(new_n3321_), .A1(new_n2615_), .B0(new_n8909_), .Y(new_n8910_));
  AOI21X1  g08654(.A0(new_n3080_), .A1(new_n2614_), .B0(new_n8910_), .Y(new_n8911_));
  XOR2X1   g08655(.A(new_n8911_), .B(\a[38] ), .Y(new_n8912_));
  XOR2X1   g08656(.A(new_n8912_), .B(new_n8908_), .Y(new_n8913_));
  XOR2X1   g08657(.A(new_n8913_), .B(new_n8826_), .Y(new_n8914_));
  AOI22X1  g08658(.A0(new_n2813_), .A1(\b[36] ), .B0(new_n2812_), .B1(\b[35] ), .Y(new_n8915_));
  OAI21X1  g08659(.A0(new_n2946_), .A1(new_n2890_), .B0(new_n8915_), .Y(new_n8916_));
  AOI21X1  g08660(.A0(new_n3015_), .A1(new_n2652_), .B0(new_n8916_), .Y(new_n8917_));
  XOR2X1   g08661(.A(new_n8917_), .B(\a[35] ), .Y(new_n8918_));
  XOR2X1   g08662(.A(new_n8918_), .B(new_n8914_), .Y(new_n8919_));
  XOR2X1   g08663(.A(new_n8919_), .B(new_n8823_), .Y(new_n8920_));
  AOI22X1  g08664(.A0(new_n2545_), .A1(\b[39] ), .B0(new_n2544_), .B1(\b[38] ), .Y(new_n8921_));
  OAI21X1  g08665(.A0(new_n2543_), .A1(new_n3413_), .B0(new_n8921_), .Y(new_n8922_));
  AOI21X1  g08666(.A0(new_n3412_), .A1(new_n2260_), .B0(new_n8922_), .Y(new_n8923_));
  XOR2X1   g08667(.A(new_n8923_), .B(\a[32] ), .Y(new_n8924_));
  INVX1    g08668(.A(new_n8723_), .Y(new_n8925_));
  AOI21X1  g08669(.A0(new_n8725_), .A1(new_n8724_), .B0(new_n8730_), .Y(new_n8926_));
  AOI21X1  g08670(.A0(new_n8731_), .A1(new_n8925_), .B0(new_n8926_), .Y(new_n8927_));
  XOR2X1   g08671(.A(new_n8927_), .B(new_n8924_), .Y(new_n8928_));
  XOR2X1   g08672(.A(new_n8928_), .B(new_n8920_), .Y(new_n8929_));
  XOR2X1   g08673(.A(new_n8929_), .B(new_n8820_), .Y(new_n8930_));
  XOR2X1   g08674(.A(new_n8930_), .B(new_n8812_), .Y(new_n8931_));
  INVX1    g08675(.A(new_n8931_), .Y(new_n8932_));
  XOR2X1   g08676(.A(new_n8932_), .B(new_n8804_), .Y(new_n8933_));
  AOI22X1  g08677(.A0(new_n1263_), .A1(\b[51] ), .B0(new_n1262_), .B1(\b[50] ), .Y(new_n8934_));
  OAI21X1  g08678(.A0(new_n1261_), .A1(new_n5237_), .B0(new_n8934_), .Y(new_n8935_));
  AOI21X1  g08679(.A0(new_n5236_), .A1(new_n1075_), .B0(new_n8935_), .Y(new_n8936_));
  XOR2X1   g08680(.A(new_n8936_), .B(\a[20] ), .Y(new_n8937_));
  NOR2X1   g08681(.A(new_n8611_), .B(new_n8609_), .Y(new_n8938_));
  INVX1    g08682(.A(new_n8744_), .Y(new_n8939_));
  AOI21X1  g08683(.A0(new_n8939_), .A1(new_n8612_), .B0(new_n8938_), .Y(new_n8940_));
  XOR2X1   g08684(.A(new_n8940_), .B(new_n8937_), .Y(new_n8941_));
  XOR2X1   g08685(.A(new_n8941_), .B(new_n8933_), .Y(new_n8942_));
  XOR2X1   g08686(.A(new_n8942_), .B(new_n8796_), .Y(new_n8943_));
  INVX1    g08687(.A(new_n8943_), .Y(new_n8944_));
  AOI22X1  g08688(.A0(new_n818_), .A1(\b[57] ), .B0(new_n817_), .B1(\b[56] ), .Y(new_n8945_));
  OAI21X1  g08689(.A0(new_n816_), .A1(new_n6523_), .B0(new_n8945_), .Y(new_n8946_));
  AOI21X1  g08690(.A0(new_n6522_), .A1(new_n668_), .B0(new_n8946_), .Y(new_n8947_));
  XOR2X1   g08691(.A(new_n8947_), .B(\a[14] ), .Y(new_n8948_));
  NOR2X1   g08692(.A(new_n8595_), .B(new_n8593_), .Y(new_n8949_));
  AOI21X1  g08693(.A0(new_n8746_), .A1(new_n8596_), .B0(new_n8949_), .Y(new_n8950_));
  XOR2X1   g08694(.A(new_n8950_), .B(new_n8948_), .Y(new_n8951_));
  XOR2X1   g08695(.A(new_n8951_), .B(new_n8944_), .Y(new_n8952_));
  XOR2X1   g08696(.A(new_n8952_), .B(new_n8786_), .Y(new_n8953_));
  XOR2X1   g08697(.A(new_n8953_), .B(new_n8778_), .Y(new_n8954_));
  XOR2X1   g08698(.A(new_n8954_), .B(new_n8771_), .Y(new_n8955_));
  XOR2X1   g08699(.A(new_n8955_), .B(new_n8769_), .Y(\f[69] ));
  OR2X1    g08700(.A(new_n8785_), .B(new_n8782_), .Y(new_n8957_));
  INVX1    g08701(.A(new_n8786_), .Y(new_n8958_));
  OAI21X1  g08702(.A0(new_n8952_), .A1(new_n8958_), .B0(new_n8957_), .Y(new_n8959_));
  OAI22X1  g08703(.A0(new_n467_), .A1(new_n7745_), .B0(new_n510_), .B1(new_n7772_), .Y(new_n8960_));
  AOI21X1  g08704(.A0(new_n7775_), .A1(new_n404_), .B0(new_n8960_), .Y(new_n8961_));
  XOR2X1   g08705(.A(new_n8961_), .B(\a[8] ), .Y(new_n8962_));
  XOR2X1   g08706(.A(new_n8962_), .B(new_n8959_), .Y(new_n8963_));
  AOI22X1  g08707(.A0(new_n603_), .A1(\b[61] ), .B0(new_n602_), .B1(\b[60] ), .Y(new_n8964_));
  OAI21X1  g08708(.A0(new_n601_), .A1(new_n7339_), .B0(new_n8964_), .Y(new_n8965_));
  AOI21X1  g08709(.A0(new_n7338_), .A1(new_n518_), .B0(new_n8965_), .Y(new_n8966_));
  XOR2X1   g08710(.A(new_n8966_), .B(\a[11] ), .Y(new_n8967_));
  INVX1    g08711(.A(new_n8967_), .Y(new_n8968_));
  NOR2X1   g08712(.A(new_n8950_), .B(new_n8948_), .Y(new_n8969_));
  AOI21X1  g08713(.A0(new_n8951_), .A1(new_n8943_), .B0(new_n8969_), .Y(new_n8970_));
  XOR2X1   g08714(.A(new_n8970_), .B(new_n8968_), .Y(new_n8971_));
  AOI21X1  g08715(.A0(new_n8790_), .A1(new_n8789_), .B0(new_n8795_), .Y(new_n8972_));
  INVX1    g08716(.A(new_n8972_), .Y(new_n8973_));
  OAI21X1  g08717(.A0(new_n8942_), .A1(new_n8796_), .B0(new_n8973_), .Y(new_n8974_));
  INVX1    g08718(.A(new_n816_), .Y(new_n8975_));
  OAI22X1  g08719(.A0(new_n875_), .A1(new_n6930_), .B0(new_n874_), .B1(new_n6933_), .Y(new_n8976_));
  AOI21X1  g08720(.A0(new_n8975_), .A1(\b[56] ), .B0(new_n8976_), .Y(new_n8977_));
  OAI21X1  g08721(.A0(new_n8540_), .A1(new_n751_), .B0(new_n8977_), .Y(new_n8978_));
  XOR2X1   g08722(.A(new_n8978_), .B(new_n665_), .Y(new_n8979_));
  INVX1    g08723(.A(new_n8979_), .Y(new_n8980_));
  XOR2X1   g08724(.A(new_n8980_), .B(new_n8974_), .Y(new_n8981_));
  INVX1    g08725(.A(new_n8981_), .Y(new_n8982_));
  AOI22X1  g08726(.A0(new_n1017_), .A1(\b[55] ), .B0(new_n1016_), .B1(\b[54] ), .Y(new_n8983_));
  OAI21X1  g08727(.A0(new_n1015_), .A1(new_n6151_), .B0(new_n8983_), .Y(new_n8984_));
  AOI21X1  g08728(.A0(new_n6150_), .A1(new_n882_), .B0(new_n8984_), .Y(new_n8985_));
  XOR2X1   g08729(.A(new_n8985_), .B(\a[17] ), .Y(new_n8986_));
  INVX1    g08730(.A(new_n8986_), .Y(new_n8987_));
  INVX1    g08731(.A(new_n8933_), .Y(new_n8988_));
  NOR2X1   g08732(.A(new_n8940_), .B(new_n8937_), .Y(new_n8989_));
  AOI21X1  g08733(.A0(new_n8941_), .A1(new_n8988_), .B0(new_n8989_), .Y(new_n8990_));
  XOR2X1   g08734(.A(new_n8990_), .B(new_n8987_), .Y(new_n8991_));
  AOI22X1  g08735(.A0(new_n1263_), .A1(\b[52] ), .B0(new_n1262_), .B1(\b[51] ), .Y(new_n8992_));
  OAI21X1  g08736(.A0(new_n1261_), .A1(new_n5234_), .B0(new_n8992_), .Y(new_n8993_));
  AOI21X1  g08737(.A0(new_n5590_), .A1(new_n1075_), .B0(new_n8993_), .Y(new_n8994_));
  XOR2X1   g08738(.A(new_n8994_), .B(\a[20] ), .Y(new_n8995_));
  NOR2X1   g08739(.A(new_n8803_), .B(new_n8800_), .Y(new_n8996_));
  AOI21X1  g08740(.A0(new_n8931_), .A1(new_n8804_), .B0(new_n8996_), .Y(new_n8997_));
  XOR2X1   g08741(.A(new_n8997_), .B(new_n8995_), .Y(new_n8998_));
  AOI22X1  g08742(.A0(new_n1526_), .A1(\b[49] ), .B0(new_n1525_), .B1(\b[48] ), .Y(new_n8999_));
  OAI21X1  g08743(.A0(new_n1524_), .A1(new_n5039_), .B0(new_n8999_), .Y(new_n9000_));
  AOI21X1  g08744(.A0(new_n5038_), .A1(new_n1347_), .B0(new_n9000_), .Y(new_n9001_));
  XOR2X1   g08745(.A(new_n9001_), .B(\a[23] ), .Y(new_n9002_));
  NOR2X1   g08746(.A(new_n8811_), .B(new_n8807_), .Y(new_n9003_));
  AOI21X1  g08747(.A0(new_n8930_), .A1(new_n8812_), .B0(new_n9003_), .Y(new_n9004_));
  XOR2X1   g08748(.A(new_n9004_), .B(new_n9002_), .Y(new_n9005_));
  AOI21X1  g08749(.A0(new_n8818_), .A1(new_n8817_), .B0(new_n8816_), .Y(new_n9006_));
  AOI21X1  g08750(.A0(new_n8929_), .A1(new_n8820_), .B0(new_n9006_), .Y(new_n9007_));
  INVX1    g08751(.A(new_n4509_), .Y(new_n9008_));
  OAI22X1  g08752(.A0(new_n1623_), .A1(new_n4693_), .B0(new_n1620_), .B1(new_n4674_), .Y(new_n9009_));
  AOI21X1  g08753(.A0(new_n1725_), .A1(\b[44] ), .B0(new_n9009_), .Y(new_n9010_));
  OAI21X1  g08754(.A0(new_n9008_), .A1(new_n1723_), .B0(new_n9010_), .Y(new_n9011_));
  XOR2X1   g08755(.A(new_n9011_), .B(new_n1621_), .Y(new_n9012_));
  XOR2X1   g08756(.A(new_n9012_), .B(new_n9007_), .Y(new_n9013_));
  AOI22X1  g08757(.A0(new_n2163_), .A1(\b[43] ), .B0(new_n2162_), .B1(\b[42] ), .Y(new_n9014_));
  OAI21X1  g08758(.A0(new_n2161_), .A1(new_n4015_), .B0(new_n9014_), .Y(new_n9015_));
  AOI21X1  g08759(.A0(new_n4014_), .A1(new_n1907_), .B0(new_n9015_), .Y(new_n9016_));
  XOR2X1   g08760(.A(new_n9016_), .B(\a[29] ), .Y(new_n9017_));
  NOR2X1   g08761(.A(new_n8927_), .B(new_n8924_), .Y(new_n9018_));
  AOI21X1  g08762(.A0(new_n8928_), .A1(new_n8920_), .B0(new_n9018_), .Y(new_n9019_));
  XOR2X1   g08763(.A(new_n9019_), .B(new_n9017_), .Y(new_n9020_));
  AOI22X1  g08764(.A0(new_n2545_), .A1(\b[40] ), .B0(new_n2544_), .B1(\b[39] ), .Y(new_n9021_));
  OAI21X1  g08765(.A0(new_n2543_), .A1(new_n3575_), .B0(new_n9021_), .Y(new_n9022_));
  AOI21X1  g08766(.A0(new_n3574_), .A1(new_n2260_), .B0(new_n9022_), .Y(new_n9023_));
  XOR2X1   g08767(.A(new_n9023_), .B(\a[32] ), .Y(new_n9024_));
  NOR2X1   g08768(.A(new_n8918_), .B(new_n8914_), .Y(new_n9025_));
  AOI21X1  g08769(.A0(new_n8919_), .A1(new_n8823_), .B0(new_n9025_), .Y(new_n9026_));
  XOR2X1   g08770(.A(new_n9026_), .B(new_n9024_), .Y(new_n9027_));
  AOI22X1  g08771(.A0(new_n2813_), .A1(\b[37] ), .B0(new_n2812_), .B1(\b[36] ), .Y(new_n9028_));
  OAI21X1  g08772(.A0(new_n2946_), .A1(new_n3156_), .B0(new_n9028_), .Y(new_n9029_));
  AOI21X1  g08773(.A0(new_n3155_), .A1(new_n2652_), .B0(new_n9029_), .Y(new_n9030_));
  XOR2X1   g08774(.A(new_n9030_), .B(\a[35] ), .Y(new_n9031_));
  INVX1    g08775(.A(new_n8826_), .Y(new_n9032_));
  INVX1    g08776(.A(new_n8912_), .Y(new_n9033_));
  NAND2X1  g08777(.A(new_n9033_), .B(new_n8908_), .Y(new_n9034_));
  OAI21X1  g08778(.A0(new_n8913_), .A1(new_n9032_), .B0(new_n9034_), .Y(new_n9035_));
  AOI22X1  g08779(.A0(new_n3204_), .A1(\b[34] ), .B0(new_n3203_), .B1(\b[33] ), .Y(new_n9036_));
  OAI21X1  g08780(.A0(new_n3321_), .A1(new_n2612_), .B0(new_n9036_), .Y(new_n9037_));
  AOI21X1  g08781(.A0(new_n3080_), .A1(new_n2759_), .B0(new_n9037_), .Y(new_n9038_));
  XOR2X1   g08782(.A(new_n9038_), .B(new_n3078_), .Y(new_n9039_));
  AND2X1   g08783(.A(new_n8849_), .B(new_n8845_), .Y(new_n9040_));
  INVX1    g08784(.A(new_n9040_), .Y(new_n9041_));
  OAI21X1  g08785(.A0(new_n8854_), .A1(new_n8850_), .B0(new_n9041_), .Y(new_n9042_));
  OR2X1    g08786(.A(\a[5] ), .B(\a[2] ), .Y(new_n9043_));
  OAI21X1  g08787(.A0(new_n8848_), .A1(new_n8847_), .B0(new_n9043_), .Y(new_n9044_));
  AOI22X1  g08788(.A0(new_n7818_), .A1(\b[6] ), .B0(new_n7817_), .B1(\b[7] ), .Y(new_n9045_));
  INVX1    g08789(.A(new_n9045_), .Y(new_n9046_));
  XOR2X1   g08790(.A(new_n9046_), .B(new_n9044_), .Y(new_n9047_));
  AOI22X1  g08791(.A0(new_n7192_), .A1(\b[10] ), .B0(new_n7189_), .B1(\b[9] ), .Y(new_n9048_));
  OAI21X1  g08792(.A0(new_n7627_), .A1(new_n489_), .B0(new_n9048_), .Y(new_n9049_));
  AOI21X1  g08793(.A0(new_n7187_), .A1(new_n543_), .B0(new_n9049_), .Y(new_n9050_));
  XOR2X1   g08794(.A(new_n9050_), .B(\a[62] ), .Y(new_n9051_));
  XOR2X1   g08795(.A(new_n9051_), .B(new_n9047_), .Y(new_n9052_));
  XOR2X1   g08796(.A(new_n9052_), .B(new_n9042_), .Y(new_n9053_));
  AOI22X1  g08797(.A0(new_n6603_), .A1(\b[13] ), .B0(new_n6600_), .B1(\b[12] ), .Y(new_n9054_));
  OAI21X1  g08798(.A0(new_n6804_), .A1(new_n716_), .B0(new_n9054_), .Y(new_n9055_));
  AOI21X1  g08799(.A0(new_n6598_), .A1(new_n715_), .B0(new_n9055_), .Y(new_n9056_));
  XOR2X1   g08800(.A(new_n9056_), .B(\a[59] ), .Y(new_n9057_));
  XOR2X1   g08801(.A(new_n9057_), .B(new_n9053_), .Y(new_n9058_));
  INVX1    g08802(.A(new_n8843_), .Y(new_n9059_));
  AND2X1   g08803(.A(new_n8855_), .B(new_n9059_), .Y(new_n9060_));
  INVX1    g08804(.A(new_n8856_), .Y(new_n9061_));
  AOI21X1  g08805(.A0(new_n9061_), .A1(new_n8839_), .B0(new_n9060_), .Y(new_n9062_));
  XOR2X1   g08806(.A(new_n9062_), .B(new_n9058_), .Y(new_n9063_));
  AOI22X1  g08807(.A0(new_n6438_), .A1(\b[16] ), .B0(new_n6437_), .B1(\b[15] ), .Y(new_n9064_));
  OAI21X1  g08808(.A0(new_n6436_), .A1(new_n792_), .B0(new_n9064_), .Y(new_n9065_));
  AOI21X1  g08809(.A0(new_n6023_), .A1(new_n842_), .B0(new_n9065_), .Y(new_n9066_));
  XOR2X1   g08810(.A(new_n9066_), .B(\a[56] ), .Y(new_n9067_));
  XOR2X1   g08811(.A(new_n9067_), .B(new_n9063_), .Y(new_n9068_));
  INVX1    g08812(.A(new_n9068_), .Y(new_n9069_));
  OR2X1    g08813(.A(new_n8861_), .B(new_n8857_), .Y(new_n9070_));
  OAI21X1  g08814(.A0(new_n8866_), .A1(new_n8863_), .B0(new_n9070_), .Y(new_n9071_));
  XOR2X1   g08815(.A(new_n9071_), .B(new_n9069_), .Y(new_n9072_));
  AOI22X1  g08816(.A0(new_n5430_), .A1(\b[19] ), .B0(new_n5427_), .B1(\b[18] ), .Y(new_n9073_));
  OAI21X1  g08817(.A0(new_n5891_), .A1(new_n1118_), .B0(new_n9073_), .Y(new_n9074_));
  AOI21X1  g08818(.A0(new_n5425_), .A1(new_n1117_), .B0(new_n9074_), .Y(new_n9075_));
  XOR2X1   g08819(.A(new_n9075_), .B(\a[53] ), .Y(new_n9076_));
  XOR2X1   g08820(.A(new_n9076_), .B(new_n9072_), .Y(new_n9077_));
  INVX1    g08821(.A(new_n8871_), .Y(new_n9078_));
  NOR2X1   g08822(.A(new_n8875_), .B(new_n8872_), .Y(new_n9079_));
  AOI21X1  g08823(.A0(new_n9078_), .A1(new_n8867_), .B0(new_n9079_), .Y(new_n9080_));
  XOR2X1   g08824(.A(new_n9080_), .B(new_n9077_), .Y(new_n9081_));
  AOI22X1  g08825(.A0(new_n4880_), .A1(\b[22] ), .B0(new_n4877_), .B1(\b[21] ), .Y(new_n9082_));
  OAI21X1  g08826(.A0(new_n5291_), .A1(new_n1297_), .B0(new_n9082_), .Y(new_n9083_));
  AOI21X1  g08827(.A0(new_n4875_), .A1(new_n1399_), .B0(new_n9083_), .Y(new_n9084_));
  XOR2X1   g08828(.A(new_n9084_), .B(\a[50] ), .Y(new_n9085_));
  XOR2X1   g08829(.A(new_n9085_), .B(new_n9081_), .Y(new_n9086_));
  XOR2X1   g08830(.A(new_n8879_), .B(new_n4873_), .Y(new_n9087_));
  AND2X1   g08831(.A(new_n9087_), .B(new_n8876_), .Y(new_n9088_));
  INVX1    g08832(.A(new_n8881_), .Y(new_n9089_));
  AOI21X1  g08833(.A0(new_n9089_), .A1(new_n8837_), .B0(new_n9088_), .Y(new_n9090_));
  XOR2X1   g08834(.A(new_n9090_), .B(new_n9086_), .Y(new_n9091_));
  AOI22X1  g08835(.A0(new_n4572_), .A1(\b[25] ), .B0(new_n4571_), .B1(\b[24] ), .Y(new_n9092_));
  OAI21X1  g08836(.A0(new_n4740_), .A1(new_n1591_), .B0(new_n9092_), .Y(new_n9093_));
  AOI21X1  g08837(.A0(new_n4375_), .A1(new_n1590_), .B0(new_n9093_), .Y(new_n9094_));
  XOR2X1   g08838(.A(new_n9094_), .B(\a[47] ), .Y(new_n9095_));
  XOR2X1   g08839(.A(new_n9095_), .B(new_n9091_), .Y(new_n9096_));
  NOR2X1   g08840(.A(new_n8886_), .B(new_n8882_), .Y(new_n9097_));
  AOI21X1  g08841(.A0(new_n8887_), .A1(new_n8835_), .B0(new_n9097_), .Y(new_n9098_));
  XOR2X1   g08842(.A(new_n9098_), .B(new_n9096_), .Y(new_n9099_));
  AOI22X1  g08843(.A0(new_n4095_), .A1(\b[28] ), .B0(new_n4094_), .B1(\b[27] ), .Y(new_n9100_));
  OAI21X1  g08844(.A0(new_n4233_), .A1(new_n1877_), .B0(new_n9100_), .Y(new_n9101_));
  AOI21X1  g08845(.A0(new_n3901_), .A1(new_n2004_), .B0(new_n9101_), .Y(new_n9102_));
  XOR2X1   g08846(.A(new_n9102_), .B(\a[44] ), .Y(new_n9103_));
  XOR2X1   g08847(.A(new_n9103_), .B(new_n9099_), .Y(new_n9104_));
  INVX1    g08848(.A(new_n9104_), .Y(new_n9105_));
  INVX1    g08849(.A(new_n8892_), .Y(new_n9106_));
  NOR2X1   g08850(.A(new_n8896_), .B(new_n8893_), .Y(new_n9107_));
  AOI21X1  g08851(.A0(new_n9106_), .A1(new_n8888_), .B0(new_n9107_), .Y(new_n9108_));
  XOR2X1   g08852(.A(new_n9108_), .B(new_n9105_), .Y(new_n9109_));
  AOI22X1  g08853(.A0(new_n3652_), .A1(\b[31] ), .B0(new_n3651_), .B1(\b[30] ), .Y(new_n9110_));
  OAI21X1  g08854(.A0(new_n3778_), .A1(new_n2359_), .B0(new_n9110_), .Y(new_n9111_));
  AOI21X1  g08855(.A0(new_n3480_), .A1(new_n2358_), .B0(new_n9111_), .Y(new_n9112_));
  XOR2X1   g08856(.A(new_n9112_), .B(\a[41] ), .Y(new_n9113_));
  XOR2X1   g08857(.A(new_n9113_), .B(new_n9109_), .Y(new_n9114_));
  XOR2X1   g08858(.A(new_n9114_), .B(new_n8907_), .Y(new_n9115_));
  XOR2X1   g08859(.A(new_n9115_), .B(new_n9039_), .Y(new_n9116_));
  XOR2X1   g08860(.A(new_n9116_), .B(new_n9035_), .Y(new_n9117_));
  XOR2X1   g08861(.A(new_n9117_), .B(new_n9031_), .Y(new_n9118_));
  XOR2X1   g08862(.A(new_n9118_), .B(new_n9027_), .Y(new_n9119_));
  XOR2X1   g08863(.A(new_n9119_), .B(new_n9020_), .Y(new_n9120_));
  XOR2X1   g08864(.A(new_n9120_), .B(new_n9013_), .Y(new_n9121_));
  XOR2X1   g08865(.A(new_n9121_), .B(new_n9005_), .Y(new_n9122_));
  XOR2X1   g08866(.A(new_n9122_), .B(new_n8998_), .Y(new_n9123_));
  XOR2X1   g08867(.A(new_n9123_), .B(new_n8991_), .Y(new_n9124_));
  XOR2X1   g08868(.A(new_n9124_), .B(new_n8982_), .Y(new_n9125_));
  XOR2X1   g08869(.A(new_n9125_), .B(new_n8971_), .Y(new_n9126_));
  INVX1    g08870(.A(new_n9126_), .Y(new_n9127_));
  XOR2X1   g08871(.A(new_n9127_), .B(new_n8963_), .Y(new_n9128_));
  NOR2X1   g08872(.A(new_n8777_), .B(new_n8773_), .Y(new_n9129_));
  INVX1    g08873(.A(new_n8953_), .Y(new_n9130_));
  AOI21X1  g08874(.A0(new_n9130_), .A1(new_n8778_), .B0(new_n9129_), .Y(new_n9131_));
  XOR2X1   g08875(.A(new_n9131_), .B(new_n9128_), .Y(new_n9132_));
  OR2X1    g08876(.A(new_n8954_), .B(new_n8771_), .Y(new_n9133_));
  OAI21X1  g08877(.A0(new_n8768_), .A1(new_n8767_), .B0(new_n8955_), .Y(new_n9134_));
  AND2X1   g08878(.A(new_n9134_), .B(new_n9133_), .Y(new_n9135_));
  XOR2X1   g08879(.A(new_n9135_), .B(new_n9132_), .Y(\f[70] ));
  INVX1    g08880(.A(new_n9128_), .Y(new_n9137_));
  NOR2X1   g08881(.A(new_n9131_), .B(new_n9137_), .Y(new_n9138_));
  AOI21X1  g08882(.A0(new_n9134_), .A1(new_n9133_), .B0(new_n9132_), .Y(new_n9139_));
  OR2X1    g08883(.A(new_n9139_), .B(new_n9138_), .Y(new_n9140_));
  INVX1    g08884(.A(new_n8962_), .Y(new_n9141_));
  NOR2X1   g08885(.A(new_n9127_), .B(new_n8963_), .Y(new_n9142_));
  AOI21X1  g08886(.A0(new_n9141_), .A1(new_n8959_), .B0(new_n9142_), .Y(new_n9143_));
  OR2X1    g08887(.A(new_n8970_), .B(new_n8967_), .Y(new_n9144_));
  OAI21X1  g08888(.A0(new_n9125_), .A1(new_n8971_), .B0(new_n9144_), .Y(new_n9145_));
  AOI22X1  g08889(.A0(new_n7774_), .A1(new_n404_), .B0(new_n8551_), .B1(\b[63] ), .Y(new_n9146_));
  XOR2X1   g08890(.A(new_n9146_), .B(\a[8] ), .Y(new_n9147_));
  INVX1    g08891(.A(new_n9147_), .Y(new_n9148_));
  XOR2X1   g08892(.A(new_n9148_), .B(new_n9145_), .Y(new_n9149_));
  AOI22X1  g08893(.A0(new_n1017_), .A1(\b[56] ), .B0(new_n1016_), .B1(\b[55] ), .Y(new_n9150_));
  OAI21X1  g08894(.A0(new_n1015_), .A1(new_n6148_), .B0(new_n9150_), .Y(new_n9151_));
  AOI21X1  g08895(.A0(new_n6342_), .A1(new_n882_), .B0(new_n9151_), .Y(new_n9152_));
  XOR2X1   g08896(.A(new_n9152_), .B(\a[17] ), .Y(new_n9153_));
  NOR2X1   g08897(.A(new_n8997_), .B(new_n8995_), .Y(new_n9154_));
  INVX1    g08898(.A(new_n9122_), .Y(new_n9155_));
  AOI21X1  g08899(.A0(new_n9155_), .A1(new_n8998_), .B0(new_n9154_), .Y(new_n9156_));
  XOR2X1   g08900(.A(new_n9156_), .B(new_n9153_), .Y(new_n9157_));
  AOI22X1  g08901(.A0(new_n1526_), .A1(\b[50] ), .B0(new_n1525_), .B1(\b[49] ), .Y(new_n9158_));
  OAI21X1  g08902(.A0(new_n1524_), .A1(new_n5036_), .B0(new_n9158_), .Y(new_n9159_));
  AOI21X1  g08903(.A0(new_n5204_), .A1(new_n1347_), .B0(new_n9159_), .Y(new_n9160_));
  XOR2X1   g08904(.A(new_n9160_), .B(\a[23] ), .Y(new_n9161_));
  NOR2X1   g08905(.A(new_n9012_), .B(new_n9007_), .Y(new_n9162_));
  INVX1    g08906(.A(new_n9120_), .Y(new_n9163_));
  AOI21X1  g08907(.A0(new_n9163_), .A1(new_n9013_), .B0(new_n9162_), .Y(new_n9164_));
  XOR2X1   g08908(.A(new_n9164_), .B(new_n9161_), .Y(new_n9165_));
  AOI22X1  g08909(.A0(new_n1814_), .A1(\b[47] ), .B0(new_n1813_), .B1(\b[46] ), .Y(new_n9166_));
  OAI21X1  g08910(.A0(new_n1812_), .A1(new_n4674_), .B0(new_n9166_), .Y(new_n9167_));
  AOI21X1  g08911(.A0(new_n4673_), .A1(new_n1617_), .B0(new_n9167_), .Y(new_n9168_));
  XOR2X1   g08912(.A(new_n9168_), .B(\a[26] ), .Y(new_n9169_));
  NOR2X1   g08913(.A(new_n9019_), .B(new_n9017_), .Y(new_n9170_));
  INVX1    g08914(.A(new_n9119_), .Y(new_n9171_));
  AOI21X1  g08915(.A0(new_n9171_), .A1(new_n9020_), .B0(new_n9170_), .Y(new_n9172_));
  XOR2X1   g08916(.A(new_n9172_), .B(new_n9169_), .Y(new_n9173_));
  AOI22X1  g08917(.A0(new_n2545_), .A1(\b[41] ), .B0(new_n2544_), .B1(\b[40] ), .Y(new_n9174_));
  OAI21X1  g08918(.A0(new_n2543_), .A1(new_n3723_), .B0(new_n9174_), .Y(new_n9175_));
  AOI21X1  g08919(.A0(new_n3722_), .A1(new_n2260_), .B0(new_n9175_), .Y(new_n9176_));
  XOR2X1   g08920(.A(new_n9176_), .B(\a[32] ), .Y(new_n9177_));
  INVX1    g08921(.A(new_n9031_), .Y(new_n9178_));
  AND2X1   g08922(.A(new_n9116_), .B(new_n9035_), .Y(new_n9179_));
  AOI21X1  g08923(.A0(new_n9117_), .A1(new_n9178_), .B0(new_n9179_), .Y(new_n9180_));
  XOR2X1   g08924(.A(new_n9180_), .B(new_n9177_), .Y(new_n9181_));
  NOR2X1   g08925(.A(new_n9080_), .B(new_n9077_), .Y(new_n9182_));
  INVX1    g08926(.A(new_n9182_), .Y(new_n9183_));
  INVX1    g08927(.A(new_n9081_), .Y(new_n9184_));
  OAI21X1  g08928(.A0(new_n9085_), .A1(new_n9184_), .B0(new_n9183_), .Y(new_n9185_));
  AOI22X1  g08929(.A0(new_n4880_), .A1(\b[23] ), .B0(new_n4877_), .B1(\b[22] ), .Y(new_n9186_));
  OAI21X1  g08930(.A0(new_n5291_), .A1(new_n1482_), .B0(new_n9186_), .Y(new_n9187_));
  AOI21X1  g08931(.A0(new_n4875_), .A1(new_n1481_), .B0(new_n9187_), .Y(new_n9188_));
  XOR2X1   g08932(.A(new_n9188_), .B(\a[50] ), .Y(new_n9189_));
  AND2X1   g08933(.A(new_n9071_), .B(new_n9069_), .Y(new_n9190_));
  INVX1    g08934(.A(new_n9190_), .Y(new_n9191_));
  INVX1    g08935(.A(new_n9072_), .Y(new_n9192_));
  OAI21X1  g08936(.A0(new_n9076_), .A1(new_n9192_), .B0(new_n9191_), .Y(new_n9193_));
  INVX1    g08937(.A(new_n9193_), .Y(new_n9194_));
  AND2X1   g08938(.A(new_n9052_), .B(new_n9042_), .Y(new_n9195_));
  INVX1    g08939(.A(new_n9195_), .Y(new_n9196_));
  INVX1    g08940(.A(new_n9053_), .Y(new_n9197_));
  OAI21X1  g08941(.A0(new_n9057_), .A1(new_n9197_), .B0(new_n9196_), .Y(new_n9198_));
  NOR2X1   g08942(.A(new_n9051_), .B(new_n9047_), .Y(new_n9199_));
  AOI21X1  g08943(.A0(new_n9045_), .A1(new_n9044_), .B0(new_n9199_), .Y(new_n9200_));
  AOI22X1  g08944(.A0(new_n7818_), .A1(\b[7] ), .B0(new_n7817_), .B1(\b[8] ), .Y(new_n9201_));
  INVX1    g08945(.A(new_n9201_), .Y(new_n9202_));
  AND2X1   g08946(.A(new_n9202_), .B(new_n9045_), .Y(new_n9203_));
  XOR2X1   g08947(.A(new_n9201_), .B(new_n9046_), .Y(new_n9204_));
  OR2X1    g08948(.A(new_n9202_), .B(new_n9045_), .Y(new_n9205_));
  OAI21X1  g08949(.A0(new_n9203_), .A1(new_n9200_), .B0(new_n9205_), .Y(new_n9206_));
  OAI22X1  g08950(.A0(new_n9206_), .A1(new_n9203_), .B0(new_n9204_), .B1(new_n9200_), .Y(new_n9207_));
  AOI22X1  g08951(.A0(new_n7192_), .A1(\b[11] ), .B0(new_n7189_), .B1(\b[10] ), .Y(new_n9208_));
  OAI21X1  g08952(.A0(new_n7627_), .A1(new_n590_), .B0(new_n9208_), .Y(new_n9209_));
  AOI21X1  g08953(.A0(new_n7187_), .A1(new_n589_), .B0(new_n9209_), .Y(new_n9210_));
  XOR2X1   g08954(.A(new_n9210_), .B(\a[62] ), .Y(new_n9211_));
  XOR2X1   g08955(.A(new_n9211_), .B(new_n9207_), .Y(new_n9212_));
  AOI22X1  g08956(.A0(new_n6603_), .A1(\b[14] ), .B0(new_n6600_), .B1(\b[13] ), .Y(new_n9213_));
  OAI21X1  g08957(.A0(new_n6804_), .A1(new_n713_), .B0(new_n9213_), .Y(new_n9214_));
  AOI21X1  g08958(.A0(new_n6598_), .A1(new_n734_), .B0(new_n9214_), .Y(new_n9215_));
  XOR2X1   g08959(.A(new_n9215_), .B(\a[59] ), .Y(new_n9216_));
  XOR2X1   g08960(.A(new_n9216_), .B(new_n9212_), .Y(new_n9217_));
  XOR2X1   g08961(.A(new_n9217_), .B(new_n9198_), .Y(new_n9218_));
  AOI22X1  g08962(.A0(new_n6438_), .A1(\b[17] ), .B0(new_n6437_), .B1(\b[16] ), .Y(new_n9219_));
  OAI21X1  g08963(.A0(new_n6436_), .A1(new_n977_), .B0(new_n9219_), .Y(new_n9220_));
  AOI21X1  g08964(.A0(new_n6023_), .A1(new_n976_), .B0(new_n9220_), .Y(new_n9221_));
  XOR2X1   g08965(.A(new_n9221_), .B(\a[56] ), .Y(new_n9222_));
  XOR2X1   g08966(.A(new_n9222_), .B(new_n9218_), .Y(new_n9223_));
  INVX1    g08967(.A(new_n9223_), .Y(new_n9224_));
  NOR2X1   g08968(.A(new_n9062_), .B(new_n9058_), .Y(new_n9225_));
  INVX1    g08969(.A(new_n9067_), .Y(new_n9226_));
  AOI21X1  g08970(.A0(new_n9226_), .A1(new_n9063_), .B0(new_n9225_), .Y(new_n9227_));
  XOR2X1   g08971(.A(new_n9227_), .B(new_n9224_), .Y(new_n9228_));
  AOI22X1  g08972(.A0(new_n5430_), .A1(\b[20] ), .B0(new_n5427_), .B1(\b[19] ), .Y(new_n9229_));
  OAI21X1  g08973(.A0(new_n5891_), .A1(new_n1115_), .B0(new_n9229_), .Y(new_n9230_));
  AOI21X1  g08974(.A0(new_n5425_), .A1(new_n1217_), .B0(new_n9230_), .Y(new_n9231_));
  XOR2X1   g08975(.A(new_n9231_), .B(\a[53] ), .Y(new_n9232_));
  XOR2X1   g08976(.A(new_n9232_), .B(new_n9228_), .Y(new_n9233_));
  XOR2X1   g08977(.A(new_n9233_), .B(new_n9194_), .Y(new_n9234_));
  XOR2X1   g08978(.A(new_n9234_), .B(new_n9189_), .Y(new_n9235_));
  XOR2X1   g08979(.A(new_n9235_), .B(new_n9185_), .Y(new_n9236_));
  AOI22X1  g08980(.A0(new_n4572_), .A1(\b[26] ), .B0(new_n4571_), .B1(\b[25] ), .Y(new_n9237_));
  OAI21X1  g08981(.A0(new_n4740_), .A1(new_n1588_), .B0(new_n9237_), .Y(new_n9238_));
  AOI21X1  g08982(.A0(new_n4375_), .A1(new_n1783_), .B0(new_n9238_), .Y(new_n9239_));
  XOR2X1   g08983(.A(new_n9239_), .B(\a[47] ), .Y(new_n9240_));
  XOR2X1   g08984(.A(new_n9240_), .B(new_n9236_), .Y(new_n9241_));
  NOR2X1   g08985(.A(new_n9090_), .B(new_n9086_), .Y(new_n9242_));
  INVX1    g08986(.A(new_n9095_), .Y(new_n9243_));
  AOI21X1  g08987(.A0(new_n9243_), .A1(new_n9091_), .B0(new_n9242_), .Y(new_n9244_));
  XOR2X1   g08988(.A(new_n9244_), .B(new_n9241_), .Y(new_n9245_));
  AOI22X1  g08989(.A0(new_n4095_), .A1(\b[29] ), .B0(new_n4094_), .B1(\b[28] ), .Y(new_n9246_));
  OAI21X1  g08990(.A0(new_n4233_), .A1(new_n2126_), .B0(new_n9246_), .Y(new_n9247_));
  AOI21X1  g08991(.A0(new_n3901_), .A1(new_n2125_), .B0(new_n9247_), .Y(new_n9248_));
  XOR2X1   g08992(.A(new_n9248_), .B(\a[44] ), .Y(new_n9249_));
  XOR2X1   g08993(.A(new_n9249_), .B(new_n9245_), .Y(new_n9250_));
  NOR2X1   g08994(.A(new_n9098_), .B(new_n9096_), .Y(new_n9251_));
  INVX1    g08995(.A(new_n9103_), .Y(new_n9252_));
  AOI21X1  g08996(.A0(new_n9252_), .A1(new_n9099_), .B0(new_n9251_), .Y(new_n9253_));
  XOR2X1   g08997(.A(new_n9253_), .B(new_n9250_), .Y(new_n9254_));
  INVX1    g08998(.A(new_n9254_), .Y(new_n9255_));
  AOI22X1  g08999(.A0(new_n3652_), .A1(\b[32] ), .B0(new_n3651_), .B1(\b[31] ), .Y(new_n9256_));
  OAI21X1  g09000(.A0(new_n3778_), .A1(new_n2356_), .B0(new_n9256_), .Y(new_n9257_));
  AOI21X1  g09001(.A0(new_n3480_), .A1(new_n2495_), .B0(new_n9257_), .Y(new_n9258_));
  XOR2X1   g09002(.A(new_n9258_), .B(\a[41] ), .Y(new_n9259_));
  XOR2X1   g09003(.A(new_n9259_), .B(new_n9255_), .Y(new_n9260_));
  INVX1    g09004(.A(new_n9260_), .Y(new_n9261_));
  OR2X1    g09005(.A(new_n9108_), .B(new_n9104_), .Y(new_n9262_));
  OR2X1    g09006(.A(new_n9113_), .B(new_n9109_), .Y(new_n9263_));
  AND2X1   g09007(.A(new_n9263_), .B(new_n9262_), .Y(new_n9264_));
  XOR2X1   g09008(.A(new_n9264_), .B(new_n9261_), .Y(new_n9265_));
  AOI22X1  g09009(.A0(new_n3204_), .A1(\b[35] ), .B0(new_n3203_), .B1(\b[34] ), .Y(new_n9266_));
  OAI21X1  g09010(.A0(new_n3321_), .A1(new_n2893_), .B0(new_n9266_), .Y(new_n9267_));
  AOI21X1  g09011(.A0(new_n3080_), .A1(new_n2892_), .B0(new_n9267_), .Y(new_n9268_));
  XOR2X1   g09012(.A(new_n9268_), .B(\a[38] ), .Y(new_n9269_));
  XOR2X1   g09013(.A(new_n9269_), .B(new_n9265_), .Y(new_n9270_));
  INVX1    g09014(.A(new_n9270_), .Y(new_n9271_));
  AND2X1   g09015(.A(new_n9114_), .B(new_n8907_), .Y(new_n9272_));
  AOI21X1  g09016(.A0(new_n9115_), .A1(new_n9039_), .B0(new_n9272_), .Y(new_n9273_));
  XOR2X1   g09017(.A(new_n9273_), .B(new_n9271_), .Y(new_n9274_));
  AOI22X1  g09018(.A0(new_n2813_), .A1(\b[38] ), .B0(new_n2812_), .B1(\b[37] ), .Y(new_n9275_));
  OAI21X1  g09019(.A0(new_n2946_), .A1(new_n3276_), .B0(new_n9275_), .Y(new_n9276_));
  AOI21X1  g09020(.A0(new_n3275_), .A1(new_n2652_), .B0(new_n9276_), .Y(new_n9277_));
  XOR2X1   g09021(.A(new_n9277_), .B(\a[35] ), .Y(new_n9278_));
  XOR2X1   g09022(.A(new_n9278_), .B(new_n9274_), .Y(new_n9279_));
  XOR2X1   g09023(.A(new_n9279_), .B(new_n9181_), .Y(new_n9280_));
  NOR2X1   g09024(.A(new_n9026_), .B(new_n9024_), .Y(new_n9281_));
  INVX1    g09025(.A(new_n9281_), .Y(new_n9282_));
  INVX1    g09026(.A(new_n9027_), .Y(new_n9283_));
  OAI21X1  g09027(.A0(new_n9118_), .A1(new_n9283_), .B0(new_n9282_), .Y(new_n9284_));
  OAI22X1  g09028(.A0(new_n1913_), .A1(new_n4336_), .B0(new_n1910_), .B1(new_n4339_), .Y(new_n9285_));
  AOI21X1  g09029(.A0(new_n2045_), .A1(\b[42] ), .B0(new_n9285_), .Y(new_n9286_));
  OAI21X1  g09030(.A0(new_n8736_), .A1(new_n2043_), .B0(new_n9286_), .Y(new_n9287_));
  XOR2X1   g09031(.A(new_n9287_), .B(new_n1911_), .Y(new_n9288_));
  XOR2X1   g09032(.A(new_n9288_), .B(new_n9284_), .Y(new_n9289_));
  XOR2X1   g09033(.A(new_n9289_), .B(new_n9280_), .Y(new_n9290_));
  XOR2X1   g09034(.A(new_n9290_), .B(new_n9173_), .Y(new_n9291_));
  INVX1    g09035(.A(new_n9291_), .Y(new_n9292_));
  XOR2X1   g09036(.A(new_n9292_), .B(new_n9165_), .Y(new_n9293_));
  NOR2X1   g09037(.A(new_n9004_), .B(new_n9002_), .Y(new_n9294_));
  INVX1    g09038(.A(new_n9121_), .Y(new_n9295_));
  AOI21X1  g09039(.A0(new_n9295_), .A1(new_n9005_), .B0(new_n9294_), .Y(new_n9296_));
  OAI22X1  g09040(.A0(new_n1080_), .A1(new_n6151_), .B0(new_n1078_), .B1(new_n5808_), .Y(new_n9297_));
  AOI21X1  g09041(.A0(new_n1167_), .A1(\b[51] ), .B0(new_n9297_), .Y(new_n9298_));
  OAI21X1  g09042(.A0(new_n8599_), .A1(new_n1165_), .B0(new_n9298_), .Y(new_n9299_));
  XOR2X1   g09043(.A(new_n9299_), .B(new_n1072_), .Y(new_n9300_));
  INVX1    g09044(.A(new_n9300_), .Y(new_n9301_));
  XOR2X1   g09045(.A(new_n9301_), .B(new_n9296_), .Y(new_n9302_));
  XOR2X1   g09046(.A(new_n9302_), .B(new_n9293_), .Y(new_n9303_));
  XOR2X1   g09047(.A(new_n9303_), .B(new_n9157_), .Y(new_n9304_));
  AOI22X1  g09048(.A0(new_n818_), .A1(\b[59] ), .B0(new_n817_), .B1(\b[58] ), .Y(new_n9305_));
  OAI21X1  g09049(.A0(new_n816_), .A1(new_n6933_), .B0(new_n9305_), .Y(new_n9306_));
  AOI21X1  g09050(.A0(new_n6932_), .A1(new_n668_), .B0(new_n9306_), .Y(new_n9307_));
  XOR2X1   g09051(.A(new_n9307_), .B(\a[14] ), .Y(new_n9308_));
  OR2X1    g09052(.A(new_n8990_), .B(new_n8986_), .Y(new_n9309_));
  OR2X1    g09053(.A(new_n9123_), .B(new_n8991_), .Y(new_n9310_));
  AND2X1   g09054(.A(new_n9310_), .B(new_n9309_), .Y(new_n9311_));
  XOR2X1   g09055(.A(new_n9311_), .B(new_n9308_), .Y(new_n9312_));
  XOR2X1   g09056(.A(new_n9312_), .B(new_n9304_), .Y(new_n9313_));
  INVX1    g09057(.A(new_n9313_), .Y(new_n9314_));
  OAI22X1  g09058(.A0(new_n661_), .A1(new_n7745_), .B0(new_n660_), .B1(new_n7748_), .Y(new_n9315_));
  AOI21X1  g09059(.A0(new_n8541_), .A1(\b[60] ), .B0(new_n9315_), .Y(new_n9316_));
  OAI21X1  g09060(.A0(new_n8753_), .A1(new_n567_), .B0(new_n9316_), .Y(new_n9317_));
  XOR2X1   g09061(.A(new_n9317_), .B(new_n515_), .Y(new_n9318_));
  AND2X1   g09062(.A(new_n8980_), .B(new_n8974_), .Y(new_n9319_));
  AOI21X1  g09063(.A0(new_n9124_), .A1(new_n8981_), .B0(new_n9319_), .Y(new_n9320_));
  NOR2X1   g09064(.A(new_n9318_), .B(new_n9320_), .Y(new_n9321_));
  OR2X1    g09065(.A(new_n9321_), .B(new_n9318_), .Y(new_n9322_));
  XOR2X1   g09066(.A(new_n9318_), .B(new_n9320_), .Y(new_n9323_));
  INVX1    g09067(.A(new_n9320_), .Y(new_n9324_));
  AOI21X1  g09068(.A0(new_n9318_), .A1(new_n9324_), .B0(new_n9314_), .Y(new_n9325_));
  AOI22X1  g09069(.A0(new_n9325_), .A1(new_n9322_), .B0(new_n9323_), .B1(new_n9314_), .Y(new_n9326_));
  XOR2X1   g09070(.A(new_n9326_), .B(new_n9149_), .Y(new_n9327_));
  INVX1    g09071(.A(new_n9327_), .Y(new_n9328_));
  XOR2X1   g09072(.A(new_n9328_), .B(new_n9143_), .Y(new_n9329_));
  XOR2X1   g09073(.A(new_n9329_), .B(new_n9140_), .Y(\f[71] ));
  OR2X1    g09074(.A(new_n9328_), .B(new_n9143_), .Y(new_n9331_));
  OAI21X1  g09075(.A0(new_n9139_), .A1(new_n9138_), .B0(new_n9329_), .Y(new_n9332_));
  AND2X1   g09076(.A(new_n9332_), .B(new_n9331_), .Y(new_n9333_));
  AND2X1   g09077(.A(new_n9148_), .B(new_n9145_), .Y(new_n9334_));
  AOI21X1  g09078(.A0(new_n9326_), .A1(new_n9149_), .B0(new_n9334_), .Y(new_n9335_));
  AOI21X1  g09079(.A0(new_n9323_), .A1(new_n9314_), .B0(new_n9321_), .Y(new_n9336_));
  AOI22X1  g09080(.A0(new_n603_), .A1(\b[63] ), .B0(new_n602_), .B1(\b[62] ), .Y(new_n9337_));
  OAI21X1  g09081(.A0(new_n601_), .A1(new_n7748_), .B0(new_n9337_), .Y(new_n9338_));
  AOI21X1  g09082(.A0(new_n7747_), .A1(new_n518_), .B0(new_n9338_), .Y(new_n9339_));
  XOR2X1   g09083(.A(new_n9339_), .B(\a[11] ), .Y(new_n9340_));
  XOR2X1   g09084(.A(new_n9340_), .B(new_n9336_), .Y(new_n9341_));
  INVX1    g09085(.A(new_n9304_), .Y(new_n9342_));
  AOI21X1  g09086(.A0(new_n9310_), .A1(new_n9309_), .B0(new_n9308_), .Y(new_n9343_));
  AOI21X1  g09087(.A0(new_n9312_), .A1(new_n9342_), .B0(new_n9343_), .Y(new_n9344_));
  AOI22X1  g09088(.A0(new_n818_), .A1(\b[60] ), .B0(new_n817_), .B1(\b[59] ), .Y(new_n9345_));
  OAI21X1  g09089(.A0(new_n816_), .A1(new_n6930_), .B0(new_n9345_), .Y(new_n9346_));
  AOI21X1  g09090(.A0(new_n6951_), .A1(new_n668_), .B0(new_n9346_), .Y(new_n9347_));
  XOR2X1   g09091(.A(new_n9347_), .B(\a[14] ), .Y(new_n9348_));
  XOR2X1   g09092(.A(new_n9348_), .B(new_n9344_), .Y(new_n9349_));
  AOI22X1  g09093(.A0(new_n1017_), .A1(\b[57] ), .B0(new_n1016_), .B1(\b[56] ), .Y(new_n9350_));
  OAI21X1  g09094(.A0(new_n1015_), .A1(new_n6523_), .B0(new_n9350_), .Y(new_n9351_));
  AOI21X1  g09095(.A0(new_n6522_), .A1(new_n882_), .B0(new_n9351_), .Y(new_n9352_));
  XOR2X1   g09096(.A(new_n9352_), .B(\a[17] ), .Y(new_n9353_));
  INVX1    g09097(.A(new_n9353_), .Y(new_n9354_));
  NOR2X1   g09098(.A(new_n9156_), .B(new_n9153_), .Y(new_n9355_));
  INVX1    g09099(.A(new_n9303_), .Y(new_n9356_));
  AOI21X1  g09100(.A0(new_n9356_), .A1(new_n9157_), .B0(new_n9355_), .Y(new_n9357_));
  XOR2X1   g09101(.A(new_n9357_), .B(new_n9354_), .Y(new_n9358_));
  INVX1    g09102(.A(new_n9293_), .Y(new_n9359_));
  NOR2X1   g09103(.A(new_n9300_), .B(new_n9296_), .Y(new_n9360_));
  INVX1    g09104(.A(new_n9360_), .Y(new_n9361_));
  OAI21X1  g09105(.A0(new_n9302_), .A1(new_n9359_), .B0(new_n9361_), .Y(new_n9362_));
  AOI22X1  g09106(.A0(new_n1263_), .A1(\b[54] ), .B0(new_n1262_), .B1(\b[53] ), .Y(new_n9363_));
  OAI21X1  g09107(.A0(new_n1261_), .A1(new_n5808_), .B0(new_n9363_), .Y(new_n9364_));
  AOI21X1  g09108(.A0(new_n5807_), .A1(new_n1075_), .B0(new_n9364_), .Y(new_n9365_));
  XOR2X1   g09109(.A(new_n9365_), .B(\a[20] ), .Y(new_n9366_));
  XOR2X1   g09110(.A(new_n9366_), .B(new_n9362_), .Y(new_n9367_));
  AOI22X1  g09111(.A0(new_n1814_), .A1(\b[48] ), .B0(new_n1813_), .B1(\b[47] ), .Y(new_n9368_));
  OAI21X1  g09112(.A0(new_n1812_), .A1(new_n4693_), .B0(new_n9368_), .Y(new_n9369_));
  AOI21X1  g09113(.A0(new_n4692_), .A1(new_n1617_), .B0(new_n9369_), .Y(new_n9370_));
  XOR2X1   g09114(.A(new_n9370_), .B(\a[26] ), .Y(new_n9371_));
  NOR2X1   g09115(.A(new_n9172_), .B(new_n9169_), .Y(new_n9372_));
  INVX1    g09116(.A(new_n9290_), .Y(new_n9373_));
  AOI21X1  g09117(.A0(new_n9373_), .A1(new_n9173_), .B0(new_n9372_), .Y(new_n9374_));
  XOR2X1   g09118(.A(new_n9374_), .B(new_n9371_), .Y(new_n9375_));
  INVX1    g09119(.A(new_n9288_), .Y(new_n9376_));
  AND2X1   g09120(.A(new_n9376_), .B(new_n9284_), .Y(new_n9377_));
  XOR2X1   g09121(.A(new_n9376_), .B(new_n9284_), .Y(new_n9378_));
  AOI21X1  g09122(.A0(new_n9378_), .A1(new_n9280_), .B0(new_n9377_), .Y(new_n9379_));
  AOI22X1  g09123(.A0(new_n2163_), .A1(\b[45] ), .B0(new_n2162_), .B1(\b[44] ), .Y(new_n9380_));
  OAI21X1  g09124(.A0(new_n2161_), .A1(new_n4339_), .B0(new_n9380_), .Y(new_n9381_));
  AOI21X1  g09125(.A0(new_n4338_), .A1(new_n1907_), .B0(new_n9381_), .Y(new_n9382_));
  XOR2X1   g09126(.A(new_n9382_), .B(\a[29] ), .Y(new_n9383_));
  XOR2X1   g09127(.A(new_n9383_), .B(new_n9379_), .Y(new_n9384_));
  NOR2X1   g09128(.A(new_n9180_), .B(new_n9177_), .Y(new_n9385_));
  AOI21X1  g09129(.A0(new_n9279_), .A1(new_n9181_), .B0(new_n9385_), .Y(new_n9386_));
  AOI22X1  g09130(.A0(new_n2545_), .A1(\b[42] ), .B0(new_n2544_), .B1(\b[41] ), .Y(new_n9387_));
  OAI21X1  g09131(.A0(new_n2543_), .A1(new_n3720_), .B0(new_n9387_), .Y(new_n9388_));
  AOI21X1  g09132(.A0(new_n3860_), .A1(new_n2260_), .B0(new_n9388_), .Y(new_n9389_));
  XOR2X1   g09133(.A(new_n9389_), .B(\a[32] ), .Y(new_n9390_));
  XOR2X1   g09134(.A(new_n9390_), .B(new_n9386_), .Y(new_n9391_));
  NOR2X1   g09135(.A(new_n9264_), .B(new_n9261_), .Y(new_n9392_));
  INVX1    g09136(.A(new_n9392_), .Y(new_n9393_));
  INVX1    g09137(.A(new_n9265_), .Y(new_n9394_));
  OAI21X1  g09138(.A0(new_n9269_), .A1(new_n9394_), .B0(new_n9393_), .Y(new_n9395_));
  NOR2X1   g09139(.A(new_n9253_), .B(new_n9250_), .Y(new_n9396_));
  INVX1    g09140(.A(new_n9396_), .Y(new_n9397_));
  OAI21X1  g09141(.A0(new_n9259_), .A1(new_n9255_), .B0(new_n9397_), .Y(new_n9398_));
  NOR2X1   g09142(.A(new_n9244_), .B(new_n9241_), .Y(new_n9399_));
  INVX1    g09143(.A(new_n9399_), .Y(new_n9400_));
  INVX1    g09144(.A(new_n9245_), .Y(new_n9401_));
  OAI21X1  g09145(.A0(new_n9249_), .A1(new_n9401_), .B0(new_n9400_), .Y(new_n9402_));
  INVX1    g09146(.A(new_n9402_), .Y(new_n9403_));
  NAND2X1  g09147(.A(new_n9233_), .B(new_n9193_), .Y(new_n9404_));
  OAI21X1  g09148(.A0(new_n9234_), .A1(new_n9189_), .B0(new_n9404_), .Y(new_n9405_));
  AOI22X1  g09149(.A0(new_n4880_), .A1(\b[24] ), .B0(new_n4877_), .B1(\b[23] ), .Y(new_n9406_));
  OAI21X1  g09150(.A0(new_n5291_), .A1(new_n1479_), .B0(new_n9406_), .Y(new_n9407_));
  AOI21X1  g09151(.A0(new_n4875_), .A1(new_n1572_), .B0(new_n9407_), .Y(new_n9408_));
  XOR2X1   g09152(.A(new_n9408_), .B(\a[50] ), .Y(new_n9409_));
  INVX1    g09153(.A(new_n9211_), .Y(new_n9410_));
  NOR2X1   g09154(.A(new_n9216_), .B(new_n9212_), .Y(new_n9411_));
  AOI21X1  g09155(.A0(new_n9410_), .A1(new_n9207_), .B0(new_n9411_), .Y(new_n9412_));
  AOI22X1  g09156(.A0(new_n7192_), .A1(\b[12] ), .B0(new_n7189_), .B1(\b[11] ), .Y(new_n9413_));
  OAI21X1  g09157(.A0(new_n7627_), .A1(new_n587_), .B0(new_n9413_), .Y(new_n9414_));
  AOI21X1  g09158(.A0(new_n7187_), .A1(new_n635_), .B0(new_n9414_), .Y(new_n9415_));
  XOR2X1   g09159(.A(new_n9415_), .B(\a[62] ), .Y(new_n9416_));
  AOI22X1  g09160(.A0(new_n7818_), .A1(\b[8] ), .B0(new_n7817_), .B1(\b[9] ), .Y(new_n9417_));
  XOR2X1   g09161(.A(new_n9201_), .B(new_n400_), .Y(new_n9418_));
  XOR2X1   g09162(.A(new_n9418_), .B(new_n9417_), .Y(new_n9419_));
  XOR2X1   g09163(.A(new_n9419_), .B(new_n9206_), .Y(new_n9420_));
  XOR2X1   g09164(.A(new_n9420_), .B(new_n9416_), .Y(new_n9421_));
  AOI22X1  g09165(.A0(new_n6603_), .A1(\b[15] ), .B0(new_n6600_), .B1(\b[14] ), .Y(new_n9422_));
  OAI21X1  g09166(.A0(new_n6804_), .A1(new_n795_), .B0(new_n9422_), .Y(new_n9423_));
  AOI21X1  g09167(.A0(new_n6598_), .A1(new_n794_), .B0(new_n9423_), .Y(new_n9424_));
  XOR2X1   g09168(.A(new_n9424_), .B(\a[59] ), .Y(new_n9425_));
  XOR2X1   g09169(.A(new_n9425_), .B(new_n9421_), .Y(new_n9426_));
  INVX1    g09170(.A(new_n9426_), .Y(new_n9427_));
  XOR2X1   g09171(.A(new_n9427_), .B(new_n9412_), .Y(new_n9428_));
  AOI22X1  g09172(.A0(new_n6438_), .A1(\b[18] ), .B0(new_n6437_), .B1(\b[17] ), .Y(new_n9429_));
  OAI21X1  g09173(.A0(new_n6436_), .A1(new_n974_), .B0(new_n9429_), .Y(new_n9430_));
  AOI21X1  g09174(.A0(new_n6023_), .A1(new_n1042_), .B0(new_n9430_), .Y(new_n9431_));
  XOR2X1   g09175(.A(new_n9431_), .B(\a[56] ), .Y(new_n9432_));
  XOR2X1   g09176(.A(new_n9432_), .B(new_n9428_), .Y(new_n9433_));
  AND2X1   g09177(.A(new_n9217_), .B(new_n9198_), .Y(new_n9434_));
  INVX1    g09178(.A(new_n9222_), .Y(new_n9435_));
  AOI21X1  g09179(.A0(new_n9435_), .A1(new_n9218_), .B0(new_n9434_), .Y(new_n9436_));
  XOR2X1   g09180(.A(new_n9436_), .B(new_n9433_), .Y(new_n9437_));
  AOI22X1  g09181(.A0(new_n5430_), .A1(\b[21] ), .B0(new_n5427_), .B1(\b[20] ), .Y(new_n9438_));
  OAI21X1  g09182(.A0(new_n5891_), .A1(new_n1300_), .B0(new_n9438_), .Y(new_n9439_));
  AOI21X1  g09183(.A0(new_n5425_), .A1(new_n1299_), .B0(new_n9439_), .Y(new_n9440_));
  XOR2X1   g09184(.A(new_n9440_), .B(\a[53] ), .Y(new_n9441_));
  XOR2X1   g09185(.A(new_n9441_), .B(new_n9437_), .Y(new_n9442_));
  OR2X1    g09186(.A(new_n9227_), .B(new_n9223_), .Y(new_n9443_));
  OR2X1    g09187(.A(new_n9232_), .B(new_n9228_), .Y(new_n9444_));
  AND2X1   g09188(.A(new_n9444_), .B(new_n9443_), .Y(new_n9445_));
  XOR2X1   g09189(.A(new_n9445_), .B(new_n9442_), .Y(new_n9446_));
  XOR2X1   g09190(.A(new_n9446_), .B(new_n9409_), .Y(new_n9447_));
  XOR2X1   g09191(.A(new_n9447_), .B(new_n9405_), .Y(new_n9448_));
  AOI22X1  g09192(.A0(new_n4572_), .A1(\b[27] ), .B0(new_n4571_), .B1(\b[26] ), .Y(new_n9449_));
  OAI21X1  g09193(.A0(new_n4740_), .A1(new_n1880_), .B0(new_n9449_), .Y(new_n9450_));
  AOI21X1  g09194(.A0(new_n4375_), .A1(new_n1879_), .B0(new_n9450_), .Y(new_n9451_));
  XOR2X1   g09195(.A(new_n9451_), .B(\a[47] ), .Y(new_n9452_));
  XOR2X1   g09196(.A(new_n9452_), .B(new_n9448_), .Y(new_n9453_));
  AND2X1   g09197(.A(new_n9235_), .B(new_n9185_), .Y(new_n9454_));
  INVX1    g09198(.A(new_n9240_), .Y(new_n9455_));
  AOI21X1  g09199(.A0(new_n9455_), .A1(new_n9236_), .B0(new_n9454_), .Y(new_n9456_));
  XOR2X1   g09200(.A(new_n9456_), .B(new_n9453_), .Y(new_n9457_));
  AOI22X1  g09201(.A0(new_n4095_), .A1(\b[30] ), .B0(new_n4094_), .B1(\b[29] ), .Y(new_n9458_));
  OAI21X1  g09202(.A0(new_n4233_), .A1(new_n2231_), .B0(new_n9458_), .Y(new_n9459_));
  AOI21X1  g09203(.A0(new_n3901_), .A1(new_n2230_), .B0(new_n9459_), .Y(new_n9460_));
  XOR2X1   g09204(.A(new_n9460_), .B(\a[44] ), .Y(new_n9461_));
  AND2X1   g09205(.A(new_n9461_), .B(new_n9457_), .Y(new_n9462_));
  NOR2X1   g09206(.A(new_n9461_), .B(new_n9457_), .Y(new_n9463_));
  NOR3X1   g09207(.A(new_n9463_), .B(new_n9462_), .C(new_n9403_), .Y(new_n9464_));
  NOR2X1   g09208(.A(new_n9464_), .B(new_n9463_), .Y(new_n9465_));
  INVX1    g09209(.A(new_n9465_), .Y(new_n9466_));
  OAI22X1  g09210(.A0(new_n9466_), .A1(new_n9462_), .B0(new_n9464_), .B1(new_n9403_), .Y(new_n9467_));
  AOI22X1  g09211(.A0(new_n3652_), .A1(\b[33] ), .B0(new_n3651_), .B1(\b[32] ), .Y(new_n9468_));
  OAI21X1  g09212(.A0(new_n3778_), .A1(new_n2615_), .B0(new_n9468_), .Y(new_n9469_));
  AOI21X1  g09213(.A0(new_n3480_), .A1(new_n2614_), .B0(new_n9469_), .Y(new_n9470_));
  XOR2X1   g09214(.A(new_n9470_), .B(\a[41] ), .Y(new_n9471_));
  XOR2X1   g09215(.A(new_n9471_), .B(new_n9467_), .Y(new_n9472_));
  XOR2X1   g09216(.A(new_n9472_), .B(new_n9398_), .Y(new_n9473_));
  AOI22X1  g09217(.A0(new_n3204_), .A1(\b[36] ), .B0(new_n3203_), .B1(\b[35] ), .Y(new_n9474_));
  OAI21X1  g09218(.A0(new_n3321_), .A1(new_n2890_), .B0(new_n9474_), .Y(new_n9475_));
  AOI21X1  g09219(.A0(new_n3080_), .A1(new_n3015_), .B0(new_n9475_), .Y(new_n9476_));
  XOR2X1   g09220(.A(new_n9476_), .B(\a[38] ), .Y(new_n9477_));
  XOR2X1   g09221(.A(new_n9477_), .B(new_n9473_), .Y(new_n9478_));
  XOR2X1   g09222(.A(new_n9478_), .B(new_n9395_), .Y(new_n9479_));
  AOI22X1  g09223(.A0(new_n2813_), .A1(\b[39] ), .B0(new_n2812_), .B1(\b[38] ), .Y(new_n9480_));
  OAI21X1  g09224(.A0(new_n2946_), .A1(new_n3413_), .B0(new_n9480_), .Y(new_n9481_));
  AOI21X1  g09225(.A0(new_n3412_), .A1(new_n2652_), .B0(new_n9481_), .Y(new_n9482_));
  XOR2X1   g09226(.A(new_n9482_), .B(\a[35] ), .Y(new_n9483_));
  XOR2X1   g09227(.A(new_n9483_), .B(new_n9479_), .Y(new_n9484_));
  OR2X1    g09228(.A(new_n9273_), .B(new_n9270_), .Y(new_n9485_));
  OAI21X1  g09229(.A0(new_n9278_), .A1(new_n9274_), .B0(new_n9485_), .Y(new_n9486_));
  XOR2X1   g09230(.A(new_n9486_), .B(new_n9484_), .Y(new_n9487_));
  XOR2X1   g09231(.A(new_n9487_), .B(new_n9391_), .Y(new_n9488_));
  XOR2X1   g09232(.A(new_n9488_), .B(new_n9384_), .Y(new_n9489_));
  XOR2X1   g09233(.A(new_n9489_), .B(new_n9375_), .Y(new_n9490_));
  AOI22X1  g09234(.A0(new_n1526_), .A1(\b[51] ), .B0(new_n1525_), .B1(\b[50] ), .Y(new_n9491_));
  OAI21X1  g09235(.A0(new_n1524_), .A1(new_n5237_), .B0(new_n9491_), .Y(new_n9492_));
  AOI21X1  g09236(.A0(new_n5236_), .A1(new_n1347_), .B0(new_n9492_), .Y(new_n9493_));
  XOR2X1   g09237(.A(new_n9493_), .B(\a[23] ), .Y(new_n9494_));
  NOR2X1   g09238(.A(new_n9164_), .B(new_n9161_), .Y(new_n9495_));
  AOI21X1  g09239(.A0(new_n9292_), .A1(new_n9165_), .B0(new_n9495_), .Y(new_n9496_));
  XOR2X1   g09240(.A(new_n9496_), .B(new_n9494_), .Y(new_n9497_));
  XOR2X1   g09241(.A(new_n9497_), .B(new_n9490_), .Y(new_n9498_));
  INVX1    g09242(.A(new_n9498_), .Y(new_n9499_));
  XOR2X1   g09243(.A(new_n9499_), .B(new_n9367_), .Y(new_n9500_));
  XOR2X1   g09244(.A(new_n9500_), .B(new_n9358_), .Y(new_n9501_));
  XOR2X1   g09245(.A(new_n9501_), .B(new_n9349_), .Y(new_n9502_));
  INVX1    g09246(.A(new_n9502_), .Y(new_n9503_));
  XOR2X1   g09247(.A(new_n9503_), .B(new_n9341_), .Y(new_n9504_));
  XOR2X1   g09248(.A(new_n9504_), .B(new_n9335_), .Y(new_n9505_));
  INVX1    g09249(.A(new_n9505_), .Y(new_n9506_));
  XOR2X1   g09250(.A(new_n9506_), .B(new_n9333_), .Y(\f[72] ));
  NOR2X1   g09251(.A(new_n9504_), .B(new_n9335_), .Y(new_n9508_));
  AOI21X1  g09252(.A0(new_n9332_), .A1(new_n9331_), .B0(new_n9506_), .Y(new_n9509_));
  OR2X1    g09253(.A(new_n9509_), .B(new_n9508_), .Y(new_n9510_));
  NOR2X1   g09254(.A(new_n9340_), .B(new_n9336_), .Y(new_n9511_));
  AOI21X1  g09255(.A0(new_n9502_), .A1(new_n9341_), .B0(new_n9511_), .Y(new_n9512_));
  INVX1    g09256(.A(new_n9512_), .Y(new_n9513_));
  OAI22X1  g09257(.A0(new_n601_), .A1(new_n7745_), .B0(new_n660_), .B1(new_n7772_), .Y(new_n9514_));
  AOI21X1  g09258(.A0(new_n7775_), .A1(new_n518_), .B0(new_n9514_), .Y(new_n9515_));
  XOR2X1   g09259(.A(new_n9515_), .B(\a[11] ), .Y(new_n9516_));
  NOR2X1   g09260(.A(new_n9348_), .B(new_n9344_), .Y(new_n9517_));
  AOI21X1  g09261(.A0(new_n9501_), .A1(new_n9349_), .B0(new_n9517_), .Y(new_n9518_));
  NOR2X1   g09262(.A(new_n9516_), .B(new_n9518_), .Y(new_n9519_));
  OR2X1    g09263(.A(new_n9519_), .B(new_n9516_), .Y(new_n9520_));
  AOI22X1  g09264(.A0(new_n818_), .A1(\b[61] ), .B0(new_n817_), .B1(\b[60] ), .Y(new_n9521_));
  OAI21X1  g09265(.A0(new_n816_), .A1(new_n7339_), .B0(new_n9521_), .Y(new_n9522_));
  AOI21X1  g09266(.A0(new_n7338_), .A1(new_n668_), .B0(new_n9522_), .Y(new_n9523_));
  XOR2X1   g09267(.A(new_n9523_), .B(\a[14] ), .Y(new_n9524_));
  OR2X1    g09268(.A(new_n9357_), .B(new_n9353_), .Y(new_n9525_));
  OR2X1    g09269(.A(new_n9500_), .B(new_n9358_), .Y(new_n9526_));
  AND2X1   g09270(.A(new_n9526_), .B(new_n9525_), .Y(new_n9527_));
  XOR2X1   g09271(.A(new_n9527_), .B(new_n9524_), .Y(new_n9528_));
  AOI22X1  g09272(.A0(new_n1263_), .A1(\b[55] ), .B0(new_n1262_), .B1(\b[54] ), .Y(new_n9529_));
  OAI21X1  g09273(.A0(new_n1261_), .A1(new_n6151_), .B0(new_n9529_), .Y(new_n9530_));
  AOI21X1  g09274(.A0(new_n6150_), .A1(new_n1075_), .B0(new_n9530_), .Y(new_n9531_));
  XOR2X1   g09275(.A(new_n9531_), .B(\a[20] ), .Y(new_n9532_));
  INVX1    g09276(.A(new_n9490_), .Y(new_n9533_));
  NOR2X1   g09277(.A(new_n9496_), .B(new_n9494_), .Y(new_n9534_));
  AOI21X1  g09278(.A0(new_n9497_), .A1(new_n9533_), .B0(new_n9534_), .Y(new_n9535_));
  XOR2X1   g09279(.A(new_n9535_), .B(new_n9532_), .Y(new_n9536_));
  AOI22X1  g09280(.A0(new_n1526_), .A1(\b[52] ), .B0(new_n1525_), .B1(\b[51] ), .Y(new_n9537_));
  OAI21X1  g09281(.A0(new_n1524_), .A1(new_n5234_), .B0(new_n9537_), .Y(new_n9538_));
  AOI21X1  g09282(.A0(new_n5590_), .A1(new_n1347_), .B0(new_n9538_), .Y(new_n9539_));
  XOR2X1   g09283(.A(new_n9539_), .B(\a[23] ), .Y(new_n9540_));
  INVX1    g09284(.A(new_n9540_), .Y(new_n9541_));
  NOR2X1   g09285(.A(new_n9374_), .B(new_n9371_), .Y(new_n9542_));
  INVX1    g09286(.A(new_n9489_), .Y(new_n9543_));
  AOI21X1  g09287(.A0(new_n9543_), .A1(new_n9375_), .B0(new_n9542_), .Y(new_n9544_));
  XOR2X1   g09288(.A(new_n9544_), .B(new_n9541_), .Y(new_n9545_));
  AOI22X1  g09289(.A0(new_n1814_), .A1(\b[49] ), .B0(new_n1813_), .B1(\b[48] ), .Y(new_n9546_));
  OAI21X1  g09290(.A0(new_n1812_), .A1(new_n5039_), .B0(new_n9546_), .Y(new_n9547_));
  AOI21X1  g09291(.A0(new_n5038_), .A1(new_n1617_), .B0(new_n9547_), .Y(new_n9548_));
  XOR2X1   g09292(.A(new_n9548_), .B(\a[26] ), .Y(new_n9549_));
  NOR2X1   g09293(.A(new_n9383_), .B(new_n9379_), .Y(new_n9550_));
  INVX1    g09294(.A(new_n9488_), .Y(new_n9551_));
  AOI21X1  g09295(.A0(new_n9551_), .A1(new_n9384_), .B0(new_n9550_), .Y(new_n9552_));
  XOR2X1   g09296(.A(new_n9552_), .B(new_n9549_), .Y(new_n9553_));
  AOI22X1  g09297(.A0(new_n2545_), .A1(\b[43] ), .B0(new_n2544_), .B1(\b[42] ), .Y(new_n9554_));
  OAI21X1  g09298(.A0(new_n2543_), .A1(new_n4015_), .B0(new_n9554_), .Y(new_n9555_));
  AOI21X1  g09299(.A0(new_n4014_), .A1(new_n2260_), .B0(new_n9555_), .Y(new_n9556_));
  XOR2X1   g09300(.A(new_n9556_), .B(\a[32] ), .Y(new_n9557_));
  XOR2X1   g09301(.A(new_n9482_), .B(new_n2650_), .Y(new_n9558_));
  AND2X1   g09302(.A(new_n9558_), .B(new_n9479_), .Y(new_n9559_));
  INVX1    g09303(.A(new_n9484_), .Y(new_n9560_));
  AOI21X1  g09304(.A0(new_n9486_), .A1(new_n9560_), .B0(new_n9559_), .Y(new_n9561_));
  XOR2X1   g09305(.A(new_n9561_), .B(new_n9557_), .Y(new_n9562_));
  AOI22X1  g09306(.A0(new_n2813_), .A1(\b[40] ), .B0(new_n2812_), .B1(\b[39] ), .Y(new_n9563_));
  OAI21X1  g09307(.A0(new_n2946_), .A1(new_n3575_), .B0(new_n9563_), .Y(new_n9564_));
  AOI21X1  g09308(.A0(new_n3574_), .A1(new_n2652_), .B0(new_n9564_), .Y(new_n9565_));
  XOR2X1   g09309(.A(new_n9565_), .B(\a[35] ), .Y(new_n9566_));
  NOR2X1   g09310(.A(new_n9477_), .B(new_n9473_), .Y(new_n9567_));
  AOI21X1  g09311(.A0(new_n9478_), .A1(new_n9395_), .B0(new_n9567_), .Y(new_n9568_));
  AOI22X1  g09312(.A0(new_n3204_), .A1(\b[37] ), .B0(new_n3203_), .B1(\b[36] ), .Y(new_n9569_));
  OAI21X1  g09313(.A0(new_n3321_), .A1(new_n3156_), .B0(new_n9569_), .Y(new_n9570_));
  AOI21X1  g09314(.A0(new_n3155_), .A1(new_n3080_), .B0(new_n9570_), .Y(new_n9571_));
  XOR2X1   g09315(.A(new_n9571_), .B(\a[38] ), .Y(new_n9572_));
  XOR2X1   g09316(.A(new_n9470_), .B(new_n3478_), .Y(new_n9573_));
  AND2X1   g09317(.A(new_n9573_), .B(new_n9467_), .Y(new_n9574_));
  INVX1    g09318(.A(new_n9398_), .Y(new_n9575_));
  NOR2X1   g09319(.A(new_n9472_), .B(new_n9575_), .Y(new_n9576_));
  NOR2X1   g09320(.A(new_n9576_), .B(new_n9574_), .Y(new_n9577_));
  AOI22X1  g09321(.A0(new_n3652_), .A1(\b[34] ), .B0(new_n3651_), .B1(\b[33] ), .Y(new_n9578_));
  OAI21X1  g09322(.A0(new_n3778_), .A1(new_n2612_), .B0(new_n9578_), .Y(new_n9579_));
  AOI21X1  g09323(.A0(new_n3480_), .A1(new_n2759_), .B0(new_n9579_), .Y(new_n9580_));
  XOR2X1   g09324(.A(new_n9580_), .B(new_n3478_), .Y(new_n9581_));
  AOI22X1  g09325(.A0(new_n7192_), .A1(\b[13] ), .B0(new_n7189_), .B1(\b[12] ), .Y(new_n9582_));
  OAI21X1  g09326(.A0(new_n7627_), .A1(new_n716_), .B0(new_n9582_), .Y(new_n9583_));
  AOI21X1  g09327(.A0(new_n7187_), .A1(new_n715_), .B0(new_n9583_), .Y(new_n9584_));
  XOR2X1   g09328(.A(new_n9584_), .B(new_n7185_), .Y(new_n9585_));
  AOI22X1  g09329(.A0(new_n7818_), .A1(\b[9] ), .B0(new_n7817_), .B1(\b[10] ), .Y(new_n9586_));
  NOR2X1   g09330(.A(new_n9418_), .B(new_n9417_), .Y(new_n9587_));
  AOI21X1  g09331(.A0(new_n9202_), .A1(new_n400_), .B0(new_n9587_), .Y(new_n9588_));
  XOR2X1   g09332(.A(new_n9588_), .B(new_n9586_), .Y(new_n9589_));
  XOR2X1   g09333(.A(new_n9589_), .B(new_n9585_), .Y(new_n9590_));
  INVX1    g09334(.A(new_n9416_), .Y(new_n9591_));
  AND2X1   g09335(.A(new_n9419_), .B(new_n9206_), .Y(new_n9592_));
  AOI21X1  g09336(.A0(new_n9420_), .A1(new_n9591_), .B0(new_n9592_), .Y(new_n9593_));
  XOR2X1   g09337(.A(new_n9593_), .B(new_n9590_), .Y(new_n9594_));
  AOI22X1  g09338(.A0(new_n6603_), .A1(\b[16] ), .B0(new_n6600_), .B1(\b[15] ), .Y(new_n9595_));
  OAI21X1  g09339(.A0(new_n6804_), .A1(new_n792_), .B0(new_n9595_), .Y(new_n9596_));
  AOI21X1  g09340(.A0(new_n6598_), .A1(new_n842_), .B0(new_n9596_), .Y(new_n9597_));
  XOR2X1   g09341(.A(new_n9597_), .B(\a[59] ), .Y(new_n9598_));
  XOR2X1   g09342(.A(new_n9598_), .B(new_n9594_), .Y(new_n9599_));
  INVX1    g09343(.A(new_n9599_), .Y(new_n9600_));
  OR2X1    g09344(.A(new_n9425_), .B(new_n9421_), .Y(new_n9601_));
  OAI21X1  g09345(.A0(new_n9427_), .A1(new_n9412_), .B0(new_n9601_), .Y(new_n9602_));
  XOR2X1   g09346(.A(new_n9602_), .B(new_n9600_), .Y(new_n9603_));
  AOI22X1  g09347(.A0(new_n6438_), .A1(\b[19] ), .B0(new_n6437_), .B1(\b[18] ), .Y(new_n9604_));
  OAI21X1  g09348(.A0(new_n6436_), .A1(new_n1118_), .B0(new_n9604_), .Y(new_n9605_));
  AOI21X1  g09349(.A0(new_n6023_), .A1(new_n1117_), .B0(new_n9605_), .Y(new_n9606_));
  XOR2X1   g09350(.A(new_n9606_), .B(\a[56] ), .Y(new_n9607_));
  XOR2X1   g09351(.A(new_n9607_), .B(new_n9603_), .Y(new_n9608_));
  INVX1    g09352(.A(new_n9432_), .Y(new_n9609_));
  NOR2X1   g09353(.A(new_n9436_), .B(new_n9433_), .Y(new_n9610_));
  AOI21X1  g09354(.A0(new_n9609_), .A1(new_n9428_), .B0(new_n9610_), .Y(new_n9611_));
  XOR2X1   g09355(.A(new_n9611_), .B(new_n9608_), .Y(new_n9612_));
  AOI22X1  g09356(.A0(new_n5430_), .A1(\b[22] ), .B0(new_n5427_), .B1(\b[21] ), .Y(new_n9613_));
  OAI21X1  g09357(.A0(new_n5891_), .A1(new_n1297_), .B0(new_n9613_), .Y(new_n9614_));
  AOI21X1  g09358(.A0(new_n5425_), .A1(new_n1399_), .B0(new_n9614_), .Y(new_n9615_));
  XOR2X1   g09359(.A(new_n9615_), .B(\a[53] ), .Y(new_n9616_));
  XOR2X1   g09360(.A(new_n9616_), .B(new_n9612_), .Y(new_n9617_));
  INVX1    g09361(.A(new_n9441_), .Y(new_n9618_));
  NOR2X1   g09362(.A(new_n9445_), .B(new_n9442_), .Y(new_n9619_));
  AOI21X1  g09363(.A0(new_n9618_), .A1(new_n9437_), .B0(new_n9619_), .Y(new_n9620_));
  XOR2X1   g09364(.A(new_n9620_), .B(new_n9617_), .Y(new_n9621_));
  AOI22X1  g09365(.A0(new_n4880_), .A1(\b[25] ), .B0(new_n4877_), .B1(\b[24] ), .Y(new_n9622_));
  OAI21X1  g09366(.A0(new_n5291_), .A1(new_n1591_), .B0(new_n9622_), .Y(new_n9623_));
  AOI21X1  g09367(.A0(new_n4875_), .A1(new_n1590_), .B0(new_n9623_), .Y(new_n9624_));
  XOR2X1   g09368(.A(new_n9624_), .B(\a[50] ), .Y(new_n9625_));
  XOR2X1   g09369(.A(new_n9625_), .B(new_n9621_), .Y(new_n9626_));
  AND2X1   g09370(.A(new_n9445_), .B(new_n9442_), .Y(new_n9627_));
  NOR3X1   g09371(.A(new_n9627_), .B(new_n9619_), .C(new_n9409_), .Y(new_n9628_));
  INVX1    g09372(.A(new_n9447_), .Y(new_n9629_));
  AOI21X1  g09373(.A0(new_n9629_), .A1(new_n9405_), .B0(new_n9628_), .Y(new_n9630_));
  XOR2X1   g09374(.A(new_n9630_), .B(new_n9626_), .Y(new_n9631_));
  AOI22X1  g09375(.A0(new_n4572_), .A1(\b[28] ), .B0(new_n4571_), .B1(\b[27] ), .Y(new_n9632_));
  OAI21X1  g09376(.A0(new_n4740_), .A1(new_n1877_), .B0(new_n9632_), .Y(new_n9633_));
  AOI21X1  g09377(.A0(new_n4375_), .A1(new_n2004_), .B0(new_n9633_), .Y(new_n9634_));
  XOR2X1   g09378(.A(new_n9634_), .B(\a[47] ), .Y(new_n9635_));
  XOR2X1   g09379(.A(new_n9635_), .B(new_n9631_), .Y(new_n9636_));
  OR2X1    g09380(.A(new_n9452_), .B(new_n9448_), .Y(new_n9637_));
  INVX1    g09381(.A(new_n9453_), .Y(new_n9638_));
  OAI21X1  g09382(.A0(new_n9456_), .A1(new_n9638_), .B0(new_n9637_), .Y(new_n9639_));
  XOR2X1   g09383(.A(new_n9639_), .B(new_n9636_), .Y(new_n9640_));
  AOI22X1  g09384(.A0(new_n4095_), .A1(\b[31] ), .B0(new_n4094_), .B1(\b[30] ), .Y(new_n9641_));
  OAI21X1  g09385(.A0(new_n4233_), .A1(new_n2359_), .B0(new_n9641_), .Y(new_n9642_));
  AOI21X1  g09386(.A0(new_n3901_), .A1(new_n2358_), .B0(new_n9642_), .Y(new_n9643_));
  XOR2X1   g09387(.A(new_n9643_), .B(\a[44] ), .Y(new_n9644_));
  XOR2X1   g09388(.A(new_n9644_), .B(new_n9640_), .Y(new_n9645_));
  XOR2X1   g09389(.A(new_n9645_), .B(new_n9466_), .Y(new_n9646_));
  XOR2X1   g09390(.A(new_n9646_), .B(new_n9581_), .Y(new_n9647_));
  XOR2X1   g09391(.A(new_n9647_), .B(new_n9577_), .Y(new_n9648_));
  XOR2X1   g09392(.A(new_n9648_), .B(new_n9572_), .Y(new_n9649_));
  XOR2X1   g09393(.A(new_n9649_), .B(new_n9568_), .Y(new_n9650_));
  XOR2X1   g09394(.A(new_n9650_), .B(new_n9566_), .Y(new_n9651_));
  INVX1    g09395(.A(new_n9651_), .Y(new_n9652_));
  XOR2X1   g09396(.A(new_n9652_), .B(new_n9562_), .Y(new_n9653_));
  INVX1    g09397(.A(new_n9653_), .Y(new_n9654_));
  NOR2X1   g09398(.A(new_n9390_), .B(new_n9386_), .Y(new_n9655_));
  INVX1    g09399(.A(new_n9655_), .Y(new_n9656_));
  INVX1    g09400(.A(new_n9391_), .Y(new_n9657_));
  OAI21X1  g09401(.A0(new_n9487_), .A1(new_n9657_), .B0(new_n9656_), .Y(new_n9658_));
  OAI22X1  g09402(.A0(new_n1913_), .A1(new_n4693_), .B0(new_n1910_), .B1(new_n4674_), .Y(new_n9659_));
  AOI21X1  g09403(.A0(new_n2045_), .A1(\b[44] ), .B0(new_n9659_), .Y(new_n9660_));
  OAI21X1  g09404(.A0(new_n9008_), .A1(new_n2043_), .B0(new_n9660_), .Y(new_n9661_));
  XOR2X1   g09405(.A(new_n9661_), .B(new_n1911_), .Y(new_n9662_));
  XOR2X1   g09406(.A(new_n9662_), .B(new_n9658_), .Y(new_n9663_));
  XOR2X1   g09407(.A(new_n9663_), .B(new_n9654_), .Y(new_n9664_));
  XOR2X1   g09408(.A(new_n9664_), .B(new_n9553_), .Y(new_n9665_));
  XOR2X1   g09409(.A(new_n9665_), .B(new_n9545_), .Y(new_n9666_));
  XOR2X1   g09410(.A(new_n9666_), .B(new_n9536_), .Y(new_n9667_));
  XOR2X1   g09411(.A(new_n9365_), .B(new_n1072_), .Y(new_n9668_));
  NOR2X1   g09412(.A(new_n9498_), .B(new_n9367_), .Y(new_n9669_));
  AOI21X1  g09413(.A0(new_n9668_), .A1(new_n9362_), .B0(new_n9669_), .Y(new_n9670_));
  OAI22X1  g09414(.A0(new_n1068_), .A1(new_n6930_), .B0(new_n1067_), .B1(new_n6933_), .Y(new_n9671_));
  AOI21X1  g09415(.A0(new_n8600_), .A1(\b[56] ), .B0(new_n9671_), .Y(new_n9672_));
  OAI21X1  g09416(.A0(new_n8540_), .A1(new_n934_), .B0(new_n9672_), .Y(new_n9673_));
  XOR2X1   g09417(.A(new_n9673_), .B(new_n879_), .Y(new_n9674_));
  INVX1    g09418(.A(new_n9674_), .Y(new_n9675_));
  XOR2X1   g09419(.A(new_n9675_), .B(new_n9670_), .Y(new_n9676_));
  XOR2X1   g09420(.A(new_n9676_), .B(new_n9667_), .Y(new_n9677_));
  XOR2X1   g09421(.A(new_n9677_), .B(new_n9528_), .Y(new_n9678_));
  INVX1    g09422(.A(new_n9518_), .Y(new_n9679_));
  XOR2X1   g09423(.A(new_n9516_), .B(new_n9679_), .Y(new_n9680_));
  NOR2X1   g09424(.A(new_n9680_), .B(new_n9678_), .Y(new_n9681_));
  NAND2X1  g09425(.A(new_n9516_), .B(new_n9679_), .Y(new_n9682_));
  AND2X1   g09426(.A(new_n9682_), .B(new_n9678_), .Y(new_n9683_));
  AOI21X1  g09427(.A0(new_n9683_), .A1(new_n9520_), .B0(new_n9681_), .Y(new_n9684_));
  XOR2X1   g09428(.A(new_n9684_), .B(new_n9513_), .Y(new_n9685_));
  XOR2X1   g09429(.A(new_n9685_), .B(new_n9510_), .Y(\f[73] ));
  NAND2X1  g09430(.A(new_n9684_), .B(new_n9513_), .Y(new_n9687_));
  OAI21X1  g09431(.A0(new_n9509_), .A1(new_n9508_), .B0(new_n9685_), .Y(new_n9688_));
  AND2X1   g09432(.A(new_n9688_), .B(new_n9687_), .Y(new_n9689_));
  NOR2X1   g09433(.A(new_n9681_), .B(new_n9519_), .Y(new_n9690_));
  AOI21X1  g09434(.A0(new_n9526_), .A1(new_n9525_), .B0(new_n9524_), .Y(new_n9691_));
  INVX1    g09435(.A(new_n9691_), .Y(new_n9692_));
  INVX1    g09436(.A(new_n9528_), .Y(new_n9693_));
  OAI21X1  g09437(.A0(new_n9677_), .A1(new_n9693_), .B0(new_n9692_), .Y(new_n9694_));
  AOI22X1  g09438(.A0(new_n7774_), .A1(new_n518_), .B0(new_n8541_), .B1(\b[63] ), .Y(new_n9695_));
  XOR2X1   g09439(.A(new_n9695_), .B(\a[11] ), .Y(new_n9696_));
  XOR2X1   g09440(.A(new_n9696_), .B(new_n9694_), .Y(new_n9697_));
  NOR2X1   g09441(.A(new_n9674_), .B(new_n9670_), .Y(new_n9698_));
  XOR2X1   g09442(.A(new_n9674_), .B(new_n9670_), .Y(new_n9699_));
  AOI21X1  g09443(.A0(new_n9699_), .A1(new_n9667_), .B0(new_n9698_), .Y(new_n9700_));
  OAI22X1  g09444(.A0(new_n875_), .A1(new_n7745_), .B0(new_n874_), .B1(new_n7748_), .Y(new_n9701_));
  AOI21X1  g09445(.A0(new_n8975_), .A1(\b[60] ), .B0(new_n9701_), .Y(new_n9702_));
  OAI21X1  g09446(.A0(new_n8753_), .A1(new_n751_), .B0(new_n9702_), .Y(new_n9703_));
  XOR2X1   g09447(.A(new_n9703_), .B(new_n665_), .Y(new_n9704_));
  XOR2X1   g09448(.A(new_n9704_), .B(new_n9700_), .Y(new_n9705_));
  AOI22X1  g09449(.A0(new_n1017_), .A1(\b[59] ), .B0(new_n1016_), .B1(\b[58] ), .Y(new_n9706_));
  OAI21X1  g09450(.A0(new_n1015_), .A1(new_n6933_), .B0(new_n9706_), .Y(new_n9707_));
  AOI21X1  g09451(.A0(new_n6932_), .A1(new_n882_), .B0(new_n9707_), .Y(new_n9708_));
  XOR2X1   g09452(.A(new_n9708_), .B(\a[17] ), .Y(new_n9709_));
  INVX1    g09453(.A(new_n9709_), .Y(new_n9710_));
  NOR2X1   g09454(.A(new_n9535_), .B(new_n9532_), .Y(new_n9711_));
  AOI21X1  g09455(.A0(new_n9666_), .A1(new_n9536_), .B0(new_n9711_), .Y(new_n9712_));
  XOR2X1   g09456(.A(new_n9712_), .B(new_n9710_), .Y(new_n9713_));
  AOI22X1  g09457(.A0(new_n1263_), .A1(\b[56] ), .B0(new_n1262_), .B1(\b[55] ), .Y(new_n9714_));
  OAI21X1  g09458(.A0(new_n1261_), .A1(new_n6148_), .B0(new_n9714_), .Y(new_n9715_));
  AOI21X1  g09459(.A0(new_n6342_), .A1(new_n1075_), .B0(new_n9715_), .Y(new_n9716_));
  XOR2X1   g09460(.A(new_n9716_), .B(\a[20] ), .Y(new_n9717_));
  OR2X1    g09461(.A(new_n9544_), .B(new_n9540_), .Y(new_n9718_));
  OR2X1    g09462(.A(new_n9665_), .B(new_n9545_), .Y(new_n9719_));
  AND2X1   g09463(.A(new_n9719_), .B(new_n9718_), .Y(new_n9720_));
  XOR2X1   g09464(.A(new_n9720_), .B(new_n9717_), .Y(new_n9721_));
  XOR2X1   g09465(.A(new_n9661_), .B(\a[29] ), .Y(new_n9722_));
  NOR2X1   g09466(.A(new_n9663_), .B(new_n9653_), .Y(new_n9723_));
  AOI21X1  g09467(.A0(new_n9722_), .A1(new_n9658_), .B0(new_n9723_), .Y(new_n9724_));
  INVX1    g09468(.A(new_n5204_), .Y(new_n9725_));
  OAI22X1  g09469(.A0(new_n1623_), .A1(new_n5234_), .B0(new_n1620_), .B1(new_n5237_), .Y(new_n9726_));
  AOI21X1  g09470(.A0(new_n1725_), .A1(\b[48] ), .B0(new_n9726_), .Y(new_n9727_));
  OAI21X1  g09471(.A0(new_n9725_), .A1(new_n1723_), .B0(new_n9727_), .Y(new_n9728_));
  XOR2X1   g09472(.A(new_n9728_), .B(new_n1621_), .Y(new_n9729_));
  XOR2X1   g09473(.A(new_n9729_), .B(new_n9724_), .Y(new_n9730_));
  AOI22X1  g09474(.A0(new_n2163_), .A1(\b[47] ), .B0(new_n2162_), .B1(\b[46] ), .Y(new_n9731_));
  OAI21X1  g09475(.A0(new_n2161_), .A1(new_n4674_), .B0(new_n9731_), .Y(new_n9732_));
  AOI21X1  g09476(.A0(new_n4673_), .A1(new_n1907_), .B0(new_n9732_), .Y(new_n9733_));
  XOR2X1   g09477(.A(new_n9733_), .B(\a[29] ), .Y(new_n9734_));
  INVX1    g09478(.A(new_n9734_), .Y(new_n9735_));
  NOR2X1   g09479(.A(new_n9561_), .B(new_n9557_), .Y(new_n9736_));
  AOI21X1  g09480(.A0(new_n9651_), .A1(new_n9562_), .B0(new_n9736_), .Y(new_n9737_));
  XOR2X1   g09481(.A(new_n9737_), .B(new_n9735_), .Y(new_n9738_));
  INVX1    g09482(.A(new_n9568_), .Y(new_n9739_));
  NOR2X1   g09483(.A(new_n9650_), .B(new_n9566_), .Y(new_n9740_));
  AOI21X1  g09484(.A0(new_n9649_), .A1(new_n9739_), .B0(new_n9740_), .Y(new_n9741_));
  OAI22X1  g09485(.A0(new_n2263_), .A1(new_n4336_), .B0(new_n2262_), .B1(new_n4339_), .Y(new_n9742_));
  AOI21X1  g09486(.A0(new_n2402_), .A1(\b[42] ), .B0(new_n9742_), .Y(new_n9743_));
  OAI21X1  g09487(.A0(new_n8736_), .A1(new_n2400_), .B0(new_n9743_), .Y(new_n9744_));
  XOR2X1   g09488(.A(new_n9744_), .B(new_n2258_), .Y(new_n9745_));
  XOR2X1   g09489(.A(new_n9745_), .B(new_n9741_), .Y(new_n9746_));
  AOI22X1  g09490(.A0(new_n2813_), .A1(\b[41] ), .B0(new_n2812_), .B1(\b[40] ), .Y(new_n9747_));
  OAI21X1  g09491(.A0(new_n2946_), .A1(new_n3723_), .B0(new_n9747_), .Y(new_n9748_));
  AOI21X1  g09492(.A0(new_n3722_), .A1(new_n2652_), .B0(new_n9748_), .Y(new_n9749_));
  XOR2X1   g09493(.A(new_n9749_), .B(\a[35] ), .Y(new_n9750_));
  OAI21X1  g09494(.A0(new_n9576_), .A1(new_n9574_), .B0(new_n9647_), .Y(new_n9751_));
  OAI21X1  g09495(.A0(new_n9648_), .A1(new_n9572_), .B0(new_n9751_), .Y(new_n9752_));
  NOR2X1   g09496(.A(new_n9620_), .B(new_n9617_), .Y(new_n9753_));
  INVX1    g09497(.A(new_n9753_), .Y(new_n9754_));
  INVX1    g09498(.A(new_n9621_), .Y(new_n9755_));
  OAI21X1  g09499(.A0(new_n9625_), .A1(new_n9755_), .B0(new_n9754_), .Y(new_n9756_));
  AOI22X1  g09500(.A0(new_n4880_), .A1(\b[26] ), .B0(new_n4877_), .B1(\b[25] ), .Y(new_n9757_));
  OAI21X1  g09501(.A0(new_n5291_), .A1(new_n1588_), .B0(new_n9757_), .Y(new_n9758_));
  AOI21X1  g09502(.A0(new_n4875_), .A1(new_n1783_), .B0(new_n9758_), .Y(new_n9759_));
  XOR2X1   g09503(.A(new_n9759_), .B(new_n4873_), .Y(new_n9760_));
  AND2X1   g09504(.A(new_n9611_), .B(new_n9608_), .Y(new_n9761_));
  OR2X1    g09505(.A(new_n9611_), .B(new_n9608_), .Y(new_n9762_));
  OAI21X1  g09506(.A0(new_n9616_), .A1(new_n9761_), .B0(new_n9762_), .Y(new_n9763_));
  AOI22X1  g09507(.A0(new_n5430_), .A1(\b[23] ), .B0(new_n5427_), .B1(\b[22] ), .Y(new_n9764_));
  OAI21X1  g09508(.A0(new_n5891_), .A1(new_n1482_), .B0(new_n9764_), .Y(new_n9765_));
  AOI21X1  g09509(.A0(new_n5425_), .A1(new_n1481_), .B0(new_n9765_), .Y(new_n9766_));
  XOR2X1   g09510(.A(new_n9766_), .B(\a[53] ), .Y(new_n9767_));
  AND2X1   g09511(.A(new_n9602_), .B(new_n9600_), .Y(new_n9768_));
  INVX1    g09512(.A(new_n9768_), .Y(new_n9769_));
  INVX1    g09513(.A(new_n9603_), .Y(new_n9770_));
  OAI21X1  g09514(.A0(new_n9607_), .A1(new_n9770_), .B0(new_n9769_), .Y(new_n9771_));
  INVX1    g09515(.A(new_n9771_), .Y(new_n9772_));
  INVX1    g09516(.A(new_n9586_), .Y(new_n9773_));
  NOR2X1   g09517(.A(new_n9588_), .B(new_n9773_), .Y(new_n9774_));
  INVX1    g09518(.A(new_n9589_), .Y(new_n9775_));
  AOI21X1  g09519(.A0(new_n9775_), .A1(new_n9585_), .B0(new_n9774_), .Y(new_n9776_));
  AOI22X1  g09520(.A0(new_n7818_), .A1(\b[10] ), .B0(new_n7817_), .B1(\b[11] ), .Y(new_n9777_));
  XOR2X1   g09521(.A(new_n9777_), .B(new_n9586_), .Y(new_n9778_));
  XOR2X1   g09522(.A(new_n9778_), .B(new_n9776_), .Y(new_n9779_));
  AOI22X1  g09523(.A0(new_n7192_), .A1(\b[14] ), .B0(new_n7189_), .B1(\b[13] ), .Y(new_n9780_));
  OAI21X1  g09524(.A0(new_n7627_), .A1(new_n713_), .B0(new_n9780_), .Y(new_n9781_));
  AOI21X1  g09525(.A0(new_n7187_), .A1(new_n734_), .B0(new_n9781_), .Y(new_n9782_));
  XOR2X1   g09526(.A(new_n9782_), .B(\a[62] ), .Y(new_n9783_));
  XOR2X1   g09527(.A(new_n9783_), .B(new_n9779_), .Y(new_n9784_));
  AOI22X1  g09528(.A0(new_n6603_), .A1(\b[17] ), .B0(new_n6600_), .B1(\b[16] ), .Y(new_n9785_));
  OAI21X1  g09529(.A0(new_n6804_), .A1(new_n977_), .B0(new_n9785_), .Y(new_n9786_));
  AOI21X1  g09530(.A0(new_n6598_), .A1(new_n976_), .B0(new_n9786_), .Y(new_n9787_));
  XOR2X1   g09531(.A(new_n9787_), .B(\a[59] ), .Y(new_n9788_));
  XOR2X1   g09532(.A(new_n9788_), .B(new_n9784_), .Y(new_n9789_));
  NOR2X1   g09533(.A(new_n9593_), .B(new_n9590_), .Y(new_n9790_));
  INVX1    g09534(.A(new_n9598_), .Y(new_n9791_));
  AOI21X1  g09535(.A0(new_n9791_), .A1(new_n9594_), .B0(new_n9790_), .Y(new_n9792_));
  XOR2X1   g09536(.A(new_n9792_), .B(new_n9789_), .Y(new_n9793_));
  AOI22X1  g09537(.A0(new_n6438_), .A1(\b[20] ), .B0(new_n6437_), .B1(\b[19] ), .Y(new_n9794_));
  OAI21X1  g09538(.A0(new_n6436_), .A1(new_n1115_), .B0(new_n9794_), .Y(new_n9795_));
  AOI21X1  g09539(.A0(new_n6023_), .A1(new_n1217_), .B0(new_n9795_), .Y(new_n9796_));
  XOR2X1   g09540(.A(new_n9796_), .B(\a[56] ), .Y(new_n9797_));
  XOR2X1   g09541(.A(new_n9797_), .B(new_n9793_), .Y(new_n9798_));
  XOR2X1   g09542(.A(new_n9798_), .B(new_n9772_), .Y(new_n9799_));
  XOR2X1   g09543(.A(new_n9799_), .B(new_n9767_), .Y(new_n9800_));
  XOR2X1   g09544(.A(new_n9800_), .B(new_n9763_), .Y(new_n9801_));
  XOR2X1   g09545(.A(new_n9801_), .B(new_n9760_), .Y(new_n9802_));
  XOR2X1   g09546(.A(new_n9802_), .B(new_n9756_), .Y(new_n9803_));
  AOI22X1  g09547(.A0(new_n4572_), .A1(\b[29] ), .B0(new_n4571_), .B1(\b[28] ), .Y(new_n9804_));
  OAI21X1  g09548(.A0(new_n4740_), .A1(new_n2126_), .B0(new_n9804_), .Y(new_n9805_));
  AOI21X1  g09549(.A0(new_n4375_), .A1(new_n2125_), .B0(new_n9805_), .Y(new_n9806_));
  XOR2X1   g09550(.A(new_n9806_), .B(\a[47] ), .Y(new_n9807_));
  XOR2X1   g09551(.A(new_n9807_), .B(new_n9803_), .Y(new_n9808_));
  NOR2X1   g09552(.A(new_n9630_), .B(new_n9626_), .Y(new_n9809_));
  INVX1    g09553(.A(new_n9635_), .Y(new_n9810_));
  AOI21X1  g09554(.A0(new_n9810_), .A1(new_n9631_), .B0(new_n9809_), .Y(new_n9811_));
  XOR2X1   g09555(.A(new_n9811_), .B(new_n9808_), .Y(new_n9812_));
  INVX1    g09556(.A(new_n9812_), .Y(new_n9813_));
  AOI22X1  g09557(.A0(new_n4095_), .A1(\b[32] ), .B0(new_n4094_), .B1(\b[31] ), .Y(new_n9814_));
  OAI21X1  g09558(.A0(new_n4233_), .A1(new_n2356_), .B0(new_n9814_), .Y(new_n9815_));
  AOI21X1  g09559(.A0(new_n3901_), .A1(new_n2495_), .B0(new_n9815_), .Y(new_n9816_));
  XOR2X1   g09560(.A(new_n9816_), .B(\a[44] ), .Y(new_n9817_));
  XOR2X1   g09561(.A(new_n9817_), .B(new_n9813_), .Y(new_n9818_));
  INVX1    g09562(.A(new_n9818_), .Y(new_n9819_));
  INVX1    g09563(.A(new_n9636_), .Y(new_n9820_));
  NOR2X1   g09564(.A(new_n9644_), .B(new_n9640_), .Y(new_n9821_));
  AOI21X1  g09565(.A0(new_n9639_), .A1(new_n9820_), .B0(new_n9821_), .Y(new_n9822_));
  XOR2X1   g09566(.A(new_n9822_), .B(new_n9819_), .Y(new_n9823_));
  AOI22X1  g09567(.A0(new_n3652_), .A1(\b[35] ), .B0(new_n3651_), .B1(\b[34] ), .Y(new_n9824_));
  OAI21X1  g09568(.A0(new_n3778_), .A1(new_n2893_), .B0(new_n9824_), .Y(new_n9825_));
  AOI21X1  g09569(.A0(new_n3480_), .A1(new_n2892_), .B0(new_n9825_), .Y(new_n9826_));
  XOR2X1   g09570(.A(new_n9826_), .B(\a[41] ), .Y(new_n9827_));
  XOR2X1   g09571(.A(new_n9827_), .B(new_n9823_), .Y(new_n9828_));
  INVX1    g09572(.A(new_n9828_), .Y(new_n9829_));
  AND2X1   g09573(.A(new_n9645_), .B(new_n9466_), .Y(new_n9830_));
  AOI21X1  g09574(.A0(new_n9646_), .A1(new_n9581_), .B0(new_n9830_), .Y(new_n9831_));
  XOR2X1   g09575(.A(new_n9831_), .B(new_n9829_), .Y(new_n9832_));
  AOI22X1  g09576(.A0(new_n3204_), .A1(\b[38] ), .B0(new_n3203_), .B1(\b[37] ), .Y(new_n9833_));
  OAI21X1  g09577(.A0(new_n3321_), .A1(new_n3276_), .B0(new_n9833_), .Y(new_n9834_));
  AOI21X1  g09578(.A0(new_n3275_), .A1(new_n3080_), .B0(new_n9834_), .Y(new_n9835_));
  XOR2X1   g09579(.A(new_n9835_), .B(\a[38] ), .Y(new_n9836_));
  XOR2X1   g09580(.A(new_n9836_), .B(new_n9832_), .Y(new_n9837_));
  XOR2X1   g09581(.A(new_n9837_), .B(new_n9752_), .Y(new_n9838_));
  XOR2X1   g09582(.A(new_n9838_), .B(new_n9750_), .Y(new_n9839_));
  XOR2X1   g09583(.A(new_n9839_), .B(new_n9746_), .Y(new_n9840_));
  XOR2X1   g09584(.A(new_n9840_), .B(new_n9738_), .Y(new_n9841_));
  XOR2X1   g09585(.A(new_n9841_), .B(new_n9730_), .Y(new_n9842_));
  NOR2X1   g09586(.A(new_n9552_), .B(new_n9549_), .Y(new_n9843_));
  INVX1    g09587(.A(new_n9843_), .Y(new_n9844_));
  INVX1    g09588(.A(new_n9553_), .Y(new_n9845_));
  OAI21X1  g09589(.A0(new_n9664_), .A1(new_n9845_), .B0(new_n9844_), .Y(new_n9846_));
  OAI22X1  g09590(.A0(new_n1353_), .A1(new_n6151_), .B0(new_n1350_), .B1(new_n5808_), .Y(new_n9847_));
  AOI21X1  g09591(.A0(new_n1430_), .A1(\b[51] ), .B0(new_n9847_), .Y(new_n9848_));
  OAI21X1  g09592(.A0(new_n8599_), .A1(new_n1428_), .B0(new_n9848_), .Y(new_n9849_));
  XOR2X1   g09593(.A(new_n9849_), .B(new_n1351_), .Y(new_n9850_));
  XOR2X1   g09594(.A(new_n9850_), .B(new_n9846_), .Y(new_n9851_));
  XOR2X1   g09595(.A(new_n9851_), .B(new_n9842_), .Y(new_n9852_));
  XOR2X1   g09596(.A(new_n9852_), .B(new_n9721_), .Y(new_n9853_));
  XOR2X1   g09597(.A(new_n9853_), .B(new_n9713_), .Y(new_n9854_));
  XOR2X1   g09598(.A(new_n9854_), .B(new_n9705_), .Y(new_n9855_));
  XOR2X1   g09599(.A(new_n9855_), .B(new_n9697_), .Y(new_n9856_));
  INVX1    g09600(.A(new_n9856_), .Y(new_n9857_));
  XOR2X1   g09601(.A(new_n9857_), .B(new_n9690_), .Y(new_n9858_));
  XOR2X1   g09602(.A(new_n9858_), .B(new_n9689_), .Y(\f[74] ));
  NOR2X1   g09603(.A(new_n9856_), .B(new_n9690_), .Y(new_n9860_));
  AOI21X1  g09604(.A0(new_n9688_), .A1(new_n9687_), .B0(new_n9858_), .Y(new_n9861_));
  OR2X1    g09605(.A(new_n9861_), .B(new_n9860_), .Y(new_n9862_));
  XOR2X1   g09606(.A(new_n9695_), .B(new_n515_), .Y(new_n9863_));
  AND2X1   g09607(.A(new_n9863_), .B(new_n9694_), .Y(new_n9864_));
  INVX1    g09608(.A(new_n9697_), .Y(new_n9865_));
  AOI21X1  g09609(.A0(new_n9855_), .A1(new_n9865_), .B0(new_n9864_), .Y(new_n9866_));
  NOR2X1   g09610(.A(new_n9704_), .B(new_n9700_), .Y(new_n9867_));
  AOI21X1  g09611(.A0(new_n9854_), .A1(new_n9705_), .B0(new_n9867_), .Y(new_n9868_));
  AOI22X1  g09612(.A0(new_n818_), .A1(\b[63] ), .B0(new_n817_), .B1(\b[62] ), .Y(new_n9869_));
  OAI21X1  g09613(.A0(new_n816_), .A1(new_n7748_), .B0(new_n9869_), .Y(new_n9870_));
  AOI21X1  g09614(.A0(new_n7747_), .A1(new_n668_), .B0(new_n9870_), .Y(new_n9871_));
  XOR2X1   g09615(.A(new_n9871_), .B(\a[14] ), .Y(new_n9872_));
  XOR2X1   g09616(.A(new_n9872_), .B(new_n9868_), .Y(new_n9873_));
  NOR2X1   g09617(.A(new_n9712_), .B(new_n9709_), .Y(new_n9874_));
  NOR2X1   g09618(.A(new_n9853_), .B(new_n9713_), .Y(new_n9875_));
  NOR2X1   g09619(.A(new_n9875_), .B(new_n9874_), .Y(new_n9876_));
  AOI22X1  g09620(.A0(new_n1017_), .A1(\b[60] ), .B0(new_n1016_), .B1(\b[59] ), .Y(new_n9877_));
  OAI21X1  g09621(.A0(new_n1015_), .A1(new_n6930_), .B0(new_n9877_), .Y(new_n9878_));
  AOI21X1  g09622(.A0(new_n6951_), .A1(new_n882_), .B0(new_n9878_), .Y(new_n9879_));
  XOR2X1   g09623(.A(new_n9879_), .B(\a[17] ), .Y(new_n9880_));
  INVX1    g09624(.A(new_n9880_), .Y(new_n9881_));
  XOR2X1   g09625(.A(new_n9881_), .B(new_n9876_), .Y(new_n9882_));
  AOI22X1  g09626(.A0(new_n1263_), .A1(\b[57] ), .B0(new_n1262_), .B1(\b[56] ), .Y(new_n9883_));
  OAI21X1  g09627(.A0(new_n1261_), .A1(new_n6523_), .B0(new_n9883_), .Y(new_n9884_));
  AOI21X1  g09628(.A0(new_n6522_), .A1(new_n1075_), .B0(new_n9884_), .Y(new_n9885_));
  XOR2X1   g09629(.A(new_n9885_), .B(\a[20] ), .Y(new_n9886_));
  INVX1    g09630(.A(new_n9886_), .Y(new_n9887_));
  AOI21X1  g09631(.A0(new_n9719_), .A1(new_n9718_), .B0(new_n9717_), .Y(new_n9888_));
  INVX1    g09632(.A(new_n9852_), .Y(new_n9889_));
  AOI21X1  g09633(.A0(new_n9889_), .A1(new_n9721_), .B0(new_n9888_), .Y(new_n9890_));
  XOR2X1   g09634(.A(new_n9890_), .B(new_n9887_), .Y(new_n9891_));
  XOR2X1   g09635(.A(new_n9849_), .B(\a[23] ), .Y(new_n9892_));
  AND2X1   g09636(.A(new_n9892_), .B(new_n9846_), .Y(new_n9893_));
  XOR2X1   g09637(.A(new_n9892_), .B(new_n9846_), .Y(new_n9894_));
  AOI21X1  g09638(.A0(new_n9894_), .A1(new_n9842_), .B0(new_n9893_), .Y(new_n9895_));
  AOI22X1  g09639(.A0(new_n1526_), .A1(\b[54] ), .B0(new_n1525_), .B1(\b[53] ), .Y(new_n9896_));
  OAI21X1  g09640(.A0(new_n1524_), .A1(new_n5808_), .B0(new_n9896_), .Y(new_n9897_));
  AOI21X1  g09641(.A0(new_n5807_), .A1(new_n1347_), .B0(new_n9897_), .Y(new_n9898_));
  XOR2X1   g09642(.A(new_n9898_), .B(\a[23] ), .Y(new_n9899_));
  XOR2X1   g09643(.A(new_n9899_), .B(new_n9895_), .Y(new_n9900_));
  INVX1    g09644(.A(new_n9900_), .Y(new_n9901_));
  AOI22X1  g09645(.A0(new_n1814_), .A1(\b[51] ), .B0(new_n1813_), .B1(\b[50] ), .Y(new_n9902_));
  OAI21X1  g09646(.A0(new_n1812_), .A1(new_n5237_), .B0(new_n9902_), .Y(new_n9903_));
  AOI21X1  g09647(.A0(new_n5236_), .A1(new_n1617_), .B0(new_n9903_), .Y(new_n9904_));
  XOR2X1   g09648(.A(new_n9904_), .B(\a[26] ), .Y(new_n9905_));
  INVX1    g09649(.A(new_n9905_), .Y(new_n9906_));
  NOR2X1   g09650(.A(new_n9729_), .B(new_n9724_), .Y(new_n9907_));
  AOI21X1  g09651(.A0(new_n9841_), .A1(new_n9730_), .B0(new_n9907_), .Y(new_n9908_));
  XOR2X1   g09652(.A(new_n9908_), .B(new_n9906_), .Y(new_n9909_));
  NOR2X1   g09653(.A(new_n9737_), .B(new_n9734_), .Y(new_n9910_));
  NOR2X1   g09654(.A(new_n9840_), .B(new_n9738_), .Y(new_n9911_));
  OR2X1    g09655(.A(new_n9911_), .B(new_n9910_), .Y(new_n9912_));
  AOI22X1  g09656(.A0(new_n2163_), .A1(\b[48] ), .B0(new_n2162_), .B1(\b[47] ), .Y(new_n9913_));
  OAI21X1  g09657(.A0(new_n2161_), .A1(new_n4693_), .B0(new_n9913_), .Y(new_n9914_));
  AOI21X1  g09658(.A0(new_n4692_), .A1(new_n1907_), .B0(new_n9914_), .Y(new_n9915_));
  XOR2X1   g09659(.A(new_n9915_), .B(\a[29] ), .Y(new_n9916_));
  XOR2X1   g09660(.A(new_n9916_), .B(new_n9912_), .Y(new_n9917_));
  INVX1    g09661(.A(new_n9750_), .Y(new_n9918_));
  AND2X1   g09662(.A(new_n9837_), .B(new_n9752_), .Y(new_n9919_));
  AOI21X1  g09663(.A0(new_n9838_), .A1(new_n9918_), .B0(new_n9919_), .Y(new_n9920_));
  NOR2X1   g09664(.A(new_n9831_), .B(new_n9828_), .Y(new_n9921_));
  NOR2X1   g09665(.A(new_n9836_), .B(new_n9832_), .Y(new_n9922_));
  NOR2X1   g09666(.A(new_n9922_), .B(new_n9921_), .Y(new_n9923_));
  NOR2X1   g09667(.A(new_n9822_), .B(new_n9819_), .Y(new_n9924_));
  INVX1    g09668(.A(new_n9924_), .Y(new_n9925_));
  INVX1    g09669(.A(new_n9823_), .Y(new_n9926_));
  OAI21X1  g09670(.A0(new_n9827_), .A1(new_n9926_), .B0(new_n9925_), .Y(new_n9927_));
  NOR2X1   g09671(.A(new_n9811_), .B(new_n9808_), .Y(new_n9928_));
  INVX1    g09672(.A(new_n9928_), .Y(new_n9929_));
  OAI21X1  g09673(.A0(new_n9817_), .A1(new_n9813_), .B0(new_n9929_), .Y(new_n9930_));
  AND2X1   g09674(.A(new_n9802_), .B(new_n9756_), .Y(new_n9931_));
  INVX1    g09675(.A(new_n9931_), .Y(new_n9932_));
  INVX1    g09676(.A(new_n9803_), .Y(new_n9933_));
  OAI21X1  g09677(.A0(new_n9807_), .A1(new_n9933_), .B0(new_n9932_), .Y(new_n9934_));
  INVX1    g09678(.A(new_n9934_), .Y(new_n9935_));
  NAND2X1  g09679(.A(new_n9798_), .B(new_n9771_), .Y(new_n9936_));
  OAI21X1  g09680(.A0(new_n9799_), .A1(new_n9767_), .B0(new_n9936_), .Y(new_n9937_));
  AOI22X1  g09681(.A0(new_n5430_), .A1(\b[24] ), .B0(new_n5427_), .B1(\b[23] ), .Y(new_n9938_));
  OAI21X1  g09682(.A0(new_n5891_), .A1(new_n1479_), .B0(new_n9938_), .Y(new_n9939_));
  AOI21X1  g09683(.A0(new_n5425_), .A1(new_n1572_), .B0(new_n9939_), .Y(new_n9940_));
  XOR2X1   g09684(.A(new_n9940_), .B(\a[53] ), .Y(new_n9941_));
  OR2X1    g09685(.A(new_n9777_), .B(new_n9773_), .Y(new_n9942_));
  OAI21X1  g09686(.A0(new_n9778_), .A1(new_n9776_), .B0(new_n9942_), .Y(new_n9943_));
  AOI22X1  g09687(.A0(new_n7192_), .A1(\b[15] ), .B0(new_n7189_), .B1(\b[14] ), .Y(new_n9944_));
  OAI21X1  g09688(.A0(new_n7627_), .A1(new_n795_), .B0(new_n9944_), .Y(new_n9945_));
  AOI21X1  g09689(.A0(new_n7187_), .A1(new_n794_), .B0(new_n9945_), .Y(new_n9946_));
  XOR2X1   g09690(.A(new_n9946_), .B(\a[62] ), .Y(new_n9947_));
  AOI22X1  g09691(.A0(new_n7818_), .A1(\b[11] ), .B0(new_n7817_), .B1(\b[12] ), .Y(new_n9948_));
  XOR2X1   g09692(.A(new_n9586_), .B(new_n515_), .Y(new_n9949_));
  XOR2X1   g09693(.A(new_n9949_), .B(new_n9948_), .Y(new_n9950_));
  XOR2X1   g09694(.A(new_n9950_), .B(new_n9947_), .Y(new_n9951_));
  XOR2X1   g09695(.A(new_n9951_), .B(new_n9943_), .Y(new_n9952_));
  AOI22X1  g09696(.A0(new_n6603_), .A1(\b[18] ), .B0(new_n6600_), .B1(\b[17] ), .Y(new_n9953_));
  OAI21X1  g09697(.A0(new_n6804_), .A1(new_n974_), .B0(new_n9953_), .Y(new_n9954_));
  AOI21X1  g09698(.A0(new_n6598_), .A1(new_n1042_), .B0(new_n9954_), .Y(new_n9955_));
  XOR2X1   g09699(.A(new_n9955_), .B(\a[59] ), .Y(new_n9956_));
  XOR2X1   g09700(.A(new_n9956_), .B(new_n9952_), .Y(new_n9957_));
  INVX1    g09701(.A(new_n9957_), .Y(new_n9958_));
  INVX1    g09702(.A(new_n9783_), .Y(new_n9959_));
  NOR2X1   g09703(.A(new_n9788_), .B(new_n9784_), .Y(new_n9960_));
  AOI21X1  g09704(.A0(new_n9959_), .A1(new_n9779_), .B0(new_n9960_), .Y(new_n9961_));
  XOR2X1   g09705(.A(new_n9961_), .B(new_n9958_), .Y(new_n9962_));
  AOI22X1  g09706(.A0(new_n6438_), .A1(\b[21] ), .B0(new_n6437_), .B1(\b[20] ), .Y(new_n9963_));
  OAI21X1  g09707(.A0(new_n6436_), .A1(new_n1300_), .B0(new_n9963_), .Y(new_n9964_));
  AOI21X1  g09708(.A0(new_n6023_), .A1(new_n1299_), .B0(new_n9964_), .Y(new_n9965_));
  XOR2X1   g09709(.A(new_n9965_), .B(\a[56] ), .Y(new_n9966_));
  XOR2X1   g09710(.A(new_n9966_), .B(new_n9962_), .Y(new_n9967_));
  AND2X1   g09711(.A(new_n9791_), .B(new_n9594_), .Y(new_n9968_));
  OAI21X1  g09712(.A0(new_n9968_), .A1(new_n9790_), .B0(new_n9789_), .Y(new_n9969_));
  OR2X1    g09713(.A(new_n9797_), .B(new_n9793_), .Y(new_n9970_));
  AND2X1   g09714(.A(new_n9970_), .B(new_n9969_), .Y(new_n9971_));
  XOR2X1   g09715(.A(new_n9971_), .B(new_n9967_), .Y(new_n9972_));
  XOR2X1   g09716(.A(new_n9972_), .B(new_n9941_), .Y(new_n9973_));
  XOR2X1   g09717(.A(new_n9973_), .B(new_n9937_), .Y(new_n9974_));
  AOI22X1  g09718(.A0(new_n4880_), .A1(\b[27] ), .B0(new_n4877_), .B1(\b[26] ), .Y(new_n9975_));
  OAI21X1  g09719(.A0(new_n5291_), .A1(new_n1880_), .B0(new_n9975_), .Y(new_n9976_));
  AOI21X1  g09720(.A0(new_n4875_), .A1(new_n1879_), .B0(new_n9976_), .Y(new_n9977_));
  XOR2X1   g09721(.A(new_n9977_), .B(\a[50] ), .Y(new_n9978_));
  XOR2X1   g09722(.A(new_n9978_), .B(new_n9974_), .Y(new_n9979_));
  AND2X1   g09723(.A(new_n9800_), .B(new_n9763_), .Y(new_n9980_));
  AOI21X1  g09724(.A0(new_n9801_), .A1(new_n9760_), .B0(new_n9980_), .Y(new_n9981_));
  XOR2X1   g09725(.A(new_n9981_), .B(new_n9979_), .Y(new_n9982_));
  AOI22X1  g09726(.A0(new_n4572_), .A1(\b[30] ), .B0(new_n4571_), .B1(\b[29] ), .Y(new_n9983_));
  OAI21X1  g09727(.A0(new_n4740_), .A1(new_n2231_), .B0(new_n9983_), .Y(new_n9984_));
  AOI21X1  g09728(.A0(new_n4375_), .A1(new_n2230_), .B0(new_n9984_), .Y(new_n9985_));
  XOR2X1   g09729(.A(new_n9985_), .B(\a[47] ), .Y(new_n9986_));
  AND2X1   g09730(.A(new_n9986_), .B(new_n9982_), .Y(new_n9987_));
  NOR2X1   g09731(.A(new_n9986_), .B(new_n9982_), .Y(new_n9988_));
  NOR3X1   g09732(.A(new_n9988_), .B(new_n9987_), .C(new_n9935_), .Y(new_n9989_));
  NOR2X1   g09733(.A(new_n9989_), .B(new_n9988_), .Y(new_n9990_));
  INVX1    g09734(.A(new_n9990_), .Y(new_n9991_));
  OAI22X1  g09735(.A0(new_n9991_), .A1(new_n9987_), .B0(new_n9989_), .B1(new_n9935_), .Y(new_n9992_));
  AOI22X1  g09736(.A0(new_n4095_), .A1(\b[33] ), .B0(new_n4094_), .B1(\b[32] ), .Y(new_n9993_));
  OAI21X1  g09737(.A0(new_n4233_), .A1(new_n2615_), .B0(new_n9993_), .Y(new_n9994_));
  AOI21X1  g09738(.A0(new_n3901_), .A1(new_n2614_), .B0(new_n9994_), .Y(new_n9995_));
  XOR2X1   g09739(.A(new_n9995_), .B(\a[44] ), .Y(new_n9996_));
  XOR2X1   g09740(.A(new_n9996_), .B(new_n9992_), .Y(new_n9997_));
  XOR2X1   g09741(.A(new_n9997_), .B(new_n9930_), .Y(new_n9998_));
  AOI22X1  g09742(.A0(new_n3652_), .A1(\b[36] ), .B0(new_n3651_), .B1(\b[35] ), .Y(new_n9999_));
  OAI21X1  g09743(.A0(new_n3778_), .A1(new_n2890_), .B0(new_n9999_), .Y(new_n10000_));
  AOI21X1  g09744(.A0(new_n3480_), .A1(new_n3015_), .B0(new_n10000_), .Y(new_n10001_));
  XOR2X1   g09745(.A(new_n10001_), .B(\a[41] ), .Y(new_n10002_));
  XOR2X1   g09746(.A(new_n10002_), .B(new_n9998_), .Y(new_n10003_));
  XOR2X1   g09747(.A(new_n10003_), .B(new_n9927_), .Y(new_n10004_));
  AOI22X1  g09748(.A0(new_n3204_), .A1(\b[39] ), .B0(new_n3203_), .B1(\b[38] ), .Y(new_n10005_));
  OAI21X1  g09749(.A0(new_n3321_), .A1(new_n3413_), .B0(new_n10005_), .Y(new_n10006_));
  AOI21X1  g09750(.A0(new_n3412_), .A1(new_n3080_), .B0(new_n10006_), .Y(new_n10007_));
  XOR2X1   g09751(.A(new_n10007_), .B(\a[38] ), .Y(new_n10008_));
  XOR2X1   g09752(.A(new_n10008_), .B(new_n10004_), .Y(new_n10009_));
  INVX1    g09753(.A(new_n10009_), .Y(new_n10010_));
  XOR2X1   g09754(.A(new_n10010_), .B(new_n9923_), .Y(new_n10011_));
  AOI22X1  g09755(.A0(new_n2813_), .A1(\b[42] ), .B0(new_n2812_), .B1(\b[41] ), .Y(new_n10012_));
  OAI21X1  g09756(.A0(new_n2946_), .A1(new_n3720_), .B0(new_n10012_), .Y(new_n10013_));
  AOI21X1  g09757(.A0(new_n3860_), .A1(new_n2652_), .B0(new_n10013_), .Y(new_n10014_));
  XOR2X1   g09758(.A(new_n10014_), .B(\a[35] ), .Y(new_n10015_));
  XOR2X1   g09759(.A(new_n10015_), .B(new_n10011_), .Y(new_n10016_));
  XOR2X1   g09760(.A(new_n10016_), .B(new_n9920_), .Y(new_n10017_));
  NOR2X1   g09761(.A(new_n9745_), .B(new_n9741_), .Y(new_n10018_));
  INVX1    g09762(.A(new_n10018_), .Y(new_n10019_));
  INVX1    g09763(.A(new_n9746_), .Y(new_n10020_));
  OAI21X1  g09764(.A0(new_n9839_), .A1(new_n10020_), .B0(new_n10019_), .Y(new_n10021_));
  AOI22X1  g09765(.A0(new_n2545_), .A1(\b[45] ), .B0(new_n2544_), .B1(\b[44] ), .Y(new_n10022_));
  OAI21X1  g09766(.A0(new_n2543_), .A1(new_n4339_), .B0(new_n10022_), .Y(new_n10023_));
  AOI21X1  g09767(.A0(new_n4338_), .A1(new_n2260_), .B0(new_n10023_), .Y(new_n10024_));
  XOR2X1   g09768(.A(new_n10024_), .B(\a[32] ), .Y(new_n10025_));
  XOR2X1   g09769(.A(new_n10025_), .B(new_n10021_), .Y(new_n10026_));
  XOR2X1   g09770(.A(new_n10026_), .B(new_n10017_), .Y(new_n10027_));
  XOR2X1   g09771(.A(new_n10027_), .B(new_n9917_), .Y(new_n10028_));
  XOR2X1   g09772(.A(new_n10028_), .B(new_n9909_), .Y(new_n10029_));
  XOR2X1   g09773(.A(new_n10029_), .B(new_n9901_), .Y(new_n10030_));
  XOR2X1   g09774(.A(new_n10030_), .B(new_n9891_), .Y(new_n10031_));
  XOR2X1   g09775(.A(new_n10031_), .B(new_n9882_), .Y(new_n10032_));
  XOR2X1   g09776(.A(new_n10032_), .B(new_n9873_), .Y(new_n10033_));
  XOR2X1   g09777(.A(new_n10033_), .B(new_n9866_), .Y(new_n10034_));
  XOR2X1   g09778(.A(new_n10034_), .B(new_n9862_), .Y(\f[75] ));
  NOR2X1   g09779(.A(new_n10033_), .B(new_n9866_), .Y(new_n10036_));
  INVX1    g09780(.A(new_n10036_), .Y(new_n10037_));
  OAI21X1  g09781(.A0(new_n9861_), .A1(new_n9860_), .B0(new_n10034_), .Y(new_n10038_));
  AND2X1   g09782(.A(new_n10038_), .B(new_n10037_), .Y(new_n10039_));
  NOR2X1   g09783(.A(new_n9872_), .B(new_n9868_), .Y(new_n10040_));
  INVX1    g09784(.A(new_n10032_), .Y(new_n10041_));
  AOI21X1  g09785(.A0(new_n10041_), .A1(new_n9873_), .B0(new_n10040_), .Y(new_n10042_));
  AOI22X1  g09786(.A0(new_n1017_), .A1(\b[61] ), .B0(new_n1016_), .B1(\b[60] ), .Y(new_n10043_));
  OAI21X1  g09787(.A0(new_n1015_), .A1(new_n7339_), .B0(new_n10043_), .Y(new_n10044_));
  AOI21X1  g09788(.A0(new_n7338_), .A1(new_n882_), .B0(new_n10044_), .Y(new_n10045_));
  XOR2X1   g09789(.A(new_n10045_), .B(\a[17] ), .Y(new_n10046_));
  OR2X1    g09790(.A(new_n9890_), .B(new_n9886_), .Y(new_n10047_));
  OR2X1    g09791(.A(new_n10030_), .B(new_n9891_), .Y(new_n10048_));
  AND2X1   g09792(.A(new_n10048_), .B(new_n10047_), .Y(new_n10049_));
  XOR2X1   g09793(.A(new_n10049_), .B(new_n10046_), .Y(new_n10050_));
  AOI22X1  g09794(.A0(new_n1526_), .A1(\b[55] ), .B0(new_n1525_), .B1(\b[54] ), .Y(new_n10051_));
  OAI21X1  g09795(.A0(new_n1524_), .A1(new_n6151_), .B0(new_n10051_), .Y(new_n10052_));
  AOI21X1  g09796(.A0(new_n6150_), .A1(new_n1347_), .B0(new_n10052_), .Y(new_n10053_));
  XOR2X1   g09797(.A(new_n10053_), .B(\a[23] ), .Y(new_n10054_));
  OR2X1    g09798(.A(new_n9908_), .B(new_n9905_), .Y(new_n10055_));
  OR2X1    g09799(.A(new_n10028_), .B(new_n9909_), .Y(new_n10056_));
  AND2X1   g09800(.A(new_n10056_), .B(new_n10055_), .Y(new_n10057_));
  XOR2X1   g09801(.A(new_n10057_), .B(new_n10054_), .Y(new_n10058_));
  AOI22X1  g09802(.A0(new_n2163_), .A1(\b[49] ), .B0(new_n2162_), .B1(\b[48] ), .Y(new_n10059_));
  OAI21X1  g09803(.A0(new_n2161_), .A1(new_n5039_), .B0(new_n10059_), .Y(new_n10060_));
  AOI21X1  g09804(.A0(new_n5038_), .A1(new_n1907_), .B0(new_n10060_), .Y(new_n10061_));
  XOR2X1   g09805(.A(new_n10061_), .B(\a[29] ), .Y(new_n10062_));
  INVX1    g09806(.A(new_n10025_), .Y(new_n10063_));
  NOR2X1   g09807(.A(new_n10026_), .B(new_n10017_), .Y(new_n10064_));
  AOI21X1  g09808(.A0(new_n10063_), .A1(new_n10021_), .B0(new_n10064_), .Y(new_n10065_));
  XOR2X1   g09809(.A(new_n10065_), .B(new_n10062_), .Y(new_n10066_));
  XOR2X1   g09810(.A(new_n10007_), .B(new_n3078_), .Y(new_n10067_));
  NOR2X1   g09811(.A(new_n10009_), .B(new_n9923_), .Y(new_n10068_));
  AOI21X1  g09812(.A0(new_n10067_), .A1(new_n10004_), .B0(new_n10068_), .Y(new_n10069_));
  INVX1    g09813(.A(new_n10069_), .Y(new_n10070_));
  AOI22X1  g09814(.A0(new_n3204_), .A1(\b[40] ), .B0(new_n3203_), .B1(\b[39] ), .Y(new_n10071_));
  OAI21X1  g09815(.A0(new_n3321_), .A1(new_n3575_), .B0(new_n10071_), .Y(new_n10072_));
  AOI21X1  g09816(.A0(new_n3574_), .A1(new_n3080_), .B0(new_n10072_), .Y(new_n10073_));
  XOR2X1   g09817(.A(new_n10073_), .B(\a[38] ), .Y(new_n10074_));
  NOR2X1   g09818(.A(new_n10002_), .B(new_n9998_), .Y(new_n10075_));
  AOI21X1  g09819(.A0(new_n10003_), .A1(new_n9927_), .B0(new_n10075_), .Y(new_n10076_));
  AOI22X1  g09820(.A0(new_n3652_), .A1(\b[37] ), .B0(new_n3651_), .B1(\b[36] ), .Y(new_n10077_));
  OAI21X1  g09821(.A0(new_n3778_), .A1(new_n3156_), .B0(new_n10077_), .Y(new_n10078_));
  AOI21X1  g09822(.A0(new_n3480_), .A1(new_n3155_), .B0(new_n10078_), .Y(new_n10079_));
  XOR2X1   g09823(.A(new_n10079_), .B(\a[41] ), .Y(new_n10080_));
  XOR2X1   g09824(.A(new_n9995_), .B(new_n3899_), .Y(new_n10081_));
  AND2X1   g09825(.A(new_n10081_), .B(new_n9992_), .Y(new_n10082_));
  INVX1    g09826(.A(new_n9930_), .Y(new_n10083_));
  NOR2X1   g09827(.A(new_n9997_), .B(new_n10083_), .Y(new_n10084_));
  NOR2X1   g09828(.A(new_n10084_), .B(new_n10082_), .Y(new_n10085_));
  AOI22X1  g09829(.A0(new_n4095_), .A1(\b[34] ), .B0(new_n4094_), .B1(\b[33] ), .Y(new_n10086_));
  OAI21X1  g09830(.A0(new_n4233_), .A1(new_n2612_), .B0(new_n10086_), .Y(new_n10087_));
  AOI21X1  g09831(.A0(new_n3901_), .A1(new_n2759_), .B0(new_n10087_), .Y(new_n10088_));
  XOR2X1   g09832(.A(new_n10088_), .B(new_n3899_), .Y(new_n10089_));
  AOI22X1  g09833(.A0(new_n4572_), .A1(\b[31] ), .B0(new_n4571_), .B1(\b[30] ), .Y(new_n10090_));
  OAI21X1  g09834(.A0(new_n4740_), .A1(new_n2359_), .B0(new_n10090_), .Y(new_n10091_));
  AOI21X1  g09835(.A0(new_n4375_), .A1(new_n2358_), .B0(new_n10091_), .Y(new_n10092_));
  XOR2X1   g09836(.A(new_n10092_), .B(\a[47] ), .Y(new_n10093_));
  NOR2X1   g09837(.A(new_n9978_), .B(new_n9974_), .Y(new_n10094_));
  INVX1    g09838(.A(new_n10094_), .Y(new_n10095_));
  INVX1    g09839(.A(new_n9979_), .Y(new_n10096_));
  OAI21X1  g09840(.A0(new_n9981_), .A1(new_n10096_), .B0(new_n10095_), .Y(new_n10097_));
  INVX1    g09841(.A(new_n10097_), .Y(new_n10098_));
  AOI22X1  g09842(.A0(new_n7818_), .A1(\b[12] ), .B0(new_n7817_), .B1(\b[13] ), .Y(new_n10099_));
  NOR2X1   g09843(.A(new_n9949_), .B(new_n9948_), .Y(new_n10100_));
  AOI21X1  g09844(.A0(new_n9773_), .A1(new_n515_), .B0(new_n10100_), .Y(new_n10101_));
  XOR2X1   g09845(.A(new_n10101_), .B(new_n10099_), .Y(new_n10102_));
  INVX1    g09846(.A(new_n10102_), .Y(new_n10103_));
  AOI22X1  g09847(.A0(new_n7192_), .A1(\b[16] ), .B0(new_n7189_), .B1(\b[15] ), .Y(new_n10104_));
  OAI21X1  g09848(.A0(new_n7627_), .A1(new_n792_), .B0(new_n10104_), .Y(new_n10105_));
  AOI21X1  g09849(.A0(new_n7187_), .A1(new_n842_), .B0(new_n10105_), .Y(new_n10106_));
  XOR2X1   g09850(.A(new_n10106_), .B(\a[62] ), .Y(new_n10107_));
  XOR2X1   g09851(.A(new_n10107_), .B(new_n10103_), .Y(new_n10108_));
  AND2X1   g09852(.A(new_n9949_), .B(new_n9948_), .Y(new_n10109_));
  NOR3X1   g09853(.A(new_n10109_), .B(new_n10100_), .C(new_n9947_), .Y(new_n10110_));
  INVX1    g09854(.A(new_n9951_), .Y(new_n10111_));
  AOI21X1  g09855(.A0(new_n10111_), .A1(new_n9943_), .B0(new_n10110_), .Y(new_n10112_));
  XOR2X1   g09856(.A(new_n10112_), .B(new_n10108_), .Y(new_n10113_));
  AOI22X1  g09857(.A0(new_n6603_), .A1(\b[19] ), .B0(new_n6600_), .B1(\b[18] ), .Y(new_n10114_));
  OAI21X1  g09858(.A0(new_n6804_), .A1(new_n1118_), .B0(new_n10114_), .Y(new_n10115_));
  AOI21X1  g09859(.A0(new_n6598_), .A1(new_n1117_), .B0(new_n10115_), .Y(new_n10116_));
  XOR2X1   g09860(.A(new_n10116_), .B(\a[59] ), .Y(new_n10117_));
  XOR2X1   g09861(.A(new_n10117_), .B(new_n10113_), .Y(new_n10118_));
  INVX1    g09862(.A(new_n10118_), .Y(new_n10119_));
  OR2X1    g09863(.A(new_n9956_), .B(new_n9952_), .Y(new_n10120_));
  OAI21X1  g09864(.A0(new_n9961_), .A1(new_n9958_), .B0(new_n10120_), .Y(new_n10121_));
  XOR2X1   g09865(.A(new_n10121_), .B(new_n10119_), .Y(new_n10122_));
  AOI22X1  g09866(.A0(new_n6438_), .A1(\b[22] ), .B0(new_n6437_), .B1(\b[21] ), .Y(new_n10123_));
  OAI21X1  g09867(.A0(new_n6436_), .A1(new_n1297_), .B0(new_n10123_), .Y(new_n10124_));
  AOI21X1  g09868(.A0(new_n6023_), .A1(new_n1399_), .B0(new_n10124_), .Y(new_n10125_));
  XOR2X1   g09869(.A(new_n10125_), .B(\a[56] ), .Y(new_n10126_));
  XOR2X1   g09870(.A(new_n10126_), .B(new_n10122_), .Y(new_n10127_));
  INVX1    g09871(.A(new_n9966_), .Y(new_n10128_));
  NOR2X1   g09872(.A(new_n9971_), .B(new_n9967_), .Y(new_n10129_));
  AOI21X1  g09873(.A0(new_n10128_), .A1(new_n9962_), .B0(new_n10129_), .Y(new_n10130_));
  XOR2X1   g09874(.A(new_n10130_), .B(new_n10127_), .Y(new_n10131_));
  AOI22X1  g09875(.A0(new_n5430_), .A1(\b[25] ), .B0(new_n5427_), .B1(\b[24] ), .Y(new_n10132_));
  OAI21X1  g09876(.A0(new_n5891_), .A1(new_n1591_), .B0(new_n10132_), .Y(new_n10133_));
  AOI21X1  g09877(.A0(new_n5425_), .A1(new_n1590_), .B0(new_n10133_), .Y(new_n10134_));
  XOR2X1   g09878(.A(new_n10134_), .B(\a[53] ), .Y(new_n10135_));
  XOR2X1   g09879(.A(new_n10135_), .B(new_n10131_), .Y(new_n10136_));
  INVX1    g09880(.A(new_n10136_), .Y(new_n10137_));
  AND2X1   g09881(.A(new_n9971_), .B(new_n9967_), .Y(new_n10138_));
  NOR3X1   g09882(.A(new_n10138_), .B(new_n10129_), .C(new_n9941_), .Y(new_n10139_));
  INVX1    g09883(.A(new_n9973_), .Y(new_n10140_));
  AOI21X1  g09884(.A0(new_n10140_), .A1(new_n9937_), .B0(new_n10139_), .Y(new_n10141_));
  XOR2X1   g09885(.A(new_n10141_), .B(new_n10137_), .Y(new_n10142_));
  AOI22X1  g09886(.A0(new_n4880_), .A1(\b[28] ), .B0(new_n4877_), .B1(\b[27] ), .Y(new_n10143_));
  OAI21X1  g09887(.A0(new_n5291_), .A1(new_n1877_), .B0(new_n10143_), .Y(new_n10144_));
  AOI21X1  g09888(.A0(new_n4875_), .A1(new_n2004_), .B0(new_n10144_), .Y(new_n10145_));
  XOR2X1   g09889(.A(new_n10145_), .B(\a[50] ), .Y(new_n10146_));
  XOR2X1   g09890(.A(new_n10146_), .B(new_n10142_), .Y(new_n10147_));
  XOR2X1   g09891(.A(new_n10147_), .B(new_n10098_), .Y(new_n10148_));
  XOR2X1   g09892(.A(new_n10148_), .B(new_n10093_), .Y(new_n10149_));
  XOR2X1   g09893(.A(new_n10149_), .B(new_n9991_), .Y(new_n10150_));
  XOR2X1   g09894(.A(new_n10150_), .B(new_n10089_), .Y(new_n10151_));
  XOR2X1   g09895(.A(new_n10151_), .B(new_n10085_), .Y(new_n10152_));
  XOR2X1   g09896(.A(new_n10152_), .B(new_n10080_), .Y(new_n10153_));
  XOR2X1   g09897(.A(new_n10153_), .B(new_n10076_), .Y(new_n10154_));
  XOR2X1   g09898(.A(new_n10154_), .B(new_n10074_), .Y(new_n10155_));
  XOR2X1   g09899(.A(new_n10155_), .B(new_n10070_), .Y(new_n10156_));
  AOI22X1  g09900(.A0(new_n2813_), .A1(\b[43] ), .B0(new_n2812_), .B1(\b[42] ), .Y(new_n10157_));
  OAI21X1  g09901(.A0(new_n2946_), .A1(new_n4015_), .B0(new_n10157_), .Y(new_n10158_));
  AOI21X1  g09902(.A0(new_n4014_), .A1(new_n2652_), .B0(new_n10158_), .Y(new_n10159_));
  XOR2X1   g09903(.A(new_n10159_), .B(\a[35] ), .Y(new_n10160_));
  XOR2X1   g09904(.A(new_n10160_), .B(new_n10156_), .Y(new_n10161_));
  INVX1    g09905(.A(new_n9920_), .Y(new_n10162_));
  NOR2X1   g09906(.A(new_n10015_), .B(new_n10011_), .Y(new_n10163_));
  AOI21X1  g09907(.A0(new_n10016_), .A1(new_n10162_), .B0(new_n10163_), .Y(new_n10164_));
  OAI22X1  g09908(.A0(new_n2263_), .A1(new_n4693_), .B0(new_n2262_), .B1(new_n4674_), .Y(new_n10165_));
  AOI21X1  g09909(.A0(new_n2402_), .A1(\b[44] ), .B0(new_n10165_), .Y(new_n10166_));
  OAI21X1  g09910(.A0(new_n9008_), .A1(new_n2400_), .B0(new_n10166_), .Y(new_n10167_));
  XOR2X1   g09911(.A(new_n10167_), .B(new_n2258_), .Y(new_n10168_));
  XOR2X1   g09912(.A(new_n10168_), .B(new_n10164_), .Y(new_n10169_));
  XOR2X1   g09913(.A(new_n10169_), .B(new_n10161_), .Y(new_n10170_));
  XOR2X1   g09914(.A(new_n10170_), .B(new_n10066_), .Y(new_n10171_));
  INVX1    g09915(.A(new_n9917_), .Y(new_n10172_));
  INVX1    g09916(.A(new_n9916_), .Y(new_n10173_));
  AND2X1   g09917(.A(new_n10173_), .B(new_n9912_), .Y(new_n10174_));
  AOI21X1  g09918(.A0(new_n10027_), .A1(new_n10172_), .B0(new_n10174_), .Y(new_n10175_));
  NOR3X1   g09919(.A(new_n1724_), .B(new_n1622_), .C(new_n5234_), .Y(new_n10176_));
  OAI22X1  g09920(.A0(new_n1623_), .A1(new_n5808_), .B0(new_n1620_), .B1(new_n5787_), .Y(new_n10177_));
  OR2X1    g09921(.A(new_n10177_), .B(new_n10176_), .Y(new_n10178_));
  AOI21X1  g09922(.A0(new_n5590_), .A1(new_n1617_), .B0(new_n10178_), .Y(new_n10179_));
  XOR2X1   g09923(.A(new_n10179_), .B(\a[26] ), .Y(new_n10180_));
  XOR2X1   g09924(.A(new_n10180_), .B(new_n10175_), .Y(new_n10181_));
  XOR2X1   g09925(.A(new_n10181_), .B(new_n10171_), .Y(new_n10182_));
  XOR2X1   g09926(.A(new_n10182_), .B(new_n10058_), .Y(new_n10183_));
  NOR2X1   g09927(.A(new_n9899_), .B(new_n9895_), .Y(new_n10184_));
  AOI21X1  g09928(.A0(new_n10029_), .A1(new_n9900_), .B0(new_n10184_), .Y(new_n10185_));
  OAI22X1  g09929(.A0(new_n1080_), .A1(new_n6930_), .B0(new_n1078_), .B1(new_n6933_), .Y(new_n10186_));
  AOI21X1  g09930(.A0(new_n1167_), .A1(\b[56] ), .B0(new_n10186_), .Y(new_n10187_));
  OAI21X1  g09931(.A0(new_n8540_), .A1(new_n1165_), .B0(new_n10187_), .Y(new_n10188_));
  XOR2X1   g09932(.A(new_n10188_), .B(new_n1072_), .Y(new_n10189_));
  INVX1    g09933(.A(new_n10189_), .Y(new_n10190_));
  XOR2X1   g09934(.A(new_n10190_), .B(new_n10185_), .Y(new_n10191_));
  XOR2X1   g09935(.A(new_n10191_), .B(new_n10183_), .Y(new_n10192_));
  INVX1    g09936(.A(new_n10192_), .Y(new_n10193_));
  XOR2X1   g09937(.A(new_n10193_), .B(new_n10050_), .Y(new_n10194_));
  INVX1    g09938(.A(new_n9882_), .Y(new_n10195_));
  NOR2X1   g09939(.A(new_n9880_), .B(new_n9876_), .Y(new_n10196_));
  AOI21X1  g09940(.A0(new_n10031_), .A1(new_n10195_), .B0(new_n10196_), .Y(new_n10197_));
  INVX1    g09941(.A(new_n10197_), .Y(new_n10198_));
  OAI22X1  g09942(.A0(new_n816_), .A1(new_n7745_), .B0(new_n874_), .B1(new_n7772_), .Y(new_n10199_));
  AOI21X1  g09943(.A0(new_n7775_), .A1(new_n668_), .B0(new_n10199_), .Y(new_n10200_));
  XOR2X1   g09944(.A(new_n10200_), .B(\a[14] ), .Y(new_n10201_));
  XOR2X1   g09945(.A(new_n10201_), .B(new_n10198_), .Y(new_n10202_));
  NOR2X1   g09946(.A(new_n10202_), .B(new_n10194_), .Y(new_n10203_));
  OR2X1    g09947(.A(new_n10201_), .B(new_n10198_), .Y(new_n10204_));
  INVX1    g09948(.A(new_n10194_), .Y(new_n10205_));
  AOI21X1  g09949(.A0(new_n10201_), .A1(new_n10198_), .B0(new_n10205_), .Y(new_n10206_));
  AND2X1   g09950(.A(new_n10206_), .B(new_n10204_), .Y(new_n10207_));
  NOR2X1   g09951(.A(new_n10207_), .B(new_n10203_), .Y(new_n10208_));
  XOR2X1   g09952(.A(new_n10208_), .B(new_n10042_), .Y(new_n10209_));
  XOR2X1   g09953(.A(new_n10209_), .B(new_n10039_), .Y(\f[76] ));
  NOR3X1   g09954(.A(new_n10207_), .B(new_n10203_), .C(new_n10042_), .Y(new_n10211_));
  AOI21X1  g09955(.A0(new_n10038_), .A1(new_n10037_), .B0(new_n10209_), .Y(new_n10212_));
  OR2X1    g09956(.A(new_n10212_), .B(new_n10211_), .Y(new_n10213_));
  OR2X1    g09957(.A(new_n10201_), .B(new_n10197_), .Y(new_n10214_));
  OAI21X1  g09958(.A0(new_n10202_), .A1(new_n10194_), .B0(new_n10214_), .Y(new_n10215_));
  AOI21X1  g09959(.A0(new_n10048_), .A1(new_n10047_), .B0(new_n10046_), .Y(new_n10216_));
  AOI21X1  g09960(.A0(new_n10192_), .A1(new_n10050_), .B0(new_n10216_), .Y(new_n10217_));
  AOI22X1  g09961(.A0(new_n7774_), .A1(new_n668_), .B0(new_n8975_), .B1(\b[63] ), .Y(new_n10218_));
  XOR2X1   g09962(.A(new_n10218_), .B(\a[14] ), .Y(new_n10219_));
  XOR2X1   g09963(.A(new_n10219_), .B(new_n10217_), .Y(new_n10220_));
  OAI22X1  g09964(.A0(new_n1068_), .A1(new_n7745_), .B0(new_n1067_), .B1(new_n7748_), .Y(new_n10221_));
  AOI21X1  g09965(.A0(new_n8600_), .A1(\b[60] ), .B0(new_n10221_), .Y(new_n10222_));
  OAI21X1  g09966(.A0(new_n8753_), .A1(new_n934_), .B0(new_n10222_), .Y(new_n10223_));
  XOR2X1   g09967(.A(new_n10223_), .B(new_n879_), .Y(new_n10224_));
  NOR2X1   g09968(.A(new_n10189_), .B(new_n10185_), .Y(new_n10225_));
  NOR2X1   g09969(.A(new_n10191_), .B(new_n10183_), .Y(new_n10226_));
  NOR2X1   g09970(.A(new_n10226_), .B(new_n10225_), .Y(new_n10227_));
  NOR2X1   g09971(.A(new_n10224_), .B(new_n10227_), .Y(new_n10228_));
  OR2X1    g09972(.A(new_n10228_), .B(new_n10224_), .Y(new_n10229_));
  AOI22X1  g09973(.A0(new_n1263_), .A1(\b[59] ), .B0(new_n1262_), .B1(\b[58] ), .Y(new_n10230_));
  OAI21X1  g09974(.A0(new_n1261_), .A1(new_n6933_), .B0(new_n10230_), .Y(new_n10231_));
  AOI21X1  g09975(.A0(new_n6932_), .A1(new_n1075_), .B0(new_n10231_), .Y(new_n10232_));
  XOR2X1   g09976(.A(new_n10232_), .B(\a[20] ), .Y(new_n10233_));
  AOI21X1  g09977(.A0(new_n10056_), .A1(new_n10055_), .B0(new_n10054_), .Y(new_n10234_));
  INVX1    g09978(.A(new_n10182_), .Y(new_n10235_));
  AOI21X1  g09979(.A0(new_n10235_), .A1(new_n10058_), .B0(new_n10234_), .Y(new_n10236_));
  XOR2X1   g09980(.A(new_n10236_), .B(new_n10233_), .Y(new_n10237_));
  AOI22X1  g09981(.A0(new_n1526_), .A1(\b[56] ), .B0(new_n1525_), .B1(\b[55] ), .Y(new_n10238_));
  OAI21X1  g09982(.A0(new_n1524_), .A1(new_n6148_), .B0(new_n10238_), .Y(new_n10239_));
  AOI21X1  g09983(.A0(new_n6342_), .A1(new_n1347_), .B0(new_n10239_), .Y(new_n10240_));
  XOR2X1   g09984(.A(new_n10240_), .B(\a[23] ), .Y(new_n10241_));
  INVX1    g09985(.A(new_n10241_), .Y(new_n10242_));
  INVX1    g09986(.A(new_n10171_), .Y(new_n10243_));
  NOR2X1   g09987(.A(new_n10180_), .B(new_n10175_), .Y(new_n10244_));
  AOI21X1  g09988(.A0(new_n10181_), .A1(new_n10243_), .B0(new_n10244_), .Y(new_n10245_));
  XOR2X1   g09989(.A(new_n10245_), .B(new_n10242_), .Y(new_n10246_));
  AOI22X1  g09990(.A0(new_n1814_), .A1(\b[53] ), .B0(new_n1813_), .B1(\b[52] ), .Y(new_n10247_));
  OAI21X1  g09991(.A0(new_n1812_), .A1(new_n5787_), .B0(new_n10247_), .Y(new_n10248_));
  AOI21X1  g09992(.A0(new_n5786_), .A1(new_n1617_), .B0(new_n10248_), .Y(new_n10249_));
  XOR2X1   g09993(.A(new_n10249_), .B(\a[26] ), .Y(new_n10250_));
  NOR2X1   g09994(.A(new_n10065_), .B(new_n10062_), .Y(new_n10251_));
  INVX1    g09995(.A(new_n10170_), .Y(new_n10252_));
  AOI21X1  g09996(.A0(new_n10252_), .A1(new_n10066_), .B0(new_n10251_), .Y(new_n10253_));
  XOR2X1   g09997(.A(new_n10253_), .B(new_n10250_), .Y(new_n10254_));
  AND2X1   g09998(.A(new_n10155_), .B(new_n10070_), .Y(new_n10255_));
  INVX1    g09999(.A(new_n10255_), .Y(new_n10256_));
  INVX1    g10000(.A(new_n10156_), .Y(new_n10257_));
  OAI21X1  g10001(.A0(new_n10160_), .A1(new_n10257_), .B0(new_n10256_), .Y(new_n10258_));
  INVX1    g10002(.A(new_n10258_), .Y(new_n10259_));
  NOR3X1   g10003(.A(new_n2401_), .B(new_n2259_), .C(new_n4674_), .Y(new_n10260_));
  OAI22X1  g10004(.A0(new_n2263_), .A1(new_n5039_), .B0(new_n2262_), .B1(new_n4693_), .Y(new_n10261_));
  OR2X1    g10005(.A(new_n10261_), .B(new_n10260_), .Y(new_n10262_));
  AOI21X1  g10006(.A0(new_n4673_), .A1(new_n2260_), .B0(new_n10262_), .Y(new_n10263_));
  XOR2X1   g10007(.A(new_n10263_), .B(\a[32] ), .Y(new_n10264_));
  XOR2X1   g10008(.A(new_n10264_), .B(new_n10259_), .Y(new_n10265_));
  AOI22X1  g10009(.A0(new_n2813_), .A1(\b[44] ), .B0(new_n2812_), .B1(\b[43] ), .Y(new_n10266_));
  OAI21X1  g10010(.A0(new_n2946_), .A1(new_n4012_), .B0(new_n10266_), .Y(new_n10267_));
  AOI21X1  g10011(.A0(new_n4178_), .A1(new_n2652_), .B0(new_n10267_), .Y(new_n10268_));
  XOR2X1   g10012(.A(new_n10268_), .B(\a[35] ), .Y(new_n10269_));
  INVX1    g10013(.A(new_n10076_), .Y(new_n10270_));
  NAND2X1  g10014(.A(new_n10153_), .B(new_n10270_), .Y(new_n10271_));
  OAI21X1  g10015(.A0(new_n10154_), .A1(new_n10074_), .B0(new_n10271_), .Y(new_n10272_));
  AOI22X1  g10016(.A0(new_n3204_), .A1(\b[41] ), .B0(new_n3203_), .B1(\b[40] ), .Y(new_n10273_));
  OAI21X1  g10017(.A0(new_n3321_), .A1(new_n3723_), .B0(new_n10273_), .Y(new_n10274_));
  AOI21X1  g10018(.A0(new_n3722_), .A1(new_n3080_), .B0(new_n10274_), .Y(new_n10275_));
  XOR2X1   g10019(.A(new_n10275_), .B(new_n3078_), .Y(new_n10276_));
  OAI21X1  g10020(.A0(new_n10084_), .A1(new_n10082_), .B0(new_n10151_), .Y(new_n10277_));
  OAI21X1  g10021(.A0(new_n10152_), .A1(new_n10080_), .B0(new_n10277_), .Y(new_n10278_));
  AND2X1   g10022(.A(new_n10147_), .B(new_n10097_), .Y(new_n10279_));
  INVX1    g10023(.A(new_n10279_), .Y(new_n10280_));
  OAI21X1  g10024(.A0(new_n10148_), .A1(new_n10093_), .B0(new_n10280_), .Y(new_n10281_));
  INVX1    g10025(.A(new_n10281_), .Y(new_n10282_));
  NOR2X1   g10026(.A(new_n10130_), .B(new_n10127_), .Y(new_n10283_));
  INVX1    g10027(.A(new_n10283_), .Y(new_n10284_));
  INVX1    g10028(.A(new_n10131_), .Y(new_n10285_));
  OAI21X1  g10029(.A0(new_n10135_), .A1(new_n10285_), .B0(new_n10284_), .Y(new_n10286_));
  AOI22X1  g10030(.A0(new_n5430_), .A1(\b[26] ), .B0(new_n5427_), .B1(\b[25] ), .Y(new_n10287_));
  OAI21X1  g10031(.A0(new_n5891_), .A1(new_n1588_), .B0(new_n10287_), .Y(new_n10288_));
  AOI21X1  g10032(.A0(new_n5425_), .A1(new_n1783_), .B0(new_n10288_), .Y(new_n10289_));
  XOR2X1   g10033(.A(new_n10289_), .B(new_n5423_), .Y(new_n10290_));
  NOR2X1   g10034(.A(new_n10121_), .B(new_n10119_), .Y(new_n10291_));
  NAND2X1  g10035(.A(new_n10121_), .B(new_n10119_), .Y(new_n10292_));
  OAI21X1  g10036(.A0(new_n10126_), .A1(new_n10291_), .B0(new_n10292_), .Y(new_n10293_));
  INVX1    g10037(.A(new_n10099_), .Y(new_n10294_));
  NOR2X1   g10038(.A(new_n10101_), .B(new_n10294_), .Y(new_n10295_));
  NOR2X1   g10039(.A(new_n10107_), .B(new_n10102_), .Y(new_n10296_));
  NOR2X1   g10040(.A(new_n10296_), .B(new_n10295_), .Y(new_n10297_));
  INVX1    g10041(.A(new_n10297_), .Y(new_n10298_));
  AOI22X1  g10042(.A0(new_n7818_), .A1(\b[13] ), .B0(new_n7817_), .B1(\b[14] ), .Y(new_n10299_));
  XOR2X1   g10043(.A(new_n10299_), .B(new_n10099_), .Y(new_n10300_));
  AOI22X1  g10044(.A0(new_n7192_), .A1(\b[17] ), .B0(new_n7189_), .B1(\b[16] ), .Y(new_n10301_));
  OAI21X1  g10045(.A0(new_n7627_), .A1(new_n977_), .B0(new_n10301_), .Y(new_n10302_));
  AOI21X1  g10046(.A0(new_n7187_), .A1(new_n976_), .B0(new_n10302_), .Y(new_n10303_));
  XOR2X1   g10047(.A(new_n10303_), .B(\a[62] ), .Y(new_n10304_));
  XOR2X1   g10048(.A(new_n10304_), .B(new_n10300_), .Y(new_n10305_));
  XOR2X1   g10049(.A(new_n10305_), .B(new_n10298_), .Y(new_n10306_));
  AOI22X1  g10050(.A0(new_n6603_), .A1(\b[20] ), .B0(new_n6600_), .B1(\b[19] ), .Y(new_n10307_));
  OAI21X1  g10051(.A0(new_n6804_), .A1(new_n1115_), .B0(new_n10307_), .Y(new_n10308_));
  AOI21X1  g10052(.A0(new_n6598_), .A1(new_n1217_), .B0(new_n10308_), .Y(new_n10309_));
  XOR2X1   g10053(.A(new_n10309_), .B(\a[59] ), .Y(new_n10310_));
  XOR2X1   g10054(.A(new_n10310_), .B(new_n10306_), .Y(new_n10311_));
  AND2X1   g10055(.A(new_n10112_), .B(new_n10108_), .Y(new_n10312_));
  OR2X1    g10056(.A(new_n10112_), .B(new_n10108_), .Y(new_n10313_));
  OAI21X1  g10057(.A0(new_n10117_), .A1(new_n10312_), .B0(new_n10313_), .Y(new_n10314_));
  XOR2X1   g10058(.A(new_n10314_), .B(new_n10311_), .Y(new_n10315_));
  AOI22X1  g10059(.A0(new_n6438_), .A1(\b[23] ), .B0(new_n6437_), .B1(\b[22] ), .Y(new_n10316_));
  OAI21X1  g10060(.A0(new_n6436_), .A1(new_n1482_), .B0(new_n10316_), .Y(new_n10317_));
  AOI21X1  g10061(.A0(new_n6023_), .A1(new_n1481_), .B0(new_n10317_), .Y(new_n10318_));
  XOR2X1   g10062(.A(new_n10318_), .B(\a[56] ), .Y(new_n10319_));
  XOR2X1   g10063(.A(new_n10319_), .B(new_n10315_), .Y(new_n10320_));
  XOR2X1   g10064(.A(new_n10320_), .B(new_n10293_), .Y(new_n10321_));
  XOR2X1   g10065(.A(new_n10321_), .B(new_n10290_), .Y(new_n10322_));
  XOR2X1   g10066(.A(new_n10322_), .B(new_n10286_), .Y(new_n10323_));
  AOI22X1  g10067(.A0(new_n4880_), .A1(\b[29] ), .B0(new_n4877_), .B1(\b[28] ), .Y(new_n10324_));
  OAI21X1  g10068(.A0(new_n5291_), .A1(new_n2126_), .B0(new_n10324_), .Y(new_n10325_));
  AOI21X1  g10069(.A0(new_n4875_), .A1(new_n2125_), .B0(new_n10325_), .Y(new_n10326_));
  XOR2X1   g10070(.A(new_n10326_), .B(\a[50] ), .Y(new_n10327_));
  XOR2X1   g10071(.A(new_n10327_), .B(new_n10323_), .Y(new_n10328_));
  OR2X1    g10072(.A(new_n10141_), .B(new_n10136_), .Y(new_n10329_));
  OR2X1    g10073(.A(new_n10146_), .B(new_n10142_), .Y(new_n10330_));
  AND2X1   g10074(.A(new_n10330_), .B(new_n10329_), .Y(new_n10331_));
  XOR2X1   g10075(.A(new_n10331_), .B(new_n10328_), .Y(new_n10332_));
  AOI22X1  g10076(.A0(new_n4572_), .A1(\b[32] ), .B0(new_n4571_), .B1(\b[31] ), .Y(new_n10333_));
  OAI21X1  g10077(.A0(new_n4740_), .A1(new_n2356_), .B0(new_n10333_), .Y(new_n10334_));
  AOI21X1  g10078(.A0(new_n4375_), .A1(new_n2495_), .B0(new_n10334_), .Y(new_n10335_));
  XOR2X1   g10079(.A(new_n10335_), .B(\a[47] ), .Y(new_n10336_));
  XOR2X1   g10080(.A(new_n10336_), .B(new_n10332_), .Y(new_n10337_));
  XOR2X1   g10081(.A(new_n10337_), .B(new_n10282_), .Y(new_n10338_));
  AOI22X1  g10082(.A0(new_n4095_), .A1(\b[35] ), .B0(new_n4094_), .B1(\b[34] ), .Y(new_n10339_));
  OAI21X1  g10083(.A0(new_n4233_), .A1(new_n2893_), .B0(new_n10339_), .Y(new_n10340_));
  AOI21X1  g10084(.A0(new_n3901_), .A1(new_n2892_), .B0(new_n10340_), .Y(new_n10341_));
  XOR2X1   g10085(.A(new_n10341_), .B(\a[44] ), .Y(new_n10342_));
  XOR2X1   g10086(.A(new_n10342_), .B(new_n10338_), .Y(new_n10343_));
  INVX1    g10087(.A(new_n10343_), .Y(new_n10344_));
  AND2X1   g10088(.A(new_n10149_), .B(new_n9991_), .Y(new_n10345_));
  AOI21X1  g10089(.A0(new_n10150_), .A1(new_n10089_), .B0(new_n10345_), .Y(new_n10346_));
  XOR2X1   g10090(.A(new_n10346_), .B(new_n10344_), .Y(new_n10347_));
  AOI22X1  g10091(.A0(new_n3652_), .A1(\b[38] ), .B0(new_n3651_), .B1(\b[37] ), .Y(new_n10348_));
  OAI21X1  g10092(.A0(new_n3778_), .A1(new_n3276_), .B0(new_n10348_), .Y(new_n10349_));
  AOI21X1  g10093(.A0(new_n3480_), .A1(new_n3275_), .B0(new_n10349_), .Y(new_n10350_));
  XOR2X1   g10094(.A(new_n10350_), .B(\a[41] ), .Y(new_n10351_));
  XOR2X1   g10095(.A(new_n10351_), .B(new_n10347_), .Y(new_n10352_));
  XOR2X1   g10096(.A(new_n10352_), .B(new_n10278_), .Y(new_n10353_));
  XOR2X1   g10097(.A(new_n10353_), .B(new_n10276_), .Y(new_n10354_));
  XOR2X1   g10098(.A(new_n10354_), .B(new_n10272_), .Y(new_n10355_));
  XOR2X1   g10099(.A(new_n10355_), .B(new_n10269_), .Y(new_n10356_));
  XOR2X1   g10100(.A(new_n10356_), .B(new_n10265_), .Y(new_n10357_));
  INVX1    g10101(.A(new_n10161_), .Y(new_n10358_));
  NOR2X1   g10102(.A(new_n10168_), .B(new_n10164_), .Y(new_n10359_));
  AOI21X1  g10103(.A0(new_n10169_), .A1(new_n10358_), .B0(new_n10359_), .Y(new_n10360_));
  OAI22X1  g10104(.A0(new_n1913_), .A1(new_n5234_), .B0(new_n1910_), .B1(new_n5237_), .Y(new_n10361_));
  AOI21X1  g10105(.A0(new_n2045_), .A1(\b[48] ), .B0(new_n10361_), .Y(new_n10362_));
  OAI21X1  g10106(.A0(new_n9725_), .A1(new_n2043_), .B0(new_n10362_), .Y(new_n10363_));
  XOR2X1   g10107(.A(new_n10363_), .B(new_n1911_), .Y(new_n10364_));
  XOR2X1   g10108(.A(new_n10364_), .B(new_n10360_), .Y(new_n10365_));
  XOR2X1   g10109(.A(new_n10365_), .B(new_n10357_), .Y(new_n10366_));
  XOR2X1   g10110(.A(new_n10366_), .B(new_n10254_), .Y(new_n10367_));
  XOR2X1   g10111(.A(new_n10367_), .B(new_n10246_), .Y(new_n10368_));
  XOR2X1   g10112(.A(new_n10368_), .B(new_n10237_), .Y(new_n10369_));
  INVX1    g10113(.A(new_n10369_), .Y(new_n10370_));
  OAI21X1  g10114(.A0(new_n10226_), .A1(new_n10225_), .B0(new_n10224_), .Y(new_n10371_));
  AOI21X1  g10115(.A0(new_n10229_), .A1(new_n10371_), .B0(new_n10370_), .Y(new_n10372_));
  AND2X1   g10116(.A(new_n10371_), .B(new_n10370_), .Y(new_n10373_));
  AOI21X1  g10117(.A0(new_n10373_), .A1(new_n10229_), .B0(new_n10372_), .Y(new_n10374_));
  XOR2X1   g10118(.A(new_n10374_), .B(new_n10220_), .Y(new_n10375_));
  XOR2X1   g10119(.A(new_n10375_), .B(new_n10215_), .Y(new_n10376_));
  XOR2X1   g10120(.A(new_n10376_), .B(new_n10213_), .Y(\f[77] ));
  NOR2X1   g10121(.A(new_n10372_), .B(new_n10228_), .Y(new_n10378_));
  AOI22X1  g10122(.A0(new_n1017_), .A1(\b[63] ), .B0(new_n1016_), .B1(\b[62] ), .Y(new_n10379_));
  OAI21X1  g10123(.A0(new_n1015_), .A1(new_n7748_), .B0(new_n10379_), .Y(new_n10380_));
  AOI21X1  g10124(.A0(new_n7747_), .A1(new_n882_), .B0(new_n10380_), .Y(new_n10381_));
  XOR2X1   g10125(.A(new_n10381_), .B(\a[17] ), .Y(new_n10382_));
  XOR2X1   g10126(.A(new_n10382_), .B(new_n10378_), .Y(new_n10383_));
  AOI22X1  g10127(.A0(new_n1263_), .A1(\b[60] ), .B0(new_n1262_), .B1(\b[59] ), .Y(new_n10384_));
  OAI21X1  g10128(.A0(new_n1261_), .A1(new_n6930_), .B0(new_n10384_), .Y(new_n10385_));
  AOI21X1  g10129(.A0(new_n6951_), .A1(new_n1075_), .B0(new_n10385_), .Y(new_n10386_));
  XOR2X1   g10130(.A(new_n10386_), .B(\a[20] ), .Y(new_n10387_));
  INVX1    g10131(.A(new_n10387_), .Y(new_n10388_));
  NOR2X1   g10132(.A(new_n10236_), .B(new_n10233_), .Y(new_n10389_));
  AOI21X1  g10133(.A0(new_n10368_), .A1(new_n10237_), .B0(new_n10389_), .Y(new_n10390_));
  XOR2X1   g10134(.A(new_n10390_), .B(new_n10388_), .Y(new_n10391_));
  NOR2X1   g10135(.A(new_n10245_), .B(new_n10241_), .Y(new_n10392_));
  NOR2X1   g10136(.A(new_n10367_), .B(new_n10246_), .Y(new_n10393_));
  OR2X1    g10137(.A(new_n10393_), .B(new_n10392_), .Y(new_n10394_));
  AOI22X1  g10138(.A0(new_n1526_), .A1(\b[57] ), .B0(new_n1525_), .B1(\b[56] ), .Y(new_n10395_));
  OAI21X1  g10139(.A0(new_n1524_), .A1(new_n6523_), .B0(new_n10395_), .Y(new_n10396_));
  AOI21X1  g10140(.A0(new_n6522_), .A1(new_n1347_), .B0(new_n10396_), .Y(new_n10397_));
  XOR2X1   g10141(.A(new_n10397_), .B(\a[23] ), .Y(new_n10398_));
  XOR2X1   g10142(.A(new_n10398_), .B(new_n10394_), .Y(new_n10399_));
  AOI22X1  g10143(.A0(new_n1814_), .A1(\b[54] ), .B0(new_n1813_), .B1(\b[53] ), .Y(new_n10400_));
  OAI21X1  g10144(.A0(new_n1812_), .A1(new_n5808_), .B0(new_n10400_), .Y(new_n10401_));
  AOI21X1  g10145(.A0(new_n5807_), .A1(new_n1617_), .B0(new_n10401_), .Y(new_n10402_));
  XOR2X1   g10146(.A(new_n10402_), .B(\a[26] ), .Y(new_n10403_));
  INVX1    g10147(.A(new_n10403_), .Y(new_n10404_));
  NOR2X1   g10148(.A(new_n10253_), .B(new_n10250_), .Y(new_n10405_));
  INVX1    g10149(.A(new_n10366_), .Y(new_n10406_));
  AOI21X1  g10150(.A0(new_n10406_), .A1(new_n10254_), .B0(new_n10405_), .Y(new_n10407_));
  XOR2X1   g10151(.A(new_n10407_), .B(new_n10404_), .Y(new_n10408_));
  AOI22X1  g10152(.A0(new_n2163_), .A1(\b[51] ), .B0(new_n2162_), .B1(\b[50] ), .Y(new_n10409_));
  OAI21X1  g10153(.A0(new_n2161_), .A1(new_n5237_), .B0(new_n10409_), .Y(new_n10410_));
  AOI21X1  g10154(.A0(new_n5236_), .A1(new_n1907_), .B0(new_n10410_), .Y(new_n10411_));
  XOR2X1   g10155(.A(new_n10411_), .B(\a[29] ), .Y(new_n10412_));
  INVX1    g10156(.A(new_n10357_), .Y(new_n10413_));
  NOR2X1   g10157(.A(new_n10364_), .B(new_n10360_), .Y(new_n10414_));
  AOI21X1  g10158(.A0(new_n10365_), .A1(new_n10413_), .B0(new_n10414_), .Y(new_n10415_));
  XOR2X1   g10159(.A(new_n10415_), .B(new_n10412_), .Y(new_n10416_));
  INVX1    g10160(.A(new_n10416_), .Y(new_n10417_));
  AND2X1   g10161(.A(new_n10352_), .B(new_n10278_), .Y(new_n10418_));
  AOI21X1  g10162(.A0(new_n10353_), .A1(new_n10276_), .B0(new_n10418_), .Y(new_n10419_));
  INVX1    g10163(.A(new_n10419_), .Y(new_n10420_));
  NOR2X1   g10164(.A(new_n10346_), .B(new_n10343_), .Y(new_n10421_));
  INVX1    g10165(.A(new_n10421_), .Y(new_n10422_));
  OAI21X1  g10166(.A0(new_n10351_), .A1(new_n10347_), .B0(new_n10422_), .Y(new_n10423_));
  NOR2X1   g10167(.A(new_n10337_), .B(new_n10282_), .Y(new_n10424_));
  INVX1    g10168(.A(new_n10424_), .Y(new_n10425_));
  INVX1    g10169(.A(new_n10338_), .Y(new_n10426_));
  OAI21X1  g10170(.A0(new_n10342_), .A1(new_n10426_), .B0(new_n10425_), .Y(new_n10427_));
  NOR2X1   g10171(.A(new_n10331_), .B(new_n10328_), .Y(new_n10428_));
  INVX1    g10172(.A(new_n10428_), .Y(new_n10429_));
  INVX1    g10173(.A(new_n10332_), .Y(new_n10430_));
  OR2X1    g10174(.A(new_n10336_), .B(new_n10430_), .Y(new_n10431_));
  AND2X1   g10175(.A(new_n10431_), .B(new_n10429_), .Y(new_n10432_));
  INVX1    g10176(.A(new_n10432_), .Y(new_n10433_));
  INVX1    g10177(.A(new_n10311_), .Y(new_n10434_));
  NOR2X1   g10178(.A(new_n10319_), .B(new_n10315_), .Y(new_n10435_));
  AOI21X1  g10179(.A0(new_n10314_), .A1(new_n10434_), .B0(new_n10435_), .Y(new_n10436_));
  AOI22X1  g10180(.A0(new_n7818_), .A1(\b[14] ), .B0(new_n7817_), .B1(\b[15] ), .Y(new_n10437_));
  XOR2X1   g10181(.A(new_n10437_), .B(new_n665_), .Y(new_n10438_));
  XOR2X1   g10182(.A(new_n10438_), .B(new_n10294_), .Y(new_n10439_));
  AOI22X1  g10183(.A0(new_n7192_), .A1(\b[18] ), .B0(new_n7189_), .B1(\b[17] ), .Y(new_n10440_));
  OAI21X1  g10184(.A0(new_n7627_), .A1(new_n974_), .B0(new_n10440_), .Y(new_n10441_));
  AOI21X1  g10185(.A0(new_n7187_), .A1(new_n1042_), .B0(new_n10441_), .Y(new_n10442_));
  XOR2X1   g10186(.A(new_n10442_), .B(\a[62] ), .Y(new_n10443_));
  XOR2X1   g10187(.A(new_n10443_), .B(new_n10439_), .Y(new_n10444_));
  OR2X1    g10188(.A(new_n10299_), .B(new_n10294_), .Y(new_n10445_));
  OAI21X1  g10189(.A0(new_n10304_), .A1(new_n10300_), .B0(new_n10445_), .Y(new_n10446_));
  XOR2X1   g10190(.A(new_n10446_), .B(new_n10444_), .Y(new_n10447_));
  AOI22X1  g10191(.A0(new_n6603_), .A1(\b[21] ), .B0(new_n6600_), .B1(\b[20] ), .Y(new_n10448_));
  OAI21X1  g10192(.A0(new_n6804_), .A1(new_n1300_), .B0(new_n10448_), .Y(new_n10449_));
  AOI21X1  g10193(.A0(new_n6598_), .A1(new_n1299_), .B0(new_n10449_), .Y(new_n10450_));
  XOR2X1   g10194(.A(new_n10450_), .B(\a[59] ), .Y(new_n10451_));
  XOR2X1   g10195(.A(new_n10451_), .B(new_n10447_), .Y(new_n10452_));
  AND2X1   g10196(.A(new_n10305_), .B(new_n10298_), .Y(new_n10453_));
  INVX1    g10197(.A(new_n10310_), .Y(new_n10454_));
  AOI21X1  g10198(.A0(new_n10454_), .A1(new_n10306_), .B0(new_n10453_), .Y(new_n10455_));
  XOR2X1   g10199(.A(new_n10455_), .B(new_n10452_), .Y(new_n10456_));
  AOI22X1  g10200(.A0(new_n6438_), .A1(\b[24] ), .B0(new_n6437_), .B1(\b[23] ), .Y(new_n10457_));
  OAI21X1  g10201(.A0(new_n6436_), .A1(new_n1479_), .B0(new_n10457_), .Y(new_n10458_));
  AOI21X1  g10202(.A0(new_n6023_), .A1(new_n1572_), .B0(new_n10458_), .Y(new_n10459_));
  XOR2X1   g10203(.A(new_n10459_), .B(new_n6019_), .Y(new_n10460_));
  NOR2X1   g10204(.A(new_n10460_), .B(new_n10456_), .Y(new_n10461_));
  AND2X1   g10205(.A(new_n10460_), .B(new_n10456_), .Y(new_n10462_));
  NOR3X1   g10206(.A(new_n10462_), .B(new_n10461_), .C(new_n10436_), .Y(new_n10463_));
  NOR2X1   g10207(.A(new_n10463_), .B(new_n10462_), .Y(new_n10464_));
  INVX1    g10208(.A(new_n10464_), .Y(new_n10465_));
  OAI22X1  g10209(.A0(new_n10465_), .A1(new_n10461_), .B0(new_n10463_), .B1(new_n10436_), .Y(new_n10466_));
  AOI22X1  g10210(.A0(new_n5430_), .A1(\b[27] ), .B0(new_n5427_), .B1(\b[26] ), .Y(new_n10467_));
  OAI21X1  g10211(.A0(new_n5891_), .A1(new_n1880_), .B0(new_n10467_), .Y(new_n10468_));
  AOI21X1  g10212(.A0(new_n5425_), .A1(new_n1879_), .B0(new_n10468_), .Y(new_n10469_));
  XOR2X1   g10213(.A(new_n10469_), .B(\a[53] ), .Y(new_n10470_));
  XOR2X1   g10214(.A(new_n10470_), .B(new_n10466_), .Y(new_n10471_));
  AND2X1   g10215(.A(new_n10320_), .B(new_n10293_), .Y(new_n10472_));
  AOI21X1  g10216(.A0(new_n10321_), .A1(new_n10290_), .B0(new_n10472_), .Y(new_n10473_));
  XOR2X1   g10217(.A(new_n10473_), .B(new_n10471_), .Y(new_n10474_));
  AOI22X1  g10218(.A0(new_n4880_), .A1(\b[30] ), .B0(new_n4877_), .B1(\b[29] ), .Y(new_n10475_));
  OAI21X1  g10219(.A0(new_n5291_), .A1(new_n2231_), .B0(new_n10475_), .Y(new_n10476_));
  AOI21X1  g10220(.A0(new_n4875_), .A1(new_n2230_), .B0(new_n10476_), .Y(new_n10477_));
  XOR2X1   g10221(.A(new_n10477_), .B(\a[50] ), .Y(new_n10478_));
  XOR2X1   g10222(.A(new_n10478_), .B(new_n10474_), .Y(new_n10479_));
  AND2X1   g10223(.A(new_n10322_), .B(new_n10286_), .Y(new_n10480_));
  INVX1    g10224(.A(new_n10327_), .Y(new_n10481_));
  AOI21X1  g10225(.A0(new_n10481_), .A1(new_n10323_), .B0(new_n10480_), .Y(new_n10482_));
  XOR2X1   g10226(.A(new_n10482_), .B(new_n10479_), .Y(new_n10483_));
  AOI22X1  g10227(.A0(new_n4572_), .A1(\b[33] ), .B0(new_n4571_), .B1(\b[32] ), .Y(new_n10484_));
  OAI21X1  g10228(.A0(new_n4740_), .A1(new_n2615_), .B0(new_n10484_), .Y(new_n10485_));
  AOI21X1  g10229(.A0(new_n4375_), .A1(new_n2614_), .B0(new_n10485_), .Y(new_n10486_));
  XOR2X1   g10230(.A(new_n10486_), .B(\a[47] ), .Y(new_n10487_));
  XOR2X1   g10231(.A(new_n10487_), .B(new_n10483_), .Y(new_n10488_));
  XOR2X1   g10232(.A(new_n10488_), .B(new_n10433_), .Y(new_n10489_));
  AOI22X1  g10233(.A0(new_n4095_), .A1(\b[36] ), .B0(new_n4094_), .B1(\b[35] ), .Y(new_n10490_));
  OAI21X1  g10234(.A0(new_n4233_), .A1(new_n2890_), .B0(new_n10490_), .Y(new_n10491_));
  AOI21X1  g10235(.A0(new_n3901_), .A1(new_n3015_), .B0(new_n10491_), .Y(new_n10492_));
  XOR2X1   g10236(.A(new_n10492_), .B(\a[44] ), .Y(new_n10493_));
  XOR2X1   g10237(.A(new_n10493_), .B(new_n10489_), .Y(new_n10494_));
  XOR2X1   g10238(.A(new_n10494_), .B(new_n10427_), .Y(new_n10495_));
  AOI22X1  g10239(.A0(new_n3652_), .A1(\b[39] ), .B0(new_n3651_), .B1(\b[38] ), .Y(new_n10496_));
  OAI21X1  g10240(.A0(new_n3778_), .A1(new_n3413_), .B0(new_n10496_), .Y(new_n10497_));
  AOI21X1  g10241(.A0(new_n3480_), .A1(new_n3412_), .B0(new_n10497_), .Y(new_n10498_));
  XOR2X1   g10242(.A(new_n10498_), .B(\a[41] ), .Y(new_n10499_));
  XOR2X1   g10243(.A(new_n10499_), .B(new_n10495_), .Y(new_n10500_));
  XOR2X1   g10244(.A(new_n10500_), .B(new_n10423_), .Y(new_n10501_));
  AOI22X1  g10245(.A0(new_n3204_), .A1(\b[42] ), .B0(new_n3203_), .B1(\b[41] ), .Y(new_n10502_));
  OAI21X1  g10246(.A0(new_n3321_), .A1(new_n3720_), .B0(new_n10502_), .Y(new_n10503_));
  AOI21X1  g10247(.A0(new_n3860_), .A1(new_n3080_), .B0(new_n10503_), .Y(new_n10504_));
  XOR2X1   g10248(.A(new_n10504_), .B(\a[38] ), .Y(new_n10505_));
  XOR2X1   g10249(.A(new_n10505_), .B(new_n10501_), .Y(new_n10506_));
  XOR2X1   g10250(.A(new_n10506_), .B(new_n10420_), .Y(new_n10507_));
  AOI22X1  g10251(.A0(new_n2813_), .A1(\b[45] ), .B0(new_n2812_), .B1(\b[44] ), .Y(new_n10508_));
  OAI21X1  g10252(.A0(new_n2946_), .A1(new_n4339_), .B0(new_n10508_), .Y(new_n10509_));
  AOI21X1  g10253(.A0(new_n4338_), .A1(new_n2652_), .B0(new_n10509_), .Y(new_n10510_));
  XOR2X1   g10254(.A(new_n10510_), .B(\a[35] ), .Y(new_n10511_));
  XOR2X1   g10255(.A(new_n10511_), .B(new_n10507_), .Y(new_n10512_));
  INVX1    g10256(.A(new_n10512_), .Y(new_n10513_));
  INVX1    g10257(.A(new_n10269_), .Y(new_n10514_));
  AND2X1   g10258(.A(new_n10354_), .B(new_n10272_), .Y(new_n10515_));
  AOI21X1  g10259(.A0(new_n10355_), .A1(new_n10514_), .B0(new_n10515_), .Y(new_n10516_));
  XOR2X1   g10260(.A(new_n10516_), .B(new_n10513_), .Y(new_n10517_));
  NOR2X1   g10261(.A(new_n10264_), .B(new_n10259_), .Y(new_n10518_));
  INVX1    g10262(.A(new_n10518_), .Y(new_n10519_));
  INVX1    g10263(.A(new_n10265_), .Y(new_n10520_));
  OAI21X1  g10264(.A0(new_n10356_), .A1(new_n10520_), .B0(new_n10519_), .Y(new_n10521_));
  AOI22X1  g10265(.A0(new_n2545_), .A1(\b[48] ), .B0(new_n2544_), .B1(\b[47] ), .Y(new_n10522_));
  OAI21X1  g10266(.A0(new_n2543_), .A1(new_n4693_), .B0(new_n10522_), .Y(new_n10523_));
  AOI21X1  g10267(.A0(new_n4692_), .A1(new_n2260_), .B0(new_n10523_), .Y(new_n10524_));
  XOR2X1   g10268(.A(new_n10524_), .B(\a[32] ), .Y(new_n10525_));
  XOR2X1   g10269(.A(new_n10525_), .B(new_n10521_), .Y(new_n10526_));
  XOR2X1   g10270(.A(new_n10526_), .B(new_n10517_), .Y(new_n10527_));
  XOR2X1   g10271(.A(new_n10527_), .B(new_n10417_), .Y(new_n10528_));
  XOR2X1   g10272(.A(new_n10528_), .B(new_n10408_), .Y(new_n10529_));
  XOR2X1   g10273(.A(new_n10529_), .B(new_n10399_), .Y(new_n10530_));
  XOR2X1   g10274(.A(new_n10530_), .B(new_n10391_), .Y(new_n10531_));
  XOR2X1   g10275(.A(new_n10531_), .B(new_n10383_), .Y(new_n10532_));
  NOR2X1   g10276(.A(new_n10219_), .B(new_n10217_), .Y(new_n10533_));
  AOI21X1  g10277(.A0(new_n10374_), .A1(new_n10220_), .B0(new_n10533_), .Y(new_n10534_));
  XOR2X1   g10278(.A(new_n10534_), .B(new_n10532_), .Y(new_n10535_));
  AND2X1   g10279(.A(new_n10375_), .B(new_n10215_), .Y(new_n10536_));
  INVX1    g10280(.A(new_n10536_), .Y(new_n10537_));
  OAI21X1  g10281(.A0(new_n10212_), .A1(new_n10211_), .B0(new_n10376_), .Y(new_n10538_));
  AND2X1   g10282(.A(new_n10538_), .B(new_n10537_), .Y(new_n10539_));
  XOR2X1   g10283(.A(new_n10539_), .B(new_n10535_), .Y(\f[78] ));
  NOR2X1   g10284(.A(new_n10390_), .B(new_n10387_), .Y(new_n10541_));
  NOR2X1   g10285(.A(new_n10530_), .B(new_n10391_), .Y(new_n10542_));
  NOR2X1   g10286(.A(new_n10542_), .B(new_n10541_), .Y(new_n10543_));
  OAI22X1  g10287(.A0(new_n1015_), .A1(new_n7745_), .B0(new_n1067_), .B1(new_n7772_), .Y(new_n10544_));
  AOI21X1  g10288(.A0(new_n7775_), .A1(new_n882_), .B0(new_n10544_), .Y(new_n10545_));
  XOR2X1   g10289(.A(new_n10545_), .B(\a[17] ), .Y(new_n10546_));
  XOR2X1   g10290(.A(new_n10546_), .B(new_n10543_), .Y(new_n10547_));
  AOI22X1  g10291(.A0(new_n1263_), .A1(\b[61] ), .B0(new_n1262_), .B1(\b[60] ), .Y(new_n10548_));
  OAI21X1  g10292(.A0(new_n1261_), .A1(new_n7339_), .B0(new_n10548_), .Y(new_n10549_));
  AOI21X1  g10293(.A0(new_n7338_), .A1(new_n1075_), .B0(new_n10549_), .Y(new_n10550_));
  XOR2X1   g10294(.A(new_n10550_), .B(\a[20] ), .Y(new_n10551_));
  INVX1    g10295(.A(new_n10551_), .Y(new_n10552_));
  INVX1    g10296(.A(new_n10398_), .Y(new_n10553_));
  NOR2X1   g10297(.A(new_n10528_), .B(new_n10408_), .Y(new_n10554_));
  AND2X1   g10298(.A(new_n10528_), .B(new_n10408_), .Y(new_n10555_));
  NOR3X1   g10299(.A(new_n10555_), .B(new_n10554_), .C(new_n10399_), .Y(new_n10556_));
  AOI21X1  g10300(.A0(new_n10553_), .A1(new_n10394_), .B0(new_n10556_), .Y(new_n10557_));
  XOR2X1   g10301(.A(new_n10557_), .B(new_n10552_), .Y(new_n10558_));
  NOR2X1   g10302(.A(new_n10407_), .B(new_n10403_), .Y(new_n10559_));
  NOR2X1   g10303(.A(new_n10554_), .B(new_n10559_), .Y(new_n10560_));
  OAI22X1  g10304(.A0(new_n1353_), .A1(new_n6930_), .B0(new_n1350_), .B1(new_n6933_), .Y(new_n10561_));
  AOI21X1  g10305(.A0(new_n1430_), .A1(\b[56] ), .B0(new_n10561_), .Y(new_n10562_));
  OAI21X1  g10306(.A0(new_n8540_), .A1(new_n1428_), .B0(new_n10562_), .Y(new_n10563_));
  XOR2X1   g10307(.A(new_n10563_), .B(new_n1351_), .Y(new_n10564_));
  XOR2X1   g10308(.A(new_n10564_), .B(new_n10560_), .Y(new_n10565_));
  INVX1    g10309(.A(new_n10565_), .Y(new_n10566_));
  AOI22X1  g10310(.A0(new_n1814_), .A1(\b[55] ), .B0(new_n1813_), .B1(\b[54] ), .Y(new_n10567_));
  OAI21X1  g10311(.A0(new_n1812_), .A1(new_n6151_), .B0(new_n10567_), .Y(new_n10568_));
  AOI21X1  g10312(.A0(new_n6150_), .A1(new_n1617_), .B0(new_n10568_), .Y(new_n10569_));
  XOR2X1   g10313(.A(new_n10569_), .B(\a[26] ), .Y(new_n10570_));
  INVX1    g10314(.A(new_n10570_), .Y(new_n10571_));
  NOR2X1   g10315(.A(new_n10415_), .B(new_n10412_), .Y(new_n10572_));
  AOI21X1  g10316(.A0(new_n10527_), .A1(new_n10416_), .B0(new_n10572_), .Y(new_n10573_));
  XOR2X1   g10317(.A(new_n10573_), .B(new_n10571_), .Y(new_n10574_));
  AOI22X1  g10318(.A0(new_n2163_), .A1(\b[52] ), .B0(new_n2162_), .B1(\b[51] ), .Y(new_n10575_));
  OAI21X1  g10319(.A0(new_n2161_), .A1(new_n5234_), .B0(new_n10575_), .Y(new_n10576_));
  AOI21X1  g10320(.A0(new_n5590_), .A1(new_n1907_), .B0(new_n10576_), .Y(new_n10577_));
  XOR2X1   g10321(.A(new_n10577_), .B(\a[29] ), .Y(new_n10578_));
  INVX1    g10322(.A(new_n10525_), .Y(new_n10579_));
  NOR2X1   g10323(.A(new_n10526_), .B(new_n10517_), .Y(new_n10580_));
  AOI21X1  g10324(.A0(new_n10579_), .A1(new_n10521_), .B0(new_n10580_), .Y(new_n10581_));
  XOR2X1   g10325(.A(new_n10581_), .B(new_n10578_), .Y(new_n10582_));
  INVX1    g10326(.A(new_n10582_), .Y(new_n10583_));
  AOI22X1  g10327(.A0(new_n2545_), .A1(\b[49] ), .B0(new_n2544_), .B1(\b[48] ), .Y(new_n10584_));
  OAI21X1  g10328(.A0(new_n2543_), .A1(new_n5039_), .B0(new_n10584_), .Y(new_n10585_));
  AOI21X1  g10329(.A0(new_n5038_), .A1(new_n2260_), .B0(new_n10585_), .Y(new_n10586_));
  XOR2X1   g10330(.A(new_n10586_), .B(\a[32] ), .Y(new_n10587_));
  INVX1    g10331(.A(new_n10587_), .Y(new_n10588_));
  INVX1    g10332(.A(new_n10511_), .Y(new_n10589_));
  NOR2X1   g10333(.A(new_n10516_), .B(new_n10512_), .Y(new_n10590_));
  AOI21X1  g10334(.A0(new_n10589_), .A1(new_n10507_), .B0(new_n10590_), .Y(new_n10591_));
  XOR2X1   g10335(.A(new_n10591_), .B(new_n10588_), .Y(new_n10592_));
  INVX1    g10336(.A(new_n10495_), .Y(new_n10593_));
  NOR2X1   g10337(.A(new_n10499_), .B(new_n10593_), .Y(new_n10594_));
  INVX1    g10338(.A(new_n10500_), .Y(new_n10595_));
  AOI21X1  g10339(.A0(new_n10595_), .A1(new_n10423_), .B0(new_n10594_), .Y(new_n10596_));
  INVX1    g10340(.A(new_n10596_), .Y(new_n10597_));
  AOI22X1  g10341(.A0(new_n3652_), .A1(\b[40] ), .B0(new_n3651_), .B1(\b[39] ), .Y(new_n10598_));
  OAI21X1  g10342(.A0(new_n3778_), .A1(new_n3575_), .B0(new_n10598_), .Y(new_n10599_));
  AOI21X1  g10343(.A0(new_n3574_), .A1(new_n3480_), .B0(new_n10599_), .Y(new_n10600_));
  XOR2X1   g10344(.A(new_n10600_), .B(\a[41] ), .Y(new_n10601_));
  NOR2X1   g10345(.A(new_n10493_), .B(new_n10489_), .Y(new_n10602_));
  AOI21X1  g10346(.A0(new_n10494_), .A1(new_n10427_), .B0(new_n10602_), .Y(new_n10603_));
  AOI22X1  g10347(.A0(new_n4095_), .A1(\b[37] ), .B0(new_n4094_), .B1(\b[36] ), .Y(new_n10604_));
  OAI21X1  g10348(.A0(new_n4233_), .A1(new_n3156_), .B0(new_n10604_), .Y(new_n10605_));
  AOI21X1  g10349(.A0(new_n3901_), .A1(new_n3155_), .B0(new_n10605_), .Y(new_n10606_));
  XOR2X1   g10350(.A(new_n10606_), .B(\a[44] ), .Y(new_n10607_));
  XOR2X1   g10351(.A(new_n10486_), .B(new_n4568_), .Y(new_n10608_));
  AND2X1   g10352(.A(new_n10608_), .B(new_n10483_), .Y(new_n10609_));
  NOR2X1   g10353(.A(new_n10488_), .B(new_n10432_), .Y(new_n10610_));
  NOR2X1   g10354(.A(new_n10610_), .B(new_n10609_), .Y(new_n10611_));
  NOR2X1   g10355(.A(new_n10443_), .B(new_n10439_), .Y(new_n10612_));
  AOI21X1  g10356(.A0(new_n10446_), .A1(new_n10444_), .B0(new_n10612_), .Y(new_n10613_));
  AOI22X1  g10357(.A0(new_n7818_), .A1(\b[15] ), .B0(new_n7817_), .B1(\b[16] ), .Y(new_n10614_));
  INVX1    g10358(.A(new_n10614_), .Y(new_n10615_));
  NOR2X1   g10359(.A(new_n10437_), .B(\a[14] ), .Y(new_n10616_));
  NOR2X1   g10360(.A(new_n10438_), .B(new_n10099_), .Y(new_n10617_));
  NOR2X1   g10361(.A(new_n10617_), .B(new_n10616_), .Y(new_n10618_));
  XOR2X1   g10362(.A(new_n10618_), .B(new_n10615_), .Y(new_n10619_));
  INVX1    g10363(.A(new_n10619_), .Y(new_n10620_));
  AOI22X1  g10364(.A0(new_n7192_), .A1(\b[19] ), .B0(new_n7189_), .B1(\b[18] ), .Y(new_n10621_));
  OAI21X1  g10365(.A0(new_n7627_), .A1(new_n1118_), .B0(new_n10621_), .Y(new_n10622_));
  AOI21X1  g10366(.A0(new_n7187_), .A1(new_n1117_), .B0(new_n10622_), .Y(new_n10623_));
  XOR2X1   g10367(.A(new_n10623_), .B(\a[62] ), .Y(new_n10624_));
  XOR2X1   g10368(.A(new_n10624_), .B(new_n10620_), .Y(new_n10625_));
  INVX1    g10369(.A(new_n10625_), .Y(new_n10626_));
  XOR2X1   g10370(.A(new_n10626_), .B(new_n10613_), .Y(new_n10627_));
  AOI22X1  g10371(.A0(new_n6603_), .A1(\b[22] ), .B0(new_n6600_), .B1(\b[21] ), .Y(new_n10628_));
  OAI21X1  g10372(.A0(new_n6804_), .A1(new_n1297_), .B0(new_n10628_), .Y(new_n10629_));
  AOI21X1  g10373(.A0(new_n6598_), .A1(new_n1399_), .B0(new_n10629_), .Y(new_n10630_));
  XOR2X1   g10374(.A(new_n10630_), .B(\a[59] ), .Y(new_n10631_));
  XOR2X1   g10375(.A(new_n10631_), .B(new_n10627_), .Y(new_n10632_));
  INVX1    g10376(.A(new_n10451_), .Y(new_n10633_));
  NOR2X1   g10377(.A(new_n10455_), .B(new_n10452_), .Y(new_n10634_));
  AOI21X1  g10378(.A0(new_n10633_), .A1(new_n10447_), .B0(new_n10634_), .Y(new_n10635_));
  XOR2X1   g10379(.A(new_n10635_), .B(new_n10632_), .Y(new_n10636_));
  AOI22X1  g10380(.A0(new_n6438_), .A1(\b[25] ), .B0(new_n6437_), .B1(\b[24] ), .Y(new_n10637_));
  OAI21X1  g10381(.A0(new_n6436_), .A1(new_n1591_), .B0(new_n10637_), .Y(new_n10638_));
  AOI21X1  g10382(.A0(new_n6023_), .A1(new_n1590_), .B0(new_n10638_), .Y(new_n10639_));
  XOR2X1   g10383(.A(new_n10639_), .B(\a[56] ), .Y(new_n10640_));
  XOR2X1   g10384(.A(new_n10640_), .B(new_n10636_), .Y(new_n10641_));
  INVX1    g10385(.A(new_n10641_), .Y(new_n10642_));
  XOR2X1   g10386(.A(new_n10642_), .B(new_n10464_), .Y(new_n10643_));
  AOI22X1  g10387(.A0(new_n5430_), .A1(\b[28] ), .B0(new_n5427_), .B1(\b[27] ), .Y(new_n10644_));
  OAI21X1  g10388(.A0(new_n5891_), .A1(new_n1877_), .B0(new_n10644_), .Y(new_n10645_));
  AOI21X1  g10389(.A0(new_n5425_), .A1(new_n2004_), .B0(new_n10645_), .Y(new_n10646_));
  XOR2X1   g10390(.A(new_n10646_), .B(\a[53] ), .Y(new_n10647_));
  XOR2X1   g10391(.A(new_n10647_), .B(new_n10643_), .Y(new_n10648_));
  INVX1    g10392(.A(new_n10648_), .Y(new_n10649_));
  INVX1    g10393(.A(new_n10470_), .Y(new_n10650_));
  NOR2X1   g10394(.A(new_n10473_), .B(new_n10471_), .Y(new_n10651_));
  AOI21X1  g10395(.A0(new_n10650_), .A1(new_n10466_), .B0(new_n10651_), .Y(new_n10652_));
  XOR2X1   g10396(.A(new_n10652_), .B(new_n10649_), .Y(new_n10653_));
  AOI22X1  g10397(.A0(new_n4880_), .A1(\b[31] ), .B0(new_n4877_), .B1(\b[30] ), .Y(new_n10654_));
  OAI21X1  g10398(.A0(new_n5291_), .A1(new_n2359_), .B0(new_n10654_), .Y(new_n10655_));
  AOI21X1  g10399(.A0(new_n4875_), .A1(new_n2358_), .B0(new_n10655_), .Y(new_n10656_));
  XOR2X1   g10400(.A(new_n10656_), .B(\a[50] ), .Y(new_n10657_));
  XOR2X1   g10401(.A(new_n10657_), .B(new_n10653_), .Y(new_n10658_));
  INVX1    g10402(.A(new_n10658_), .Y(new_n10659_));
  INVX1    g10403(.A(new_n10478_), .Y(new_n10660_));
  NOR2X1   g10404(.A(new_n10482_), .B(new_n10479_), .Y(new_n10661_));
  AOI21X1  g10405(.A0(new_n10660_), .A1(new_n10474_), .B0(new_n10661_), .Y(new_n10662_));
  XOR2X1   g10406(.A(new_n10662_), .B(new_n10659_), .Y(new_n10663_));
  AOI22X1  g10407(.A0(new_n4572_), .A1(\b[34] ), .B0(new_n4571_), .B1(\b[33] ), .Y(new_n10664_));
  OAI21X1  g10408(.A0(new_n4740_), .A1(new_n2612_), .B0(new_n10664_), .Y(new_n10665_));
  AOI21X1  g10409(.A0(new_n4375_), .A1(new_n2759_), .B0(new_n10665_), .Y(new_n10666_));
  XOR2X1   g10410(.A(new_n10666_), .B(\a[47] ), .Y(new_n10667_));
  XOR2X1   g10411(.A(new_n10667_), .B(new_n10663_), .Y(new_n10668_));
  XOR2X1   g10412(.A(new_n10668_), .B(new_n10611_), .Y(new_n10669_));
  XOR2X1   g10413(.A(new_n10669_), .B(new_n10607_), .Y(new_n10670_));
  XOR2X1   g10414(.A(new_n10670_), .B(new_n10603_), .Y(new_n10671_));
  XOR2X1   g10415(.A(new_n10671_), .B(new_n10601_), .Y(new_n10672_));
  XOR2X1   g10416(.A(new_n10672_), .B(new_n10597_), .Y(new_n10673_));
  AOI22X1  g10417(.A0(new_n3204_), .A1(\b[43] ), .B0(new_n3203_), .B1(\b[42] ), .Y(new_n10674_));
  OAI21X1  g10418(.A0(new_n3321_), .A1(new_n4015_), .B0(new_n10674_), .Y(new_n10675_));
  AOI21X1  g10419(.A0(new_n4014_), .A1(new_n3080_), .B0(new_n10675_), .Y(new_n10676_));
  XOR2X1   g10420(.A(new_n10676_), .B(\a[38] ), .Y(new_n10677_));
  XOR2X1   g10421(.A(new_n10677_), .B(new_n10673_), .Y(new_n10678_));
  NOR2X1   g10422(.A(new_n10505_), .B(new_n10501_), .Y(new_n10679_));
  AOI21X1  g10423(.A0(new_n10506_), .A1(new_n10420_), .B0(new_n10679_), .Y(new_n10680_));
  XOR2X1   g10424(.A(new_n10680_), .B(new_n10678_), .Y(new_n10681_));
  AOI22X1  g10425(.A0(new_n2813_), .A1(\b[46] ), .B0(new_n2812_), .B1(\b[45] ), .Y(new_n10682_));
  OAI21X1  g10426(.A0(new_n2946_), .A1(new_n4336_), .B0(new_n10682_), .Y(new_n10683_));
  AOI21X1  g10427(.A0(new_n4509_), .A1(new_n2652_), .B0(new_n10683_), .Y(new_n10684_));
  XOR2X1   g10428(.A(new_n10684_), .B(\a[35] ), .Y(new_n10685_));
  XOR2X1   g10429(.A(new_n10685_), .B(new_n10681_), .Y(new_n10686_));
  XOR2X1   g10430(.A(new_n10686_), .B(new_n10592_), .Y(new_n10687_));
  XOR2X1   g10431(.A(new_n10687_), .B(new_n10583_), .Y(new_n10688_));
  XOR2X1   g10432(.A(new_n10688_), .B(new_n10574_), .Y(new_n10689_));
  XOR2X1   g10433(.A(new_n10689_), .B(new_n10566_), .Y(new_n10690_));
  XOR2X1   g10434(.A(new_n10690_), .B(new_n10558_), .Y(new_n10691_));
  XOR2X1   g10435(.A(new_n10691_), .B(new_n10547_), .Y(new_n10692_));
  INVX1    g10436(.A(new_n10692_), .Y(new_n10693_));
  NOR2X1   g10437(.A(new_n10382_), .B(new_n10378_), .Y(new_n10694_));
  AOI21X1  g10438(.A0(new_n10531_), .A1(new_n10383_), .B0(new_n10694_), .Y(new_n10695_));
  XOR2X1   g10439(.A(new_n10695_), .B(new_n10693_), .Y(new_n10696_));
  INVX1    g10440(.A(new_n10532_), .Y(new_n10697_));
  NOR2X1   g10441(.A(new_n10534_), .B(new_n10697_), .Y(new_n10698_));
  AOI21X1  g10442(.A0(new_n10538_), .A1(new_n10537_), .B0(new_n10535_), .Y(new_n10699_));
  OR2X1    g10443(.A(new_n10699_), .B(new_n10698_), .Y(new_n10700_));
  XOR2X1   g10444(.A(new_n10700_), .B(new_n10696_), .Y(\f[79] ));
  NOR2X1   g10445(.A(new_n10695_), .B(new_n10693_), .Y(new_n10702_));
  INVX1    g10446(.A(new_n10702_), .Y(new_n10703_));
  OAI21X1  g10447(.A0(new_n10699_), .A1(new_n10698_), .B0(new_n10696_), .Y(new_n10704_));
  AND2X1   g10448(.A(new_n10704_), .B(new_n10703_), .Y(new_n10705_));
  NOR2X1   g10449(.A(new_n10546_), .B(new_n10543_), .Y(new_n10706_));
  AOI21X1  g10450(.A0(new_n10691_), .A1(new_n10547_), .B0(new_n10706_), .Y(new_n10707_));
  OR2X1    g10451(.A(new_n10557_), .B(new_n10551_), .Y(new_n10708_));
  OR2X1    g10452(.A(new_n10690_), .B(new_n10558_), .Y(new_n10709_));
  AND2X1   g10453(.A(new_n10709_), .B(new_n10708_), .Y(new_n10710_));
  AOI22X1  g10454(.A0(new_n7774_), .A1(new_n882_), .B0(new_n8600_), .B1(\b[63] ), .Y(new_n10711_));
  XOR2X1   g10455(.A(new_n10711_), .B(\a[17] ), .Y(new_n10712_));
  XOR2X1   g10456(.A(new_n10712_), .B(new_n10710_), .Y(new_n10713_));
  AOI22X1  g10457(.A0(new_n1263_), .A1(\b[62] ), .B0(new_n1262_), .B1(\b[61] ), .Y(new_n10714_));
  OAI21X1  g10458(.A0(new_n1261_), .A1(new_n7559_), .B0(new_n10714_), .Y(new_n10715_));
  AOI21X1  g10459(.A0(new_n7558_), .A1(new_n1075_), .B0(new_n10715_), .Y(new_n10716_));
  XOR2X1   g10460(.A(new_n10716_), .B(\a[20] ), .Y(new_n10717_));
  INVX1    g10461(.A(new_n10717_), .Y(new_n10718_));
  NOR2X1   g10462(.A(new_n10564_), .B(new_n10560_), .Y(new_n10719_));
  AOI21X1  g10463(.A0(new_n10689_), .A1(new_n10565_), .B0(new_n10719_), .Y(new_n10720_));
  XOR2X1   g10464(.A(new_n10720_), .B(new_n10718_), .Y(new_n10721_));
  AOI22X1  g10465(.A0(new_n1526_), .A1(\b[59] ), .B0(new_n1525_), .B1(\b[58] ), .Y(new_n10722_));
  OAI21X1  g10466(.A0(new_n1524_), .A1(new_n6933_), .B0(new_n10722_), .Y(new_n10723_));
  AOI21X1  g10467(.A0(new_n6932_), .A1(new_n1347_), .B0(new_n10723_), .Y(new_n10724_));
  XOR2X1   g10468(.A(new_n10724_), .B(\a[23] ), .Y(new_n10725_));
  OR2X1    g10469(.A(new_n10573_), .B(new_n10570_), .Y(new_n10726_));
  OR2X1    g10470(.A(new_n10688_), .B(new_n10574_), .Y(new_n10727_));
  AND2X1   g10471(.A(new_n10727_), .B(new_n10726_), .Y(new_n10728_));
  XOR2X1   g10472(.A(new_n10728_), .B(new_n10725_), .Y(new_n10729_));
  INVX1    g10473(.A(new_n10729_), .Y(new_n10730_));
  AOI22X1  g10474(.A0(new_n1814_), .A1(\b[56] ), .B0(new_n1813_), .B1(\b[55] ), .Y(new_n10731_));
  OAI21X1  g10475(.A0(new_n1812_), .A1(new_n6148_), .B0(new_n10731_), .Y(new_n10732_));
  AOI21X1  g10476(.A0(new_n6342_), .A1(new_n1617_), .B0(new_n10732_), .Y(new_n10733_));
  XOR2X1   g10477(.A(new_n10733_), .B(\a[26] ), .Y(new_n10734_));
  INVX1    g10478(.A(new_n10734_), .Y(new_n10735_));
  NOR2X1   g10479(.A(new_n10581_), .B(new_n10578_), .Y(new_n10736_));
  AOI21X1  g10480(.A0(new_n10687_), .A1(new_n10582_), .B0(new_n10736_), .Y(new_n10737_));
  XOR2X1   g10481(.A(new_n10737_), .B(new_n10735_), .Y(new_n10738_));
  AOI22X1  g10482(.A0(new_n2163_), .A1(\b[53] ), .B0(new_n2162_), .B1(\b[52] ), .Y(new_n10739_));
  OAI21X1  g10483(.A0(new_n2161_), .A1(new_n5787_), .B0(new_n10739_), .Y(new_n10740_));
  AOI21X1  g10484(.A0(new_n5786_), .A1(new_n1907_), .B0(new_n10740_), .Y(new_n10741_));
  XOR2X1   g10485(.A(new_n10741_), .B(\a[29] ), .Y(new_n10742_));
  OR2X1    g10486(.A(new_n10591_), .B(new_n10587_), .Y(new_n10743_));
  OR2X1    g10487(.A(new_n10686_), .B(new_n10592_), .Y(new_n10744_));
  AND2X1   g10488(.A(new_n10744_), .B(new_n10743_), .Y(new_n10745_));
  XOR2X1   g10489(.A(new_n10745_), .B(new_n10742_), .Y(new_n10746_));
  INVX1    g10490(.A(new_n10746_), .Y(new_n10747_));
  AOI22X1  g10491(.A0(new_n2545_), .A1(\b[50] ), .B0(new_n2544_), .B1(\b[49] ), .Y(new_n10748_));
  OAI21X1  g10492(.A0(new_n2543_), .A1(new_n5036_), .B0(new_n10748_), .Y(new_n10749_));
  AOI21X1  g10493(.A0(new_n5204_), .A1(new_n2260_), .B0(new_n10749_), .Y(new_n10750_));
  XOR2X1   g10494(.A(new_n10750_), .B(\a[32] ), .Y(new_n10751_));
  INVX1    g10495(.A(new_n10751_), .Y(new_n10752_));
  NOR2X1   g10496(.A(new_n10680_), .B(new_n10678_), .Y(new_n10753_));
  INVX1    g10497(.A(new_n10685_), .Y(new_n10754_));
  AOI21X1  g10498(.A0(new_n10754_), .A1(new_n10681_), .B0(new_n10753_), .Y(new_n10755_));
  XOR2X1   g10499(.A(new_n10755_), .B(new_n10752_), .Y(new_n10756_));
  AND2X1   g10500(.A(new_n10672_), .B(new_n10597_), .Y(new_n10757_));
  INVX1    g10501(.A(new_n10757_), .Y(new_n10758_));
  INVX1    g10502(.A(new_n10673_), .Y(new_n10759_));
  OAI21X1  g10503(.A0(new_n10677_), .A1(new_n10759_), .B0(new_n10758_), .Y(new_n10760_));
  AOI22X1  g10504(.A0(new_n3204_), .A1(\b[44] ), .B0(new_n3203_), .B1(\b[43] ), .Y(new_n10761_));
  OAI21X1  g10505(.A0(new_n3321_), .A1(new_n4012_), .B0(new_n10761_), .Y(new_n10762_));
  AOI21X1  g10506(.A0(new_n4178_), .A1(new_n3080_), .B0(new_n10762_), .Y(new_n10763_));
  XOR2X1   g10507(.A(new_n10763_), .B(new_n3078_), .Y(new_n10764_));
  INVX1    g10508(.A(new_n10603_), .Y(new_n10765_));
  NAND2X1  g10509(.A(new_n10670_), .B(new_n10765_), .Y(new_n10766_));
  OAI21X1  g10510(.A0(new_n10671_), .A1(new_n10601_), .B0(new_n10766_), .Y(new_n10767_));
  AOI22X1  g10511(.A0(new_n3652_), .A1(\b[41] ), .B0(new_n3651_), .B1(\b[40] ), .Y(new_n10768_));
  OAI21X1  g10512(.A0(new_n3778_), .A1(new_n3723_), .B0(new_n10768_), .Y(new_n10769_));
  AOI21X1  g10513(.A0(new_n3722_), .A1(new_n3480_), .B0(new_n10769_), .Y(new_n10770_));
  XOR2X1   g10514(.A(new_n10770_), .B(new_n3478_), .Y(new_n10771_));
  OAI21X1  g10515(.A0(new_n10610_), .A1(new_n10609_), .B0(new_n10668_), .Y(new_n10772_));
  OR2X1    g10516(.A(new_n10669_), .B(new_n10607_), .Y(new_n10773_));
  AND2X1   g10517(.A(new_n10773_), .B(new_n10772_), .Y(new_n10774_));
  NOR2X1   g10518(.A(new_n10635_), .B(new_n10632_), .Y(new_n10775_));
  INVX1    g10519(.A(new_n10775_), .Y(new_n10776_));
  INVX1    g10520(.A(new_n10636_), .Y(new_n10777_));
  OAI21X1  g10521(.A0(new_n10640_), .A1(new_n10777_), .B0(new_n10776_), .Y(new_n10778_));
  AOI22X1  g10522(.A0(new_n6438_), .A1(\b[26] ), .B0(new_n6437_), .B1(\b[25] ), .Y(new_n10779_));
  OAI21X1  g10523(.A0(new_n6436_), .A1(new_n1588_), .B0(new_n10779_), .Y(new_n10780_));
  AOI21X1  g10524(.A0(new_n6023_), .A1(new_n1783_), .B0(new_n10780_), .Y(new_n10781_));
  XOR2X1   g10525(.A(new_n10781_), .B(new_n6019_), .Y(new_n10782_));
  OR2X1    g10526(.A(new_n10626_), .B(new_n10613_), .Y(new_n10783_));
  AND2X1   g10527(.A(new_n10626_), .B(new_n10613_), .Y(new_n10784_));
  OAI21X1  g10528(.A0(new_n10631_), .A1(new_n10784_), .B0(new_n10783_), .Y(new_n10785_));
  AOI22X1  g10529(.A0(new_n7192_), .A1(\b[20] ), .B0(new_n7189_), .B1(\b[19] ), .Y(new_n10786_));
  OAI21X1  g10530(.A0(new_n7627_), .A1(new_n1115_), .B0(new_n10786_), .Y(new_n10787_));
  AOI21X1  g10531(.A0(new_n7187_), .A1(new_n1217_), .B0(new_n10787_), .Y(new_n10788_));
  XOR2X1   g10532(.A(new_n10788_), .B(\a[62] ), .Y(new_n10789_));
  AOI22X1  g10533(.A0(new_n7818_), .A1(\b[16] ), .B0(new_n7817_), .B1(\b[17] ), .Y(new_n10790_));
  NOR2X1   g10534(.A(new_n10790_), .B(new_n10615_), .Y(new_n10791_));
  XOR2X1   g10535(.A(new_n10790_), .B(new_n10615_), .Y(new_n10792_));
  INVX1    g10536(.A(new_n10792_), .Y(new_n10793_));
  NOR2X1   g10537(.A(new_n10793_), .B(new_n10789_), .Y(new_n10794_));
  AOI21X1  g10538(.A0(new_n10790_), .A1(new_n10615_), .B0(new_n10794_), .Y(new_n10795_));
  INVX1    g10539(.A(new_n10795_), .Y(new_n10796_));
  OAI22X1  g10540(.A0(new_n10796_), .A1(new_n10791_), .B0(new_n10792_), .B1(new_n10789_), .Y(new_n10797_));
  NOR2X1   g10541(.A(new_n10618_), .B(new_n10615_), .Y(new_n10798_));
  XOR2X1   g10542(.A(new_n10623_), .B(new_n7185_), .Y(new_n10799_));
  AOI21X1  g10543(.A0(new_n10799_), .A1(new_n10619_), .B0(new_n10798_), .Y(new_n10800_));
  XOR2X1   g10544(.A(new_n10800_), .B(new_n10797_), .Y(new_n10801_));
  AOI22X1  g10545(.A0(new_n6603_), .A1(\b[23] ), .B0(new_n6600_), .B1(\b[22] ), .Y(new_n10802_));
  OAI21X1  g10546(.A0(new_n6804_), .A1(new_n1482_), .B0(new_n10802_), .Y(new_n10803_));
  AOI21X1  g10547(.A0(new_n6598_), .A1(new_n1481_), .B0(new_n10803_), .Y(new_n10804_));
  XOR2X1   g10548(.A(new_n10804_), .B(\a[59] ), .Y(new_n10805_));
  XOR2X1   g10549(.A(new_n10805_), .B(new_n10801_), .Y(new_n10806_));
  XOR2X1   g10550(.A(new_n10806_), .B(new_n10785_), .Y(new_n10807_));
  XOR2X1   g10551(.A(new_n10807_), .B(new_n10782_), .Y(new_n10808_));
  XOR2X1   g10552(.A(new_n10808_), .B(new_n10778_), .Y(new_n10809_));
  AOI22X1  g10553(.A0(new_n5430_), .A1(\b[29] ), .B0(new_n5427_), .B1(\b[28] ), .Y(new_n10810_));
  OAI21X1  g10554(.A0(new_n5891_), .A1(new_n2126_), .B0(new_n10810_), .Y(new_n10811_));
  AOI21X1  g10555(.A0(new_n5425_), .A1(new_n2125_), .B0(new_n10811_), .Y(new_n10812_));
  XOR2X1   g10556(.A(new_n10812_), .B(\a[53] ), .Y(new_n10813_));
  XOR2X1   g10557(.A(new_n10813_), .B(new_n10809_), .Y(new_n10814_));
  NOR2X1   g10558(.A(new_n10647_), .B(new_n10643_), .Y(new_n10815_));
  AOI21X1  g10559(.A0(new_n10642_), .A1(new_n10465_), .B0(new_n10815_), .Y(new_n10816_));
  XOR2X1   g10560(.A(new_n10816_), .B(new_n10814_), .Y(new_n10817_));
  AOI22X1  g10561(.A0(new_n4880_), .A1(\b[32] ), .B0(new_n4877_), .B1(\b[31] ), .Y(new_n10818_));
  OAI21X1  g10562(.A0(new_n5291_), .A1(new_n2356_), .B0(new_n10818_), .Y(new_n10819_));
  AOI21X1  g10563(.A0(new_n4875_), .A1(new_n2495_), .B0(new_n10819_), .Y(new_n10820_));
  XOR2X1   g10564(.A(new_n10820_), .B(\a[50] ), .Y(new_n10821_));
  XOR2X1   g10565(.A(new_n10821_), .B(new_n10817_), .Y(new_n10822_));
  NOR2X1   g10566(.A(new_n10652_), .B(new_n10649_), .Y(new_n10823_));
  INVX1    g10567(.A(new_n10657_), .Y(new_n10824_));
  AOI21X1  g10568(.A0(new_n10824_), .A1(new_n10653_), .B0(new_n10823_), .Y(new_n10825_));
  XOR2X1   g10569(.A(new_n10825_), .B(new_n10822_), .Y(new_n10826_));
  AOI22X1  g10570(.A0(new_n4572_), .A1(\b[35] ), .B0(new_n4571_), .B1(\b[34] ), .Y(new_n10827_));
  OAI21X1  g10571(.A0(new_n4740_), .A1(new_n2893_), .B0(new_n10827_), .Y(new_n10828_));
  AOI21X1  g10572(.A0(new_n4375_), .A1(new_n2892_), .B0(new_n10828_), .Y(new_n10829_));
  XOR2X1   g10573(.A(new_n10829_), .B(\a[47] ), .Y(new_n10830_));
  XOR2X1   g10574(.A(new_n10830_), .B(new_n10826_), .Y(new_n10831_));
  OR2X1    g10575(.A(new_n10662_), .B(new_n10658_), .Y(new_n10832_));
  OR2X1    g10576(.A(new_n10667_), .B(new_n10663_), .Y(new_n10833_));
  AND2X1   g10577(.A(new_n10833_), .B(new_n10832_), .Y(new_n10834_));
  XOR2X1   g10578(.A(new_n10834_), .B(new_n10831_), .Y(new_n10835_));
  AOI22X1  g10579(.A0(new_n4095_), .A1(\b[38] ), .B0(new_n4094_), .B1(\b[37] ), .Y(new_n10836_));
  OAI21X1  g10580(.A0(new_n4233_), .A1(new_n3276_), .B0(new_n10836_), .Y(new_n10837_));
  AOI21X1  g10581(.A0(new_n3901_), .A1(new_n3275_), .B0(new_n10837_), .Y(new_n10838_));
  XOR2X1   g10582(.A(new_n10838_), .B(\a[44] ), .Y(new_n10839_));
  XOR2X1   g10583(.A(new_n10839_), .B(new_n10835_), .Y(new_n10840_));
  XOR2X1   g10584(.A(new_n10840_), .B(new_n10774_), .Y(new_n10841_));
  XOR2X1   g10585(.A(new_n10841_), .B(new_n10771_), .Y(new_n10842_));
  XOR2X1   g10586(.A(new_n10842_), .B(new_n10767_), .Y(new_n10843_));
  XOR2X1   g10587(.A(new_n10843_), .B(new_n10764_), .Y(new_n10844_));
  XOR2X1   g10588(.A(new_n10844_), .B(new_n10760_), .Y(new_n10845_));
  AOI22X1  g10589(.A0(new_n2813_), .A1(\b[47] ), .B0(new_n2812_), .B1(\b[46] ), .Y(new_n10846_));
  OAI21X1  g10590(.A0(new_n2946_), .A1(new_n4674_), .B0(new_n10846_), .Y(new_n10847_));
  AOI21X1  g10591(.A0(new_n4673_), .A1(new_n2652_), .B0(new_n10847_), .Y(new_n10848_));
  XOR2X1   g10592(.A(new_n10848_), .B(\a[35] ), .Y(new_n10849_));
  XOR2X1   g10593(.A(new_n10849_), .B(new_n10845_), .Y(new_n10850_));
  XOR2X1   g10594(.A(new_n10850_), .B(new_n10756_), .Y(new_n10851_));
  XOR2X1   g10595(.A(new_n10851_), .B(new_n10747_), .Y(new_n10852_));
  XOR2X1   g10596(.A(new_n10852_), .B(new_n10738_), .Y(new_n10853_));
  XOR2X1   g10597(.A(new_n10853_), .B(new_n10730_), .Y(new_n10854_));
  XOR2X1   g10598(.A(new_n10854_), .B(new_n10721_), .Y(new_n10855_));
  XOR2X1   g10599(.A(new_n10855_), .B(new_n10713_), .Y(new_n10856_));
  XOR2X1   g10600(.A(new_n10856_), .B(new_n10707_), .Y(new_n10857_));
  XOR2X1   g10601(.A(new_n10857_), .B(new_n10705_), .Y(\f[80] ));
  INVX1    g10602(.A(new_n10707_), .Y(new_n10859_));
  AND2X1   g10603(.A(new_n10856_), .B(new_n10859_), .Y(new_n10860_));
  AOI21X1  g10604(.A0(new_n10704_), .A1(new_n10703_), .B0(new_n10857_), .Y(new_n10861_));
  OR2X1    g10605(.A(new_n10861_), .B(new_n10860_), .Y(new_n10862_));
  AOI21X1  g10606(.A0(new_n10709_), .A1(new_n10708_), .B0(new_n10712_), .Y(new_n10863_));
  AOI21X1  g10607(.A0(new_n10855_), .A1(new_n10713_), .B0(new_n10863_), .Y(new_n10864_));
  NOR2X1   g10608(.A(new_n10720_), .B(new_n10717_), .Y(new_n10865_));
  INVX1    g10609(.A(new_n10865_), .Y(new_n10866_));
  OAI21X1  g10610(.A0(new_n10854_), .A1(new_n10721_), .B0(new_n10866_), .Y(new_n10867_));
  AOI22X1  g10611(.A0(new_n1263_), .A1(\b[63] ), .B0(new_n1262_), .B1(\b[62] ), .Y(new_n10868_));
  OAI21X1  g10612(.A0(new_n1261_), .A1(new_n7748_), .B0(new_n10868_), .Y(new_n10869_));
  AOI21X1  g10613(.A0(new_n7747_), .A1(new_n1075_), .B0(new_n10869_), .Y(new_n10870_));
  XOR2X1   g10614(.A(new_n10870_), .B(\a[20] ), .Y(new_n10871_));
  XOR2X1   g10615(.A(new_n10871_), .B(new_n10867_), .Y(new_n10872_));
  AOI22X1  g10616(.A0(new_n1526_), .A1(\b[60] ), .B0(new_n1525_), .B1(\b[59] ), .Y(new_n10873_));
  OAI21X1  g10617(.A0(new_n1524_), .A1(new_n6930_), .B0(new_n10873_), .Y(new_n10874_));
  AOI21X1  g10618(.A0(new_n6951_), .A1(new_n1347_), .B0(new_n10874_), .Y(new_n10875_));
  XOR2X1   g10619(.A(new_n10875_), .B(\a[23] ), .Y(new_n10876_));
  AOI21X1  g10620(.A0(new_n10727_), .A1(new_n10726_), .B0(new_n10725_), .Y(new_n10877_));
  AOI21X1  g10621(.A0(new_n10853_), .A1(new_n10729_), .B0(new_n10877_), .Y(new_n10878_));
  XOR2X1   g10622(.A(new_n10878_), .B(new_n10876_), .Y(new_n10879_));
  AOI22X1  g10623(.A0(new_n2163_), .A1(\b[54] ), .B0(new_n2162_), .B1(\b[53] ), .Y(new_n10880_));
  OAI21X1  g10624(.A0(new_n2161_), .A1(new_n5808_), .B0(new_n10880_), .Y(new_n10881_));
  AOI21X1  g10625(.A0(new_n5807_), .A1(new_n1907_), .B0(new_n10881_), .Y(new_n10882_));
  XOR2X1   g10626(.A(new_n10882_), .B(\a[29] ), .Y(new_n10883_));
  NOR2X1   g10627(.A(new_n10745_), .B(new_n10742_), .Y(new_n10884_));
  AOI21X1  g10628(.A0(new_n10851_), .A1(new_n10746_), .B0(new_n10884_), .Y(new_n10885_));
  XOR2X1   g10629(.A(new_n10885_), .B(new_n10883_), .Y(new_n10886_));
  NOR2X1   g10630(.A(new_n10840_), .B(new_n10774_), .Y(new_n10887_));
  AOI21X1  g10631(.A0(new_n10841_), .A1(new_n10771_), .B0(new_n10887_), .Y(new_n10888_));
  INVX1    g10632(.A(new_n10888_), .Y(new_n10889_));
  AOI21X1  g10633(.A0(new_n10833_), .A1(new_n10832_), .B0(new_n10831_), .Y(new_n10890_));
  INVX1    g10634(.A(new_n10839_), .Y(new_n10891_));
  AOI21X1  g10635(.A0(new_n10891_), .A1(new_n10835_), .B0(new_n10890_), .Y(new_n10892_));
  INVX1    g10636(.A(new_n10892_), .Y(new_n10893_));
  NOR2X1   g10637(.A(new_n10825_), .B(new_n10822_), .Y(new_n10894_));
  INVX1    g10638(.A(new_n10894_), .Y(new_n10895_));
  INVX1    g10639(.A(new_n10826_), .Y(new_n10896_));
  OAI21X1  g10640(.A0(new_n10830_), .A1(new_n10896_), .B0(new_n10895_), .Y(new_n10897_));
  INVX1    g10641(.A(new_n10797_), .Y(new_n10898_));
  NOR2X1   g10642(.A(new_n10800_), .B(new_n10898_), .Y(new_n10899_));
  NOR2X1   g10643(.A(new_n10805_), .B(new_n10801_), .Y(new_n10900_));
  NOR2X1   g10644(.A(new_n10900_), .B(new_n10899_), .Y(new_n10901_));
  INVX1    g10645(.A(new_n10901_), .Y(new_n10902_));
  AOI22X1  g10646(.A0(new_n7192_), .A1(\b[21] ), .B0(new_n7189_), .B1(\b[20] ), .Y(new_n10903_));
  OAI21X1  g10647(.A0(new_n7627_), .A1(new_n1300_), .B0(new_n10903_), .Y(new_n10904_));
  AOI21X1  g10648(.A0(new_n7187_), .A1(new_n1299_), .B0(new_n10904_), .Y(new_n10905_));
  XOR2X1   g10649(.A(new_n10905_), .B(\a[62] ), .Y(new_n10906_));
  INVX1    g10650(.A(new_n10790_), .Y(new_n10907_));
  AOI22X1  g10651(.A0(new_n7818_), .A1(\b[17] ), .B0(new_n7817_), .B1(\b[18] ), .Y(new_n10908_));
  XOR2X1   g10652(.A(new_n10908_), .B(\a[17] ), .Y(new_n10909_));
  XOR2X1   g10653(.A(new_n10909_), .B(new_n10907_), .Y(new_n10910_));
  XOR2X1   g10654(.A(new_n10910_), .B(new_n10906_), .Y(new_n10911_));
  XOR2X1   g10655(.A(new_n10911_), .B(new_n10796_), .Y(new_n10912_));
  AOI22X1  g10656(.A0(new_n6603_), .A1(\b[24] ), .B0(new_n6600_), .B1(\b[23] ), .Y(new_n10913_));
  OAI21X1  g10657(.A0(new_n6804_), .A1(new_n1479_), .B0(new_n10913_), .Y(new_n10914_));
  AOI21X1  g10658(.A0(new_n6598_), .A1(new_n1572_), .B0(new_n10914_), .Y(new_n10915_));
  XOR2X1   g10659(.A(new_n10915_), .B(\a[59] ), .Y(new_n10916_));
  XOR2X1   g10660(.A(new_n10916_), .B(new_n10912_), .Y(new_n10917_));
  XOR2X1   g10661(.A(new_n10917_), .B(new_n10902_), .Y(new_n10918_));
  AOI22X1  g10662(.A0(new_n6438_), .A1(\b[27] ), .B0(new_n6437_), .B1(\b[26] ), .Y(new_n10919_));
  OAI21X1  g10663(.A0(new_n6436_), .A1(new_n1880_), .B0(new_n10919_), .Y(new_n10920_));
  AOI21X1  g10664(.A0(new_n6023_), .A1(new_n1879_), .B0(new_n10920_), .Y(new_n10921_));
  XOR2X1   g10665(.A(new_n10921_), .B(\a[56] ), .Y(new_n10922_));
  XOR2X1   g10666(.A(new_n10922_), .B(new_n10918_), .Y(new_n10923_));
  AND2X1   g10667(.A(new_n10806_), .B(new_n10785_), .Y(new_n10924_));
  AOI21X1  g10668(.A0(new_n10807_), .A1(new_n10782_), .B0(new_n10924_), .Y(new_n10925_));
  XOR2X1   g10669(.A(new_n10925_), .B(new_n10923_), .Y(new_n10926_));
  AOI22X1  g10670(.A0(new_n5430_), .A1(\b[30] ), .B0(new_n5427_), .B1(\b[29] ), .Y(new_n10927_));
  OAI21X1  g10671(.A0(new_n5891_), .A1(new_n2231_), .B0(new_n10927_), .Y(new_n10928_));
  AOI21X1  g10672(.A0(new_n5425_), .A1(new_n2230_), .B0(new_n10928_), .Y(new_n10929_));
  XOR2X1   g10673(.A(new_n10929_), .B(\a[53] ), .Y(new_n10930_));
  XOR2X1   g10674(.A(new_n10930_), .B(new_n10926_), .Y(new_n10931_));
  AND2X1   g10675(.A(new_n10808_), .B(new_n10778_), .Y(new_n10932_));
  INVX1    g10676(.A(new_n10813_), .Y(new_n10933_));
  AOI21X1  g10677(.A0(new_n10933_), .A1(new_n10809_), .B0(new_n10932_), .Y(new_n10934_));
  XOR2X1   g10678(.A(new_n10934_), .B(new_n10931_), .Y(new_n10935_));
  INVX1    g10679(.A(new_n10935_), .Y(new_n10936_));
  AOI22X1  g10680(.A0(new_n4880_), .A1(\b[33] ), .B0(new_n4877_), .B1(\b[32] ), .Y(new_n10937_));
  OAI21X1  g10681(.A0(new_n5291_), .A1(new_n2615_), .B0(new_n10937_), .Y(new_n10938_));
  AOI21X1  g10682(.A0(new_n4875_), .A1(new_n2614_), .B0(new_n10938_), .Y(new_n10939_));
  XOR2X1   g10683(.A(new_n10939_), .B(\a[50] ), .Y(new_n10940_));
  NOR2X1   g10684(.A(new_n10816_), .B(new_n10814_), .Y(new_n10941_));
  INVX1    g10685(.A(new_n10821_), .Y(new_n10942_));
  AOI21X1  g10686(.A0(new_n10942_), .A1(new_n10817_), .B0(new_n10941_), .Y(new_n10943_));
  XOR2X1   g10687(.A(new_n10943_), .B(new_n10940_), .Y(new_n10944_));
  XOR2X1   g10688(.A(new_n10944_), .B(new_n10936_), .Y(new_n10945_));
  AOI22X1  g10689(.A0(new_n4572_), .A1(\b[36] ), .B0(new_n4571_), .B1(\b[35] ), .Y(new_n10946_));
  OAI21X1  g10690(.A0(new_n4740_), .A1(new_n2890_), .B0(new_n10946_), .Y(new_n10947_));
  AOI21X1  g10691(.A0(new_n4375_), .A1(new_n3015_), .B0(new_n10947_), .Y(new_n10948_));
  XOR2X1   g10692(.A(new_n10948_), .B(\a[47] ), .Y(new_n10949_));
  XOR2X1   g10693(.A(new_n10949_), .B(new_n10945_), .Y(new_n10950_));
  XOR2X1   g10694(.A(new_n10950_), .B(new_n10897_), .Y(new_n10951_));
  AOI22X1  g10695(.A0(new_n4095_), .A1(\b[39] ), .B0(new_n4094_), .B1(\b[38] ), .Y(new_n10952_));
  OAI21X1  g10696(.A0(new_n4233_), .A1(new_n3413_), .B0(new_n10952_), .Y(new_n10953_));
  AOI21X1  g10697(.A0(new_n3901_), .A1(new_n3412_), .B0(new_n10953_), .Y(new_n10954_));
  XOR2X1   g10698(.A(new_n10954_), .B(\a[44] ), .Y(new_n10955_));
  XOR2X1   g10699(.A(new_n10955_), .B(new_n10951_), .Y(new_n10956_));
  XOR2X1   g10700(.A(new_n10956_), .B(new_n10893_), .Y(new_n10957_));
  AOI22X1  g10701(.A0(new_n3652_), .A1(\b[42] ), .B0(new_n3651_), .B1(\b[41] ), .Y(new_n10958_));
  OAI21X1  g10702(.A0(new_n3778_), .A1(new_n3720_), .B0(new_n10958_), .Y(new_n10959_));
  AOI21X1  g10703(.A0(new_n3860_), .A1(new_n3480_), .B0(new_n10959_), .Y(new_n10960_));
  XOR2X1   g10704(.A(new_n10960_), .B(\a[41] ), .Y(new_n10961_));
  XOR2X1   g10705(.A(new_n10961_), .B(new_n10957_), .Y(new_n10962_));
  XOR2X1   g10706(.A(new_n10962_), .B(new_n10889_), .Y(new_n10963_));
  AOI22X1  g10707(.A0(new_n3204_), .A1(\b[45] ), .B0(new_n3203_), .B1(\b[44] ), .Y(new_n10964_));
  OAI21X1  g10708(.A0(new_n3321_), .A1(new_n4339_), .B0(new_n10964_), .Y(new_n10965_));
  AOI21X1  g10709(.A0(new_n4338_), .A1(new_n3080_), .B0(new_n10965_), .Y(new_n10966_));
  XOR2X1   g10710(.A(new_n10966_), .B(\a[38] ), .Y(new_n10967_));
  XOR2X1   g10711(.A(new_n10967_), .B(new_n10963_), .Y(new_n10968_));
  AND2X1   g10712(.A(new_n10842_), .B(new_n10767_), .Y(new_n10969_));
  AOI21X1  g10713(.A0(new_n10843_), .A1(new_n10764_), .B0(new_n10969_), .Y(new_n10970_));
  XOR2X1   g10714(.A(new_n10970_), .B(new_n10968_), .Y(new_n10971_));
  AOI22X1  g10715(.A0(new_n2813_), .A1(\b[48] ), .B0(new_n2812_), .B1(\b[47] ), .Y(new_n10972_));
  OAI21X1  g10716(.A0(new_n2946_), .A1(new_n4693_), .B0(new_n10972_), .Y(new_n10973_));
  AOI21X1  g10717(.A0(new_n4692_), .A1(new_n2652_), .B0(new_n10973_), .Y(new_n10974_));
  XOR2X1   g10718(.A(new_n10974_), .B(\a[35] ), .Y(new_n10975_));
  XOR2X1   g10719(.A(new_n10975_), .B(new_n10971_), .Y(new_n10976_));
  AND2X1   g10720(.A(new_n10844_), .B(new_n10760_), .Y(new_n10977_));
  INVX1    g10721(.A(new_n10849_), .Y(new_n10978_));
  AOI21X1  g10722(.A0(new_n10978_), .A1(new_n10845_), .B0(new_n10977_), .Y(new_n10979_));
  XOR2X1   g10723(.A(new_n10979_), .B(new_n10976_), .Y(new_n10980_));
  AOI22X1  g10724(.A0(new_n2545_), .A1(\b[51] ), .B0(new_n2544_), .B1(\b[50] ), .Y(new_n10981_));
  OAI21X1  g10725(.A0(new_n2543_), .A1(new_n5237_), .B0(new_n10981_), .Y(new_n10982_));
  AOI21X1  g10726(.A0(new_n5236_), .A1(new_n2260_), .B0(new_n10982_), .Y(new_n10983_));
  XOR2X1   g10727(.A(new_n10983_), .B(\a[32] ), .Y(new_n10984_));
  OR2X1    g10728(.A(new_n10755_), .B(new_n10751_), .Y(new_n10985_));
  OR2X1    g10729(.A(new_n10850_), .B(new_n10756_), .Y(new_n10986_));
  AND2X1   g10730(.A(new_n10986_), .B(new_n10985_), .Y(new_n10987_));
  XOR2X1   g10731(.A(new_n10987_), .B(new_n10984_), .Y(new_n10988_));
  XOR2X1   g10732(.A(new_n10988_), .B(new_n10980_), .Y(new_n10989_));
  INVX1    g10733(.A(new_n10989_), .Y(new_n10990_));
  XOR2X1   g10734(.A(new_n10990_), .B(new_n10886_), .Y(new_n10991_));
  AOI22X1  g10735(.A0(new_n1814_), .A1(\b[57] ), .B0(new_n1813_), .B1(\b[56] ), .Y(new_n10992_));
  OAI21X1  g10736(.A0(new_n1812_), .A1(new_n6523_), .B0(new_n10992_), .Y(new_n10993_));
  AOI21X1  g10737(.A0(new_n6522_), .A1(new_n1617_), .B0(new_n10993_), .Y(new_n10994_));
  XOR2X1   g10738(.A(new_n10994_), .B(\a[26] ), .Y(new_n10995_));
  OR2X1    g10739(.A(new_n10737_), .B(new_n10734_), .Y(new_n10996_));
  OR2X1    g10740(.A(new_n10852_), .B(new_n10738_), .Y(new_n10997_));
  AND2X1   g10741(.A(new_n10997_), .B(new_n10996_), .Y(new_n10998_));
  XOR2X1   g10742(.A(new_n10998_), .B(new_n10995_), .Y(new_n10999_));
  XOR2X1   g10743(.A(new_n10999_), .B(new_n10991_), .Y(new_n11000_));
  XOR2X1   g10744(.A(new_n11000_), .B(new_n10879_), .Y(new_n11001_));
  INVX1    g10745(.A(new_n11001_), .Y(new_n11002_));
  XOR2X1   g10746(.A(new_n11002_), .B(new_n10872_), .Y(new_n11003_));
  XOR2X1   g10747(.A(new_n11003_), .B(new_n10864_), .Y(new_n11004_));
  XOR2X1   g10748(.A(new_n11004_), .B(new_n10862_), .Y(\f[81] ));
  OR2X1    g10749(.A(new_n11003_), .B(new_n10864_), .Y(new_n11006_));
  OAI21X1  g10750(.A0(new_n10861_), .A1(new_n10860_), .B0(new_n11004_), .Y(new_n11007_));
  AND2X1   g10751(.A(new_n11007_), .B(new_n11006_), .Y(new_n11008_));
  XOR2X1   g10752(.A(new_n10870_), .B(new_n1072_), .Y(new_n11009_));
  AND2X1   g10753(.A(new_n11009_), .B(new_n10867_), .Y(new_n11010_));
  NOR2X1   g10754(.A(new_n11001_), .B(new_n10872_), .Y(new_n11011_));
  NOR2X1   g10755(.A(new_n11011_), .B(new_n11010_), .Y(new_n11012_));
  NOR2X1   g10756(.A(new_n10878_), .B(new_n10876_), .Y(new_n11013_));
  INVX1    g10757(.A(new_n11013_), .Y(new_n11014_));
  INVX1    g10758(.A(new_n10879_), .Y(new_n11015_));
  OAI21X1  g10759(.A0(new_n11000_), .A1(new_n11015_), .B0(new_n11014_), .Y(new_n11016_));
  OAI22X1  g10760(.A0(new_n1261_), .A1(new_n7745_), .B0(new_n1078_), .B1(new_n7772_), .Y(new_n11017_));
  AOI21X1  g10761(.A0(new_n7775_), .A1(new_n1075_), .B0(new_n11017_), .Y(new_n11018_));
  XOR2X1   g10762(.A(new_n11018_), .B(\a[20] ), .Y(new_n11019_));
  OR2X1    g10763(.A(new_n11019_), .B(new_n11016_), .Y(new_n11020_));
  AOI22X1  g10764(.A0(new_n1526_), .A1(\b[61] ), .B0(new_n1525_), .B1(\b[60] ), .Y(new_n11021_));
  OAI21X1  g10765(.A0(new_n1524_), .A1(new_n7339_), .B0(new_n11021_), .Y(new_n11022_));
  AOI21X1  g10766(.A0(new_n7338_), .A1(new_n1347_), .B0(new_n11022_), .Y(new_n11023_));
  XOR2X1   g10767(.A(new_n11023_), .B(\a[23] ), .Y(new_n11024_));
  INVX1    g10768(.A(new_n10991_), .Y(new_n11025_));
  AOI21X1  g10769(.A0(new_n10997_), .A1(new_n10996_), .B0(new_n10995_), .Y(new_n11026_));
  AOI21X1  g10770(.A0(new_n10999_), .A1(new_n11025_), .B0(new_n11026_), .Y(new_n11027_));
  XOR2X1   g10771(.A(new_n11027_), .B(new_n11024_), .Y(new_n11028_));
  AOI22X1  g10772(.A0(new_n1814_), .A1(\b[58] ), .B0(new_n1813_), .B1(\b[57] ), .Y(new_n11029_));
  OAI21X1  g10773(.A0(new_n1812_), .A1(new_n6520_), .B0(new_n11029_), .Y(new_n11030_));
  AOI21X1  g10774(.A0(new_n6732_), .A1(new_n1617_), .B0(new_n11030_), .Y(new_n11031_));
  XOR2X1   g10775(.A(new_n11031_), .B(\a[26] ), .Y(new_n11032_));
  INVX1    g10776(.A(new_n11032_), .Y(new_n11033_));
  NOR2X1   g10777(.A(new_n10885_), .B(new_n10883_), .Y(new_n11034_));
  AOI21X1  g10778(.A0(new_n10989_), .A1(new_n10886_), .B0(new_n11034_), .Y(new_n11035_));
  XOR2X1   g10779(.A(new_n11035_), .B(new_n11033_), .Y(new_n11036_));
  AOI22X1  g10780(.A0(new_n2163_), .A1(\b[55] ), .B0(new_n2162_), .B1(\b[54] ), .Y(new_n11037_));
  OAI21X1  g10781(.A0(new_n2161_), .A1(new_n6151_), .B0(new_n11037_), .Y(new_n11038_));
  AOI21X1  g10782(.A0(new_n6150_), .A1(new_n1907_), .B0(new_n11038_), .Y(new_n11039_));
  XOR2X1   g10783(.A(new_n11039_), .B(\a[29] ), .Y(new_n11040_));
  AOI21X1  g10784(.A0(new_n10986_), .A1(new_n10985_), .B0(new_n10984_), .Y(new_n11041_));
  AOI21X1  g10785(.A0(new_n10988_), .A1(new_n10980_), .B0(new_n11041_), .Y(new_n11042_));
  XOR2X1   g10786(.A(new_n11042_), .B(new_n11040_), .Y(new_n11043_));
  INVX1    g10787(.A(new_n11043_), .Y(new_n11044_));
  AOI22X1  g10788(.A0(new_n2545_), .A1(\b[52] ), .B0(new_n2544_), .B1(\b[51] ), .Y(new_n11045_));
  OAI21X1  g10789(.A0(new_n2543_), .A1(new_n5234_), .B0(new_n11045_), .Y(new_n11046_));
  AOI21X1  g10790(.A0(new_n5590_), .A1(new_n2260_), .B0(new_n11046_), .Y(new_n11047_));
  XOR2X1   g10791(.A(new_n11047_), .B(\a[32] ), .Y(new_n11048_));
  INVX1    g10792(.A(new_n11048_), .Y(new_n11049_));
  INVX1    g10793(.A(new_n10975_), .Y(new_n11050_));
  NOR2X1   g10794(.A(new_n10979_), .B(new_n10976_), .Y(new_n11051_));
  AOI21X1  g10795(.A0(new_n11050_), .A1(new_n10971_), .B0(new_n11051_), .Y(new_n11052_));
  XOR2X1   g10796(.A(new_n11052_), .B(new_n11049_), .Y(new_n11053_));
  XOR2X1   g10797(.A(new_n10954_), .B(new_n3899_), .Y(new_n11054_));
  NOR2X1   g10798(.A(new_n10956_), .B(new_n10892_), .Y(new_n11055_));
  AOI21X1  g10799(.A0(new_n11054_), .A1(new_n10951_), .B0(new_n11055_), .Y(new_n11056_));
  INVX1    g10800(.A(new_n11056_), .Y(new_n11057_));
  AOI22X1  g10801(.A0(new_n4095_), .A1(\b[40] ), .B0(new_n4094_), .B1(\b[39] ), .Y(new_n11058_));
  OAI21X1  g10802(.A0(new_n4233_), .A1(new_n3575_), .B0(new_n11058_), .Y(new_n11059_));
  AOI21X1  g10803(.A0(new_n3901_), .A1(new_n3574_), .B0(new_n11059_), .Y(new_n11060_));
  XOR2X1   g10804(.A(new_n11060_), .B(\a[44] ), .Y(new_n11061_));
  NOR2X1   g10805(.A(new_n10949_), .B(new_n10945_), .Y(new_n11062_));
  AOI21X1  g10806(.A0(new_n10950_), .A1(new_n10897_), .B0(new_n11062_), .Y(new_n11063_));
  NOR2X1   g10807(.A(new_n10916_), .B(new_n10912_), .Y(new_n11064_));
  AOI21X1  g10808(.A0(new_n10917_), .A1(new_n10902_), .B0(new_n11064_), .Y(new_n11065_));
  AOI22X1  g10809(.A0(new_n7818_), .A1(\b[18] ), .B0(new_n7817_), .B1(\b[19] ), .Y(new_n11066_));
  INVX1    g10810(.A(new_n11066_), .Y(new_n11067_));
  NOR2X1   g10811(.A(new_n10908_), .B(\a[17] ), .Y(new_n11068_));
  AOI21X1  g10812(.A0(new_n10909_), .A1(new_n10907_), .B0(new_n11068_), .Y(new_n11069_));
  XOR2X1   g10813(.A(new_n11069_), .B(new_n11067_), .Y(new_n11070_));
  INVX1    g10814(.A(new_n11070_), .Y(new_n11071_));
  AOI22X1  g10815(.A0(new_n7192_), .A1(\b[22] ), .B0(new_n7189_), .B1(\b[21] ), .Y(new_n11072_));
  OAI21X1  g10816(.A0(new_n7627_), .A1(new_n1297_), .B0(new_n11072_), .Y(new_n11073_));
  AOI21X1  g10817(.A0(new_n7187_), .A1(new_n1399_), .B0(new_n11073_), .Y(new_n11074_));
  XOR2X1   g10818(.A(new_n11074_), .B(\a[62] ), .Y(new_n11075_));
  XOR2X1   g10819(.A(new_n11075_), .B(new_n11071_), .Y(new_n11076_));
  INVX1    g10820(.A(new_n11076_), .Y(new_n11077_));
  INVX1    g10821(.A(new_n10906_), .Y(new_n11078_));
  NOR2X1   g10822(.A(new_n10911_), .B(new_n10795_), .Y(new_n11079_));
  AOI21X1  g10823(.A0(new_n10910_), .A1(new_n11078_), .B0(new_n11079_), .Y(new_n11080_));
  XOR2X1   g10824(.A(new_n11080_), .B(new_n11077_), .Y(new_n11081_));
  AOI22X1  g10825(.A0(new_n6603_), .A1(\b[25] ), .B0(new_n6600_), .B1(\b[24] ), .Y(new_n11082_));
  OAI21X1  g10826(.A0(new_n6804_), .A1(new_n1591_), .B0(new_n11082_), .Y(new_n11083_));
  AOI21X1  g10827(.A0(new_n6598_), .A1(new_n1590_), .B0(new_n11083_), .Y(new_n11084_));
  XOR2X1   g10828(.A(new_n11084_), .B(\a[59] ), .Y(new_n11085_));
  XOR2X1   g10829(.A(new_n11085_), .B(new_n11081_), .Y(new_n11086_));
  INVX1    g10830(.A(new_n11086_), .Y(new_n11087_));
  XOR2X1   g10831(.A(new_n11087_), .B(new_n11065_), .Y(new_n11088_));
  AOI22X1  g10832(.A0(new_n6438_), .A1(\b[28] ), .B0(new_n6437_), .B1(\b[27] ), .Y(new_n11089_));
  OAI21X1  g10833(.A0(new_n6436_), .A1(new_n1877_), .B0(new_n11089_), .Y(new_n11090_));
  AOI21X1  g10834(.A0(new_n6023_), .A1(new_n2004_), .B0(new_n11090_), .Y(new_n11091_));
  XOR2X1   g10835(.A(new_n11091_), .B(\a[56] ), .Y(new_n11092_));
  XOR2X1   g10836(.A(new_n11092_), .B(new_n11088_), .Y(new_n11093_));
  INVX1    g10837(.A(new_n11093_), .Y(new_n11094_));
  INVX1    g10838(.A(new_n10922_), .Y(new_n11095_));
  NOR2X1   g10839(.A(new_n10925_), .B(new_n10923_), .Y(new_n11096_));
  AOI21X1  g10840(.A0(new_n11095_), .A1(new_n10918_), .B0(new_n11096_), .Y(new_n11097_));
  XOR2X1   g10841(.A(new_n11097_), .B(new_n11094_), .Y(new_n11098_));
  AOI22X1  g10842(.A0(new_n5430_), .A1(\b[31] ), .B0(new_n5427_), .B1(\b[30] ), .Y(new_n11099_));
  OAI21X1  g10843(.A0(new_n5891_), .A1(new_n2359_), .B0(new_n11099_), .Y(new_n11100_));
  AOI21X1  g10844(.A0(new_n5425_), .A1(new_n2358_), .B0(new_n11100_), .Y(new_n11101_));
  XOR2X1   g10845(.A(new_n11101_), .B(\a[53] ), .Y(new_n11102_));
  XOR2X1   g10846(.A(new_n11102_), .B(new_n11098_), .Y(new_n11103_));
  INVX1    g10847(.A(new_n10930_), .Y(new_n11104_));
  NOR2X1   g10848(.A(new_n10934_), .B(new_n10931_), .Y(new_n11105_));
  AOI21X1  g10849(.A0(new_n11104_), .A1(new_n10926_), .B0(new_n11105_), .Y(new_n11106_));
  XOR2X1   g10850(.A(new_n11106_), .B(new_n11103_), .Y(new_n11107_));
  AOI22X1  g10851(.A0(new_n4880_), .A1(\b[34] ), .B0(new_n4877_), .B1(\b[33] ), .Y(new_n11108_));
  OAI21X1  g10852(.A0(new_n5291_), .A1(new_n2612_), .B0(new_n11108_), .Y(new_n11109_));
  AOI21X1  g10853(.A0(new_n4875_), .A1(new_n2759_), .B0(new_n11109_), .Y(new_n11110_));
  XOR2X1   g10854(.A(new_n11110_), .B(\a[50] ), .Y(new_n11111_));
  XOR2X1   g10855(.A(new_n11111_), .B(new_n11107_), .Y(new_n11112_));
  INVX1    g10856(.A(new_n11112_), .Y(new_n11113_));
  NOR2X1   g10857(.A(new_n10943_), .B(new_n10940_), .Y(new_n11114_));
  AOI21X1  g10858(.A0(new_n10944_), .A1(new_n10935_), .B0(new_n11114_), .Y(new_n11115_));
  XOR2X1   g10859(.A(new_n11115_), .B(new_n11113_), .Y(new_n11116_));
  AOI22X1  g10860(.A0(new_n4572_), .A1(\b[37] ), .B0(new_n4571_), .B1(\b[36] ), .Y(new_n11117_));
  OAI21X1  g10861(.A0(new_n4740_), .A1(new_n3156_), .B0(new_n11117_), .Y(new_n11118_));
  AOI21X1  g10862(.A0(new_n4375_), .A1(new_n3155_), .B0(new_n11118_), .Y(new_n11119_));
  XOR2X1   g10863(.A(new_n11119_), .B(\a[47] ), .Y(new_n11120_));
  XOR2X1   g10864(.A(new_n11120_), .B(new_n11116_), .Y(new_n11121_));
  XOR2X1   g10865(.A(new_n11121_), .B(new_n11063_), .Y(new_n11122_));
  XOR2X1   g10866(.A(new_n11122_), .B(new_n11061_), .Y(new_n11123_));
  XOR2X1   g10867(.A(new_n11123_), .B(new_n11057_), .Y(new_n11124_));
  AOI22X1  g10868(.A0(new_n3652_), .A1(\b[43] ), .B0(new_n3651_), .B1(\b[42] ), .Y(new_n11125_));
  OAI21X1  g10869(.A0(new_n3778_), .A1(new_n4015_), .B0(new_n11125_), .Y(new_n11126_));
  AOI21X1  g10870(.A0(new_n4014_), .A1(new_n3480_), .B0(new_n11126_), .Y(new_n11127_));
  XOR2X1   g10871(.A(new_n11127_), .B(\a[41] ), .Y(new_n11128_));
  XOR2X1   g10872(.A(new_n11128_), .B(new_n11124_), .Y(new_n11129_));
  NOR2X1   g10873(.A(new_n10961_), .B(new_n10957_), .Y(new_n11130_));
  AOI21X1  g10874(.A0(new_n10962_), .A1(new_n10889_), .B0(new_n11130_), .Y(new_n11131_));
  XOR2X1   g10875(.A(new_n11131_), .B(new_n11129_), .Y(new_n11132_));
  AOI22X1  g10876(.A0(new_n3204_), .A1(\b[46] ), .B0(new_n3203_), .B1(\b[45] ), .Y(new_n11133_));
  OAI21X1  g10877(.A0(new_n3321_), .A1(new_n4336_), .B0(new_n11133_), .Y(new_n11134_));
  AOI21X1  g10878(.A0(new_n4509_), .A1(new_n3080_), .B0(new_n11134_), .Y(new_n11135_));
  XOR2X1   g10879(.A(new_n11135_), .B(\a[38] ), .Y(new_n11136_));
  XOR2X1   g10880(.A(new_n11136_), .B(new_n11132_), .Y(new_n11137_));
  INVX1    g10881(.A(new_n10967_), .Y(new_n11138_));
  NOR2X1   g10882(.A(new_n10970_), .B(new_n10968_), .Y(new_n11139_));
  AOI21X1  g10883(.A0(new_n11138_), .A1(new_n10963_), .B0(new_n11139_), .Y(new_n11140_));
  XOR2X1   g10884(.A(new_n11140_), .B(new_n11137_), .Y(new_n11141_));
  AOI22X1  g10885(.A0(new_n2813_), .A1(\b[49] ), .B0(new_n2812_), .B1(\b[48] ), .Y(new_n11142_));
  OAI21X1  g10886(.A0(new_n2946_), .A1(new_n5039_), .B0(new_n11142_), .Y(new_n11143_));
  AOI21X1  g10887(.A0(new_n5038_), .A1(new_n2652_), .B0(new_n11143_), .Y(new_n11144_));
  XOR2X1   g10888(.A(new_n11144_), .B(\a[35] ), .Y(new_n11145_));
  XOR2X1   g10889(.A(new_n11145_), .B(new_n11141_), .Y(new_n11146_));
  XOR2X1   g10890(.A(new_n11146_), .B(new_n11053_), .Y(new_n11147_));
  XOR2X1   g10891(.A(new_n11147_), .B(new_n11044_), .Y(new_n11148_));
  XOR2X1   g10892(.A(new_n11148_), .B(new_n11036_), .Y(new_n11149_));
  XOR2X1   g10893(.A(new_n11149_), .B(new_n11028_), .Y(new_n11150_));
  INVX1    g10894(.A(new_n11150_), .Y(new_n11151_));
  XOR2X1   g10895(.A(new_n11019_), .B(new_n11016_), .Y(new_n11152_));
  NOR2X1   g10896(.A(new_n11152_), .B(new_n11151_), .Y(new_n11153_));
  AOI21X1  g10897(.A0(new_n11019_), .A1(new_n11016_), .B0(new_n11150_), .Y(new_n11154_));
  AOI21X1  g10898(.A0(new_n11154_), .A1(new_n11020_), .B0(new_n11153_), .Y(new_n11155_));
  XOR2X1   g10899(.A(new_n11155_), .B(new_n11012_), .Y(new_n11156_));
  XOR2X1   g10900(.A(new_n11156_), .B(new_n11008_), .Y(\f[82] ));
  OAI21X1  g10901(.A0(new_n11011_), .A1(new_n11010_), .B0(new_n11155_), .Y(new_n11158_));
  INVX1    g10902(.A(new_n11158_), .Y(new_n11159_));
  AOI21X1  g10903(.A0(new_n11007_), .A1(new_n11006_), .B0(new_n11156_), .Y(new_n11160_));
  OR2X1    g10904(.A(new_n11160_), .B(new_n11159_), .Y(new_n11161_));
  XOR2X1   g10905(.A(new_n11018_), .B(new_n1072_), .Y(new_n11162_));
  AND2X1   g10906(.A(new_n11162_), .B(new_n11016_), .Y(new_n11163_));
  OR2X1    g10907(.A(new_n11153_), .B(new_n11163_), .Y(new_n11164_));
  NOR2X1   g10908(.A(new_n11027_), .B(new_n11024_), .Y(new_n11165_));
  AOI21X1  g10909(.A0(new_n11149_), .A1(new_n11028_), .B0(new_n11165_), .Y(new_n11166_));
  AOI22X1  g10910(.A0(new_n7774_), .A1(new_n1075_), .B0(new_n1167_), .B1(\b[63] ), .Y(new_n11167_));
  XOR2X1   g10911(.A(new_n11167_), .B(new_n1072_), .Y(new_n11168_));
  XOR2X1   g10912(.A(new_n11168_), .B(new_n11166_), .Y(new_n11169_));
  AOI22X1  g10913(.A0(new_n1526_), .A1(\b[62] ), .B0(new_n1525_), .B1(\b[61] ), .Y(new_n11170_));
  OAI21X1  g10914(.A0(new_n1524_), .A1(new_n7559_), .B0(new_n11170_), .Y(new_n11171_));
  AOI21X1  g10915(.A0(new_n7558_), .A1(new_n1347_), .B0(new_n11171_), .Y(new_n11172_));
  XOR2X1   g10916(.A(new_n11172_), .B(\a[23] ), .Y(new_n11173_));
  OR2X1    g10917(.A(new_n11035_), .B(new_n11032_), .Y(new_n11174_));
  OR2X1    g10918(.A(new_n11148_), .B(new_n11036_), .Y(new_n11175_));
  AND2X1   g10919(.A(new_n11175_), .B(new_n11174_), .Y(new_n11176_));
  XOR2X1   g10920(.A(new_n11176_), .B(new_n11173_), .Y(new_n11177_));
  AOI22X1  g10921(.A0(new_n1814_), .A1(\b[59] ), .B0(new_n1813_), .B1(\b[58] ), .Y(new_n11178_));
  OAI21X1  g10922(.A0(new_n1812_), .A1(new_n6933_), .B0(new_n11178_), .Y(new_n11179_));
  AOI21X1  g10923(.A0(new_n6932_), .A1(new_n1617_), .B0(new_n11179_), .Y(new_n11180_));
  XOR2X1   g10924(.A(new_n11180_), .B(\a[26] ), .Y(new_n11181_));
  NOR2X1   g10925(.A(new_n11042_), .B(new_n11040_), .Y(new_n11182_));
  AOI21X1  g10926(.A0(new_n11147_), .A1(new_n11043_), .B0(new_n11182_), .Y(new_n11183_));
  XOR2X1   g10927(.A(new_n11183_), .B(new_n11181_), .Y(new_n11184_));
  AOI22X1  g10928(.A0(new_n2163_), .A1(\b[56] ), .B0(new_n2162_), .B1(\b[55] ), .Y(new_n11185_));
  OAI21X1  g10929(.A0(new_n2161_), .A1(new_n6148_), .B0(new_n11185_), .Y(new_n11186_));
  AOI21X1  g10930(.A0(new_n6342_), .A1(new_n1907_), .B0(new_n11186_), .Y(new_n11187_));
  XOR2X1   g10931(.A(new_n11187_), .B(\a[29] ), .Y(new_n11188_));
  OR2X1    g10932(.A(new_n11052_), .B(new_n11048_), .Y(new_n11189_));
  OR2X1    g10933(.A(new_n11146_), .B(new_n11053_), .Y(new_n11190_));
  AND2X1   g10934(.A(new_n11190_), .B(new_n11189_), .Y(new_n11191_));
  XOR2X1   g10935(.A(new_n11191_), .B(new_n11188_), .Y(new_n11192_));
  AOI22X1  g10936(.A0(new_n2545_), .A1(\b[53] ), .B0(new_n2544_), .B1(\b[52] ), .Y(new_n11193_));
  OAI21X1  g10937(.A0(new_n2543_), .A1(new_n5787_), .B0(new_n11193_), .Y(new_n11194_));
  AOI21X1  g10938(.A0(new_n5786_), .A1(new_n2260_), .B0(new_n11194_), .Y(new_n11195_));
  XOR2X1   g10939(.A(new_n11195_), .B(\a[32] ), .Y(new_n11196_));
  NOR2X1   g10940(.A(new_n11140_), .B(new_n11137_), .Y(new_n11197_));
  INVX1    g10941(.A(new_n11145_), .Y(new_n11198_));
  AOI21X1  g10942(.A0(new_n11198_), .A1(new_n11141_), .B0(new_n11197_), .Y(new_n11199_));
  XOR2X1   g10943(.A(new_n11199_), .B(new_n11196_), .Y(new_n11200_));
  AND2X1   g10944(.A(new_n11123_), .B(new_n11057_), .Y(new_n11201_));
  INVX1    g10945(.A(new_n11201_), .Y(new_n11202_));
  INVX1    g10946(.A(new_n11124_), .Y(new_n11203_));
  OAI21X1  g10947(.A0(new_n11128_), .A1(new_n11203_), .B0(new_n11202_), .Y(new_n11204_));
  AOI22X1  g10948(.A0(new_n3652_), .A1(\b[44] ), .B0(new_n3651_), .B1(\b[43] ), .Y(new_n11205_));
  OAI21X1  g10949(.A0(new_n3778_), .A1(new_n4012_), .B0(new_n11205_), .Y(new_n11206_));
  AOI21X1  g10950(.A0(new_n4178_), .A1(new_n3480_), .B0(new_n11206_), .Y(new_n11207_));
  XOR2X1   g10951(.A(new_n11207_), .B(new_n3478_), .Y(new_n11208_));
  INVX1    g10952(.A(new_n11063_), .Y(new_n11209_));
  NAND2X1  g10953(.A(new_n11121_), .B(new_n11209_), .Y(new_n11210_));
  OAI21X1  g10954(.A0(new_n11122_), .A1(new_n11061_), .B0(new_n11210_), .Y(new_n11211_));
  AOI22X1  g10955(.A0(new_n4095_), .A1(\b[41] ), .B0(new_n4094_), .B1(\b[40] ), .Y(new_n11212_));
  OAI21X1  g10956(.A0(new_n4233_), .A1(new_n3723_), .B0(new_n11212_), .Y(new_n11213_));
  AOI21X1  g10957(.A0(new_n3901_), .A1(new_n3722_), .B0(new_n11213_), .Y(new_n11214_));
  XOR2X1   g10958(.A(new_n11214_), .B(new_n3899_), .Y(new_n11215_));
  OR2X1    g10959(.A(new_n11115_), .B(new_n11112_), .Y(new_n11216_));
  OAI21X1  g10960(.A0(new_n11120_), .A1(new_n11116_), .B0(new_n11216_), .Y(new_n11217_));
  AOI22X1  g10961(.A0(new_n4572_), .A1(\b[38] ), .B0(new_n4571_), .B1(\b[37] ), .Y(new_n11218_));
  OAI21X1  g10962(.A0(new_n4740_), .A1(new_n3276_), .B0(new_n11218_), .Y(new_n11219_));
  AOI21X1  g10963(.A0(new_n4375_), .A1(new_n3275_), .B0(new_n11219_), .Y(new_n11220_));
  XOR2X1   g10964(.A(new_n11220_), .B(new_n4568_), .Y(new_n11221_));
  AND2X1   g10965(.A(new_n11106_), .B(new_n11103_), .Y(new_n11222_));
  OR2X1    g10966(.A(new_n11106_), .B(new_n11103_), .Y(new_n11223_));
  OAI21X1  g10967(.A0(new_n11111_), .A1(new_n11222_), .B0(new_n11223_), .Y(new_n11224_));
  AOI22X1  g10968(.A0(new_n4880_), .A1(\b[35] ), .B0(new_n4877_), .B1(\b[34] ), .Y(new_n11225_));
  OAI21X1  g10969(.A0(new_n5291_), .A1(new_n2893_), .B0(new_n11225_), .Y(new_n11226_));
  AOI21X1  g10970(.A0(new_n4875_), .A1(new_n2892_), .B0(new_n11226_), .Y(new_n11227_));
  XOR2X1   g10971(.A(new_n11227_), .B(new_n4873_), .Y(new_n11228_));
  NOR2X1   g10972(.A(new_n11097_), .B(new_n11094_), .Y(new_n11229_));
  INVX1    g10973(.A(new_n11102_), .Y(new_n11230_));
  AOI21X1  g10974(.A0(new_n11230_), .A1(new_n11098_), .B0(new_n11229_), .Y(new_n11231_));
  NOR2X1   g10975(.A(new_n11080_), .B(new_n11077_), .Y(new_n11232_));
  INVX1    g10976(.A(new_n11232_), .Y(new_n11233_));
  INVX1    g10977(.A(new_n11081_), .Y(new_n11234_));
  OAI21X1  g10978(.A0(new_n11085_), .A1(new_n11234_), .B0(new_n11233_), .Y(new_n11235_));
  AOI22X1  g10979(.A0(new_n6603_), .A1(\b[26] ), .B0(new_n6600_), .B1(\b[25] ), .Y(new_n11236_));
  OAI21X1  g10980(.A0(new_n6804_), .A1(new_n1588_), .B0(new_n11236_), .Y(new_n11237_));
  AOI21X1  g10981(.A0(new_n6598_), .A1(new_n1783_), .B0(new_n11237_), .Y(new_n11238_));
  XOR2X1   g10982(.A(new_n11238_), .B(new_n6596_), .Y(new_n11239_));
  OR2X1    g10983(.A(new_n11069_), .B(new_n11067_), .Y(new_n11240_));
  OAI21X1  g10984(.A0(new_n11075_), .A1(new_n11071_), .B0(new_n11240_), .Y(new_n11241_));
  AOI22X1  g10985(.A0(new_n7818_), .A1(\b[19] ), .B0(new_n7817_), .B1(\b[20] ), .Y(new_n11242_));
  XOR2X1   g10986(.A(new_n11242_), .B(new_n11066_), .Y(new_n11243_));
  AOI22X1  g10987(.A0(new_n7192_), .A1(\b[23] ), .B0(new_n7189_), .B1(\b[22] ), .Y(new_n11244_));
  OAI21X1  g10988(.A0(new_n7627_), .A1(new_n1482_), .B0(new_n11244_), .Y(new_n11245_));
  AOI21X1  g10989(.A0(new_n7187_), .A1(new_n1481_), .B0(new_n11245_), .Y(new_n11246_));
  XOR2X1   g10990(.A(new_n11246_), .B(\a[62] ), .Y(new_n11247_));
  XOR2X1   g10991(.A(new_n11247_), .B(new_n11243_), .Y(new_n11248_));
  XOR2X1   g10992(.A(new_n11248_), .B(new_n11241_), .Y(new_n11249_));
  XOR2X1   g10993(.A(new_n11249_), .B(new_n11239_), .Y(new_n11250_));
  XOR2X1   g10994(.A(new_n11250_), .B(new_n11235_), .Y(new_n11251_));
  AOI22X1  g10995(.A0(new_n6438_), .A1(\b[29] ), .B0(new_n6437_), .B1(\b[28] ), .Y(new_n11252_));
  OAI21X1  g10996(.A0(new_n6436_), .A1(new_n2126_), .B0(new_n11252_), .Y(new_n11253_));
  AOI21X1  g10997(.A0(new_n6023_), .A1(new_n2125_), .B0(new_n11253_), .Y(new_n11254_));
  XOR2X1   g10998(.A(new_n11254_), .B(\a[56] ), .Y(new_n11255_));
  XOR2X1   g10999(.A(new_n11255_), .B(new_n11251_), .Y(new_n11256_));
  OR2X1    g11000(.A(new_n11092_), .B(new_n11088_), .Y(new_n11257_));
  OR2X1    g11001(.A(new_n11086_), .B(new_n11065_), .Y(new_n11258_));
  AND2X1   g11002(.A(new_n11258_), .B(new_n11257_), .Y(new_n11259_));
  XOR2X1   g11003(.A(new_n11259_), .B(new_n11256_), .Y(new_n11260_));
  AOI22X1  g11004(.A0(new_n5430_), .A1(\b[32] ), .B0(new_n5427_), .B1(\b[31] ), .Y(new_n11261_));
  OAI21X1  g11005(.A0(new_n5891_), .A1(new_n2356_), .B0(new_n11261_), .Y(new_n11262_));
  AOI21X1  g11006(.A0(new_n5425_), .A1(new_n2495_), .B0(new_n11262_), .Y(new_n11263_));
  XOR2X1   g11007(.A(new_n11263_), .B(\a[53] ), .Y(new_n11264_));
  XOR2X1   g11008(.A(new_n11264_), .B(new_n11260_), .Y(new_n11265_));
  XOR2X1   g11009(.A(new_n11265_), .B(new_n11231_), .Y(new_n11266_));
  XOR2X1   g11010(.A(new_n11266_), .B(new_n11228_), .Y(new_n11267_));
  XOR2X1   g11011(.A(new_n11267_), .B(new_n11224_), .Y(new_n11268_));
  XOR2X1   g11012(.A(new_n11268_), .B(new_n11221_), .Y(new_n11269_));
  XOR2X1   g11013(.A(new_n11269_), .B(new_n11217_), .Y(new_n11270_));
  XOR2X1   g11014(.A(new_n11270_), .B(new_n11215_), .Y(new_n11271_));
  XOR2X1   g11015(.A(new_n11271_), .B(new_n11211_), .Y(new_n11272_));
  XOR2X1   g11016(.A(new_n11272_), .B(new_n11208_), .Y(new_n11273_));
  XOR2X1   g11017(.A(new_n11273_), .B(new_n11204_), .Y(new_n11274_));
  AOI22X1  g11018(.A0(new_n3204_), .A1(\b[47] ), .B0(new_n3203_), .B1(\b[46] ), .Y(new_n11275_));
  OAI21X1  g11019(.A0(new_n3321_), .A1(new_n4674_), .B0(new_n11275_), .Y(new_n11276_));
  AOI21X1  g11020(.A0(new_n4673_), .A1(new_n3080_), .B0(new_n11276_), .Y(new_n11277_));
  XOR2X1   g11021(.A(new_n11277_), .B(\a[38] ), .Y(new_n11278_));
  XOR2X1   g11022(.A(new_n11278_), .B(new_n11274_), .Y(new_n11279_));
  INVX1    g11023(.A(new_n11279_), .Y(new_n11280_));
  NOR2X1   g11024(.A(new_n11131_), .B(new_n11129_), .Y(new_n11281_));
  INVX1    g11025(.A(new_n11136_), .Y(new_n11282_));
  AOI21X1  g11026(.A0(new_n11282_), .A1(new_n11132_), .B0(new_n11281_), .Y(new_n11283_));
  XOR2X1   g11027(.A(new_n11283_), .B(new_n11280_), .Y(new_n11284_));
  AOI22X1  g11028(.A0(new_n2813_), .A1(\b[50] ), .B0(new_n2812_), .B1(\b[49] ), .Y(new_n11285_));
  OAI21X1  g11029(.A0(new_n2946_), .A1(new_n5036_), .B0(new_n11285_), .Y(new_n11286_));
  AOI21X1  g11030(.A0(new_n5204_), .A1(new_n2652_), .B0(new_n11286_), .Y(new_n11287_));
  XOR2X1   g11031(.A(new_n11287_), .B(\a[35] ), .Y(new_n11288_));
  XOR2X1   g11032(.A(new_n11288_), .B(new_n11284_), .Y(new_n11289_));
  XOR2X1   g11033(.A(new_n11289_), .B(new_n11200_), .Y(new_n11290_));
  XOR2X1   g11034(.A(new_n11290_), .B(new_n11192_), .Y(new_n11291_));
  INVX1    g11035(.A(new_n11291_), .Y(new_n11292_));
  XOR2X1   g11036(.A(new_n11292_), .B(new_n11184_), .Y(new_n11293_));
  XOR2X1   g11037(.A(new_n11293_), .B(new_n11177_), .Y(new_n11294_));
  XOR2X1   g11038(.A(new_n11294_), .B(new_n11169_), .Y(new_n11295_));
  XOR2X1   g11039(.A(new_n11295_), .B(new_n11164_), .Y(new_n11296_));
  XOR2X1   g11040(.A(new_n11296_), .B(new_n11161_), .Y(\f[83] ));
  NOR2X1   g11041(.A(new_n11176_), .B(new_n11173_), .Y(new_n11298_));
  INVX1    g11042(.A(new_n11293_), .Y(new_n11299_));
  AOI21X1  g11043(.A0(new_n11299_), .A1(new_n11177_), .B0(new_n11298_), .Y(new_n11300_));
  AOI22X1  g11044(.A0(new_n1526_), .A1(\b[63] ), .B0(new_n1525_), .B1(\b[62] ), .Y(new_n11301_));
  OAI21X1  g11045(.A0(new_n1524_), .A1(new_n7748_), .B0(new_n11301_), .Y(new_n11302_));
  AOI21X1  g11046(.A0(new_n7747_), .A1(new_n1347_), .B0(new_n11302_), .Y(new_n11303_));
  XOR2X1   g11047(.A(new_n11303_), .B(\a[23] ), .Y(new_n11304_));
  XOR2X1   g11048(.A(new_n11304_), .B(new_n11300_), .Y(new_n11305_));
  AOI22X1  g11049(.A0(new_n1814_), .A1(\b[60] ), .B0(new_n1813_), .B1(\b[59] ), .Y(new_n11306_));
  OAI21X1  g11050(.A0(new_n1812_), .A1(new_n6930_), .B0(new_n11306_), .Y(new_n11307_));
  AOI21X1  g11051(.A0(new_n6951_), .A1(new_n1617_), .B0(new_n11307_), .Y(new_n11308_));
  XOR2X1   g11052(.A(new_n11308_), .B(\a[26] ), .Y(new_n11309_));
  INVX1    g11053(.A(new_n11309_), .Y(new_n11310_));
  NOR2X1   g11054(.A(new_n11183_), .B(new_n11181_), .Y(new_n11311_));
  AOI21X1  g11055(.A0(new_n11291_), .A1(new_n11184_), .B0(new_n11311_), .Y(new_n11312_));
  XOR2X1   g11056(.A(new_n11312_), .B(new_n11310_), .Y(new_n11313_));
  NOR2X1   g11057(.A(new_n11191_), .B(new_n11188_), .Y(new_n11314_));
  AOI21X1  g11058(.A0(new_n11290_), .A1(new_n11192_), .B0(new_n11314_), .Y(new_n11315_));
  AOI22X1  g11059(.A0(new_n2163_), .A1(\b[57] ), .B0(new_n2162_), .B1(\b[56] ), .Y(new_n11316_));
  OAI21X1  g11060(.A0(new_n2161_), .A1(new_n6523_), .B0(new_n11316_), .Y(new_n11317_));
  AOI21X1  g11061(.A0(new_n6522_), .A1(new_n1907_), .B0(new_n11317_), .Y(new_n11318_));
  XOR2X1   g11062(.A(new_n11318_), .B(\a[29] ), .Y(new_n11319_));
  INVX1    g11063(.A(new_n11319_), .Y(new_n11320_));
  XOR2X1   g11064(.A(new_n11320_), .B(new_n11315_), .Y(new_n11321_));
  AOI22X1  g11065(.A0(new_n2545_), .A1(\b[54] ), .B0(new_n2544_), .B1(\b[53] ), .Y(new_n11322_));
  OAI21X1  g11066(.A0(new_n2543_), .A1(new_n5808_), .B0(new_n11322_), .Y(new_n11323_));
  AOI21X1  g11067(.A0(new_n5807_), .A1(new_n2260_), .B0(new_n11323_), .Y(new_n11324_));
  XOR2X1   g11068(.A(new_n11324_), .B(\a[32] ), .Y(new_n11325_));
  INVX1    g11069(.A(new_n11325_), .Y(new_n11326_));
  NOR2X1   g11070(.A(new_n11199_), .B(new_n11196_), .Y(new_n11327_));
  AOI21X1  g11071(.A0(new_n11289_), .A1(new_n11200_), .B0(new_n11327_), .Y(new_n11328_));
  XOR2X1   g11072(.A(new_n11328_), .B(new_n11326_), .Y(new_n11329_));
  NOR2X1   g11073(.A(new_n11283_), .B(new_n11279_), .Y(new_n11330_));
  INVX1    g11074(.A(new_n11330_), .Y(new_n11331_));
  OAI21X1  g11075(.A0(new_n11288_), .A1(new_n11284_), .B0(new_n11331_), .Y(new_n11332_));
  NOR2X1   g11076(.A(new_n11265_), .B(new_n11231_), .Y(new_n11333_));
  AOI21X1  g11077(.A0(new_n11266_), .A1(new_n11228_), .B0(new_n11333_), .Y(new_n11334_));
  INVX1    g11078(.A(new_n11334_), .Y(new_n11335_));
  INVX1    g11079(.A(new_n11242_), .Y(new_n11336_));
  AOI22X1  g11080(.A0(new_n7818_), .A1(\b[20] ), .B0(new_n7817_), .B1(\b[21] ), .Y(new_n11337_));
  XOR2X1   g11081(.A(new_n11337_), .B(\a[20] ), .Y(new_n11338_));
  XOR2X1   g11082(.A(new_n11338_), .B(new_n11336_), .Y(new_n11339_));
  AOI22X1  g11083(.A0(new_n7192_), .A1(\b[24] ), .B0(new_n7189_), .B1(\b[23] ), .Y(new_n11340_));
  OAI21X1  g11084(.A0(new_n7627_), .A1(new_n1479_), .B0(new_n11340_), .Y(new_n11341_));
  AOI21X1  g11085(.A0(new_n7187_), .A1(new_n1572_), .B0(new_n11341_), .Y(new_n11342_));
  XOR2X1   g11086(.A(new_n11342_), .B(\a[62] ), .Y(new_n11343_));
  XOR2X1   g11087(.A(new_n11343_), .B(new_n11339_), .Y(new_n11344_));
  NOR2X1   g11088(.A(new_n11247_), .B(new_n11243_), .Y(new_n11345_));
  AOI21X1  g11089(.A0(new_n11242_), .A1(new_n11067_), .B0(new_n11345_), .Y(new_n11346_));
  XOR2X1   g11090(.A(new_n11346_), .B(new_n11344_), .Y(new_n11347_));
  AOI22X1  g11091(.A0(new_n6603_), .A1(\b[27] ), .B0(new_n6600_), .B1(\b[26] ), .Y(new_n11348_));
  OAI21X1  g11092(.A0(new_n6804_), .A1(new_n1880_), .B0(new_n11348_), .Y(new_n11349_));
  AOI21X1  g11093(.A0(new_n6598_), .A1(new_n1879_), .B0(new_n11349_), .Y(new_n11350_));
  XOR2X1   g11094(.A(new_n11350_), .B(\a[59] ), .Y(new_n11351_));
  XOR2X1   g11095(.A(new_n11351_), .B(new_n11347_), .Y(new_n11352_));
  AND2X1   g11096(.A(new_n11248_), .B(new_n11241_), .Y(new_n11353_));
  AOI21X1  g11097(.A0(new_n11249_), .A1(new_n11239_), .B0(new_n11353_), .Y(new_n11354_));
  XOR2X1   g11098(.A(new_n11354_), .B(new_n11352_), .Y(new_n11355_));
  AOI22X1  g11099(.A0(new_n6438_), .A1(\b[30] ), .B0(new_n6437_), .B1(\b[29] ), .Y(new_n11356_));
  OAI21X1  g11100(.A0(new_n6436_), .A1(new_n2231_), .B0(new_n11356_), .Y(new_n11357_));
  AOI21X1  g11101(.A0(new_n6023_), .A1(new_n2230_), .B0(new_n11357_), .Y(new_n11358_));
  XOR2X1   g11102(.A(new_n11358_), .B(\a[56] ), .Y(new_n11359_));
  XOR2X1   g11103(.A(new_n11359_), .B(new_n11355_), .Y(new_n11360_));
  AND2X1   g11104(.A(new_n11250_), .B(new_n11235_), .Y(new_n11361_));
  INVX1    g11105(.A(new_n11255_), .Y(new_n11362_));
  AOI21X1  g11106(.A0(new_n11362_), .A1(new_n11251_), .B0(new_n11361_), .Y(new_n11363_));
  XOR2X1   g11107(.A(new_n11363_), .B(new_n11360_), .Y(new_n11364_));
  INVX1    g11108(.A(new_n11364_), .Y(new_n11365_));
  AOI22X1  g11109(.A0(new_n5430_), .A1(\b[33] ), .B0(new_n5427_), .B1(\b[32] ), .Y(new_n11366_));
  OAI21X1  g11110(.A0(new_n5891_), .A1(new_n2615_), .B0(new_n11366_), .Y(new_n11367_));
  AOI21X1  g11111(.A0(new_n5425_), .A1(new_n2614_), .B0(new_n11367_), .Y(new_n11368_));
  XOR2X1   g11112(.A(new_n11368_), .B(\a[53] ), .Y(new_n11369_));
  AOI21X1  g11113(.A0(new_n11258_), .A1(new_n11257_), .B0(new_n11256_), .Y(new_n11370_));
  INVX1    g11114(.A(new_n11264_), .Y(new_n11371_));
  AOI21X1  g11115(.A0(new_n11371_), .A1(new_n11260_), .B0(new_n11370_), .Y(new_n11372_));
  XOR2X1   g11116(.A(new_n11372_), .B(new_n11369_), .Y(new_n11373_));
  XOR2X1   g11117(.A(new_n11373_), .B(new_n11365_), .Y(new_n11374_));
  AOI22X1  g11118(.A0(new_n4880_), .A1(\b[36] ), .B0(new_n4877_), .B1(\b[35] ), .Y(new_n11375_));
  OAI21X1  g11119(.A0(new_n5291_), .A1(new_n2890_), .B0(new_n11375_), .Y(new_n11376_));
  AOI21X1  g11120(.A0(new_n4875_), .A1(new_n3015_), .B0(new_n11376_), .Y(new_n11377_));
  XOR2X1   g11121(.A(new_n11377_), .B(\a[50] ), .Y(new_n11378_));
  XOR2X1   g11122(.A(new_n11378_), .B(new_n11374_), .Y(new_n11379_));
  XOR2X1   g11123(.A(new_n11379_), .B(new_n11335_), .Y(new_n11380_));
  AOI22X1  g11124(.A0(new_n4572_), .A1(\b[39] ), .B0(new_n4571_), .B1(\b[38] ), .Y(new_n11381_));
  OAI21X1  g11125(.A0(new_n4740_), .A1(new_n3413_), .B0(new_n11381_), .Y(new_n11382_));
  AOI21X1  g11126(.A0(new_n4375_), .A1(new_n3412_), .B0(new_n11382_), .Y(new_n11383_));
  XOR2X1   g11127(.A(new_n11383_), .B(\a[47] ), .Y(new_n11384_));
  XOR2X1   g11128(.A(new_n11384_), .B(new_n11380_), .Y(new_n11385_));
  AND2X1   g11129(.A(new_n11267_), .B(new_n11224_), .Y(new_n11386_));
  AOI21X1  g11130(.A0(new_n11268_), .A1(new_n11221_), .B0(new_n11386_), .Y(new_n11387_));
  XOR2X1   g11131(.A(new_n11387_), .B(new_n11385_), .Y(new_n11388_));
  AOI22X1  g11132(.A0(new_n4095_), .A1(\b[42] ), .B0(new_n4094_), .B1(\b[41] ), .Y(new_n11389_));
  OAI21X1  g11133(.A0(new_n4233_), .A1(new_n3720_), .B0(new_n11389_), .Y(new_n11390_));
  AOI21X1  g11134(.A0(new_n3901_), .A1(new_n3860_), .B0(new_n11390_), .Y(new_n11391_));
  XOR2X1   g11135(.A(new_n11391_), .B(\a[44] ), .Y(new_n11392_));
  XOR2X1   g11136(.A(new_n11392_), .B(new_n11388_), .Y(new_n11393_));
  AND2X1   g11137(.A(new_n11269_), .B(new_n11217_), .Y(new_n11394_));
  AOI21X1  g11138(.A0(new_n11270_), .A1(new_n11215_), .B0(new_n11394_), .Y(new_n11395_));
  XOR2X1   g11139(.A(new_n11395_), .B(new_n11393_), .Y(new_n11396_));
  AOI22X1  g11140(.A0(new_n3652_), .A1(\b[45] ), .B0(new_n3651_), .B1(\b[44] ), .Y(new_n11397_));
  OAI21X1  g11141(.A0(new_n3778_), .A1(new_n4339_), .B0(new_n11397_), .Y(new_n11398_));
  AOI21X1  g11142(.A0(new_n4338_), .A1(new_n3480_), .B0(new_n11398_), .Y(new_n11399_));
  XOR2X1   g11143(.A(new_n11399_), .B(\a[41] ), .Y(new_n11400_));
  XOR2X1   g11144(.A(new_n11400_), .B(new_n11396_), .Y(new_n11401_));
  AND2X1   g11145(.A(new_n11271_), .B(new_n11211_), .Y(new_n11402_));
  AOI21X1  g11146(.A0(new_n11272_), .A1(new_n11208_), .B0(new_n11402_), .Y(new_n11403_));
  XOR2X1   g11147(.A(new_n11403_), .B(new_n11401_), .Y(new_n11404_));
  AOI22X1  g11148(.A0(new_n3204_), .A1(\b[48] ), .B0(new_n3203_), .B1(\b[47] ), .Y(new_n11405_));
  OAI21X1  g11149(.A0(new_n3321_), .A1(new_n4693_), .B0(new_n11405_), .Y(new_n11406_));
  AOI21X1  g11150(.A0(new_n4692_), .A1(new_n3080_), .B0(new_n11406_), .Y(new_n11407_));
  XOR2X1   g11151(.A(new_n11407_), .B(\a[38] ), .Y(new_n11408_));
  XOR2X1   g11152(.A(new_n11408_), .B(new_n11404_), .Y(new_n11409_));
  AND2X1   g11153(.A(new_n11273_), .B(new_n11204_), .Y(new_n11410_));
  INVX1    g11154(.A(new_n11278_), .Y(new_n11411_));
  AOI21X1  g11155(.A0(new_n11411_), .A1(new_n11274_), .B0(new_n11410_), .Y(new_n11412_));
  XOR2X1   g11156(.A(new_n11412_), .B(new_n11409_), .Y(new_n11413_));
  INVX1    g11157(.A(new_n11413_), .Y(new_n11414_));
  AOI22X1  g11158(.A0(new_n2813_), .A1(\b[51] ), .B0(new_n2812_), .B1(\b[50] ), .Y(new_n11415_));
  OAI21X1  g11159(.A0(new_n2946_), .A1(new_n5237_), .B0(new_n11415_), .Y(new_n11416_));
  AOI21X1  g11160(.A0(new_n5236_), .A1(new_n2652_), .B0(new_n11416_), .Y(new_n11417_));
  XOR2X1   g11161(.A(new_n11417_), .B(\a[35] ), .Y(new_n11418_));
  AND2X1   g11162(.A(new_n11418_), .B(new_n11414_), .Y(new_n11419_));
  INVX1    g11163(.A(new_n11419_), .Y(new_n11420_));
  OAI21X1  g11164(.A0(new_n11418_), .A1(new_n11414_), .B0(new_n11332_), .Y(new_n11421_));
  OR2X1    g11165(.A(new_n11421_), .B(new_n11419_), .Y(new_n11422_));
  NOR2X1   g11166(.A(new_n11418_), .B(new_n11414_), .Y(new_n11423_));
  AOI21X1  g11167(.A0(new_n11420_), .A1(new_n11332_), .B0(new_n11423_), .Y(new_n11424_));
  AOI22X1  g11168(.A0(new_n11424_), .A1(new_n11420_), .B0(new_n11422_), .B1(new_n11332_), .Y(new_n11425_));
  XOR2X1   g11169(.A(new_n11425_), .B(new_n11329_), .Y(new_n11426_));
  XOR2X1   g11170(.A(new_n11426_), .B(new_n11321_), .Y(new_n11427_));
  XOR2X1   g11171(.A(new_n11427_), .B(new_n11313_), .Y(new_n11428_));
  XOR2X1   g11172(.A(new_n11428_), .B(new_n11305_), .Y(new_n11429_));
  INVX1    g11173(.A(new_n11429_), .Y(new_n11430_));
  INVX1    g11174(.A(new_n11166_), .Y(new_n11431_));
  NOR2X1   g11175(.A(new_n11294_), .B(new_n11169_), .Y(new_n11432_));
  AOI21X1  g11176(.A0(new_n11168_), .A1(new_n11431_), .B0(new_n11432_), .Y(new_n11433_));
  XOR2X1   g11177(.A(new_n11433_), .B(new_n11430_), .Y(new_n11434_));
  INVX1    g11178(.A(new_n11434_), .Y(new_n11435_));
  AND2X1   g11179(.A(new_n11295_), .B(new_n11164_), .Y(new_n11436_));
  INVX1    g11180(.A(new_n11436_), .Y(new_n11437_));
  OAI21X1  g11181(.A0(new_n11160_), .A1(new_n11159_), .B0(new_n11296_), .Y(new_n11438_));
  AND2X1   g11182(.A(new_n11438_), .B(new_n11437_), .Y(new_n11439_));
  XOR2X1   g11183(.A(new_n11439_), .B(new_n11435_), .Y(\f[84] ));
  NOR2X1   g11184(.A(new_n11312_), .B(new_n11309_), .Y(new_n11441_));
  NOR2X1   g11185(.A(new_n11427_), .B(new_n11313_), .Y(new_n11442_));
  NOR2X1   g11186(.A(new_n11442_), .B(new_n11441_), .Y(new_n11443_));
  OAI22X1  g11187(.A0(new_n1524_), .A1(new_n7745_), .B0(new_n1350_), .B1(new_n7772_), .Y(new_n11444_));
  AOI21X1  g11188(.A0(new_n7775_), .A1(new_n1347_), .B0(new_n11444_), .Y(new_n11445_));
  XOR2X1   g11189(.A(new_n11445_), .B(\a[23] ), .Y(new_n11446_));
  XOR2X1   g11190(.A(new_n11446_), .B(new_n11443_), .Y(new_n11447_));
  AOI22X1  g11191(.A0(new_n1814_), .A1(\b[61] ), .B0(new_n1813_), .B1(\b[60] ), .Y(new_n11448_));
  OAI21X1  g11192(.A0(new_n1812_), .A1(new_n7339_), .B0(new_n11448_), .Y(new_n11449_));
  AOI21X1  g11193(.A0(new_n7338_), .A1(new_n1617_), .B0(new_n11449_), .Y(new_n11450_));
  XOR2X1   g11194(.A(new_n11450_), .B(\a[26] ), .Y(new_n11451_));
  INVX1    g11195(.A(new_n11451_), .Y(new_n11452_));
  INVX1    g11196(.A(new_n11321_), .Y(new_n11453_));
  NOR2X1   g11197(.A(new_n11319_), .B(new_n11315_), .Y(new_n11454_));
  AOI21X1  g11198(.A0(new_n11426_), .A1(new_n11453_), .B0(new_n11454_), .Y(new_n11455_));
  XOR2X1   g11199(.A(new_n11455_), .B(new_n11452_), .Y(new_n11456_));
  NOR2X1   g11200(.A(new_n11328_), .B(new_n11325_), .Y(new_n11457_));
  NOR2X1   g11201(.A(new_n11425_), .B(new_n11329_), .Y(new_n11458_));
  NOR2X1   g11202(.A(new_n11458_), .B(new_n11457_), .Y(new_n11459_));
  OAI22X1  g11203(.A0(new_n1913_), .A1(new_n6930_), .B0(new_n1910_), .B1(new_n6933_), .Y(new_n11460_));
  AOI21X1  g11204(.A0(new_n2045_), .A1(\b[56] ), .B0(new_n11460_), .Y(new_n11461_));
  OAI21X1  g11205(.A0(new_n8540_), .A1(new_n2043_), .B0(new_n11461_), .Y(new_n11462_));
  XOR2X1   g11206(.A(new_n11462_), .B(new_n1911_), .Y(new_n11463_));
  XOR2X1   g11207(.A(new_n11463_), .B(new_n11459_), .Y(new_n11464_));
  INVX1    g11208(.A(new_n11464_), .Y(new_n11465_));
  INVX1    g11209(.A(new_n11424_), .Y(new_n11466_));
  AOI22X1  g11210(.A0(new_n2545_), .A1(\b[55] ), .B0(new_n2544_), .B1(\b[54] ), .Y(new_n11467_));
  OAI21X1  g11211(.A0(new_n2543_), .A1(new_n6151_), .B0(new_n11467_), .Y(new_n11468_));
  AOI21X1  g11212(.A0(new_n6150_), .A1(new_n2260_), .B0(new_n11468_), .Y(new_n11469_));
  XOR2X1   g11213(.A(new_n11469_), .B(\a[32] ), .Y(new_n11470_));
  XOR2X1   g11214(.A(new_n11470_), .B(new_n11466_), .Y(new_n11471_));
  XOR2X1   g11215(.A(new_n11383_), .B(new_n4568_), .Y(new_n11472_));
  NOR2X1   g11216(.A(new_n11387_), .B(new_n11385_), .Y(new_n11473_));
  AOI21X1  g11217(.A0(new_n11472_), .A1(new_n11380_), .B0(new_n11473_), .Y(new_n11474_));
  INVX1    g11218(.A(new_n11474_), .Y(new_n11475_));
  AOI22X1  g11219(.A0(new_n4572_), .A1(\b[40] ), .B0(new_n4571_), .B1(\b[39] ), .Y(new_n11476_));
  OAI21X1  g11220(.A0(new_n4740_), .A1(new_n3575_), .B0(new_n11476_), .Y(new_n11477_));
  AOI21X1  g11221(.A0(new_n4375_), .A1(new_n3574_), .B0(new_n11477_), .Y(new_n11478_));
  XOR2X1   g11222(.A(new_n11478_), .B(\a[47] ), .Y(new_n11479_));
  NOR2X1   g11223(.A(new_n11378_), .B(new_n11374_), .Y(new_n11480_));
  AOI21X1  g11224(.A0(new_n11379_), .A1(new_n11335_), .B0(new_n11480_), .Y(new_n11481_));
  INVX1    g11225(.A(new_n11347_), .Y(new_n11482_));
  NOR2X1   g11226(.A(new_n11351_), .B(new_n11482_), .Y(new_n11483_));
  NOR2X1   g11227(.A(new_n11354_), .B(new_n11352_), .Y(new_n11484_));
  NOR2X1   g11228(.A(new_n11484_), .B(new_n11483_), .Y(new_n11485_));
  INVX1    g11229(.A(new_n11485_), .Y(new_n11486_));
  AOI22X1  g11230(.A0(new_n6603_), .A1(\b[28] ), .B0(new_n6600_), .B1(\b[27] ), .Y(new_n11487_));
  OAI21X1  g11231(.A0(new_n6804_), .A1(new_n1877_), .B0(new_n11487_), .Y(new_n11488_));
  AOI21X1  g11232(.A0(new_n6598_), .A1(new_n2004_), .B0(new_n11488_), .Y(new_n11489_));
  XOR2X1   g11233(.A(new_n11489_), .B(new_n6596_), .Y(new_n11490_));
  INVX1    g11234(.A(new_n11339_), .Y(new_n11491_));
  OR2X1    g11235(.A(new_n11343_), .B(new_n11491_), .Y(new_n11492_));
  OAI21X1  g11236(.A0(new_n11346_), .A1(new_n11344_), .B0(new_n11492_), .Y(new_n11493_));
  AOI22X1  g11237(.A0(new_n7818_), .A1(\b[21] ), .B0(new_n7817_), .B1(\b[22] ), .Y(new_n11494_));
  NOR2X1   g11238(.A(new_n11337_), .B(\a[20] ), .Y(new_n11495_));
  AOI21X1  g11239(.A0(new_n11338_), .A1(new_n11336_), .B0(new_n11495_), .Y(new_n11496_));
  XOR2X1   g11240(.A(new_n11496_), .B(new_n11494_), .Y(new_n11497_));
  AOI22X1  g11241(.A0(new_n7192_), .A1(\b[25] ), .B0(new_n7189_), .B1(\b[24] ), .Y(new_n11498_));
  OAI21X1  g11242(.A0(new_n7627_), .A1(new_n1591_), .B0(new_n11498_), .Y(new_n11499_));
  AOI21X1  g11243(.A0(new_n7187_), .A1(new_n1590_), .B0(new_n11499_), .Y(new_n11500_));
  XOR2X1   g11244(.A(new_n11500_), .B(\a[62] ), .Y(new_n11501_));
  XOR2X1   g11245(.A(new_n11501_), .B(new_n11497_), .Y(new_n11502_));
  XOR2X1   g11246(.A(new_n11502_), .B(new_n11493_), .Y(new_n11503_));
  XOR2X1   g11247(.A(new_n11503_), .B(new_n11490_), .Y(new_n11504_));
  XOR2X1   g11248(.A(new_n11504_), .B(new_n11486_), .Y(new_n11505_));
  AOI22X1  g11249(.A0(new_n6438_), .A1(\b[31] ), .B0(new_n6437_), .B1(\b[30] ), .Y(new_n11506_));
  OAI21X1  g11250(.A0(new_n6436_), .A1(new_n2359_), .B0(new_n11506_), .Y(new_n11507_));
  AOI21X1  g11251(.A0(new_n6023_), .A1(new_n2358_), .B0(new_n11507_), .Y(new_n11508_));
  XOR2X1   g11252(.A(new_n11508_), .B(\a[56] ), .Y(new_n11509_));
  XOR2X1   g11253(.A(new_n11509_), .B(new_n11505_), .Y(new_n11510_));
  INVX1    g11254(.A(new_n11359_), .Y(new_n11511_));
  NOR2X1   g11255(.A(new_n11363_), .B(new_n11360_), .Y(new_n11512_));
  AOI21X1  g11256(.A0(new_n11511_), .A1(new_n11355_), .B0(new_n11512_), .Y(new_n11513_));
  XOR2X1   g11257(.A(new_n11513_), .B(new_n11510_), .Y(new_n11514_));
  AOI22X1  g11258(.A0(new_n5430_), .A1(\b[34] ), .B0(new_n5427_), .B1(\b[33] ), .Y(new_n11515_));
  OAI21X1  g11259(.A0(new_n5891_), .A1(new_n2612_), .B0(new_n11515_), .Y(new_n11516_));
  AOI21X1  g11260(.A0(new_n5425_), .A1(new_n2759_), .B0(new_n11516_), .Y(new_n11517_));
  XOR2X1   g11261(.A(new_n11517_), .B(\a[53] ), .Y(new_n11518_));
  XOR2X1   g11262(.A(new_n11518_), .B(new_n11514_), .Y(new_n11519_));
  INVX1    g11263(.A(new_n11519_), .Y(new_n11520_));
  NOR2X1   g11264(.A(new_n11372_), .B(new_n11369_), .Y(new_n11521_));
  AOI21X1  g11265(.A0(new_n11373_), .A1(new_n11364_), .B0(new_n11521_), .Y(new_n11522_));
  XOR2X1   g11266(.A(new_n11522_), .B(new_n11520_), .Y(new_n11523_));
  AOI22X1  g11267(.A0(new_n4880_), .A1(\b[37] ), .B0(new_n4877_), .B1(\b[36] ), .Y(new_n11524_));
  OAI21X1  g11268(.A0(new_n5291_), .A1(new_n3156_), .B0(new_n11524_), .Y(new_n11525_));
  AOI21X1  g11269(.A0(new_n4875_), .A1(new_n3155_), .B0(new_n11525_), .Y(new_n11526_));
  XOR2X1   g11270(.A(new_n11526_), .B(\a[50] ), .Y(new_n11527_));
  XOR2X1   g11271(.A(new_n11527_), .B(new_n11523_), .Y(new_n11528_));
  XOR2X1   g11272(.A(new_n11528_), .B(new_n11481_), .Y(new_n11529_));
  XOR2X1   g11273(.A(new_n11529_), .B(new_n11479_), .Y(new_n11530_));
  XOR2X1   g11274(.A(new_n11530_), .B(new_n11475_), .Y(new_n11531_));
  AOI22X1  g11275(.A0(new_n4095_), .A1(\b[43] ), .B0(new_n4094_), .B1(\b[42] ), .Y(new_n11532_));
  OAI21X1  g11276(.A0(new_n4233_), .A1(new_n4015_), .B0(new_n11532_), .Y(new_n11533_));
  AOI21X1  g11277(.A0(new_n4014_), .A1(new_n3901_), .B0(new_n11533_), .Y(new_n11534_));
  XOR2X1   g11278(.A(new_n11534_), .B(\a[44] ), .Y(new_n11535_));
  XOR2X1   g11279(.A(new_n11535_), .B(new_n11531_), .Y(new_n11536_));
  INVX1    g11280(.A(new_n11392_), .Y(new_n11537_));
  NOR2X1   g11281(.A(new_n11395_), .B(new_n11393_), .Y(new_n11538_));
  AOI21X1  g11282(.A0(new_n11537_), .A1(new_n11388_), .B0(new_n11538_), .Y(new_n11539_));
  XOR2X1   g11283(.A(new_n11539_), .B(new_n11536_), .Y(new_n11540_));
  AOI22X1  g11284(.A0(new_n3652_), .A1(\b[46] ), .B0(new_n3651_), .B1(\b[45] ), .Y(new_n11541_));
  OAI21X1  g11285(.A0(new_n3778_), .A1(new_n4336_), .B0(new_n11541_), .Y(new_n11542_));
  AOI21X1  g11286(.A0(new_n4509_), .A1(new_n3480_), .B0(new_n11542_), .Y(new_n11543_));
  XOR2X1   g11287(.A(new_n11543_), .B(\a[41] ), .Y(new_n11544_));
  XOR2X1   g11288(.A(new_n11544_), .B(new_n11540_), .Y(new_n11545_));
  INVX1    g11289(.A(new_n11400_), .Y(new_n11546_));
  NOR2X1   g11290(.A(new_n11403_), .B(new_n11401_), .Y(new_n11547_));
  AOI21X1  g11291(.A0(new_n11546_), .A1(new_n11396_), .B0(new_n11547_), .Y(new_n11548_));
  XOR2X1   g11292(.A(new_n11548_), .B(new_n11545_), .Y(new_n11549_));
  AOI22X1  g11293(.A0(new_n3204_), .A1(\b[49] ), .B0(new_n3203_), .B1(\b[48] ), .Y(new_n11550_));
  OAI21X1  g11294(.A0(new_n3321_), .A1(new_n5039_), .B0(new_n11550_), .Y(new_n11551_));
  AOI21X1  g11295(.A0(new_n5038_), .A1(new_n3080_), .B0(new_n11551_), .Y(new_n11552_));
  XOR2X1   g11296(.A(new_n11552_), .B(\a[38] ), .Y(new_n11553_));
  XOR2X1   g11297(.A(new_n11553_), .B(new_n11549_), .Y(new_n11554_));
  INVX1    g11298(.A(new_n11408_), .Y(new_n11555_));
  NOR2X1   g11299(.A(new_n11412_), .B(new_n11409_), .Y(new_n11556_));
  AOI21X1  g11300(.A0(new_n11555_), .A1(new_n11404_), .B0(new_n11556_), .Y(new_n11557_));
  XOR2X1   g11301(.A(new_n11557_), .B(new_n11554_), .Y(new_n11558_));
  AOI22X1  g11302(.A0(new_n2813_), .A1(\b[52] ), .B0(new_n2812_), .B1(\b[51] ), .Y(new_n11559_));
  OAI21X1  g11303(.A0(new_n2946_), .A1(new_n5234_), .B0(new_n11559_), .Y(new_n11560_));
  AOI21X1  g11304(.A0(new_n5590_), .A1(new_n2652_), .B0(new_n11560_), .Y(new_n11561_));
  XOR2X1   g11305(.A(new_n11561_), .B(\a[35] ), .Y(new_n11562_));
  XOR2X1   g11306(.A(new_n11562_), .B(new_n11558_), .Y(new_n11563_));
  XOR2X1   g11307(.A(new_n11563_), .B(new_n11471_), .Y(new_n11564_));
  XOR2X1   g11308(.A(new_n11564_), .B(new_n11465_), .Y(new_n11565_));
  XOR2X1   g11309(.A(new_n11565_), .B(new_n11456_), .Y(new_n11566_));
  XOR2X1   g11310(.A(new_n11566_), .B(new_n11447_), .Y(new_n11567_));
  INVX1    g11311(.A(new_n11567_), .Y(new_n11568_));
  NOR2X1   g11312(.A(new_n11304_), .B(new_n11300_), .Y(new_n11569_));
  AOI21X1  g11313(.A0(new_n11428_), .A1(new_n11305_), .B0(new_n11569_), .Y(new_n11570_));
  XOR2X1   g11314(.A(new_n11570_), .B(new_n11568_), .Y(new_n11571_));
  NOR2X1   g11315(.A(new_n11433_), .B(new_n11430_), .Y(new_n11572_));
  AOI21X1  g11316(.A0(new_n11438_), .A1(new_n11437_), .B0(new_n11435_), .Y(new_n11573_));
  OR2X1    g11317(.A(new_n11573_), .B(new_n11572_), .Y(new_n11574_));
  XOR2X1   g11318(.A(new_n11574_), .B(new_n11571_), .Y(\f[85] ));
  OR2X1    g11319(.A(new_n11570_), .B(new_n11568_), .Y(new_n11576_));
  OAI21X1  g11320(.A0(new_n11573_), .A1(new_n11572_), .B0(new_n11571_), .Y(new_n11577_));
  AND2X1   g11321(.A(new_n11577_), .B(new_n11576_), .Y(new_n11578_));
  NOR2X1   g11322(.A(new_n11446_), .B(new_n11443_), .Y(new_n11579_));
  AOI21X1  g11323(.A0(new_n11566_), .A1(new_n11447_), .B0(new_n11579_), .Y(new_n11580_));
  NOR2X1   g11324(.A(new_n11455_), .B(new_n11451_), .Y(new_n11581_));
  INVX1    g11325(.A(new_n11581_), .Y(new_n11582_));
  OAI21X1  g11326(.A0(new_n11565_), .A1(new_n11456_), .B0(new_n11582_), .Y(new_n11583_));
  AOI22X1  g11327(.A0(new_n7774_), .A1(new_n1347_), .B0(new_n1430_), .B1(\b[63] ), .Y(new_n11584_));
  XOR2X1   g11328(.A(new_n11584_), .B(\a[23] ), .Y(new_n11585_));
  XOR2X1   g11329(.A(new_n11585_), .B(new_n11583_), .Y(new_n11586_));
  AOI22X1  g11330(.A0(new_n1814_), .A1(\b[62] ), .B0(new_n1813_), .B1(\b[61] ), .Y(new_n11587_));
  OAI21X1  g11331(.A0(new_n1812_), .A1(new_n7559_), .B0(new_n11587_), .Y(new_n11588_));
  AOI21X1  g11332(.A0(new_n7558_), .A1(new_n1617_), .B0(new_n11588_), .Y(new_n11589_));
  XOR2X1   g11333(.A(new_n11589_), .B(\a[26] ), .Y(new_n11590_));
  NOR2X1   g11334(.A(new_n11463_), .B(new_n11459_), .Y(new_n11591_));
  AOI21X1  g11335(.A0(new_n11564_), .A1(new_n11464_), .B0(new_n11591_), .Y(new_n11592_));
  XOR2X1   g11336(.A(new_n11592_), .B(new_n11590_), .Y(new_n11593_));
  AOI22X1  g11337(.A0(new_n2163_), .A1(\b[59] ), .B0(new_n2162_), .B1(\b[58] ), .Y(new_n11594_));
  OAI21X1  g11338(.A0(new_n2161_), .A1(new_n6933_), .B0(new_n11594_), .Y(new_n11595_));
  AOI21X1  g11339(.A0(new_n6932_), .A1(new_n1907_), .B0(new_n11595_), .Y(new_n11596_));
  XOR2X1   g11340(.A(new_n11596_), .B(\a[29] ), .Y(new_n11597_));
  OR2X1    g11341(.A(new_n11563_), .B(new_n11471_), .Y(new_n11598_));
  OR2X1    g11342(.A(new_n11470_), .B(new_n11424_), .Y(new_n11599_));
  AND2X1   g11343(.A(new_n11599_), .B(new_n11598_), .Y(new_n11600_));
  XOR2X1   g11344(.A(new_n11600_), .B(new_n11597_), .Y(new_n11601_));
  AOI22X1  g11345(.A0(new_n2545_), .A1(\b[56] ), .B0(new_n2544_), .B1(\b[55] ), .Y(new_n11602_));
  OAI21X1  g11346(.A0(new_n2543_), .A1(new_n6148_), .B0(new_n11602_), .Y(new_n11603_));
  AOI21X1  g11347(.A0(new_n6342_), .A1(new_n2260_), .B0(new_n11603_), .Y(new_n11604_));
  XOR2X1   g11348(.A(new_n11604_), .B(\a[32] ), .Y(new_n11605_));
  NOR2X1   g11349(.A(new_n11557_), .B(new_n11554_), .Y(new_n11606_));
  INVX1    g11350(.A(new_n11562_), .Y(new_n11607_));
  AOI21X1  g11351(.A0(new_n11607_), .A1(new_n11558_), .B0(new_n11606_), .Y(new_n11608_));
  XOR2X1   g11352(.A(new_n11608_), .B(new_n11605_), .Y(new_n11609_));
  AOI22X1  g11353(.A0(new_n2813_), .A1(\b[53] ), .B0(new_n2812_), .B1(\b[52] ), .Y(new_n11610_));
  OAI21X1  g11354(.A0(new_n2946_), .A1(new_n5787_), .B0(new_n11610_), .Y(new_n11611_));
  AOI21X1  g11355(.A0(new_n5786_), .A1(new_n2652_), .B0(new_n11611_), .Y(new_n11612_));
  XOR2X1   g11356(.A(new_n11612_), .B(\a[35] ), .Y(new_n11613_));
  NOR2X1   g11357(.A(new_n11548_), .B(new_n11545_), .Y(new_n11614_));
  INVX1    g11358(.A(new_n11614_), .Y(new_n11615_));
  INVX1    g11359(.A(new_n11549_), .Y(new_n11616_));
  OAI21X1  g11360(.A0(new_n11553_), .A1(new_n11616_), .B0(new_n11615_), .Y(new_n11617_));
  AND2X1   g11361(.A(new_n11530_), .B(new_n11475_), .Y(new_n11618_));
  INVX1    g11362(.A(new_n11618_), .Y(new_n11619_));
  INVX1    g11363(.A(new_n11531_), .Y(new_n11620_));
  OAI21X1  g11364(.A0(new_n11535_), .A1(new_n11620_), .B0(new_n11619_), .Y(new_n11621_));
  AOI22X1  g11365(.A0(new_n4095_), .A1(\b[44] ), .B0(new_n4094_), .B1(\b[43] ), .Y(new_n11622_));
  OAI21X1  g11366(.A0(new_n4233_), .A1(new_n4012_), .B0(new_n11622_), .Y(new_n11623_));
  AOI21X1  g11367(.A0(new_n4178_), .A1(new_n3901_), .B0(new_n11623_), .Y(new_n11624_));
  XOR2X1   g11368(.A(new_n11624_), .B(new_n3899_), .Y(new_n11625_));
  INVX1    g11369(.A(new_n11481_), .Y(new_n11626_));
  NOR2X1   g11370(.A(new_n11529_), .B(new_n11479_), .Y(new_n11627_));
  AOI21X1  g11371(.A0(new_n11528_), .A1(new_n11626_), .B0(new_n11627_), .Y(new_n11628_));
  NOR2X1   g11372(.A(new_n11513_), .B(new_n11510_), .Y(new_n11629_));
  INVX1    g11373(.A(new_n11629_), .Y(new_n11630_));
  INVX1    g11374(.A(new_n11514_), .Y(new_n11631_));
  OAI21X1  g11375(.A0(new_n11518_), .A1(new_n11631_), .B0(new_n11630_), .Y(new_n11632_));
  AOI22X1  g11376(.A0(new_n5430_), .A1(\b[35] ), .B0(new_n5427_), .B1(\b[34] ), .Y(new_n11633_));
  OAI21X1  g11377(.A0(new_n5891_), .A1(new_n2893_), .B0(new_n11633_), .Y(new_n11634_));
  AOI21X1  g11378(.A0(new_n5425_), .A1(new_n2892_), .B0(new_n11634_), .Y(new_n11635_));
  XOR2X1   g11379(.A(new_n11635_), .B(new_n5423_), .Y(new_n11636_));
  OAI21X1  g11380(.A0(new_n11484_), .A1(new_n11483_), .B0(new_n11504_), .Y(new_n11637_));
  NOR3X1   g11381(.A(new_n11504_), .B(new_n11484_), .C(new_n11483_), .Y(new_n11638_));
  OAI21X1  g11382(.A0(new_n11509_), .A1(new_n11638_), .B0(new_n11637_), .Y(new_n11639_));
  INVX1    g11383(.A(new_n11494_), .Y(new_n11640_));
  NOR2X1   g11384(.A(new_n11496_), .B(new_n11640_), .Y(new_n11641_));
  INVX1    g11385(.A(new_n11641_), .Y(new_n11642_));
  OAI21X1  g11386(.A0(new_n11501_), .A1(new_n11497_), .B0(new_n11642_), .Y(new_n11643_));
  AOI22X1  g11387(.A0(new_n7818_), .A1(\b[22] ), .B0(new_n7817_), .B1(\b[23] ), .Y(new_n11644_));
  XOR2X1   g11388(.A(new_n11644_), .B(new_n11494_), .Y(new_n11645_));
  AOI22X1  g11389(.A0(new_n7192_), .A1(\b[26] ), .B0(new_n7189_), .B1(\b[25] ), .Y(new_n11646_));
  OAI21X1  g11390(.A0(new_n7627_), .A1(new_n1588_), .B0(new_n11646_), .Y(new_n11647_));
  AOI21X1  g11391(.A0(new_n7187_), .A1(new_n1783_), .B0(new_n11647_), .Y(new_n11648_));
  XOR2X1   g11392(.A(new_n11648_), .B(\a[62] ), .Y(new_n11649_));
  XOR2X1   g11393(.A(new_n11649_), .B(new_n11645_), .Y(new_n11650_));
  XOR2X1   g11394(.A(new_n11650_), .B(new_n11643_), .Y(new_n11651_));
  AOI22X1  g11395(.A0(new_n6603_), .A1(\b[29] ), .B0(new_n6600_), .B1(\b[28] ), .Y(new_n11652_));
  OAI21X1  g11396(.A0(new_n6804_), .A1(new_n2126_), .B0(new_n11652_), .Y(new_n11653_));
  AOI21X1  g11397(.A0(new_n6598_), .A1(new_n2125_), .B0(new_n11653_), .Y(new_n11654_));
  XOR2X1   g11398(.A(new_n11654_), .B(\a[59] ), .Y(new_n11655_));
  XOR2X1   g11399(.A(new_n11655_), .B(new_n11651_), .Y(new_n11656_));
  INVX1    g11400(.A(new_n11656_), .Y(new_n11657_));
  AND2X1   g11401(.A(new_n11502_), .B(new_n11493_), .Y(new_n11658_));
  AOI21X1  g11402(.A0(new_n11503_), .A1(new_n11490_), .B0(new_n11658_), .Y(new_n11659_));
  XOR2X1   g11403(.A(new_n11659_), .B(new_n11657_), .Y(new_n11660_));
  AOI22X1  g11404(.A0(new_n6438_), .A1(\b[32] ), .B0(new_n6437_), .B1(\b[31] ), .Y(new_n11661_));
  OAI21X1  g11405(.A0(new_n6436_), .A1(new_n2356_), .B0(new_n11661_), .Y(new_n11662_));
  AOI21X1  g11406(.A0(new_n6023_), .A1(new_n2495_), .B0(new_n11662_), .Y(new_n11663_));
  XOR2X1   g11407(.A(new_n11663_), .B(\a[56] ), .Y(new_n11664_));
  XOR2X1   g11408(.A(new_n11664_), .B(new_n11660_), .Y(new_n11665_));
  XOR2X1   g11409(.A(new_n11665_), .B(new_n11639_), .Y(new_n11666_));
  XOR2X1   g11410(.A(new_n11666_), .B(new_n11636_), .Y(new_n11667_));
  XOR2X1   g11411(.A(new_n11667_), .B(new_n11632_), .Y(new_n11668_));
  AOI22X1  g11412(.A0(new_n4880_), .A1(\b[38] ), .B0(new_n4877_), .B1(\b[37] ), .Y(new_n11669_));
  OAI21X1  g11413(.A0(new_n5291_), .A1(new_n3276_), .B0(new_n11669_), .Y(new_n11670_));
  AOI21X1  g11414(.A0(new_n4875_), .A1(new_n3275_), .B0(new_n11670_), .Y(new_n11671_));
  XOR2X1   g11415(.A(new_n11671_), .B(\a[50] ), .Y(new_n11672_));
  XOR2X1   g11416(.A(new_n11672_), .B(new_n11668_), .Y(new_n11673_));
  OR2X1    g11417(.A(new_n11522_), .B(new_n11519_), .Y(new_n11674_));
  OR2X1    g11418(.A(new_n11527_), .B(new_n11523_), .Y(new_n11675_));
  AND2X1   g11419(.A(new_n11675_), .B(new_n11674_), .Y(new_n11676_));
  XOR2X1   g11420(.A(new_n11676_), .B(new_n11673_), .Y(new_n11677_));
  AOI22X1  g11421(.A0(new_n4572_), .A1(\b[41] ), .B0(new_n4571_), .B1(\b[40] ), .Y(new_n11678_));
  OAI21X1  g11422(.A0(new_n4740_), .A1(new_n3723_), .B0(new_n11678_), .Y(new_n11679_));
  AOI21X1  g11423(.A0(new_n4375_), .A1(new_n3722_), .B0(new_n11679_), .Y(new_n11680_));
  XOR2X1   g11424(.A(new_n11680_), .B(\a[47] ), .Y(new_n11681_));
  XOR2X1   g11425(.A(new_n11681_), .B(new_n11677_), .Y(new_n11682_));
  XOR2X1   g11426(.A(new_n11682_), .B(new_n11628_), .Y(new_n11683_));
  XOR2X1   g11427(.A(new_n11683_), .B(new_n11625_), .Y(new_n11684_));
  XOR2X1   g11428(.A(new_n11684_), .B(new_n11621_), .Y(new_n11685_));
  AOI22X1  g11429(.A0(new_n3652_), .A1(\b[47] ), .B0(new_n3651_), .B1(\b[46] ), .Y(new_n11686_));
  OAI21X1  g11430(.A0(new_n3778_), .A1(new_n4674_), .B0(new_n11686_), .Y(new_n11687_));
  AOI21X1  g11431(.A0(new_n4673_), .A1(new_n3480_), .B0(new_n11687_), .Y(new_n11688_));
  XOR2X1   g11432(.A(new_n11688_), .B(\a[41] ), .Y(new_n11689_));
  XOR2X1   g11433(.A(new_n11689_), .B(new_n11685_), .Y(new_n11690_));
  INVX1    g11434(.A(new_n11690_), .Y(new_n11691_));
  NOR2X1   g11435(.A(new_n11539_), .B(new_n11536_), .Y(new_n11692_));
  INVX1    g11436(.A(new_n11544_), .Y(new_n11693_));
  AOI21X1  g11437(.A0(new_n11693_), .A1(new_n11540_), .B0(new_n11692_), .Y(new_n11694_));
  XOR2X1   g11438(.A(new_n11694_), .B(new_n11691_), .Y(new_n11695_));
  AOI22X1  g11439(.A0(new_n3204_), .A1(\b[50] ), .B0(new_n3203_), .B1(\b[49] ), .Y(new_n11696_));
  OAI21X1  g11440(.A0(new_n3321_), .A1(new_n5036_), .B0(new_n11696_), .Y(new_n11697_));
  AOI21X1  g11441(.A0(new_n5204_), .A1(new_n3080_), .B0(new_n11697_), .Y(new_n11698_));
  XOR2X1   g11442(.A(new_n11698_), .B(\a[38] ), .Y(new_n11699_));
  XOR2X1   g11443(.A(new_n11699_), .B(new_n11695_), .Y(new_n11700_));
  XOR2X1   g11444(.A(new_n11700_), .B(new_n11617_), .Y(new_n11701_));
  XOR2X1   g11445(.A(new_n11701_), .B(new_n11613_), .Y(new_n11702_));
  XOR2X1   g11446(.A(new_n11702_), .B(new_n11609_), .Y(new_n11703_));
  XOR2X1   g11447(.A(new_n11703_), .B(new_n11601_), .Y(new_n11704_));
  XOR2X1   g11448(.A(new_n11704_), .B(new_n11593_), .Y(new_n11705_));
  XOR2X1   g11449(.A(new_n11705_), .B(new_n11586_), .Y(new_n11706_));
  XOR2X1   g11450(.A(new_n11706_), .B(new_n11580_), .Y(new_n11707_));
  XOR2X1   g11451(.A(new_n11707_), .B(new_n11578_), .Y(\f[86] ));
  INVX1    g11452(.A(new_n11706_), .Y(new_n11709_));
  NOR2X1   g11453(.A(new_n11709_), .B(new_n11580_), .Y(new_n11710_));
  AOI21X1  g11454(.A0(new_n11577_), .A1(new_n11576_), .B0(new_n11707_), .Y(new_n11711_));
  OR2X1    g11455(.A(new_n11711_), .B(new_n11710_), .Y(new_n11712_));
  XOR2X1   g11456(.A(new_n11584_), .B(new_n1351_), .Y(new_n11713_));
  NOR2X1   g11457(.A(new_n11705_), .B(new_n11586_), .Y(new_n11714_));
  AOI21X1  g11458(.A0(new_n11713_), .A1(new_n11583_), .B0(new_n11714_), .Y(new_n11715_));
  NOR2X1   g11459(.A(new_n11592_), .B(new_n11590_), .Y(new_n11716_));
  INVX1    g11460(.A(new_n11716_), .Y(new_n11717_));
  INVX1    g11461(.A(new_n11593_), .Y(new_n11718_));
  OAI21X1  g11462(.A0(new_n11704_), .A1(new_n11718_), .B0(new_n11717_), .Y(new_n11719_));
  AOI22X1  g11463(.A0(new_n1814_), .A1(\b[63] ), .B0(new_n1813_), .B1(\b[62] ), .Y(new_n11720_));
  OAI21X1  g11464(.A0(new_n1812_), .A1(new_n7748_), .B0(new_n11720_), .Y(new_n11721_));
  AOI21X1  g11465(.A0(new_n7747_), .A1(new_n1617_), .B0(new_n11721_), .Y(new_n11722_));
  XOR2X1   g11466(.A(new_n11722_), .B(\a[26] ), .Y(new_n11723_));
  XOR2X1   g11467(.A(new_n11723_), .B(new_n11719_), .Y(new_n11724_));
  NOR2X1   g11468(.A(new_n11600_), .B(new_n11597_), .Y(new_n11725_));
  INVX1    g11469(.A(new_n11703_), .Y(new_n11726_));
  AOI21X1  g11470(.A0(new_n11726_), .A1(new_n11601_), .B0(new_n11725_), .Y(new_n11727_));
  AOI22X1  g11471(.A0(new_n2163_), .A1(\b[60] ), .B0(new_n2162_), .B1(\b[59] ), .Y(new_n11728_));
  OAI21X1  g11472(.A0(new_n2161_), .A1(new_n6930_), .B0(new_n11728_), .Y(new_n11729_));
  AOI21X1  g11473(.A0(new_n6951_), .A1(new_n1907_), .B0(new_n11729_), .Y(new_n11730_));
  XOR2X1   g11474(.A(new_n11730_), .B(\a[29] ), .Y(new_n11731_));
  INVX1    g11475(.A(new_n11731_), .Y(new_n11732_));
  XOR2X1   g11476(.A(new_n11732_), .B(new_n11727_), .Y(new_n11733_));
  AOI22X1  g11477(.A0(new_n2545_), .A1(\b[57] ), .B0(new_n2544_), .B1(\b[56] ), .Y(new_n11734_));
  OAI21X1  g11478(.A0(new_n2543_), .A1(new_n6523_), .B0(new_n11734_), .Y(new_n11735_));
  AOI21X1  g11479(.A0(new_n6522_), .A1(new_n2260_), .B0(new_n11735_), .Y(new_n11736_));
  XOR2X1   g11480(.A(new_n11736_), .B(\a[32] ), .Y(new_n11737_));
  NOR2X1   g11481(.A(new_n11608_), .B(new_n11605_), .Y(new_n11738_));
  INVX1    g11482(.A(new_n11702_), .Y(new_n11739_));
  AOI21X1  g11483(.A0(new_n11739_), .A1(new_n11609_), .B0(new_n11738_), .Y(new_n11740_));
  XOR2X1   g11484(.A(new_n11740_), .B(new_n11737_), .Y(new_n11741_));
  NAND2X1  g11485(.A(new_n11700_), .B(new_n11617_), .Y(new_n11742_));
  INVX1    g11486(.A(new_n11701_), .Y(new_n11743_));
  OAI21X1  g11487(.A0(new_n11743_), .A1(new_n11613_), .B0(new_n11742_), .Y(new_n11744_));
  NOR2X1   g11488(.A(new_n11694_), .B(new_n11690_), .Y(new_n11745_));
  INVX1    g11489(.A(new_n11745_), .Y(new_n11746_));
  OAI21X1  g11490(.A0(new_n11699_), .A1(new_n11695_), .B0(new_n11746_), .Y(new_n11747_));
  NOR2X1   g11491(.A(new_n11682_), .B(new_n11628_), .Y(new_n11748_));
  AOI21X1  g11492(.A0(new_n11683_), .A1(new_n11625_), .B0(new_n11748_), .Y(new_n11749_));
  INVX1    g11493(.A(new_n11749_), .Y(new_n11750_));
  OR2X1    g11494(.A(new_n11676_), .B(new_n11673_), .Y(new_n11751_));
  INVX1    g11495(.A(new_n11677_), .Y(new_n11752_));
  OAI21X1  g11496(.A0(new_n11681_), .A1(new_n11752_), .B0(new_n11751_), .Y(new_n11753_));
  AND2X1   g11497(.A(new_n11650_), .B(new_n11643_), .Y(new_n11754_));
  INVX1    g11498(.A(new_n11754_), .Y(new_n11755_));
  INVX1    g11499(.A(new_n11651_), .Y(new_n11756_));
  OAI21X1  g11500(.A0(new_n11655_), .A1(new_n11756_), .B0(new_n11755_), .Y(new_n11757_));
  NOR2X1   g11501(.A(new_n11649_), .B(new_n11645_), .Y(new_n11758_));
  AOI21X1  g11502(.A0(new_n11644_), .A1(new_n11640_), .B0(new_n11758_), .Y(new_n11759_));
  INVX1    g11503(.A(new_n11759_), .Y(new_n11760_));
  INVX1    g11504(.A(new_n11644_), .Y(new_n11761_));
  AOI22X1  g11505(.A0(new_n7818_), .A1(\b[23] ), .B0(new_n7817_), .B1(\b[24] ), .Y(new_n11762_));
  XOR2X1   g11506(.A(new_n11762_), .B(\a[23] ), .Y(new_n11763_));
  XOR2X1   g11507(.A(new_n11763_), .B(new_n11761_), .Y(new_n11764_));
  AOI22X1  g11508(.A0(new_n7192_), .A1(\b[27] ), .B0(new_n7189_), .B1(\b[26] ), .Y(new_n11765_));
  OAI21X1  g11509(.A0(new_n7627_), .A1(new_n1880_), .B0(new_n11765_), .Y(new_n11766_));
  AOI21X1  g11510(.A0(new_n7187_), .A1(new_n1879_), .B0(new_n11766_), .Y(new_n11767_));
  XOR2X1   g11511(.A(new_n11767_), .B(\a[62] ), .Y(new_n11768_));
  XOR2X1   g11512(.A(new_n11768_), .B(new_n11764_), .Y(new_n11769_));
  XOR2X1   g11513(.A(new_n11769_), .B(new_n11760_), .Y(new_n11770_));
  AOI22X1  g11514(.A0(new_n6603_), .A1(\b[30] ), .B0(new_n6600_), .B1(\b[29] ), .Y(new_n11771_));
  OAI21X1  g11515(.A0(new_n6804_), .A1(new_n2231_), .B0(new_n11771_), .Y(new_n11772_));
  AOI21X1  g11516(.A0(new_n6598_), .A1(new_n2230_), .B0(new_n11772_), .Y(new_n11773_));
  XOR2X1   g11517(.A(new_n11773_), .B(\a[59] ), .Y(new_n11774_));
  XOR2X1   g11518(.A(new_n11774_), .B(new_n11770_), .Y(new_n11775_));
  XOR2X1   g11519(.A(new_n11775_), .B(new_n11757_), .Y(new_n11776_));
  AOI22X1  g11520(.A0(new_n6438_), .A1(\b[33] ), .B0(new_n6437_), .B1(\b[32] ), .Y(new_n11777_));
  OAI21X1  g11521(.A0(new_n6436_), .A1(new_n2615_), .B0(new_n11777_), .Y(new_n11778_));
  AOI21X1  g11522(.A0(new_n6023_), .A1(new_n2614_), .B0(new_n11778_), .Y(new_n11779_));
  XOR2X1   g11523(.A(new_n11779_), .B(\a[56] ), .Y(new_n11780_));
  OR2X1    g11524(.A(new_n11659_), .B(new_n11656_), .Y(new_n11781_));
  OR2X1    g11525(.A(new_n11664_), .B(new_n11660_), .Y(new_n11782_));
  AND2X1   g11526(.A(new_n11782_), .B(new_n11781_), .Y(new_n11783_));
  XOR2X1   g11527(.A(new_n11783_), .B(new_n11780_), .Y(new_n11784_));
  XOR2X1   g11528(.A(new_n11784_), .B(new_n11776_), .Y(new_n11785_));
  AOI22X1  g11529(.A0(new_n5430_), .A1(\b[36] ), .B0(new_n5427_), .B1(\b[35] ), .Y(new_n11786_));
  OAI21X1  g11530(.A0(new_n5891_), .A1(new_n2890_), .B0(new_n11786_), .Y(new_n11787_));
  AOI21X1  g11531(.A0(new_n5425_), .A1(new_n3015_), .B0(new_n11787_), .Y(new_n11788_));
  XOR2X1   g11532(.A(new_n11788_), .B(\a[53] ), .Y(new_n11789_));
  XOR2X1   g11533(.A(new_n11789_), .B(new_n11785_), .Y(new_n11790_));
  AND2X1   g11534(.A(new_n11665_), .B(new_n11639_), .Y(new_n11791_));
  AOI21X1  g11535(.A0(new_n11666_), .A1(new_n11636_), .B0(new_n11791_), .Y(new_n11792_));
  XOR2X1   g11536(.A(new_n11792_), .B(new_n11790_), .Y(new_n11793_));
  AOI22X1  g11537(.A0(new_n4880_), .A1(\b[39] ), .B0(new_n4877_), .B1(\b[38] ), .Y(new_n11794_));
  OAI21X1  g11538(.A0(new_n5291_), .A1(new_n3413_), .B0(new_n11794_), .Y(new_n11795_));
  AOI21X1  g11539(.A0(new_n4875_), .A1(new_n3412_), .B0(new_n11795_), .Y(new_n11796_));
  XOR2X1   g11540(.A(new_n11796_), .B(\a[50] ), .Y(new_n11797_));
  XOR2X1   g11541(.A(new_n11797_), .B(new_n11793_), .Y(new_n11798_));
  AND2X1   g11542(.A(new_n11667_), .B(new_n11632_), .Y(new_n11799_));
  INVX1    g11543(.A(new_n11672_), .Y(new_n11800_));
  AOI21X1  g11544(.A0(new_n11800_), .A1(new_n11668_), .B0(new_n11799_), .Y(new_n11801_));
  XOR2X1   g11545(.A(new_n11801_), .B(new_n11798_), .Y(new_n11802_));
  AOI22X1  g11546(.A0(new_n4572_), .A1(\b[42] ), .B0(new_n4571_), .B1(\b[41] ), .Y(new_n11803_));
  OAI21X1  g11547(.A0(new_n4740_), .A1(new_n3720_), .B0(new_n11803_), .Y(new_n11804_));
  AOI21X1  g11548(.A0(new_n4375_), .A1(new_n3860_), .B0(new_n11804_), .Y(new_n11805_));
  XOR2X1   g11549(.A(new_n11805_), .B(\a[47] ), .Y(new_n11806_));
  XOR2X1   g11550(.A(new_n11806_), .B(new_n11802_), .Y(new_n11807_));
  XOR2X1   g11551(.A(new_n11807_), .B(new_n11753_), .Y(new_n11808_));
  AOI22X1  g11552(.A0(new_n4095_), .A1(\b[45] ), .B0(new_n4094_), .B1(\b[44] ), .Y(new_n11809_));
  OAI21X1  g11553(.A0(new_n4233_), .A1(new_n4339_), .B0(new_n11809_), .Y(new_n11810_));
  AOI21X1  g11554(.A0(new_n4338_), .A1(new_n3901_), .B0(new_n11810_), .Y(new_n11811_));
  XOR2X1   g11555(.A(new_n11811_), .B(\a[44] ), .Y(new_n11812_));
  XOR2X1   g11556(.A(new_n11812_), .B(new_n11808_), .Y(new_n11813_));
  XOR2X1   g11557(.A(new_n11813_), .B(new_n11750_), .Y(new_n11814_));
  AOI22X1  g11558(.A0(new_n3652_), .A1(\b[48] ), .B0(new_n3651_), .B1(\b[47] ), .Y(new_n11815_));
  OAI21X1  g11559(.A0(new_n3778_), .A1(new_n4693_), .B0(new_n11815_), .Y(new_n11816_));
  AOI21X1  g11560(.A0(new_n4692_), .A1(new_n3480_), .B0(new_n11816_), .Y(new_n11817_));
  XOR2X1   g11561(.A(new_n11817_), .B(\a[41] ), .Y(new_n11818_));
  XOR2X1   g11562(.A(new_n11818_), .B(new_n11814_), .Y(new_n11819_));
  AND2X1   g11563(.A(new_n11684_), .B(new_n11621_), .Y(new_n11820_));
  INVX1    g11564(.A(new_n11689_), .Y(new_n11821_));
  AOI21X1  g11565(.A0(new_n11821_), .A1(new_n11685_), .B0(new_n11820_), .Y(new_n11822_));
  XOR2X1   g11566(.A(new_n11822_), .B(new_n11819_), .Y(new_n11823_));
  INVX1    g11567(.A(new_n11823_), .Y(new_n11824_));
  AOI22X1  g11568(.A0(new_n3204_), .A1(\b[51] ), .B0(new_n3203_), .B1(\b[50] ), .Y(new_n11825_));
  OAI21X1  g11569(.A0(new_n3321_), .A1(new_n5237_), .B0(new_n11825_), .Y(new_n11826_));
  AOI21X1  g11570(.A0(new_n5236_), .A1(new_n3080_), .B0(new_n11826_), .Y(new_n11827_));
  XOR2X1   g11571(.A(new_n11827_), .B(\a[38] ), .Y(new_n11828_));
  AND2X1   g11572(.A(new_n11828_), .B(new_n11824_), .Y(new_n11829_));
  INVX1    g11573(.A(new_n11829_), .Y(new_n11830_));
  OAI21X1  g11574(.A0(new_n11828_), .A1(new_n11824_), .B0(new_n11747_), .Y(new_n11831_));
  OR2X1    g11575(.A(new_n11831_), .B(new_n11829_), .Y(new_n11832_));
  NOR2X1   g11576(.A(new_n11828_), .B(new_n11824_), .Y(new_n11833_));
  AOI21X1  g11577(.A0(new_n11830_), .A1(new_n11747_), .B0(new_n11833_), .Y(new_n11834_));
  AOI22X1  g11578(.A0(new_n11834_), .A1(new_n11830_), .B0(new_n11832_), .B1(new_n11747_), .Y(new_n11835_));
  AOI22X1  g11579(.A0(new_n2813_), .A1(\b[54] ), .B0(new_n2812_), .B1(\b[53] ), .Y(new_n11836_));
  OAI21X1  g11580(.A0(new_n2946_), .A1(new_n5808_), .B0(new_n11836_), .Y(new_n11837_));
  AOI21X1  g11581(.A0(new_n5807_), .A1(new_n2652_), .B0(new_n11837_), .Y(new_n11838_));
  XOR2X1   g11582(.A(new_n11838_), .B(\a[35] ), .Y(new_n11839_));
  XOR2X1   g11583(.A(new_n11839_), .B(new_n11835_), .Y(new_n11840_));
  XOR2X1   g11584(.A(new_n11840_), .B(new_n11744_), .Y(new_n11841_));
  XOR2X1   g11585(.A(new_n11841_), .B(new_n11741_), .Y(new_n11842_));
  XOR2X1   g11586(.A(new_n11842_), .B(new_n11733_), .Y(new_n11843_));
  INVX1    g11587(.A(new_n11843_), .Y(new_n11844_));
  XOR2X1   g11588(.A(new_n11844_), .B(new_n11724_), .Y(new_n11845_));
  XOR2X1   g11589(.A(new_n11845_), .B(new_n11715_), .Y(new_n11846_));
  XOR2X1   g11590(.A(new_n11846_), .B(new_n11712_), .Y(\f[87] ));
  NOR2X1   g11591(.A(new_n11845_), .B(new_n11715_), .Y(new_n11848_));
  INVX1    g11592(.A(new_n11848_), .Y(new_n11849_));
  OAI21X1  g11593(.A0(new_n11711_), .A1(new_n11710_), .B0(new_n11846_), .Y(new_n11850_));
  AND2X1   g11594(.A(new_n11850_), .B(new_n11849_), .Y(new_n11851_));
  XOR2X1   g11595(.A(new_n11722_), .B(new_n1621_), .Y(new_n11852_));
  NOR2X1   g11596(.A(new_n11843_), .B(new_n11724_), .Y(new_n11853_));
  AOI21X1  g11597(.A0(new_n11852_), .A1(new_n11719_), .B0(new_n11853_), .Y(new_n11854_));
  OAI22X1  g11598(.A0(new_n1812_), .A1(new_n7745_), .B0(new_n1620_), .B1(new_n7772_), .Y(new_n11855_));
  AOI21X1  g11599(.A0(new_n7775_), .A1(new_n1617_), .B0(new_n11855_), .Y(new_n11856_));
  XOR2X1   g11600(.A(new_n11856_), .B(\a[26] ), .Y(new_n11857_));
  INVX1    g11601(.A(new_n11733_), .Y(new_n11858_));
  NOR2X1   g11602(.A(new_n11731_), .B(new_n11727_), .Y(new_n11859_));
  AOI21X1  g11603(.A0(new_n11842_), .A1(new_n11858_), .B0(new_n11859_), .Y(new_n11860_));
  NOR2X1   g11604(.A(new_n11857_), .B(new_n11860_), .Y(new_n11861_));
  OR2X1    g11605(.A(new_n11861_), .B(new_n11857_), .Y(new_n11862_));
  AOI22X1  g11606(.A0(new_n2163_), .A1(\b[61] ), .B0(new_n2162_), .B1(\b[60] ), .Y(new_n11863_));
  OAI21X1  g11607(.A0(new_n2161_), .A1(new_n7339_), .B0(new_n11863_), .Y(new_n11864_));
  AOI21X1  g11608(.A0(new_n7338_), .A1(new_n1907_), .B0(new_n11864_), .Y(new_n11865_));
  XOR2X1   g11609(.A(new_n11865_), .B(\a[29] ), .Y(new_n11866_));
  NOR2X1   g11610(.A(new_n11740_), .B(new_n11737_), .Y(new_n11867_));
  AOI21X1  g11611(.A0(new_n11841_), .A1(new_n11741_), .B0(new_n11867_), .Y(new_n11868_));
  XOR2X1   g11612(.A(new_n11868_), .B(new_n11866_), .Y(new_n11869_));
  INVX1    g11613(.A(new_n11869_), .Y(new_n11870_));
  NOR2X1   g11614(.A(new_n11839_), .B(new_n11835_), .Y(new_n11871_));
  AOI21X1  g11615(.A0(new_n11840_), .A1(new_n11744_), .B0(new_n11871_), .Y(new_n11872_));
  OAI22X1  g11616(.A0(new_n2263_), .A1(new_n6930_), .B0(new_n2262_), .B1(new_n6933_), .Y(new_n11873_));
  AOI21X1  g11617(.A0(new_n2402_), .A1(\b[56] ), .B0(new_n11873_), .Y(new_n11874_));
  OAI21X1  g11618(.A0(new_n8540_), .A1(new_n2400_), .B0(new_n11874_), .Y(new_n11875_));
  XOR2X1   g11619(.A(new_n11875_), .B(new_n2258_), .Y(new_n11876_));
  XOR2X1   g11620(.A(new_n11876_), .B(new_n11872_), .Y(new_n11877_));
  XOR2X1   g11621(.A(new_n11796_), .B(new_n4873_), .Y(new_n11878_));
  NOR2X1   g11622(.A(new_n11801_), .B(new_n11798_), .Y(new_n11879_));
  AOI21X1  g11623(.A0(new_n11878_), .A1(new_n11793_), .B0(new_n11879_), .Y(new_n11880_));
  INVX1    g11624(.A(new_n11880_), .Y(new_n11881_));
  AOI22X1  g11625(.A0(new_n4880_), .A1(\b[40] ), .B0(new_n4877_), .B1(\b[39] ), .Y(new_n11882_));
  OAI21X1  g11626(.A0(new_n5291_), .A1(new_n3575_), .B0(new_n11882_), .Y(new_n11883_));
  AOI21X1  g11627(.A0(new_n4875_), .A1(new_n3574_), .B0(new_n11883_), .Y(new_n11884_));
  XOR2X1   g11628(.A(new_n11884_), .B(\a[50] ), .Y(new_n11885_));
  XOR2X1   g11629(.A(new_n11788_), .B(new_n5423_), .Y(new_n11886_));
  AND2X1   g11630(.A(new_n11886_), .B(new_n11785_), .Y(new_n11887_));
  NOR2X1   g11631(.A(new_n11792_), .B(new_n11790_), .Y(new_n11888_));
  NOR2X1   g11632(.A(new_n11888_), .B(new_n11887_), .Y(new_n11889_));
  INVX1    g11633(.A(new_n11764_), .Y(new_n11890_));
  NOR2X1   g11634(.A(new_n11768_), .B(new_n11890_), .Y(new_n11891_));
  NOR2X1   g11635(.A(new_n11769_), .B(new_n11759_), .Y(new_n11892_));
  NOR2X1   g11636(.A(new_n11892_), .B(new_n11891_), .Y(new_n11893_));
  INVX1    g11637(.A(new_n11893_), .Y(new_n11894_));
  AOI22X1  g11638(.A0(new_n7818_), .A1(\b[24] ), .B0(new_n7817_), .B1(\b[25] ), .Y(new_n11895_));
  NOR2X1   g11639(.A(new_n11762_), .B(\a[23] ), .Y(new_n11896_));
  AOI21X1  g11640(.A0(new_n11763_), .A1(new_n11761_), .B0(new_n11896_), .Y(new_n11897_));
  XOR2X1   g11641(.A(new_n11897_), .B(new_n11895_), .Y(new_n11898_));
  AOI22X1  g11642(.A0(new_n7192_), .A1(\b[28] ), .B0(new_n7189_), .B1(\b[27] ), .Y(new_n11899_));
  OAI21X1  g11643(.A0(new_n7627_), .A1(new_n1877_), .B0(new_n11899_), .Y(new_n11900_));
  AOI21X1  g11644(.A0(new_n7187_), .A1(new_n2004_), .B0(new_n11900_), .Y(new_n11901_));
  XOR2X1   g11645(.A(new_n11901_), .B(\a[62] ), .Y(new_n11902_));
  XOR2X1   g11646(.A(new_n11902_), .B(new_n11898_), .Y(new_n11903_));
  XOR2X1   g11647(.A(new_n11903_), .B(new_n11894_), .Y(new_n11904_));
  AOI22X1  g11648(.A0(new_n6603_), .A1(\b[31] ), .B0(new_n6600_), .B1(\b[30] ), .Y(new_n11905_));
  OAI21X1  g11649(.A0(new_n6804_), .A1(new_n2359_), .B0(new_n11905_), .Y(new_n11906_));
  AOI21X1  g11650(.A0(new_n6598_), .A1(new_n2358_), .B0(new_n11906_), .Y(new_n11907_));
  XOR2X1   g11651(.A(new_n11907_), .B(\a[59] ), .Y(new_n11908_));
  XOR2X1   g11652(.A(new_n11908_), .B(new_n11904_), .Y(new_n11909_));
  NOR2X1   g11653(.A(new_n11774_), .B(new_n11770_), .Y(new_n11910_));
  AOI21X1  g11654(.A0(new_n11775_), .A1(new_n11757_), .B0(new_n11910_), .Y(new_n11911_));
  XOR2X1   g11655(.A(new_n11911_), .B(new_n11909_), .Y(new_n11912_));
  AOI22X1  g11656(.A0(new_n6438_), .A1(\b[34] ), .B0(new_n6437_), .B1(\b[33] ), .Y(new_n11913_));
  OAI21X1  g11657(.A0(new_n6436_), .A1(new_n2612_), .B0(new_n11913_), .Y(new_n11914_));
  AOI21X1  g11658(.A0(new_n6023_), .A1(new_n2759_), .B0(new_n11914_), .Y(new_n11915_));
  XOR2X1   g11659(.A(new_n11915_), .B(\a[56] ), .Y(new_n11916_));
  XOR2X1   g11660(.A(new_n11916_), .B(new_n11912_), .Y(new_n11917_));
  INVX1    g11661(.A(new_n11917_), .Y(new_n11918_));
  AOI21X1  g11662(.A0(new_n11782_), .A1(new_n11781_), .B0(new_n11780_), .Y(new_n11919_));
  AOI21X1  g11663(.A0(new_n11784_), .A1(new_n11776_), .B0(new_n11919_), .Y(new_n11920_));
  XOR2X1   g11664(.A(new_n11920_), .B(new_n11918_), .Y(new_n11921_));
  AOI22X1  g11665(.A0(new_n5430_), .A1(\b[37] ), .B0(new_n5427_), .B1(\b[36] ), .Y(new_n11922_));
  OAI21X1  g11666(.A0(new_n5891_), .A1(new_n3156_), .B0(new_n11922_), .Y(new_n11923_));
  AOI21X1  g11667(.A0(new_n5425_), .A1(new_n3155_), .B0(new_n11923_), .Y(new_n11924_));
  XOR2X1   g11668(.A(new_n11924_), .B(\a[53] ), .Y(new_n11925_));
  XOR2X1   g11669(.A(new_n11925_), .B(new_n11921_), .Y(new_n11926_));
  XOR2X1   g11670(.A(new_n11926_), .B(new_n11889_), .Y(new_n11927_));
  XOR2X1   g11671(.A(new_n11927_), .B(new_n11885_), .Y(new_n11928_));
  XOR2X1   g11672(.A(new_n11928_), .B(new_n11881_), .Y(new_n11929_));
  AOI22X1  g11673(.A0(new_n4572_), .A1(\b[43] ), .B0(new_n4571_), .B1(\b[42] ), .Y(new_n11930_));
  OAI21X1  g11674(.A0(new_n4740_), .A1(new_n4015_), .B0(new_n11930_), .Y(new_n11931_));
  AOI21X1  g11675(.A0(new_n4375_), .A1(new_n4014_), .B0(new_n11931_), .Y(new_n11932_));
  XOR2X1   g11676(.A(new_n11932_), .B(\a[47] ), .Y(new_n11933_));
  XOR2X1   g11677(.A(new_n11933_), .B(new_n11929_), .Y(new_n11934_));
  INVX1    g11678(.A(new_n11802_), .Y(new_n11935_));
  NOR2X1   g11679(.A(new_n11806_), .B(new_n11935_), .Y(new_n11936_));
  INVX1    g11680(.A(new_n11807_), .Y(new_n11937_));
  AOI21X1  g11681(.A0(new_n11937_), .A1(new_n11753_), .B0(new_n11936_), .Y(new_n11938_));
  XOR2X1   g11682(.A(new_n11938_), .B(new_n11934_), .Y(new_n11939_));
  AOI22X1  g11683(.A0(new_n4095_), .A1(\b[46] ), .B0(new_n4094_), .B1(\b[45] ), .Y(new_n11940_));
  OAI21X1  g11684(.A0(new_n4233_), .A1(new_n4336_), .B0(new_n11940_), .Y(new_n11941_));
  AOI21X1  g11685(.A0(new_n4509_), .A1(new_n3901_), .B0(new_n11941_), .Y(new_n11942_));
  XOR2X1   g11686(.A(new_n11942_), .B(\a[44] ), .Y(new_n11943_));
  XOR2X1   g11687(.A(new_n11943_), .B(new_n11939_), .Y(new_n11944_));
  NOR2X1   g11688(.A(new_n11812_), .B(new_n11808_), .Y(new_n11945_));
  AOI21X1  g11689(.A0(new_n11813_), .A1(new_n11750_), .B0(new_n11945_), .Y(new_n11946_));
  XOR2X1   g11690(.A(new_n11946_), .B(new_n11944_), .Y(new_n11947_));
  AOI22X1  g11691(.A0(new_n3652_), .A1(\b[49] ), .B0(new_n3651_), .B1(\b[48] ), .Y(new_n11948_));
  OAI21X1  g11692(.A0(new_n3778_), .A1(new_n5039_), .B0(new_n11948_), .Y(new_n11949_));
  AOI21X1  g11693(.A0(new_n5038_), .A1(new_n3480_), .B0(new_n11949_), .Y(new_n11950_));
  XOR2X1   g11694(.A(new_n11950_), .B(\a[41] ), .Y(new_n11951_));
  XOR2X1   g11695(.A(new_n11951_), .B(new_n11947_), .Y(new_n11952_));
  INVX1    g11696(.A(new_n11818_), .Y(new_n11953_));
  NOR2X1   g11697(.A(new_n11822_), .B(new_n11819_), .Y(new_n11954_));
  AOI21X1  g11698(.A0(new_n11953_), .A1(new_n11814_), .B0(new_n11954_), .Y(new_n11955_));
  XOR2X1   g11699(.A(new_n11955_), .B(new_n11952_), .Y(new_n11956_));
  AOI22X1  g11700(.A0(new_n3204_), .A1(\b[52] ), .B0(new_n3203_), .B1(\b[51] ), .Y(new_n11957_));
  OAI21X1  g11701(.A0(new_n3321_), .A1(new_n5234_), .B0(new_n11957_), .Y(new_n11958_));
  AOI21X1  g11702(.A0(new_n5590_), .A1(new_n3080_), .B0(new_n11958_), .Y(new_n11959_));
  XOR2X1   g11703(.A(new_n11959_), .B(\a[38] ), .Y(new_n11960_));
  XOR2X1   g11704(.A(new_n11960_), .B(new_n11956_), .Y(new_n11961_));
  INVX1    g11705(.A(new_n11961_), .Y(new_n11962_));
  XOR2X1   g11706(.A(new_n11962_), .B(new_n11834_), .Y(new_n11963_));
  AOI22X1  g11707(.A0(new_n2813_), .A1(\b[55] ), .B0(new_n2812_), .B1(\b[54] ), .Y(new_n11964_));
  OAI21X1  g11708(.A0(new_n2946_), .A1(new_n6151_), .B0(new_n11964_), .Y(new_n11965_));
  AOI21X1  g11709(.A0(new_n6150_), .A1(new_n2652_), .B0(new_n11965_), .Y(new_n11966_));
  XOR2X1   g11710(.A(new_n11966_), .B(\a[35] ), .Y(new_n11967_));
  XOR2X1   g11711(.A(new_n11967_), .B(new_n11963_), .Y(new_n11968_));
  XOR2X1   g11712(.A(new_n11968_), .B(new_n11877_), .Y(new_n11969_));
  XOR2X1   g11713(.A(new_n11969_), .B(new_n11870_), .Y(new_n11970_));
  OR2X1    g11714(.A(new_n11861_), .B(new_n11860_), .Y(new_n11971_));
  AOI21X1  g11715(.A0(new_n11862_), .A1(new_n11971_), .B0(new_n11970_), .Y(new_n11972_));
  AND2X1   g11716(.A(new_n11971_), .B(new_n11970_), .Y(new_n11973_));
  AOI21X1  g11717(.A0(new_n11973_), .A1(new_n11862_), .B0(new_n11972_), .Y(new_n11974_));
  XOR2X1   g11718(.A(new_n11974_), .B(new_n11854_), .Y(new_n11975_));
  XOR2X1   g11719(.A(new_n11975_), .B(new_n11851_), .Y(\f[88] ));
  AND2X1   g11720(.A(new_n11973_), .B(new_n11862_), .Y(new_n11977_));
  NOR3X1   g11721(.A(new_n11977_), .B(new_n11972_), .C(new_n11854_), .Y(new_n11978_));
  AOI21X1  g11722(.A0(new_n11850_), .A1(new_n11849_), .B0(new_n11975_), .Y(new_n11979_));
  OR2X1    g11723(.A(new_n11979_), .B(new_n11978_), .Y(new_n11980_));
  OR2X1    g11724(.A(new_n11972_), .B(new_n11861_), .Y(new_n11981_));
  NOR2X1   g11725(.A(new_n11868_), .B(new_n11866_), .Y(new_n11982_));
  AOI21X1  g11726(.A0(new_n11969_), .A1(new_n11869_), .B0(new_n11982_), .Y(new_n11983_));
  AOI22X1  g11727(.A0(new_n7774_), .A1(new_n1617_), .B0(new_n1725_), .B1(\b[63] ), .Y(new_n11984_));
  XOR2X1   g11728(.A(new_n11984_), .B(\a[26] ), .Y(new_n11985_));
  XOR2X1   g11729(.A(new_n11985_), .B(new_n11983_), .Y(new_n11986_));
  AOI22X1  g11730(.A0(new_n2163_), .A1(\b[62] ), .B0(new_n2162_), .B1(\b[61] ), .Y(new_n11987_));
  OAI21X1  g11731(.A0(new_n2161_), .A1(new_n7559_), .B0(new_n11987_), .Y(new_n11988_));
  AOI21X1  g11732(.A0(new_n7558_), .A1(new_n1907_), .B0(new_n11988_), .Y(new_n11989_));
  XOR2X1   g11733(.A(new_n11989_), .B(\a[29] ), .Y(new_n11990_));
  INVX1    g11734(.A(new_n11990_), .Y(new_n11991_));
  NOR2X1   g11735(.A(new_n11876_), .B(new_n11872_), .Y(new_n11992_));
  AOI21X1  g11736(.A0(new_n11968_), .A1(new_n11877_), .B0(new_n11992_), .Y(new_n11993_));
  XOR2X1   g11737(.A(new_n11993_), .B(new_n11991_), .Y(new_n11994_));
  AOI22X1  g11738(.A0(new_n2545_), .A1(\b[59] ), .B0(new_n2544_), .B1(\b[58] ), .Y(new_n11995_));
  OAI21X1  g11739(.A0(new_n2543_), .A1(new_n6933_), .B0(new_n11995_), .Y(new_n11996_));
  AOI21X1  g11740(.A0(new_n6932_), .A1(new_n2260_), .B0(new_n11996_), .Y(new_n11997_));
  XOR2X1   g11741(.A(new_n11997_), .B(\a[32] ), .Y(new_n11998_));
  OR2X1    g11742(.A(new_n11967_), .B(new_n11963_), .Y(new_n11999_));
  OR2X1    g11743(.A(new_n11961_), .B(new_n11834_), .Y(new_n12000_));
  AND2X1   g11744(.A(new_n12000_), .B(new_n11999_), .Y(new_n12001_));
  XOR2X1   g11745(.A(new_n12001_), .B(new_n11998_), .Y(new_n12002_));
  AOI22X1  g11746(.A0(new_n2813_), .A1(\b[56] ), .B0(new_n2812_), .B1(\b[55] ), .Y(new_n12003_));
  OAI21X1  g11747(.A0(new_n2946_), .A1(new_n6148_), .B0(new_n12003_), .Y(new_n12004_));
  AOI21X1  g11748(.A0(new_n6342_), .A1(new_n2652_), .B0(new_n12004_), .Y(new_n12005_));
  XOR2X1   g11749(.A(new_n12005_), .B(\a[35] ), .Y(new_n12006_));
  AND2X1   g11750(.A(new_n11955_), .B(new_n11952_), .Y(new_n12007_));
  OR2X1    g11751(.A(new_n11955_), .B(new_n11952_), .Y(new_n12008_));
  OAI21X1  g11752(.A0(new_n11960_), .A1(new_n12007_), .B0(new_n12008_), .Y(new_n12009_));
  AOI22X1  g11753(.A0(new_n3204_), .A1(\b[53] ), .B0(new_n3203_), .B1(\b[52] ), .Y(new_n12010_));
  OAI21X1  g11754(.A0(new_n3321_), .A1(new_n5787_), .B0(new_n12010_), .Y(new_n12011_));
  AOI21X1  g11755(.A0(new_n5786_), .A1(new_n3080_), .B0(new_n12011_), .Y(new_n12012_));
  XOR2X1   g11756(.A(new_n12012_), .B(\a[38] ), .Y(new_n12013_));
  NOR2X1   g11757(.A(new_n11946_), .B(new_n11944_), .Y(new_n12014_));
  INVX1    g11758(.A(new_n12014_), .Y(new_n12015_));
  INVX1    g11759(.A(new_n11947_), .Y(new_n12016_));
  OAI21X1  g11760(.A0(new_n11951_), .A1(new_n12016_), .B0(new_n12015_), .Y(new_n12017_));
  INVX1    g11761(.A(new_n12017_), .Y(new_n12018_));
  AND2X1   g11762(.A(new_n11928_), .B(new_n11881_), .Y(new_n12019_));
  INVX1    g11763(.A(new_n12019_), .Y(new_n12020_));
  INVX1    g11764(.A(new_n11929_), .Y(new_n12021_));
  OAI21X1  g11765(.A0(new_n11933_), .A1(new_n12021_), .B0(new_n12020_), .Y(new_n12022_));
  AOI22X1  g11766(.A0(new_n4572_), .A1(\b[44] ), .B0(new_n4571_), .B1(\b[43] ), .Y(new_n12023_));
  OAI21X1  g11767(.A0(new_n4740_), .A1(new_n4012_), .B0(new_n12023_), .Y(new_n12024_));
  AOI21X1  g11768(.A0(new_n4375_), .A1(new_n4178_), .B0(new_n12024_), .Y(new_n12025_));
  XOR2X1   g11769(.A(new_n12025_), .B(new_n4568_), .Y(new_n12026_));
  OAI21X1  g11770(.A0(new_n11888_), .A1(new_n11887_), .B0(new_n11926_), .Y(new_n12027_));
  OR2X1    g11771(.A(new_n11927_), .B(new_n11885_), .Y(new_n12028_));
  AND2X1   g11772(.A(new_n12028_), .B(new_n12027_), .Y(new_n12029_));
  NOR2X1   g11773(.A(new_n11911_), .B(new_n11909_), .Y(new_n12030_));
  INVX1    g11774(.A(new_n12030_), .Y(new_n12031_));
  INVX1    g11775(.A(new_n11912_), .Y(new_n12032_));
  OAI21X1  g11776(.A0(new_n11916_), .A1(new_n12032_), .B0(new_n12031_), .Y(new_n12033_));
  AOI22X1  g11777(.A0(new_n6438_), .A1(\b[35] ), .B0(new_n6437_), .B1(\b[34] ), .Y(new_n12034_));
  OAI21X1  g11778(.A0(new_n6436_), .A1(new_n2893_), .B0(new_n12034_), .Y(new_n12035_));
  AOI21X1  g11779(.A0(new_n6023_), .A1(new_n2892_), .B0(new_n12035_), .Y(new_n12036_));
  XOR2X1   g11780(.A(new_n12036_), .B(new_n6019_), .Y(new_n12037_));
  OAI21X1  g11781(.A0(new_n11892_), .A1(new_n11891_), .B0(new_n11903_), .Y(new_n12038_));
  NOR3X1   g11782(.A(new_n11903_), .B(new_n11892_), .C(new_n11891_), .Y(new_n12039_));
  OAI21X1  g11783(.A0(new_n11908_), .A1(new_n12039_), .B0(new_n12038_), .Y(new_n12040_));
  AOI22X1  g11784(.A0(new_n6603_), .A1(\b[32] ), .B0(new_n6600_), .B1(\b[31] ), .Y(new_n12041_));
  OAI21X1  g11785(.A0(new_n6804_), .A1(new_n2356_), .B0(new_n12041_), .Y(new_n12042_));
  AOI21X1  g11786(.A0(new_n6598_), .A1(new_n2495_), .B0(new_n12042_), .Y(new_n12043_));
  XOR2X1   g11787(.A(new_n12043_), .B(new_n6596_), .Y(new_n12044_));
  INVX1    g11788(.A(new_n11895_), .Y(new_n12045_));
  OR2X1    g11789(.A(new_n11897_), .B(new_n12045_), .Y(new_n12046_));
  OAI21X1  g11790(.A0(new_n11902_), .A1(new_n11898_), .B0(new_n12046_), .Y(new_n12047_));
  AOI22X1  g11791(.A0(new_n7818_), .A1(\b[25] ), .B0(new_n7817_), .B1(\b[26] ), .Y(new_n12048_));
  XOR2X1   g11792(.A(new_n12048_), .B(new_n11895_), .Y(new_n12049_));
  AOI22X1  g11793(.A0(new_n7192_), .A1(\b[29] ), .B0(new_n7189_), .B1(\b[28] ), .Y(new_n12050_));
  OAI21X1  g11794(.A0(new_n7627_), .A1(new_n2126_), .B0(new_n12050_), .Y(new_n12051_));
  AOI21X1  g11795(.A0(new_n7187_), .A1(new_n2125_), .B0(new_n12051_), .Y(new_n12052_));
  XOR2X1   g11796(.A(new_n12052_), .B(\a[62] ), .Y(new_n12053_));
  XOR2X1   g11797(.A(new_n12053_), .B(new_n12049_), .Y(new_n12054_));
  XOR2X1   g11798(.A(new_n12054_), .B(new_n12047_), .Y(new_n12055_));
  XOR2X1   g11799(.A(new_n12055_), .B(new_n12044_), .Y(new_n12056_));
  XOR2X1   g11800(.A(new_n12056_), .B(new_n12040_), .Y(new_n12057_));
  XOR2X1   g11801(.A(new_n12057_), .B(new_n12037_), .Y(new_n12058_));
  XOR2X1   g11802(.A(new_n12058_), .B(new_n12033_), .Y(new_n12059_));
  AOI22X1  g11803(.A0(new_n5430_), .A1(\b[38] ), .B0(new_n5427_), .B1(\b[37] ), .Y(new_n12060_));
  OAI21X1  g11804(.A0(new_n5891_), .A1(new_n3276_), .B0(new_n12060_), .Y(new_n12061_));
  AOI21X1  g11805(.A0(new_n5425_), .A1(new_n3275_), .B0(new_n12061_), .Y(new_n12062_));
  XOR2X1   g11806(.A(new_n12062_), .B(\a[53] ), .Y(new_n12063_));
  XOR2X1   g11807(.A(new_n12063_), .B(new_n12059_), .Y(new_n12064_));
  OR2X1    g11808(.A(new_n11920_), .B(new_n11917_), .Y(new_n12065_));
  OR2X1    g11809(.A(new_n11925_), .B(new_n11921_), .Y(new_n12066_));
  AND2X1   g11810(.A(new_n12066_), .B(new_n12065_), .Y(new_n12067_));
  XOR2X1   g11811(.A(new_n12067_), .B(new_n12064_), .Y(new_n12068_));
  AOI22X1  g11812(.A0(new_n4880_), .A1(\b[41] ), .B0(new_n4877_), .B1(\b[40] ), .Y(new_n12069_));
  OAI21X1  g11813(.A0(new_n5291_), .A1(new_n3723_), .B0(new_n12069_), .Y(new_n12070_));
  AOI21X1  g11814(.A0(new_n4875_), .A1(new_n3722_), .B0(new_n12070_), .Y(new_n12071_));
  XOR2X1   g11815(.A(new_n12071_), .B(\a[50] ), .Y(new_n12072_));
  XOR2X1   g11816(.A(new_n12072_), .B(new_n12068_), .Y(new_n12073_));
  XOR2X1   g11817(.A(new_n12073_), .B(new_n12029_), .Y(new_n12074_));
  XOR2X1   g11818(.A(new_n12074_), .B(new_n12026_), .Y(new_n12075_));
  XOR2X1   g11819(.A(new_n12075_), .B(new_n12022_), .Y(new_n12076_));
  AOI22X1  g11820(.A0(new_n4095_), .A1(\b[47] ), .B0(new_n4094_), .B1(\b[46] ), .Y(new_n12077_));
  OAI21X1  g11821(.A0(new_n4233_), .A1(new_n4674_), .B0(new_n12077_), .Y(new_n12078_));
  AOI21X1  g11822(.A0(new_n4673_), .A1(new_n3901_), .B0(new_n12078_), .Y(new_n12079_));
  XOR2X1   g11823(.A(new_n12079_), .B(\a[44] ), .Y(new_n12080_));
  XOR2X1   g11824(.A(new_n12080_), .B(new_n12076_), .Y(new_n12081_));
  INVX1    g11825(.A(new_n12081_), .Y(new_n12082_));
  NOR2X1   g11826(.A(new_n11938_), .B(new_n11934_), .Y(new_n12083_));
  INVX1    g11827(.A(new_n11943_), .Y(new_n12084_));
  AOI21X1  g11828(.A0(new_n12084_), .A1(new_n11939_), .B0(new_n12083_), .Y(new_n12085_));
  XOR2X1   g11829(.A(new_n12085_), .B(new_n12082_), .Y(new_n12086_));
  AOI22X1  g11830(.A0(new_n3652_), .A1(\b[50] ), .B0(new_n3651_), .B1(\b[49] ), .Y(new_n12087_));
  OAI21X1  g11831(.A0(new_n3778_), .A1(new_n5036_), .B0(new_n12087_), .Y(new_n12088_));
  AOI21X1  g11832(.A0(new_n5204_), .A1(new_n3480_), .B0(new_n12088_), .Y(new_n12089_));
  XOR2X1   g11833(.A(new_n12089_), .B(\a[41] ), .Y(new_n12090_));
  XOR2X1   g11834(.A(new_n12090_), .B(new_n12086_), .Y(new_n12091_));
  XOR2X1   g11835(.A(new_n12091_), .B(new_n12018_), .Y(new_n12092_));
  XOR2X1   g11836(.A(new_n12092_), .B(new_n12013_), .Y(new_n12093_));
  XOR2X1   g11837(.A(new_n12093_), .B(new_n12009_), .Y(new_n12094_));
  XOR2X1   g11838(.A(new_n12094_), .B(new_n12006_), .Y(new_n12095_));
  XOR2X1   g11839(.A(new_n12095_), .B(new_n12002_), .Y(new_n12096_));
  XOR2X1   g11840(.A(new_n12096_), .B(new_n11994_), .Y(new_n12097_));
  XOR2X1   g11841(.A(new_n12097_), .B(new_n11986_), .Y(new_n12098_));
  XOR2X1   g11842(.A(new_n12098_), .B(new_n11981_), .Y(new_n12099_));
  XOR2X1   g11843(.A(new_n12099_), .B(new_n11980_), .Y(\f[89] ));
  NOR2X1   g11844(.A(new_n11985_), .B(new_n11983_), .Y(new_n12101_));
  AOI21X1  g11845(.A0(new_n12097_), .A1(new_n11986_), .B0(new_n12101_), .Y(new_n12102_));
  NOR2X1   g11846(.A(new_n11993_), .B(new_n11990_), .Y(new_n12103_));
  INVX1    g11847(.A(new_n12103_), .Y(new_n12104_));
  OAI21X1  g11848(.A0(new_n12096_), .A1(new_n11994_), .B0(new_n12104_), .Y(new_n12105_));
  AOI22X1  g11849(.A0(new_n2163_), .A1(\b[63] ), .B0(new_n2162_), .B1(\b[62] ), .Y(new_n12106_));
  OAI21X1  g11850(.A0(new_n2161_), .A1(new_n7748_), .B0(new_n12106_), .Y(new_n12107_));
  AOI21X1  g11851(.A0(new_n7747_), .A1(new_n1907_), .B0(new_n12107_), .Y(new_n12108_));
  XOR2X1   g11852(.A(new_n12108_), .B(\a[29] ), .Y(new_n12109_));
  XOR2X1   g11853(.A(new_n12109_), .B(new_n12105_), .Y(new_n12110_));
  AND2X1   g11854(.A(new_n12091_), .B(new_n12017_), .Y(new_n12111_));
  INVX1    g11855(.A(new_n12111_), .Y(new_n12112_));
  OAI21X1  g11856(.A0(new_n12092_), .A1(new_n12013_), .B0(new_n12112_), .Y(new_n12113_));
  NOR2X1   g11857(.A(new_n12085_), .B(new_n12081_), .Y(new_n12114_));
  INVX1    g11858(.A(new_n12114_), .Y(new_n12115_));
  OAI21X1  g11859(.A0(new_n12090_), .A1(new_n12086_), .B0(new_n12115_), .Y(new_n12116_));
  NOR2X1   g11860(.A(new_n12073_), .B(new_n12029_), .Y(new_n12117_));
  AOI21X1  g11861(.A0(new_n12074_), .A1(new_n12026_), .B0(new_n12117_), .Y(new_n12118_));
  INVX1    g11862(.A(new_n12118_), .Y(new_n12119_));
  OR2X1    g11863(.A(new_n12067_), .B(new_n12064_), .Y(new_n12120_));
  INVX1    g11864(.A(new_n12068_), .Y(new_n12121_));
  OAI21X1  g11865(.A0(new_n12072_), .A1(new_n12121_), .B0(new_n12120_), .Y(new_n12122_));
  AOI22X1  g11866(.A0(new_n6603_), .A1(\b[33] ), .B0(new_n6600_), .B1(\b[32] ), .Y(new_n12123_));
  OAI21X1  g11867(.A0(new_n6804_), .A1(new_n2615_), .B0(new_n12123_), .Y(new_n12124_));
  AOI21X1  g11868(.A0(new_n6598_), .A1(new_n2614_), .B0(new_n12124_), .Y(new_n12125_));
  XOR2X1   g11869(.A(new_n12125_), .B(\a[59] ), .Y(new_n12126_));
  AND2X1   g11870(.A(new_n12054_), .B(new_n12047_), .Y(new_n12127_));
  AOI21X1  g11871(.A0(new_n12055_), .A1(new_n12044_), .B0(new_n12127_), .Y(new_n12128_));
  XOR2X1   g11872(.A(new_n12128_), .B(new_n12126_), .Y(new_n12129_));
  INVX1    g11873(.A(new_n12129_), .Y(new_n12130_));
  NOR2X1   g11874(.A(new_n12053_), .B(new_n12049_), .Y(new_n12131_));
  AOI21X1  g11875(.A0(new_n12048_), .A1(new_n12045_), .B0(new_n12131_), .Y(new_n12132_));
  INVX1    g11876(.A(new_n12132_), .Y(new_n12133_));
  INVX1    g11877(.A(new_n12048_), .Y(new_n12134_));
  AOI22X1  g11878(.A0(new_n7818_), .A1(\b[26] ), .B0(new_n7817_), .B1(\b[27] ), .Y(new_n12135_));
  XOR2X1   g11879(.A(new_n12135_), .B(\a[26] ), .Y(new_n12136_));
  XOR2X1   g11880(.A(new_n12136_), .B(new_n12134_), .Y(new_n12137_));
  XOR2X1   g11881(.A(new_n12137_), .B(new_n12133_), .Y(new_n12138_));
  AOI22X1  g11882(.A0(new_n7192_), .A1(\b[30] ), .B0(new_n7189_), .B1(\b[29] ), .Y(new_n12139_));
  OAI21X1  g11883(.A0(new_n7627_), .A1(new_n2231_), .B0(new_n12139_), .Y(new_n12140_));
  AOI21X1  g11884(.A0(new_n7187_), .A1(new_n2230_), .B0(new_n12140_), .Y(new_n12141_));
  XOR2X1   g11885(.A(new_n12141_), .B(\a[62] ), .Y(new_n12142_));
  XOR2X1   g11886(.A(new_n12142_), .B(new_n12138_), .Y(new_n12143_));
  XOR2X1   g11887(.A(new_n12143_), .B(new_n12130_), .Y(new_n12144_));
  AOI22X1  g11888(.A0(new_n6438_), .A1(\b[36] ), .B0(new_n6437_), .B1(\b[35] ), .Y(new_n12145_));
  OAI21X1  g11889(.A0(new_n6436_), .A1(new_n2890_), .B0(new_n12145_), .Y(new_n12146_));
  AOI21X1  g11890(.A0(new_n6023_), .A1(new_n3015_), .B0(new_n12146_), .Y(new_n12147_));
  XOR2X1   g11891(.A(new_n12147_), .B(\a[56] ), .Y(new_n12148_));
  XOR2X1   g11892(.A(new_n12148_), .B(new_n12144_), .Y(new_n12149_));
  AND2X1   g11893(.A(new_n12056_), .B(new_n12040_), .Y(new_n12150_));
  AOI21X1  g11894(.A0(new_n12057_), .A1(new_n12037_), .B0(new_n12150_), .Y(new_n12151_));
  XOR2X1   g11895(.A(new_n12151_), .B(new_n12149_), .Y(new_n12152_));
  AOI22X1  g11896(.A0(new_n5430_), .A1(\b[39] ), .B0(new_n5427_), .B1(\b[38] ), .Y(new_n12153_));
  OAI21X1  g11897(.A0(new_n5891_), .A1(new_n3413_), .B0(new_n12153_), .Y(new_n12154_));
  AOI21X1  g11898(.A0(new_n5425_), .A1(new_n3412_), .B0(new_n12154_), .Y(new_n12155_));
  XOR2X1   g11899(.A(new_n12155_), .B(\a[53] ), .Y(new_n12156_));
  XOR2X1   g11900(.A(new_n12156_), .B(new_n12152_), .Y(new_n12157_));
  AND2X1   g11901(.A(new_n12058_), .B(new_n12033_), .Y(new_n12158_));
  INVX1    g11902(.A(new_n12063_), .Y(new_n12159_));
  AOI21X1  g11903(.A0(new_n12159_), .A1(new_n12059_), .B0(new_n12158_), .Y(new_n12160_));
  XOR2X1   g11904(.A(new_n12160_), .B(new_n12157_), .Y(new_n12161_));
  AOI22X1  g11905(.A0(new_n4880_), .A1(\b[42] ), .B0(new_n4877_), .B1(\b[41] ), .Y(new_n12162_));
  OAI21X1  g11906(.A0(new_n5291_), .A1(new_n3720_), .B0(new_n12162_), .Y(new_n12163_));
  AOI21X1  g11907(.A0(new_n4875_), .A1(new_n3860_), .B0(new_n12163_), .Y(new_n12164_));
  XOR2X1   g11908(.A(new_n12164_), .B(\a[50] ), .Y(new_n12165_));
  XOR2X1   g11909(.A(new_n12165_), .B(new_n12161_), .Y(new_n12166_));
  XOR2X1   g11910(.A(new_n12166_), .B(new_n12122_), .Y(new_n12167_));
  AOI22X1  g11911(.A0(new_n4572_), .A1(\b[45] ), .B0(new_n4571_), .B1(\b[44] ), .Y(new_n12168_));
  OAI21X1  g11912(.A0(new_n4740_), .A1(new_n4339_), .B0(new_n12168_), .Y(new_n12169_));
  AOI21X1  g11913(.A0(new_n4375_), .A1(new_n4338_), .B0(new_n12169_), .Y(new_n12170_));
  XOR2X1   g11914(.A(new_n12170_), .B(\a[47] ), .Y(new_n12171_));
  XOR2X1   g11915(.A(new_n12171_), .B(new_n12167_), .Y(new_n12172_));
  XOR2X1   g11916(.A(new_n12172_), .B(new_n12119_), .Y(new_n12173_));
  AOI22X1  g11917(.A0(new_n4095_), .A1(\b[48] ), .B0(new_n4094_), .B1(\b[47] ), .Y(new_n12174_));
  OAI21X1  g11918(.A0(new_n4233_), .A1(new_n4693_), .B0(new_n12174_), .Y(new_n12175_));
  AOI21X1  g11919(.A0(new_n4692_), .A1(new_n3901_), .B0(new_n12175_), .Y(new_n12176_));
  XOR2X1   g11920(.A(new_n12176_), .B(\a[44] ), .Y(new_n12177_));
  XOR2X1   g11921(.A(new_n12177_), .B(new_n12173_), .Y(new_n12178_));
  AND2X1   g11922(.A(new_n12075_), .B(new_n12022_), .Y(new_n12179_));
  INVX1    g11923(.A(new_n12080_), .Y(new_n12180_));
  AOI21X1  g11924(.A0(new_n12180_), .A1(new_n12076_), .B0(new_n12179_), .Y(new_n12181_));
  XOR2X1   g11925(.A(new_n12181_), .B(new_n12178_), .Y(new_n12182_));
  INVX1    g11926(.A(new_n12182_), .Y(new_n12183_));
  AOI22X1  g11927(.A0(new_n3652_), .A1(\b[51] ), .B0(new_n3651_), .B1(\b[50] ), .Y(new_n12184_));
  OAI21X1  g11928(.A0(new_n3778_), .A1(new_n5237_), .B0(new_n12184_), .Y(new_n12185_));
  AOI21X1  g11929(.A0(new_n5236_), .A1(new_n3480_), .B0(new_n12185_), .Y(new_n12186_));
  XOR2X1   g11930(.A(new_n12186_), .B(\a[41] ), .Y(new_n12187_));
  AND2X1   g11931(.A(new_n12187_), .B(new_n12183_), .Y(new_n12188_));
  INVX1    g11932(.A(new_n12188_), .Y(new_n12189_));
  OAI21X1  g11933(.A0(new_n12187_), .A1(new_n12183_), .B0(new_n12116_), .Y(new_n12190_));
  OR2X1    g11934(.A(new_n12190_), .B(new_n12188_), .Y(new_n12191_));
  NOR2X1   g11935(.A(new_n12187_), .B(new_n12183_), .Y(new_n12192_));
  AOI21X1  g11936(.A0(new_n12189_), .A1(new_n12116_), .B0(new_n12192_), .Y(new_n12193_));
  AOI22X1  g11937(.A0(new_n12193_), .A1(new_n12189_), .B0(new_n12191_), .B1(new_n12116_), .Y(new_n12194_));
  AOI22X1  g11938(.A0(new_n3204_), .A1(\b[54] ), .B0(new_n3203_), .B1(\b[53] ), .Y(new_n12195_));
  OAI21X1  g11939(.A0(new_n3321_), .A1(new_n5808_), .B0(new_n12195_), .Y(new_n12196_));
  AOI21X1  g11940(.A0(new_n5807_), .A1(new_n3080_), .B0(new_n12196_), .Y(new_n12197_));
  XOR2X1   g11941(.A(new_n12197_), .B(\a[38] ), .Y(new_n12198_));
  XOR2X1   g11942(.A(new_n12198_), .B(new_n12194_), .Y(new_n12199_));
  XOR2X1   g11943(.A(new_n12199_), .B(new_n12113_), .Y(new_n12200_));
  AOI22X1  g11944(.A0(new_n2813_), .A1(\b[57] ), .B0(new_n2812_), .B1(\b[56] ), .Y(new_n12201_));
  OAI21X1  g11945(.A0(new_n2946_), .A1(new_n6523_), .B0(new_n12201_), .Y(new_n12202_));
  AOI21X1  g11946(.A0(new_n6522_), .A1(new_n2652_), .B0(new_n12202_), .Y(new_n12203_));
  XOR2X1   g11947(.A(new_n12203_), .B(\a[35] ), .Y(new_n12204_));
  XOR2X1   g11948(.A(new_n12204_), .B(new_n12200_), .Y(new_n12205_));
  INVX1    g11949(.A(new_n12006_), .Y(new_n12206_));
  AND2X1   g11950(.A(new_n12093_), .B(new_n12009_), .Y(new_n12207_));
  AOI21X1  g11951(.A0(new_n12094_), .A1(new_n12206_), .B0(new_n12207_), .Y(new_n12208_));
  XOR2X1   g11952(.A(new_n12208_), .B(new_n12205_), .Y(new_n12209_));
  INVX1    g11953(.A(new_n12209_), .Y(new_n12210_));
  AOI22X1  g11954(.A0(new_n2545_), .A1(\b[60] ), .B0(new_n2544_), .B1(\b[59] ), .Y(new_n12211_));
  OAI21X1  g11955(.A0(new_n2543_), .A1(new_n6930_), .B0(new_n12211_), .Y(new_n12212_));
  AOI21X1  g11956(.A0(new_n6951_), .A1(new_n2260_), .B0(new_n12212_), .Y(new_n12213_));
  XOR2X1   g11957(.A(new_n12213_), .B(\a[32] ), .Y(new_n12214_));
  NOR2X1   g11958(.A(new_n12001_), .B(new_n11998_), .Y(new_n12215_));
  INVX1    g11959(.A(new_n12095_), .Y(new_n12216_));
  AOI21X1  g11960(.A0(new_n12216_), .A1(new_n12002_), .B0(new_n12215_), .Y(new_n12217_));
  XOR2X1   g11961(.A(new_n12217_), .B(new_n12214_), .Y(new_n12218_));
  XOR2X1   g11962(.A(new_n12218_), .B(new_n12210_), .Y(new_n12219_));
  XOR2X1   g11963(.A(new_n12219_), .B(new_n12110_), .Y(new_n12220_));
  XOR2X1   g11964(.A(new_n12220_), .B(new_n12102_), .Y(new_n12221_));
  AND2X1   g11965(.A(new_n12098_), .B(new_n11981_), .Y(new_n12222_));
  INVX1    g11966(.A(new_n12222_), .Y(new_n12223_));
  OAI21X1  g11967(.A0(new_n11979_), .A1(new_n11978_), .B0(new_n12099_), .Y(new_n12224_));
  AND2X1   g11968(.A(new_n12224_), .B(new_n12223_), .Y(new_n12225_));
  XOR2X1   g11969(.A(new_n12225_), .B(new_n12221_), .Y(\f[90] ));
  NOR2X1   g11970(.A(new_n12217_), .B(new_n12214_), .Y(new_n12227_));
  AOI21X1  g11971(.A0(new_n12218_), .A1(new_n12209_), .B0(new_n12227_), .Y(new_n12228_));
  OAI22X1  g11972(.A0(new_n2161_), .A1(new_n7745_), .B0(new_n1910_), .B1(new_n7772_), .Y(new_n12229_));
  AOI21X1  g11973(.A0(new_n7775_), .A1(new_n1907_), .B0(new_n12229_), .Y(new_n12230_));
  XOR2X1   g11974(.A(new_n12230_), .B(\a[29] ), .Y(new_n12231_));
  XOR2X1   g11975(.A(new_n12231_), .B(new_n12228_), .Y(new_n12232_));
  AOI22X1  g11976(.A0(new_n2545_), .A1(\b[61] ), .B0(new_n2544_), .B1(\b[60] ), .Y(new_n12233_));
  OAI21X1  g11977(.A0(new_n2543_), .A1(new_n7339_), .B0(new_n12233_), .Y(new_n12234_));
  AOI21X1  g11978(.A0(new_n7338_), .A1(new_n2260_), .B0(new_n12234_), .Y(new_n12235_));
  XOR2X1   g11979(.A(new_n12235_), .B(\a[32] ), .Y(new_n12236_));
  INVX1    g11980(.A(new_n12236_), .Y(new_n12237_));
  INVX1    g11981(.A(new_n12204_), .Y(new_n12238_));
  NOR2X1   g11982(.A(new_n12208_), .B(new_n12205_), .Y(new_n12239_));
  AOI21X1  g11983(.A0(new_n12238_), .A1(new_n12200_), .B0(new_n12239_), .Y(new_n12240_));
  XOR2X1   g11984(.A(new_n12240_), .B(new_n12237_), .Y(new_n12241_));
  NOR2X1   g11985(.A(new_n12198_), .B(new_n12194_), .Y(new_n12242_));
  AOI21X1  g11986(.A0(new_n12199_), .A1(new_n12113_), .B0(new_n12242_), .Y(new_n12243_));
  INVX1    g11987(.A(new_n12243_), .Y(new_n12244_));
  XOR2X1   g11988(.A(new_n12155_), .B(new_n5423_), .Y(new_n12245_));
  NOR2X1   g11989(.A(new_n12160_), .B(new_n12157_), .Y(new_n12246_));
  AOI21X1  g11990(.A0(new_n12245_), .A1(new_n12152_), .B0(new_n12246_), .Y(new_n12247_));
  INVX1    g11991(.A(new_n12247_), .Y(new_n12248_));
  AOI22X1  g11992(.A0(new_n5430_), .A1(\b[40] ), .B0(new_n5427_), .B1(\b[39] ), .Y(new_n12249_));
  OAI21X1  g11993(.A0(new_n5891_), .A1(new_n3575_), .B0(new_n12249_), .Y(new_n12250_));
  AOI21X1  g11994(.A0(new_n5425_), .A1(new_n3574_), .B0(new_n12250_), .Y(new_n12251_));
  XOR2X1   g11995(.A(new_n12251_), .B(\a[53] ), .Y(new_n12252_));
  XOR2X1   g11996(.A(new_n12147_), .B(new_n6019_), .Y(new_n12253_));
  AND2X1   g11997(.A(new_n12253_), .B(new_n12144_), .Y(new_n12254_));
  NOR2X1   g11998(.A(new_n12151_), .B(new_n12149_), .Y(new_n12255_));
  NOR2X1   g11999(.A(new_n12255_), .B(new_n12254_), .Y(new_n12256_));
  AOI22X1  g12000(.A0(new_n7818_), .A1(\b[27] ), .B0(new_n7817_), .B1(\b[28] ), .Y(new_n12257_));
  INVX1    g12001(.A(new_n12257_), .Y(new_n12258_));
  NOR2X1   g12002(.A(new_n12135_), .B(\a[26] ), .Y(new_n12259_));
  AOI21X1  g12003(.A0(new_n12136_), .A1(new_n12134_), .B0(new_n12259_), .Y(new_n12260_));
  XOR2X1   g12004(.A(new_n12260_), .B(new_n12258_), .Y(new_n12261_));
  INVX1    g12005(.A(new_n12261_), .Y(new_n12262_));
  AOI22X1  g12006(.A0(new_n7192_), .A1(\b[31] ), .B0(new_n7189_), .B1(\b[30] ), .Y(new_n12263_));
  OAI21X1  g12007(.A0(new_n7627_), .A1(new_n2359_), .B0(new_n12263_), .Y(new_n12264_));
  AOI21X1  g12008(.A0(new_n7187_), .A1(new_n2358_), .B0(new_n12264_), .Y(new_n12265_));
  XOR2X1   g12009(.A(new_n12265_), .B(\a[62] ), .Y(new_n12266_));
  XOR2X1   g12010(.A(new_n12266_), .B(new_n12262_), .Y(new_n12267_));
  INVX1    g12011(.A(new_n12267_), .Y(new_n12268_));
  AND2X1   g12012(.A(new_n12137_), .B(new_n12133_), .Y(new_n12269_));
  INVX1    g12013(.A(new_n12142_), .Y(new_n12270_));
  AOI21X1  g12014(.A0(new_n12270_), .A1(new_n12138_), .B0(new_n12269_), .Y(new_n12271_));
  XOR2X1   g12015(.A(new_n12271_), .B(new_n12268_), .Y(new_n12272_));
  AOI22X1  g12016(.A0(new_n6603_), .A1(\b[34] ), .B0(new_n6600_), .B1(\b[33] ), .Y(new_n12273_));
  OAI21X1  g12017(.A0(new_n6804_), .A1(new_n2612_), .B0(new_n12273_), .Y(new_n12274_));
  AOI21X1  g12018(.A0(new_n6598_), .A1(new_n2759_), .B0(new_n12274_), .Y(new_n12275_));
  XOR2X1   g12019(.A(new_n12275_), .B(\a[59] ), .Y(new_n12276_));
  XOR2X1   g12020(.A(new_n12276_), .B(new_n12272_), .Y(new_n12277_));
  NOR2X1   g12021(.A(new_n12128_), .B(new_n12126_), .Y(new_n12278_));
  INVX1    g12022(.A(new_n12143_), .Y(new_n12279_));
  AOI21X1  g12023(.A0(new_n12279_), .A1(new_n12129_), .B0(new_n12278_), .Y(new_n12280_));
  XOR2X1   g12024(.A(new_n12280_), .B(new_n12277_), .Y(new_n12281_));
  AOI22X1  g12025(.A0(new_n6438_), .A1(\b[37] ), .B0(new_n6437_), .B1(\b[36] ), .Y(new_n12282_));
  OAI21X1  g12026(.A0(new_n6436_), .A1(new_n3156_), .B0(new_n12282_), .Y(new_n12283_));
  AOI21X1  g12027(.A0(new_n6023_), .A1(new_n3155_), .B0(new_n12283_), .Y(new_n12284_));
  XOR2X1   g12028(.A(new_n12284_), .B(\a[56] ), .Y(new_n12285_));
  INVX1    g12029(.A(new_n12285_), .Y(new_n12286_));
  XOR2X1   g12030(.A(new_n12286_), .B(new_n12281_), .Y(new_n12287_));
  XOR2X1   g12031(.A(new_n12287_), .B(new_n12256_), .Y(new_n12288_));
  XOR2X1   g12032(.A(new_n12288_), .B(new_n12252_), .Y(new_n12289_));
  XOR2X1   g12033(.A(new_n12289_), .B(new_n12248_), .Y(new_n12290_));
  AOI22X1  g12034(.A0(new_n4880_), .A1(\b[43] ), .B0(new_n4877_), .B1(\b[42] ), .Y(new_n12291_));
  OAI21X1  g12035(.A0(new_n5291_), .A1(new_n4015_), .B0(new_n12291_), .Y(new_n12292_));
  AOI21X1  g12036(.A0(new_n4875_), .A1(new_n4014_), .B0(new_n12292_), .Y(new_n12293_));
  XOR2X1   g12037(.A(new_n12293_), .B(\a[50] ), .Y(new_n12294_));
  XOR2X1   g12038(.A(new_n12294_), .B(new_n12290_), .Y(new_n12295_));
  INVX1    g12039(.A(new_n12161_), .Y(new_n12296_));
  NOR2X1   g12040(.A(new_n12165_), .B(new_n12296_), .Y(new_n12297_));
  INVX1    g12041(.A(new_n12166_), .Y(new_n12298_));
  AOI21X1  g12042(.A0(new_n12298_), .A1(new_n12122_), .B0(new_n12297_), .Y(new_n12299_));
  XOR2X1   g12043(.A(new_n12299_), .B(new_n12295_), .Y(new_n12300_));
  AOI22X1  g12044(.A0(new_n4572_), .A1(\b[46] ), .B0(new_n4571_), .B1(\b[45] ), .Y(new_n12301_));
  OAI21X1  g12045(.A0(new_n4740_), .A1(new_n4336_), .B0(new_n12301_), .Y(new_n12302_));
  AOI21X1  g12046(.A0(new_n4509_), .A1(new_n4375_), .B0(new_n12302_), .Y(new_n12303_));
  XOR2X1   g12047(.A(new_n12303_), .B(\a[47] ), .Y(new_n12304_));
  XOR2X1   g12048(.A(new_n12304_), .B(new_n12300_), .Y(new_n12305_));
  NOR2X1   g12049(.A(new_n12171_), .B(new_n12167_), .Y(new_n12306_));
  AOI21X1  g12050(.A0(new_n12172_), .A1(new_n12119_), .B0(new_n12306_), .Y(new_n12307_));
  XOR2X1   g12051(.A(new_n12307_), .B(new_n12305_), .Y(new_n12308_));
  AOI22X1  g12052(.A0(new_n4095_), .A1(\b[49] ), .B0(new_n4094_), .B1(\b[48] ), .Y(new_n12309_));
  OAI21X1  g12053(.A0(new_n4233_), .A1(new_n5039_), .B0(new_n12309_), .Y(new_n12310_));
  AOI21X1  g12054(.A0(new_n5038_), .A1(new_n3901_), .B0(new_n12310_), .Y(new_n12311_));
  XOR2X1   g12055(.A(new_n12311_), .B(\a[44] ), .Y(new_n12312_));
  XOR2X1   g12056(.A(new_n12312_), .B(new_n12308_), .Y(new_n12313_));
  INVX1    g12057(.A(new_n12177_), .Y(new_n12314_));
  NOR2X1   g12058(.A(new_n12181_), .B(new_n12178_), .Y(new_n12315_));
  AOI21X1  g12059(.A0(new_n12314_), .A1(new_n12173_), .B0(new_n12315_), .Y(new_n12316_));
  XOR2X1   g12060(.A(new_n12316_), .B(new_n12313_), .Y(new_n12317_));
  AOI22X1  g12061(.A0(new_n3652_), .A1(\b[52] ), .B0(new_n3651_), .B1(\b[51] ), .Y(new_n12318_));
  OAI21X1  g12062(.A0(new_n3778_), .A1(new_n5234_), .B0(new_n12318_), .Y(new_n12319_));
  AOI21X1  g12063(.A0(new_n5590_), .A1(new_n3480_), .B0(new_n12319_), .Y(new_n12320_));
  XOR2X1   g12064(.A(new_n12320_), .B(\a[41] ), .Y(new_n12321_));
  XOR2X1   g12065(.A(new_n12321_), .B(new_n12317_), .Y(new_n12322_));
  INVX1    g12066(.A(new_n12322_), .Y(new_n12323_));
  XOR2X1   g12067(.A(new_n12323_), .B(new_n12193_), .Y(new_n12324_));
  AOI22X1  g12068(.A0(new_n3204_), .A1(\b[55] ), .B0(new_n3203_), .B1(\b[54] ), .Y(new_n12325_));
  OAI21X1  g12069(.A0(new_n3321_), .A1(new_n6151_), .B0(new_n12325_), .Y(new_n12326_));
  AOI21X1  g12070(.A0(new_n6150_), .A1(new_n3080_), .B0(new_n12326_), .Y(new_n12327_));
  XOR2X1   g12071(.A(new_n12327_), .B(\a[38] ), .Y(new_n12328_));
  XOR2X1   g12072(.A(new_n12328_), .B(new_n12324_), .Y(new_n12329_));
  XOR2X1   g12073(.A(new_n12329_), .B(new_n12244_), .Y(new_n12330_));
  AOI22X1  g12074(.A0(new_n2813_), .A1(\b[58] ), .B0(new_n2812_), .B1(\b[57] ), .Y(new_n12331_));
  OAI21X1  g12075(.A0(new_n2946_), .A1(new_n6520_), .B0(new_n12331_), .Y(new_n12332_));
  AOI21X1  g12076(.A0(new_n6732_), .A1(new_n2652_), .B0(new_n12332_), .Y(new_n12333_));
  XOR2X1   g12077(.A(new_n12333_), .B(\a[35] ), .Y(new_n12334_));
  XOR2X1   g12078(.A(new_n12334_), .B(new_n12330_), .Y(new_n12335_));
  XOR2X1   g12079(.A(new_n12335_), .B(new_n12241_), .Y(new_n12336_));
  XOR2X1   g12080(.A(new_n12336_), .B(new_n12232_), .Y(new_n12337_));
  INVX1    g12081(.A(new_n12337_), .Y(new_n12338_));
  INVX1    g12082(.A(new_n12109_), .Y(new_n12339_));
  NOR2X1   g12083(.A(new_n12219_), .B(new_n12110_), .Y(new_n12340_));
  AOI21X1  g12084(.A0(new_n12339_), .A1(new_n12105_), .B0(new_n12340_), .Y(new_n12341_));
  XOR2X1   g12085(.A(new_n12341_), .B(new_n12338_), .Y(new_n12342_));
  INVX1    g12086(.A(new_n12102_), .Y(new_n12343_));
  AND2X1   g12087(.A(new_n12220_), .B(new_n12343_), .Y(new_n12344_));
  AOI21X1  g12088(.A0(new_n12224_), .A1(new_n12223_), .B0(new_n12221_), .Y(new_n12345_));
  OR2X1    g12089(.A(new_n12345_), .B(new_n12344_), .Y(new_n12346_));
  XOR2X1   g12090(.A(new_n12346_), .B(new_n12342_), .Y(\f[91] ));
  NOR2X1   g12091(.A(new_n12341_), .B(new_n12338_), .Y(new_n12348_));
  INVX1    g12092(.A(new_n12348_), .Y(new_n12349_));
  OAI21X1  g12093(.A0(new_n12345_), .A1(new_n12344_), .B0(new_n12342_), .Y(new_n12350_));
  AND2X1   g12094(.A(new_n12350_), .B(new_n12349_), .Y(new_n12351_));
  NOR2X1   g12095(.A(new_n12231_), .B(new_n12228_), .Y(new_n12352_));
  AOI21X1  g12096(.A0(new_n12336_), .A1(new_n12232_), .B0(new_n12352_), .Y(new_n12353_));
  OR2X1    g12097(.A(new_n12240_), .B(new_n12236_), .Y(new_n12354_));
  OR2X1    g12098(.A(new_n12335_), .B(new_n12241_), .Y(new_n12355_));
  AND2X1   g12099(.A(new_n12355_), .B(new_n12354_), .Y(new_n12356_));
  AOI22X1  g12100(.A0(new_n7774_), .A1(new_n1907_), .B0(new_n2045_), .B1(\b[63] ), .Y(new_n12357_));
  XOR2X1   g12101(.A(new_n12357_), .B(\a[29] ), .Y(new_n12358_));
  XOR2X1   g12102(.A(new_n12358_), .B(new_n12356_), .Y(new_n12359_));
  AOI22X1  g12103(.A0(new_n2545_), .A1(\b[62] ), .B0(new_n2544_), .B1(\b[61] ), .Y(new_n12360_));
  OAI21X1  g12104(.A0(new_n2543_), .A1(new_n7559_), .B0(new_n12360_), .Y(new_n12361_));
  AOI21X1  g12105(.A0(new_n7558_), .A1(new_n2260_), .B0(new_n12361_), .Y(new_n12362_));
  XOR2X1   g12106(.A(new_n12362_), .B(\a[32] ), .Y(new_n12363_));
  INVX1    g12107(.A(new_n12363_), .Y(new_n12364_));
  AND2X1   g12108(.A(new_n12329_), .B(new_n12244_), .Y(new_n12365_));
  INVX1    g12109(.A(new_n12334_), .Y(new_n12366_));
  AOI21X1  g12110(.A0(new_n12366_), .A1(new_n12330_), .B0(new_n12365_), .Y(new_n12367_));
  XOR2X1   g12111(.A(new_n12367_), .B(new_n12364_), .Y(new_n12368_));
  OR2X1    g12112(.A(new_n12322_), .B(new_n12193_), .Y(new_n12369_));
  OAI21X1  g12113(.A0(new_n12328_), .A1(new_n12324_), .B0(new_n12369_), .Y(new_n12370_));
  AOI22X1  g12114(.A0(new_n3204_), .A1(\b[56] ), .B0(new_n3203_), .B1(\b[55] ), .Y(new_n12371_));
  OAI21X1  g12115(.A0(new_n3321_), .A1(new_n6148_), .B0(new_n12371_), .Y(new_n12372_));
  AOI21X1  g12116(.A0(new_n6342_), .A1(new_n3080_), .B0(new_n12372_), .Y(new_n12373_));
  XOR2X1   g12117(.A(new_n12373_), .B(new_n3078_), .Y(new_n12374_));
  AND2X1   g12118(.A(new_n12316_), .B(new_n12313_), .Y(new_n12375_));
  OR2X1    g12119(.A(new_n12316_), .B(new_n12313_), .Y(new_n12376_));
  OAI21X1  g12120(.A0(new_n12321_), .A1(new_n12375_), .B0(new_n12376_), .Y(new_n12377_));
  AOI22X1  g12121(.A0(new_n3652_), .A1(\b[53] ), .B0(new_n3651_), .B1(\b[52] ), .Y(new_n12378_));
  OAI21X1  g12122(.A0(new_n3778_), .A1(new_n5787_), .B0(new_n12378_), .Y(new_n12379_));
  AOI21X1  g12123(.A0(new_n5786_), .A1(new_n3480_), .B0(new_n12379_), .Y(new_n12380_));
  XOR2X1   g12124(.A(new_n12380_), .B(\a[41] ), .Y(new_n12381_));
  NOR2X1   g12125(.A(new_n12307_), .B(new_n12305_), .Y(new_n12382_));
  INVX1    g12126(.A(new_n12382_), .Y(new_n12383_));
  INVX1    g12127(.A(new_n12308_), .Y(new_n12384_));
  OAI21X1  g12128(.A0(new_n12312_), .A1(new_n12384_), .B0(new_n12383_), .Y(new_n12385_));
  INVX1    g12129(.A(new_n12385_), .Y(new_n12386_));
  AND2X1   g12130(.A(new_n12289_), .B(new_n12248_), .Y(new_n12387_));
  INVX1    g12131(.A(new_n12387_), .Y(new_n12388_));
  INVX1    g12132(.A(new_n12290_), .Y(new_n12389_));
  OAI21X1  g12133(.A0(new_n12294_), .A1(new_n12389_), .B0(new_n12388_), .Y(new_n12390_));
  AOI22X1  g12134(.A0(new_n4880_), .A1(\b[44] ), .B0(new_n4877_), .B1(\b[43] ), .Y(new_n12391_));
  OAI21X1  g12135(.A0(new_n5291_), .A1(new_n4012_), .B0(new_n12391_), .Y(new_n12392_));
  AOI21X1  g12136(.A0(new_n4875_), .A1(new_n4178_), .B0(new_n12392_), .Y(new_n12393_));
  XOR2X1   g12137(.A(new_n12393_), .B(new_n4873_), .Y(new_n12394_));
  OAI21X1  g12138(.A0(new_n12255_), .A1(new_n12254_), .B0(new_n12287_), .Y(new_n12395_));
  OR2X1    g12139(.A(new_n12288_), .B(new_n12252_), .Y(new_n12396_));
  AND2X1   g12140(.A(new_n12396_), .B(new_n12395_), .Y(new_n12397_));
  NOR2X1   g12141(.A(new_n12271_), .B(new_n12268_), .Y(new_n12398_));
  INVX1    g12142(.A(new_n12398_), .Y(new_n12399_));
  INVX1    g12143(.A(new_n12272_), .Y(new_n12400_));
  OAI21X1  g12144(.A0(new_n12276_), .A1(new_n12400_), .B0(new_n12399_), .Y(new_n12401_));
  AOI22X1  g12145(.A0(new_n6603_), .A1(\b[35] ), .B0(new_n6600_), .B1(\b[34] ), .Y(new_n12402_));
  OAI21X1  g12146(.A0(new_n6804_), .A1(new_n2893_), .B0(new_n12402_), .Y(new_n12403_));
  AOI21X1  g12147(.A0(new_n6598_), .A1(new_n2892_), .B0(new_n12403_), .Y(new_n12404_));
  XOR2X1   g12148(.A(new_n12404_), .B(\a[59] ), .Y(new_n12405_));
  NOR2X1   g12149(.A(new_n12260_), .B(new_n12258_), .Y(new_n12406_));
  INVX1    g12150(.A(new_n12406_), .Y(new_n12407_));
  OAI21X1  g12151(.A0(new_n12266_), .A1(new_n12262_), .B0(new_n12407_), .Y(new_n12408_));
  AOI22X1  g12152(.A0(new_n7818_), .A1(\b[28] ), .B0(new_n7817_), .B1(\b[29] ), .Y(new_n12409_));
  NOR2X1   g12153(.A(new_n12409_), .B(new_n12258_), .Y(new_n12410_));
  INVX1    g12154(.A(new_n12410_), .Y(new_n12411_));
  XOR2X1   g12155(.A(new_n12409_), .B(new_n12258_), .Y(new_n12412_));
  INVX1    g12156(.A(new_n12412_), .Y(new_n12413_));
  AND2X1   g12157(.A(new_n12409_), .B(new_n12258_), .Y(new_n12414_));
  AOI21X1  g12158(.A0(new_n12411_), .A1(new_n12408_), .B0(new_n12414_), .Y(new_n12415_));
  AOI22X1  g12159(.A0(new_n12415_), .A1(new_n12411_), .B0(new_n12413_), .B1(new_n12408_), .Y(new_n12416_));
  AOI22X1  g12160(.A0(new_n7192_), .A1(\b[32] ), .B0(new_n7189_), .B1(\b[31] ), .Y(new_n12417_));
  OAI21X1  g12161(.A0(new_n7627_), .A1(new_n2356_), .B0(new_n12417_), .Y(new_n12418_));
  AOI21X1  g12162(.A0(new_n7187_), .A1(new_n2495_), .B0(new_n12418_), .Y(new_n12419_));
  XOR2X1   g12163(.A(new_n12419_), .B(\a[62] ), .Y(new_n12420_));
  INVX1    g12164(.A(new_n12420_), .Y(new_n12421_));
  XOR2X1   g12165(.A(new_n12421_), .B(new_n12416_), .Y(new_n12422_));
  XOR2X1   g12166(.A(new_n12422_), .B(new_n12405_), .Y(new_n12423_));
  XOR2X1   g12167(.A(new_n12423_), .B(new_n12401_), .Y(new_n12424_));
  AOI22X1  g12168(.A0(new_n6438_), .A1(\b[38] ), .B0(new_n6437_), .B1(\b[37] ), .Y(new_n12425_));
  OAI21X1  g12169(.A0(new_n6436_), .A1(new_n3276_), .B0(new_n12425_), .Y(new_n12426_));
  AOI21X1  g12170(.A0(new_n6023_), .A1(new_n3275_), .B0(new_n12426_), .Y(new_n12427_));
  XOR2X1   g12171(.A(new_n12427_), .B(\a[56] ), .Y(new_n12428_));
  XOR2X1   g12172(.A(new_n12428_), .B(new_n12424_), .Y(new_n12429_));
  NOR2X1   g12173(.A(new_n12280_), .B(new_n12277_), .Y(new_n12430_));
  AOI21X1  g12174(.A0(new_n12286_), .A1(new_n12281_), .B0(new_n12430_), .Y(new_n12431_));
  XOR2X1   g12175(.A(new_n12431_), .B(new_n12429_), .Y(new_n12432_));
  AOI22X1  g12176(.A0(new_n5430_), .A1(\b[41] ), .B0(new_n5427_), .B1(\b[40] ), .Y(new_n12433_));
  OAI21X1  g12177(.A0(new_n5891_), .A1(new_n3723_), .B0(new_n12433_), .Y(new_n12434_));
  AOI21X1  g12178(.A0(new_n5425_), .A1(new_n3722_), .B0(new_n12434_), .Y(new_n12435_));
  XOR2X1   g12179(.A(new_n12435_), .B(\a[53] ), .Y(new_n12436_));
  XOR2X1   g12180(.A(new_n12436_), .B(new_n12432_), .Y(new_n12437_));
  XOR2X1   g12181(.A(new_n12437_), .B(new_n12397_), .Y(new_n12438_));
  XOR2X1   g12182(.A(new_n12438_), .B(new_n12394_), .Y(new_n12439_));
  XOR2X1   g12183(.A(new_n12439_), .B(new_n12390_), .Y(new_n12440_));
  AOI22X1  g12184(.A0(new_n4572_), .A1(\b[47] ), .B0(new_n4571_), .B1(\b[46] ), .Y(new_n12441_));
  OAI21X1  g12185(.A0(new_n4740_), .A1(new_n4674_), .B0(new_n12441_), .Y(new_n12442_));
  AOI21X1  g12186(.A0(new_n4673_), .A1(new_n4375_), .B0(new_n12442_), .Y(new_n12443_));
  XOR2X1   g12187(.A(new_n12443_), .B(\a[47] ), .Y(new_n12444_));
  XOR2X1   g12188(.A(new_n12444_), .B(new_n12440_), .Y(new_n12445_));
  INVX1    g12189(.A(new_n12445_), .Y(new_n12446_));
  NOR2X1   g12190(.A(new_n12299_), .B(new_n12295_), .Y(new_n12447_));
  INVX1    g12191(.A(new_n12304_), .Y(new_n12448_));
  AOI21X1  g12192(.A0(new_n12448_), .A1(new_n12300_), .B0(new_n12447_), .Y(new_n12449_));
  XOR2X1   g12193(.A(new_n12449_), .B(new_n12446_), .Y(new_n12450_));
  AOI22X1  g12194(.A0(new_n4095_), .A1(\b[50] ), .B0(new_n4094_), .B1(\b[49] ), .Y(new_n12451_));
  OAI21X1  g12195(.A0(new_n4233_), .A1(new_n5036_), .B0(new_n12451_), .Y(new_n12452_));
  AOI21X1  g12196(.A0(new_n5204_), .A1(new_n3901_), .B0(new_n12452_), .Y(new_n12453_));
  XOR2X1   g12197(.A(new_n12453_), .B(\a[44] ), .Y(new_n12454_));
  XOR2X1   g12198(.A(new_n12454_), .B(new_n12450_), .Y(new_n12455_));
  XOR2X1   g12199(.A(new_n12455_), .B(new_n12386_), .Y(new_n12456_));
  XOR2X1   g12200(.A(new_n12456_), .B(new_n12381_), .Y(new_n12457_));
  XOR2X1   g12201(.A(new_n12457_), .B(new_n12377_), .Y(new_n12458_));
  XOR2X1   g12202(.A(new_n12458_), .B(new_n12374_), .Y(new_n12459_));
  XOR2X1   g12203(.A(new_n12459_), .B(new_n12370_), .Y(new_n12460_));
  AOI22X1  g12204(.A0(new_n2813_), .A1(\b[59] ), .B0(new_n2812_), .B1(\b[58] ), .Y(new_n12461_));
  OAI21X1  g12205(.A0(new_n2946_), .A1(new_n6933_), .B0(new_n12461_), .Y(new_n12462_));
  AOI21X1  g12206(.A0(new_n6932_), .A1(new_n2652_), .B0(new_n12462_), .Y(new_n12463_));
  XOR2X1   g12207(.A(new_n12463_), .B(\a[35] ), .Y(new_n12464_));
  XOR2X1   g12208(.A(new_n12464_), .B(new_n12460_), .Y(new_n12465_));
  XOR2X1   g12209(.A(new_n12465_), .B(new_n12368_), .Y(new_n12466_));
  XOR2X1   g12210(.A(new_n12466_), .B(new_n12359_), .Y(new_n12467_));
  XOR2X1   g12211(.A(new_n12467_), .B(new_n12353_), .Y(new_n12468_));
  XOR2X1   g12212(.A(new_n12468_), .B(new_n12351_), .Y(\f[92] ));
  INVX1    g12213(.A(new_n12353_), .Y(new_n12470_));
  AND2X1   g12214(.A(new_n12467_), .B(new_n12470_), .Y(new_n12471_));
  AOI21X1  g12215(.A0(new_n12350_), .A1(new_n12349_), .B0(new_n12468_), .Y(new_n12472_));
  OR2X1    g12216(.A(new_n12472_), .B(new_n12471_), .Y(new_n12473_));
  NAND2X1  g12217(.A(new_n12466_), .B(new_n12359_), .Y(new_n12474_));
  OAI21X1  g12218(.A0(new_n12358_), .A1(new_n12356_), .B0(new_n12474_), .Y(new_n12475_));
  AND2X1   g12219(.A(new_n12455_), .B(new_n12385_), .Y(new_n12476_));
  INVX1    g12220(.A(new_n12476_), .Y(new_n12477_));
  OAI21X1  g12221(.A0(new_n12456_), .A1(new_n12381_), .B0(new_n12477_), .Y(new_n12478_));
  NOR2X1   g12222(.A(new_n12449_), .B(new_n12445_), .Y(new_n12479_));
  INVX1    g12223(.A(new_n12479_), .Y(new_n12480_));
  OAI21X1  g12224(.A0(new_n12454_), .A1(new_n12450_), .B0(new_n12480_), .Y(new_n12481_));
  NOR2X1   g12225(.A(new_n12437_), .B(new_n12397_), .Y(new_n12482_));
  AOI21X1  g12226(.A0(new_n12438_), .A1(new_n12394_), .B0(new_n12482_), .Y(new_n12483_));
  INVX1    g12227(.A(new_n12483_), .Y(new_n12484_));
  OR2X1    g12228(.A(new_n12431_), .B(new_n12429_), .Y(new_n12485_));
  INVX1    g12229(.A(new_n12432_), .Y(new_n12486_));
  OAI21X1  g12230(.A0(new_n12436_), .A1(new_n12486_), .B0(new_n12485_), .Y(new_n12487_));
  OR2X1    g12231(.A(new_n12420_), .B(new_n12416_), .Y(new_n12488_));
  OAI21X1  g12232(.A0(new_n12422_), .A1(new_n12405_), .B0(new_n12488_), .Y(new_n12489_));
  AOI22X1  g12233(.A0(new_n7818_), .A1(\b[29] ), .B0(new_n7817_), .B1(\b[30] ), .Y(new_n12490_));
  XOR2X1   g12234(.A(new_n12490_), .B(\a[29] ), .Y(new_n12491_));
  XOR2X1   g12235(.A(new_n12491_), .B(new_n12409_), .Y(new_n12492_));
  XOR2X1   g12236(.A(new_n12492_), .B(new_n12415_), .Y(new_n12493_));
  AOI22X1  g12237(.A0(new_n7192_), .A1(\b[33] ), .B0(new_n7189_), .B1(\b[32] ), .Y(new_n12494_));
  OAI21X1  g12238(.A0(new_n7627_), .A1(new_n2615_), .B0(new_n12494_), .Y(new_n12495_));
  AOI21X1  g12239(.A0(new_n7187_), .A1(new_n2614_), .B0(new_n12495_), .Y(new_n12496_));
  XOR2X1   g12240(.A(new_n12496_), .B(\a[62] ), .Y(new_n12497_));
  XOR2X1   g12241(.A(new_n12497_), .B(new_n12493_), .Y(new_n12498_));
  AOI22X1  g12242(.A0(new_n6603_), .A1(\b[36] ), .B0(new_n6600_), .B1(\b[35] ), .Y(new_n12499_));
  OAI21X1  g12243(.A0(new_n6804_), .A1(new_n2890_), .B0(new_n12499_), .Y(new_n12500_));
  AOI21X1  g12244(.A0(new_n6598_), .A1(new_n3015_), .B0(new_n12500_), .Y(new_n12501_));
  XOR2X1   g12245(.A(new_n12501_), .B(\a[59] ), .Y(new_n12502_));
  XOR2X1   g12246(.A(new_n12502_), .B(new_n12498_), .Y(new_n12503_));
  XOR2X1   g12247(.A(new_n12503_), .B(new_n12489_), .Y(new_n12504_));
  AOI22X1  g12248(.A0(new_n6438_), .A1(\b[39] ), .B0(new_n6437_), .B1(\b[38] ), .Y(new_n12505_));
  OAI21X1  g12249(.A0(new_n6436_), .A1(new_n3413_), .B0(new_n12505_), .Y(new_n12506_));
  AOI21X1  g12250(.A0(new_n6023_), .A1(new_n3412_), .B0(new_n12506_), .Y(new_n12507_));
  XOR2X1   g12251(.A(new_n12507_), .B(\a[56] ), .Y(new_n12508_));
  XOR2X1   g12252(.A(new_n12508_), .B(new_n12504_), .Y(new_n12509_));
  AND2X1   g12253(.A(new_n12423_), .B(new_n12401_), .Y(new_n12510_));
  INVX1    g12254(.A(new_n12428_), .Y(new_n12511_));
  AOI21X1  g12255(.A0(new_n12511_), .A1(new_n12424_), .B0(new_n12510_), .Y(new_n12512_));
  XOR2X1   g12256(.A(new_n12512_), .B(new_n12509_), .Y(new_n12513_));
  AOI22X1  g12257(.A0(new_n5430_), .A1(\b[42] ), .B0(new_n5427_), .B1(\b[41] ), .Y(new_n12514_));
  OAI21X1  g12258(.A0(new_n5891_), .A1(new_n3720_), .B0(new_n12514_), .Y(new_n12515_));
  AOI21X1  g12259(.A0(new_n5425_), .A1(new_n3860_), .B0(new_n12515_), .Y(new_n12516_));
  XOR2X1   g12260(.A(new_n12516_), .B(\a[53] ), .Y(new_n12517_));
  XOR2X1   g12261(.A(new_n12517_), .B(new_n12513_), .Y(new_n12518_));
  XOR2X1   g12262(.A(new_n12518_), .B(new_n12487_), .Y(new_n12519_));
  AOI22X1  g12263(.A0(new_n4880_), .A1(\b[45] ), .B0(new_n4877_), .B1(\b[44] ), .Y(new_n12520_));
  OAI21X1  g12264(.A0(new_n5291_), .A1(new_n4339_), .B0(new_n12520_), .Y(new_n12521_));
  AOI21X1  g12265(.A0(new_n4875_), .A1(new_n4338_), .B0(new_n12521_), .Y(new_n12522_));
  XOR2X1   g12266(.A(new_n12522_), .B(\a[50] ), .Y(new_n12523_));
  XOR2X1   g12267(.A(new_n12523_), .B(new_n12519_), .Y(new_n12524_));
  XOR2X1   g12268(.A(new_n12524_), .B(new_n12484_), .Y(new_n12525_));
  AOI22X1  g12269(.A0(new_n4572_), .A1(\b[48] ), .B0(new_n4571_), .B1(\b[47] ), .Y(new_n12526_));
  OAI21X1  g12270(.A0(new_n4740_), .A1(new_n4693_), .B0(new_n12526_), .Y(new_n12527_));
  AOI21X1  g12271(.A0(new_n4692_), .A1(new_n4375_), .B0(new_n12527_), .Y(new_n12528_));
  XOR2X1   g12272(.A(new_n12528_), .B(\a[47] ), .Y(new_n12529_));
  XOR2X1   g12273(.A(new_n12529_), .B(new_n12525_), .Y(new_n12530_));
  AND2X1   g12274(.A(new_n12439_), .B(new_n12390_), .Y(new_n12531_));
  INVX1    g12275(.A(new_n12444_), .Y(new_n12532_));
  AOI21X1  g12276(.A0(new_n12532_), .A1(new_n12440_), .B0(new_n12531_), .Y(new_n12533_));
  XOR2X1   g12277(.A(new_n12533_), .B(new_n12530_), .Y(new_n12534_));
  INVX1    g12278(.A(new_n12534_), .Y(new_n12535_));
  AOI22X1  g12279(.A0(new_n4095_), .A1(\b[51] ), .B0(new_n4094_), .B1(\b[50] ), .Y(new_n12536_));
  OAI21X1  g12280(.A0(new_n4233_), .A1(new_n5237_), .B0(new_n12536_), .Y(new_n12537_));
  AOI21X1  g12281(.A0(new_n5236_), .A1(new_n3901_), .B0(new_n12537_), .Y(new_n12538_));
  XOR2X1   g12282(.A(new_n12538_), .B(\a[44] ), .Y(new_n12539_));
  AND2X1   g12283(.A(new_n12539_), .B(new_n12535_), .Y(new_n12540_));
  INVX1    g12284(.A(new_n12540_), .Y(new_n12541_));
  OAI21X1  g12285(.A0(new_n12539_), .A1(new_n12535_), .B0(new_n12481_), .Y(new_n12542_));
  OR2X1    g12286(.A(new_n12542_), .B(new_n12540_), .Y(new_n12543_));
  NOR2X1   g12287(.A(new_n12539_), .B(new_n12535_), .Y(new_n12544_));
  AOI21X1  g12288(.A0(new_n12541_), .A1(new_n12481_), .B0(new_n12544_), .Y(new_n12545_));
  AOI22X1  g12289(.A0(new_n12545_), .A1(new_n12541_), .B0(new_n12543_), .B1(new_n12481_), .Y(new_n12546_));
  AOI22X1  g12290(.A0(new_n3652_), .A1(\b[54] ), .B0(new_n3651_), .B1(\b[53] ), .Y(new_n12547_));
  OAI21X1  g12291(.A0(new_n3778_), .A1(new_n5808_), .B0(new_n12547_), .Y(new_n12548_));
  AOI21X1  g12292(.A0(new_n5807_), .A1(new_n3480_), .B0(new_n12548_), .Y(new_n12549_));
  XOR2X1   g12293(.A(new_n12549_), .B(\a[41] ), .Y(new_n12550_));
  XOR2X1   g12294(.A(new_n12550_), .B(new_n12546_), .Y(new_n12551_));
  XOR2X1   g12295(.A(new_n12551_), .B(new_n12478_), .Y(new_n12552_));
  AOI22X1  g12296(.A0(new_n3204_), .A1(\b[57] ), .B0(new_n3203_), .B1(\b[56] ), .Y(new_n12553_));
  OAI21X1  g12297(.A0(new_n3321_), .A1(new_n6523_), .B0(new_n12553_), .Y(new_n12554_));
  AOI21X1  g12298(.A0(new_n6522_), .A1(new_n3080_), .B0(new_n12554_), .Y(new_n12555_));
  XOR2X1   g12299(.A(new_n12555_), .B(\a[38] ), .Y(new_n12556_));
  XOR2X1   g12300(.A(new_n12556_), .B(new_n12552_), .Y(new_n12557_));
  AND2X1   g12301(.A(new_n12457_), .B(new_n12377_), .Y(new_n12558_));
  AOI21X1  g12302(.A0(new_n12458_), .A1(new_n12374_), .B0(new_n12558_), .Y(new_n12559_));
  XOR2X1   g12303(.A(new_n12559_), .B(new_n12557_), .Y(new_n12560_));
  AOI22X1  g12304(.A0(new_n2813_), .A1(\b[60] ), .B0(new_n2812_), .B1(\b[59] ), .Y(new_n12561_));
  OAI21X1  g12305(.A0(new_n2946_), .A1(new_n6930_), .B0(new_n12561_), .Y(new_n12562_));
  AOI21X1  g12306(.A0(new_n6951_), .A1(new_n2652_), .B0(new_n12562_), .Y(new_n12563_));
  XOR2X1   g12307(.A(new_n12563_), .B(\a[35] ), .Y(new_n12564_));
  XOR2X1   g12308(.A(new_n12564_), .B(new_n12560_), .Y(new_n12565_));
  INVX1    g12309(.A(new_n12565_), .Y(new_n12566_));
  AND2X1   g12310(.A(new_n12459_), .B(new_n12370_), .Y(new_n12567_));
  INVX1    g12311(.A(new_n12464_), .Y(new_n12568_));
  AOI21X1  g12312(.A0(new_n12568_), .A1(new_n12460_), .B0(new_n12567_), .Y(new_n12569_));
  XOR2X1   g12313(.A(new_n12569_), .B(new_n12566_), .Y(new_n12570_));
  NOR2X1   g12314(.A(new_n12367_), .B(new_n12363_), .Y(new_n12571_));
  INVX1    g12315(.A(new_n12571_), .Y(new_n12572_));
  OAI21X1  g12316(.A0(new_n12465_), .A1(new_n12368_), .B0(new_n12572_), .Y(new_n12573_));
  AOI22X1  g12317(.A0(new_n2545_), .A1(\b[63] ), .B0(new_n2544_), .B1(\b[62] ), .Y(new_n12574_));
  OAI21X1  g12318(.A0(new_n2543_), .A1(new_n7748_), .B0(new_n12574_), .Y(new_n12575_));
  AOI21X1  g12319(.A0(new_n7747_), .A1(new_n2260_), .B0(new_n12575_), .Y(new_n12576_));
  XOR2X1   g12320(.A(new_n12576_), .B(\a[32] ), .Y(new_n12577_));
  XOR2X1   g12321(.A(new_n12577_), .B(new_n12573_), .Y(new_n12578_));
  XOR2X1   g12322(.A(new_n12578_), .B(new_n12570_), .Y(new_n12579_));
  XOR2X1   g12323(.A(new_n12579_), .B(new_n12475_), .Y(new_n12580_));
  XOR2X1   g12324(.A(new_n12580_), .B(new_n12473_), .Y(\f[93] ));
  XOR2X1   g12325(.A(new_n12563_), .B(new_n2650_), .Y(new_n12582_));
  NOR2X1   g12326(.A(new_n12569_), .B(new_n12565_), .Y(new_n12583_));
  AOI21X1  g12327(.A0(new_n12582_), .A1(new_n12560_), .B0(new_n12583_), .Y(new_n12584_));
  OAI22X1  g12328(.A0(new_n2543_), .A1(new_n7745_), .B0(new_n2262_), .B1(new_n7772_), .Y(new_n12585_));
  AOI21X1  g12329(.A0(new_n7775_), .A1(new_n2260_), .B0(new_n12585_), .Y(new_n12586_));
  XOR2X1   g12330(.A(new_n12586_), .B(\a[32] ), .Y(new_n12587_));
  XOR2X1   g12331(.A(new_n12587_), .B(new_n12584_), .Y(new_n12588_));
  NOR2X1   g12332(.A(new_n12550_), .B(new_n12546_), .Y(new_n12589_));
  AOI21X1  g12333(.A0(new_n12551_), .A1(new_n12478_), .B0(new_n12589_), .Y(new_n12590_));
  INVX1    g12334(.A(new_n12590_), .Y(new_n12591_));
  XOR2X1   g12335(.A(new_n12507_), .B(new_n6019_), .Y(new_n12592_));
  NOR2X1   g12336(.A(new_n12512_), .B(new_n12509_), .Y(new_n12593_));
  AOI21X1  g12337(.A0(new_n12592_), .A1(new_n12504_), .B0(new_n12593_), .Y(new_n12594_));
  INVX1    g12338(.A(new_n12594_), .Y(new_n12595_));
  AOI22X1  g12339(.A0(new_n6438_), .A1(\b[40] ), .B0(new_n6437_), .B1(\b[39] ), .Y(new_n12596_));
  OAI21X1  g12340(.A0(new_n6436_), .A1(new_n3575_), .B0(new_n12596_), .Y(new_n12597_));
  AOI21X1  g12341(.A0(new_n6023_), .A1(new_n3574_), .B0(new_n12597_), .Y(new_n12598_));
  XOR2X1   g12342(.A(new_n12598_), .B(\a[56] ), .Y(new_n12599_));
  NOR2X1   g12343(.A(new_n12502_), .B(new_n12498_), .Y(new_n12600_));
  AOI21X1  g12344(.A0(new_n12503_), .A1(new_n12489_), .B0(new_n12600_), .Y(new_n12601_));
  AOI22X1  g12345(.A0(new_n6603_), .A1(\b[37] ), .B0(new_n6600_), .B1(\b[36] ), .Y(new_n12602_));
  OAI21X1  g12346(.A0(new_n6804_), .A1(new_n3156_), .B0(new_n12602_), .Y(new_n12603_));
  AOI21X1  g12347(.A0(new_n6598_), .A1(new_n3155_), .B0(new_n12603_), .Y(new_n12604_));
  XOR2X1   g12348(.A(new_n12604_), .B(\a[59] ), .Y(new_n12605_));
  NOR2X1   g12349(.A(new_n12492_), .B(new_n12415_), .Y(new_n12606_));
  INVX1    g12350(.A(new_n12497_), .Y(new_n12607_));
  AOI21X1  g12351(.A0(new_n12607_), .A1(new_n12493_), .B0(new_n12606_), .Y(new_n12608_));
  AOI22X1  g12352(.A0(new_n7818_), .A1(\b[30] ), .B0(new_n7817_), .B1(\b[31] ), .Y(new_n12609_));
  INVX1    g12353(.A(new_n12409_), .Y(new_n12610_));
  NOR2X1   g12354(.A(new_n12490_), .B(\a[29] ), .Y(new_n12611_));
  AOI21X1  g12355(.A0(new_n12491_), .A1(new_n12610_), .B0(new_n12611_), .Y(new_n12612_));
  XOR2X1   g12356(.A(new_n12612_), .B(new_n12609_), .Y(new_n12613_));
  AOI22X1  g12357(.A0(new_n7192_), .A1(\b[34] ), .B0(new_n7189_), .B1(\b[33] ), .Y(new_n12614_));
  OAI21X1  g12358(.A0(new_n7627_), .A1(new_n2612_), .B0(new_n12614_), .Y(new_n12615_));
  AOI21X1  g12359(.A0(new_n7187_), .A1(new_n2759_), .B0(new_n12615_), .Y(new_n12616_));
  XOR2X1   g12360(.A(new_n12616_), .B(\a[62] ), .Y(new_n12617_));
  XOR2X1   g12361(.A(new_n12617_), .B(new_n12613_), .Y(new_n12618_));
  XOR2X1   g12362(.A(new_n12618_), .B(new_n12608_), .Y(new_n12619_));
  XOR2X1   g12363(.A(new_n12619_), .B(new_n12605_), .Y(new_n12620_));
  XOR2X1   g12364(.A(new_n12620_), .B(new_n12601_), .Y(new_n12621_));
  XOR2X1   g12365(.A(new_n12621_), .B(new_n12599_), .Y(new_n12622_));
  XOR2X1   g12366(.A(new_n12622_), .B(new_n12595_), .Y(new_n12623_));
  AOI22X1  g12367(.A0(new_n5430_), .A1(\b[43] ), .B0(new_n5427_), .B1(\b[42] ), .Y(new_n12624_));
  OAI21X1  g12368(.A0(new_n5891_), .A1(new_n4015_), .B0(new_n12624_), .Y(new_n12625_));
  AOI21X1  g12369(.A0(new_n5425_), .A1(new_n4014_), .B0(new_n12625_), .Y(new_n12626_));
  XOR2X1   g12370(.A(new_n12626_), .B(\a[53] ), .Y(new_n12627_));
  XOR2X1   g12371(.A(new_n12627_), .B(new_n12623_), .Y(new_n12628_));
  INVX1    g12372(.A(new_n12513_), .Y(new_n12629_));
  NOR2X1   g12373(.A(new_n12517_), .B(new_n12629_), .Y(new_n12630_));
  INVX1    g12374(.A(new_n12518_), .Y(new_n12631_));
  AOI21X1  g12375(.A0(new_n12631_), .A1(new_n12487_), .B0(new_n12630_), .Y(new_n12632_));
  XOR2X1   g12376(.A(new_n12632_), .B(new_n12628_), .Y(new_n12633_));
  AOI22X1  g12377(.A0(new_n4880_), .A1(\b[46] ), .B0(new_n4877_), .B1(\b[45] ), .Y(new_n12634_));
  OAI21X1  g12378(.A0(new_n5291_), .A1(new_n4336_), .B0(new_n12634_), .Y(new_n12635_));
  AOI21X1  g12379(.A0(new_n4875_), .A1(new_n4509_), .B0(new_n12635_), .Y(new_n12636_));
  XOR2X1   g12380(.A(new_n12636_), .B(\a[50] ), .Y(new_n12637_));
  XOR2X1   g12381(.A(new_n12637_), .B(new_n12633_), .Y(new_n12638_));
  NOR2X1   g12382(.A(new_n12523_), .B(new_n12519_), .Y(new_n12639_));
  AOI21X1  g12383(.A0(new_n12524_), .A1(new_n12484_), .B0(new_n12639_), .Y(new_n12640_));
  XOR2X1   g12384(.A(new_n12640_), .B(new_n12638_), .Y(new_n12641_));
  AOI22X1  g12385(.A0(new_n4572_), .A1(\b[49] ), .B0(new_n4571_), .B1(\b[48] ), .Y(new_n12642_));
  OAI21X1  g12386(.A0(new_n4740_), .A1(new_n5039_), .B0(new_n12642_), .Y(new_n12643_));
  AOI21X1  g12387(.A0(new_n5038_), .A1(new_n4375_), .B0(new_n12643_), .Y(new_n12644_));
  XOR2X1   g12388(.A(new_n12644_), .B(\a[47] ), .Y(new_n12645_));
  XOR2X1   g12389(.A(new_n12645_), .B(new_n12641_), .Y(new_n12646_));
  INVX1    g12390(.A(new_n12529_), .Y(new_n12647_));
  NOR2X1   g12391(.A(new_n12533_), .B(new_n12530_), .Y(new_n12648_));
  AOI21X1  g12392(.A0(new_n12647_), .A1(new_n12525_), .B0(new_n12648_), .Y(new_n12649_));
  XOR2X1   g12393(.A(new_n12649_), .B(new_n12646_), .Y(new_n12650_));
  AOI22X1  g12394(.A0(new_n4095_), .A1(\b[52] ), .B0(new_n4094_), .B1(\b[51] ), .Y(new_n12651_));
  OAI21X1  g12395(.A0(new_n4233_), .A1(new_n5234_), .B0(new_n12651_), .Y(new_n12652_));
  AOI21X1  g12396(.A0(new_n5590_), .A1(new_n3901_), .B0(new_n12652_), .Y(new_n12653_));
  XOR2X1   g12397(.A(new_n12653_), .B(\a[44] ), .Y(new_n12654_));
  XOR2X1   g12398(.A(new_n12654_), .B(new_n12650_), .Y(new_n12655_));
  INVX1    g12399(.A(new_n12655_), .Y(new_n12656_));
  XOR2X1   g12400(.A(new_n12656_), .B(new_n12545_), .Y(new_n12657_));
  AOI22X1  g12401(.A0(new_n3652_), .A1(\b[55] ), .B0(new_n3651_), .B1(\b[54] ), .Y(new_n12658_));
  OAI21X1  g12402(.A0(new_n3778_), .A1(new_n6151_), .B0(new_n12658_), .Y(new_n12659_));
  AOI21X1  g12403(.A0(new_n6150_), .A1(new_n3480_), .B0(new_n12659_), .Y(new_n12660_));
  XOR2X1   g12404(.A(new_n12660_), .B(\a[41] ), .Y(new_n12661_));
  XOR2X1   g12405(.A(new_n12661_), .B(new_n12657_), .Y(new_n12662_));
  XOR2X1   g12406(.A(new_n12662_), .B(new_n12591_), .Y(new_n12663_));
  AOI22X1  g12407(.A0(new_n3204_), .A1(\b[58] ), .B0(new_n3203_), .B1(\b[57] ), .Y(new_n12664_));
  OAI21X1  g12408(.A0(new_n3321_), .A1(new_n6520_), .B0(new_n12664_), .Y(new_n12665_));
  AOI21X1  g12409(.A0(new_n6732_), .A1(new_n3080_), .B0(new_n12665_), .Y(new_n12666_));
  XOR2X1   g12410(.A(new_n12666_), .B(\a[38] ), .Y(new_n12667_));
  XOR2X1   g12411(.A(new_n12667_), .B(new_n12663_), .Y(new_n12668_));
  INVX1    g12412(.A(new_n12668_), .Y(new_n12669_));
  INVX1    g12413(.A(new_n12556_), .Y(new_n12670_));
  NOR2X1   g12414(.A(new_n12559_), .B(new_n12557_), .Y(new_n12671_));
  AOI21X1  g12415(.A0(new_n12670_), .A1(new_n12552_), .B0(new_n12671_), .Y(new_n12672_));
  XOR2X1   g12416(.A(new_n12672_), .B(new_n12669_), .Y(new_n12673_));
  AOI22X1  g12417(.A0(new_n2813_), .A1(\b[61] ), .B0(new_n2812_), .B1(\b[60] ), .Y(new_n12674_));
  OAI21X1  g12418(.A0(new_n2946_), .A1(new_n7339_), .B0(new_n12674_), .Y(new_n12675_));
  AOI21X1  g12419(.A0(new_n7338_), .A1(new_n2652_), .B0(new_n12675_), .Y(new_n12676_));
  XOR2X1   g12420(.A(new_n12676_), .B(\a[35] ), .Y(new_n12677_));
  XOR2X1   g12421(.A(new_n12677_), .B(new_n12673_), .Y(new_n12678_));
  XOR2X1   g12422(.A(new_n12678_), .B(new_n12588_), .Y(new_n12679_));
  INVX1    g12423(.A(new_n12577_), .Y(new_n12680_));
  NOR2X1   g12424(.A(new_n12578_), .B(new_n12570_), .Y(new_n12681_));
  AOI21X1  g12425(.A0(new_n12680_), .A1(new_n12573_), .B0(new_n12681_), .Y(new_n12682_));
  XOR2X1   g12426(.A(new_n12682_), .B(new_n12679_), .Y(new_n12683_));
  AND2X1   g12427(.A(new_n12579_), .B(new_n12475_), .Y(new_n12684_));
  INVX1    g12428(.A(new_n12684_), .Y(new_n12685_));
  OAI21X1  g12429(.A0(new_n12472_), .A1(new_n12471_), .B0(new_n12580_), .Y(new_n12686_));
  AND2X1   g12430(.A(new_n12686_), .B(new_n12685_), .Y(new_n12687_));
  XOR2X1   g12431(.A(new_n12687_), .B(new_n12683_), .Y(\f[94] ));
  INVX1    g12432(.A(new_n12679_), .Y(new_n12689_));
  NOR2X1   g12433(.A(new_n12682_), .B(new_n12689_), .Y(new_n12690_));
  AOI21X1  g12434(.A0(new_n12686_), .A1(new_n12685_), .B0(new_n12683_), .Y(new_n12691_));
  OR2X1    g12435(.A(new_n12691_), .B(new_n12690_), .Y(new_n12692_));
  NOR2X1   g12436(.A(new_n12587_), .B(new_n12584_), .Y(new_n12693_));
  AOI21X1  g12437(.A0(new_n12678_), .A1(new_n12588_), .B0(new_n12693_), .Y(new_n12694_));
  NOR2X1   g12438(.A(new_n12672_), .B(new_n12668_), .Y(new_n12695_));
  INVX1    g12439(.A(new_n12695_), .Y(new_n12696_));
  OAI21X1  g12440(.A0(new_n12677_), .A1(new_n12673_), .B0(new_n12696_), .Y(new_n12697_));
  AOI22X1  g12441(.A0(new_n7774_), .A1(new_n2260_), .B0(new_n2402_), .B1(\b[63] ), .Y(new_n12698_));
  XOR2X1   g12442(.A(new_n12698_), .B(\a[32] ), .Y(new_n12699_));
  XOR2X1   g12443(.A(new_n12699_), .B(new_n12697_), .Y(new_n12700_));
  OR2X1    g12444(.A(new_n12655_), .B(new_n12545_), .Y(new_n12701_));
  OAI21X1  g12445(.A0(new_n12661_), .A1(new_n12657_), .B0(new_n12701_), .Y(new_n12702_));
  AOI22X1  g12446(.A0(new_n3652_), .A1(\b[56] ), .B0(new_n3651_), .B1(\b[55] ), .Y(new_n12703_));
  OAI21X1  g12447(.A0(new_n3778_), .A1(new_n6148_), .B0(new_n12703_), .Y(new_n12704_));
  AOI21X1  g12448(.A0(new_n6342_), .A1(new_n3480_), .B0(new_n12704_), .Y(new_n12705_));
  XOR2X1   g12449(.A(new_n12705_), .B(new_n3478_), .Y(new_n12706_));
  AND2X1   g12450(.A(new_n12649_), .B(new_n12646_), .Y(new_n12707_));
  OR2X1    g12451(.A(new_n12649_), .B(new_n12646_), .Y(new_n12708_));
  OAI21X1  g12452(.A0(new_n12654_), .A1(new_n12707_), .B0(new_n12708_), .Y(new_n12709_));
  AOI22X1  g12453(.A0(new_n4095_), .A1(\b[53] ), .B0(new_n4094_), .B1(\b[52] ), .Y(new_n12710_));
  OAI21X1  g12454(.A0(new_n4233_), .A1(new_n5787_), .B0(new_n12710_), .Y(new_n12711_));
  AOI21X1  g12455(.A0(new_n5786_), .A1(new_n3901_), .B0(new_n12711_), .Y(new_n12712_));
  XOR2X1   g12456(.A(new_n12712_), .B(\a[44] ), .Y(new_n12713_));
  NOR2X1   g12457(.A(new_n12640_), .B(new_n12638_), .Y(new_n12714_));
  INVX1    g12458(.A(new_n12714_), .Y(new_n12715_));
  INVX1    g12459(.A(new_n12641_), .Y(new_n12716_));
  OAI21X1  g12460(.A0(new_n12645_), .A1(new_n12716_), .B0(new_n12715_), .Y(new_n12717_));
  INVX1    g12461(.A(new_n12717_), .Y(new_n12718_));
  AND2X1   g12462(.A(new_n12622_), .B(new_n12595_), .Y(new_n12719_));
  INVX1    g12463(.A(new_n12719_), .Y(new_n12720_));
  INVX1    g12464(.A(new_n12623_), .Y(new_n12721_));
  OAI21X1  g12465(.A0(new_n12627_), .A1(new_n12721_), .B0(new_n12720_), .Y(new_n12722_));
  AOI22X1  g12466(.A0(new_n5430_), .A1(\b[44] ), .B0(new_n5427_), .B1(\b[43] ), .Y(new_n12723_));
  OAI21X1  g12467(.A0(new_n5891_), .A1(new_n4012_), .B0(new_n12723_), .Y(new_n12724_));
  AOI21X1  g12468(.A0(new_n5425_), .A1(new_n4178_), .B0(new_n12724_), .Y(new_n12725_));
  XOR2X1   g12469(.A(new_n12725_), .B(new_n5423_), .Y(new_n12726_));
  AND2X1   g12470(.A(new_n12503_), .B(new_n12489_), .Y(new_n12727_));
  OAI21X1  g12471(.A0(new_n12727_), .A1(new_n12600_), .B0(new_n12620_), .Y(new_n12728_));
  OAI21X1  g12472(.A0(new_n12621_), .A1(new_n12599_), .B0(new_n12728_), .Y(new_n12729_));
  AOI22X1  g12473(.A0(new_n6438_), .A1(\b[41] ), .B0(new_n6437_), .B1(\b[40] ), .Y(new_n12730_));
  OAI21X1  g12474(.A0(new_n6436_), .A1(new_n3723_), .B0(new_n12730_), .Y(new_n12731_));
  AOI21X1  g12475(.A0(new_n6023_), .A1(new_n3722_), .B0(new_n12731_), .Y(new_n12732_));
  XOR2X1   g12476(.A(new_n12732_), .B(new_n6019_), .Y(new_n12733_));
  INVX1    g12477(.A(new_n12608_), .Y(new_n12734_));
  NOR2X1   g12478(.A(new_n12619_), .B(new_n12605_), .Y(new_n12735_));
  AOI21X1  g12479(.A0(new_n12618_), .A1(new_n12734_), .B0(new_n12735_), .Y(new_n12736_));
  INVX1    g12480(.A(new_n12609_), .Y(new_n12737_));
  NOR2X1   g12481(.A(new_n12612_), .B(new_n12737_), .Y(new_n12738_));
  INVX1    g12482(.A(new_n12738_), .Y(new_n12739_));
  OAI21X1  g12483(.A0(new_n12617_), .A1(new_n12613_), .B0(new_n12739_), .Y(new_n12740_));
  AOI22X1  g12484(.A0(new_n7818_), .A1(\b[31] ), .B0(new_n7817_), .B1(\b[32] ), .Y(new_n12741_));
  NOR2X1   g12485(.A(new_n12741_), .B(new_n12737_), .Y(new_n12742_));
  INVX1    g12486(.A(new_n12742_), .Y(new_n12743_));
  XOR2X1   g12487(.A(new_n12741_), .B(new_n12737_), .Y(new_n12744_));
  INVX1    g12488(.A(new_n12744_), .Y(new_n12745_));
  AND2X1   g12489(.A(new_n12741_), .B(new_n12737_), .Y(new_n12746_));
  AOI21X1  g12490(.A0(new_n12743_), .A1(new_n12740_), .B0(new_n12746_), .Y(new_n12747_));
  AOI22X1  g12491(.A0(new_n12747_), .A1(new_n12743_), .B0(new_n12745_), .B1(new_n12740_), .Y(new_n12748_));
  AOI22X1  g12492(.A0(new_n7192_), .A1(\b[35] ), .B0(new_n7189_), .B1(\b[34] ), .Y(new_n12749_));
  OAI21X1  g12493(.A0(new_n7627_), .A1(new_n2893_), .B0(new_n12749_), .Y(new_n12750_));
  AOI21X1  g12494(.A0(new_n7187_), .A1(new_n2892_), .B0(new_n12750_), .Y(new_n12751_));
  XOR2X1   g12495(.A(new_n12751_), .B(\a[62] ), .Y(new_n12752_));
  XOR2X1   g12496(.A(new_n12752_), .B(new_n12748_), .Y(new_n12753_));
  AOI22X1  g12497(.A0(new_n6603_), .A1(\b[38] ), .B0(new_n6600_), .B1(\b[37] ), .Y(new_n12754_));
  OAI21X1  g12498(.A0(new_n6804_), .A1(new_n3276_), .B0(new_n12754_), .Y(new_n12755_));
  AOI21X1  g12499(.A0(new_n6598_), .A1(new_n3275_), .B0(new_n12755_), .Y(new_n12756_));
  XOR2X1   g12500(.A(new_n12756_), .B(\a[59] ), .Y(new_n12757_));
  XOR2X1   g12501(.A(new_n12757_), .B(new_n12753_), .Y(new_n12758_));
  XOR2X1   g12502(.A(new_n12758_), .B(new_n12736_), .Y(new_n12759_));
  XOR2X1   g12503(.A(new_n12759_), .B(new_n12733_), .Y(new_n12760_));
  XOR2X1   g12504(.A(new_n12760_), .B(new_n12729_), .Y(new_n12761_));
  XOR2X1   g12505(.A(new_n12761_), .B(new_n12726_), .Y(new_n12762_));
  XOR2X1   g12506(.A(new_n12762_), .B(new_n12722_), .Y(new_n12763_));
  AOI22X1  g12507(.A0(new_n4880_), .A1(\b[47] ), .B0(new_n4877_), .B1(\b[46] ), .Y(new_n12764_));
  OAI21X1  g12508(.A0(new_n5291_), .A1(new_n4674_), .B0(new_n12764_), .Y(new_n12765_));
  AOI21X1  g12509(.A0(new_n4875_), .A1(new_n4673_), .B0(new_n12765_), .Y(new_n12766_));
  XOR2X1   g12510(.A(new_n12766_), .B(\a[50] ), .Y(new_n12767_));
  XOR2X1   g12511(.A(new_n12767_), .B(new_n12763_), .Y(new_n12768_));
  INVX1    g12512(.A(new_n12768_), .Y(new_n12769_));
  NOR2X1   g12513(.A(new_n12632_), .B(new_n12628_), .Y(new_n12770_));
  INVX1    g12514(.A(new_n12637_), .Y(new_n12771_));
  AOI21X1  g12515(.A0(new_n12771_), .A1(new_n12633_), .B0(new_n12770_), .Y(new_n12772_));
  XOR2X1   g12516(.A(new_n12772_), .B(new_n12769_), .Y(new_n12773_));
  AOI22X1  g12517(.A0(new_n4572_), .A1(\b[50] ), .B0(new_n4571_), .B1(\b[49] ), .Y(new_n12774_));
  OAI21X1  g12518(.A0(new_n4740_), .A1(new_n5036_), .B0(new_n12774_), .Y(new_n12775_));
  AOI21X1  g12519(.A0(new_n5204_), .A1(new_n4375_), .B0(new_n12775_), .Y(new_n12776_));
  XOR2X1   g12520(.A(new_n12776_), .B(\a[47] ), .Y(new_n12777_));
  XOR2X1   g12521(.A(new_n12777_), .B(new_n12773_), .Y(new_n12778_));
  XOR2X1   g12522(.A(new_n12778_), .B(new_n12718_), .Y(new_n12779_));
  XOR2X1   g12523(.A(new_n12779_), .B(new_n12713_), .Y(new_n12780_));
  XOR2X1   g12524(.A(new_n12780_), .B(new_n12709_), .Y(new_n12781_));
  XOR2X1   g12525(.A(new_n12781_), .B(new_n12706_), .Y(new_n12782_));
  XOR2X1   g12526(.A(new_n12782_), .B(new_n12702_), .Y(new_n12783_));
  AOI22X1  g12527(.A0(new_n3204_), .A1(\b[59] ), .B0(new_n3203_), .B1(\b[58] ), .Y(new_n12784_));
  OAI21X1  g12528(.A0(new_n3321_), .A1(new_n6933_), .B0(new_n12784_), .Y(new_n12785_));
  AOI21X1  g12529(.A0(new_n6932_), .A1(new_n3080_), .B0(new_n12785_), .Y(new_n12786_));
  XOR2X1   g12530(.A(new_n12786_), .B(\a[38] ), .Y(new_n12787_));
  XOR2X1   g12531(.A(new_n12787_), .B(new_n12783_), .Y(new_n12788_));
  AND2X1   g12532(.A(new_n12662_), .B(new_n12591_), .Y(new_n12789_));
  INVX1    g12533(.A(new_n12667_), .Y(new_n12790_));
  AOI21X1  g12534(.A0(new_n12790_), .A1(new_n12663_), .B0(new_n12789_), .Y(new_n12791_));
  XOR2X1   g12535(.A(new_n12791_), .B(new_n12788_), .Y(new_n12792_));
  AOI22X1  g12536(.A0(new_n2813_), .A1(\b[62] ), .B0(new_n2812_), .B1(\b[61] ), .Y(new_n12793_));
  OAI21X1  g12537(.A0(new_n2946_), .A1(new_n7559_), .B0(new_n12793_), .Y(new_n12794_));
  AOI21X1  g12538(.A0(new_n7558_), .A1(new_n2652_), .B0(new_n12794_), .Y(new_n12795_));
  XOR2X1   g12539(.A(new_n12795_), .B(\a[35] ), .Y(new_n12796_));
  XOR2X1   g12540(.A(new_n12796_), .B(new_n12792_), .Y(new_n12797_));
  INVX1    g12541(.A(new_n12797_), .Y(new_n12798_));
  XOR2X1   g12542(.A(new_n12798_), .B(new_n12700_), .Y(new_n12799_));
  XOR2X1   g12543(.A(new_n12799_), .B(new_n12694_), .Y(new_n12800_));
  XOR2X1   g12544(.A(new_n12800_), .B(new_n12692_), .Y(\f[95] ));
  NOR2X1   g12545(.A(new_n12799_), .B(new_n12694_), .Y(new_n12802_));
  INVX1    g12546(.A(new_n12802_), .Y(new_n12803_));
  OAI21X1  g12547(.A0(new_n12691_), .A1(new_n12690_), .B0(new_n12800_), .Y(new_n12804_));
  NAND2X1  g12548(.A(new_n12804_), .B(new_n12803_), .Y(new_n12805_));
  XOR2X1   g12549(.A(new_n12698_), .B(new_n2258_), .Y(new_n12806_));
  NOR2X1   g12550(.A(new_n12797_), .B(new_n12700_), .Y(new_n12807_));
  AOI21X1  g12551(.A0(new_n12806_), .A1(new_n12697_), .B0(new_n12807_), .Y(new_n12808_));
  INVX1    g12552(.A(new_n12808_), .Y(new_n12809_));
  AND2X1   g12553(.A(new_n12778_), .B(new_n12717_), .Y(new_n12810_));
  INVX1    g12554(.A(new_n12810_), .Y(new_n12811_));
  OAI21X1  g12555(.A0(new_n12779_), .A1(new_n12713_), .B0(new_n12811_), .Y(new_n12812_));
  NOR2X1   g12556(.A(new_n12772_), .B(new_n12768_), .Y(new_n12813_));
  INVX1    g12557(.A(new_n12813_), .Y(new_n12814_));
  OAI21X1  g12558(.A0(new_n12777_), .A1(new_n12773_), .B0(new_n12814_), .Y(new_n12815_));
  NOR2X1   g12559(.A(new_n12752_), .B(new_n12748_), .Y(new_n12816_));
  INVX1    g12560(.A(new_n12757_), .Y(new_n12817_));
  AOI21X1  g12561(.A0(new_n12817_), .A1(new_n12753_), .B0(new_n12816_), .Y(new_n12818_));
  INVX1    g12562(.A(new_n12818_), .Y(new_n12819_));
  AOI22X1  g12563(.A0(new_n7818_), .A1(\b[32] ), .B0(new_n7817_), .B1(\b[33] ), .Y(new_n12820_));
  XOR2X1   g12564(.A(new_n12820_), .B(\a[32] ), .Y(new_n12821_));
  XOR2X1   g12565(.A(new_n12821_), .B(new_n12741_), .Y(new_n12822_));
  XOR2X1   g12566(.A(new_n12822_), .B(new_n12747_), .Y(new_n12823_));
  AOI22X1  g12567(.A0(new_n7192_), .A1(\b[36] ), .B0(new_n7189_), .B1(\b[35] ), .Y(new_n12824_));
  OAI21X1  g12568(.A0(new_n7627_), .A1(new_n2890_), .B0(new_n12824_), .Y(new_n12825_));
  AOI21X1  g12569(.A0(new_n7187_), .A1(new_n3015_), .B0(new_n12825_), .Y(new_n12826_));
  XOR2X1   g12570(.A(new_n12826_), .B(\a[62] ), .Y(new_n12827_));
  XOR2X1   g12571(.A(new_n12827_), .B(new_n12823_), .Y(new_n12828_));
  AOI22X1  g12572(.A0(new_n6603_), .A1(\b[39] ), .B0(new_n6600_), .B1(\b[38] ), .Y(new_n12829_));
  OAI21X1  g12573(.A0(new_n6804_), .A1(new_n3413_), .B0(new_n12829_), .Y(new_n12830_));
  AOI21X1  g12574(.A0(new_n6598_), .A1(new_n3412_), .B0(new_n12830_), .Y(new_n12831_));
  XOR2X1   g12575(.A(new_n12831_), .B(\a[59] ), .Y(new_n12832_));
  XOR2X1   g12576(.A(new_n12832_), .B(new_n12828_), .Y(new_n12833_));
  XOR2X1   g12577(.A(new_n12833_), .B(new_n12819_), .Y(new_n12834_));
  AOI22X1  g12578(.A0(new_n6438_), .A1(\b[42] ), .B0(new_n6437_), .B1(\b[41] ), .Y(new_n12835_));
  OAI21X1  g12579(.A0(new_n6436_), .A1(new_n3720_), .B0(new_n12835_), .Y(new_n12836_));
  AOI21X1  g12580(.A0(new_n6023_), .A1(new_n3860_), .B0(new_n12836_), .Y(new_n12837_));
  XOR2X1   g12581(.A(new_n12837_), .B(\a[56] ), .Y(new_n12838_));
  XOR2X1   g12582(.A(new_n12838_), .B(new_n12834_), .Y(new_n12839_));
  NOR2X1   g12583(.A(new_n12758_), .B(new_n12736_), .Y(new_n12840_));
  AOI21X1  g12584(.A0(new_n12759_), .A1(new_n12733_), .B0(new_n12840_), .Y(new_n12841_));
  XOR2X1   g12585(.A(new_n12841_), .B(new_n12839_), .Y(new_n12842_));
  AOI22X1  g12586(.A0(new_n5430_), .A1(\b[45] ), .B0(new_n5427_), .B1(\b[44] ), .Y(new_n12843_));
  OAI21X1  g12587(.A0(new_n5891_), .A1(new_n4339_), .B0(new_n12843_), .Y(new_n12844_));
  AOI21X1  g12588(.A0(new_n5425_), .A1(new_n4338_), .B0(new_n12844_), .Y(new_n12845_));
  XOR2X1   g12589(.A(new_n12845_), .B(\a[53] ), .Y(new_n12846_));
  XOR2X1   g12590(.A(new_n12846_), .B(new_n12842_), .Y(new_n12847_));
  AND2X1   g12591(.A(new_n12760_), .B(new_n12729_), .Y(new_n12848_));
  AOI21X1  g12592(.A0(new_n12761_), .A1(new_n12726_), .B0(new_n12848_), .Y(new_n12849_));
  XOR2X1   g12593(.A(new_n12849_), .B(new_n12847_), .Y(new_n12850_));
  AOI22X1  g12594(.A0(new_n4880_), .A1(\b[48] ), .B0(new_n4877_), .B1(\b[47] ), .Y(new_n12851_));
  OAI21X1  g12595(.A0(new_n5291_), .A1(new_n4693_), .B0(new_n12851_), .Y(new_n12852_));
  AOI21X1  g12596(.A0(new_n4875_), .A1(new_n4692_), .B0(new_n12852_), .Y(new_n12853_));
  XOR2X1   g12597(.A(new_n12853_), .B(\a[50] ), .Y(new_n12854_));
  XOR2X1   g12598(.A(new_n12854_), .B(new_n12850_), .Y(new_n12855_));
  AND2X1   g12599(.A(new_n12762_), .B(new_n12722_), .Y(new_n12856_));
  INVX1    g12600(.A(new_n12767_), .Y(new_n12857_));
  AOI21X1  g12601(.A0(new_n12857_), .A1(new_n12763_), .B0(new_n12856_), .Y(new_n12858_));
  XOR2X1   g12602(.A(new_n12858_), .B(new_n12855_), .Y(new_n12859_));
  INVX1    g12603(.A(new_n12859_), .Y(new_n12860_));
  AOI22X1  g12604(.A0(new_n4572_), .A1(\b[51] ), .B0(new_n4571_), .B1(\b[50] ), .Y(new_n12861_));
  OAI21X1  g12605(.A0(new_n4740_), .A1(new_n5237_), .B0(new_n12861_), .Y(new_n12862_));
  AOI21X1  g12606(.A0(new_n5236_), .A1(new_n4375_), .B0(new_n12862_), .Y(new_n12863_));
  XOR2X1   g12607(.A(new_n12863_), .B(\a[47] ), .Y(new_n12864_));
  AND2X1   g12608(.A(new_n12864_), .B(new_n12860_), .Y(new_n12865_));
  INVX1    g12609(.A(new_n12865_), .Y(new_n12866_));
  OAI21X1  g12610(.A0(new_n12864_), .A1(new_n12860_), .B0(new_n12815_), .Y(new_n12867_));
  OR2X1    g12611(.A(new_n12867_), .B(new_n12865_), .Y(new_n12868_));
  NOR2X1   g12612(.A(new_n12864_), .B(new_n12860_), .Y(new_n12869_));
  AOI21X1  g12613(.A0(new_n12866_), .A1(new_n12815_), .B0(new_n12869_), .Y(new_n12870_));
  AOI22X1  g12614(.A0(new_n12870_), .A1(new_n12866_), .B0(new_n12868_), .B1(new_n12815_), .Y(new_n12871_));
  AOI22X1  g12615(.A0(new_n4095_), .A1(\b[54] ), .B0(new_n4094_), .B1(\b[53] ), .Y(new_n12872_));
  OAI21X1  g12616(.A0(new_n4233_), .A1(new_n5808_), .B0(new_n12872_), .Y(new_n12873_));
  AOI21X1  g12617(.A0(new_n5807_), .A1(new_n3901_), .B0(new_n12873_), .Y(new_n12874_));
  XOR2X1   g12618(.A(new_n12874_), .B(\a[44] ), .Y(new_n12875_));
  XOR2X1   g12619(.A(new_n12875_), .B(new_n12871_), .Y(new_n12876_));
  XOR2X1   g12620(.A(new_n12876_), .B(new_n12812_), .Y(new_n12877_));
  AOI22X1  g12621(.A0(new_n3652_), .A1(\b[57] ), .B0(new_n3651_), .B1(\b[56] ), .Y(new_n12878_));
  OAI21X1  g12622(.A0(new_n3778_), .A1(new_n6523_), .B0(new_n12878_), .Y(new_n12879_));
  AOI21X1  g12623(.A0(new_n6522_), .A1(new_n3480_), .B0(new_n12879_), .Y(new_n12880_));
  XOR2X1   g12624(.A(new_n12880_), .B(\a[41] ), .Y(new_n12881_));
  XOR2X1   g12625(.A(new_n12881_), .B(new_n12877_), .Y(new_n12882_));
  AND2X1   g12626(.A(new_n12780_), .B(new_n12709_), .Y(new_n12883_));
  AOI21X1  g12627(.A0(new_n12781_), .A1(new_n12706_), .B0(new_n12883_), .Y(new_n12884_));
  XOR2X1   g12628(.A(new_n12884_), .B(new_n12882_), .Y(new_n12885_));
  AOI22X1  g12629(.A0(new_n3204_), .A1(\b[60] ), .B0(new_n3203_), .B1(\b[59] ), .Y(new_n12886_));
  OAI21X1  g12630(.A0(new_n3321_), .A1(new_n6930_), .B0(new_n12886_), .Y(new_n12887_));
  AOI21X1  g12631(.A0(new_n6951_), .A1(new_n3080_), .B0(new_n12887_), .Y(new_n12888_));
  XOR2X1   g12632(.A(new_n12888_), .B(\a[38] ), .Y(new_n12889_));
  XOR2X1   g12633(.A(new_n12889_), .B(new_n12885_), .Y(new_n12890_));
  INVX1    g12634(.A(new_n12890_), .Y(new_n12891_));
  AND2X1   g12635(.A(new_n12782_), .B(new_n12702_), .Y(new_n12892_));
  INVX1    g12636(.A(new_n12787_), .Y(new_n12893_));
  AOI21X1  g12637(.A0(new_n12893_), .A1(new_n12783_), .B0(new_n12892_), .Y(new_n12894_));
  XOR2X1   g12638(.A(new_n12894_), .B(new_n12891_), .Y(new_n12895_));
  NOR2X1   g12639(.A(new_n12791_), .B(new_n12788_), .Y(new_n12896_));
  INVX1    g12640(.A(new_n12896_), .Y(new_n12897_));
  INVX1    g12641(.A(new_n12792_), .Y(new_n12898_));
  OAI21X1  g12642(.A0(new_n12796_), .A1(new_n12898_), .B0(new_n12897_), .Y(new_n12899_));
  AOI22X1  g12643(.A0(new_n2813_), .A1(\b[63] ), .B0(new_n2812_), .B1(\b[62] ), .Y(new_n12900_));
  OAI21X1  g12644(.A0(new_n2946_), .A1(new_n7748_), .B0(new_n12900_), .Y(new_n12901_));
  AOI21X1  g12645(.A0(new_n7747_), .A1(new_n2652_), .B0(new_n12901_), .Y(new_n12902_));
  XOR2X1   g12646(.A(new_n12902_), .B(\a[35] ), .Y(new_n12903_));
  XOR2X1   g12647(.A(new_n12903_), .B(new_n12899_), .Y(new_n12904_));
  XOR2X1   g12648(.A(new_n12904_), .B(new_n12895_), .Y(new_n12905_));
  XOR2X1   g12649(.A(new_n12905_), .B(new_n12809_), .Y(new_n12906_));
  XOR2X1   g12650(.A(new_n12906_), .B(new_n12805_), .Y(\f[96] ));
  XOR2X1   g12651(.A(new_n12888_), .B(new_n3078_), .Y(new_n12908_));
  NOR2X1   g12652(.A(new_n12894_), .B(new_n12890_), .Y(new_n12909_));
  AOI21X1  g12653(.A0(new_n12908_), .A1(new_n12885_), .B0(new_n12909_), .Y(new_n12910_));
  OAI22X1  g12654(.A0(new_n2946_), .A1(new_n7745_), .B0(new_n2654_), .B1(new_n7772_), .Y(new_n12911_));
  AOI21X1  g12655(.A0(new_n7775_), .A1(new_n2652_), .B0(new_n12911_), .Y(new_n12912_));
  XOR2X1   g12656(.A(new_n12912_), .B(\a[35] ), .Y(new_n12913_));
  XOR2X1   g12657(.A(new_n12913_), .B(new_n12910_), .Y(new_n12914_));
  NOR2X1   g12658(.A(new_n12875_), .B(new_n12871_), .Y(new_n12915_));
  AOI21X1  g12659(.A0(new_n12876_), .A1(new_n12812_), .B0(new_n12915_), .Y(new_n12916_));
  INVX1    g12660(.A(new_n12916_), .Y(new_n12917_));
  NOR2X1   g12661(.A(new_n12832_), .B(new_n12828_), .Y(new_n12918_));
  AOI21X1  g12662(.A0(new_n12833_), .A1(new_n12819_), .B0(new_n12918_), .Y(new_n12919_));
  INVX1    g12663(.A(new_n12919_), .Y(new_n12920_));
  AOI22X1  g12664(.A0(new_n6603_), .A1(\b[40] ), .B0(new_n6600_), .B1(\b[39] ), .Y(new_n12921_));
  OAI21X1  g12665(.A0(new_n6804_), .A1(new_n3575_), .B0(new_n12921_), .Y(new_n12922_));
  AOI21X1  g12666(.A0(new_n6598_), .A1(new_n3574_), .B0(new_n12922_), .Y(new_n12923_));
  XOR2X1   g12667(.A(new_n12923_), .B(\a[59] ), .Y(new_n12924_));
  NOR2X1   g12668(.A(new_n12822_), .B(new_n12747_), .Y(new_n12925_));
  INVX1    g12669(.A(new_n12827_), .Y(new_n12926_));
  AOI21X1  g12670(.A0(new_n12926_), .A1(new_n12823_), .B0(new_n12925_), .Y(new_n12927_));
  AOI22X1  g12671(.A0(new_n7818_), .A1(\b[33] ), .B0(new_n7817_), .B1(\b[34] ), .Y(new_n12928_));
  INVX1    g12672(.A(new_n12741_), .Y(new_n12929_));
  NOR2X1   g12673(.A(new_n12820_), .B(\a[32] ), .Y(new_n12930_));
  AOI21X1  g12674(.A0(new_n12821_), .A1(new_n12929_), .B0(new_n12930_), .Y(new_n12931_));
  XOR2X1   g12675(.A(new_n12931_), .B(new_n12928_), .Y(new_n12932_));
  AOI22X1  g12676(.A0(new_n7192_), .A1(\b[37] ), .B0(new_n7189_), .B1(\b[36] ), .Y(new_n12933_));
  OAI21X1  g12677(.A0(new_n7627_), .A1(new_n3156_), .B0(new_n12933_), .Y(new_n12934_));
  AOI21X1  g12678(.A0(new_n7187_), .A1(new_n3155_), .B0(new_n12934_), .Y(new_n12935_));
  XOR2X1   g12679(.A(new_n12935_), .B(\a[62] ), .Y(new_n12936_));
  XOR2X1   g12680(.A(new_n12936_), .B(new_n12932_), .Y(new_n12937_));
  XOR2X1   g12681(.A(new_n12937_), .B(new_n12927_), .Y(new_n12938_));
  XOR2X1   g12682(.A(new_n12938_), .B(new_n12924_), .Y(new_n12939_));
  XOR2X1   g12683(.A(new_n12939_), .B(new_n12920_), .Y(new_n12940_));
  AOI22X1  g12684(.A0(new_n6438_), .A1(\b[43] ), .B0(new_n6437_), .B1(\b[42] ), .Y(new_n12941_));
  OAI21X1  g12685(.A0(new_n6436_), .A1(new_n4015_), .B0(new_n12941_), .Y(new_n12942_));
  AOI21X1  g12686(.A0(new_n6023_), .A1(new_n4014_), .B0(new_n12942_), .Y(new_n12943_));
  XOR2X1   g12687(.A(new_n12943_), .B(\a[56] ), .Y(new_n12944_));
  XOR2X1   g12688(.A(new_n12944_), .B(new_n12940_), .Y(new_n12945_));
  INVX1    g12689(.A(new_n12838_), .Y(new_n12946_));
  NOR2X1   g12690(.A(new_n12841_), .B(new_n12839_), .Y(new_n12947_));
  AOI21X1  g12691(.A0(new_n12946_), .A1(new_n12834_), .B0(new_n12947_), .Y(new_n12948_));
  XOR2X1   g12692(.A(new_n12948_), .B(new_n12945_), .Y(new_n12949_));
  AOI22X1  g12693(.A0(new_n5430_), .A1(\b[46] ), .B0(new_n5427_), .B1(\b[45] ), .Y(new_n12950_));
  OAI21X1  g12694(.A0(new_n5891_), .A1(new_n4336_), .B0(new_n12950_), .Y(new_n12951_));
  AOI21X1  g12695(.A0(new_n5425_), .A1(new_n4509_), .B0(new_n12951_), .Y(new_n12952_));
  XOR2X1   g12696(.A(new_n12952_), .B(\a[53] ), .Y(new_n12953_));
  XOR2X1   g12697(.A(new_n12953_), .B(new_n12949_), .Y(new_n12954_));
  INVX1    g12698(.A(new_n12846_), .Y(new_n12955_));
  NOR2X1   g12699(.A(new_n12849_), .B(new_n12847_), .Y(new_n12956_));
  AOI21X1  g12700(.A0(new_n12955_), .A1(new_n12842_), .B0(new_n12956_), .Y(new_n12957_));
  XOR2X1   g12701(.A(new_n12957_), .B(new_n12954_), .Y(new_n12958_));
  AOI22X1  g12702(.A0(new_n4880_), .A1(\b[49] ), .B0(new_n4877_), .B1(\b[48] ), .Y(new_n12959_));
  OAI21X1  g12703(.A0(new_n5291_), .A1(new_n5039_), .B0(new_n12959_), .Y(new_n12960_));
  AOI21X1  g12704(.A0(new_n5038_), .A1(new_n4875_), .B0(new_n12960_), .Y(new_n12961_));
  XOR2X1   g12705(.A(new_n12961_), .B(\a[50] ), .Y(new_n12962_));
  XOR2X1   g12706(.A(new_n12962_), .B(new_n12958_), .Y(new_n12963_));
  INVX1    g12707(.A(new_n12854_), .Y(new_n12964_));
  NOR2X1   g12708(.A(new_n12858_), .B(new_n12855_), .Y(new_n12965_));
  AOI21X1  g12709(.A0(new_n12964_), .A1(new_n12850_), .B0(new_n12965_), .Y(new_n12966_));
  XOR2X1   g12710(.A(new_n12966_), .B(new_n12963_), .Y(new_n12967_));
  AOI22X1  g12711(.A0(new_n4572_), .A1(\b[52] ), .B0(new_n4571_), .B1(\b[51] ), .Y(new_n12968_));
  OAI21X1  g12712(.A0(new_n4740_), .A1(new_n5234_), .B0(new_n12968_), .Y(new_n12969_));
  AOI21X1  g12713(.A0(new_n5590_), .A1(new_n4375_), .B0(new_n12969_), .Y(new_n12970_));
  XOR2X1   g12714(.A(new_n12970_), .B(\a[47] ), .Y(new_n12971_));
  XOR2X1   g12715(.A(new_n12971_), .B(new_n12967_), .Y(new_n12972_));
  INVX1    g12716(.A(new_n12972_), .Y(new_n12973_));
  XOR2X1   g12717(.A(new_n12973_), .B(new_n12870_), .Y(new_n12974_));
  AOI22X1  g12718(.A0(new_n4095_), .A1(\b[55] ), .B0(new_n4094_), .B1(\b[54] ), .Y(new_n12975_));
  OAI21X1  g12719(.A0(new_n4233_), .A1(new_n6151_), .B0(new_n12975_), .Y(new_n12976_));
  AOI21X1  g12720(.A0(new_n6150_), .A1(new_n3901_), .B0(new_n12976_), .Y(new_n12977_));
  XOR2X1   g12721(.A(new_n12977_), .B(\a[44] ), .Y(new_n12978_));
  XOR2X1   g12722(.A(new_n12978_), .B(new_n12974_), .Y(new_n12979_));
  XOR2X1   g12723(.A(new_n12979_), .B(new_n12917_), .Y(new_n12980_));
  AOI22X1  g12724(.A0(new_n3652_), .A1(\b[58] ), .B0(new_n3651_), .B1(\b[57] ), .Y(new_n12981_));
  OAI21X1  g12725(.A0(new_n3778_), .A1(new_n6520_), .B0(new_n12981_), .Y(new_n12982_));
  AOI21X1  g12726(.A0(new_n6732_), .A1(new_n3480_), .B0(new_n12982_), .Y(new_n12983_));
  XOR2X1   g12727(.A(new_n12983_), .B(\a[41] ), .Y(new_n12984_));
  XOR2X1   g12728(.A(new_n12984_), .B(new_n12980_), .Y(new_n12985_));
  INVX1    g12729(.A(new_n12985_), .Y(new_n12986_));
  INVX1    g12730(.A(new_n12881_), .Y(new_n12987_));
  NOR2X1   g12731(.A(new_n12884_), .B(new_n12882_), .Y(new_n12988_));
  AOI21X1  g12732(.A0(new_n12987_), .A1(new_n12877_), .B0(new_n12988_), .Y(new_n12989_));
  XOR2X1   g12733(.A(new_n12989_), .B(new_n12986_), .Y(new_n12990_));
  AOI22X1  g12734(.A0(new_n3204_), .A1(\b[61] ), .B0(new_n3203_), .B1(\b[60] ), .Y(new_n12991_));
  OAI21X1  g12735(.A0(new_n3321_), .A1(new_n7339_), .B0(new_n12991_), .Y(new_n12992_));
  AOI21X1  g12736(.A0(new_n7338_), .A1(new_n3080_), .B0(new_n12992_), .Y(new_n12993_));
  XOR2X1   g12737(.A(new_n12993_), .B(\a[38] ), .Y(new_n12994_));
  XOR2X1   g12738(.A(new_n12994_), .B(new_n12990_), .Y(new_n12995_));
  XOR2X1   g12739(.A(new_n12995_), .B(new_n12914_), .Y(new_n12996_));
  INVX1    g12740(.A(new_n12903_), .Y(new_n12997_));
  NOR2X1   g12741(.A(new_n12904_), .B(new_n12895_), .Y(new_n12998_));
  AOI21X1  g12742(.A0(new_n12997_), .A1(new_n12899_), .B0(new_n12998_), .Y(new_n12999_));
  XOR2X1   g12743(.A(new_n12999_), .B(new_n12996_), .Y(new_n13000_));
  AND2X1   g12744(.A(new_n12905_), .B(new_n12809_), .Y(new_n13001_));
  INVX1    g12745(.A(new_n12906_), .Y(new_n13002_));
  AOI21X1  g12746(.A0(new_n12804_), .A1(new_n12803_), .B0(new_n13002_), .Y(new_n13003_));
  NOR2X1   g12747(.A(new_n13003_), .B(new_n13001_), .Y(new_n13004_));
  XOR2X1   g12748(.A(new_n13004_), .B(new_n13000_), .Y(\f[97] ));
  INVX1    g12749(.A(new_n12996_), .Y(new_n13006_));
  NOR2X1   g12750(.A(new_n12999_), .B(new_n13006_), .Y(new_n13007_));
  INVX1    g12751(.A(new_n13007_), .Y(new_n13008_));
  INVX1    g12752(.A(new_n13000_), .Y(new_n13009_));
  OAI21X1  g12753(.A0(new_n13003_), .A1(new_n13001_), .B0(new_n13009_), .Y(new_n13010_));
  NAND2X1  g12754(.A(new_n13010_), .B(new_n13008_), .Y(new_n13011_));
  NOR2X1   g12755(.A(new_n12913_), .B(new_n12910_), .Y(new_n13012_));
  AOI21X1  g12756(.A0(new_n12995_), .A1(new_n12914_), .B0(new_n13012_), .Y(new_n13013_));
  OR2X1    g12757(.A(new_n12989_), .B(new_n12985_), .Y(new_n13014_));
  OR2X1    g12758(.A(new_n12994_), .B(new_n12990_), .Y(new_n13015_));
  AND2X1   g12759(.A(new_n13015_), .B(new_n13014_), .Y(new_n13016_));
  NOR3X1   g12760(.A(new_n2945_), .B(new_n2651_), .C(new_n7772_), .Y(new_n13017_));
  AOI21X1  g12761(.A0(new_n7774_), .A1(new_n2652_), .B0(new_n13017_), .Y(new_n13018_));
  XOR2X1   g12762(.A(new_n13018_), .B(\a[35] ), .Y(new_n13019_));
  XOR2X1   g12763(.A(new_n13019_), .B(new_n13016_), .Y(new_n13020_));
  OR2X1    g12764(.A(new_n12972_), .B(new_n12870_), .Y(new_n13021_));
  OAI21X1  g12765(.A0(new_n12978_), .A1(new_n12974_), .B0(new_n13021_), .Y(new_n13022_));
  AOI22X1  g12766(.A0(new_n4095_), .A1(\b[56] ), .B0(new_n4094_), .B1(\b[55] ), .Y(new_n13023_));
  OAI21X1  g12767(.A0(new_n4233_), .A1(new_n6148_), .B0(new_n13023_), .Y(new_n13024_));
  AOI21X1  g12768(.A0(new_n6342_), .A1(new_n3901_), .B0(new_n13024_), .Y(new_n13025_));
  XOR2X1   g12769(.A(new_n13025_), .B(new_n3899_), .Y(new_n13026_));
  AND2X1   g12770(.A(new_n12966_), .B(new_n12963_), .Y(new_n13027_));
  OR2X1    g12771(.A(new_n12966_), .B(new_n12963_), .Y(new_n13028_));
  OAI21X1  g12772(.A0(new_n12971_), .A1(new_n13027_), .B0(new_n13028_), .Y(new_n13029_));
  AOI22X1  g12773(.A0(new_n4572_), .A1(\b[53] ), .B0(new_n4571_), .B1(\b[52] ), .Y(new_n13030_));
  OAI21X1  g12774(.A0(new_n4740_), .A1(new_n5787_), .B0(new_n13030_), .Y(new_n13031_));
  AOI21X1  g12775(.A0(new_n5786_), .A1(new_n4375_), .B0(new_n13031_), .Y(new_n13032_));
  XOR2X1   g12776(.A(new_n13032_), .B(\a[47] ), .Y(new_n13033_));
  NOR2X1   g12777(.A(new_n12957_), .B(new_n12954_), .Y(new_n13034_));
  INVX1    g12778(.A(new_n13034_), .Y(new_n13035_));
  INVX1    g12779(.A(new_n12958_), .Y(new_n13036_));
  OAI21X1  g12780(.A0(new_n12962_), .A1(new_n13036_), .B0(new_n13035_), .Y(new_n13037_));
  INVX1    g12781(.A(new_n13037_), .Y(new_n13038_));
  AND2X1   g12782(.A(new_n12939_), .B(new_n12920_), .Y(new_n13039_));
  INVX1    g12783(.A(new_n13039_), .Y(new_n13040_));
  INVX1    g12784(.A(new_n12940_), .Y(new_n13041_));
  OAI21X1  g12785(.A0(new_n12944_), .A1(new_n13041_), .B0(new_n13040_), .Y(new_n13042_));
  AOI22X1  g12786(.A0(new_n6438_), .A1(\b[44] ), .B0(new_n6437_), .B1(\b[43] ), .Y(new_n13043_));
  OAI21X1  g12787(.A0(new_n6436_), .A1(new_n4012_), .B0(new_n13043_), .Y(new_n13044_));
  AOI21X1  g12788(.A0(new_n6023_), .A1(new_n4178_), .B0(new_n13044_), .Y(new_n13045_));
  XOR2X1   g12789(.A(new_n13045_), .B(new_n6019_), .Y(new_n13046_));
  INVX1    g12790(.A(new_n12927_), .Y(new_n13047_));
  NOR2X1   g12791(.A(new_n12938_), .B(new_n12924_), .Y(new_n13048_));
  AOI21X1  g12792(.A0(new_n12937_), .A1(new_n13047_), .B0(new_n13048_), .Y(new_n13049_));
  INVX1    g12793(.A(new_n12928_), .Y(new_n13050_));
  OR2X1    g12794(.A(new_n12931_), .B(new_n13050_), .Y(new_n13051_));
  OR2X1    g12795(.A(new_n12936_), .B(new_n12932_), .Y(new_n13052_));
  AND2X1   g12796(.A(new_n13052_), .B(new_n13051_), .Y(new_n13053_));
  AOI22X1  g12797(.A0(new_n7818_), .A1(\b[34] ), .B0(new_n7817_), .B1(\b[35] ), .Y(new_n13054_));
  NOR2X1   g12798(.A(new_n13054_), .B(new_n13050_), .Y(new_n13055_));
  XOR2X1   g12799(.A(new_n13054_), .B(new_n13050_), .Y(new_n13056_));
  NAND2X1  g12800(.A(new_n13054_), .B(new_n13050_), .Y(new_n13057_));
  OAI21X1  g12801(.A0(new_n13055_), .A1(new_n13053_), .B0(new_n13057_), .Y(new_n13058_));
  OAI22X1  g12802(.A0(new_n13058_), .A1(new_n13055_), .B0(new_n13056_), .B1(new_n13053_), .Y(new_n13059_));
  AOI22X1  g12803(.A0(new_n7192_), .A1(\b[38] ), .B0(new_n7189_), .B1(\b[37] ), .Y(new_n13060_));
  OAI21X1  g12804(.A0(new_n7627_), .A1(new_n3276_), .B0(new_n13060_), .Y(new_n13061_));
  AOI21X1  g12805(.A0(new_n7187_), .A1(new_n3275_), .B0(new_n13061_), .Y(new_n13062_));
  XOR2X1   g12806(.A(new_n13062_), .B(\a[62] ), .Y(new_n13063_));
  XOR2X1   g12807(.A(new_n13063_), .B(new_n13059_), .Y(new_n13064_));
  AOI22X1  g12808(.A0(new_n6603_), .A1(\b[41] ), .B0(new_n6600_), .B1(\b[40] ), .Y(new_n13065_));
  OAI21X1  g12809(.A0(new_n6804_), .A1(new_n3723_), .B0(new_n13065_), .Y(new_n13066_));
  AOI21X1  g12810(.A0(new_n6598_), .A1(new_n3722_), .B0(new_n13066_), .Y(new_n13067_));
  XOR2X1   g12811(.A(new_n13067_), .B(\a[59] ), .Y(new_n13068_));
  INVX1    g12812(.A(new_n13068_), .Y(new_n13069_));
  XOR2X1   g12813(.A(new_n13069_), .B(new_n13064_), .Y(new_n13070_));
  XOR2X1   g12814(.A(new_n13070_), .B(new_n13049_), .Y(new_n13071_));
  XOR2X1   g12815(.A(new_n13071_), .B(new_n13046_), .Y(new_n13072_));
  XOR2X1   g12816(.A(new_n13072_), .B(new_n13042_), .Y(new_n13073_));
  AOI22X1  g12817(.A0(new_n5430_), .A1(\b[47] ), .B0(new_n5427_), .B1(\b[46] ), .Y(new_n13074_));
  OAI21X1  g12818(.A0(new_n5891_), .A1(new_n4674_), .B0(new_n13074_), .Y(new_n13075_));
  AOI21X1  g12819(.A0(new_n5425_), .A1(new_n4673_), .B0(new_n13075_), .Y(new_n13076_));
  XOR2X1   g12820(.A(new_n13076_), .B(\a[53] ), .Y(new_n13077_));
  XOR2X1   g12821(.A(new_n13077_), .B(new_n13073_), .Y(new_n13078_));
  INVX1    g12822(.A(new_n13078_), .Y(new_n13079_));
  NOR2X1   g12823(.A(new_n12948_), .B(new_n12945_), .Y(new_n13080_));
  INVX1    g12824(.A(new_n12953_), .Y(new_n13081_));
  AOI21X1  g12825(.A0(new_n13081_), .A1(new_n12949_), .B0(new_n13080_), .Y(new_n13082_));
  XOR2X1   g12826(.A(new_n13082_), .B(new_n13079_), .Y(new_n13083_));
  AOI22X1  g12827(.A0(new_n4880_), .A1(\b[50] ), .B0(new_n4877_), .B1(\b[49] ), .Y(new_n13084_));
  OAI21X1  g12828(.A0(new_n5291_), .A1(new_n5036_), .B0(new_n13084_), .Y(new_n13085_));
  AOI21X1  g12829(.A0(new_n5204_), .A1(new_n4875_), .B0(new_n13085_), .Y(new_n13086_));
  XOR2X1   g12830(.A(new_n13086_), .B(\a[50] ), .Y(new_n13087_));
  XOR2X1   g12831(.A(new_n13087_), .B(new_n13083_), .Y(new_n13088_));
  XOR2X1   g12832(.A(new_n13088_), .B(new_n13038_), .Y(new_n13089_));
  XOR2X1   g12833(.A(new_n13089_), .B(new_n13033_), .Y(new_n13090_));
  XOR2X1   g12834(.A(new_n13090_), .B(new_n13029_), .Y(new_n13091_));
  XOR2X1   g12835(.A(new_n13091_), .B(new_n13026_), .Y(new_n13092_));
  XOR2X1   g12836(.A(new_n13092_), .B(new_n13022_), .Y(new_n13093_));
  AOI22X1  g12837(.A0(new_n3652_), .A1(\b[59] ), .B0(new_n3651_), .B1(\b[58] ), .Y(new_n13094_));
  OAI21X1  g12838(.A0(new_n3778_), .A1(new_n6933_), .B0(new_n13094_), .Y(new_n13095_));
  AOI21X1  g12839(.A0(new_n6932_), .A1(new_n3480_), .B0(new_n13095_), .Y(new_n13096_));
  XOR2X1   g12840(.A(new_n13096_), .B(\a[41] ), .Y(new_n13097_));
  XOR2X1   g12841(.A(new_n13097_), .B(new_n13093_), .Y(new_n13098_));
  AND2X1   g12842(.A(new_n12979_), .B(new_n12917_), .Y(new_n13099_));
  INVX1    g12843(.A(new_n12984_), .Y(new_n13100_));
  AOI21X1  g12844(.A0(new_n13100_), .A1(new_n12980_), .B0(new_n13099_), .Y(new_n13101_));
  XOR2X1   g12845(.A(new_n13101_), .B(new_n13098_), .Y(new_n13102_));
  AOI22X1  g12846(.A0(new_n3204_), .A1(\b[62] ), .B0(new_n3203_), .B1(\b[61] ), .Y(new_n13103_));
  OAI21X1  g12847(.A0(new_n3321_), .A1(new_n7559_), .B0(new_n13103_), .Y(new_n13104_));
  AOI21X1  g12848(.A0(new_n7558_), .A1(new_n3080_), .B0(new_n13104_), .Y(new_n13105_));
  XOR2X1   g12849(.A(new_n13105_), .B(\a[38] ), .Y(new_n13106_));
  XOR2X1   g12850(.A(new_n13106_), .B(new_n13102_), .Y(new_n13107_));
  XOR2X1   g12851(.A(new_n13107_), .B(new_n13020_), .Y(new_n13108_));
  XOR2X1   g12852(.A(new_n13108_), .B(new_n13013_), .Y(new_n13109_));
  XOR2X1   g12853(.A(new_n13109_), .B(new_n13011_), .Y(\f[98] ));
  NOR2X1   g12854(.A(new_n13108_), .B(new_n13013_), .Y(new_n13111_));
  INVX1    g12855(.A(new_n13109_), .Y(new_n13112_));
  AOI21X1  g12856(.A0(new_n13010_), .A1(new_n13008_), .B0(new_n13112_), .Y(new_n13113_));
  OR2X1    g12857(.A(new_n13113_), .B(new_n13111_), .Y(new_n13114_));
  AND2X1   g12858(.A(new_n13088_), .B(new_n13037_), .Y(new_n13115_));
  INVX1    g12859(.A(new_n13115_), .Y(new_n13116_));
  OAI21X1  g12860(.A0(new_n13089_), .A1(new_n13033_), .B0(new_n13116_), .Y(new_n13117_));
  AOI22X1  g12861(.A0(new_n4572_), .A1(\b[54] ), .B0(new_n4571_), .B1(\b[53] ), .Y(new_n13118_));
  OAI21X1  g12862(.A0(new_n4740_), .A1(new_n5808_), .B0(new_n13118_), .Y(new_n13119_));
  AOI21X1  g12863(.A0(new_n5807_), .A1(new_n4375_), .B0(new_n13119_), .Y(new_n13120_));
  XOR2X1   g12864(.A(new_n13120_), .B(new_n4568_), .Y(new_n13121_));
  OR2X1    g12865(.A(new_n13082_), .B(new_n13078_), .Y(new_n13122_));
  OAI21X1  g12866(.A0(new_n13087_), .A1(new_n13083_), .B0(new_n13122_), .Y(new_n13123_));
  AOI22X1  g12867(.A0(new_n7818_), .A1(\b[35] ), .B0(new_n7817_), .B1(\b[36] ), .Y(new_n13124_));
  XOR2X1   g12868(.A(new_n13054_), .B(new_n2650_), .Y(new_n13125_));
  XOR2X1   g12869(.A(new_n13125_), .B(new_n13124_), .Y(new_n13126_));
  XOR2X1   g12870(.A(new_n13126_), .B(new_n13058_), .Y(new_n13127_));
  AOI22X1  g12871(.A0(new_n7192_), .A1(\b[39] ), .B0(new_n7189_), .B1(\b[38] ), .Y(new_n13128_));
  OAI21X1  g12872(.A0(new_n7627_), .A1(new_n3413_), .B0(new_n13128_), .Y(new_n13129_));
  AOI21X1  g12873(.A0(new_n7187_), .A1(new_n3412_), .B0(new_n13129_), .Y(new_n13130_));
  XOR2X1   g12874(.A(new_n13130_), .B(\a[62] ), .Y(new_n13131_));
  XOR2X1   g12875(.A(new_n13131_), .B(new_n13127_), .Y(new_n13132_));
  AOI22X1  g12876(.A0(new_n6603_), .A1(\b[42] ), .B0(new_n6600_), .B1(\b[41] ), .Y(new_n13133_));
  OAI21X1  g12877(.A0(new_n6804_), .A1(new_n3720_), .B0(new_n13133_), .Y(new_n13134_));
  AOI21X1  g12878(.A0(new_n6598_), .A1(new_n3860_), .B0(new_n13134_), .Y(new_n13135_));
  XOR2X1   g12879(.A(new_n13135_), .B(\a[59] ), .Y(new_n13136_));
  XOR2X1   g12880(.A(new_n13136_), .B(new_n13132_), .Y(new_n13137_));
  INVX1    g12881(.A(new_n13063_), .Y(new_n13138_));
  AND2X1   g12882(.A(new_n13138_), .B(new_n13059_), .Y(new_n13139_));
  NOR2X1   g12883(.A(new_n13068_), .B(new_n13064_), .Y(new_n13140_));
  NOR2X1   g12884(.A(new_n13140_), .B(new_n13139_), .Y(new_n13141_));
  XOR2X1   g12885(.A(new_n13141_), .B(new_n13137_), .Y(new_n13142_));
  AOI22X1  g12886(.A0(new_n6438_), .A1(\b[45] ), .B0(new_n6437_), .B1(\b[44] ), .Y(new_n13143_));
  OAI21X1  g12887(.A0(new_n6436_), .A1(new_n4339_), .B0(new_n13143_), .Y(new_n13144_));
  AOI21X1  g12888(.A0(new_n6023_), .A1(new_n4338_), .B0(new_n13144_), .Y(new_n13145_));
  XOR2X1   g12889(.A(new_n13145_), .B(\a[56] ), .Y(new_n13146_));
  XOR2X1   g12890(.A(new_n13146_), .B(new_n13142_), .Y(new_n13147_));
  INVX1    g12891(.A(new_n13147_), .Y(new_n13148_));
  NOR2X1   g12892(.A(new_n13070_), .B(new_n13049_), .Y(new_n13149_));
  AOI21X1  g12893(.A0(new_n13071_), .A1(new_n13046_), .B0(new_n13149_), .Y(new_n13150_));
  XOR2X1   g12894(.A(new_n13150_), .B(new_n13148_), .Y(new_n13151_));
  AOI22X1  g12895(.A0(new_n5430_), .A1(\b[48] ), .B0(new_n5427_), .B1(\b[47] ), .Y(new_n13152_));
  OAI21X1  g12896(.A0(new_n5891_), .A1(new_n4693_), .B0(new_n13152_), .Y(new_n13153_));
  AOI21X1  g12897(.A0(new_n5425_), .A1(new_n4692_), .B0(new_n13153_), .Y(new_n13154_));
  XOR2X1   g12898(.A(new_n13154_), .B(\a[53] ), .Y(new_n13155_));
  XOR2X1   g12899(.A(new_n13155_), .B(new_n13151_), .Y(new_n13156_));
  INVX1    g12900(.A(new_n13156_), .Y(new_n13157_));
  AND2X1   g12901(.A(new_n13072_), .B(new_n13042_), .Y(new_n13158_));
  INVX1    g12902(.A(new_n13077_), .Y(new_n13159_));
  AOI21X1  g12903(.A0(new_n13159_), .A1(new_n13073_), .B0(new_n13158_), .Y(new_n13160_));
  XOR2X1   g12904(.A(new_n13160_), .B(new_n13157_), .Y(new_n13161_));
  AOI22X1  g12905(.A0(new_n4880_), .A1(\b[51] ), .B0(new_n4877_), .B1(\b[50] ), .Y(new_n13162_));
  OAI21X1  g12906(.A0(new_n5291_), .A1(new_n5237_), .B0(new_n13162_), .Y(new_n13163_));
  AOI21X1  g12907(.A0(new_n5236_), .A1(new_n4875_), .B0(new_n13163_), .Y(new_n13164_));
  XOR2X1   g12908(.A(new_n13164_), .B(\a[50] ), .Y(new_n13165_));
  XOR2X1   g12909(.A(new_n13165_), .B(new_n13161_), .Y(new_n13166_));
  XOR2X1   g12910(.A(new_n13166_), .B(new_n13123_), .Y(new_n13167_));
  XOR2X1   g12911(.A(new_n13167_), .B(new_n13121_), .Y(new_n13168_));
  XOR2X1   g12912(.A(new_n13168_), .B(new_n13117_), .Y(new_n13169_));
  AOI22X1  g12913(.A0(new_n4095_), .A1(\b[57] ), .B0(new_n4094_), .B1(\b[56] ), .Y(new_n13170_));
  OAI21X1  g12914(.A0(new_n4233_), .A1(new_n6523_), .B0(new_n13170_), .Y(new_n13171_));
  AOI21X1  g12915(.A0(new_n6522_), .A1(new_n3901_), .B0(new_n13171_), .Y(new_n13172_));
  XOR2X1   g12916(.A(new_n13172_), .B(\a[44] ), .Y(new_n13173_));
  XOR2X1   g12917(.A(new_n13173_), .B(new_n13169_), .Y(new_n13174_));
  AND2X1   g12918(.A(new_n13090_), .B(new_n13029_), .Y(new_n13175_));
  AOI21X1  g12919(.A0(new_n13091_), .A1(new_n13026_), .B0(new_n13175_), .Y(new_n13176_));
  XOR2X1   g12920(.A(new_n13176_), .B(new_n13174_), .Y(new_n13177_));
  AOI22X1  g12921(.A0(new_n3652_), .A1(\b[60] ), .B0(new_n3651_), .B1(\b[59] ), .Y(new_n13178_));
  OAI21X1  g12922(.A0(new_n3778_), .A1(new_n6930_), .B0(new_n13178_), .Y(new_n13179_));
  AOI21X1  g12923(.A0(new_n6951_), .A1(new_n3480_), .B0(new_n13179_), .Y(new_n13180_));
  XOR2X1   g12924(.A(new_n13180_), .B(\a[41] ), .Y(new_n13181_));
  XOR2X1   g12925(.A(new_n13181_), .B(new_n13177_), .Y(new_n13182_));
  AND2X1   g12926(.A(new_n13092_), .B(new_n13022_), .Y(new_n13183_));
  INVX1    g12927(.A(new_n13097_), .Y(new_n13184_));
  AOI21X1  g12928(.A0(new_n13184_), .A1(new_n13093_), .B0(new_n13183_), .Y(new_n13185_));
  XOR2X1   g12929(.A(new_n13185_), .B(new_n13182_), .Y(new_n13186_));
  AOI22X1  g12930(.A0(new_n3204_), .A1(\b[63] ), .B0(new_n3203_), .B1(\b[62] ), .Y(new_n13187_));
  OAI21X1  g12931(.A0(new_n3321_), .A1(new_n7748_), .B0(new_n13187_), .Y(new_n13188_));
  AOI21X1  g12932(.A0(new_n7747_), .A1(new_n3080_), .B0(new_n13188_), .Y(new_n13189_));
  XOR2X1   g12933(.A(new_n13189_), .B(\a[38] ), .Y(new_n13190_));
  XOR2X1   g12934(.A(new_n13190_), .B(new_n13186_), .Y(new_n13191_));
  INVX1    g12935(.A(new_n13191_), .Y(new_n13192_));
  NOR2X1   g12936(.A(new_n13101_), .B(new_n13098_), .Y(new_n13193_));
  INVX1    g12937(.A(new_n13106_), .Y(new_n13194_));
  AOI21X1  g12938(.A0(new_n13194_), .A1(new_n13102_), .B0(new_n13193_), .Y(new_n13195_));
  XOR2X1   g12939(.A(new_n13195_), .B(new_n13192_), .Y(new_n13196_));
  AOI21X1  g12940(.A0(new_n13015_), .A1(new_n13014_), .B0(new_n13019_), .Y(new_n13197_));
  INVX1    g12941(.A(new_n13107_), .Y(new_n13198_));
  AOI21X1  g12942(.A0(new_n13198_), .A1(new_n13020_), .B0(new_n13197_), .Y(new_n13199_));
  XOR2X1   g12943(.A(new_n13199_), .B(new_n13196_), .Y(new_n13200_));
  XOR2X1   g12944(.A(new_n13200_), .B(new_n13114_), .Y(\f[99] ));
  XOR2X1   g12945(.A(new_n13180_), .B(new_n3478_), .Y(new_n13202_));
  NOR2X1   g12946(.A(new_n13185_), .B(new_n13182_), .Y(new_n13203_));
  AOI21X1  g12947(.A0(new_n13202_), .A1(new_n13177_), .B0(new_n13203_), .Y(new_n13204_));
  OAI22X1  g12948(.A0(new_n3321_), .A1(new_n7745_), .B0(new_n3082_), .B1(new_n7772_), .Y(new_n13205_));
  AOI21X1  g12949(.A0(new_n7775_), .A1(new_n3080_), .B0(new_n13205_), .Y(new_n13206_));
  XOR2X1   g12950(.A(new_n13206_), .B(\a[38] ), .Y(new_n13207_));
  XOR2X1   g12951(.A(new_n13207_), .B(new_n13204_), .Y(new_n13208_));
  AOI22X1  g12952(.A0(new_n7192_), .A1(\b[40] ), .B0(new_n7189_), .B1(\b[39] ), .Y(new_n13209_));
  OAI21X1  g12953(.A0(new_n7627_), .A1(new_n3575_), .B0(new_n13209_), .Y(new_n13210_));
  AOI21X1  g12954(.A0(new_n7187_), .A1(new_n3574_), .B0(new_n13210_), .Y(new_n13211_));
  XOR2X1   g12955(.A(new_n13211_), .B(new_n7185_), .Y(new_n13212_));
  AOI22X1  g12956(.A0(new_n7818_), .A1(\b[36] ), .B0(new_n7817_), .B1(\b[37] ), .Y(new_n13213_));
  OR2X1    g12957(.A(new_n13125_), .B(new_n13124_), .Y(new_n13214_));
  OR2X1    g12958(.A(new_n13054_), .B(\a[35] ), .Y(new_n13215_));
  AND2X1   g12959(.A(new_n13215_), .B(new_n13214_), .Y(new_n13216_));
  XOR2X1   g12960(.A(new_n13216_), .B(new_n13213_), .Y(new_n13217_));
  XOR2X1   g12961(.A(new_n13217_), .B(new_n13212_), .Y(new_n13218_));
  AND2X1   g12962(.A(new_n13126_), .B(new_n13058_), .Y(new_n13219_));
  INVX1    g12963(.A(new_n13131_), .Y(new_n13220_));
  AOI21X1  g12964(.A0(new_n13220_), .A1(new_n13127_), .B0(new_n13219_), .Y(new_n13221_));
  XOR2X1   g12965(.A(new_n13221_), .B(new_n13218_), .Y(new_n13222_));
  AOI22X1  g12966(.A0(new_n6603_), .A1(\b[43] ), .B0(new_n6600_), .B1(\b[42] ), .Y(new_n13223_));
  OAI21X1  g12967(.A0(new_n6804_), .A1(new_n4015_), .B0(new_n13223_), .Y(new_n13224_));
  AOI21X1  g12968(.A0(new_n6598_), .A1(new_n4014_), .B0(new_n13224_), .Y(new_n13225_));
  XOR2X1   g12969(.A(new_n13225_), .B(\a[59] ), .Y(new_n13226_));
  XOR2X1   g12970(.A(new_n13226_), .B(new_n13222_), .Y(new_n13227_));
  OR2X1    g12971(.A(new_n13136_), .B(new_n13132_), .Y(new_n13228_));
  OAI21X1  g12972(.A0(new_n13140_), .A1(new_n13139_), .B0(new_n13137_), .Y(new_n13229_));
  AND2X1   g12973(.A(new_n13229_), .B(new_n13228_), .Y(new_n13230_));
  XOR2X1   g12974(.A(new_n13230_), .B(new_n13227_), .Y(new_n13231_));
  AOI22X1  g12975(.A0(new_n6438_), .A1(\b[46] ), .B0(new_n6437_), .B1(\b[45] ), .Y(new_n13232_));
  OAI21X1  g12976(.A0(new_n6436_), .A1(new_n4336_), .B0(new_n13232_), .Y(new_n13233_));
  AOI21X1  g12977(.A0(new_n6023_), .A1(new_n4509_), .B0(new_n13233_), .Y(new_n13234_));
  XOR2X1   g12978(.A(new_n13234_), .B(\a[56] ), .Y(new_n13235_));
  XOR2X1   g12979(.A(new_n13235_), .B(new_n13231_), .Y(new_n13236_));
  INVX1    g12980(.A(new_n13236_), .Y(new_n13237_));
  OR2X1    g12981(.A(new_n13146_), .B(new_n13142_), .Y(new_n13238_));
  OAI21X1  g12982(.A0(new_n13150_), .A1(new_n13148_), .B0(new_n13238_), .Y(new_n13239_));
  XOR2X1   g12983(.A(new_n13239_), .B(new_n13237_), .Y(new_n13240_));
  AOI22X1  g12984(.A0(new_n5430_), .A1(\b[49] ), .B0(new_n5427_), .B1(\b[48] ), .Y(new_n13241_));
  OAI21X1  g12985(.A0(new_n5891_), .A1(new_n5039_), .B0(new_n13241_), .Y(new_n13242_));
  AOI21X1  g12986(.A0(new_n5425_), .A1(new_n5038_), .B0(new_n13242_), .Y(new_n13243_));
  XOR2X1   g12987(.A(new_n13243_), .B(\a[53] ), .Y(new_n13244_));
  XOR2X1   g12988(.A(new_n13244_), .B(new_n13240_), .Y(new_n13245_));
  INVX1    g12989(.A(new_n13155_), .Y(new_n13246_));
  NOR2X1   g12990(.A(new_n13160_), .B(new_n13156_), .Y(new_n13247_));
  AOI21X1  g12991(.A0(new_n13246_), .A1(new_n13151_), .B0(new_n13247_), .Y(new_n13248_));
  XOR2X1   g12992(.A(new_n13248_), .B(new_n13245_), .Y(new_n13249_));
  AOI22X1  g12993(.A0(new_n4880_), .A1(\b[52] ), .B0(new_n4877_), .B1(\b[51] ), .Y(new_n13250_));
  OAI21X1  g12994(.A0(new_n5291_), .A1(new_n5234_), .B0(new_n13250_), .Y(new_n13251_));
  AOI21X1  g12995(.A0(new_n5590_), .A1(new_n4875_), .B0(new_n13251_), .Y(new_n13252_));
  XOR2X1   g12996(.A(new_n13252_), .B(\a[50] ), .Y(new_n13253_));
  XOR2X1   g12997(.A(new_n13253_), .B(new_n13249_), .Y(new_n13254_));
  NOR2X1   g12998(.A(new_n13165_), .B(new_n13161_), .Y(new_n13255_));
  AOI21X1  g12999(.A0(new_n13166_), .A1(new_n13123_), .B0(new_n13255_), .Y(new_n13256_));
  XOR2X1   g13000(.A(new_n13256_), .B(new_n13254_), .Y(new_n13257_));
  AOI22X1  g13001(.A0(new_n4572_), .A1(\b[55] ), .B0(new_n4571_), .B1(\b[54] ), .Y(new_n13258_));
  OAI21X1  g13002(.A0(new_n4740_), .A1(new_n6151_), .B0(new_n13258_), .Y(new_n13259_));
  AOI21X1  g13003(.A0(new_n6150_), .A1(new_n4375_), .B0(new_n13259_), .Y(new_n13260_));
  XOR2X1   g13004(.A(new_n13260_), .B(\a[47] ), .Y(new_n13261_));
  XOR2X1   g13005(.A(new_n13261_), .B(new_n13257_), .Y(new_n13262_));
  AND2X1   g13006(.A(new_n13167_), .B(new_n13121_), .Y(new_n13263_));
  AOI21X1  g13007(.A0(new_n13168_), .A1(new_n13117_), .B0(new_n13263_), .Y(new_n13264_));
  XOR2X1   g13008(.A(new_n13264_), .B(new_n13262_), .Y(new_n13265_));
  AOI22X1  g13009(.A0(new_n4095_), .A1(\b[58] ), .B0(new_n4094_), .B1(\b[57] ), .Y(new_n13266_));
  OAI21X1  g13010(.A0(new_n4233_), .A1(new_n6520_), .B0(new_n13266_), .Y(new_n13267_));
  AOI21X1  g13011(.A0(new_n6732_), .A1(new_n3901_), .B0(new_n13267_), .Y(new_n13268_));
  XOR2X1   g13012(.A(new_n13268_), .B(\a[44] ), .Y(new_n13269_));
  XOR2X1   g13013(.A(new_n13269_), .B(new_n13265_), .Y(new_n13270_));
  INVX1    g13014(.A(new_n13270_), .Y(new_n13271_));
  INVX1    g13015(.A(new_n13173_), .Y(new_n13272_));
  NOR2X1   g13016(.A(new_n13176_), .B(new_n13174_), .Y(new_n13273_));
  AOI21X1  g13017(.A0(new_n13272_), .A1(new_n13169_), .B0(new_n13273_), .Y(new_n13274_));
  XOR2X1   g13018(.A(new_n13274_), .B(new_n13271_), .Y(new_n13275_));
  AOI22X1  g13019(.A0(new_n3652_), .A1(\b[61] ), .B0(new_n3651_), .B1(\b[60] ), .Y(new_n13276_));
  OAI21X1  g13020(.A0(new_n3778_), .A1(new_n7339_), .B0(new_n13276_), .Y(new_n13277_));
  AOI21X1  g13021(.A0(new_n7338_), .A1(new_n3480_), .B0(new_n13277_), .Y(new_n13278_));
  XOR2X1   g13022(.A(new_n13278_), .B(\a[41] ), .Y(new_n13279_));
  XOR2X1   g13023(.A(new_n13279_), .B(new_n13275_), .Y(new_n13280_));
  XOR2X1   g13024(.A(new_n13280_), .B(new_n13208_), .Y(new_n13281_));
  INVX1    g13025(.A(new_n13190_), .Y(new_n13282_));
  NOR2X1   g13026(.A(new_n13195_), .B(new_n13191_), .Y(new_n13283_));
  AOI21X1  g13027(.A0(new_n13282_), .A1(new_n13186_), .B0(new_n13283_), .Y(new_n13284_));
  XOR2X1   g13028(.A(new_n13284_), .B(new_n13281_), .Y(new_n13285_));
  OR2X1    g13029(.A(new_n13199_), .B(new_n13196_), .Y(new_n13286_));
  OAI21X1  g13030(.A0(new_n13113_), .A1(new_n13111_), .B0(new_n13200_), .Y(new_n13287_));
  AND2X1   g13031(.A(new_n13287_), .B(new_n13286_), .Y(new_n13288_));
  XOR2X1   g13032(.A(new_n13288_), .B(new_n13285_), .Y(\f[100] ));
  INVX1    g13033(.A(new_n13281_), .Y(new_n13290_));
  NOR2X1   g13034(.A(new_n13284_), .B(new_n13290_), .Y(new_n13291_));
  AOI21X1  g13035(.A0(new_n13287_), .A1(new_n13286_), .B0(new_n13285_), .Y(new_n13292_));
  OR2X1    g13036(.A(new_n13292_), .B(new_n13291_), .Y(new_n13293_));
  NOR2X1   g13037(.A(new_n13207_), .B(new_n13204_), .Y(new_n13294_));
  AOI21X1  g13038(.A0(new_n13280_), .A1(new_n13208_), .B0(new_n13294_), .Y(new_n13295_));
  OR2X1    g13039(.A(new_n13274_), .B(new_n13270_), .Y(new_n13296_));
  OR2X1    g13040(.A(new_n13279_), .B(new_n13275_), .Y(new_n13297_));
  AND2X1   g13041(.A(new_n13297_), .B(new_n13296_), .Y(new_n13298_));
  NOR3X1   g13042(.A(new_n3320_), .B(new_n3079_), .C(new_n7772_), .Y(new_n13299_));
  AOI21X1  g13043(.A0(new_n7774_), .A1(new_n3080_), .B0(new_n13299_), .Y(new_n13300_));
  XOR2X1   g13044(.A(new_n13300_), .B(\a[38] ), .Y(new_n13301_));
  XOR2X1   g13045(.A(new_n13301_), .B(new_n13298_), .Y(new_n13302_));
  NOR2X1   g13046(.A(new_n13256_), .B(new_n13254_), .Y(new_n13303_));
  INVX1    g13047(.A(new_n13303_), .Y(new_n13304_));
  INVX1    g13048(.A(new_n13257_), .Y(new_n13305_));
  OAI21X1  g13049(.A0(new_n13261_), .A1(new_n13305_), .B0(new_n13304_), .Y(new_n13306_));
  AOI22X1  g13050(.A0(new_n4572_), .A1(\b[56] ), .B0(new_n4571_), .B1(\b[55] ), .Y(new_n13307_));
  OAI21X1  g13051(.A0(new_n4740_), .A1(new_n6148_), .B0(new_n13307_), .Y(new_n13308_));
  AOI21X1  g13052(.A0(new_n6342_), .A1(new_n4375_), .B0(new_n13308_), .Y(new_n13309_));
  XOR2X1   g13053(.A(new_n13309_), .B(new_n4568_), .Y(new_n13310_));
  AND2X1   g13054(.A(new_n13248_), .B(new_n13245_), .Y(new_n13311_));
  OR2X1    g13055(.A(new_n13248_), .B(new_n13245_), .Y(new_n13312_));
  OAI21X1  g13056(.A0(new_n13253_), .A1(new_n13311_), .B0(new_n13312_), .Y(new_n13313_));
  AOI22X1  g13057(.A0(new_n4880_), .A1(\b[53] ), .B0(new_n4877_), .B1(\b[52] ), .Y(new_n13314_));
  OAI21X1  g13058(.A0(new_n5291_), .A1(new_n5787_), .B0(new_n13314_), .Y(new_n13315_));
  AOI21X1  g13059(.A0(new_n5786_), .A1(new_n4875_), .B0(new_n13315_), .Y(new_n13316_));
  XOR2X1   g13060(.A(new_n13316_), .B(\a[50] ), .Y(new_n13317_));
  AND2X1   g13061(.A(new_n13239_), .B(new_n13237_), .Y(new_n13318_));
  INVX1    g13062(.A(new_n13318_), .Y(new_n13319_));
  INVX1    g13063(.A(new_n13240_), .Y(new_n13320_));
  OAI21X1  g13064(.A0(new_n13244_), .A1(new_n13320_), .B0(new_n13319_), .Y(new_n13321_));
  INVX1    g13065(.A(new_n13321_), .Y(new_n13322_));
  INVX1    g13066(.A(new_n13213_), .Y(new_n13323_));
  AOI21X1  g13067(.A0(new_n13215_), .A1(new_n13214_), .B0(new_n13323_), .Y(new_n13324_));
  INVX1    g13068(.A(new_n13217_), .Y(new_n13325_));
  AOI21X1  g13069(.A0(new_n13325_), .A1(new_n13212_), .B0(new_n13324_), .Y(new_n13326_));
  AOI22X1  g13070(.A0(new_n7818_), .A1(\b[37] ), .B0(new_n7817_), .B1(\b[38] ), .Y(new_n13327_));
  XOR2X1   g13071(.A(new_n13327_), .B(new_n13213_), .Y(new_n13328_));
  XOR2X1   g13072(.A(new_n13328_), .B(new_n13326_), .Y(new_n13329_));
  AOI22X1  g13073(.A0(new_n7192_), .A1(\b[41] ), .B0(new_n7189_), .B1(\b[40] ), .Y(new_n13330_));
  OAI21X1  g13074(.A0(new_n7627_), .A1(new_n3723_), .B0(new_n13330_), .Y(new_n13331_));
  AOI21X1  g13075(.A0(new_n7187_), .A1(new_n3722_), .B0(new_n13331_), .Y(new_n13332_));
  XOR2X1   g13076(.A(new_n13332_), .B(\a[62] ), .Y(new_n13333_));
  XOR2X1   g13077(.A(new_n13333_), .B(new_n13329_), .Y(new_n13334_));
  INVX1    g13078(.A(new_n13334_), .Y(new_n13335_));
  AOI22X1  g13079(.A0(new_n6603_), .A1(\b[44] ), .B0(new_n6600_), .B1(\b[43] ), .Y(new_n13336_));
  OAI21X1  g13080(.A0(new_n6804_), .A1(new_n4012_), .B0(new_n13336_), .Y(new_n13337_));
  AOI21X1  g13081(.A0(new_n6598_), .A1(new_n4178_), .B0(new_n13337_), .Y(new_n13338_));
  XOR2X1   g13082(.A(new_n13338_), .B(\a[59] ), .Y(new_n13339_));
  XOR2X1   g13083(.A(new_n13339_), .B(new_n13335_), .Y(new_n13340_));
  NOR2X1   g13084(.A(new_n13221_), .B(new_n13218_), .Y(new_n13341_));
  INVX1    g13085(.A(new_n13226_), .Y(new_n13342_));
  AOI21X1  g13086(.A0(new_n13342_), .A1(new_n13222_), .B0(new_n13341_), .Y(new_n13343_));
  XOR2X1   g13087(.A(new_n13343_), .B(new_n13340_), .Y(new_n13344_));
  AOI22X1  g13088(.A0(new_n6438_), .A1(\b[47] ), .B0(new_n6437_), .B1(\b[46] ), .Y(new_n13345_));
  OAI21X1  g13089(.A0(new_n6436_), .A1(new_n4674_), .B0(new_n13345_), .Y(new_n13346_));
  AOI21X1  g13090(.A0(new_n6023_), .A1(new_n4673_), .B0(new_n13346_), .Y(new_n13347_));
  XOR2X1   g13091(.A(new_n13347_), .B(\a[56] ), .Y(new_n13348_));
  XOR2X1   g13092(.A(new_n13348_), .B(new_n13344_), .Y(new_n13349_));
  INVX1    g13093(.A(new_n13349_), .Y(new_n13350_));
  AOI21X1  g13094(.A0(new_n13229_), .A1(new_n13228_), .B0(new_n13227_), .Y(new_n13351_));
  INVX1    g13095(.A(new_n13235_), .Y(new_n13352_));
  AOI21X1  g13096(.A0(new_n13352_), .A1(new_n13231_), .B0(new_n13351_), .Y(new_n13353_));
  XOR2X1   g13097(.A(new_n13353_), .B(new_n13350_), .Y(new_n13354_));
  AOI22X1  g13098(.A0(new_n5430_), .A1(\b[50] ), .B0(new_n5427_), .B1(\b[49] ), .Y(new_n13355_));
  OAI21X1  g13099(.A0(new_n5891_), .A1(new_n5036_), .B0(new_n13355_), .Y(new_n13356_));
  AOI21X1  g13100(.A0(new_n5425_), .A1(new_n5204_), .B0(new_n13356_), .Y(new_n13357_));
  XOR2X1   g13101(.A(new_n13357_), .B(\a[53] ), .Y(new_n13358_));
  XOR2X1   g13102(.A(new_n13358_), .B(new_n13354_), .Y(new_n13359_));
  XOR2X1   g13103(.A(new_n13359_), .B(new_n13322_), .Y(new_n13360_));
  XOR2X1   g13104(.A(new_n13360_), .B(new_n13317_), .Y(new_n13361_));
  XOR2X1   g13105(.A(new_n13361_), .B(new_n13313_), .Y(new_n13362_));
  XOR2X1   g13106(.A(new_n13362_), .B(new_n13310_), .Y(new_n13363_));
  XOR2X1   g13107(.A(new_n13363_), .B(new_n13306_), .Y(new_n13364_));
  AOI22X1  g13108(.A0(new_n4095_), .A1(\b[59] ), .B0(new_n4094_), .B1(\b[58] ), .Y(new_n13365_));
  OAI21X1  g13109(.A0(new_n4233_), .A1(new_n6933_), .B0(new_n13365_), .Y(new_n13366_));
  AOI21X1  g13110(.A0(new_n6932_), .A1(new_n3901_), .B0(new_n13366_), .Y(new_n13367_));
  XOR2X1   g13111(.A(new_n13367_), .B(\a[44] ), .Y(new_n13368_));
  XOR2X1   g13112(.A(new_n13368_), .B(new_n13364_), .Y(new_n13369_));
  NOR2X1   g13113(.A(new_n13264_), .B(new_n13262_), .Y(new_n13370_));
  INVX1    g13114(.A(new_n13269_), .Y(new_n13371_));
  AOI21X1  g13115(.A0(new_n13371_), .A1(new_n13265_), .B0(new_n13370_), .Y(new_n13372_));
  XOR2X1   g13116(.A(new_n13372_), .B(new_n13369_), .Y(new_n13373_));
  AOI22X1  g13117(.A0(new_n3652_), .A1(\b[62] ), .B0(new_n3651_), .B1(\b[61] ), .Y(new_n13374_));
  OAI21X1  g13118(.A0(new_n3778_), .A1(new_n7559_), .B0(new_n13374_), .Y(new_n13375_));
  AOI21X1  g13119(.A0(new_n7558_), .A1(new_n3480_), .B0(new_n13375_), .Y(new_n13376_));
  XOR2X1   g13120(.A(new_n13376_), .B(\a[41] ), .Y(new_n13377_));
  XOR2X1   g13121(.A(new_n13377_), .B(new_n13373_), .Y(new_n13378_));
  XOR2X1   g13122(.A(new_n13378_), .B(new_n13302_), .Y(new_n13379_));
  XOR2X1   g13123(.A(new_n13379_), .B(new_n13295_), .Y(new_n13380_));
  XOR2X1   g13124(.A(new_n13380_), .B(new_n13293_), .Y(\f[101] ));
  NOR2X1   g13125(.A(new_n13379_), .B(new_n13295_), .Y(new_n13382_));
  INVX1    g13126(.A(new_n13382_), .Y(new_n13383_));
  OAI21X1  g13127(.A0(new_n13292_), .A1(new_n13291_), .B0(new_n13380_), .Y(new_n13384_));
  NAND2X1  g13128(.A(new_n13384_), .B(new_n13383_), .Y(new_n13385_));
  AND2X1   g13129(.A(new_n13359_), .B(new_n13321_), .Y(new_n13386_));
  INVX1    g13130(.A(new_n13386_), .Y(new_n13387_));
  OAI21X1  g13131(.A0(new_n13360_), .A1(new_n13317_), .B0(new_n13387_), .Y(new_n13388_));
  AOI22X1  g13132(.A0(new_n4880_), .A1(\b[54] ), .B0(new_n4877_), .B1(\b[53] ), .Y(new_n13389_));
  OAI21X1  g13133(.A0(new_n5291_), .A1(new_n5808_), .B0(new_n13389_), .Y(new_n13390_));
  AOI21X1  g13134(.A0(new_n5807_), .A1(new_n4875_), .B0(new_n13390_), .Y(new_n13391_));
  XOR2X1   g13135(.A(new_n13391_), .B(new_n4873_), .Y(new_n13392_));
  OR2X1    g13136(.A(new_n13353_), .B(new_n13349_), .Y(new_n13393_));
  OAI21X1  g13137(.A0(new_n13358_), .A1(new_n13354_), .B0(new_n13393_), .Y(new_n13394_));
  OR2X1    g13138(.A(new_n13327_), .B(new_n13323_), .Y(new_n13395_));
  OAI21X1  g13139(.A0(new_n13328_), .A1(new_n13326_), .B0(new_n13395_), .Y(new_n13396_));
  AOI22X1  g13140(.A0(new_n7818_), .A1(\b[38] ), .B0(new_n7817_), .B1(\b[39] ), .Y(new_n13397_));
  XOR2X1   g13141(.A(new_n13213_), .B(new_n3078_), .Y(new_n13398_));
  XOR2X1   g13142(.A(new_n13398_), .B(new_n13397_), .Y(new_n13399_));
  XOR2X1   g13143(.A(new_n13399_), .B(new_n13396_), .Y(new_n13400_));
  AOI22X1  g13144(.A0(new_n7192_), .A1(\b[42] ), .B0(new_n7189_), .B1(\b[41] ), .Y(new_n13401_));
  OAI21X1  g13145(.A0(new_n7627_), .A1(new_n3720_), .B0(new_n13401_), .Y(new_n13402_));
  AOI21X1  g13146(.A0(new_n7187_), .A1(new_n3860_), .B0(new_n13402_), .Y(new_n13403_));
  XOR2X1   g13147(.A(new_n13403_), .B(\a[62] ), .Y(new_n13404_));
  XOR2X1   g13148(.A(new_n13404_), .B(new_n13400_), .Y(new_n13405_));
  AOI22X1  g13149(.A0(new_n6603_), .A1(\b[45] ), .B0(new_n6600_), .B1(\b[44] ), .Y(new_n13406_));
  OAI21X1  g13150(.A0(new_n6804_), .A1(new_n4339_), .B0(new_n13406_), .Y(new_n13407_));
  AOI21X1  g13151(.A0(new_n6598_), .A1(new_n4338_), .B0(new_n13407_), .Y(new_n13408_));
  XOR2X1   g13152(.A(new_n13408_), .B(\a[59] ), .Y(new_n13409_));
  XOR2X1   g13153(.A(new_n13409_), .B(new_n13405_), .Y(new_n13410_));
  XOR2X1   g13154(.A(new_n13332_), .B(new_n7185_), .Y(new_n13411_));
  AND2X1   g13155(.A(new_n13411_), .B(new_n13329_), .Y(new_n13412_));
  NOR2X1   g13156(.A(new_n13339_), .B(new_n13334_), .Y(new_n13413_));
  NOR2X1   g13157(.A(new_n13413_), .B(new_n13412_), .Y(new_n13414_));
  XOR2X1   g13158(.A(new_n13414_), .B(new_n13410_), .Y(new_n13415_));
  AOI22X1  g13159(.A0(new_n6438_), .A1(\b[48] ), .B0(new_n6437_), .B1(\b[47] ), .Y(new_n13416_));
  OAI21X1  g13160(.A0(new_n6436_), .A1(new_n4693_), .B0(new_n13416_), .Y(new_n13417_));
  AOI21X1  g13161(.A0(new_n6023_), .A1(new_n4692_), .B0(new_n13417_), .Y(new_n13418_));
  XOR2X1   g13162(.A(new_n13418_), .B(\a[56] ), .Y(new_n13419_));
  XOR2X1   g13163(.A(new_n13419_), .B(new_n13415_), .Y(new_n13420_));
  NOR2X1   g13164(.A(new_n13343_), .B(new_n13340_), .Y(new_n13421_));
  INVX1    g13165(.A(new_n13348_), .Y(new_n13422_));
  AOI21X1  g13166(.A0(new_n13422_), .A1(new_n13344_), .B0(new_n13421_), .Y(new_n13423_));
  XOR2X1   g13167(.A(new_n13423_), .B(new_n13420_), .Y(new_n13424_));
  AOI22X1  g13168(.A0(new_n5430_), .A1(\b[51] ), .B0(new_n5427_), .B1(\b[50] ), .Y(new_n13425_));
  OAI21X1  g13169(.A0(new_n5891_), .A1(new_n5237_), .B0(new_n13425_), .Y(new_n13426_));
  AOI21X1  g13170(.A0(new_n5425_), .A1(new_n5236_), .B0(new_n13426_), .Y(new_n13427_));
  XOR2X1   g13171(.A(new_n13427_), .B(\a[53] ), .Y(new_n13428_));
  XOR2X1   g13172(.A(new_n13428_), .B(new_n13424_), .Y(new_n13429_));
  XOR2X1   g13173(.A(new_n13429_), .B(new_n13394_), .Y(new_n13430_));
  XOR2X1   g13174(.A(new_n13430_), .B(new_n13392_), .Y(new_n13431_));
  XOR2X1   g13175(.A(new_n13431_), .B(new_n13388_), .Y(new_n13432_));
  AOI22X1  g13176(.A0(new_n4572_), .A1(\b[57] ), .B0(new_n4571_), .B1(\b[56] ), .Y(new_n13433_));
  OAI21X1  g13177(.A0(new_n4740_), .A1(new_n6523_), .B0(new_n13433_), .Y(new_n13434_));
  AOI21X1  g13178(.A0(new_n6522_), .A1(new_n4375_), .B0(new_n13434_), .Y(new_n13435_));
  XOR2X1   g13179(.A(new_n13435_), .B(\a[47] ), .Y(new_n13436_));
  XOR2X1   g13180(.A(new_n13436_), .B(new_n13432_), .Y(new_n13437_));
  AND2X1   g13181(.A(new_n13361_), .B(new_n13313_), .Y(new_n13438_));
  AOI21X1  g13182(.A0(new_n13362_), .A1(new_n13310_), .B0(new_n13438_), .Y(new_n13439_));
  XOR2X1   g13183(.A(new_n13439_), .B(new_n13437_), .Y(new_n13440_));
  AOI22X1  g13184(.A0(new_n4095_), .A1(\b[60] ), .B0(new_n4094_), .B1(\b[59] ), .Y(new_n13441_));
  OAI21X1  g13185(.A0(new_n4233_), .A1(new_n6930_), .B0(new_n13441_), .Y(new_n13442_));
  AOI21X1  g13186(.A0(new_n6951_), .A1(new_n3901_), .B0(new_n13442_), .Y(new_n13443_));
  XOR2X1   g13187(.A(new_n13443_), .B(\a[44] ), .Y(new_n13444_));
  XOR2X1   g13188(.A(new_n13444_), .B(new_n13440_), .Y(new_n13445_));
  AND2X1   g13189(.A(new_n13363_), .B(new_n13306_), .Y(new_n13446_));
  INVX1    g13190(.A(new_n13368_), .Y(new_n13447_));
  AOI21X1  g13191(.A0(new_n13447_), .A1(new_n13364_), .B0(new_n13446_), .Y(new_n13448_));
  XOR2X1   g13192(.A(new_n13448_), .B(new_n13445_), .Y(new_n13449_));
  AOI22X1  g13193(.A0(new_n3652_), .A1(\b[63] ), .B0(new_n3651_), .B1(\b[62] ), .Y(new_n13450_));
  OAI21X1  g13194(.A0(new_n3778_), .A1(new_n7748_), .B0(new_n13450_), .Y(new_n13451_));
  AOI21X1  g13195(.A0(new_n7747_), .A1(new_n3480_), .B0(new_n13451_), .Y(new_n13452_));
  XOR2X1   g13196(.A(new_n13452_), .B(\a[41] ), .Y(new_n13453_));
  XOR2X1   g13197(.A(new_n13453_), .B(new_n13449_), .Y(new_n13454_));
  NOR2X1   g13198(.A(new_n13372_), .B(new_n13369_), .Y(new_n13455_));
  INVX1    g13199(.A(new_n13377_), .Y(new_n13456_));
  AOI21X1  g13200(.A0(new_n13456_), .A1(new_n13373_), .B0(new_n13455_), .Y(new_n13457_));
  XOR2X1   g13201(.A(new_n13457_), .B(new_n13454_), .Y(new_n13458_));
  INVX1    g13202(.A(new_n13458_), .Y(new_n13459_));
  NOR2X1   g13203(.A(new_n13301_), .B(new_n13298_), .Y(new_n13460_));
  INVX1    g13204(.A(new_n13378_), .Y(new_n13461_));
  AOI21X1  g13205(.A0(new_n13461_), .A1(new_n13302_), .B0(new_n13460_), .Y(new_n13462_));
  XOR2X1   g13206(.A(new_n13462_), .B(new_n13459_), .Y(new_n13463_));
  XOR2X1   g13207(.A(new_n13463_), .B(new_n13385_), .Y(\f[102] ));
  XOR2X1   g13208(.A(new_n13443_), .B(new_n3899_), .Y(new_n13465_));
  NOR2X1   g13209(.A(new_n13448_), .B(new_n13445_), .Y(new_n13466_));
  AOI21X1  g13210(.A0(new_n13465_), .A1(new_n13440_), .B0(new_n13466_), .Y(new_n13467_));
  OAI22X1  g13211(.A0(new_n3778_), .A1(new_n7745_), .B0(new_n3482_), .B1(new_n7772_), .Y(new_n13468_));
  AOI21X1  g13212(.A0(new_n7775_), .A1(new_n3480_), .B0(new_n13468_), .Y(new_n13469_));
  XOR2X1   g13213(.A(new_n13469_), .B(\a[41] ), .Y(new_n13470_));
  XOR2X1   g13214(.A(new_n13470_), .B(new_n13467_), .Y(new_n13471_));
  AND2X1   g13215(.A(new_n13399_), .B(new_n13396_), .Y(new_n13472_));
  INVX1    g13216(.A(new_n13404_), .Y(new_n13473_));
  AOI21X1  g13217(.A0(new_n13473_), .A1(new_n13400_), .B0(new_n13472_), .Y(new_n13474_));
  AOI22X1  g13218(.A0(new_n7818_), .A1(\b[39] ), .B0(new_n7817_), .B1(\b[40] ), .Y(new_n13475_));
  INVX1    g13219(.A(new_n13475_), .Y(new_n13476_));
  NOR2X1   g13220(.A(new_n13398_), .B(new_n13397_), .Y(new_n13477_));
  AOI21X1  g13221(.A0(new_n13323_), .A1(new_n3078_), .B0(new_n13477_), .Y(new_n13478_));
  XOR2X1   g13222(.A(new_n13478_), .B(new_n13476_), .Y(new_n13479_));
  INVX1    g13223(.A(new_n13479_), .Y(new_n13480_));
  AOI22X1  g13224(.A0(new_n7192_), .A1(\b[43] ), .B0(new_n7189_), .B1(\b[42] ), .Y(new_n13481_));
  OAI21X1  g13225(.A0(new_n7627_), .A1(new_n4015_), .B0(new_n13481_), .Y(new_n13482_));
  AOI21X1  g13226(.A0(new_n7187_), .A1(new_n4014_), .B0(new_n13482_), .Y(new_n13483_));
  XOR2X1   g13227(.A(new_n13483_), .B(\a[62] ), .Y(new_n13484_));
  XOR2X1   g13228(.A(new_n13484_), .B(new_n13480_), .Y(new_n13485_));
  INVX1    g13229(.A(new_n13485_), .Y(new_n13486_));
  XOR2X1   g13230(.A(new_n13486_), .B(new_n13474_), .Y(new_n13487_));
  AOI22X1  g13231(.A0(new_n6603_), .A1(\b[46] ), .B0(new_n6600_), .B1(\b[45] ), .Y(new_n13488_));
  OAI21X1  g13232(.A0(new_n6804_), .A1(new_n4336_), .B0(new_n13488_), .Y(new_n13489_));
  AOI21X1  g13233(.A0(new_n6598_), .A1(new_n4509_), .B0(new_n13489_), .Y(new_n13490_));
  XOR2X1   g13234(.A(new_n13490_), .B(\a[59] ), .Y(new_n13491_));
  XOR2X1   g13235(.A(new_n13491_), .B(new_n13487_), .Y(new_n13492_));
  OR2X1    g13236(.A(new_n13409_), .B(new_n13405_), .Y(new_n13493_));
  OAI21X1  g13237(.A0(new_n13413_), .A1(new_n13412_), .B0(new_n13410_), .Y(new_n13494_));
  AND2X1   g13238(.A(new_n13494_), .B(new_n13493_), .Y(new_n13495_));
  XOR2X1   g13239(.A(new_n13495_), .B(new_n13492_), .Y(new_n13496_));
  AOI22X1  g13240(.A0(new_n6438_), .A1(\b[49] ), .B0(new_n6437_), .B1(\b[48] ), .Y(new_n13497_));
  OAI21X1  g13241(.A0(new_n6436_), .A1(new_n5039_), .B0(new_n13497_), .Y(new_n13498_));
  AOI21X1  g13242(.A0(new_n6023_), .A1(new_n5038_), .B0(new_n13498_), .Y(new_n13499_));
  XOR2X1   g13243(.A(new_n13499_), .B(\a[56] ), .Y(new_n13500_));
  XOR2X1   g13244(.A(new_n13500_), .B(new_n13496_), .Y(new_n13501_));
  INVX1    g13245(.A(new_n13501_), .Y(new_n13502_));
  OR2X1    g13246(.A(new_n13419_), .B(new_n13415_), .Y(new_n13503_));
  INVX1    g13247(.A(new_n13420_), .Y(new_n13504_));
  OAI21X1  g13248(.A0(new_n13423_), .A1(new_n13504_), .B0(new_n13503_), .Y(new_n13505_));
  XOR2X1   g13249(.A(new_n13505_), .B(new_n13502_), .Y(new_n13506_));
  AOI22X1  g13250(.A0(new_n5430_), .A1(\b[52] ), .B0(new_n5427_), .B1(\b[51] ), .Y(new_n13507_));
  OAI21X1  g13251(.A0(new_n5891_), .A1(new_n5234_), .B0(new_n13507_), .Y(new_n13508_));
  AOI21X1  g13252(.A0(new_n5590_), .A1(new_n5425_), .B0(new_n13508_), .Y(new_n13509_));
  XOR2X1   g13253(.A(new_n13509_), .B(\a[53] ), .Y(new_n13510_));
  XOR2X1   g13254(.A(new_n13510_), .B(new_n13506_), .Y(new_n13511_));
  NOR2X1   g13255(.A(new_n13428_), .B(new_n13424_), .Y(new_n13512_));
  AOI21X1  g13256(.A0(new_n13429_), .A1(new_n13394_), .B0(new_n13512_), .Y(new_n13513_));
  XOR2X1   g13257(.A(new_n13513_), .B(new_n13511_), .Y(new_n13514_));
  AOI22X1  g13258(.A0(new_n4880_), .A1(\b[55] ), .B0(new_n4877_), .B1(\b[54] ), .Y(new_n13515_));
  OAI21X1  g13259(.A0(new_n5291_), .A1(new_n6151_), .B0(new_n13515_), .Y(new_n13516_));
  AOI21X1  g13260(.A0(new_n6150_), .A1(new_n4875_), .B0(new_n13516_), .Y(new_n13517_));
  XOR2X1   g13261(.A(new_n13517_), .B(\a[50] ), .Y(new_n13518_));
  XOR2X1   g13262(.A(new_n13518_), .B(new_n13514_), .Y(new_n13519_));
  AND2X1   g13263(.A(new_n13430_), .B(new_n13392_), .Y(new_n13520_));
  AOI21X1  g13264(.A0(new_n13431_), .A1(new_n13388_), .B0(new_n13520_), .Y(new_n13521_));
  XOR2X1   g13265(.A(new_n13521_), .B(new_n13519_), .Y(new_n13522_));
  AOI22X1  g13266(.A0(new_n4572_), .A1(\b[58] ), .B0(new_n4571_), .B1(\b[57] ), .Y(new_n13523_));
  OAI21X1  g13267(.A0(new_n4740_), .A1(new_n6520_), .B0(new_n13523_), .Y(new_n13524_));
  AOI21X1  g13268(.A0(new_n6732_), .A1(new_n4375_), .B0(new_n13524_), .Y(new_n13525_));
  XOR2X1   g13269(.A(new_n13525_), .B(\a[47] ), .Y(new_n13526_));
  XOR2X1   g13270(.A(new_n13526_), .B(new_n13522_), .Y(new_n13527_));
  INVX1    g13271(.A(new_n13527_), .Y(new_n13528_));
  INVX1    g13272(.A(new_n13436_), .Y(new_n13529_));
  NOR2X1   g13273(.A(new_n13439_), .B(new_n13437_), .Y(new_n13530_));
  AOI21X1  g13274(.A0(new_n13529_), .A1(new_n13432_), .B0(new_n13530_), .Y(new_n13531_));
  XOR2X1   g13275(.A(new_n13531_), .B(new_n13528_), .Y(new_n13532_));
  AOI22X1  g13276(.A0(new_n4095_), .A1(\b[61] ), .B0(new_n4094_), .B1(\b[60] ), .Y(new_n13533_));
  OAI21X1  g13277(.A0(new_n4233_), .A1(new_n7339_), .B0(new_n13533_), .Y(new_n13534_));
  AOI21X1  g13278(.A0(new_n7338_), .A1(new_n3901_), .B0(new_n13534_), .Y(new_n13535_));
  XOR2X1   g13279(.A(new_n13535_), .B(\a[44] ), .Y(new_n13536_));
  XOR2X1   g13280(.A(new_n13536_), .B(new_n13532_), .Y(new_n13537_));
  XOR2X1   g13281(.A(new_n13537_), .B(new_n13471_), .Y(new_n13538_));
  INVX1    g13282(.A(new_n13538_), .Y(new_n13539_));
  INVX1    g13283(.A(new_n13453_), .Y(new_n13540_));
  NOR2X1   g13284(.A(new_n13457_), .B(new_n13454_), .Y(new_n13541_));
  AOI21X1  g13285(.A0(new_n13540_), .A1(new_n13449_), .B0(new_n13541_), .Y(new_n13542_));
  XOR2X1   g13286(.A(new_n13542_), .B(new_n13539_), .Y(new_n13543_));
  NOR2X1   g13287(.A(new_n13462_), .B(new_n13459_), .Y(new_n13544_));
  INVX1    g13288(.A(new_n13463_), .Y(new_n13545_));
  AOI21X1  g13289(.A0(new_n13384_), .A1(new_n13383_), .B0(new_n13545_), .Y(new_n13546_));
  OR2X1    g13290(.A(new_n13546_), .B(new_n13544_), .Y(new_n13547_));
  XOR2X1   g13291(.A(new_n13547_), .B(new_n13543_), .Y(\f[103] ));
  NOR2X1   g13292(.A(new_n13542_), .B(new_n13539_), .Y(new_n13549_));
  INVX1    g13293(.A(new_n13549_), .Y(new_n13550_));
  OAI21X1  g13294(.A0(new_n13546_), .A1(new_n13544_), .B0(new_n13543_), .Y(new_n13551_));
  NAND2X1  g13295(.A(new_n13551_), .B(new_n13550_), .Y(new_n13552_));
  NOR2X1   g13296(.A(new_n13470_), .B(new_n13467_), .Y(new_n13553_));
  AOI21X1  g13297(.A0(new_n13537_), .A1(new_n13471_), .B0(new_n13553_), .Y(new_n13554_));
  OR2X1    g13298(.A(new_n13531_), .B(new_n13527_), .Y(new_n13555_));
  OR2X1    g13299(.A(new_n13536_), .B(new_n13532_), .Y(new_n13556_));
  AND2X1   g13300(.A(new_n13556_), .B(new_n13555_), .Y(new_n13557_));
  NOR3X1   g13301(.A(new_n3777_), .B(new_n3479_), .C(new_n7772_), .Y(new_n13558_));
  AOI21X1  g13302(.A0(new_n7774_), .A1(new_n3480_), .B0(new_n13558_), .Y(new_n13559_));
  XOR2X1   g13303(.A(new_n13559_), .B(\a[41] ), .Y(new_n13560_));
  XOR2X1   g13304(.A(new_n13560_), .B(new_n13557_), .Y(new_n13561_));
  NOR2X1   g13305(.A(new_n13513_), .B(new_n13511_), .Y(new_n13562_));
  INVX1    g13306(.A(new_n13562_), .Y(new_n13563_));
  INVX1    g13307(.A(new_n13514_), .Y(new_n13564_));
  OAI21X1  g13308(.A0(new_n13518_), .A1(new_n13564_), .B0(new_n13563_), .Y(new_n13565_));
  AOI22X1  g13309(.A0(new_n4880_), .A1(\b[56] ), .B0(new_n4877_), .B1(\b[55] ), .Y(new_n13566_));
  OAI21X1  g13310(.A0(new_n5291_), .A1(new_n6148_), .B0(new_n13566_), .Y(new_n13567_));
  AOI21X1  g13311(.A0(new_n6342_), .A1(new_n4875_), .B0(new_n13567_), .Y(new_n13568_));
  XOR2X1   g13312(.A(new_n13568_), .B(\a[50] ), .Y(new_n13569_));
  AND2X1   g13313(.A(new_n13505_), .B(new_n13502_), .Y(new_n13570_));
  INVX1    g13314(.A(new_n13570_), .Y(new_n13571_));
  INVX1    g13315(.A(new_n13506_), .Y(new_n13572_));
  OAI21X1  g13316(.A0(new_n13510_), .A1(new_n13572_), .B0(new_n13571_), .Y(new_n13573_));
  INVX1    g13317(.A(new_n13573_), .Y(new_n13574_));
  AOI22X1  g13318(.A0(new_n5430_), .A1(\b[53] ), .B0(new_n5427_), .B1(\b[52] ), .Y(new_n13575_));
  OAI21X1  g13319(.A0(new_n5891_), .A1(new_n5787_), .B0(new_n13575_), .Y(new_n13576_));
  AOI21X1  g13320(.A0(new_n5786_), .A1(new_n5425_), .B0(new_n13576_), .Y(new_n13577_));
  XOR2X1   g13321(.A(new_n13577_), .B(\a[53] ), .Y(new_n13578_));
  AOI21X1  g13322(.A0(new_n13494_), .A1(new_n13493_), .B0(new_n13492_), .Y(new_n13579_));
  INVX1    g13323(.A(new_n13579_), .Y(new_n13580_));
  INVX1    g13324(.A(new_n13496_), .Y(new_n13581_));
  OAI21X1  g13325(.A0(new_n13500_), .A1(new_n13581_), .B0(new_n13580_), .Y(new_n13582_));
  INVX1    g13326(.A(new_n13582_), .Y(new_n13583_));
  NOR2X1   g13327(.A(new_n13486_), .B(new_n13474_), .Y(new_n13584_));
  INVX1    g13328(.A(new_n13584_), .Y(new_n13585_));
  INVX1    g13329(.A(new_n13487_), .Y(new_n13586_));
  OAI21X1  g13330(.A0(new_n13491_), .A1(new_n13586_), .B0(new_n13585_), .Y(new_n13587_));
  INVX1    g13331(.A(new_n13587_), .Y(new_n13588_));
  NOR2X1   g13332(.A(new_n13478_), .B(new_n13476_), .Y(new_n13589_));
  XOR2X1   g13333(.A(new_n13483_), .B(new_n7185_), .Y(new_n13590_));
  AOI21X1  g13334(.A0(new_n13590_), .A1(new_n13479_), .B0(new_n13589_), .Y(new_n13591_));
  AOI22X1  g13335(.A0(new_n7818_), .A1(\b[40] ), .B0(new_n7817_), .B1(\b[41] ), .Y(new_n13592_));
  XOR2X1   g13336(.A(new_n13592_), .B(new_n13475_), .Y(new_n13593_));
  XOR2X1   g13337(.A(new_n13593_), .B(new_n13591_), .Y(new_n13594_));
  AOI22X1  g13338(.A0(new_n7192_), .A1(\b[44] ), .B0(new_n7189_), .B1(\b[43] ), .Y(new_n13595_));
  OAI21X1  g13339(.A0(new_n7627_), .A1(new_n4012_), .B0(new_n13595_), .Y(new_n13596_));
  AOI21X1  g13340(.A0(new_n7187_), .A1(new_n4178_), .B0(new_n13596_), .Y(new_n13597_));
  XOR2X1   g13341(.A(new_n13597_), .B(\a[62] ), .Y(new_n13598_));
  XOR2X1   g13342(.A(new_n13598_), .B(new_n13594_), .Y(new_n13599_));
  AOI22X1  g13343(.A0(new_n6603_), .A1(\b[47] ), .B0(new_n6600_), .B1(\b[46] ), .Y(new_n13600_));
  OAI21X1  g13344(.A0(new_n6804_), .A1(new_n4674_), .B0(new_n13600_), .Y(new_n13601_));
  AOI21X1  g13345(.A0(new_n6598_), .A1(new_n4673_), .B0(new_n13601_), .Y(new_n13602_));
  XOR2X1   g13346(.A(new_n13602_), .B(\a[59] ), .Y(new_n13603_));
  XOR2X1   g13347(.A(new_n13603_), .B(new_n13599_), .Y(new_n13604_));
  XOR2X1   g13348(.A(new_n13604_), .B(new_n13588_), .Y(new_n13605_));
  AOI22X1  g13349(.A0(new_n6438_), .A1(\b[50] ), .B0(new_n6437_), .B1(\b[49] ), .Y(new_n13606_));
  OAI21X1  g13350(.A0(new_n6436_), .A1(new_n5036_), .B0(new_n13606_), .Y(new_n13607_));
  AOI21X1  g13351(.A0(new_n6023_), .A1(new_n5204_), .B0(new_n13607_), .Y(new_n13608_));
  XOR2X1   g13352(.A(new_n13608_), .B(\a[56] ), .Y(new_n13609_));
  XOR2X1   g13353(.A(new_n13609_), .B(new_n13605_), .Y(new_n13610_));
  XOR2X1   g13354(.A(new_n13610_), .B(new_n13583_), .Y(new_n13611_));
  XOR2X1   g13355(.A(new_n13611_), .B(new_n13578_), .Y(new_n13612_));
  XOR2X1   g13356(.A(new_n13612_), .B(new_n13574_), .Y(new_n13613_));
  XOR2X1   g13357(.A(new_n13613_), .B(new_n13569_), .Y(new_n13614_));
  XOR2X1   g13358(.A(new_n13614_), .B(new_n13565_), .Y(new_n13615_));
  AOI22X1  g13359(.A0(new_n4572_), .A1(\b[59] ), .B0(new_n4571_), .B1(\b[58] ), .Y(new_n13616_));
  OAI21X1  g13360(.A0(new_n4740_), .A1(new_n6933_), .B0(new_n13616_), .Y(new_n13617_));
  AOI21X1  g13361(.A0(new_n6932_), .A1(new_n4375_), .B0(new_n13617_), .Y(new_n13618_));
  XOR2X1   g13362(.A(new_n13618_), .B(\a[47] ), .Y(new_n13619_));
  XOR2X1   g13363(.A(new_n13619_), .B(new_n13615_), .Y(new_n13620_));
  NOR2X1   g13364(.A(new_n13521_), .B(new_n13519_), .Y(new_n13621_));
  INVX1    g13365(.A(new_n13526_), .Y(new_n13622_));
  AOI21X1  g13366(.A0(new_n13622_), .A1(new_n13522_), .B0(new_n13621_), .Y(new_n13623_));
  XOR2X1   g13367(.A(new_n13623_), .B(new_n13620_), .Y(new_n13624_));
  AOI22X1  g13368(.A0(new_n4095_), .A1(\b[62] ), .B0(new_n4094_), .B1(\b[61] ), .Y(new_n13625_));
  OAI21X1  g13369(.A0(new_n4233_), .A1(new_n7559_), .B0(new_n13625_), .Y(new_n13626_));
  AOI21X1  g13370(.A0(new_n7558_), .A1(new_n3901_), .B0(new_n13626_), .Y(new_n13627_));
  XOR2X1   g13371(.A(new_n13627_), .B(\a[44] ), .Y(new_n13628_));
  XOR2X1   g13372(.A(new_n13628_), .B(new_n13624_), .Y(new_n13629_));
  XOR2X1   g13373(.A(new_n13629_), .B(new_n13561_), .Y(new_n13630_));
  XOR2X1   g13374(.A(new_n13630_), .B(new_n13554_), .Y(new_n13631_));
  XOR2X1   g13375(.A(new_n13631_), .B(new_n13552_), .Y(\f[104] ));
  NOR2X1   g13376(.A(new_n13630_), .B(new_n13554_), .Y(new_n13633_));
  INVX1    g13377(.A(new_n13631_), .Y(new_n13634_));
  AOI21X1  g13378(.A0(new_n13551_), .A1(new_n13550_), .B0(new_n13634_), .Y(new_n13635_));
  OR2X1    g13379(.A(new_n13635_), .B(new_n13633_), .Y(new_n13636_));
  AND2X1   g13380(.A(new_n13612_), .B(new_n13573_), .Y(new_n13637_));
  INVX1    g13381(.A(new_n13637_), .Y(new_n13638_));
  OAI21X1  g13382(.A0(new_n13613_), .A1(new_n13569_), .B0(new_n13638_), .Y(new_n13639_));
  AOI22X1  g13383(.A0(new_n4880_), .A1(\b[57] ), .B0(new_n4877_), .B1(\b[56] ), .Y(new_n13640_));
  OAI21X1  g13384(.A0(new_n5291_), .A1(new_n6523_), .B0(new_n13640_), .Y(new_n13641_));
  AOI21X1  g13385(.A0(new_n6522_), .A1(new_n4875_), .B0(new_n13641_), .Y(new_n13642_));
  XOR2X1   g13386(.A(new_n13642_), .B(new_n4873_), .Y(new_n13643_));
  NAND2X1  g13387(.A(new_n13610_), .B(new_n13582_), .Y(new_n13644_));
  OAI21X1  g13388(.A0(new_n13611_), .A1(new_n13578_), .B0(new_n13644_), .Y(new_n13645_));
  NAND2X1  g13389(.A(new_n13604_), .B(new_n13587_), .Y(new_n13646_));
  OAI21X1  g13390(.A0(new_n13609_), .A1(new_n13605_), .B0(new_n13646_), .Y(new_n13647_));
  AOI22X1  g13391(.A0(new_n6438_), .A1(\b[51] ), .B0(new_n6437_), .B1(\b[50] ), .Y(new_n13648_));
  OAI21X1  g13392(.A0(new_n6436_), .A1(new_n5237_), .B0(new_n13648_), .Y(new_n13649_));
  AOI21X1  g13393(.A0(new_n6023_), .A1(new_n5236_), .B0(new_n13649_), .Y(new_n13650_));
  XOR2X1   g13394(.A(new_n13650_), .B(\a[56] ), .Y(new_n13651_));
  XOR2X1   g13395(.A(new_n13475_), .B(new_n3478_), .Y(new_n13652_));
  AOI22X1  g13396(.A0(new_n7818_), .A1(\b[41] ), .B0(new_n7817_), .B1(\b[42] ), .Y(new_n13653_));
  XOR2X1   g13397(.A(new_n13653_), .B(new_n13652_), .Y(new_n13654_));
  AOI22X1  g13398(.A0(new_n7192_), .A1(\b[45] ), .B0(new_n7189_), .B1(\b[44] ), .Y(new_n13655_));
  OAI21X1  g13399(.A0(new_n7627_), .A1(new_n4339_), .B0(new_n13655_), .Y(new_n13656_));
  AOI21X1  g13400(.A0(new_n7187_), .A1(new_n4338_), .B0(new_n13656_), .Y(new_n13657_));
  XOR2X1   g13401(.A(new_n13657_), .B(\a[62] ), .Y(new_n13658_));
  XOR2X1   g13402(.A(new_n13658_), .B(new_n13654_), .Y(new_n13659_));
  INVX1    g13403(.A(new_n13659_), .Y(new_n13660_));
  OR2X1    g13404(.A(new_n13592_), .B(new_n13476_), .Y(new_n13661_));
  OAI21X1  g13405(.A0(new_n13593_), .A1(new_n13591_), .B0(new_n13661_), .Y(new_n13662_));
  XOR2X1   g13406(.A(new_n13662_), .B(new_n13660_), .Y(new_n13663_));
  AOI22X1  g13407(.A0(new_n6603_), .A1(\b[48] ), .B0(new_n6600_), .B1(\b[47] ), .Y(new_n13664_));
  OAI21X1  g13408(.A0(new_n6804_), .A1(new_n4693_), .B0(new_n13664_), .Y(new_n13665_));
  AOI21X1  g13409(.A0(new_n6598_), .A1(new_n4692_), .B0(new_n13665_), .Y(new_n13666_));
  XOR2X1   g13410(.A(new_n13666_), .B(\a[59] ), .Y(new_n13667_));
  XOR2X1   g13411(.A(new_n13667_), .B(new_n13663_), .Y(new_n13668_));
  INVX1    g13412(.A(new_n13598_), .Y(new_n13669_));
  NOR2X1   g13413(.A(new_n13603_), .B(new_n13599_), .Y(new_n13670_));
  AOI21X1  g13414(.A0(new_n13669_), .A1(new_n13594_), .B0(new_n13670_), .Y(new_n13671_));
  XOR2X1   g13415(.A(new_n13671_), .B(new_n13668_), .Y(new_n13672_));
  XOR2X1   g13416(.A(new_n13672_), .B(new_n13651_), .Y(new_n13673_));
  XOR2X1   g13417(.A(new_n13673_), .B(new_n13647_), .Y(new_n13674_));
  AOI22X1  g13418(.A0(new_n5430_), .A1(\b[54] ), .B0(new_n5427_), .B1(\b[53] ), .Y(new_n13675_));
  OAI21X1  g13419(.A0(new_n5891_), .A1(new_n5808_), .B0(new_n13675_), .Y(new_n13676_));
  AOI21X1  g13420(.A0(new_n5807_), .A1(new_n5425_), .B0(new_n13676_), .Y(new_n13677_));
  XOR2X1   g13421(.A(new_n13677_), .B(\a[53] ), .Y(new_n13678_));
  XOR2X1   g13422(.A(new_n13678_), .B(new_n13674_), .Y(new_n13679_));
  XOR2X1   g13423(.A(new_n13679_), .B(new_n13645_), .Y(new_n13680_));
  XOR2X1   g13424(.A(new_n13680_), .B(new_n13643_), .Y(new_n13681_));
  XOR2X1   g13425(.A(new_n13681_), .B(new_n13639_), .Y(new_n13682_));
  AOI22X1  g13426(.A0(new_n4572_), .A1(\b[60] ), .B0(new_n4571_), .B1(\b[59] ), .Y(new_n13683_));
  OAI21X1  g13427(.A0(new_n4740_), .A1(new_n6930_), .B0(new_n13683_), .Y(new_n13684_));
  AOI21X1  g13428(.A0(new_n6951_), .A1(new_n4375_), .B0(new_n13684_), .Y(new_n13685_));
  XOR2X1   g13429(.A(new_n13685_), .B(\a[47] ), .Y(new_n13686_));
  XOR2X1   g13430(.A(new_n13686_), .B(new_n13682_), .Y(new_n13687_));
  AND2X1   g13431(.A(new_n13614_), .B(new_n13565_), .Y(new_n13688_));
  INVX1    g13432(.A(new_n13619_), .Y(new_n13689_));
  AOI21X1  g13433(.A0(new_n13689_), .A1(new_n13615_), .B0(new_n13688_), .Y(new_n13690_));
  XOR2X1   g13434(.A(new_n13690_), .B(new_n13687_), .Y(new_n13691_));
  AOI22X1  g13435(.A0(new_n4095_), .A1(\b[63] ), .B0(new_n4094_), .B1(\b[62] ), .Y(new_n13692_));
  OAI21X1  g13436(.A0(new_n4233_), .A1(new_n7748_), .B0(new_n13692_), .Y(new_n13693_));
  AOI21X1  g13437(.A0(new_n7747_), .A1(new_n3901_), .B0(new_n13693_), .Y(new_n13694_));
  XOR2X1   g13438(.A(new_n13694_), .B(\a[44] ), .Y(new_n13695_));
  XOR2X1   g13439(.A(new_n13695_), .B(new_n13691_), .Y(new_n13696_));
  NOR2X1   g13440(.A(new_n13623_), .B(new_n13620_), .Y(new_n13697_));
  INVX1    g13441(.A(new_n13628_), .Y(new_n13698_));
  AOI21X1  g13442(.A0(new_n13698_), .A1(new_n13624_), .B0(new_n13697_), .Y(new_n13699_));
  XOR2X1   g13443(.A(new_n13699_), .B(new_n13696_), .Y(new_n13700_));
  INVX1    g13444(.A(new_n13700_), .Y(new_n13701_));
  NOR2X1   g13445(.A(new_n13560_), .B(new_n13557_), .Y(new_n13702_));
  INVX1    g13446(.A(new_n13629_), .Y(new_n13703_));
  AOI21X1  g13447(.A0(new_n13703_), .A1(new_n13561_), .B0(new_n13702_), .Y(new_n13704_));
  XOR2X1   g13448(.A(new_n13704_), .B(new_n13701_), .Y(new_n13705_));
  XOR2X1   g13449(.A(new_n13705_), .B(new_n13636_), .Y(\f[105] ));
  XOR2X1   g13450(.A(new_n13685_), .B(new_n4568_), .Y(new_n13707_));
  NOR2X1   g13451(.A(new_n13690_), .B(new_n13687_), .Y(new_n13708_));
  AOI21X1  g13452(.A0(new_n13707_), .A1(new_n13682_), .B0(new_n13708_), .Y(new_n13709_));
  OAI22X1  g13453(.A0(new_n4233_), .A1(new_n7745_), .B0(new_n3903_), .B1(new_n7772_), .Y(new_n13710_));
  AOI21X1  g13454(.A0(new_n7775_), .A1(new_n3901_), .B0(new_n13710_), .Y(new_n13711_));
  XOR2X1   g13455(.A(new_n13711_), .B(\a[44] ), .Y(new_n13712_));
  XOR2X1   g13456(.A(new_n13712_), .B(new_n13709_), .Y(new_n13713_));
  AOI22X1  g13457(.A0(new_n4572_), .A1(\b[61] ), .B0(new_n4571_), .B1(\b[60] ), .Y(new_n13714_));
  OAI21X1  g13458(.A0(new_n4740_), .A1(new_n7339_), .B0(new_n13714_), .Y(new_n13715_));
  AOI21X1  g13459(.A0(new_n7338_), .A1(new_n4375_), .B0(new_n13715_), .Y(new_n13716_));
  XOR2X1   g13460(.A(new_n13716_), .B(\a[47] ), .Y(new_n13717_));
  AND2X1   g13461(.A(new_n13680_), .B(new_n13643_), .Y(new_n13718_));
  AOI21X1  g13462(.A0(new_n13681_), .A1(new_n13639_), .B0(new_n13718_), .Y(new_n13719_));
  NAND2X1  g13463(.A(new_n13679_), .B(new_n13645_), .Y(new_n13720_));
  OAI21X1  g13464(.A0(new_n13678_), .A1(new_n13674_), .B0(new_n13720_), .Y(new_n13721_));
  INVX1    g13465(.A(new_n13654_), .Y(new_n13722_));
  NOR2X1   g13466(.A(new_n13658_), .B(new_n13722_), .Y(new_n13723_));
  AOI21X1  g13467(.A0(new_n13662_), .A1(new_n13660_), .B0(new_n13723_), .Y(new_n13724_));
  AOI22X1  g13468(.A0(new_n7818_), .A1(\b[42] ), .B0(new_n7817_), .B1(\b[43] ), .Y(new_n13725_));
  NOR2X1   g13469(.A(new_n13653_), .B(new_n13652_), .Y(new_n13726_));
  AOI21X1  g13470(.A0(new_n13476_), .A1(new_n3478_), .B0(new_n13726_), .Y(new_n13727_));
  XOR2X1   g13471(.A(new_n13727_), .B(new_n13725_), .Y(new_n13728_));
  AOI22X1  g13472(.A0(new_n7192_), .A1(\b[46] ), .B0(new_n7189_), .B1(\b[45] ), .Y(new_n13729_));
  OAI21X1  g13473(.A0(new_n7627_), .A1(new_n4336_), .B0(new_n13729_), .Y(new_n13730_));
  AOI21X1  g13474(.A0(new_n7187_), .A1(new_n4509_), .B0(new_n13730_), .Y(new_n13731_));
  XOR2X1   g13475(.A(new_n13731_), .B(\a[62] ), .Y(new_n13732_));
  XOR2X1   g13476(.A(new_n13732_), .B(new_n13728_), .Y(new_n13733_));
  INVX1    g13477(.A(new_n13733_), .Y(new_n13734_));
  XOR2X1   g13478(.A(new_n13734_), .B(new_n13724_), .Y(new_n13735_));
  AOI22X1  g13479(.A0(new_n6603_), .A1(\b[49] ), .B0(new_n6600_), .B1(\b[48] ), .Y(new_n13736_));
  OAI21X1  g13480(.A0(new_n6804_), .A1(new_n5039_), .B0(new_n13736_), .Y(new_n13737_));
  AOI21X1  g13481(.A0(new_n6598_), .A1(new_n5038_), .B0(new_n13737_), .Y(new_n13738_));
  XOR2X1   g13482(.A(new_n13738_), .B(\a[59] ), .Y(new_n13739_));
  XOR2X1   g13483(.A(new_n13739_), .B(new_n13735_), .Y(new_n13740_));
  INVX1    g13484(.A(new_n13667_), .Y(new_n13741_));
  NOR2X1   g13485(.A(new_n13671_), .B(new_n13668_), .Y(new_n13742_));
  AOI21X1  g13486(.A0(new_n13741_), .A1(new_n13663_), .B0(new_n13742_), .Y(new_n13743_));
  XOR2X1   g13487(.A(new_n13743_), .B(new_n13740_), .Y(new_n13744_));
  AOI22X1  g13488(.A0(new_n6438_), .A1(\b[52] ), .B0(new_n6437_), .B1(\b[51] ), .Y(new_n13745_));
  OAI21X1  g13489(.A0(new_n6436_), .A1(new_n5234_), .B0(new_n13745_), .Y(new_n13746_));
  AOI21X1  g13490(.A0(new_n6023_), .A1(new_n5590_), .B0(new_n13746_), .Y(new_n13747_));
  XOR2X1   g13491(.A(new_n13747_), .B(\a[56] ), .Y(new_n13748_));
  XOR2X1   g13492(.A(new_n13748_), .B(new_n13744_), .Y(new_n13749_));
  AND2X1   g13493(.A(new_n13671_), .B(new_n13668_), .Y(new_n13750_));
  NOR3X1   g13494(.A(new_n13750_), .B(new_n13742_), .C(new_n13651_), .Y(new_n13751_));
  INVX1    g13495(.A(new_n13673_), .Y(new_n13752_));
  AOI21X1  g13496(.A0(new_n13752_), .A1(new_n13647_), .B0(new_n13751_), .Y(new_n13753_));
  XOR2X1   g13497(.A(new_n13753_), .B(new_n13749_), .Y(new_n13754_));
  AOI22X1  g13498(.A0(new_n5430_), .A1(\b[55] ), .B0(new_n5427_), .B1(\b[54] ), .Y(new_n13755_));
  OAI21X1  g13499(.A0(new_n5891_), .A1(new_n6151_), .B0(new_n13755_), .Y(new_n13756_));
  AOI21X1  g13500(.A0(new_n6150_), .A1(new_n5425_), .B0(new_n13756_), .Y(new_n13757_));
  XOR2X1   g13501(.A(new_n13757_), .B(\a[53] ), .Y(new_n13758_));
  XOR2X1   g13502(.A(new_n13758_), .B(new_n13754_), .Y(new_n13759_));
  XOR2X1   g13503(.A(new_n13759_), .B(new_n13721_), .Y(new_n13760_));
  AOI22X1  g13504(.A0(new_n4880_), .A1(\b[58] ), .B0(new_n4877_), .B1(\b[57] ), .Y(new_n13761_));
  OAI21X1  g13505(.A0(new_n5291_), .A1(new_n6520_), .B0(new_n13761_), .Y(new_n13762_));
  AOI21X1  g13506(.A0(new_n6732_), .A1(new_n4875_), .B0(new_n13762_), .Y(new_n13763_));
  XOR2X1   g13507(.A(new_n13763_), .B(\a[50] ), .Y(new_n13764_));
  XOR2X1   g13508(.A(new_n13764_), .B(new_n13760_), .Y(new_n13765_));
  XOR2X1   g13509(.A(new_n13765_), .B(new_n13719_), .Y(new_n13766_));
  XOR2X1   g13510(.A(new_n13766_), .B(new_n13717_), .Y(new_n13767_));
  INVX1    g13511(.A(new_n13767_), .Y(new_n13768_));
  XOR2X1   g13512(.A(new_n13768_), .B(new_n13713_), .Y(new_n13769_));
  INVX1    g13513(.A(new_n13695_), .Y(new_n13770_));
  NOR2X1   g13514(.A(new_n13699_), .B(new_n13696_), .Y(new_n13771_));
  AOI21X1  g13515(.A0(new_n13770_), .A1(new_n13691_), .B0(new_n13771_), .Y(new_n13772_));
  XOR2X1   g13516(.A(new_n13772_), .B(new_n13769_), .Y(new_n13773_));
  INVX1    g13517(.A(new_n13773_), .Y(new_n13774_));
  NOR2X1   g13518(.A(new_n13704_), .B(new_n13701_), .Y(new_n13775_));
  INVX1    g13519(.A(new_n13775_), .Y(new_n13776_));
  OAI21X1  g13520(.A0(new_n13635_), .A1(new_n13633_), .B0(new_n13705_), .Y(new_n13777_));
  AND2X1   g13521(.A(new_n13777_), .B(new_n13776_), .Y(new_n13778_));
  XOR2X1   g13522(.A(new_n13778_), .B(new_n13774_), .Y(\f[106] ));
  NOR2X1   g13523(.A(new_n13772_), .B(new_n13769_), .Y(new_n13780_));
  AOI21X1  g13524(.A0(new_n13777_), .A1(new_n13776_), .B0(new_n13774_), .Y(new_n13781_));
  OR2X1    g13525(.A(new_n13781_), .B(new_n13780_), .Y(new_n13782_));
  NOR2X1   g13526(.A(new_n13712_), .B(new_n13709_), .Y(new_n13783_));
  AOI21X1  g13527(.A0(new_n13767_), .A1(new_n13713_), .B0(new_n13783_), .Y(new_n13784_));
  INVX1    g13528(.A(new_n13719_), .Y(new_n13785_));
  NOR2X1   g13529(.A(new_n13766_), .B(new_n13717_), .Y(new_n13786_));
  AOI21X1  g13530(.A0(new_n13765_), .A1(new_n13785_), .B0(new_n13786_), .Y(new_n13787_));
  NOR3X1   g13531(.A(new_n4232_), .B(new_n3900_), .C(new_n7772_), .Y(new_n13788_));
  AOI21X1  g13532(.A0(new_n7774_), .A1(new_n3901_), .B0(new_n13788_), .Y(new_n13789_));
  XOR2X1   g13533(.A(new_n13789_), .B(\a[44] ), .Y(new_n13790_));
  XOR2X1   g13534(.A(new_n13790_), .B(new_n13787_), .Y(new_n13791_));
  NOR2X1   g13535(.A(new_n13753_), .B(new_n13749_), .Y(new_n13792_));
  INVX1    g13536(.A(new_n13792_), .Y(new_n13793_));
  INVX1    g13537(.A(new_n13754_), .Y(new_n13794_));
  OAI21X1  g13538(.A0(new_n13758_), .A1(new_n13794_), .B0(new_n13793_), .Y(new_n13795_));
  AOI22X1  g13539(.A0(new_n5430_), .A1(\b[56] ), .B0(new_n5427_), .B1(\b[55] ), .Y(new_n13796_));
  OAI21X1  g13540(.A0(new_n5891_), .A1(new_n6148_), .B0(new_n13796_), .Y(new_n13797_));
  AOI21X1  g13541(.A0(new_n6342_), .A1(new_n5425_), .B0(new_n13797_), .Y(new_n13798_));
  XOR2X1   g13542(.A(new_n13798_), .B(\a[53] ), .Y(new_n13799_));
  NOR2X1   g13543(.A(new_n13743_), .B(new_n13740_), .Y(new_n13800_));
  INVX1    g13544(.A(new_n13800_), .Y(new_n13801_));
  INVX1    g13545(.A(new_n13744_), .Y(new_n13802_));
  OAI21X1  g13546(.A0(new_n13748_), .A1(new_n13802_), .B0(new_n13801_), .Y(new_n13803_));
  INVX1    g13547(.A(new_n13803_), .Y(new_n13804_));
  AOI22X1  g13548(.A0(new_n6438_), .A1(\b[53] ), .B0(new_n6437_), .B1(\b[52] ), .Y(new_n13805_));
  OAI21X1  g13549(.A0(new_n6436_), .A1(new_n5787_), .B0(new_n13805_), .Y(new_n13806_));
  AOI21X1  g13550(.A0(new_n6023_), .A1(new_n5786_), .B0(new_n13806_), .Y(new_n13807_));
  XOR2X1   g13551(.A(new_n13807_), .B(\a[56] ), .Y(new_n13808_));
  NOR2X1   g13552(.A(new_n13734_), .B(new_n13724_), .Y(new_n13809_));
  INVX1    g13553(.A(new_n13809_), .Y(new_n13810_));
  INVX1    g13554(.A(new_n13735_), .Y(new_n13811_));
  OAI21X1  g13555(.A0(new_n13739_), .A1(new_n13811_), .B0(new_n13810_), .Y(new_n13812_));
  INVX1    g13556(.A(new_n13812_), .Y(new_n13813_));
  AOI22X1  g13557(.A0(new_n6603_), .A1(\b[50] ), .B0(new_n6600_), .B1(\b[49] ), .Y(new_n13814_));
  OAI21X1  g13558(.A0(new_n6804_), .A1(new_n5036_), .B0(new_n13814_), .Y(new_n13815_));
  AOI21X1  g13559(.A0(new_n6598_), .A1(new_n5204_), .B0(new_n13815_), .Y(new_n13816_));
  XOR2X1   g13560(.A(new_n13816_), .B(\a[59] ), .Y(new_n13817_));
  INVX1    g13561(.A(new_n13725_), .Y(new_n13818_));
  NOR2X1   g13562(.A(new_n13727_), .B(new_n13818_), .Y(new_n13819_));
  INVX1    g13563(.A(new_n13819_), .Y(new_n13820_));
  OAI21X1  g13564(.A0(new_n13732_), .A1(new_n13728_), .B0(new_n13820_), .Y(new_n13821_));
  INVX1    g13565(.A(new_n13821_), .Y(new_n13822_));
  AOI22X1  g13566(.A0(new_n7818_), .A1(\b[43] ), .B0(new_n7817_), .B1(\b[44] ), .Y(new_n13823_));
  XOR2X1   g13567(.A(new_n13823_), .B(new_n13725_), .Y(new_n13824_));
  AOI22X1  g13568(.A0(new_n7192_), .A1(\b[47] ), .B0(new_n7189_), .B1(\b[46] ), .Y(new_n13825_));
  OAI21X1  g13569(.A0(new_n7627_), .A1(new_n4674_), .B0(new_n13825_), .Y(new_n13826_));
  AOI21X1  g13570(.A0(new_n7187_), .A1(new_n4673_), .B0(new_n13826_), .Y(new_n13827_));
  XOR2X1   g13571(.A(new_n13827_), .B(\a[62] ), .Y(new_n13828_));
  XOR2X1   g13572(.A(new_n13828_), .B(new_n13824_), .Y(new_n13829_));
  XOR2X1   g13573(.A(new_n13829_), .B(new_n13822_), .Y(new_n13830_));
  XOR2X1   g13574(.A(new_n13830_), .B(new_n13817_), .Y(new_n13831_));
  XOR2X1   g13575(.A(new_n13831_), .B(new_n13813_), .Y(new_n13832_));
  XOR2X1   g13576(.A(new_n13832_), .B(new_n13808_), .Y(new_n13833_));
  XOR2X1   g13577(.A(new_n13833_), .B(new_n13804_), .Y(new_n13834_));
  XOR2X1   g13578(.A(new_n13834_), .B(new_n13799_), .Y(new_n13835_));
  XOR2X1   g13579(.A(new_n13835_), .B(new_n13795_), .Y(new_n13836_));
  AOI22X1  g13580(.A0(new_n4880_), .A1(\b[59] ), .B0(new_n4877_), .B1(\b[58] ), .Y(new_n13837_));
  OAI21X1  g13581(.A0(new_n5291_), .A1(new_n6933_), .B0(new_n13837_), .Y(new_n13838_));
  AOI21X1  g13582(.A0(new_n6932_), .A1(new_n4875_), .B0(new_n13838_), .Y(new_n13839_));
  XOR2X1   g13583(.A(new_n13839_), .B(\a[50] ), .Y(new_n13840_));
  XOR2X1   g13584(.A(new_n13840_), .B(new_n13836_), .Y(new_n13841_));
  INVX1    g13585(.A(new_n13759_), .Y(new_n13842_));
  NOR2X1   g13586(.A(new_n13764_), .B(new_n13760_), .Y(new_n13843_));
  AOI21X1  g13587(.A0(new_n13842_), .A1(new_n13721_), .B0(new_n13843_), .Y(new_n13844_));
  XOR2X1   g13588(.A(new_n13844_), .B(new_n13841_), .Y(new_n13845_));
  AOI22X1  g13589(.A0(new_n4572_), .A1(\b[62] ), .B0(new_n4571_), .B1(\b[61] ), .Y(new_n13846_));
  OAI21X1  g13590(.A0(new_n4740_), .A1(new_n7559_), .B0(new_n13846_), .Y(new_n13847_));
  AOI21X1  g13591(.A0(new_n7558_), .A1(new_n4375_), .B0(new_n13847_), .Y(new_n13848_));
  XOR2X1   g13592(.A(new_n13848_), .B(\a[47] ), .Y(new_n13849_));
  XOR2X1   g13593(.A(new_n13849_), .B(new_n13845_), .Y(new_n13850_));
  XOR2X1   g13594(.A(new_n13850_), .B(new_n13791_), .Y(new_n13851_));
  XOR2X1   g13595(.A(new_n13851_), .B(new_n13784_), .Y(new_n13852_));
  XOR2X1   g13596(.A(new_n13852_), .B(new_n13782_), .Y(\f[107] ));
  OR2X1    g13597(.A(new_n13851_), .B(new_n13784_), .Y(new_n13854_));
  OAI21X1  g13598(.A0(new_n13781_), .A1(new_n13780_), .B0(new_n13852_), .Y(new_n13855_));
  NAND2X1  g13599(.A(new_n13855_), .B(new_n13854_), .Y(new_n13856_));
  AND2X1   g13600(.A(new_n13835_), .B(new_n13795_), .Y(new_n13857_));
  INVX1    g13601(.A(new_n13857_), .Y(new_n13858_));
  INVX1    g13602(.A(new_n13836_), .Y(new_n13859_));
  OAI21X1  g13603(.A0(new_n13840_), .A1(new_n13859_), .B0(new_n13858_), .Y(new_n13860_));
  AOI22X1  g13604(.A0(new_n4880_), .A1(\b[60] ), .B0(new_n4877_), .B1(\b[59] ), .Y(new_n13861_));
  OAI21X1  g13605(.A0(new_n5291_), .A1(new_n6930_), .B0(new_n13861_), .Y(new_n13862_));
  AOI21X1  g13606(.A0(new_n6951_), .A1(new_n4875_), .B0(new_n13862_), .Y(new_n13863_));
  XOR2X1   g13607(.A(new_n13863_), .B(new_n4873_), .Y(new_n13864_));
  NAND2X1  g13608(.A(new_n13833_), .B(new_n13803_), .Y(new_n13865_));
  OAI21X1  g13609(.A0(new_n13834_), .A1(new_n13799_), .B0(new_n13865_), .Y(new_n13866_));
  AOI22X1  g13610(.A0(new_n5430_), .A1(\b[57] ), .B0(new_n5427_), .B1(\b[56] ), .Y(new_n13867_));
  OAI21X1  g13611(.A0(new_n5891_), .A1(new_n6523_), .B0(new_n13867_), .Y(new_n13868_));
  AOI21X1  g13612(.A0(new_n6522_), .A1(new_n5425_), .B0(new_n13868_), .Y(new_n13869_));
  XOR2X1   g13613(.A(new_n13869_), .B(new_n5423_), .Y(new_n13870_));
  NAND2X1  g13614(.A(new_n13831_), .B(new_n13812_), .Y(new_n13871_));
  OAI21X1  g13615(.A0(new_n13832_), .A1(new_n13808_), .B0(new_n13871_), .Y(new_n13872_));
  AOI22X1  g13616(.A0(new_n6438_), .A1(\b[54] ), .B0(new_n6437_), .B1(\b[53] ), .Y(new_n13873_));
  OAI21X1  g13617(.A0(new_n6436_), .A1(new_n5808_), .B0(new_n13873_), .Y(new_n13874_));
  AOI21X1  g13618(.A0(new_n6023_), .A1(new_n5807_), .B0(new_n13874_), .Y(new_n13875_));
  XOR2X1   g13619(.A(new_n13875_), .B(new_n6019_), .Y(new_n13876_));
  NAND2X1  g13620(.A(new_n13829_), .B(new_n13821_), .Y(new_n13877_));
  OAI21X1  g13621(.A0(new_n13830_), .A1(new_n13817_), .B0(new_n13877_), .Y(new_n13878_));
  OR2X1    g13622(.A(new_n13823_), .B(new_n13818_), .Y(new_n13879_));
  OAI21X1  g13623(.A0(new_n13828_), .A1(new_n13824_), .B0(new_n13879_), .Y(new_n13880_));
  AOI22X1  g13624(.A0(new_n7818_), .A1(\b[44] ), .B0(new_n7817_), .B1(\b[45] ), .Y(new_n13881_));
  XOR2X1   g13625(.A(new_n13881_), .B(\a[44] ), .Y(new_n13882_));
  XOR2X1   g13626(.A(new_n13882_), .B(new_n13725_), .Y(new_n13883_));
  XOR2X1   g13627(.A(new_n13883_), .B(new_n13880_), .Y(new_n13884_));
  AOI22X1  g13628(.A0(new_n7192_), .A1(\b[48] ), .B0(new_n7189_), .B1(\b[47] ), .Y(new_n13885_));
  OAI21X1  g13629(.A0(new_n7627_), .A1(new_n4693_), .B0(new_n13885_), .Y(new_n13886_));
  AOI21X1  g13630(.A0(new_n7187_), .A1(new_n4692_), .B0(new_n13886_), .Y(new_n13887_));
  XOR2X1   g13631(.A(new_n13887_), .B(\a[62] ), .Y(new_n13888_));
  INVX1    g13632(.A(new_n13888_), .Y(new_n13889_));
  XOR2X1   g13633(.A(new_n13889_), .B(new_n13884_), .Y(new_n13890_));
  AOI22X1  g13634(.A0(new_n6603_), .A1(\b[51] ), .B0(new_n6600_), .B1(\b[50] ), .Y(new_n13891_));
  OAI21X1  g13635(.A0(new_n6804_), .A1(new_n5237_), .B0(new_n13891_), .Y(new_n13892_));
  AOI21X1  g13636(.A0(new_n6598_), .A1(new_n5236_), .B0(new_n13892_), .Y(new_n13893_));
  XOR2X1   g13637(.A(new_n13893_), .B(\a[59] ), .Y(new_n13894_));
  XOR2X1   g13638(.A(new_n13894_), .B(new_n13890_), .Y(new_n13895_));
  XOR2X1   g13639(.A(new_n13895_), .B(new_n13878_), .Y(new_n13896_));
  XOR2X1   g13640(.A(new_n13896_), .B(new_n13876_), .Y(new_n13897_));
  XOR2X1   g13641(.A(new_n13897_), .B(new_n13872_), .Y(new_n13898_));
  XOR2X1   g13642(.A(new_n13898_), .B(new_n13870_), .Y(new_n13899_));
  XOR2X1   g13643(.A(new_n13899_), .B(new_n13866_), .Y(new_n13900_));
  XOR2X1   g13644(.A(new_n13900_), .B(new_n13864_), .Y(new_n13901_));
  XOR2X1   g13645(.A(new_n13901_), .B(new_n13860_), .Y(new_n13902_));
  AOI22X1  g13646(.A0(new_n4572_), .A1(\b[63] ), .B0(new_n4571_), .B1(\b[62] ), .Y(new_n13903_));
  OAI21X1  g13647(.A0(new_n4740_), .A1(new_n7748_), .B0(new_n13903_), .Y(new_n13904_));
  AOI21X1  g13648(.A0(new_n7747_), .A1(new_n4375_), .B0(new_n13904_), .Y(new_n13905_));
  XOR2X1   g13649(.A(new_n13905_), .B(\a[47] ), .Y(new_n13906_));
  XOR2X1   g13650(.A(new_n13906_), .B(new_n13902_), .Y(new_n13907_));
  NOR2X1   g13651(.A(new_n13844_), .B(new_n13841_), .Y(new_n13908_));
  INVX1    g13652(.A(new_n13849_), .Y(new_n13909_));
  AOI21X1  g13653(.A0(new_n13909_), .A1(new_n13845_), .B0(new_n13908_), .Y(new_n13910_));
  XOR2X1   g13654(.A(new_n13910_), .B(new_n13907_), .Y(new_n13911_));
  INVX1    g13655(.A(new_n13911_), .Y(new_n13912_));
  NOR2X1   g13656(.A(new_n13790_), .B(new_n13787_), .Y(new_n13913_));
  INVX1    g13657(.A(new_n13850_), .Y(new_n13914_));
  AOI21X1  g13658(.A0(new_n13914_), .A1(new_n13791_), .B0(new_n13913_), .Y(new_n13915_));
  XOR2X1   g13659(.A(new_n13915_), .B(new_n13912_), .Y(new_n13916_));
  XOR2X1   g13660(.A(new_n13916_), .B(new_n13856_), .Y(\f[108] ));
  AND2X1   g13661(.A(new_n13900_), .B(new_n13864_), .Y(new_n13918_));
  AOI21X1  g13662(.A0(new_n13901_), .A1(new_n13860_), .B0(new_n13918_), .Y(new_n13919_));
  OAI22X1  g13663(.A0(new_n4740_), .A1(new_n7745_), .B0(new_n4378_), .B1(new_n7772_), .Y(new_n13920_));
  AOI21X1  g13664(.A0(new_n7775_), .A1(new_n4375_), .B0(new_n13920_), .Y(new_n13921_));
  XOR2X1   g13665(.A(new_n13921_), .B(\a[47] ), .Y(new_n13922_));
  XOR2X1   g13666(.A(new_n13922_), .B(new_n13919_), .Y(new_n13923_));
  AOI22X1  g13667(.A0(new_n4880_), .A1(\b[61] ), .B0(new_n4877_), .B1(\b[60] ), .Y(new_n13924_));
  OAI21X1  g13668(.A0(new_n5291_), .A1(new_n7339_), .B0(new_n13924_), .Y(new_n13925_));
  AOI21X1  g13669(.A0(new_n7338_), .A1(new_n4875_), .B0(new_n13925_), .Y(new_n13926_));
  XOR2X1   g13670(.A(new_n13926_), .B(\a[50] ), .Y(new_n13927_));
  AND2X1   g13671(.A(new_n13898_), .B(new_n13870_), .Y(new_n13928_));
  AOI21X1  g13672(.A0(new_n13899_), .A1(new_n13866_), .B0(new_n13928_), .Y(new_n13929_));
  AND2X1   g13673(.A(new_n13896_), .B(new_n13876_), .Y(new_n13930_));
  AND2X1   g13674(.A(new_n13897_), .B(new_n13872_), .Y(new_n13931_));
  OR2X1    g13675(.A(new_n13931_), .B(new_n13930_), .Y(new_n13932_));
  NOR2X1   g13676(.A(new_n13894_), .B(new_n13890_), .Y(new_n13933_));
  AOI21X1  g13677(.A0(new_n13895_), .A1(new_n13878_), .B0(new_n13933_), .Y(new_n13934_));
  INVX1    g13678(.A(new_n13934_), .Y(new_n13935_));
  AOI22X1  g13679(.A0(new_n6603_), .A1(\b[52] ), .B0(new_n6600_), .B1(\b[51] ), .Y(new_n13936_));
  OAI21X1  g13680(.A0(new_n6804_), .A1(new_n5234_), .B0(new_n13936_), .Y(new_n13937_));
  AOI21X1  g13681(.A0(new_n6598_), .A1(new_n5590_), .B0(new_n13937_), .Y(new_n13938_));
  XOR2X1   g13682(.A(new_n13938_), .B(\a[59] ), .Y(new_n13939_));
  INVX1    g13683(.A(new_n13883_), .Y(new_n13940_));
  AND2X1   g13684(.A(new_n13940_), .B(new_n13880_), .Y(new_n13941_));
  NOR2X1   g13685(.A(new_n13888_), .B(new_n13884_), .Y(new_n13942_));
  NOR2X1   g13686(.A(new_n13942_), .B(new_n13941_), .Y(new_n13943_));
  AOI22X1  g13687(.A0(new_n7818_), .A1(\b[45] ), .B0(new_n7817_), .B1(\b[46] ), .Y(new_n13944_));
  NOR2X1   g13688(.A(new_n13881_), .B(\a[44] ), .Y(new_n13945_));
  AOI21X1  g13689(.A0(new_n13882_), .A1(new_n13818_), .B0(new_n13945_), .Y(new_n13946_));
  XOR2X1   g13690(.A(new_n13946_), .B(new_n13944_), .Y(new_n13947_));
  AOI22X1  g13691(.A0(new_n7192_), .A1(\b[49] ), .B0(new_n7189_), .B1(\b[48] ), .Y(new_n13948_));
  OAI21X1  g13692(.A0(new_n7627_), .A1(new_n5039_), .B0(new_n13948_), .Y(new_n13949_));
  AOI21X1  g13693(.A0(new_n7187_), .A1(new_n5038_), .B0(new_n13949_), .Y(new_n13950_));
  XOR2X1   g13694(.A(new_n13950_), .B(\a[62] ), .Y(new_n13951_));
  XOR2X1   g13695(.A(new_n13951_), .B(new_n13947_), .Y(new_n13952_));
  XOR2X1   g13696(.A(new_n13952_), .B(new_n13943_), .Y(new_n13953_));
  XOR2X1   g13697(.A(new_n13953_), .B(new_n13939_), .Y(new_n13954_));
  XOR2X1   g13698(.A(new_n13954_), .B(new_n13935_), .Y(new_n13955_));
  AOI22X1  g13699(.A0(new_n6438_), .A1(\b[55] ), .B0(new_n6437_), .B1(\b[54] ), .Y(new_n13956_));
  OAI21X1  g13700(.A0(new_n6436_), .A1(new_n6151_), .B0(new_n13956_), .Y(new_n13957_));
  AOI21X1  g13701(.A0(new_n6150_), .A1(new_n6023_), .B0(new_n13957_), .Y(new_n13958_));
  XOR2X1   g13702(.A(new_n13958_), .B(\a[56] ), .Y(new_n13959_));
  XOR2X1   g13703(.A(new_n13959_), .B(new_n13955_), .Y(new_n13960_));
  XOR2X1   g13704(.A(new_n13960_), .B(new_n13932_), .Y(new_n13961_));
  AOI22X1  g13705(.A0(new_n5430_), .A1(\b[58] ), .B0(new_n5427_), .B1(\b[57] ), .Y(new_n13962_));
  OAI21X1  g13706(.A0(new_n5891_), .A1(new_n6520_), .B0(new_n13962_), .Y(new_n13963_));
  AOI21X1  g13707(.A0(new_n6732_), .A1(new_n5425_), .B0(new_n13963_), .Y(new_n13964_));
  XOR2X1   g13708(.A(new_n13964_), .B(\a[53] ), .Y(new_n13965_));
  XOR2X1   g13709(.A(new_n13965_), .B(new_n13961_), .Y(new_n13966_));
  XOR2X1   g13710(.A(new_n13966_), .B(new_n13929_), .Y(new_n13967_));
  XOR2X1   g13711(.A(new_n13967_), .B(new_n13927_), .Y(new_n13968_));
  INVX1    g13712(.A(new_n13968_), .Y(new_n13969_));
  XOR2X1   g13713(.A(new_n13969_), .B(new_n13923_), .Y(new_n13970_));
  INVX1    g13714(.A(new_n13906_), .Y(new_n13971_));
  NOR2X1   g13715(.A(new_n13910_), .B(new_n13907_), .Y(new_n13972_));
  AOI21X1  g13716(.A0(new_n13971_), .A1(new_n13902_), .B0(new_n13972_), .Y(new_n13973_));
  XOR2X1   g13717(.A(new_n13973_), .B(new_n13970_), .Y(new_n13974_));
  NOR2X1   g13718(.A(new_n13915_), .B(new_n13912_), .Y(new_n13975_));
  INVX1    g13719(.A(new_n13916_), .Y(new_n13976_));
  AOI21X1  g13720(.A0(new_n13855_), .A1(new_n13854_), .B0(new_n13976_), .Y(new_n13977_));
  OR2X1    g13721(.A(new_n13977_), .B(new_n13975_), .Y(new_n13978_));
  XOR2X1   g13722(.A(new_n13978_), .B(new_n13974_), .Y(\f[109] ));
  AND2X1   g13723(.A(new_n13954_), .B(new_n13935_), .Y(new_n13980_));
  INVX1    g13724(.A(new_n13980_), .Y(new_n13981_));
  INVX1    g13725(.A(new_n13955_), .Y(new_n13982_));
  OAI21X1  g13726(.A0(new_n13959_), .A1(new_n13982_), .B0(new_n13981_), .Y(new_n13983_));
  AOI22X1  g13727(.A0(new_n6438_), .A1(\b[56] ), .B0(new_n6437_), .B1(\b[55] ), .Y(new_n13984_));
  OAI21X1  g13728(.A0(new_n6436_), .A1(new_n6148_), .B0(new_n13984_), .Y(new_n13985_));
  AOI21X1  g13729(.A0(new_n6342_), .A1(new_n6023_), .B0(new_n13985_), .Y(new_n13986_));
  XOR2X1   g13730(.A(new_n13986_), .B(\a[56] ), .Y(new_n13987_));
  OAI21X1  g13731(.A0(new_n13942_), .A1(new_n13941_), .B0(new_n13952_), .Y(new_n13988_));
  OAI21X1  g13732(.A0(new_n13953_), .A1(new_n13939_), .B0(new_n13988_), .Y(new_n13989_));
  INVX1    g13733(.A(new_n13989_), .Y(new_n13990_));
  AOI22X1  g13734(.A0(new_n6603_), .A1(\b[53] ), .B0(new_n6600_), .B1(\b[52] ), .Y(new_n13991_));
  OAI21X1  g13735(.A0(new_n6804_), .A1(new_n5787_), .B0(new_n13991_), .Y(new_n13992_));
  AOI21X1  g13736(.A0(new_n6598_), .A1(new_n5786_), .B0(new_n13992_), .Y(new_n13993_));
  XOR2X1   g13737(.A(new_n13993_), .B(\a[59] ), .Y(new_n13994_));
  INVX1    g13738(.A(new_n13944_), .Y(new_n13995_));
  OR2X1    g13739(.A(new_n13946_), .B(new_n13995_), .Y(new_n13996_));
  OR2X1    g13740(.A(new_n13951_), .B(new_n13947_), .Y(new_n13997_));
  AND2X1   g13741(.A(new_n13997_), .B(new_n13996_), .Y(new_n13998_));
  AOI22X1  g13742(.A0(new_n7818_), .A1(\b[46] ), .B0(new_n7817_), .B1(\b[47] ), .Y(new_n13999_));
  NOR2X1   g13743(.A(new_n13999_), .B(new_n13995_), .Y(new_n14000_));
  XOR2X1   g13744(.A(new_n13999_), .B(new_n13995_), .Y(new_n14001_));
  NAND2X1  g13745(.A(new_n13999_), .B(new_n13995_), .Y(new_n14002_));
  OAI21X1  g13746(.A0(new_n14000_), .A1(new_n13998_), .B0(new_n14002_), .Y(new_n14003_));
  OAI22X1  g13747(.A0(new_n14003_), .A1(new_n14000_), .B0(new_n14001_), .B1(new_n13998_), .Y(new_n14004_));
  AOI22X1  g13748(.A0(new_n7192_), .A1(\b[50] ), .B0(new_n7189_), .B1(\b[49] ), .Y(new_n14005_));
  OAI21X1  g13749(.A0(new_n7627_), .A1(new_n5036_), .B0(new_n14005_), .Y(new_n14006_));
  AOI21X1  g13750(.A0(new_n7187_), .A1(new_n5204_), .B0(new_n14006_), .Y(new_n14007_));
  XOR2X1   g13751(.A(new_n14007_), .B(\a[62] ), .Y(new_n14008_));
  XOR2X1   g13752(.A(new_n14008_), .B(new_n14004_), .Y(new_n14009_));
  XOR2X1   g13753(.A(new_n14009_), .B(new_n13994_), .Y(new_n14010_));
  XOR2X1   g13754(.A(new_n14010_), .B(new_n13990_), .Y(new_n14011_));
  XOR2X1   g13755(.A(new_n14011_), .B(new_n13987_), .Y(new_n14012_));
  XOR2X1   g13756(.A(new_n14012_), .B(new_n13983_), .Y(new_n14013_));
  AOI22X1  g13757(.A0(new_n5430_), .A1(\b[59] ), .B0(new_n5427_), .B1(\b[58] ), .Y(new_n14014_));
  OAI21X1  g13758(.A0(new_n5891_), .A1(new_n6933_), .B0(new_n14014_), .Y(new_n14015_));
  AOI21X1  g13759(.A0(new_n6932_), .A1(new_n5425_), .B0(new_n14015_), .Y(new_n14016_));
  XOR2X1   g13760(.A(new_n14016_), .B(\a[53] ), .Y(new_n14017_));
  XOR2X1   g13761(.A(new_n14017_), .B(new_n14013_), .Y(new_n14018_));
  INVX1    g13762(.A(new_n13960_), .Y(new_n14019_));
  NOR2X1   g13763(.A(new_n13965_), .B(new_n13961_), .Y(new_n14020_));
  AOI21X1  g13764(.A0(new_n14019_), .A1(new_n13932_), .B0(new_n14020_), .Y(new_n14021_));
  XOR2X1   g13765(.A(new_n14021_), .B(new_n14018_), .Y(new_n14022_));
  AOI22X1  g13766(.A0(new_n4880_), .A1(\b[62] ), .B0(new_n4877_), .B1(\b[61] ), .Y(new_n14023_));
  OAI21X1  g13767(.A0(new_n5291_), .A1(new_n7559_), .B0(new_n14023_), .Y(new_n14024_));
  AOI21X1  g13768(.A0(new_n7558_), .A1(new_n4875_), .B0(new_n14024_), .Y(new_n14025_));
  XOR2X1   g13769(.A(new_n14025_), .B(\a[50] ), .Y(new_n14026_));
  XOR2X1   g13770(.A(new_n14026_), .B(new_n14022_), .Y(new_n14027_));
  INVX1    g13771(.A(new_n13929_), .Y(new_n14028_));
  NOR2X1   g13772(.A(new_n13967_), .B(new_n13927_), .Y(new_n14029_));
  AOI21X1  g13773(.A0(new_n13966_), .A1(new_n14028_), .B0(new_n14029_), .Y(new_n14030_));
  NOR3X1   g13774(.A(new_n4739_), .B(new_n4379_), .C(new_n7772_), .Y(new_n14031_));
  AOI21X1  g13775(.A0(new_n7774_), .A1(new_n4375_), .B0(new_n14031_), .Y(new_n14032_));
  XOR2X1   g13776(.A(new_n14032_), .B(\a[47] ), .Y(new_n14033_));
  XOR2X1   g13777(.A(new_n14033_), .B(new_n14030_), .Y(new_n14034_));
  XOR2X1   g13778(.A(new_n14034_), .B(new_n14027_), .Y(new_n14035_));
  NOR2X1   g13779(.A(new_n13922_), .B(new_n13919_), .Y(new_n14036_));
  AOI21X1  g13780(.A0(new_n13968_), .A1(new_n13923_), .B0(new_n14036_), .Y(new_n14037_));
  XOR2X1   g13781(.A(new_n14037_), .B(new_n14035_), .Y(new_n14038_));
  INVX1    g13782(.A(new_n14038_), .Y(new_n14039_));
  NOR2X1   g13783(.A(new_n13973_), .B(new_n13970_), .Y(new_n14040_));
  INVX1    g13784(.A(new_n14040_), .Y(new_n14041_));
  OAI21X1  g13785(.A0(new_n13977_), .A1(new_n13975_), .B0(new_n13974_), .Y(new_n14042_));
  AND2X1   g13786(.A(new_n14042_), .B(new_n14041_), .Y(new_n14043_));
  XOR2X1   g13787(.A(new_n14043_), .B(new_n14039_), .Y(\f[110] ));
  AND2X1   g13788(.A(new_n14012_), .B(new_n13983_), .Y(new_n14045_));
  INVX1    g13789(.A(new_n14045_), .Y(new_n14046_));
  INVX1    g13790(.A(new_n14013_), .Y(new_n14047_));
  OAI21X1  g13791(.A0(new_n14017_), .A1(new_n14047_), .B0(new_n14046_), .Y(new_n14048_));
  AOI22X1  g13792(.A0(new_n5430_), .A1(\b[60] ), .B0(new_n5427_), .B1(\b[59] ), .Y(new_n14049_));
  OAI21X1  g13793(.A0(new_n5891_), .A1(new_n6930_), .B0(new_n14049_), .Y(new_n14050_));
  AOI21X1  g13794(.A0(new_n6951_), .A1(new_n5425_), .B0(new_n14050_), .Y(new_n14051_));
  XOR2X1   g13795(.A(new_n14051_), .B(new_n5423_), .Y(new_n14052_));
  NAND2X1  g13796(.A(new_n14010_), .B(new_n13989_), .Y(new_n14053_));
  OAI21X1  g13797(.A0(new_n14011_), .A1(new_n13987_), .B0(new_n14053_), .Y(new_n14054_));
  AOI22X1  g13798(.A0(new_n6438_), .A1(\b[57] ), .B0(new_n6437_), .B1(\b[56] ), .Y(new_n14055_));
  OAI21X1  g13799(.A0(new_n6436_), .A1(new_n6523_), .B0(new_n14055_), .Y(new_n14056_));
  AOI21X1  g13800(.A0(new_n6522_), .A1(new_n6023_), .B0(new_n14056_), .Y(new_n14057_));
  XOR2X1   g13801(.A(new_n14057_), .B(new_n6019_), .Y(new_n14058_));
  INVX1    g13802(.A(new_n14008_), .Y(new_n14059_));
  NOR2X1   g13803(.A(new_n14009_), .B(new_n13994_), .Y(new_n14060_));
  AOI21X1  g13804(.A0(new_n14059_), .A1(new_n14004_), .B0(new_n14060_), .Y(new_n14061_));
  AOI22X1  g13805(.A0(new_n7192_), .A1(\b[51] ), .B0(new_n7189_), .B1(\b[50] ), .Y(new_n14062_));
  OAI21X1  g13806(.A0(new_n7627_), .A1(new_n5237_), .B0(new_n14062_), .Y(new_n14063_));
  AOI21X1  g13807(.A0(new_n7187_), .A1(new_n5236_), .B0(new_n14063_), .Y(new_n14064_));
  XOR2X1   g13808(.A(new_n14064_), .B(\a[62] ), .Y(new_n14065_));
  AOI22X1  g13809(.A0(new_n7818_), .A1(\b[47] ), .B0(new_n7817_), .B1(\b[48] ), .Y(new_n14066_));
  XOR2X1   g13810(.A(new_n13999_), .B(new_n4568_), .Y(new_n14067_));
  XOR2X1   g13811(.A(new_n14067_), .B(new_n14066_), .Y(new_n14068_));
  XOR2X1   g13812(.A(new_n14068_), .B(new_n14065_), .Y(new_n14069_));
  XOR2X1   g13813(.A(new_n14069_), .B(new_n14003_), .Y(new_n14070_));
  INVX1    g13814(.A(new_n14070_), .Y(new_n14071_));
  AOI22X1  g13815(.A0(new_n6603_), .A1(\b[54] ), .B0(new_n6600_), .B1(\b[53] ), .Y(new_n14072_));
  OAI21X1  g13816(.A0(new_n6804_), .A1(new_n5808_), .B0(new_n14072_), .Y(new_n14073_));
  AOI21X1  g13817(.A0(new_n6598_), .A1(new_n5807_), .B0(new_n14073_), .Y(new_n14074_));
  XOR2X1   g13818(.A(new_n14074_), .B(\a[59] ), .Y(new_n14075_));
  XOR2X1   g13819(.A(new_n14075_), .B(new_n14071_), .Y(new_n14076_));
  XOR2X1   g13820(.A(new_n14076_), .B(new_n14061_), .Y(new_n14077_));
  XOR2X1   g13821(.A(new_n14077_), .B(new_n14058_), .Y(new_n14078_));
  XOR2X1   g13822(.A(new_n14078_), .B(new_n14054_), .Y(new_n14079_));
  XOR2X1   g13823(.A(new_n14079_), .B(new_n14052_), .Y(new_n14080_));
  XOR2X1   g13824(.A(new_n14080_), .B(new_n14048_), .Y(new_n14081_));
  AOI22X1  g13825(.A0(new_n4880_), .A1(\b[63] ), .B0(new_n4877_), .B1(\b[62] ), .Y(new_n14082_));
  OAI21X1  g13826(.A0(new_n5291_), .A1(new_n7748_), .B0(new_n14082_), .Y(new_n14083_));
  AOI21X1  g13827(.A0(new_n7747_), .A1(new_n4875_), .B0(new_n14083_), .Y(new_n14084_));
  XOR2X1   g13828(.A(new_n14084_), .B(\a[50] ), .Y(new_n14085_));
  XOR2X1   g13829(.A(new_n14085_), .B(new_n14081_), .Y(new_n14086_));
  NOR2X1   g13830(.A(new_n14021_), .B(new_n14018_), .Y(new_n14087_));
  INVX1    g13831(.A(new_n14026_), .Y(new_n14088_));
  AOI21X1  g13832(.A0(new_n14088_), .A1(new_n14022_), .B0(new_n14087_), .Y(new_n14089_));
  XOR2X1   g13833(.A(new_n14089_), .B(new_n14086_), .Y(new_n14090_));
  INVX1    g13834(.A(new_n14090_), .Y(new_n14091_));
  INVX1    g13835(.A(new_n14027_), .Y(new_n14092_));
  NOR2X1   g13836(.A(new_n14033_), .B(new_n14030_), .Y(new_n14093_));
  AOI21X1  g13837(.A0(new_n14034_), .A1(new_n14092_), .B0(new_n14093_), .Y(new_n14094_));
  XOR2X1   g13838(.A(new_n14094_), .B(new_n14091_), .Y(new_n14095_));
  NOR2X1   g13839(.A(new_n14037_), .B(new_n14035_), .Y(new_n14096_));
  AOI21X1  g13840(.A0(new_n14042_), .A1(new_n14041_), .B0(new_n14039_), .Y(new_n14097_));
  OR2X1    g13841(.A(new_n14097_), .B(new_n14096_), .Y(new_n14098_));
  XOR2X1   g13842(.A(new_n14098_), .B(new_n14095_), .Y(\f[111] ));
  AND2X1   g13843(.A(new_n14079_), .B(new_n14052_), .Y(new_n14100_));
  AOI21X1  g13844(.A0(new_n14080_), .A1(new_n14048_), .B0(new_n14100_), .Y(new_n14101_));
  INVX1    g13845(.A(new_n14101_), .Y(new_n14102_));
  AOI22X1  g13846(.A0(new_n5430_), .A1(\b[61] ), .B0(new_n5427_), .B1(\b[60] ), .Y(new_n14103_));
  OAI21X1  g13847(.A0(new_n5891_), .A1(new_n7339_), .B0(new_n14103_), .Y(new_n14104_));
  AOI21X1  g13848(.A0(new_n7338_), .A1(new_n5425_), .B0(new_n14104_), .Y(new_n14105_));
  XOR2X1   g13849(.A(new_n14105_), .B(\a[53] ), .Y(new_n14106_));
  AND2X1   g13850(.A(new_n14077_), .B(new_n14058_), .Y(new_n14107_));
  AOI21X1  g13851(.A0(new_n14078_), .A1(new_n14054_), .B0(new_n14107_), .Y(new_n14108_));
  AOI22X1  g13852(.A0(new_n6438_), .A1(\b[58] ), .B0(new_n6437_), .B1(\b[57] ), .Y(new_n14109_));
  OAI21X1  g13853(.A0(new_n6436_), .A1(new_n6520_), .B0(new_n14109_), .Y(new_n14110_));
  AOI21X1  g13854(.A0(new_n6732_), .A1(new_n6023_), .B0(new_n14110_), .Y(new_n14111_));
  XOR2X1   g13855(.A(new_n14111_), .B(new_n6019_), .Y(new_n14112_));
  OR2X1    g13856(.A(new_n14075_), .B(new_n14070_), .Y(new_n14113_));
  OAI21X1  g13857(.A0(new_n14076_), .A1(new_n14061_), .B0(new_n14113_), .Y(new_n14114_));
  AOI22X1  g13858(.A0(new_n6603_), .A1(\b[55] ), .B0(new_n6600_), .B1(\b[54] ), .Y(new_n14115_));
  OAI21X1  g13859(.A0(new_n6804_), .A1(new_n6151_), .B0(new_n14115_), .Y(new_n14116_));
  AOI21X1  g13860(.A0(new_n6598_), .A1(new_n6150_), .B0(new_n14116_), .Y(new_n14117_));
  XOR2X1   g13861(.A(new_n14117_), .B(\a[59] ), .Y(new_n14118_));
  INVX1    g13862(.A(new_n14065_), .Y(new_n14119_));
  AND2X1   g13863(.A(new_n14068_), .B(new_n14119_), .Y(new_n14120_));
  INVX1    g13864(.A(new_n14069_), .Y(new_n14121_));
  AOI21X1  g13865(.A0(new_n14121_), .A1(new_n14003_), .B0(new_n14120_), .Y(new_n14122_));
  AOI22X1  g13866(.A0(new_n7818_), .A1(\b[48] ), .B0(new_n7817_), .B1(\b[49] ), .Y(new_n14123_));
  INVX1    g13867(.A(new_n14123_), .Y(new_n14124_));
  OR2X1    g13868(.A(new_n14067_), .B(new_n14066_), .Y(new_n14125_));
  OR2X1    g13869(.A(new_n13999_), .B(\a[47] ), .Y(new_n14126_));
  AND2X1   g13870(.A(new_n14126_), .B(new_n14125_), .Y(new_n14127_));
  XOR2X1   g13871(.A(new_n14127_), .B(new_n14124_), .Y(new_n14128_));
  INVX1    g13872(.A(new_n14128_), .Y(new_n14129_));
  AOI22X1  g13873(.A0(new_n7192_), .A1(\b[52] ), .B0(new_n7189_), .B1(\b[51] ), .Y(new_n14130_));
  OAI21X1  g13874(.A0(new_n7627_), .A1(new_n5234_), .B0(new_n14130_), .Y(new_n14131_));
  AOI21X1  g13875(.A0(new_n7187_), .A1(new_n5590_), .B0(new_n14131_), .Y(new_n14132_));
  XOR2X1   g13876(.A(new_n14132_), .B(\a[62] ), .Y(new_n14133_));
  XOR2X1   g13877(.A(new_n14133_), .B(new_n14129_), .Y(new_n14134_));
  XOR2X1   g13878(.A(new_n14134_), .B(new_n14122_), .Y(new_n14135_));
  XOR2X1   g13879(.A(new_n14135_), .B(new_n14118_), .Y(new_n14136_));
  XOR2X1   g13880(.A(new_n14136_), .B(new_n14114_), .Y(new_n14137_));
  XOR2X1   g13881(.A(new_n14137_), .B(new_n14112_), .Y(new_n14138_));
  XOR2X1   g13882(.A(new_n14138_), .B(new_n14108_), .Y(new_n14139_));
  XOR2X1   g13883(.A(new_n14139_), .B(new_n14106_), .Y(new_n14140_));
  XOR2X1   g13884(.A(new_n14140_), .B(new_n14102_), .Y(new_n14141_));
  OAI22X1  g13885(.A0(new_n5291_), .A1(new_n7745_), .B0(new_n4878_), .B1(new_n7772_), .Y(new_n14142_));
  AOI21X1  g13886(.A0(new_n7775_), .A1(new_n4875_), .B0(new_n14142_), .Y(new_n14143_));
  XOR2X1   g13887(.A(new_n14143_), .B(\a[50] ), .Y(new_n14144_));
  XOR2X1   g13888(.A(new_n14144_), .B(new_n14141_), .Y(new_n14145_));
  INVX1    g13889(.A(new_n14085_), .Y(new_n14146_));
  NOR2X1   g13890(.A(new_n14089_), .B(new_n14086_), .Y(new_n14147_));
  AOI21X1  g13891(.A0(new_n14146_), .A1(new_n14081_), .B0(new_n14147_), .Y(new_n14148_));
  XOR2X1   g13892(.A(new_n14148_), .B(new_n14145_), .Y(new_n14149_));
  INVX1    g13893(.A(new_n14149_), .Y(new_n14150_));
  NOR2X1   g13894(.A(new_n14094_), .B(new_n14091_), .Y(new_n14151_));
  INVX1    g13895(.A(new_n14151_), .Y(new_n14152_));
  OAI21X1  g13896(.A0(new_n14097_), .A1(new_n14096_), .B0(new_n14095_), .Y(new_n14153_));
  AND2X1   g13897(.A(new_n14153_), .B(new_n14152_), .Y(new_n14154_));
  XOR2X1   g13898(.A(new_n14154_), .B(new_n14150_), .Y(\f[112] ));
  INVX1    g13899(.A(new_n14134_), .Y(new_n14156_));
  NOR2X1   g13900(.A(new_n14156_), .B(new_n14122_), .Y(new_n14157_));
  NOR2X1   g13901(.A(new_n14135_), .B(new_n14118_), .Y(new_n14158_));
  NOR2X1   g13902(.A(new_n14158_), .B(new_n14157_), .Y(new_n14159_));
  INVX1    g13903(.A(new_n14159_), .Y(new_n14160_));
  AOI22X1  g13904(.A0(new_n7192_), .A1(\b[53] ), .B0(new_n7189_), .B1(\b[52] ), .Y(new_n14161_));
  OAI21X1  g13905(.A0(new_n7627_), .A1(new_n5787_), .B0(new_n14161_), .Y(new_n14162_));
  AOI21X1  g13906(.A0(new_n7187_), .A1(new_n5786_), .B0(new_n14162_), .Y(new_n14163_));
  XOR2X1   g13907(.A(new_n14163_), .B(\a[62] ), .Y(new_n14164_));
  AOI22X1  g13908(.A0(new_n7818_), .A1(\b[49] ), .B0(new_n7817_), .B1(\b[50] ), .Y(new_n14165_));
  XOR2X1   g13909(.A(new_n14165_), .B(new_n14123_), .Y(new_n14166_));
  XOR2X1   g13910(.A(new_n14166_), .B(new_n14164_), .Y(new_n14167_));
  INVX1    g13911(.A(new_n14167_), .Y(new_n14168_));
  OR2X1    g13912(.A(new_n14127_), .B(new_n14124_), .Y(new_n14169_));
  OAI21X1  g13913(.A0(new_n14133_), .A1(new_n14129_), .B0(new_n14169_), .Y(new_n14170_));
  XOR2X1   g13914(.A(new_n14170_), .B(new_n14168_), .Y(new_n14171_));
  AOI22X1  g13915(.A0(new_n6603_), .A1(\b[56] ), .B0(new_n6600_), .B1(\b[55] ), .Y(new_n14172_));
  OAI21X1  g13916(.A0(new_n6804_), .A1(new_n6148_), .B0(new_n14172_), .Y(new_n14173_));
  AOI21X1  g13917(.A0(new_n6598_), .A1(new_n6342_), .B0(new_n14173_), .Y(new_n14174_));
  XOR2X1   g13918(.A(new_n14174_), .B(\a[59] ), .Y(new_n14175_));
  XOR2X1   g13919(.A(new_n14175_), .B(new_n14171_), .Y(new_n14176_));
  XOR2X1   g13920(.A(new_n14176_), .B(new_n14160_), .Y(new_n14177_));
  AOI22X1  g13921(.A0(new_n6438_), .A1(\b[59] ), .B0(new_n6437_), .B1(\b[58] ), .Y(new_n14178_));
  OAI21X1  g13922(.A0(new_n6436_), .A1(new_n6933_), .B0(new_n14178_), .Y(new_n14179_));
  AOI21X1  g13923(.A0(new_n6932_), .A1(new_n6023_), .B0(new_n14179_), .Y(new_n14180_));
  XOR2X1   g13924(.A(new_n14180_), .B(\a[56] ), .Y(new_n14181_));
  XOR2X1   g13925(.A(new_n14181_), .B(new_n14177_), .Y(new_n14182_));
  AND2X1   g13926(.A(new_n14136_), .B(new_n14114_), .Y(new_n14183_));
  AOI21X1  g13927(.A0(new_n14137_), .A1(new_n14112_), .B0(new_n14183_), .Y(new_n14184_));
  XOR2X1   g13928(.A(new_n14184_), .B(new_n14182_), .Y(new_n14185_));
  AOI22X1  g13929(.A0(new_n5430_), .A1(\b[62] ), .B0(new_n5427_), .B1(\b[61] ), .Y(new_n14186_));
  OAI21X1  g13930(.A0(new_n5891_), .A1(new_n7559_), .B0(new_n14186_), .Y(new_n14187_));
  AOI21X1  g13931(.A0(new_n7558_), .A1(new_n5425_), .B0(new_n14187_), .Y(new_n14188_));
  XOR2X1   g13932(.A(new_n14188_), .B(\a[53] ), .Y(new_n14189_));
  XOR2X1   g13933(.A(new_n14189_), .B(new_n14185_), .Y(new_n14190_));
  INVX1    g13934(.A(new_n14108_), .Y(new_n14191_));
  NOR2X1   g13935(.A(new_n14139_), .B(new_n14106_), .Y(new_n14192_));
  AOI21X1  g13936(.A0(new_n14138_), .A1(new_n14191_), .B0(new_n14192_), .Y(new_n14193_));
  NOR4X1   g13937(.A(new_n4876_), .B(new_n4874_), .C(new_n4879_), .D(new_n7772_), .Y(new_n14194_));
  AOI21X1  g13938(.A0(new_n7774_), .A1(new_n4875_), .B0(new_n14194_), .Y(new_n14195_));
  XOR2X1   g13939(.A(new_n14195_), .B(\a[50] ), .Y(new_n14196_));
  XOR2X1   g13940(.A(new_n14196_), .B(new_n14193_), .Y(new_n14197_));
  XOR2X1   g13941(.A(new_n14197_), .B(new_n14190_), .Y(new_n14198_));
  AND2X1   g13942(.A(new_n14140_), .B(new_n14102_), .Y(new_n14199_));
  INVX1    g13943(.A(new_n14144_), .Y(new_n14200_));
  AOI21X1  g13944(.A0(new_n14200_), .A1(new_n14141_), .B0(new_n14199_), .Y(new_n14201_));
  XOR2X1   g13945(.A(new_n14201_), .B(new_n14198_), .Y(new_n14202_));
  NOR2X1   g13946(.A(new_n14148_), .B(new_n14145_), .Y(new_n14203_));
  AOI21X1  g13947(.A0(new_n14153_), .A1(new_n14152_), .B0(new_n14150_), .Y(new_n14204_));
  OR2X1    g13948(.A(new_n14204_), .B(new_n14203_), .Y(new_n14205_));
  XOR2X1   g13949(.A(new_n14205_), .B(new_n14202_), .Y(\f[113] ));
  AND2X1   g13950(.A(new_n14176_), .B(new_n14160_), .Y(new_n14207_));
  INVX1    g13951(.A(new_n14207_), .Y(new_n14208_));
  INVX1    g13952(.A(new_n14177_), .Y(new_n14209_));
  OAI21X1  g13953(.A0(new_n14181_), .A1(new_n14209_), .B0(new_n14208_), .Y(new_n14210_));
  AOI22X1  g13954(.A0(new_n6438_), .A1(\b[60] ), .B0(new_n6437_), .B1(\b[59] ), .Y(new_n14211_));
  OAI21X1  g13955(.A0(new_n6436_), .A1(new_n6930_), .B0(new_n14211_), .Y(new_n14212_));
  AOI21X1  g13956(.A0(new_n6951_), .A1(new_n6023_), .B0(new_n14212_), .Y(new_n14213_));
  XOR2X1   g13957(.A(new_n14213_), .B(\a[56] ), .Y(new_n14214_));
  NOR2X1   g13958(.A(new_n14175_), .B(new_n14171_), .Y(new_n14215_));
  AOI21X1  g13959(.A0(new_n14170_), .A1(new_n14167_), .B0(new_n14215_), .Y(new_n14216_));
  AOI22X1  g13960(.A0(new_n6603_), .A1(\b[57] ), .B0(new_n6600_), .B1(\b[56] ), .Y(new_n14217_));
  OAI21X1  g13961(.A0(new_n6804_), .A1(new_n6523_), .B0(new_n14217_), .Y(new_n14218_));
  AOI21X1  g13962(.A0(new_n6598_), .A1(new_n6522_), .B0(new_n14218_), .Y(new_n14219_));
  XOR2X1   g13963(.A(new_n14219_), .B(\a[59] ), .Y(new_n14220_));
  AOI22X1  g13964(.A0(new_n7192_), .A1(\b[54] ), .B0(new_n7189_), .B1(\b[53] ), .Y(new_n14221_));
  OAI21X1  g13965(.A0(new_n7627_), .A1(new_n5808_), .B0(new_n14221_), .Y(new_n14222_));
  AOI21X1  g13966(.A0(new_n7187_), .A1(new_n5807_), .B0(new_n14222_), .Y(new_n14223_));
  XOR2X1   g13967(.A(new_n14223_), .B(new_n7185_), .Y(new_n14224_));
  OR2X1    g13968(.A(new_n14165_), .B(new_n14124_), .Y(new_n14225_));
  OAI21X1  g13969(.A0(new_n14166_), .A1(new_n14164_), .B0(new_n14225_), .Y(new_n14226_));
  AOI22X1  g13970(.A0(new_n7818_), .A1(\b[50] ), .B0(new_n7817_), .B1(\b[51] ), .Y(new_n14227_));
  XOR2X1   g13971(.A(new_n14227_), .B(\a[50] ), .Y(new_n14228_));
  XOR2X1   g13972(.A(new_n14228_), .B(new_n14124_), .Y(new_n14229_));
  INVX1    g13973(.A(new_n14229_), .Y(new_n14230_));
  OR2X1    g13974(.A(new_n14230_), .B(new_n14226_), .Y(new_n14231_));
  XOR2X1   g13975(.A(new_n14229_), .B(new_n14226_), .Y(new_n14232_));
  AOI21X1  g13976(.A0(new_n14230_), .A1(new_n14226_), .B0(new_n14224_), .Y(new_n14233_));
  AOI22X1  g13977(.A0(new_n14233_), .A1(new_n14231_), .B0(new_n14232_), .B1(new_n14224_), .Y(new_n14234_));
  AND2X1   g13978(.A(new_n14234_), .B(new_n14220_), .Y(new_n14235_));
  XOR2X1   g13979(.A(new_n14234_), .B(new_n14220_), .Y(new_n14236_));
  OAI21X1  g13980(.A0(new_n14234_), .A1(new_n14220_), .B0(new_n14216_), .Y(new_n14237_));
  OAI22X1  g13981(.A0(new_n14237_), .A1(new_n14235_), .B0(new_n14236_), .B1(new_n14216_), .Y(new_n14238_));
  XOR2X1   g13982(.A(new_n14238_), .B(new_n14214_), .Y(new_n14239_));
  XOR2X1   g13983(.A(new_n14239_), .B(new_n14210_), .Y(new_n14240_));
  AOI22X1  g13984(.A0(new_n5430_), .A1(\b[63] ), .B0(new_n5427_), .B1(\b[62] ), .Y(new_n14241_));
  OAI21X1  g13985(.A0(new_n5891_), .A1(new_n7748_), .B0(new_n14241_), .Y(new_n14242_));
  AOI21X1  g13986(.A0(new_n7747_), .A1(new_n5425_), .B0(new_n14242_), .Y(new_n14243_));
  XOR2X1   g13987(.A(new_n14243_), .B(\a[53] ), .Y(new_n14244_));
  XOR2X1   g13988(.A(new_n14244_), .B(new_n14240_), .Y(new_n14245_));
  NOR2X1   g13989(.A(new_n14184_), .B(new_n14182_), .Y(new_n14246_));
  INVX1    g13990(.A(new_n14189_), .Y(new_n14247_));
  AOI21X1  g13991(.A0(new_n14247_), .A1(new_n14185_), .B0(new_n14246_), .Y(new_n14248_));
  XOR2X1   g13992(.A(new_n14248_), .B(new_n14245_), .Y(new_n14249_));
  INVX1    g13993(.A(new_n14190_), .Y(new_n14250_));
  NOR2X1   g13994(.A(new_n14196_), .B(new_n14193_), .Y(new_n14251_));
  AOI21X1  g13995(.A0(new_n14197_), .A1(new_n14250_), .B0(new_n14251_), .Y(new_n14252_));
  XOR2X1   g13996(.A(new_n14252_), .B(new_n14249_), .Y(new_n14253_));
  OR2X1    g13997(.A(new_n14201_), .B(new_n14198_), .Y(new_n14254_));
  OAI21X1  g13998(.A0(new_n14204_), .A1(new_n14203_), .B0(new_n14202_), .Y(new_n14255_));
  AND2X1   g13999(.A(new_n14255_), .B(new_n14254_), .Y(new_n14256_));
  XOR2X1   g14000(.A(new_n14256_), .B(new_n14253_), .Y(\f[114] ));
  NOR2X1   g14001(.A(new_n14238_), .B(new_n14214_), .Y(new_n14258_));
  AOI21X1  g14002(.A0(new_n14239_), .A1(new_n14210_), .B0(new_n14258_), .Y(new_n14259_));
  INVX1    g14003(.A(new_n14259_), .Y(new_n14260_));
  AOI22X1  g14004(.A0(new_n6438_), .A1(\b[61] ), .B0(new_n6437_), .B1(\b[60] ), .Y(new_n14261_));
  OAI21X1  g14005(.A0(new_n6436_), .A1(new_n7339_), .B0(new_n14261_), .Y(new_n14262_));
  AOI21X1  g14006(.A0(new_n7338_), .A1(new_n6023_), .B0(new_n14262_), .Y(new_n14263_));
  XOR2X1   g14007(.A(new_n14263_), .B(\a[56] ), .Y(new_n14264_));
  INVX1    g14008(.A(new_n14220_), .Y(new_n14265_));
  AND2X1   g14009(.A(new_n14234_), .B(new_n14265_), .Y(new_n14266_));
  NOR2X1   g14010(.A(new_n14236_), .B(new_n14216_), .Y(new_n14267_));
  NOR2X1   g14011(.A(new_n14267_), .B(new_n14266_), .Y(new_n14268_));
  AOI22X1  g14012(.A0(new_n6603_), .A1(\b[58] ), .B0(new_n6600_), .B1(\b[57] ), .Y(new_n14269_));
  OAI21X1  g14013(.A0(new_n6804_), .A1(new_n6520_), .B0(new_n14269_), .Y(new_n14270_));
  AOI21X1  g14014(.A0(new_n6732_), .A1(new_n6598_), .B0(new_n14270_), .Y(new_n14271_));
  XOR2X1   g14015(.A(new_n14271_), .B(new_n6596_), .Y(new_n14272_));
  AND2X1   g14016(.A(new_n14229_), .B(new_n14226_), .Y(new_n14273_));
  AOI21X1  g14017(.A0(new_n14232_), .A1(new_n14224_), .B0(new_n14273_), .Y(new_n14274_));
  AOI22X1  g14018(.A0(new_n7818_), .A1(\b[51] ), .B0(new_n7817_), .B1(\b[52] ), .Y(new_n14275_));
  INVX1    g14019(.A(new_n14275_), .Y(new_n14276_));
  NOR2X1   g14020(.A(new_n14227_), .B(\a[50] ), .Y(new_n14277_));
  AOI21X1  g14021(.A0(new_n14228_), .A1(new_n14124_), .B0(new_n14277_), .Y(new_n14278_));
  XOR2X1   g14022(.A(new_n14278_), .B(new_n14276_), .Y(new_n14279_));
  AOI22X1  g14023(.A0(new_n7192_), .A1(\b[55] ), .B0(new_n7189_), .B1(\b[54] ), .Y(new_n14280_));
  OAI21X1  g14024(.A0(new_n7627_), .A1(new_n6151_), .B0(new_n14280_), .Y(new_n14281_));
  AOI21X1  g14025(.A0(new_n7187_), .A1(new_n6150_), .B0(new_n14281_), .Y(new_n14282_));
  XOR2X1   g14026(.A(new_n14282_), .B(\a[62] ), .Y(new_n14283_));
  XOR2X1   g14027(.A(new_n14283_), .B(new_n14279_), .Y(new_n14284_));
  XOR2X1   g14028(.A(new_n14284_), .B(new_n14274_), .Y(new_n14285_));
  XOR2X1   g14029(.A(new_n14285_), .B(new_n14272_), .Y(new_n14286_));
  XOR2X1   g14030(.A(new_n14286_), .B(new_n14268_), .Y(new_n14287_));
  XOR2X1   g14031(.A(new_n14287_), .B(new_n14264_), .Y(new_n14288_));
  XOR2X1   g14032(.A(new_n14288_), .B(new_n14260_), .Y(new_n14289_));
  OAI22X1  g14033(.A0(new_n5891_), .A1(new_n7745_), .B0(new_n5428_), .B1(new_n7772_), .Y(new_n14290_));
  AOI21X1  g14034(.A0(new_n7775_), .A1(new_n5425_), .B0(new_n14290_), .Y(new_n14291_));
  XOR2X1   g14035(.A(new_n14291_), .B(\a[53] ), .Y(new_n14292_));
  XOR2X1   g14036(.A(new_n14292_), .B(new_n14289_), .Y(new_n14293_));
  INVX1    g14037(.A(new_n14244_), .Y(new_n14294_));
  NOR2X1   g14038(.A(new_n14248_), .B(new_n14245_), .Y(new_n14295_));
  AOI21X1  g14039(.A0(new_n14294_), .A1(new_n14240_), .B0(new_n14295_), .Y(new_n14296_));
  XOR2X1   g14040(.A(new_n14296_), .B(new_n14293_), .Y(new_n14297_));
  AND2X1   g14041(.A(new_n14248_), .B(new_n14245_), .Y(new_n14298_));
  NOR3X1   g14042(.A(new_n14252_), .B(new_n14295_), .C(new_n14298_), .Y(new_n14299_));
  AOI21X1  g14043(.A0(new_n14255_), .A1(new_n14254_), .B0(new_n14253_), .Y(new_n14300_));
  OR2X1    g14044(.A(new_n14300_), .B(new_n14299_), .Y(new_n14301_));
  XOR2X1   g14045(.A(new_n14301_), .B(new_n14297_), .Y(\f[115] ));
  NOR2X1   g14046(.A(new_n14284_), .B(new_n14274_), .Y(new_n14303_));
  AOI21X1  g14047(.A0(new_n14285_), .A1(new_n14272_), .B0(new_n14303_), .Y(new_n14304_));
  INVX1    g14048(.A(new_n14304_), .Y(new_n14305_));
  NOR2X1   g14049(.A(new_n14278_), .B(new_n14276_), .Y(new_n14306_));
  INVX1    g14050(.A(new_n14283_), .Y(new_n14307_));
  AOI21X1  g14051(.A0(new_n14307_), .A1(new_n14279_), .B0(new_n14306_), .Y(new_n14308_));
  AOI22X1  g14052(.A0(new_n7818_), .A1(\b[52] ), .B0(new_n7817_), .B1(\b[53] ), .Y(new_n14309_));
  NOR2X1   g14053(.A(new_n14309_), .B(new_n14276_), .Y(new_n14310_));
  XOR2X1   g14054(.A(new_n14309_), .B(new_n14276_), .Y(new_n14311_));
  NAND2X1  g14055(.A(new_n14309_), .B(new_n14276_), .Y(new_n14312_));
  OAI21X1  g14056(.A0(new_n14310_), .A1(new_n14308_), .B0(new_n14312_), .Y(new_n14313_));
  OAI22X1  g14057(.A0(new_n14313_), .A1(new_n14310_), .B0(new_n14311_), .B1(new_n14308_), .Y(new_n14314_));
  AOI22X1  g14058(.A0(new_n7192_), .A1(\b[56] ), .B0(new_n7189_), .B1(\b[55] ), .Y(new_n14315_));
  OAI21X1  g14059(.A0(new_n7627_), .A1(new_n6148_), .B0(new_n14315_), .Y(new_n14316_));
  AOI21X1  g14060(.A0(new_n7187_), .A1(new_n6342_), .B0(new_n14316_), .Y(new_n14317_));
  XOR2X1   g14061(.A(new_n14317_), .B(\a[62] ), .Y(new_n14318_));
  XOR2X1   g14062(.A(new_n14318_), .B(new_n14314_), .Y(new_n14319_));
  AOI22X1  g14063(.A0(new_n6603_), .A1(\b[59] ), .B0(new_n6600_), .B1(\b[58] ), .Y(new_n14320_));
  OAI21X1  g14064(.A0(new_n6804_), .A1(new_n6933_), .B0(new_n14320_), .Y(new_n14321_));
  AOI21X1  g14065(.A0(new_n6932_), .A1(new_n6598_), .B0(new_n14321_), .Y(new_n14322_));
  XOR2X1   g14066(.A(new_n14322_), .B(\a[59] ), .Y(new_n14323_));
  XOR2X1   g14067(.A(new_n14323_), .B(new_n14319_), .Y(new_n14324_));
  XOR2X1   g14068(.A(new_n14324_), .B(new_n14305_), .Y(new_n14325_));
  AOI22X1  g14069(.A0(new_n6438_), .A1(\b[62] ), .B0(new_n6437_), .B1(\b[61] ), .Y(new_n14326_));
  OAI21X1  g14070(.A0(new_n6436_), .A1(new_n7559_), .B0(new_n14326_), .Y(new_n14327_));
  AOI21X1  g14071(.A0(new_n7558_), .A1(new_n6023_), .B0(new_n14327_), .Y(new_n14328_));
  XOR2X1   g14072(.A(new_n14328_), .B(\a[56] ), .Y(new_n14329_));
  XOR2X1   g14073(.A(new_n14329_), .B(new_n14325_), .Y(new_n14330_));
  OAI21X1  g14074(.A0(new_n14267_), .A1(new_n14266_), .B0(new_n14286_), .Y(new_n14331_));
  OR2X1    g14075(.A(new_n14287_), .B(new_n14264_), .Y(new_n14332_));
  AND2X1   g14076(.A(new_n14332_), .B(new_n14331_), .Y(new_n14333_));
  AOI22X1  g14077(.A0(new_n7774_), .A1(new_n5425_), .B0(new_n5890_), .B1(\b[63] ), .Y(new_n14334_));
  XOR2X1   g14078(.A(new_n14334_), .B(\a[53] ), .Y(new_n14335_));
  XOR2X1   g14079(.A(new_n14335_), .B(new_n14333_), .Y(new_n14336_));
  XOR2X1   g14080(.A(new_n14336_), .B(new_n14330_), .Y(new_n14337_));
  INVX1    g14081(.A(new_n14337_), .Y(new_n14338_));
  AND2X1   g14082(.A(new_n14288_), .B(new_n14260_), .Y(new_n14339_));
  INVX1    g14083(.A(new_n14292_), .Y(new_n14340_));
  AOI21X1  g14084(.A0(new_n14340_), .A1(new_n14289_), .B0(new_n14339_), .Y(new_n14341_));
  XOR2X1   g14085(.A(new_n14341_), .B(new_n14338_), .Y(new_n14342_));
  NOR2X1   g14086(.A(new_n14296_), .B(new_n14293_), .Y(new_n14343_));
  INVX1    g14087(.A(new_n14343_), .Y(new_n14344_));
  OAI21X1  g14088(.A0(new_n14300_), .A1(new_n14299_), .B0(new_n14297_), .Y(new_n14345_));
  AND2X1   g14089(.A(new_n14345_), .B(new_n14344_), .Y(new_n14346_));
  XOR2X1   g14090(.A(new_n14346_), .B(new_n14342_), .Y(\f[116] ));
  NOR2X1   g14091(.A(new_n14341_), .B(new_n14337_), .Y(new_n14348_));
  AOI21X1  g14092(.A0(new_n14345_), .A1(new_n14344_), .B0(new_n14342_), .Y(new_n14349_));
  OR2X1    g14093(.A(new_n14349_), .B(new_n14348_), .Y(new_n14350_));
  INVX1    g14094(.A(new_n14330_), .Y(new_n14351_));
  NOR2X1   g14095(.A(new_n14335_), .B(new_n14333_), .Y(new_n14352_));
  AOI21X1  g14096(.A0(new_n14336_), .A1(new_n14351_), .B0(new_n14352_), .Y(new_n14353_));
  AND2X1   g14097(.A(new_n14324_), .B(new_n14305_), .Y(new_n14354_));
  INVX1    g14098(.A(new_n14329_), .Y(new_n14355_));
  AOI21X1  g14099(.A0(new_n14355_), .A1(new_n14325_), .B0(new_n14354_), .Y(new_n14356_));
  AOI22X1  g14100(.A0(new_n6438_), .A1(\b[63] ), .B0(new_n6437_), .B1(\b[62] ), .Y(new_n14357_));
  OAI21X1  g14101(.A0(new_n6436_), .A1(new_n7748_), .B0(new_n14357_), .Y(new_n14358_));
  AOI21X1  g14102(.A0(new_n7747_), .A1(new_n6023_), .B0(new_n14358_), .Y(new_n14359_));
  XOR2X1   g14103(.A(new_n14359_), .B(\a[56] ), .Y(new_n14360_));
  XOR2X1   g14104(.A(new_n14360_), .B(new_n14356_), .Y(new_n14361_));
  INVX1    g14105(.A(new_n14318_), .Y(new_n14362_));
  NOR2X1   g14106(.A(new_n14323_), .B(new_n14319_), .Y(new_n14363_));
  AOI21X1  g14107(.A0(new_n14362_), .A1(new_n14314_), .B0(new_n14363_), .Y(new_n14364_));
  AOI22X1  g14108(.A0(new_n6603_), .A1(\b[60] ), .B0(new_n6600_), .B1(\b[59] ), .Y(new_n14365_));
  OAI21X1  g14109(.A0(new_n6804_), .A1(new_n6930_), .B0(new_n14365_), .Y(new_n14366_));
  AOI21X1  g14110(.A0(new_n6951_), .A1(new_n6598_), .B0(new_n14366_), .Y(new_n14367_));
  XOR2X1   g14111(.A(new_n14367_), .B(\a[59] ), .Y(new_n14368_));
  XOR2X1   g14112(.A(new_n14309_), .B(new_n5423_), .Y(new_n14369_));
  NAND3X1  g14113(.A(\b[53] ), .B(\a[63] ), .C(\a[62] ), .Y(new_n14370_));
  OAI21X1  g14114(.A0(new_n7624_), .A1(new_n6148_), .B0(new_n14370_), .Y(new_n14371_));
  XOR2X1   g14115(.A(new_n14371_), .B(new_n14369_), .Y(new_n14372_));
  AOI22X1  g14116(.A0(new_n7192_), .A1(\b[57] ), .B0(new_n7189_), .B1(\b[56] ), .Y(new_n14373_));
  OAI21X1  g14117(.A0(new_n7627_), .A1(new_n6523_), .B0(new_n14373_), .Y(new_n14374_));
  AOI21X1  g14118(.A0(new_n7187_), .A1(new_n6522_), .B0(new_n14374_), .Y(new_n14375_));
  XOR2X1   g14119(.A(new_n14375_), .B(\a[62] ), .Y(new_n14376_));
  XOR2X1   g14120(.A(new_n14376_), .B(new_n14372_), .Y(new_n14377_));
  XOR2X1   g14121(.A(new_n14377_), .B(new_n14313_), .Y(new_n14378_));
  XOR2X1   g14122(.A(new_n14378_), .B(new_n14368_), .Y(new_n14379_));
  XOR2X1   g14123(.A(new_n14379_), .B(new_n14364_), .Y(new_n14380_));
  INVX1    g14124(.A(new_n14380_), .Y(new_n14381_));
  XOR2X1   g14125(.A(new_n14381_), .B(new_n14361_), .Y(new_n14382_));
  XOR2X1   g14126(.A(new_n14382_), .B(new_n14353_), .Y(new_n14383_));
  XOR2X1   g14127(.A(new_n14383_), .B(new_n14350_), .Y(\f[117] ));
  AND2X1   g14128(.A(new_n14377_), .B(new_n14313_), .Y(new_n14385_));
  NOR2X1   g14129(.A(new_n14377_), .B(new_n14313_), .Y(new_n14386_));
  NOR3X1   g14130(.A(new_n14386_), .B(new_n14385_), .C(new_n14368_), .Y(new_n14387_));
  NOR2X1   g14131(.A(new_n14379_), .B(new_n14364_), .Y(new_n14388_));
  NOR2X1   g14132(.A(new_n14388_), .B(new_n14387_), .Y(new_n14389_));
  AOI22X1  g14133(.A0(new_n6603_), .A1(\b[61] ), .B0(new_n6600_), .B1(\b[60] ), .Y(new_n14390_));
  OAI21X1  g14134(.A0(new_n6804_), .A1(new_n7339_), .B0(new_n14390_), .Y(new_n14391_));
  AOI21X1  g14135(.A0(new_n7338_), .A1(new_n6598_), .B0(new_n14391_), .Y(new_n14392_));
  XOR2X1   g14136(.A(new_n14392_), .B(\a[59] ), .Y(new_n14393_));
  NOR2X1   g14137(.A(new_n14376_), .B(new_n14372_), .Y(new_n14394_));
  AOI21X1  g14138(.A0(new_n14377_), .A1(new_n14313_), .B0(new_n14394_), .Y(new_n14395_));
  AOI22X1  g14139(.A0(new_n7818_), .A1(\b[54] ), .B0(new_n7817_), .B1(\b[55] ), .Y(new_n14396_));
  INVX1    g14140(.A(new_n14396_), .Y(new_n14397_));
  INVX1    g14141(.A(new_n14369_), .Y(new_n14398_));
  NOR2X1   g14142(.A(new_n14309_), .B(\a[53] ), .Y(new_n14399_));
  AOI21X1  g14143(.A0(new_n14371_), .A1(new_n14398_), .B0(new_n14399_), .Y(new_n14400_));
  XOR2X1   g14144(.A(new_n14400_), .B(new_n14397_), .Y(new_n14401_));
  INVX1    g14145(.A(new_n14401_), .Y(new_n14402_));
  AOI22X1  g14146(.A0(new_n7192_), .A1(\b[58] ), .B0(new_n7189_), .B1(\b[57] ), .Y(new_n14403_));
  OAI21X1  g14147(.A0(new_n7627_), .A1(new_n6520_), .B0(new_n14403_), .Y(new_n14404_));
  AOI21X1  g14148(.A0(new_n7187_), .A1(new_n6732_), .B0(new_n14404_), .Y(new_n14405_));
  XOR2X1   g14149(.A(new_n14405_), .B(\a[62] ), .Y(new_n14406_));
  XOR2X1   g14150(.A(new_n14406_), .B(new_n14402_), .Y(new_n14407_));
  XOR2X1   g14151(.A(new_n14407_), .B(new_n14395_), .Y(new_n14408_));
  XOR2X1   g14152(.A(new_n14408_), .B(new_n14393_), .Y(new_n14409_));
  XOR2X1   g14153(.A(new_n14409_), .B(new_n14389_), .Y(new_n14410_));
  OAI22X1  g14154(.A0(new_n6436_), .A1(new_n7745_), .B0(new_n6025_), .B1(new_n7772_), .Y(new_n14411_));
  AOI21X1  g14155(.A0(new_n7775_), .A1(new_n6023_), .B0(new_n14411_), .Y(new_n14412_));
  XOR2X1   g14156(.A(new_n14412_), .B(\a[56] ), .Y(new_n14413_));
  XOR2X1   g14157(.A(new_n14413_), .B(new_n14410_), .Y(new_n14414_));
  NOR2X1   g14158(.A(new_n14360_), .B(new_n14356_), .Y(new_n14415_));
  AOI21X1  g14159(.A0(new_n14380_), .A1(new_n14361_), .B0(new_n14415_), .Y(new_n14416_));
  XOR2X1   g14160(.A(new_n14416_), .B(new_n14414_), .Y(new_n14417_));
  NOR2X1   g14161(.A(new_n14382_), .B(new_n14353_), .Y(new_n14418_));
  INVX1    g14162(.A(new_n14418_), .Y(new_n14419_));
  OAI21X1  g14163(.A0(new_n14349_), .A1(new_n14348_), .B0(new_n14383_), .Y(new_n14420_));
  AND2X1   g14164(.A(new_n14420_), .B(new_n14419_), .Y(new_n14421_));
  XOR2X1   g14165(.A(new_n14421_), .B(new_n14417_), .Y(\f[118] ));
  AOI22X1  g14166(.A0(new_n7192_), .A1(\b[59] ), .B0(new_n7189_), .B1(\b[58] ), .Y(new_n14423_));
  OAI21X1  g14167(.A0(new_n7627_), .A1(new_n6933_), .B0(new_n14423_), .Y(new_n14424_));
  AOI21X1  g14168(.A0(new_n7187_), .A1(new_n6932_), .B0(new_n14424_), .Y(new_n14425_));
  XOR2X1   g14169(.A(new_n14425_), .B(\a[62] ), .Y(new_n14426_));
  AOI22X1  g14170(.A0(new_n7818_), .A1(\b[55] ), .B0(new_n7817_), .B1(\b[56] ), .Y(new_n14427_));
  XOR2X1   g14171(.A(new_n14427_), .B(new_n14396_), .Y(new_n14428_));
  XOR2X1   g14172(.A(new_n14428_), .B(new_n14426_), .Y(new_n14429_));
  INVX1    g14173(.A(new_n14429_), .Y(new_n14430_));
  NOR2X1   g14174(.A(new_n14400_), .B(new_n14397_), .Y(new_n14431_));
  XOR2X1   g14175(.A(new_n14405_), .B(new_n7185_), .Y(new_n14432_));
  AOI21X1  g14176(.A0(new_n14432_), .A1(new_n14401_), .B0(new_n14431_), .Y(new_n14433_));
  XOR2X1   g14177(.A(new_n14433_), .B(new_n14430_), .Y(new_n14434_));
  AOI22X1  g14178(.A0(new_n6603_), .A1(\b[62] ), .B0(new_n6600_), .B1(\b[61] ), .Y(new_n14435_));
  OAI21X1  g14179(.A0(new_n6804_), .A1(new_n7559_), .B0(new_n14435_), .Y(new_n14436_));
  AOI21X1  g14180(.A0(new_n7558_), .A1(new_n6598_), .B0(new_n14436_), .Y(new_n14437_));
  XOR2X1   g14181(.A(new_n14437_), .B(\a[59] ), .Y(new_n14438_));
  XOR2X1   g14182(.A(new_n14438_), .B(new_n14434_), .Y(new_n14439_));
  OAI21X1  g14183(.A0(new_n14385_), .A1(new_n14394_), .B0(new_n14407_), .Y(new_n14440_));
  OR2X1    g14184(.A(new_n14408_), .B(new_n14393_), .Y(new_n14441_));
  AND2X1   g14185(.A(new_n14441_), .B(new_n14440_), .Y(new_n14442_));
  AOI22X1  g14186(.A0(new_n7774_), .A1(new_n6023_), .B0(new_n6214_), .B1(\b[63] ), .Y(new_n14443_));
  XOR2X1   g14187(.A(new_n14443_), .B(\a[56] ), .Y(new_n14444_));
  XOR2X1   g14188(.A(new_n14444_), .B(new_n14442_), .Y(new_n14445_));
  XOR2X1   g14189(.A(new_n14445_), .B(new_n14439_), .Y(new_n14446_));
  OAI21X1  g14190(.A0(new_n14388_), .A1(new_n14387_), .B0(new_n14409_), .Y(new_n14447_));
  OR2X1    g14191(.A(new_n14413_), .B(new_n14410_), .Y(new_n14448_));
  AND2X1   g14192(.A(new_n14448_), .B(new_n14447_), .Y(new_n14449_));
  XOR2X1   g14193(.A(new_n14449_), .B(new_n14446_), .Y(new_n14450_));
  INVX1    g14194(.A(new_n14414_), .Y(new_n14451_));
  NOR2X1   g14195(.A(new_n14416_), .B(new_n14451_), .Y(new_n14452_));
  AOI21X1  g14196(.A0(new_n14420_), .A1(new_n14419_), .B0(new_n14417_), .Y(new_n14453_));
  OR2X1    g14197(.A(new_n14453_), .B(new_n14452_), .Y(new_n14454_));
  XOR2X1   g14198(.A(new_n14454_), .B(new_n14450_), .Y(\f[119] ));
  NOR2X1   g14199(.A(new_n14433_), .B(new_n14430_), .Y(new_n14456_));
  INVX1    g14200(.A(new_n14456_), .Y(new_n14457_));
  INVX1    g14201(.A(new_n14434_), .Y(new_n14458_));
  OAI21X1  g14202(.A0(new_n14438_), .A1(new_n14458_), .B0(new_n14457_), .Y(new_n14459_));
  AOI22X1  g14203(.A0(new_n6603_), .A1(\b[63] ), .B0(new_n6600_), .B1(\b[62] ), .Y(new_n14460_));
  OAI21X1  g14204(.A0(new_n6804_), .A1(new_n7748_), .B0(new_n14460_), .Y(new_n14461_));
  AOI21X1  g14205(.A0(new_n7747_), .A1(new_n6598_), .B0(new_n14461_), .Y(new_n14462_));
  XOR2X1   g14206(.A(new_n14462_), .B(\a[59] ), .Y(new_n14463_));
  XOR2X1   g14207(.A(new_n14463_), .B(new_n14459_), .Y(new_n14464_));
  AOI22X1  g14208(.A0(new_n7818_), .A1(\b[56] ), .B0(new_n7817_), .B1(\b[57] ), .Y(new_n14465_));
  XOR2X1   g14209(.A(new_n14465_), .B(new_n6019_), .Y(new_n14466_));
  XOR2X1   g14210(.A(new_n14466_), .B(new_n14397_), .Y(new_n14467_));
  OR2X1    g14211(.A(new_n14427_), .B(new_n14397_), .Y(new_n14468_));
  OAI21X1  g14212(.A0(new_n14428_), .A1(new_n14426_), .B0(new_n14468_), .Y(new_n14469_));
  XOR2X1   g14213(.A(new_n14469_), .B(new_n14467_), .Y(new_n14470_));
  AOI22X1  g14214(.A0(new_n7192_), .A1(\b[60] ), .B0(new_n7189_), .B1(\b[59] ), .Y(new_n14471_));
  OAI21X1  g14215(.A0(new_n7627_), .A1(new_n6930_), .B0(new_n14471_), .Y(new_n14472_));
  AOI21X1  g14216(.A0(new_n7187_), .A1(new_n6951_), .B0(new_n14472_), .Y(new_n14473_));
  XOR2X1   g14217(.A(new_n14473_), .B(\a[62] ), .Y(new_n14474_));
  XOR2X1   g14218(.A(new_n14474_), .B(new_n14470_), .Y(new_n14475_));
  XOR2X1   g14219(.A(new_n14475_), .B(new_n14464_), .Y(new_n14476_));
  INVX1    g14220(.A(new_n14439_), .Y(new_n14477_));
  NOR2X1   g14221(.A(new_n14444_), .B(new_n14442_), .Y(new_n14478_));
  AOI21X1  g14222(.A0(new_n14445_), .A1(new_n14477_), .B0(new_n14478_), .Y(new_n14479_));
  XOR2X1   g14223(.A(new_n14479_), .B(new_n14476_), .Y(new_n14480_));
  INVX1    g14224(.A(new_n14480_), .Y(new_n14481_));
  AOI21X1  g14225(.A0(new_n14448_), .A1(new_n14447_), .B0(new_n14446_), .Y(new_n14482_));
  INVX1    g14226(.A(new_n14482_), .Y(new_n14483_));
  OAI21X1  g14227(.A0(new_n14453_), .A1(new_n14452_), .B0(new_n14450_), .Y(new_n14484_));
  AND2X1   g14228(.A(new_n14484_), .B(new_n14483_), .Y(new_n14485_));
  XOR2X1   g14229(.A(new_n14485_), .B(new_n14481_), .Y(\f[120] ));
  INVX1    g14230(.A(new_n14467_), .Y(new_n14487_));
  NOR2X1   g14231(.A(new_n14474_), .B(new_n14470_), .Y(new_n14488_));
  AOI21X1  g14232(.A0(new_n14469_), .A1(new_n14487_), .B0(new_n14488_), .Y(new_n14489_));
  AOI22X1  g14233(.A0(new_n7818_), .A1(\b[57] ), .B0(new_n7817_), .B1(\b[58] ), .Y(new_n14490_));
  OR2X1    g14234(.A(new_n14465_), .B(\a[56] ), .Y(new_n14491_));
  OAI21X1  g14235(.A0(new_n14466_), .A1(new_n14396_), .B0(new_n14491_), .Y(new_n14492_));
  XOR2X1   g14236(.A(new_n14492_), .B(new_n14490_), .Y(new_n14493_));
  AOI22X1  g14237(.A0(new_n7192_), .A1(\b[61] ), .B0(new_n7189_), .B1(\b[60] ), .Y(new_n14494_));
  OAI21X1  g14238(.A0(new_n7627_), .A1(new_n7339_), .B0(new_n14494_), .Y(new_n14495_));
  AOI21X1  g14239(.A0(new_n7338_), .A1(new_n7187_), .B0(new_n14495_), .Y(new_n14496_));
  XOR2X1   g14240(.A(new_n14496_), .B(\a[62] ), .Y(new_n14497_));
  INVX1    g14241(.A(new_n14497_), .Y(new_n14498_));
  XOR2X1   g14242(.A(new_n14498_), .B(new_n14493_), .Y(new_n14499_));
  INVX1    g14243(.A(new_n14499_), .Y(new_n14500_));
  XOR2X1   g14244(.A(new_n14500_), .B(new_n14489_), .Y(new_n14501_));
  OAI22X1  g14245(.A0(new_n6804_), .A1(new_n7745_), .B0(new_n6601_), .B1(new_n7772_), .Y(new_n14502_));
  AOI21X1  g14246(.A0(new_n7775_), .A1(new_n6598_), .B0(new_n14502_), .Y(new_n14503_));
  XOR2X1   g14247(.A(new_n14503_), .B(\a[59] ), .Y(new_n14504_));
  XOR2X1   g14248(.A(new_n14504_), .B(new_n14501_), .Y(new_n14505_));
  XOR2X1   g14249(.A(new_n14462_), .B(new_n6596_), .Y(new_n14506_));
  AND2X1   g14250(.A(new_n14506_), .B(new_n14459_), .Y(new_n14507_));
  INVX1    g14251(.A(new_n14464_), .Y(new_n14508_));
  AOI21X1  g14252(.A0(new_n14475_), .A1(new_n14508_), .B0(new_n14507_), .Y(new_n14509_));
  XOR2X1   g14253(.A(new_n14509_), .B(new_n14505_), .Y(new_n14510_));
  NOR2X1   g14254(.A(new_n14479_), .B(new_n14476_), .Y(new_n14511_));
  AOI21X1  g14255(.A0(new_n14484_), .A1(new_n14483_), .B0(new_n14481_), .Y(new_n14512_));
  OR2X1    g14256(.A(new_n14512_), .B(new_n14511_), .Y(new_n14513_));
  XOR2X1   g14257(.A(new_n14513_), .B(new_n14510_), .Y(\f[121] ));
  OR2X1    g14258(.A(new_n14509_), .B(new_n14505_), .Y(new_n14515_));
  OAI21X1  g14259(.A0(new_n14512_), .A1(new_n14511_), .B0(new_n14510_), .Y(new_n14516_));
  AND2X1   g14260(.A(new_n14516_), .B(new_n14515_), .Y(new_n14517_));
  NOR2X1   g14261(.A(new_n14500_), .B(new_n14489_), .Y(new_n14518_));
  INVX1    g14262(.A(new_n14518_), .Y(new_n14519_));
  INVX1    g14263(.A(new_n14501_), .Y(new_n14520_));
  OAI21X1  g14264(.A0(new_n14504_), .A1(new_n14520_), .B0(new_n14519_), .Y(new_n14521_));
  AND2X1   g14265(.A(new_n14492_), .B(new_n14490_), .Y(new_n14522_));
  AOI21X1  g14266(.A0(new_n14498_), .A1(new_n14493_), .B0(new_n14522_), .Y(new_n14523_));
  INVX1    g14267(.A(new_n14490_), .Y(new_n14524_));
  AOI22X1  g14268(.A0(new_n7818_), .A1(\b[58] ), .B0(new_n7817_), .B1(\b[59] ), .Y(new_n14525_));
  NOR2X1   g14269(.A(new_n14525_), .B(new_n14524_), .Y(new_n14526_));
  XOR2X1   g14270(.A(new_n14525_), .B(new_n14524_), .Y(new_n14527_));
  NAND2X1  g14271(.A(new_n14525_), .B(new_n14524_), .Y(new_n14528_));
  OAI21X1  g14272(.A0(new_n14526_), .A1(new_n14523_), .B0(new_n14528_), .Y(new_n14529_));
  OAI22X1  g14273(.A0(new_n14529_), .A1(new_n14526_), .B0(new_n14527_), .B1(new_n14523_), .Y(new_n14530_));
  AOI22X1  g14274(.A0(new_n7192_), .A1(\b[62] ), .B0(new_n7189_), .B1(\b[61] ), .Y(new_n14531_));
  OAI21X1  g14275(.A0(new_n7627_), .A1(new_n7559_), .B0(new_n14531_), .Y(new_n14532_));
  AOI21X1  g14276(.A0(new_n7558_), .A1(new_n7187_), .B0(new_n14532_), .Y(new_n14533_));
  XOR2X1   g14277(.A(new_n14533_), .B(new_n7185_), .Y(new_n14534_));
  AOI22X1  g14278(.A0(new_n7774_), .A1(new_n6598_), .B0(new_n6803_), .B1(\b[63] ), .Y(new_n14535_));
  XOR2X1   g14279(.A(new_n14535_), .B(\a[59] ), .Y(new_n14536_));
  XOR2X1   g14280(.A(new_n14536_), .B(new_n14534_), .Y(new_n14537_));
  XOR2X1   g14281(.A(new_n14537_), .B(new_n14530_), .Y(new_n14538_));
  XOR2X1   g14282(.A(new_n14538_), .B(new_n14521_), .Y(new_n14539_));
  XOR2X1   g14283(.A(new_n14539_), .B(new_n14517_), .Y(\f[122] ));
  INVX1    g14284(.A(new_n14537_), .Y(new_n14541_));
  XOR2X1   g14285(.A(new_n14541_), .B(new_n14530_), .Y(new_n14542_));
  AND2X1   g14286(.A(new_n14542_), .B(new_n14521_), .Y(new_n14543_));
  AOI21X1  g14287(.A0(new_n14516_), .A1(new_n14515_), .B0(new_n14539_), .Y(new_n14544_));
  NOR2X1   g14288(.A(new_n14544_), .B(new_n14543_), .Y(new_n14545_));
  XOR2X1   g14289(.A(new_n14533_), .B(\a[62] ), .Y(new_n14546_));
  NOR2X1   g14290(.A(new_n14536_), .B(new_n14546_), .Y(new_n14547_));
  AOI21X1  g14291(.A0(new_n14541_), .A1(new_n14530_), .B0(new_n14547_), .Y(new_n14548_));
  XOR2X1   g14292(.A(new_n14525_), .B(new_n6596_), .Y(new_n14549_));
  AOI22X1  g14293(.A0(new_n7818_), .A1(\b[59] ), .B0(new_n7817_), .B1(\b[60] ), .Y(new_n14550_));
  XOR2X1   g14294(.A(new_n14550_), .B(new_n14549_), .Y(new_n14551_));
  AOI22X1  g14295(.A0(new_n7192_), .A1(\b[63] ), .B0(new_n7189_), .B1(\b[62] ), .Y(new_n14552_));
  OAI21X1  g14296(.A0(new_n7627_), .A1(new_n7748_), .B0(new_n14552_), .Y(new_n14553_));
  AOI21X1  g14297(.A0(new_n7747_), .A1(new_n7187_), .B0(new_n14553_), .Y(new_n14554_));
  XOR2X1   g14298(.A(new_n14554_), .B(\a[62] ), .Y(new_n14555_));
  XOR2X1   g14299(.A(new_n14555_), .B(new_n14551_), .Y(new_n14556_));
  INVX1    g14300(.A(new_n14556_), .Y(new_n14557_));
  XOR2X1   g14301(.A(new_n14557_), .B(new_n14529_), .Y(new_n14558_));
  XOR2X1   g14302(.A(new_n14558_), .B(new_n14548_), .Y(new_n14559_));
  XOR2X1   g14303(.A(new_n14559_), .B(new_n14545_), .Y(\f[123] ));
  INVX1    g14304(.A(new_n14558_), .Y(new_n14561_));
  NOR2X1   g14305(.A(new_n14561_), .B(new_n14548_), .Y(new_n14562_));
  INVX1    g14306(.A(new_n14562_), .Y(new_n14563_));
  INVX1    g14307(.A(new_n14559_), .Y(new_n14564_));
  OAI21X1  g14308(.A0(new_n14544_), .A1(new_n14543_), .B0(new_n14564_), .Y(new_n14565_));
  AND2X1   g14309(.A(new_n14565_), .B(new_n14563_), .Y(new_n14566_));
  INVX1    g14310(.A(new_n14551_), .Y(new_n14567_));
  NOR2X1   g14311(.A(new_n14555_), .B(new_n14567_), .Y(new_n14568_));
  AOI21X1  g14312(.A0(new_n14557_), .A1(new_n14529_), .B0(new_n14568_), .Y(new_n14569_));
  AOI22X1  g14313(.A0(new_n7818_), .A1(\b[60] ), .B0(new_n7817_), .B1(\b[61] ), .Y(new_n14570_));
  INVX1    g14314(.A(new_n14570_), .Y(new_n14571_));
  OR2X1    g14315(.A(new_n14550_), .B(new_n14549_), .Y(new_n14572_));
  OR2X1    g14316(.A(new_n14525_), .B(\a[59] ), .Y(new_n14573_));
  AND2X1   g14317(.A(new_n14573_), .B(new_n14572_), .Y(new_n14574_));
  XOR2X1   g14318(.A(new_n14574_), .B(new_n14571_), .Y(new_n14575_));
  INVX1    g14319(.A(new_n14575_), .Y(new_n14576_));
  OAI22X1  g14320(.A0(new_n7627_), .A1(new_n7745_), .B0(new_n7190_), .B1(new_n7772_), .Y(new_n14577_));
  AOI21X1  g14321(.A0(new_n7775_), .A1(new_n7187_), .B0(new_n14577_), .Y(new_n14578_));
  XOR2X1   g14322(.A(new_n14578_), .B(\a[62] ), .Y(new_n14579_));
  XOR2X1   g14323(.A(new_n14579_), .B(new_n14576_), .Y(new_n14580_));
  XOR2X1   g14324(.A(new_n14580_), .B(new_n14569_), .Y(new_n14581_));
  XOR2X1   g14325(.A(new_n14581_), .B(new_n14566_), .Y(\f[124] ));
  INVX1    g14326(.A(new_n14580_), .Y(new_n14583_));
  NOR2X1   g14327(.A(new_n14583_), .B(new_n14569_), .Y(new_n14584_));
  AOI21X1  g14328(.A0(new_n14565_), .A1(new_n14563_), .B0(new_n14581_), .Y(new_n14585_));
  NOR2X1   g14329(.A(new_n14585_), .B(new_n14584_), .Y(new_n14586_));
  OR2X1    g14330(.A(new_n14574_), .B(new_n14571_), .Y(new_n14587_));
  OAI21X1  g14331(.A0(new_n14579_), .A1(new_n14576_), .B0(new_n14587_), .Y(new_n14588_));
  AOI22X1  g14332(.A0(new_n7818_), .A1(\b[61] ), .B0(new_n7817_), .B1(\b[62] ), .Y(new_n14589_));
  XOR2X1   g14333(.A(new_n14589_), .B(new_n14571_), .Y(new_n14590_));
  INVX1    g14334(.A(new_n14590_), .Y(new_n14591_));
  AOI22X1  g14335(.A0(new_n7774_), .A1(new_n7187_), .B0(new_n7411_), .B1(\b[63] ), .Y(new_n14592_));
  XOR2X1   g14336(.A(new_n14592_), .B(\a[62] ), .Y(new_n14593_));
  XOR2X1   g14337(.A(new_n14593_), .B(new_n14591_), .Y(new_n14594_));
  INVX1    g14338(.A(new_n14594_), .Y(new_n14595_));
  XOR2X1   g14339(.A(new_n14595_), .B(new_n14588_), .Y(new_n14596_));
  XOR2X1   g14340(.A(new_n14596_), .B(new_n14586_), .Y(\f[125] ));
  NAND2X1  g14341(.A(new_n14594_), .B(new_n14588_), .Y(new_n14598_));
  OAI21X1  g14342(.A0(new_n14596_), .A1(new_n14586_), .B0(new_n14598_), .Y(new_n14599_));
  OR2X1    g14343(.A(new_n14589_), .B(new_n14571_), .Y(new_n14600_));
  OAI21X1  g14344(.A0(new_n14593_), .A1(new_n14591_), .B0(new_n14600_), .Y(new_n14601_));
  AOI22X1  g14345(.A0(new_n7818_), .A1(\b[62] ), .B0(new_n7817_), .B1(\b[63] ), .Y(new_n14602_));
  XOR2X1   g14346(.A(new_n14602_), .B(\a[62] ), .Y(new_n14603_));
  XOR2X1   g14347(.A(new_n14603_), .B(new_n14571_), .Y(new_n14604_));
  XOR2X1   g14348(.A(new_n14604_), .B(new_n14601_), .Y(new_n14605_));
  XOR2X1   g14349(.A(new_n14605_), .B(new_n14599_), .Y(\f[126] ));
  NOR2X1   g14350(.A(new_n14602_), .B(\a[62] ), .Y(new_n14607_));
  AOI21X1  g14351(.A0(new_n14603_), .A1(new_n14571_), .B0(new_n14607_), .Y(new_n14608_));
  NAND3X1  g14352(.A(\b[63] ), .B(\a[63] ), .C(\a[62] ), .Y(new_n14609_));
  XOR2X1   g14353(.A(new_n14609_), .B(new_n14608_), .Y(new_n14610_));
  AND2X1   g14354(.A(new_n14604_), .B(new_n14601_), .Y(new_n14611_));
  AOI21X1  g14355(.A0(new_n14605_), .A1(new_n14599_), .B0(new_n14611_), .Y(new_n14612_));
  XOR2X1   g14356(.A(new_n14612_), .B(new_n14610_), .Y(\f[127] ));
endmodule


