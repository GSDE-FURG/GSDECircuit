//Converted to Combinational , Module name: s832 , Timestamp: 2018-12-03T15:51:02.061896 
module s832 ( G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G18, G38, G39, G40, G41, G42, G327, G325, G300, G322, G45, G312, G53, G49, G47, G296, G290, G292, G298, G288, G315, G55, G43, G310, G302, n75, n80, n85, n90, n95 );
input G0, G1, G2, G3, G4, G5, G6, G7, G8, G9, G10, G11, G12, G13, G14, G15, G16, G18, G38, G39, G40, G41, G42;
output G327, G325, G300, G322, G45, G312, G53, G49, G47, G296, G290, G292, G298, G288, G315, G55, G43, G310, G302, n75, n80, n85, n90, n95;
wire n52, n53, n54, n55, n57, n58, n60, n61, n62, n63, n64, n66, n67, n68, n70, n71, n72, n73, n74, n76, n77, n78, n80_1, n81, n83, n84, n85_1, n86, n87, n88, n89, n92, n95_1, n96, n97, n101, n102, n103, n104, n107, n109, n111, n113, n114, n115, n116, n117, n118, n119, n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249;
INVX1    g000(.A(G15), .Y(n52));
INVX1    g001(.A(G39), .Y(n53));
INVX1    g002(.A(G42), .Y(n54));
OR2X1    g003(.A(G41), .B(G40), .Y(n55));
NOR4X1   g004(.A(n54), .B(n53), .C(n52), .D(n55), .Y(G327));
AND2X1   g005(.A(G40), .B(G39), .Y(n57));
INVX1    g006(.A(n57), .Y(n58));
NOR4X1   g007(.A(n54), .B(G41), .C(G38), .D(n58), .Y(G325));
OR2X1    g008(.A(G42), .B(G41), .Y(n60));
INVX1    g009(.A(G1), .Y(n61));
INVX1    g010(.A(G16), .Y(n62));
NOR2X1   g011(.A(G39), .B(G38), .Y(n63));
NAND4X1  g012(.A(n62), .B(G3), .C(n61), .D(n63), .Y(n64));
NOR3X1   g013(.A(n64), .B(n60), .C(G40), .Y(G300));
NOR2X1   g014(.A(G40), .B(G39), .Y(n66));
INVX1    g015(.A(n66), .Y(n67));
MX2X1    g016(.A(n58), .B(n67), .S0(n54), .Y(n68));
NOR4X1   g017(.A(G41), .B(G38), .C(n61), .D(n68), .Y(G322));
OAI21X1  g018(.A0(G12), .A1(G10), .B0(n63), .Y(n70));
AOI21X1  g019(.A0(G12), .A1(G10), .B0(G11), .Y(n71));
NAND3X1  g020(.A(n54), .B(G41), .C(G40), .Y(n72));
INVX1    g021(.A(G4), .Y(n73));
NAND3X1  g022(.A(G16), .B(G15), .C(n73), .Y(n74));
NOR4X1   g023(.A(n72), .B(n71), .C(n70), .D(n74), .Y(G45));
INVX1    g024(.A(G38), .Y(n76));
NAND2X1  g025(.A(n57), .B(n76), .Y(n77));
NAND2X1  g026(.A(G42), .B(G41), .Y(n78));
NOR3X1   g027(.A(n78), .B(n77), .C(n62), .Y(G312));
INVX1    g028(.A(G41), .Y(n80_1));
OR2X1    g029(.A(G42), .B(G38), .Y(n81));
NOR4X1   g030(.A(n80_1), .B(G40), .C(G39), .D(n81), .Y(G53));
NOR2X1   g031(.A(G40), .B(n76), .Y(n83));
AND2X1   g032(.A(G42), .B(G41), .Y(n84));
NAND2X1  g033(.A(n84), .B(n53), .Y(n85_1));
NAND2X1  g034(.A(G39), .B(G38), .Y(n86));
NOR2X1   g035(.A(n86), .B(n60), .Y(n87));
MX2X1    g036(.A(G39), .B(n63), .S0(G40), .Y(n88));
NOR2X1   g037(.A(n88), .B(n87), .Y(n89));
OAI21X1  g038(.A0(n85_1), .A1(n83), .B0(n89), .Y(G49));
NOR3X1   g039(.A(n77), .B(n60), .C(G5), .Y(G47));
NAND2X1  g040(.A(G41), .B(G40), .Y(n92));
NOR3X1   g041(.A(n92), .B(n81), .C(n53), .Y(G296));
NOR4X1   g042(.A(G42), .B(n53), .C(n52), .D(n55), .Y(G290));
NAND2X1  g043(.A(G38), .B(G15), .Y(n95_1));
NAND4X1  g044(.A(G8), .B(G7), .C(G6), .D(G9), .Y(n96));
OAI21X1  g045(.A0(n96), .A1(n95_1), .B0(G16), .Y(n97));
AND2X1   g046(.A(n169), .B(n97), .Y(G292));
NOR3X1   g047(.A(G42), .B(n80_1), .C(G40), .Y(n101));
INVX1    g048(.A(G14), .Y(n102));
OR2X1    g049(.A(G39), .B(G38), .Y(n103));
NOR3X1   g050(.A(n103), .B(n52), .C(n102), .Y(n104));
AND2X1   g051(.A(n104), .B(n101), .Y(G298));
NOR4X1   g052(.A(G42), .B(G41), .C(G38), .D(n58), .Y(G288));
NAND4X1  g053(.A(n54), .B(n80_1), .C(n76), .D(n66), .Y(n107));
OAI21X1  g054(.A0(n78), .A1(n77), .B0(n107), .Y(G315));
INVX1    g055(.A(G5), .Y(n109));
NOR3X1   g056(.A(n77), .B(n60), .C(n109), .Y(G55));
NAND3X1  g057(.A(n54), .B(G41), .C(G15), .Y(n111));
NOR3X1   g058(.A(n111), .B(n67), .C(G38), .Y(G43));
NOR4X1   g059(.A(G40), .B(n62), .C(G1), .D(n60), .Y(n113));
INVX1    g060(.A(G40), .Y(n114));
AOI21X1  g061(.A0(G16), .A1(n73), .B0(n114), .Y(n115));
OAI21X1  g062(.A0(n115), .A1(n113), .B0(n63), .Y(n116));
OAI21X1  g063(.A0(n60), .A1(n76), .B0(G40), .Y(n117));
NAND3X1  g064(.A(n117), .B(G39), .C(G4), .Y(n118));
OAI22X1  g065(.A0(n76), .A1(G40), .B0(n62), .B1(G4), .Y(n119));
OR2X1    g066(.A(n119), .B(n85_1), .Y(n120));
NAND4X1  g067(.A(n114), .B(G39), .C(n62), .D(n78), .Y(n121));
NAND4X1  g068(.A(n120), .B(n118), .C(n116), .D(n121), .Y(G302));
NAND4X1  g069(.A(G39), .B(n76), .C(G1), .D(n80_1), .Y(n123));
INVX1    g070(.A(G0), .Y(n124));
NAND3X1  g071(.A(G39), .B(G38), .C(n124), .Y(n125));
AND2X1   g072(.A(G42), .B(G40), .Y(n126));
OAI21X1  g073(.A0(G41), .A1(n76), .B0(n126), .Y(n127));
AOI21X1  g074(.A0(n125), .A1(n123), .B0(n127), .Y(n128));
NAND2X1  g075(.A(G16), .B(n73), .Y(n129));
AOI21X1  g076(.A0(G41), .A1(G40), .B0(G39), .Y(n130));
AND2X1   g077(.A(G41), .B(G40), .Y(n131));
MX2X1    g078(.A(n57), .B(n131), .S0(n54), .Y(n132));
NOR4X1   g079(.A(n130), .B(n129), .C(n76), .D(n132), .Y(n133));
OAI21X1  g080(.A0(n54), .A1(G16), .B0(n53), .Y(n134));
NOR2X1   g081(.A(G41), .B(G40), .Y(n135));
OAI21X1  g082(.A0(n54), .A1(G38), .B0(n135), .Y(n136));
NOR3X1   g083(.A(G42), .B(n76), .C(n124), .Y(n137));
NOR3X1   g084(.A(G38), .B(G16), .C(G1), .Y(n138));
NOR4X1   g085(.A(n137), .B(n136), .C(n134), .D(n138), .Y(n139));
OR2X1    g086(.A(G11), .B(G10), .Y(n140));
OR2X1    g087(.A(G12), .B(G11), .Y(n141));
NAND3X1  g088(.A(n141), .B(n140), .C(n63), .Y(n142));
NOR4X1   g089(.A(n129), .B(n72), .C(n52), .D(n142), .Y(n143));
NOR4X1   g090(.A(n139), .B(n133), .C(n128), .D(n143), .Y(n144));
NOR2X1   g091(.A(n144), .B(G18), .Y(n75));
NOR2X1   g092(.A(n60), .B(n109), .Y(n146));
INVX1    g093(.A(G3), .Y(n147));
OAI21X1  g094(.A0(n54), .A1(n147), .B0(n76), .Y(n148));
AOI21X1  g095(.A0(n80_1), .A1(n61), .B0(n54), .Y(n149));
NOR3X1   g096(.A(n149), .B(n148), .C(n146), .Y(n150));
NAND3X1  g097(.A(n84), .B(G38), .C(n124), .Y(n151));
NAND3X1  g098(.A(n80_1), .B(G38), .C(n73), .Y(n152));
AOI22X1  g099(.A0(n151), .A1(n152), .B0(G42), .B1(n80_1), .Y(n153));
OAI21X1  g100(.A0(n153), .A1(n150), .B0(n57), .Y(n154));
NAND4X1  g101(.A(G16), .B(G15), .C(n73), .D(n53), .Y(n155));
OAI21X1  g102(.A0(G42), .A1(n76), .B0(n131), .Y(n156));
INVX1    g103(.A(G10), .Y(n157));
NOR4X1   g104(.A(G12), .B(G11), .C(n157), .D(G42), .Y(n158));
NAND2X1  g105(.A(n54), .B(G11), .Y(n159));
NOR3X1   g106(.A(n159), .B(G12), .C(G10), .Y(n160));
NOR4X1   g107(.A(n158), .B(n156), .C(n155), .D(n160), .Y(n161));
NAND4X1  g108(.A(n147), .B(G2), .C(n61), .D(n62), .Y(n162));
NOR4X1   g109(.A(n103), .B(n60), .C(G40), .D(n162), .Y(n163));
AOI21X1  g110(.A0(G42), .A1(G41), .B0(G16), .Y(n164));
NOR4X1   g111(.A(G40), .B(n53), .C(G4), .D(n164), .Y(n165));
NOR3X1   g112(.A(n165), .B(n163), .C(n161), .Y(n166));
AOI21X1  g113(.A0(n166), .A1(n154), .B0(G18), .Y(n80));
INVX1    g114(.A(G18), .Y(n168));
NOR4X1   g115(.A(G40), .B(n53), .C(G4), .D(n78), .Y(n169));
NAND2X1  g116(.A(n169), .B(n97), .Y(n170));
NAND2X1  g117(.A(n162), .B(n80_1), .Y(n171));
NAND2X1  g118(.A(G15), .B(n102), .Y(n172));
AOI21X1  g119(.A0(n172), .A1(G41), .B0(n103), .Y(n173));
NOR2X1   g120(.A(G42), .B(G40), .Y(n174));
NAND3X1  g121(.A(n174), .B(n173), .C(n171), .Y(n175));
AOI21X1  g122(.A0(n54), .A1(G10), .B0(n92), .Y(n176));
NAND3X1  g123(.A(n176), .B(n159), .C(G15), .Y(n177));
NAND3X1  g124(.A(n84), .B(n76), .C(G15), .Y(n178));
NAND2X1  g125(.A(n178), .B(n114), .Y(n179));
NAND3X1  g126(.A(n53), .B(G16), .C(n73), .Y(n180));
AOI21X1  g127(.A0(n78), .A1(G38), .B0(n180), .Y(n181));
NAND3X1  g128(.A(n181), .B(n179), .C(n177), .Y(n182));
NAND4X1  g129(.A(n175), .B(n170), .C(n154), .D(n182), .Y(n183));
AND2X1   g130(.A(n183), .B(n168), .Y(n85));
NOR4X1   g131(.A(G41), .B(n114), .C(n52), .D(n54), .Y(n185));
NOR3X1   g132(.A(n185), .B(n174), .C(n62), .Y(n186));
NOR3X1   g133(.A(G42), .B(G41), .C(G40), .Y(n187));
OAI21X1  g134(.A0(n114), .A1(n73), .B0(n53), .Y(n188));
OR2X1    g135(.A(G42), .B(G40), .Y(n189));
OAI22X1  g136(.A0(n172), .A1(n189), .B0(n78), .B1(n73), .Y(n190));
NOR4X1   g137(.A(n188), .B(n187), .C(n186), .D(n190), .Y(n191));
NOR3X1   g138(.A(G42), .B(n80_1), .C(G4), .Y(n192));
NOR2X1   g139(.A(n192), .B(G39), .Y(n193));
AOI21X1  g140(.A0(n80_1), .A1(n109), .B0(n114), .Y(n194));
OAI21X1  g141(.A0(n80_1), .A1(G16), .B0(G42), .Y(n195));
NAND2X1  g142(.A(n195), .B(n194), .Y(n196));
AOI22X1  g143(.A0(n57), .A1(G42), .B0(n62), .B1(n66), .Y(n197));
NAND4X1  g144(.A(n147), .B(G2), .C(n61), .D(n80_1), .Y(n198));
OAI22X1  g145(.A0(n197), .A1(n198), .B0(n196), .B1(n193), .Y(n199));
OAI21X1  g146(.A0(n199), .A1(n191), .B0(n76), .Y(n200));
AOI21X1  g147(.A0(G38), .A1(G15), .B0(n80_1), .Y(n201));
NOR2X1   g148(.A(n201), .B(n96), .Y(n202));
NOR2X1   g149(.A(G40), .B(n62), .Y(n203));
OAI21X1  g150(.A0(G39), .A1(n76), .B0(n203), .Y(n204));
AOI21X1  g151(.A0(G42), .A1(G15), .B0(G41), .Y(n205));
AOI21X1  g152(.A0(n53), .A1(G15), .B0(G4), .Y(n206));
OAI21X1  g153(.A0(n95_1), .A1(G42), .B0(n206), .Y(n207));
NOR4X1   g154(.A(n205), .B(n204), .C(n202), .D(n207), .Y(n208));
NAND3X1  g155(.A(G42), .B(G41), .C(G40), .Y(n209));
NAND3X1  g156(.A(G16), .B(G15), .C(G13), .Y(n210));
NAND3X1  g157(.A(n210), .B(n53), .C(n73), .Y(n211));
NOR2X1   g158(.A(n211), .B(n209), .Y(n212));
NOR3X1   g159(.A(n209), .B(n86), .C(G0), .Y(n213));
NAND4X1  g160(.A(n114), .B(G39), .C(n73), .D(n78), .Y(n214));
NOR2X1   g161(.A(n60), .B(n62), .Y(n215));
NOR3X1   g162(.A(G41), .B(n62), .C(G15), .Y(n216));
NOR3X1   g163(.A(n216), .B(n215), .C(n214), .Y(n217));
NOR4X1   g164(.A(n213), .B(n212), .C(n208), .D(n217), .Y(n218));
AOI21X1  g165(.A0(n218), .A1(n200), .B0(G18), .Y(n90));
NAND2X1  g166(.A(n54), .B(G38), .Y(n220));
NAND3X1  g167(.A(G42), .B(G15), .C(G13), .Y(n221));
OR2X1    g168(.A(G42), .B(G15), .Y(n222));
NAND4X1  g169(.A(n221), .B(n220), .C(G40), .D(n222), .Y(n223));
AOI21X1  g170(.A0(n96), .A1(n114), .B0(n86), .Y(n224));
OAI21X1  g171(.A0(G40), .A1(G15), .B0(G41), .Y(n225));
OR2X1    g172(.A(n225), .B(n224), .Y(n226));
AOI21X1  g173(.A0(n223), .A1(n53), .B0(n226), .Y(n227));
NAND3X1  g174(.A(G42), .B(G39), .C(G15), .Y(n228));
OAI21X1  g175(.A0(n54), .A1(G41), .B0(n53), .Y(n229));
NAND4X1  g176(.A(n228), .B(n222), .C(n114), .D(n229), .Y(n230));
NOR3X1   g177(.A(G42), .B(n114), .C(n52), .Y(n231));
INVX1    g178(.A(G6), .Y(n232));
INVX1    g179(.A(G9), .Y(n233));
NOR4X1   g180(.A(G8), .B(G7), .C(n232), .D(n233), .Y(n234));
OAI22X1  g181(.A0(n54), .A1(G15), .B0(G1), .B1(n55), .Y(n235));
AOI21X1  g182(.A0(n234), .A1(n231), .B0(n235), .Y(n236));
OAI21X1  g183(.A0(n236), .A1(n103), .B0(n230), .Y(n237));
OAI21X1  g184(.A0(n237), .A1(n227), .B0(G16), .Y(n238));
OR2X1    g185(.A(G3), .B(G1), .Y(n239));
NOR4X1   g186(.A(n54), .B(G41), .C(G2), .D(n239), .Y(n240));
AOI21X1  g187(.A0(n80_1), .A1(G5), .B0(G42), .Y(n241));
OAI21X1  g188(.A0(n241), .A1(n240), .B0(n57), .Y(n242));
NAND4X1  g189(.A(n53), .B(G15), .C(G14), .D(n101), .Y(n243));
NAND4X1  g190(.A(n55), .B(n53), .C(G4), .D(n189), .Y(n244));
NAND3X1  g191(.A(n244), .B(n243), .C(n242), .Y(n245));
OAI21X1  g192(.A0(n76), .A1(G0), .B0(G39), .Y(n246));
OAI21X1  g193(.A0(G39), .A1(G4), .B0(n246), .Y(n247));
OAI21X1  g194(.A0(n247), .A1(n209), .B0(n118), .Y(n248));
AOI21X1  g195(.A0(n245), .A1(n76), .B0(n248), .Y(n249));
AOI21X1  g196(.A0(n249), .A1(n238), .B0(G18), .Y(n95));
NOR4X1   g197(.A(n54), .B(G41), .C(G38), .D(n58), .Y(G310));
endmodule
