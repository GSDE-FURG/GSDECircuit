// Benchmark "mem_ctrl" written by ABC on Fri Sep 18 14:36:54 2020

module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire new_n2436_, new_n2437_, new_n2438_, new_n2439_, new_n2440_,
    new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_, new_n2446_,
    new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_, new_n2452_,
    new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_, new_n2458_,
    new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_, new_n2464_,
    new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_, new_n2470_,
    new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_, new_n2476_,
    new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_, new_n2482_,
    new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_, new_n2488_,
    new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_, new_n2494_,
    new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_, new_n2500_,
    new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_, new_n2506_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2584_,
    new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_,
    new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_,
    new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_,
    new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_,
    new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_,
    new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_,
    new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_,
    new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_,
    new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_,
    new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_,
    new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_, new_n2650_,
    new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_, new_n2656_,
    new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_, new_n2662_,
    new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_, new_n2668_,
    new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_, new_n2674_,
    new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_, new_n2680_,
    new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_, new_n2686_,
    new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_, new_n2692_,
    new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_, new_n2698_,
    new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_, new_n2704_,
    new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_, new_n2710_,
    new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_, new_n2716_,
    new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_, new_n2722_,
    new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_, new_n2728_,
    new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_, new_n2734_,
    new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_, new_n2740_,
    new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_, new_n2746_,
    new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_, new_n2752_,
    new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_, new_n2758_,
    new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_, new_n2764_,
    new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_, new_n2770_,
    new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_, new_n2776_,
    new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_, new_n2782_,
    new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_, new_n2788_,
    new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_, new_n2794_,
    new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_, new_n2800_,
    new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_, new_n2806_,
    new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_, new_n2812_,
    new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_, new_n2818_,
    new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_, new_n2824_,
    new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_, new_n2830_,
    new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_, new_n2836_,
    new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_, new_n2842_,
    new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_, new_n2848_,
    new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_, new_n2854_,
    new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_, new_n2860_,
    new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_, new_n2866_,
    new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_, new_n2872_,
    new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_, new_n2878_,
    new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_, new_n2884_,
    new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_, new_n2890_,
    new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_, new_n2896_,
    new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_, new_n2902_,
    new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2974_,
    new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_,
    new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_,
    new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_,
    new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_,
    new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_,
    new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_,
    new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_,
    new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_,
    new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_,
    new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_, new_n3034_,
    new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_, new_n3040_,
    new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_, new_n3046_,
    new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_, new_n3052_,
    new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_, new_n3058_,
    new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_, new_n3064_,
    new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_, new_n3070_,
    new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_, new_n3076_,
    new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_, new_n3082_,
    new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_, new_n3088_,
    new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_, new_n3094_,
    new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_, new_n3100_,
    new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_, new_n3106_,
    new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_, new_n3112_,
    new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_, new_n3118_,
    new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_, new_n3124_,
    new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3130_, new_n3131_,
    new_n3132_, new_n3133_, new_n3134_, new_n3135_, new_n3136_, new_n3137_,
    new_n3138_, new_n3139_, new_n3140_, new_n3141_, new_n3142_, new_n3143_,
    new_n3144_, new_n3145_, new_n3146_, new_n3147_, new_n3148_, new_n3149_,
    new_n3150_, new_n3151_, new_n3152_, new_n3153_, new_n3154_, new_n3155_,
    new_n3156_, new_n3157_, new_n3158_, new_n3159_, new_n3160_, new_n3161_,
    new_n3162_, new_n3163_, new_n3164_, new_n3165_, new_n3166_, new_n3167_,
    new_n3168_, new_n3169_, new_n3170_, new_n3171_, new_n3172_, new_n3173_,
    new_n3174_, new_n3175_, new_n3176_, new_n3177_, new_n3178_, new_n3179_,
    new_n3180_, new_n3181_, new_n3182_, new_n3183_, new_n3184_, new_n3185_,
    new_n3186_, new_n3187_, new_n3188_, new_n3189_, new_n3190_, new_n3191_,
    new_n3192_, new_n3193_, new_n3194_, new_n3195_, new_n3196_, new_n3197_,
    new_n3198_, new_n3199_, new_n3200_, new_n3201_, new_n3202_, new_n3203_,
    new_n3204_, new_n3205_, new_n3206_, new_n3207_, new_n3208_, new_n3209_,
    new_n3210_, new_n3211_, new_n3212_, new_n3213_, new_n3214_, new_n3215_,
    new_n3216_, new_n3217_, new_n3218_, new_n3219_, new_n3220_, new_n3221_,
    new_n3222_, new_n3223_, new_n3224_, new_n3225_, new_n3226_, new_n3227_,
    new_n3228_, new_n3229_, new_n3230_, new_n3231_, new_n3232_, new_n3233_,
    new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_, new_n3239_,
    new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_, new_n3245_,
    new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_, new_n3251_,
    new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_, new_n3257_,
    new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_, new_n3263_,
    new_n3264_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3298_, new_n3299_, new_n3300_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3348_,
    new_n3349_, new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_,
    new_n3355_, new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3360_,
    new_n3361_, new_n3362_, new_n3363_, new_n3364_, new_n3365_, new_n3366_,
    new_n3367_, new_n3368_, new_n3369_, new_n3370_, new_n3371_, new_n3372_,
    new_n3373_, new_n3374_, new_n3375_, new_n3376_, new_n3377_, new_n3378_,
    new_n3379_, new_n3380_, new_n3381_, new_n3382_, new_n3383_, new_n3384_,
    new_n3385_, new_n3386_, new_n3387_, new_n3388_, new_n3389_, new_n3390_,
    new_n3391_, new_n3392_, new_n3393_, new_n3394_, new_n3395_, new_n3396_,
    new_n3397_, new_n3398_, new_n3399_, new_n3400_, new_n3401_, new_n3402_,
    new_n3403_, new_n3404_, new_n3405_, new_n3406_, new_n3407_, new_n3408_,
    new_n3409_, new_n3410_, new_n3411_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3417_, new_n3418_, new_n3419_, new_n3420_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3427_,
    new_n3428_, new_n3429_, new_n3430_, new_n3431_, new_n3432_, new_n3433_,
    new_n3434_, new_n3435_, new_n3436_, new_n3437_, new_n3438_, new_n3439_,
    new_n3440_, new_n3441_, new_n3442_, new_n3443_, new_n3444_, new_n3445_,
    new_n3446_, new_n3447_, new_n3448_, new_n3449_, new_n3450_, new_n3451_,
    new_n3452_, new_n3453_, new_n3454_, new_n3455_, new_n3456_, new_n3457_,
    new_n3458_, new_n3459_, new_n3460_, new_n3461_, new_n3462_, new_n3463_,
    new_n3464_, new_n3465_, new_n3466_, new_n3467_, new_n3468_, new_n3469_,
    new_n3470_, new_n3471_, new_n3472_, new_n3473_, new_n3474_, new_n3475_,
    new_n3476_, new_n3477_, new_n3478_, new_n3479_, new_n3480_, new_n3481_,
    new_n3482_, new_n3483_, new_n3484_, new_n3485_, new_n3486_, new_n3487_,
    new_n3488_, new_n3489_, new_n3490_, new_n3491_, new_n3492_, new_n3493_,
    new_n3494_, new_n3495_, new_n3496_, new_n3497_, new_n3498_, new_n3499_,
    new_n3500_, new_n3501_, new_n3502_, new_n3503_, new_n3504_, new_n3505_,
    new_n3506_, new_n3507_, new_n3508_, new_n3509_, new_n3510_, new_n3511_,
    new_n3512_, new_n3513_, new_n3514_, new_n3515_, new_n3516_, new_n3517_,
    new_n3518_, new_n3519_, new_n3520_, new_n3521_, new_n3522_, new_n3523_,
    new_n3524_, new_n3525_, new_n3526_, new_n3527_, new_n3528_, new_n3529_,
    new_n3530_, new_n3531_, new_n3532_, new_n3533_, new_n3534_, new_n3535_,
    new_n3536_, new_n3537_, new_n3538_, new_n3539_, new_n3540_, new_n3541_,
    new_n3542_, new_n3543_, new_n3544_, new_n3545_, new_n3546_, new_n3547_,
    new_n3548_, new_n3549_, new_n3550_, new_n3551_, new_n3552_, new_n3553_,
    new_n3554_, new_n3555_, new_n3556_, new_n3557_, new_n3559_, new_n3560_,
    new_n3561_, new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_,
    new_n3567_, new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_,
    new_n3573_, new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_,
    new_n3579_, new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_,
    new_n3585_, new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_,
    new_n3591_, new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_,
    new_n3597_, new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_,
    new_n3603_, new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_,
    new_n3609_, new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_,
    new_n3615_, new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_,
    new_n3621_, new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_,
    new_n3627_, new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_,
    new_n3633_, new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_,
    new_n3639_, new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_,
    new_n3645_, new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_,
    new_n3651_, new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_,
    new_n3657_, new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_,
    new_n3663_, new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_,
    new_n3669_, new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_,
    new_n3675_, new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_,
    new_n3681_, new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_,
    new_n3687_, new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_,
    new_n3693_, new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_,
    new_n3699_, new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_,
    new_n3705_, new_n3706_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3858_, new_n3859_, new_n3860_, new_n3861_, new_n3862_,
    new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_, new_n3868_,
    new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_, new_n3874_,
    new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_, new_n3880_,
    new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_, new_n3886_,
    new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_, new_n3892_,
    new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_, new_n3898_,
    new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_, new_n3904_,
    new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_, new_n3910_,
    new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_, new_n3916_,
    new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_, new_n3922_,
    new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_, new_n3928_,
    new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_, new_n3934_,
    new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_, new_n3940_,
    new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_, new_n3946_,
    new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_, new_n3952_,
    new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_, new_n3958_,
    new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_, new_n3964_,
    new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_, new_n3970_,
    new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_, new_n3976_,
    new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_, new_n3982_,
    new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_, new_n3988_,
    new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_, new_n3994_,
    new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_, new_n4000_,
    new_n4001_, new_n4002_, new_n4004_, new_n4005_, new_n4006_, new_n4007_,
    new_n4008_, new_n4009_, new_n4010_, new_n4011_, new_n4012_, new_n4013_,
    new_n4014_, new_n4015_, new_n4016_, new_n4017_, new_n4018_, new_n4019_,
    new_n4020_, new_n4021_, new_n4022_, new_n4023_, new_n4024_, new_n4025_,
    new_n4026_, new_n4027_, new_n4028_, new_n4029_, new_n4030_, new_n4031_,
    new_n4032_, new_n4033_, new_n4034_, new_n4035_, new_n4036_, new_n4037_,
    new_n4038_, new_n4039_, new_n4040_, new_n4041_, new_n4042_, new_n4043_,
    new_n4044_, new_n4045_, new_n4046_, new_n4047_, new_n4048_, new_n4049_,
    new_n4050_, new_n4051_, new_n4052_, new_n4053_, new_n4054_, new_n4055_,
    new_n4056_, new_n4057_, new_n4058_, new_n4059_, new_n4060_, new_n4061_,
    new_n4062_, new_n4063_, new_n4064_, new_n4065_, new_n4066_, new_n4067_,
    new_n4068_, new_n4069_, new_n4070_, new_n4071_, new_n4072_, new_n4073_,
    new_n4074_, new_n4075_, new_n4076_, new_n4077_, new_n4078_, new_n4079_,
    new_n4080_, new_n4081_, new_n4082_, new_n4083_, new_n4084_, new_n4085_,
    new_n4086_, new_n4087_, new_n4088_, new_n4089_, new_n4090_, new_n4091_,
    new_n4092_, new_n4093_, new_n4094_, new_n4095_, new_n4096_, new_n4097_,
    new_n4098_, new_n4099_, new_n4100_, new_n4101_, new_n4102_, new_n4103_,
    new_n4104_, new_n4105_, new_n4106_, new_n4107_, new_n4108_, new_n4109_,
    new_n4110_, new_n4111_, new_n4112_, new_n4113_, new_n4114_, new_n4115_,
    new_n4116_, new_n4117_, new_n4118_, new_n4119_, new_n4120_, new_n4121_,
    new_n4122_, new_n4123_, new_n4124_, new_n4125_, new_n4126_, new_n4127_,
    new_n4128_, new_n4129_, new_n4130_, new_n4131_, new_n4132_, new_n4133_,
    new_n4134_, new_n4135_, new_n4136_, new_n4137_, new_n4138_, new_n4139_,
    new_n4140_, new_n4141_, new_n4142_, new_n4143_, new_n4144_, new_n4145_,
    new_n4146_, new_n4147_, new_n4148_, new_n4149_, new_n4150_, new_n4151_,
    new_n4152_, new_n4153_, new_n4155_, new_n4156_, new_n4157_, new_n4158_,
    new_n4159_, new_n4160_, new_n4161_, new_n4162_, new_n4163_, new_n4164_,
    new_n4165_, new_n4166_, new_n4167_, new_n4168_, new_n4169_, new_n4170_,
    new_n4171_, new_n4172_, new_n4173_, new_n4174_, new_n4175_, new_n4176_,
    new_n4177_, new_n4178_, new_n4179_, new_n4180_, new_n4181_, new_n4182_,
    new_n4183_, new_n4184_, new_n4185_, new_n4186_, new_n4187_, new_n4188_,
    new_n4189_, new_n4190_, new_n4191_, new_n4192_, new_n4193_, new_n4194_,
    new_n4195_, new_n4196_, new_n4197_, new_n4198_, new_n4199_, new_n4200_,
    new_n4201_, new_n4202_, new_n4203_, new_n4204_, new_n4205_, new_n4206_,
    new_n4207_, new_n4208_, new_n4209_, new_n4210_, new_n4211_, new_n4212_,
    new_n4213_, new_n4214_, new_n4215_, new_n4216_, new_n4217_, new_n4218_,
    new_n4219_, new_n4220_, new_n4221_, new_n4222_, new_n4223_, new_n4224_,
    new_n4225_, new_n4226_, new_n4227_, new_n4228_, new_n4229_, new_n4230_,
    new_n4231_, new_n4232_, new_n4233_, new_n4234_, new_n4235_, new_n4236_,
    new_n4237_, new_n4238_, new_n4239_, new_n4240_, new_n4241_, new_n4242_,
    new_n4243_, new_n4244_, new_n4245_, new_n4246_, new_n4247_, new_n4248_,
    new_n4249_, new_n4250_, new_n4251_, new_n4252_, new_n4253_, new_n4254_,
    new_n4255_, new_n4256_, new_n4257_, new_n4258_, new_n4259_, new_n4260_,
    new_n4261_, new_n4262_, new_n4263_, new_n4264_, new_n4265_, new_n4266_,
    new_n4267_, new_n4268_, new_n4269_, new_n4270_, new_n4271_, new_n4272_,
    new_n4273_, new_n4274_, new_n4275_, new_n4276_, new_n4277_, new_n4278_,
    new_n4279_, new_n4280_, new_n4281_, new_n4282_, new_n4283_, new_n4284_,
    new_n4285_, new_n4286_, new_n4287_, new_n4288_, new_n4289_, new_n4290_,
    new_n4291_, new_n4292_, new_n4293_, new_n4294_, new_n4295_, new_n4296_,
    new_n4297_, new_n4298_, new_n4299_, new_n4301_, new_n4302_, new_n4303_,
    new_n4304_, new_n4305_, new_n4306_, new_n4307_, new_n4308_, new_n4309_,
    new_n4310_, new_n4311_, new_n4312_, new_n4313_, new_n4314_, new_n4315_,
    new_n4316_, new_n4317_, new_n4318_, new_n4319_, new_n4320_, new_n4321_,
    new_n4322_, new_n4323_, new_n4324_, new_n4325_, new_n4326_, new_n4327_,
    new_n4328_, new_n4329_, new_n4330_, new_n4331_, new_n4332_, new_n4333_,
    new_n4334_, new_n4335_, new_n4336_, new_n4337_, new_n4338_, new_n4339_,
    new_n4340_, new_n4341_, new_n4342_, new_n4343_, new_n4344_, new_n4345_,
    new_n4346_, new_n4347_, new_n4348_, new_n4349_, new_n4350_, new_n4351_,
    new_n4352_, new_n4353_, new_n4354_, new_n4355_, new_n4356_, new_n4357_,
    new_n4358_, new_n4359_, new_n4360_, new_n4361_, new_n4362_, new_n4363_,
    new_n4364_, new_n4365_, new_n4366_, new_n4367_, new_n4368_, new_n4369_,
    new_n4370_, new_n4371_, new_n4372_, new_n4373_, new_n4374_, new_n4375_,
    new_n4376_, new_n4377_, new_n4378_, new_n4379_, new_n4380_, new_n4381_,
    new_n4382_, new_n4383_, new_n4384_, new_n4385_, new_n4386_, new_n4387_,
    new_n4388_, new_n4389_, new_n4390_, new_n4391_, new_n4392_, new_n4393_,
    new_n4394_, new_n4395_, new_n4396_, new_n4397_, new_n4398_, new_n4399_,
    new_n4400_, new_n4401_, new_n4402_, new_n4403_, new_n4404_, new_n4405_,
    new_n4406_, new_n4407_, new_n4408_, new_n4409_, new_n4410_, new_n4411_,
    new_n4412_, new_n4413_, new_n4414_, new_n4415_, new_n4416_, new_n4417_,
    new_n4418_, new_n4419_, new_n4420_, new_n4421_, new_n4422_, new_n4423_,
    new_n4424_, new_n4425_, new_n4426_, new_n4427_, new_n4428_, new_n4429_,
    new_n4430_, new_n4431_, new_n4432_, new_n4433_, new_n4434_, new_n4435_,
    new_n4436_, new_n4437_, new_n4438_, new_n4439_, new_n4440_, new_n4441_,
    new_n4442_, new_n4443_, new_n4444_, new_n4445_, new_n4447_, new_n4448_,
    new_n4449_, new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_,
    new_n4455_, new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_,
    new_n4461_, new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_,
    new_n4467_, new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_,
    new_n4473_, new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_,
    new_n4479_, new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_,
    new_n4485_, new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_,
    new_n4491_, new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_,
    new_n4497_, new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_,
    new_n4503_, new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_,
    new_n4509_, new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_,
    new_n4515_, new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_,
    new_n4521_, new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_,
    new_n4527_, new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_,
    new_n4533_, new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_,
    new_n4539_, new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_,
    new_n4545_, new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_,
    new_n4551_, new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_,
    new_n4557_, new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_,
    new_n4563_, new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_,
    new_n4569_, new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_,
    new_n4575_, new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_,
    new_n4581_, new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_,
    new_n4587_, new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_,
    new_n4593_, new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4747_, new_n4748_, new_n4749_, new_n4750_,
    new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_, new_n4756_,
    new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_, new_n4762_,
    new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_, new_n4768_,
    new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_, new_n4774_,
    new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_, new_n4780_,
    new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_, new_n4786_,
    new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_, new_n4792_,
    new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_, new_n4798_,
    new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_, new_n4804_,
    new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_, new_n4810_,
    new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_, new_n4816_,
    new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_, new_n4822_,
    new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_, new_n4828_,
    new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_, new_n4834_,
    new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_, new_n4840_,
    new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_, new_n4846_,
    new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_, new_n4852_,
    new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_, new_n4858_,
    new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_, new_n4864_,
    new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_, new_n4870_,
    new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_, new_n4876_,
    new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_, new_n4882_,
    new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_, new_n4888_,
    new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_, new_n4894_,
    new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_, new_n4900_,
    new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_, new_n4906_,
    new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_, new_n4912_,
    new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_, new_n4918_,
    new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_, new_n4924_,
    new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_, new_n4930_,
    new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_, new_n4936_,
    new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_, new_n4942_,
    new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_, new_n4948_,
    new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_, new_n4954_,
    new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_, new_n4960_,
    new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_, new_n4966_,
    new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4973_, new_n4974_,
    new_n4975_, new_n4976_, new_n4977_, new_n4978_, new_n4979_, new_n4980_,
    new_n4981_, new_n4982_, new_n4983_, new_n4984_, new_n4985_, new_n4986_,
    new_n4987_, new_n4988_, new_n4989_, new_n4990_, new_n4991_, new_n4992_,
    new_n4993_, new_n4994_, new_n4995_, new_n4996_, new_n4997_, new_n4998_,
    new_n4999_, new_n5000_, new_n5001_, new_n5002_, new_n5003_, new_n5004_,
    new_n5005_, new_n5006_, new_n5007_, new_n5008_, new_n5009_, new_n5010_,
    new_n5011_, new_n5012_, new_n5013_, new_n5014_, new_n5015_, new_n5016_,
    new_n5017_, new_n5018_, new_n5019_, new_n5020_, new_n5021_, new_n5023_,
    new_n5024_, new_n5025_, new_n5026_, new_n5027_, new_n5028_, new_n5029_,
    new_n5030_, new_n5031_, new_n5032_, new_n5033_, new_n5034_, new_n5035_,
    new_n5036_, new_n5037_, new_n5038_, new_n5039_, new_n5040_, new_n5041_,
    new_n5042_, new_n5043_, new_n5044_, new_n5045_, new_n5046_, new_n5047_,
    new_n5048_, new_n5049_, new_n5050_, new_n5051_, new_n5052_, new_n5053_,
    new_n5054_, new_n5055_, new_n5056_, new_n5057_, new_n5058_, new_n5059_,
    new_n5060_, new_n5061_, new_n5062_, new_n5063_, new_n5064_, new_n5065_,
    new_n5066_, new_n5067_, new_n5068_, new_n5069_, new_n5070_, new_n5071_,
    new_n5072_, new_n5073_, new_n5074_, new_n5075_, new_n5076_, new_n5077_,
    new_n5078_, new_n5079_, new_n5080_, new_n5081_, new_n5082_, new_n5083_,
    new_n5084_, new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_,
    new_n5091_, new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_,
    new_n5097_, new_n5098_, new_n5099_, new_n5102_, new_n5103_, new_n5104_,
    new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_, new_n5110_,
    new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_, new_n5116_,
    new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_, new_n5122_,
    new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_, new_n5128_,
    new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_, new_n5134_,
    new_n5136_, new_n5137_, new_n5138_, new_n5139_, new_n5140_, new_n5141_,
    new_n5142_, new_n5143_, new_n5144_, new_n5145_, new_n5146_, new_n5147_,
    new_n5148_, new_n5149_, new_n5150_, new_n5151_, new_n5152_, new_n5153_,
    new_n5154_, new_n5155_, new_n5156_, new_n5157_, new_n5158_, new_n5159_,
    new_n5160_, new_n5161_, new_n5162_, new_n5163_, new_n5164_, new_n5165_,
    new_n5166_, new_n5167_, new_n5168_, new_n5169_, new_n5170_, new_n5171_,
    new_n5172_, new_n5173_, new_n5174_, new_n5175_, new_n5176_, new_n5177_,
    new_n5178_, new_n5179_, new_n5180_, new_n5181_, new_n5182_, new_n5183_,
    new_n5184_, new_n5185_, new_n5186_, new_n5187_, new_n5188_, new_n5189_,
    new_n5190_, new_n5191_, new_n5192_, new_n5193_, new_n5194_, new_n5195_,
    new_n5196_, new_n5197_, new_n5198_, new_n5199_, new_n5200_, new_n5201_,
    new_n5202_, new_n5203_, new_n5204_, new_n5205_, new_n5206_, new_n5207_,
    new_n5208_, new_n5209_, new_n5210_, new_n5211_, new_n5212_, new_n5213_,
    new_n5214_, new_n5215_, new_n5216_, new_n5217_, new_n5218_, new_n5219_,
    new_n5220_, new_n5221_, new_n5222_, new_n5223_, new_n5224_, new_n5225_,
    new_n5226_, new_n5227_, new_n5228_, new_n5229_, new_n5230_, new_n5231_,
    new_n5232_, new_n5233_, new_n5234_, new_n5235_, new_n5236_, new_n5237_,
    new_n5238_, new_n5239_, new_n5240_, new_n5241_, new_n5242_, new_n5243_,
    new_n5244_, new_n5245_, new_n5246_, new_n5247_, new_n5248_, new_n5249_,
    new_n5250_, new_n5251_, new_n5252_, new_n5253_, new_n5254_, new_n5255_,
    new_n5256_, new_n5257_, new_n5258_, new_n5259_, new_n5260_, new_n5261_,
    new_n5262_, new_n5263_, new_n5264_, new_n5265_, new_n5266_, new_n5267_,
    new_n5268_, new_n5269_, new_n5270_, new_n5271_, new_n5272_, new_n5273_,
    new_n5274_, new_n5275_, new_n5276_, new_n5277_, new_n5278_, new_n5279_,
    new_n5280_, new_n5281_, new_n5282_, new_n5283_, new_n5284_, new_n5285_,
    new_n5286_, new_n5287_, new_n5288_, new_n5289_, new_n5290_, new_n5291_,
    new_n5292_, new_n5293_, new_n5294_, new_n5295_, new_n5296_, new_n5297_,
    new_n5298_, new_n5299_, new_n5300_, new_n5301_, new_n5302_, new_n5303_,
    new_n5304_, new_n5305_, new_n5306_, new_n5307_, new_n5308_, new_n5310_,
    new_n5311_, new_n5312_, new_n5313_, new_n5314_, new_n5315_, new_n5316_,
    new_n5317_, new_n5318_, new_n5319_, new_n5320_, new_n5321_, new_n5322_,
    new_n5323_, new_n5324_, new_n5325_, new_n5326_, new_n5327_, new_n5328_,
    new_n5329_, new_n5330_, new_n5331_, new_n5332_, new_n5333_, new_n5334_,
    new_n5335_, new_n5336_, new_n5337_, new_n5338_, new_n5339_, new_n5340_,
    new_n5341_, new_n5342_, new_n5343_, new_n5344_, new_n5345_, new_n5346_,
    new_n5347_, new_n5348_, new_n5349_, new_n5350_, new_n5351_, new_n5352_,
    new_n5353_, new_n5354_, new_n5355_, new_n5356_, new_n5357_, new_n5358_,
    new_n5359_, new_n5360_, new_n5361_, new_n5362_, new_n5363_, new_n5364_,
    new_n5365_, new_n5366_, new_n5367_, new_n5368_, new_n5369_, new_n5370_,
    new_n5371_, new_n5372_, new_n5373_, new_n5374_, new_n5375_, new_n5376_,
    new_n5377_, new_n5378_, new_n5379_, new_n5380_, new_n5381_, new_n5382_,
    new_n5383_, new_n5384_, new_n5385_, new_n5386_, new_n5387_, new_n5388_,
    new_n5389_, new_n5390_, new_n5391_, new_n5393_, new_n5394_, new_n5395_,
    new_n5396_, new_n5397_, new_n5398_, new_n5399_, new_n5400_, new_n5401_,
    new_n5402_, new_n5403_, new_n5404_, new_n5405_, new_n5406_, new_n5407_,
    new_n5408_, new_n5409_, new_n5410_, new_n5411_, new_n5412_, new_n5413_,
    new_n5414_, new_n5415_, new_n5416_, new_n5417_, new_n5418_, new_n5419_,
    new_n5420_, new_n5421_, new_n5422_, new_n5423_, new_n5424_, new_n5425_,
    new_n5426_, new_n5427_, new_n5428_, new_n5429_, new_n5430_, new_n5431_,
    new_n5432_, new_n5433_, new_n5434_, new_n5435_, new_n5436_, new_n5437_,
    new_n5438_, new_n5439_, new_n5440_, new_n5441_, new_n5442_, new_n5443_,
    new_n5444_, new_n5445_, new_n5446_, new_n5447_, new_n5448_, new_n5449_,
    new_n5450_, new_n5451_, new_n5452_, new_n5453_, new_n5454_, new_n5455_,
    new_n5456_, new_n5457_, new_n5458_, new_n5459_, new_n5460_, new_n5461_,
    new_n5462_, new_n5463_, new_n5464_, new_n5465_, new_n5466_, new_n5467_,
    new_n5468_, new_n5469_, new_n5470_, new_n5471_, new_n5472_, new_n5473_,
    new_n5474_, new_n5475_, new_n5477_, new_n5478_, new_n5479_, new_n5480_,
    new_n5481_, new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_,
    new_n5487_, new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_,
    new_n5493_, new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_,
    new_n5499_, new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_,
    new_n5505_, new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_,
    new_n5511_, new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_,
    new_n5517_, new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_,
    new_n5523_, new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_,
    new_n5529_, new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_,
    new_n5535_, new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_,
    new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_,
    new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_,
    new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_,
    new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_,
    new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_,
    new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_,
    new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_, new_n5602_,
    new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_, new_n5608_,
    new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_, new_n5614_,
    new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_, new_n5620_,
    new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_, new_n5626_,
    new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_, new_n5632_,
    new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_, new_n5638_,
    new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_, new_n5644_,
    new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_, new_n5650_,
    new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_, new_n5657_,
    new_n5658_, new_n5659_, new_n5660_, new_n5661_, new_n5662_, new_n5663_,
    new_n5664_, new_n5665_, new_n5666_, new_n5667_, new_n5668_, new_n5669_,
    new_n5670_, new_n5671_, new_n5672_, new_n5673_, new_n5674_, new_n5675_,
    new_n5676_, new_n5677_, new_n5678_, new_n5679_, new_n5680_, new_n5681_,
    new_n5682_, new_n5683_, new_n5684_, new_n5685_, new_n5686_, new_n5687_,
    new_n5688_, new_n5689_, new_n5690_, new_n5691_, new_n5692_, new_n5693_,
    new_n5694_, new_n5695_, new_n5696_, new_n5697_, new_n5698_, new_n5699_,
    new_n5700_, new_n5701_, new_n5702_, new_n5703_, new_n5704_, new_n5705_,
    new_n5706_, new_n5707_, new_n5708_, new_n5709_, new_n5710_, new_n5711_,
    new_n5712_, new_n5713_, new_n5714_, new_n5715_, new_n5717_, new_n5718_,
    new_n5719_, new_n5720_, new_n5721_, new_n5722_, new_n5723_, new_n5724_,
    new_n5725_, new_n5726_, new_n5727_, new_n5728_, new_n5729_, new_n5730_,
    new_n5731_, new_n5732_, new_n5733_, new_n5734_, new_n5735_, new_n5736_,
    new_n5737_, new_n5738_, new_n5739_, new_n5740_, new_n5741_, new_n5742_,
    new_n5743_, new_n5744_, new_n5745_, new_n5746_, new_n5747_, new_n5748_,
    new_n5749_, new_n5750_, new_n5751_, new_n5752_, new_n5753_, new_n5754_,
    new_n5755_, new_n5756_, new_n5757_, new_n5758_, new_n5759_, new_n5760_,
    new_n5761_, new_n5762_, new_n5763_, new_n5764_, new_n5765_, new_n5766_,
    new_n5767_, new_n5768_, new_n5769_, new_n5770_, new_n5771_, new_n5772_,
    new_n5773_, new_n5774_, new_n5775_, new_n5777_, new_n5778_, new_n5779_,
    new_n5780_, new_n5781_, new_n5782_, new_n5783_, new_n5784_, new_n5785_,
    new_n5786_, new_n5787_, new_n5788_, new_n5789_, new_n5790_, new_n5791_,
    new_n5792_, new_n5793_, new_n5794_, new_n5795_, new_n5796_, new_n5797_,
    new_n5798_, new_n5799_, new_n5800_, new_n5801_, new_n5802_, new_n5803_,
    new_n5804_, new_n5805_, new_n5806_, new_n5807_, new_n5808_, new_n5809_,
    new_n5810_, new_n5811_, new_n5812_, new_n5813_, new_n5814_, new_n5815_,
    new_n5816_, new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_,
    new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_,
    new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_,
    new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5850_, new_n5851_, new_n5853_, new_n5855_, new_n5857_,
    new_n5859_, new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_,
    new_n5865_, new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_,
    new_n5871_, new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_,
    new_n5877_, new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_,
    new_n5883_, new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_,
    new_n5889_, new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_,
    new_n5895_, new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_,
    new_n5901_, new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_,
    new_n5907_, new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_,
    new_n5913_, new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_,
    new_n5919_, new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_,
    new_n5925_, new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_,
    new_n5931_, new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_,
    new_n5937_, new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_,
    new_n5943_, new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_,
    new_n5949_, new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_,
    new_n5955_, new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_,
    new_n5961_, new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_,
    new_n5967_, new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_,
    new_n5973_, new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_,
    new_n5979_, new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_,
    new_n5985_, new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_,
    new_n5991_, new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_,
    new_n5997_, new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_,
    new_n6003_, new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_,
    new_n6009_, new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_,
    new_n6015_, new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_,
    new_n6021_, new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_,
    new_n6027_, new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_,
    new_n6033_, new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_,
    new_n6039_, new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_,
    new_n6045_, new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_,
    new_n6051_, new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_,
    new_n6057_, new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_,
    new_n6063_, new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_,
    new_n6069_, new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_,
    new_n6075_, new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_,
    new_n6081_, new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_,
    new_n6087_, new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_,
    new_n6093_, new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_,
    new_n6099_, new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_,
    new_n6105_, new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_,
    new_n6111_, new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_,
    new_n6117_, new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_,
    new_n6123_, new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_,
    new_n6129_, new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_,
    new_n6135_, new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_,
    new_n6141_, new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_,
    new_n6147_, new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_,
    new_n6153_, new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_,
    new_n6159_, new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_,
    new_n6165_, new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_,
    new_n6171_, new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_,
    new_n6177_, new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_,
    new_n6183_, new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_,
    new_n6189_, new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_,
    new_n6195_, new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_,
    new_n6201_, new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_,
    new_n6207_, new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_,
    new_n6213_, new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_,
    new_n6219_, new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_,
    new_n6225_, new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_,
    new_n6231_, new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_,
    new_n6237_, new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_,
    new_n6243_, new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_,
    new_n6249_, new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_,
    new_n6255_, new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_,
    new_n6261_, new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_,
    new_n6267_, new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_,
    new_n6273_, new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_,
    new_n6279_, new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_,
    new_n6285_, new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_,
    new_n6291_, new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_,
    new_n6297_, new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_,
    new_n6303_, new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_,
    new_n6309_, new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_,
    new_n6315_, new_n6316_, new_n6317_, new_n6318_, new_n6319_, new_n6320_,
    new_n6321_, new_n6322_, new_n6323_, new_n6324_, new_n6325_, new_n6326_,
    new_n6327_, new_n6328_, new_n6329_, new_n6330_, new_n6331_, new_n6332_,
    new_n6333_, new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_,
    new_n6339_, new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_,
    new_n6345_, new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_,
    new_n6351_, new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_,
    new_n6357_, new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_,
    new_n6363_, new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_,
    new_n6369_, new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_,
    new_n6375_, new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_,
    new_n6381_, new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_,
    new_n6387_, new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_,
    new_n6393_, new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_,
    new_n6399_, new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_,
    new_n6405_, new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_,
    new_n6411_, new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_,
    new_n6417_, new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_,
    new_n6423_, new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_,
    new_n6429_, new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_,
    new_n6435_, new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_,
    new_n6441_, new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_,
    new_n6447_, new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_,
    new_n6453_, new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_,
    new_n6459_, new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_,
    new_n6465_, new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_,
    new_n6471_, new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_,
    new_n6477_, new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_,
    new_n6483_, new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_,
    new_n6489_, new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_,
    new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_,
    new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_,
    new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_,
    new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_,
    new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_,
    new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_,
    new_n6574_, new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_,
    new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_,
    new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_,
    new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_,
    new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_,
    new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_,
    new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_,
    new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_,
    new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_,
    new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_,
    new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_,
    new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_,
    new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_,
    new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_,
    new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_,
    new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_,
    new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_,
    new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_,
    new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_,
    new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_,
    new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_,
    new_n6718_, new_n6720_, new_n6721_, new_n6722_, new_n6723_, new_n6725_,
    new_n6726_, new_n6727_, new_n6728_, new_n6729_, new_n6730_, new_n6731_,
    new_n6732_, new_n6733_, new_n6734_, new_n6735_, new_n6736_, new_n6737_,
    new_n6738_, new_n6739_, new_n6740_, new_n6741_, new_n6742_, new_n6743_,
    new_n6744_, new_n6745_, new_n6746_, new_n6747_, new_n6748_, new_n6749_,
    new_n6750_, new_n6751_, new_n6752_, new_n6753_, new_n6754_, new_n6755_,
    new_n6756_, new_n6757_, new_n6758_, new_n6759_, new_n6760_, new_n6761_,
    new_n6762_, new_n6763_, new_n6764_, new_n6765_, new_n6766_, new_n6767_,
    new_n6768_, new_n6769_, new_n6770_, new_n6772_, new_n6773_, new_n6774_,
    new_n6775_, new_n6776_, new_n6777_, new_n6778_, new_n6779_, new_n6780_,
    new_n6781_, new_n6783_, new_n6784_, new_n6785_, new_n6786_, new_n6787_,
    new_n6788_, new_n6789_, new_n6790_, new_n6791_, new_n6792_, new_n6793_,
    new_n6794_, new_n6795_, new_n6796_, new_n6797_, new_n6798_, new_n6799_,
    new_n6800_, new_n6801_, new_n6802_, new_n6803_, new_n6804_, new_n6805_,
    new_n6806_, new_n6807_, new_n6808_, new_n6809_, new_n6810_, new_n6811_,
    new_n6812_, new_n6813_, new_n6814_, new_n6815_, new_n6816_, new_n6817_,
    new_n6818_, new_n6819_, new_n6820_, new_n6821_, new_n6822_, new_n6823_,
    new_n6824_, new_n6825_, new_n6826_, new_n6827_, new_n6828_, new_n6829_,
    new_n6830_, new_n6831_, new_n6832_, new_n6833_, new_n6834_, new_n6835_,
    new_n6836_, new_n6837_, new_n6838_, new_n6839_, new_n6840_, new_n6841_,
    new_n6842_, new_n6843_, new_n6844_, new_n6845_, new_n6846_, new_n6847_,
    new_n6848_, new_n6849_, new_n6850_, new_n6851_, new_n6852_, new_n6853_,
    new_n6854_, new_n6855_, new_n6856_, new_n6857_, new_n6858_, new_n6859_,
    new_n6860_, new_n6861_, new_n6862_, new_n6863_, new_n6864_, new_n6865_,
    new_n6866_, new_n6867_, new_n6868_, new_n6869_, new_n6870_, new_n6871_,
    new_n6872_, new_n6873_, new_n6874_, new_n6875_, new_n6876_, new_n6877_,
    new_n6878_, new_n6879_, new_n6880_, new_n6881_, new_n6882_, new_n6883_,
    new_n6884_, new_n6885_, new_n6886_, new_n6887_, new_n6888_, new_n6889_,
    new_n6890_, new_n6891_, new_n6892_, new_n6893_, new_n6894_, new_n6895_,
    new_n6896_, new_n6897_, new_n6898_, new_n6899_, new_n6900_, new_n6901_,
    new_n6902_, new_n6903_, new_n6904_, new_n6905_, new_n6906_, new_n6907_,
    new_n6908_, new_n6909_, new_n6910_, new_n6911_, new_n6912_, new_n6913_,
    new_n6914_, new_n6915_, new_n6916_, new_n6917_, new_n6918_, new_n6919_,
    new_n6920_, new_n6921_, new_n6922_, new_n6923_, new_n6924_, new_n6925_,
    new_n6926_, new_n6927_, new_n6928_, new_n6929_, new_n6930_, new_n6931_,
    new_n6932_, new_n6933_, new_n6934_, new_n6935_, new_n6936_, new_n6937_,
    new_n6938_, new_n6939_, new_n6940_, new_n6941_, new_n6942_, new_n6943_,
    new_n6944_, new_n6945_, new_n6946_, new_n6947_, new_n6948_, new_n6949_,
    new_n6950_, new_n6951_, new_n6952_, new_n6953_, new_n6954_, new_n6955_,
    new_n6956_, new_n6957_, new_n6958_, new_n6959_, new_n6960_, new_n6961_,
    new_n6962_, new_n6963_, new_n6964_, new_n6965_, new_n6966_, new_n6967_,
    new_n6968_, new_n6969_, new_n6970_, new_n6971_, new_n6972_, new_n6973_,
    new_n6974_, new_n6975_, new_n6976_, new_n6977_, new_n6978_, new_n6979_,
    new_n6980_, new_n6981_, new_n6982_, new_n6983_, new_n6984_, new_n6985_,
    new_n6986_, new_n6987_, new_n6988_, new_n6989_, new_n6990_, new_n6991_,
    new_n6992_, new_n6993_, new_n6994_, new_n6995_, new_n6996_, new_n6997_,
    new_n6998_, new_n6999_, new_n7000_, new_n7001_, new_n7002_, new_n7003_,
    new_n7004_, new_n7005_, new_n7006_, new_n7007_, new_n7008_, new_n7009_,
    new_n7010_, new_n7011_, new_n7012_, new_n7013_, new_n7014_, new_n7015_,
    new_n7016_, new_n7017_, new_n7018_, new_n7019_, new_n7020_, new_n7021_,
    new_n7022_, new_n7023_, new_n7024_, new_n7025_, new_n7026_, new_n7027_,
    new_n7028_, new_n7029_, new_n7030_, new_n7031_, new_n7032_, new_n7033_,
    new_n7034_, new_n7035_, new_n7036_, new_n7037_, new_n7038_, new_n7039_,
    new_n7040_, new_n7041_, new_n7042_, new_n7043_, new_n7044_, new_n7045_,
    new_n7046_, new_n7047_, new_n7048_, new_n7049_, new_n7050_, new_n7051_,
    new_n7052_, new_n7053_, new_n7054_, new_n7055_, new_n7056_, new_n7057_,
    new_n7058_, new_n7059_, new_n7060_, new_n7061_, new_n7062_, new_n7063_,
    new_n7064_, new_n7065_, new_n7066_, new_n7067_, new_n7068_, new_n7069_,
    new_n7070_, new_n7071_, new_n7072_, new_n7073_, new_n7074_, new_n7075_,
    new_n7076_, new_n7077_, new_n7078_, new_n7079_, new_n7080_, new_n7081_,
    new_n7082_, new_n7083_, new_n7084_, new_n7085_, new_n7086_, new_n7087_,
    new_n7088_, new_n7089_, new_n7090_, new_n7091_, new_n7092_, new_n7093_,
    new_n7094_, new_n7095_, new_n7096_, new_n7097_, new_n7098_, new_n7099_,
    new_n7100_, new_n7101_, new_n7102_, new_n7103_, new_n7104_, new_n7105_,
    new_n7106_, new_n7107_, new_n7108_, new_n7109_, new_n7110_, new_n7111_,
    new_n7112_, new_n7113_, new_n7114_, new_n7115_, new_n7116_, new_n7117_,
    new_n7118_, new_n7119_, new_n7120_, new_n7121_, new_n7122_, new_n7123_,
    new_n7124_, new_n7125_, new_n7126_, new_n7127_, new_n7128_, new_n7129_,
    new_n7130_, new_n7131_, new_n7132_, new_n7133_, new_n7134_, new_n7135_,
    new_n7136_, new_n7137_, new_n7138_, new_n7139_, new_n7140_, new_n7141_,
    new_n7142_, new_n7143_, new_n7144_, new_n7145_, new_n7146_, new_n7147_,
    new_n7148_, new_n7149_, new_n7150_, new_n7151_, new_n7152_, new_n7153_,
    new_n7154_, new_n7155_, new_n7156_, new_n7157_, new_n7158_, new_n7159_,
    new_n7160_, new_n7161_, new_n7162_, new_n7163_, new_n7164_, new_n7165_,
    new_n7166_, new_n7167_, new_n7168_, new_n7169_, new_n7170_, new_n7171_,
    new_n7172_, new_n7173_, new_n7174_, new_n7175_, new_n7176_, new_n7177_,
    new_n7178_, new_n7179_, new_n7180_, new_n7181_, new_n7182_, new_n7183_,
    new_n7184_, new_n7185_, new_n7186_, new_n7187_, new_n7188_, new_n7189_,
    new_n7190_, new_n7191_, new_n7192_, new_n7193_, new_n7194_, new_n7195_,
    new_n7196_, new_n7197_, new_n7198_, new_n7199_, new_n7200_, new_n7201_,
    new_n7202_, new_n7203_, new_n7204_, new_n7205_, new_n7206_, new_n7207_,
    new_n7208_, new_n7209_, new_n7210_, new_n7211_, new_n7212_, new_n7213_,
    new_n7214_, new_n7215_, new_n7216_, new_n7217_, new_n7218_, new_n7219_,
    new_n7220_, new_n7221_, new_n7222_, new_n7223_, new_n7224_, new_n7225_,
    new_n7226_, new_n7227_, new_n7228_, new_n7229_, new_n7230_, new_n7231_,
    new_n7232_, new_n7233_, new_n7234_, new_n7235_, new_n7236_, new_n7237_,
    new_n7238_, new_n7239_, new_n7240_, new_n7241_, new_n7242_, new_n7243_,
    new_n7244_, new_n7245_, new_n7246_, new_n7247_, new_n7248_, new_n7249_,
    new_n7250_, new_n7251_, new_n7252_, new_n7253_, new_n7254_, new_n7255_,
    new_n7256_, new_n7257_, new_n7258_, new_n7259_, new_n7260_, new_n7261_,
    new_n7262_, new_n7263_, new_n7264_, new_n7265_, new_n7266_, new_n7267_,
    new_n7268_, new_n7269_, new_n7270_, new_n7271_, new_n7272_, new_n7273_,
    new_n7274_, new_n7275_, new_n7276_, new_n7277_, new_n7278_, new_n7279_,
    new_n7280_, new_n7281_, new_n7282_, new_n7283_, new_n7284_, new_n7285_,
    new_n7286_, new_n7287_, new_n7288_, new_n7289_, new_n7290_, new_n7291_,
    new_n7292_, new_n7293_, new_n7294_, new_n7295_, new_n7296_, new_n7297_,
    new_n7298_, new_n7299_, new_n7301_, new_n7303_, new_n7304_, new_n7305_,
    new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_,
    new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_,
    new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7552_,
    new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_, new_n7558_,
    new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_, new_n7564_,
    new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_, new_n7570_,
    new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_, new_n7576_,
    new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_, new_n7582_,
    new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_, new_n7588_,
    new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_, new_n7594_,
    new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7600_, new_n7601_,
    new_n7602_, new_n7603_, new_n7604_, new_n7605_, new_n7606_, new_n7607_,
    new_n7608_, new_n7609_, new_n7611_, new_n7612_, new_n7613_, new_n7614_,
    new_n7615_, new_n7616_, new_n7617_, new_n7618_, new_n7619_, new_n7620_,
    new_n7621_, new_n7622_, new_n7623_, new_n7624_, new_n7625_, new_n7626_,
    new_n7628_, new_n7629_, new_n7630_, new_n7631_, new_n7632_, new_n7633_,
    new_n7634_, new_n7635_, new_n7636_, new_n7637_, new_n7638_, new_n7639_,
    new_n7640_, new_n7641_, new_n7642_, new_n7643_, new_n7644_, new_n7645_,
    new_n7646_, new_n7647_, new_n7648_, new_n7649_, new_n7650_, new_n7651_,
    new_n7652_, new_n7653_, new_n7654_, new_n7655_, new_n7656_, new_n7657_,
    new_n7658_, new_n7659_, new_n7660_, new_n7661_, new_n7662_, new_n7663_,
    new_n7664_, new_n7665_, new_n7666_, new_n7667_, new_n7668_, new_n7669_,
    new_n7670_, new_n7671_, new_n7672_, new_n7673_, new_n7674_, new_n7675_,
    new_n7676_, new_n7677_, new_n7678_, new_n7679_, new_n7680_, new_n7682_,
    new_n7683_, new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_,
    new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_,
    new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_,
    new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_,
    new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_,
    new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7826_, new_n7827_, new_n7828_,
    new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_, new_n7834_,
    new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_, new_n7840_,
    new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_, new_n7846_,
    new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_, new_n7852_,
    new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_, new_n7858_,
    new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_, new_n7864_,
    new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_, new_n7870_,
    new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_, new_n7876_,
    new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_, new_n7882_,
    new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_, new_n7888_,
    new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_, new_n7894_,
    new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_, new_n7900_,
    new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_, new_n7906_,
    new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_, new_n7912_,
    new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_, new_n7918_,
    new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_, new_n7924_,
    new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_, new_n7930_,
    new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_, new_n7936_,
    new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_, new_n7942_,
    new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_, new_n7948_,
    new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_, new_n7954_,
    new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_, new_n7960_,
    new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_, new_n7966_,
    new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_, new_n7972_,
    new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_, new_n7978_,
    new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_, new_n7984_,
    new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_, new_n7990_,
    new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7996_, new_n7997_,
    new_n7998_, new_n7999_, new_n8000_, new_n8001_, new_n8002_, new_n8003_,
    new_n8004_, new_n8005_, new_n8006_, new_n8007_, new_n8008_, new_n8009_,
    new_n8010_, new_n8011_, new_n8012_, new_n8013_, new_n8014_, new_n8015_,
    new_n8016_, new_n8017_, new_n8018_, new_n8019_, new_n8020_, new_n8021_,
    new_n8022_, new_n8023_, new_n8024_, new_n8025_, new_n8026_, new_n8027_,
    new_n8028_, new_n8029_, new_n8030_, new_n8031_, new_n8032_, new_n8033_,
    new_n8034_, new_n8035_, new_n8036_, new_n8037_, new_n8038_, new_n8039_,
    new_n8040_, new_n8041_, new_n8042_, new_n8043_, new_n8044_, new_n8045_,
    new_n8046_, new_n8047_, new_n8048_, new_n8049_, new_n8050_, new_n8051_,
    new_n8052_, new_n8053_, new_n8054_, new_n8055_, new_n8056_, new_n8057_,
    new_n8058_, new_n8059_, new_n8060_, new_n8061_, new_n8062_, new_n8063_,
    new_n8064_, new_n8065_, new_n8066_, new_n8067_, new_n8068_, new_n8069_,
    new_n8070_, new_n8071_, new_n8072_, new_n8073_, new_n8074_, new_n8075_,
    new_n8076_, new_n8077_, new_n8078_, new_n8079_, new_n8080_, new_n8081_,
    new_n8082_, new_n8083_, new_n8084_, new_n8085_, new_n8086_, new_n8087_,
    new_n8088_, new_n8089_, new_n8090_, new_n8091_, new_n8092_, new_n8093_,
    new_n8094_, new_n8095_, new_n8096_, new_n8097_, new_n8098_, new_n8099_,
    new_n8100_, new_n8101_, new_n8102_, new_n8103_, new_n8104_, new_n8105_,
    new_n8106_, new_n8107_, new_n8108_, new_n8109_, new_n8110_, new_n8111_,
    new_n8112_, new_n8113_, new_n8114_, new_n8116_, new_n8117_, new_n8118_,
    new_n8119_, new_n8120_, new_n8121_, new_n8122_, new_n8123_, new_n8124_,
    new_n8125_, new_n8126_, new_n8127_, new_n8128_, new_n8129_, new_n8130_,
    new_n8131_, new_n8132_, new_n8133_, new_n8134_, new_n8135_, new_n8136_,
    new_n8137_, new_n8138_, new_n8139_, new_n8140_, new_n8141_, new_n8142_,
    new_n8143_, new_n8144_, new_n8145_, new_n8146_, new_n8147_, new_n8148_,
    new_n8149_, new_n8150_, new_n8151_, new_n8152_, new_n8153_, new_n8154_,
    new_n8155_, new_n8156_, new_n8157_, new_n8158_, new_n8159_, new_n8160_,
    new_n8161_, new_n8162_, new_n8163_, new_n8164_, new_n8165_, new_n8166_,
    new_n8167_, new_n8169_, new_n8170_, new_n8172_, new_n8173_, new_n8174_,
    new_n8175_, new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_,
    new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_,
    new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_,
    new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_,
    new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_,
    new_n8213_, new_n8214_, new_n8216_, new_n8217_, new_n8218_, new_n8219_,
    new_n8220_, new_n8221_, new_n8222_, new_n8223_, new_n8224_, new_n8225_,
    new_n8227_, new_n8228_, new_n8229_, new_n8230_, new_n8231_, new_n8232_,
    new_n8233_, new_n8234_, new_n8235_, new_n8236_, new_n8237_, new_n8238_,
    new_n8239_, new_n8240_, new_n8241_, new_n8243_, new_n8244_, new_n8245_,
    new_n8246_, new_n8247_, new_n8249_, new_n8250_, new_n8251_, new_n8252_,
    new_n8253_, new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_,
    new_n8259_, new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_,
    new_n8265_, new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_,
    new_n8271_, new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_,
    new_n8277_, new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_,
    new_n8283_, new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_,
    new_n8289_, new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_,
    new_n8295_, new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_,
    new_n8301_, new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_,
    new_n8307_, new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_,
    new_n8313_, new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_,
    new_n8319_, new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_,
    new_n8325_, new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_,
    new_n8331_, new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_,
    new_n8337_, new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_,
    new_n8343_, new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8349_,
    new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8355_, new_n8356_,
    new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_, new_n8362_,
    new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8368_, new_n8369_,
    new_n8370_, new_n8371_, new_n8372_, new_n8373_, new_n8375_, new_n8376_,
    new_n8377_, new_n8378_, new_n8379_, new_n8381_, new_n8382_, new_n8383_,
    new_n8384_, new_n8385_, new_n8386_, new_n8387_, new_n8388_, new_n8390_,
    new_n8391_, new_n8393_, new_n8394_, new_n8395_, new_n8397_, new_n8398_,
    new_n8399_, new_n8400_, new_n8402_, new_n8403_, new_n8405_, new_n8406_,
    new_n8407_, new_n8409_, new_n8410_, new_n8411_, new_n8413_, new_n8414_,
    new_n8415_, new_n8416_, new_n8417_, new_n8419_, new_n8420_, new_n8422_,
    new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_, new_n8428_,
    new_n8429_, new_n8430_, new_n8432_, new_n8434_, new_n8435_, new_n8436_,
    new_n8437_, new_n8438_, new_n8440_, new_n8441_, new_n8442_, new_n8443_,
    new_n8444_, new_n8445_, new_n8446_, new_n8447_, new_n8449_, new_n8450_,
    new_n8451_, new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_,
    new_n8457_, new_n8458_, new_n8459_, new_n8460_, new_n8462_, new_n8463_,
    new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_,
    new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_,
    new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_, new_n8482_,
    new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_, new_n8489_,
    new_n8490_, new_n8491_, new_n8492_, new_n8493_, new_n8494_, new_n8495_,
    new_n8496_, new_n8498_, new_n8499_, new_n8500_, new_n8501_, new_n8502_,
    new_n8503_, new_n8504_, new_n8505_, new_n8507_, new_n8508_, new_n8509_,
    new_n8510_, new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_,
    new_n8517_, new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_,
    new_n8523_, new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_,
    new_n8529_, new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_,
    new_n8535_, new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_,
    new_n8541_, new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_,
    new_n8547_, new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_,
    new_n8553_, new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_,
    new_n8559_, new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_,
    new_n8565_, new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_,
    new_n8571_, new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_,
    new_n8577_, new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_,
    new_n8583_, new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_,
    new_n8589_, new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_,
    new_n8595_, new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_,
    new_n8601_, new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_,
    new_n8607_, new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8621_, new_n8623_, new_n8624_, new_n8625_, new_n8626_, new_n8627_,
    new_n8628_, new_n8629_, new_n8630_, new_n8631_, new_n8632_, new_n8633_,
    new_n8634_, new_n8635_, new_n8636_, new_n8637_, new_n8638_, new_n8639_,
    new_n8640_, new_n8641_, new_n8642_, new_n8643_, new_n8644_, new_n8645_,
    new_n8646_, new_n8647_, new_n8648_, new_n8649_, new_n8650_, new_n8651_,
    new_n8652_, new_n8653_, new_n8654_, new_n8655_, new_n8656_, new_n8657_,
    new_n8658_, new_n8659_, new_n8660_, new_n8661_, new_n8662_, new_n8663_,
    new_n8664_, new_n8665_, new_n8666_, new_n8667_, new_n8668_, new_n8669_,
    new_n8670_, new_n8671_, new_n8672_, new_n8673_, new_n8674_, new_n8675_,
    new_n8676_, new_n8677_, new_n8678_, new_n8679_, new_n8680_, new_n8681_,
    new_n8682_, new_n8683_, new_n8684_, new_n8685_, new_n8686_, new_n8687_,
    new_n8688_, new_n8689_, new_n8690_, new_n8691_, new_n8692_, new_n8693_,
    new_n8694_, new_n8695_, new_n8696_, new_n8697_, new_n8698_, new_n8699_,
    new_n8700_, new_n8701_, new_n8702_, new_n8703_, new_n8704_, new_n8705_,
    new_n8706_, new_n8707_, new_n8708_, new_n8709_, new_n8710_, new_n8711_,
    new_n8712_, new_n8713_, new_n8714_, new_n8715_, new_n8716_, new_n8717_,
    new_n8718_, new_n8719_, new_n8720_, new_n8721_, new_n8722_, new_n8723_,
    new_n8724_, new_n8725_, new_n8726_, new_n8727_, new_n8728_, new_n8729_,
    new_n8730_, new_n8731_, new_n8732_, new_n8733_, new_n8734_, new_n8735_,
    new_n8736_, new_n8737_, new_n8738_, new_n8739_, new_n8740_, new_n8741_,
    new_n8742_, new_n8743_, new_n8744_, new_n8745_, new_n8746_, new_n8747_,
    new_n8748_, new_n8749_, new_n8750_, new_n8751_, new_n8752_, new_n8753_,
    new_n8754_, new_n8755_, new_n8756_, new_n8757_, new_n8758_, new_n8759_,
    new_n8760_, new_n8761_, new_n8762_, new_n8763_, new_n8764_, new_n8765_,
    new_n8766_, new_n8767_, new_n8768_, new_n8769_, new_n8770_, new_n8771_,
    new_n8772_, new_n8773_, new_n8774_, new_n8775_, new_n8776_, new_n8777_,
    new_n8778_, new_n8779_, new_n8780_, new_n8781_, new_n8782_, new_n8783_,
    new_n8784_, new_n8785_, new_n8786_, new_n8787_, new_n8788_, new_n8789_,
    new_n8790_, new_n8791_, new_n8792_, new_n8793_, new_n8794_, new_n8795_,
    new_n8796_, new_n8797_, new_n8798_, new_n8799_, new_n8800_, new_n8801_,
    new_n8802_, new_n8803_, new_n8804_, new_n8805_, new_n8806_, new_n8807_,
    new_n8808_, new_n8809_, new_n8810_, new_n8811_, new_n8812_, new_n8813_,
    new_n8814_, new_n8815_, new_n8816_, new_n8817_, new_n8818_, new_n8819_,
    new_n8820_, new_n8821_, new_n8822_, new_n8823_, new_n8824_, new_n8825_,
    new_n8826_, new_n8827_, new_n8828_, new_n8829_, new_n8830_, new_n8831_,
    new_n8832_, new_n8833_, new_n8834_, new_n8835_, new_n8836_, new_n8837_,
    new_n8838_, new_n8839_, new_n8840_, new_n8841_, new_n8842_, new_n8843_,
    new_n8844_, new_n8845_, new_n8846_, new_n8847_, new_n8848_, new_n8849_,
    new_n8850_, new_n8851_, new_n8852_, new_n8853_, new_n8854_, new_n8855_,
    new_n8856_, new_n8857_, new_n8858_, new_n8859_, new_n8860_, new_n8861_,
    new_n8862_, new_n8863_, new_n8864_, new_n8865_, new_n8866_, new_n8867_,
    new_n8868_, new_n8869_, new_n8870_, new_n8871_, new_n8872_, new_n8873_,
    new_n8874_, new_n8875_, new_n8876_, new_n8877_, new_n8878_, new_n8879_,
    new_n8880_, new_n8881_, new_n8882_, new_n8883_, new_n8884_, new_n8885_,
    new_n8886_, new_n8887_, new_n8888_, new_n8889_, new_n8890_, new_n8891_,
    new_n8892_, new_n8893_, new_n8894_, new_n8895_, new_n8896_, new_n8897_,
    new_n8898_, new_n8899_, new_n8900_, new_n8901_, new_n8902_, new_n8903_,
    new_n8904_, new_n8905_, new_n8906_, new_n8907_, new_n8908_, new_n8909_,
    new_n8910_, new_n8911_, new_n8912_, new_n8913_, new_n8914_, new_n8915_,
    new_n8916_, new_n8917_, new_n8918_, new_n8919_, new_n8920_, new_n8921_,
    new_n8922_, new_n8923_, new_n8924_, new_n8925_, new_n8926_, new_n8927_,
    new_n8928_, new_n8929_, new_n8930_, new_n8931_, new_n8932_, new_n8933_,
    new_n8934_, new_n8935_, new_n8936_, new_n8937_, new_n8938_, new_n8939_,
    new_n8940_, new_n8941_, new_n8943_, new_n8944_, new_n8945_, new_n8946_,
    new_n8947_, new_n8948_, new_n8949_, new_n8950_, new_n8951_, new_n8952_,
    new_n8953_, new_n8954_, new_n8955_, new_n8956_, new_n8957_, new_n8958_,
    new_n8959_, new_n8960_, new_n8961_, new_n8962_, new_n8963_, new_n8964_,
    new_n8965_, new_n8966_, new_n8967_, new_n8968_, new_n8969_, new_n8970_,
    new_n8971_, new_n8972_, new_n8973_, new_n8974_, new_n8975_, new_n8976_,
    new_n8977_, new_n8978_, new_n8979_, new_n8980_, new_n8981_, new_n8982_,
    new_n8983_, new_n8984_, new_n8985_, new_n8986_, new_n8987_, new_n8988_,
    new_n8989_, new_n8990_, new_n8991_, new_n8992_, new_n8993_, new_n8994_,
    new_n8995_, new_n8996_, new_n8997_, new_n8998_, new_n8999_, new_n9000_,
    new_n9001_, new_n9002_, new_n9003_, new_n9004_, new_n9005_, new_n9006_,
    new_n9007_, new_n9008_, new_n9009_, new_n9010_, new_n9011_, new_n9012_,
    new_n9013_, new_n9014_, new_n9015_, new_n9016_, new_n9017_, new_n9018_,
    new_n9019_, new_n9020_, new_n9021_, new_n9022_, new_n9023_, new_n9024_,
    new_n9025_, new_n9026_, new_n9027_, new_n9028_, new_n9029_, new_n9030_,
    new_n9031_, new_n9032_, new_n9033_, new_n9034_, new_n9035_, new_n9036_,
    new_n9037_, new_n9038_, new_n9039_, new_n9040_, new_n9041_, new_n9042_,
    new_n9043_, new_n9044_, new_n9045_, new_n9046_, new_n9047_, new_n9048_,
    new_n9049_, new_n9050_, new_n9051_, new_n9052_, new_n9053_, new_n9054_,
    new_n9055_, new_n9056_, new_n9057_, new_n9058_, new_n9059_, new_n9060_,
    new_n9061_, new_n9062_, new_n9063_, new_n9064_, new_n9065_, new_n9066_,
    new_n9067_, new_n9068_, new_n9069_, new_n9070_, new_n9071_, new_n9072_,
    new_n9073_, new_n9074_, new_n9075_, new_n9076_, new_n9077_, new_n9078_,
    new_n9079_, new_n9080_, new_n9081_, new_n9082_, new_n9083_, new_n9084_,
    new_n9085_, new_n9086_, new_n9087_, new_n9088_, new_n9089_, new_n9090_,
    new_n9091_, new_n9092_, new_n9093_, new_n9094_, new_n9095_, new_n9096_,
    new_n9097_, new_n9098_, new_n9099_, new_n9100_, new_n9101_, new_n9102_,
    new_n9103_, new_n9104_, new_n9105_, new_n9106_, new_n9107_, new_n9108_,
    new_n9109_, new_n9110_, new_n9111_, new_n9112_, new_n9113_, new_n9114_,
    new_n9115_, new_n9116_, new_n9117_, new_n9118_, new_n9119_, new_n9120_,
    new_n9121_, new_n9122_, new_n9123_, new_n9124_, new_n9125_, new_n9126_,
    new_n9127_, new_n9128_, new_n9129_, new_n9130_, new_n9131_, new_n9132_,
    new_n9133_, new_n9134_, new_n9135_, new_n9136_, new_n9137_, new_n9138_,
    new_n9139_, new_n9140_, new_n9141_, new_n9142_, new_n9143_, new_n9144_,
    new_n9145_, new_n9146_, new_n9147_, new_n9148_, new_n9149_, new_n9150_,
    new_n9151_, new_n9152_, new_n9153_, new_n9154_, new_n9155_, new_n9156_,
    new_n9157_, new_n9158_, new_n9159_, new_n9160_, new_n9161_, new_n9162_,
    new_n9163_, new_n9164_, new_n9165_, new_n9166_, new_n9167_, new_n9168_,
    new_n9169_, new_n9170_, new_n9171_, new_n9172_, new_n9173_, new_n9174_,
    new_n9175_, new_n9176_, new_n9177_, new_n9178_, new_n9179_, new_n9180_,
    new_n9181_, new_n9182_, new_n9183_, new_n9184_, new_n9185_, new_n9186_,
    new_n9187_, new_n9188_, new_n9189_, new_n9190_, new_n9191_, new_n9192_,
    new_n9193_, new_n9194_, new_n9195_, new_n9196_, new_n9197_, new_n9198_,
    new_n9199_, new_n9200_, new_n9201_, new_n9202_, new_n9203_, new_n9204_,
    new_n9205_, new_n9206_, new_n9207_, new_n9208_, new_n9209_, new_n9210_,
    new_n9211_, new_n9212_, new_n9213_, new_n9214_, new_n9215_, new_n9216_,
    new_n9217_, new_n9218_, new_n9219_, new_n9220_, new_n9221_, new_n9222_,
    new_n9223_, new_n9224_, new_n9225_, new_n9226_, new_n9227_, new_n9228_,
    new_n9229_, new_n9230_, new_n9231_, new_n9232_, new_n9233_, new_n9234_,
    new_n9235_, new_n9236_, new_n9237_, new_n9238_, new_n9239_, new_n9240_,
    new_n9241_, new_n9242_, new_n9243_, new_n9244_, new_n9245_, new_n9246_,
    new_n9247_, new_n9248_, new_n9249_, new_n9250_, new_n9251_, new_n9252_,
    new_n9253_, new_n9254_, new_n9255_, new_n9256_, new_n9257_, new_n9258_,
    new_n9259_, new_n9260_, new_n9261_, new_n9262_, new_n9263_, new_n9264_,
    new_n9265_, new_n9266_, new_n9267_, new_n9268_, new_n9269_, new_n9270_,
    new_n9271_, new_n9272_, new_n9273_, new_n9274_, new_n9275_, new_n9276_,
    new_n9277_, new_n9278_, new_n9279_, new_n9280_, new_n9281_, new_n9282_,
    new_n9283_, new_n9284_, new_n9285_, new_n9286_, new_n9287_, new_n9288_,
    new_n9289_, new_n9290_, new_n9291_, new_n9292_, new_n9293_, new_n9294_,
    new_n9295_, new_n9296_, new_n9297_, new_n9298_, new_n9299_, new_n9300_,
    new_n9301_, new_n9302_, new_n9303_, new_n9304_, new_n9305_, new_n9306_,
    new_n9307_, new_n9308_, new_n9309_, new_n9310_, new_n9311_, new_n9312_,
    new_n9313_, new_n9314_, new_n9315_, new_n9316_, new_n9317_, new_n9318_,
    new_n9319_, new_n9320_, new_n9321_, new_n9322_, new_n9323_, new_n9324_,
    new_n9325_, new_n9326_, new_n9327_, new_n9328_, new_n9329_, new_n9330_,
    new_n9331_, new_n9332_, new_n9333_, new_n9334_, new_n9335_, new_n9336_,
    new_n9337_, new_n9338_, new_n9339_, new_n9340_, new_n9341_, new_n9342_,
    new_n9343_, new_n9344_, new_n9345_, new_n9346_, new_n9347_, new_n9348_,
    new_n9349_, new_n9350_, new_n9351_, new_n9352_, new_n9353_, new_n9354_,
    new_n9355_, new_n9356_, new_n9357_, new_n9358_, new_n9359_, new_n9360_,
    new_n9361_, new_n9362_, new_n9363_, new_n9364_, new_n9365_, new_n9366_,
    new_n9367_, new_n9368_, new_n9369_, new_n9370_, new_n9371_, new_n9372_,
    new_n9373_, new_n9374_, new_n9375_, new_n9376_, new_n9377_, new_n9378_,
    new_n9379_, new_n9380_, new_n9381_, new_n9382_, new_n9383_, new_n9384_,
    new_n9385_, new_n9386_, new_n9387_, new_n9388_, new_n9389_, new_n9390_,
    new_n9391_, new_n9392_, new_n9393_, new_n9394_, new_n9395_, new_n9396_,
    new_n9397_, new_n9398_, new_n9399_, new_n9400_, new_n9401_, new_n9402_,
    new_n9403_, new_n9404_, new_n9405_, new_n9406_, new_n9407_, new_n9408_,
    new_n9409_, new_n9410_, new_n9411_, new_n9412_, new_n9413_, new_n9414_,
    new_n9415_, new_n9416_, new_n9417_, new_n9418_, new_n9419_, new_n9420_,
    new_n9421_, new_n9422_, new_n9423_, new_n9424_, new_n9426_, new_n9427_,
    new_n9428_, new_n9429_, new_n9430_, new_n9431_, new_n9433_, new_n9434_,
    new_n9435_, new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_,
    new_n9442_, new_n9443_, new_n9445_, new_n9446_, new_n9447_, new_n9448_,
    new_n9449_, new_n9451_, new_n9452_, new_n9453_, new_n9454_, new_n9456_,
    new_n9457_, new_n9459_, new_n9461_, new_n9462_, new_n9463_, new_n9464_,
    new_n9465_, new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_,
    new_n9471_, new_n9472_, new_n9474_, new_n9475_, new_n9476_, new_n9477_,
    new_n9478_, new_n9479_, new_n9481_, new_n9483_, new_n9484_, new_n9485_,
    new_n9486_, new_n9487_, new_n9488_, new_n9489_, new_n9491_, new_n9492_,
    new_n9493_, new_n9494_, new_n9495_, new_n9496_, new_n9498_, new_n9499_,
    new_n9500_, new_n9501_, new_n9503_, new_n9504_, new_n9505_, new_n9506_,
    new_n9507_, new_n9508_, new_n9509_, new_n9510_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9523_, new_n9524_, new_n9525_, new_n9526_,
    new_n9527_, new_n9528_, new_n9529_, new_n9531_, new_n9532_, new_n9533_,
    new_n9534_, new_n9536_, new_n9537_, new_n9539_, new_n9540_, new_n9541_,
    new_n9542_, new_n9543_, new_n9544_, new_n9545_, new_n9546_, new_n9547_,
    new_n9548_, new_n9549_, new_n9550_, new_n9551_, new_n9552_, new_n9553_,
    new_n9554_, new_n9555_, new_n9556_, new_n9557_, new_n9558_, new_n9559_,
    new_n9560_, new_n9561_, new_n9562_, new_n9563_, new_n9564_, new_n9565_,
    new_n9566_, new_n9567_, new_n9568_, new_n9569_, new_n9570_, new_n9571_,
    new_n9572_, new_n9573_, new_n9574_, new_n9575_, new_n9576_, new_n9577_,
    new_n9578_, new_n9579_, new_n9580_, new_n9581_, new_n9582_, new_n9583_,
    new_n9584_, new_n9585_, new_n9586_, new_n9587_, new_n9588_, new_n9590_,
    new_n9591_, new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_,
    new_n9597_, new_n9598_, new_n9599_, new_n9600_, new_n9602_, new_n9603_,
    new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_,
    new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_,
    new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_,
    new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9655_, new_n9657_, new_n9658_, new_n9659_,
    new_n9660_, new_n9661_, new_n9663_, new_n9664_, new_n9665_, new_n9666_,
    new_n9667_, new_n9668_, new_n9669_, new_n9670_, new_n9671_, new_n9672_,
    new_n9673_, new_n9674_, new_n9676_, new_n9677_, new_n9678_, new_n9679_,
    new_n9680_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9695_, new_n9697_, new_n9698_, new_n9699_, new_n9700_, new_n9701_,
    new_n9703_, new_n9704_, new_n9705_, new_n9708_, new_n9709_, new_n9710_,
    new_n9711_, new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_,
    new_n9717_, new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_,
    new_n9723_, new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_,
    new_n9729_, new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_,
    new_n9735_, new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9769_, new_n9770_, new_n9771_, new_n9772_,
    new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_, new_n9778_,
    new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_, new_n9784_,
    new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_, new_n9790_,
    new_n9791_, new_n9792_, new_n9794_, new_n9795_, new_n9796_, new_n9797_,
    new_n9798_, new_n9799_, new_n9800_, new_n9801_, new_n9802_, new_n9803_,
    new_n9804_, new_n9805_, new_n9806_, new_n9807_, new_n9808_, new_n9809_,
    new_n9810_, new_n9811_, new_n9812_, new_n9813_, new_n9814_, new_n9815_,
    new_n9816_, new_n9817_, new_n9818_, new_n9819_, new_n9820_, new_n9821_,
    new_n9822_, new_n9823_, new_n9824_, new_n9825_, new_n9827_, new_n9828_,
    new_n9829_, new_n9830_, new_n9831_, new_n9832_, new_n9833_, new_n9834_,
    new_n9836_, new_n9837_, new_n9838_, new_n9839_, new_n9840_, new_n9841_,
    new_n9842_, new_n9843_, new_n9844_, new_n9845_, new_n9846_, new_n9847_,
    new_n9848_, new_n9849_, new_n9850_, new_n9851_, new_n9852_, new_n9853_,
    new_n9854_, new_n9855_, new_n9856_, new_n9857_, new_n9858_, new_n9859_,
    new_n9860_, new_n9861_, new_n9862_, new_n9863_, new_n9864_, new_n9865_,
    new_n9866_, new_n9867_, new_n9868_, new_n9869_, new_n9870_, new_n9871_,
    new_n9872_, new_n9873_, new_n9874_, new_n9875_, new_n9876_, new_n9877_,
    new_n9878_, new_n9879_, new_n9880_, new_n9881_, new_n9882_, new_n9883_,
    new_n9884_, new_n9885_, new_n9886_, new_n9887_, new_n9888_, new_n9889_,
    new_n9890_, new_n9891_, new_n9892_, new_n9893_, new_n9894_, new_n9895_,
    new_n9896_, new_n9897_, new_n9898_, new_n9899_, new_n9900_, new_n9901_,
    new_n9902_, new_n9903_, new_n9904_, new_n9905_, new_n9906_, new_n9907_,
    new_n9908_, new_n9909_, new_n9910_, new_n9911_, new_n9912_, new_n9913_,
    new_n9914_, new_n9915_, new_n9916_, new_n9917_, new_n9918_, new_n9919_,
    new_n9920_, new_n9921_, new_n9922_, new_n9923_, new_n9924_, new_n9925_,
    new_n9926_, new_n9927_, new_n9928_, new_n9929_, new_n9930_, new_n9931_,
    new_n9932_, new_n9933_, new_n9934_, new_n9935_, new_n9936_, new_n9937_,
    new_n9938_, new_n9939_, new_n9940_, new_n9941_, new_n9942_, new_n9943_,
    new_n9944_, new_n9945_, new_n9946_, new_n9947_, new_n9948_, new_n9949_,
    new_n9950_, new_n9951_, new_n9952_, new_n9953_, new_n9954_, new_n9955_,
    new_n9956_, new_n9957_, new_n9958_, new_n9959_, new_n9960_, new_n9961_,
    new_n9962_, new_n9963_, new_n9964_, new_n9965_, new_n9966_, new_n9967_,
    new_n9968_, new_n9969_, new_n9970_, new_n9971_, new_n9972_, new_n9973_,
    new_n9974_, new_n9975_, new_n9976_, new_n9977_, new_n9978_, new_n9979_,
    new_n9980_, new_n9981_, new_n9982_, new_n9983_, new_n9984_, new_n9985_,
    new_n9986_, new_n9987_, new_n9988_, new_n9989_, new_n9990_, new_n9991_,
    new_n9992_, new_n9993_, new_n9994_, new_n9995_, new_n9996_, new_n9997_,
    new_n9998_, new_n9999_, new_n10000_, new_n10001_, new_n10002_,
    new_n10003_, new_n10004_, new_n10005_, new_n10006_, new_n10007_,
    new_n10008_, new_n10009_, new_n10010_, new_n10011_, new_n10012_,
    new_n10013_, new_n10014_, new_n10015_, new_n10016_, new_n10017_,
    new_n10018_, new_n10019_, new_n10020_, new_n10021_, new_n10022_,
    new_n10023_, new_n10024_, new_n10025_, new_n10026_, new_n10027_,
    new_n10028_, new_n10029_, new_n10030_, new_n10031_, new_n10032_,
    new_n10033_, new_n10034_, new_n10035_, new_n10036_, new_n10037_,
    new_n10038_, new_n10039_, new_n10041_, new_n10042_, new_n10043_,
    new_n10044_, new_n10045_, new_n10046_, new_n10047_, new_n10048_,
    new_n10049_, new_n10050_, new_n10051_, new_n10052_, new_n10053_,
    new_n10054_, new_n10055_, new_n10056_, new_n10057_, new_n10058_,
    new_n10059_, new_n10060_, new_n10061_, new_n10062_, new_n10063_,
    new_n10064_, new_n10065_, new_n10066_, new_n10067_, new_n10068_,
    new_n10069_, new_n10070_, new_n10071_, new_n10072_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10334_, new_n10335_,
    new_n10336_, new_n10337_, new_n10338_, new_n10339_, new_n10340_,
    new_n10341_, new_n10342_, new_n10343_, new_n10344_, new_n10345_,
    new_n10346_, new_n10347_, new_n10348_, new_n10349_, new_n10350_,
    new_n10351_, new_n10352_, new_n10353_, new_n10354_, new_n10355_,
    new_n10356_, new_n10357_, new_n10358_, new_n10359_, new_n10360_,
    new_n10361_, new_n10362_, new_n10363_, new_n10364_, new_n10365_,
    new_n10366_, new_n10367_, new_n10368_, new_n10369_, new_n10370_,
    new_n10371_, new_n10372_, new_n10373_, new_n10374_, new_n10375_,
    new_n10376_, new_n10377_, new_n10378_, new_n10379_, new_n10380_,
    new_n10381_, new_n10382_, new_n10383_, new_n10384_, new_n10385_,
    new_n10386_, new_n10387_, new_n10388_, new_n10389_, new_n10390_,
    new_n10391_, new_n10392_, new_n10393_, new_n10394_, new_n10395_,
    new_n10396_, new_n10397_, new_n10398_, new_n10399_, new_n10400_,
    new_n10401_, new_n10402_, new_n10403_, new_n10404_, new_n10405_,
    new_n10406_, new_n10407_, new_n10408_, new_n10409_, new_n10410_,
    new_n10411_, new_n10412_, new_n10413_, new_n10414_, new_n10415_,
    new_n10416_, new_n10417_, new_n10418_, new_n10419_, new_n10420_,
    new_n10421_, new_n10422_, new_n10423_, new_n10424_, new_n10425_,
    new_n10426_, new_n10427_, new_n10428_, new_n10429_, new_n10430_,
    new_n10431_, new_n10432_, new_n10433_, new_n10434_, new_n10435_,
    new_n10436_, new_n10437_, new_n10438_, new_n10439_, new_n10440_,
    new_n10441_, new_n10442_, new_n10443_, new_n10444_, new_n10445_,
    new_n10446_, new_n10447_, new_n10448_, new_n10449_, new_n10450_,
    new_n10451_, new_n10452_, new_n10453_, new_n10454_, new_n10455_,
    new_n10456_, new_n10457_, new_n10458_, new_n10459_, new_n10460_,
    new_n10461_, new_n10462_, new_n10463_, new_n10464_, new_n10465_,
    new_n10466_, new_n10467_, new_n10468_, new_n10469_, new_n10470_,
    new_n10471_, new_n10472_, new_n10473_, new_n10474_, new_n10475_,
    new_n10476_, new_n10477_, new_n10478_, new_n10479_, new_n10480_,
    new_n10481_, new_n10482_, new_n10483_, new_n10484_, new_n10485_,
    new_n10486_, new_n10487_, new_n10488_, new_n10489_, new_n10490_,
    new_n10491_, new_n10492_, new_n10493_, new_n10494_, new_n10495_,
    new_n10496_, new_n10497_, new_n10498_, new_n10499_, new_n10500_,
    new_n10501_, new_n10502_, new_n10503_, new_n10504_, new_n10505_,
    new_n10506_, new_n10507_, new_n10508_, new_n10509_, new_n10510_,
    new_n10511_, new_n10512_, new_n10513_, new_n10514_, new_n10515_,
    new_n10516_, new_n10517_, new_n10518_, new_n10519_, new_n10520_,
    new_n10521_, new_n10522_, new_n10523_, new_n10524_, new_n10525_,
    new_n10526_, new_n10527_, new_n10528_, new_n10529_, new_n10530_,
    new_n10531_, new_n10532_, new_n10533_, new_n10534_, new_n10535_,
    new_n10536_, new_n10537_, new_n10538_, new_n10539_, new_n10540_,
    new_n10541_, new_n10542_, new_n10543_, new_n10544_, new_n10545_,
    new_n10546_, new_n10547_, new_n10548_, new_n10549_, new_n10550_,
    new_n10551_, new_n10552_, new_n10553_, new_n10554_, new_n10555_,
    new_n10556_, new_n10557_, new_n10558_, new_n10559_, new_n10560_,
    new_n10561_, new_n10562_, new_n10563_, new_n10564_, new_n10565_,
    new_n10566_, new_n10567_, new_n10568_, new_n10569_, new_n10570_,
    new_n10571_, new_n10572_, new_n10573_, new_n10574_, new_n10575_,
    new_n10576_, new_n10577_, new_n10578_, new_n10579_, new_n10580_,
    new_n10581_, new_n10582_, new_n10583_, new_n10584_, new_n10585_,
    new_n10586_, new_n10587_, new_n10588_, new_n10589_, new_n10590_,
    new_n10591_, new_n10592_, new_n10593_, new_n10594_, new_n10595_,
    new_n10596_, new_n10597_, new_n10598_, new_n10599_, new_n10600_,
    new_n10601_, new_n10602_, new_n10603_, new_n10604_, new_n10605_,
    new_n10606_, new_n10607_, new_n10608_, new_n10609_, new_n10610_,
    new_n10611_, new_n10612_, new_n10613_, new_n10614_, new_n10615_,
    new_n10616_, new_n10617_, new_n10619_, new_n10620_, new_n10621_,
    new_n10623_, new_n10624_, new_n10625_, new_n10626_, new_n10627_,
    new_n10628_, new_n10629_, new_n10630_, new_n10631_, new_n10632_,
    new_n10633_, new_n10634_, new_n10635_, new_n10636_, new_n10637_,
    new_n10638_, new_n10639_, new_n10640_, new_n10641_, new_n10642_,
    new_n10643_, new_n10644_, new_n10645_, new_n10646_, new_n10647_,
    new_n10648_, new_n10649_, new_n10650_, new_n10651_, new_n10652_,
    new_n10653_, new_n10654_, new_n10655_, new_n10656_, new_n10657_,
    new_n10658_, new_n10660_, new_n10661_, new_n10662_, new_n10663_,
    new_n10664_, new_n10665_, new_n10666_, new_n10667_, new_n10668_,
    new_n10669_, new_n10670_, new_n10671_, new_n10672_, new_n10673_,
    new_n10674_, new_n10675_, new_n10676_, new_n10677_, new_n10678_,
    new_n10679_, new_n10680_, new_n10681_, new_n10682_, new_n10683_,
    new_n10684_, new_n10685_, new_n10686_, new_n10687_, new_n10688_,
    new_n10689_, new_n10690_, new_n10691_, new_n10692_, new_n10693_,
    new_n10694_, new_n10695_, new_n10696_, new_n10697_, new_n10698_,
    new_n10699_, new_n10700_, new_n10701_, new_n10702_, new_n10703_,
    new_n10704_, new_n10705_, new_n10706_, new_n10707_, new_n10708_,
    new_n10709_, new_n10710_, new_n10711_, new_n10712_, new_n10713_,
    new_n10714_, new_n10715_, new_n10716_, new_n10717_, new_n10718_,
    new_n10719_, new_n10720_, new_n10721_, new_n10722_, new_n10723_,
    new_n10724_, new_n10725_, new_n10726_, new_n10727_, new_n10728_,
    new_n10729_, new_n10730_, new_n10731_, new_n10732_, new_n10733_,
    new_n10734_, new_n10735_, new_n10736_, new_n10737_, new_n10738_,
    new_n10739_, new_n10740_, new_n10741_, new_n10742_, new_n10743_,
    new_n10744_, new_n10745_, new_n10746_, new_n10747_, new_n10748_,
    new_n10749_, new_n10750_, new_n10751_, new_n10752_, new_n10753_,
    new_n10754_, new_n10755_, new_n10756_, new_n10757_, new_n10758_,
    new_n10759_, new_n10760_, new_n10761_, new_n10762_, new_n10763_,
    new_n10764_, new_n10765_, new_n10766_, new_n10767_, new_n10768_,
    new_n10769_, new_n10770_, new_n10771_, new_n10772_, new_n10773_,
    new_n10774_, new_n10775_, new_n10776_, new_n10777_, new_n10778_,
    new_n10779_, new_n10780_, new_n10781_, new_n10782_, new_n10783_,
    new_n10784_, new_n10785_, new_n10786_, new_n10787_, new_n10788_,
    new_n10789_, new_n10790_, new_n10791_, new_n10792_, new_n10793_,
    new_n10794_, new_n10795_, new_n10796_, new_n10797_, new_n10798_,
    new_n10799_, new_n10800_, new_n10801_, new_n10802_, new_n10803_,
    new_n10804_, new_n10805_, new_n10806_, new_n10807_, new_n10808_,
    new_n10809_, new_n10810_, new_n10811_, new_n10812_, new_n10813_,
    new_n10814_, new_n10815_, new_n10816_, new_n10817_, new_n10818_,
    new_n10819_, new_n10820_, new_n10821_, new_n10822_, new_n10823_,
    new_n10824_, new_n10825_, new_n10826_, new_n10827_, new_n10828_,
    new_n10829_, new_n10830_, new_n10831_, new_n10832_, new_n10833_,
    new_n10834_, new_n10835_, new_n10836_, new_n10837_, new_n10838_,
    new_n10839_, new_n10840_, new_n10841_, new_n10842_, new_n10843_,
    new_n10844_, new_n10845_, new_n10846_, new_n10847_, new_n10848_,
    new_n10849_, new_n10850_, new_n10851_, new_n10852_, new_n10853_,
    new_n10854_, new_n10855_, new_n10856_, new_n10857_, new_n10858_,
    new_n10859_, new_n10860_, new_n10861_, new_n10862_, new_n10863_,
    new_n10864_, new_n10865_, new_n10866_, new_n10867_, new_n10868_,
    new_n10869_, new_n10870_, new_n10871_, new_n10872_, new_n10873_,
    new_n10874_, new_n10875_, new_n10876_, new_n10877_, new_n10878_,
    new_n10879_, new_n10880_, new_n10881_, new_n10882_, new_n10883_,
    new_n10884_, new_n10885_, new_n10886_, new_n10887_, new_n10888_,
    new_n10889_, new_n10890_, new_n10891_, new_n10892_, new_n10893_,
    new_n10894_, new_n10895_, new_n10896_, new_n10897_, new_n10898_,
    new_n10899_, new_n10900_, new_n10901_, new_n10902_, new_n10903_,
    new_n10904_, new_n10905_, new_n10906_, new_n10907_, new_n10908_,
    new_n10909_, new_n10910_, new_n10911_, new_n10912_, new_n10913_,
    new_n10914_, new_n10915_, new_n10916_, new_n10917_, new_n10918_,
    new_n10919_, new_n10920_, new_n10921_, new_n10922_, new_n10923_,
    new_n10924_, new_n10925_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10933_, new_n10934_,
    new_n10935_, new_n10936_, new_n10937_, new_n10938_, new_n10939_,
    new_n10940_, new_n10941_, new_n10942_, new_n10943_, new_n10944_,
    new_n10945_, new_n10946_, new_n10947_, new_n10948_, new_n10949_,
    new_n10950_, new_n10951_, new_n10952_, new_n10953_, new_n10954_,
    new_n10955_, new_n10956_, new_n10957_, new_n10958_, new_n10959_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10974_,
    new_n10975_, new_n10976_, new_n10977_, new_n10978_, new_n10979_,
    new_n10980_, new_n10981_, new_n10982_, new_n10983_, new_n10984_,
    new_n10985_, new_n10986_, new_n10987_, new_n10988_, new_n10989_,
    new_n10990_, new_n10991_, new_n10992_, new_n10993_, new_n10994_,
    new_n10995_, new_n10996_, new_n10997_, new_n10998_, new_n10999_,
    new_n11000_, new_n11001_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11050_, new_n11051_, new_n11052_, new_n11053_, new_n11054_,
    new_n11055_, new_n11056_, new_n11057_, new_n11058_, new_n11059_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11073_, new_n11074_,
    new_n11075_, new_n11076_, new_n11077_, new_n11078_, new_n11079_,
    new_n11080_, new_n11081_, new_n11082_, new_n11083_, new_n11084_,
    new_n11085_, new_n11086_, new_n11087_, new_n11088_, new_n11089_,
    new_n11090_, new_n11091_, new_n11092_, new_n11093_, new_n11094_,
    new_n11095_, new_n11096_, new_n11097_, new_n11098_, new_n11099_,
    new_n11100_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11106_, new_n11108_, new_n11109_, new_n11110_,
    new_n11111_, new_n11112_, new_n11113_, new_n11114_, new_n11115_,
    new_n11116_, new_n11117_, new_n11118_, new_n11119_, new_n11120_,
    new_n11121_, new_n11122_, new_n11123_, new_n11124_, new_n11125_,
    new_n11126_, new_n11127_, new_n11128_, new_n11129_, new_n11130_,
    new_n11131_, new_n11132_, new_n11133_, new_n11134_, new_n11135_,
    new_n11136_, new_n11137_, new_n11138_, new_n11139_, new_n11140_,
    new_n11141_, new_n11142_, new_n11143_, new_n11144_, new_n11145_,
    new_n11146_, new_n11147_, new_n11148_, new_n11149_, new_n11150_,
    new_n11151_, new_n11152_, new_n11153_, new_n11154_, new_n11155_,
    new_n11156_, new_n11157_, new_n11158_, new_n11159_, new_n11160_,
    new_n11161_, new_n11162_, new_n11163_, new_n11164_, new_n11165_,
    new_n11167_, new_n11168_, new_n11169_, new_n11170_, new_n11171_,
    new_n11172_, new_n11173_, new_n11174_, new_n11175_, new_n11176_,
    new_n11177_, new_n11178_, new_n11179_, new_n11180_, new_n11181_,
    new_n11183_, new_n11184_, new_n11185_, new_n11186_, new_n11187_,
    new_n11188_, new_n11189_, new_n11190_, new_n11191_, new_n11192_,
    new_n11193_, new_n11194_, new_n11195_, new_n11196_, new_n11197_,
    new_n11198_, new_n11199_, new_n11200_, new_n11201_, new_n11202_,
    new_n11203_, new_n11204_, new_n11205_, new_n11206_, new_n11207_,
    new_n11208_, new_n11209_, new_n11210_, new_n11211_, new_n11212_,
    new_n11213_, new_n11214_, new_n11215_, new_n11216_, new_n11217_,
    new_n11218_, new_n11219_, new_n11220_, new_n11221_, new_n11222_,
    new_n11223_, new_n11224_, new_n11225_, new_n11226_, new_n11227_,
    new_n11228_, new_n11229_, new_n11230_, new_n11231_, new_n11232_,
    new_n11233_, new_n11234_, new_n11235_, new_n11236_, new_n11237_,
    new_n11238_, new_n11239_, new_n11240_, new_n11241_, new_n11242_,
    new_n11243_, new_n11244_, new_n11245_, new_n11246_, new_n11247_,
    new_n11248_, new_n11249_, new_n11250_, new_n11251_, new_n11252_,
    new_n11253_, new_n11254_, new_n11255_, new_n11256_, new_n11257_,
    new_n11258_, new_n11259_, new_n11260_, new_n11261_, new_n11262_,
    new_n11263_, new_n11264_, new_n11265_, new_n11266_, new_n11267_,
    new_n11268_, new_n11269_, new_n11271_, new_n11272_, new_n11273_,
    new_n11274_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11286_, new_n11287_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11298_, new_n11299_,
    new_n11300_, new_n11301_, new_n11302_, new_n11303_, new_n11304_,
    new_n11305_, new_n11306_, new_n11307_, new_n11308_, new_n11309_,
    new_n11310_, new_n11311_, new_n11312_, new_n11313_, new_n11314_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11324_,
    new_n11325_, new_n11326_, new_n11327_, new_n11328_, new_n11329_,
    new_n11330_, new_n11331_, new_n11332_, new_n11333_, new_n11334_,
    new_n11335_, new_n11336_, new_n11337_, new_n11338_, new_n11339_,
    new_n11340_, new_n11341_, new_n11342_, new_n11343_, new_n11344_,
    new_n11345_, new_n11346_, new_n11347_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11352_, new_n11353_, new_n11354_,
    new_n11355_, new_n11356_, new_n11357_, new_n11358_, new_n11359_,
    new_n11360_, new_n11361_, new_n11362_, new_n11363_, new_n11364_,
    new_n11365_, new_n11366_, new_n11367_, new_n11368_, new_n11369_,
    new_n11370_, new_n11371_, new_n11372_, new_n11373_, new_n11374_,
    new_n11375_, new_n11376_, new_n11377_, new_n11378_, new_n11379_,
    new_n11380_, new_n11381_, new_n11382_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11409_, new_n11410_,
    new_n11411_, new_n11412_, new_n11413_, new_n11414_, new_n11415_,
    new_n11416_, new_n11417_, new_n11418_, new_n11419_, new_n11420_,
    new_n11421_, new_n11422_, new_n11423_, new_n11424_, new_n11425_,
    new_n11426_, new_n11427_, new_n11428_, new_n11429_, new_n11430_,
    new_n11431_, new_n11432_, new_n11433_, new_n11434_, new_n11435_,
    new_n11436_, new_n11437_, new_n11438_, new_n11439_, new_n11440_,
    new_n11441_, new_n11442_, new_n11443_, new_n11444_, new_n11445_,
    new_n11446_, new_n11448_, new_n11449_, new_n11450_, new_n11451_,
    new_n11452_, new_n11453_, new_n11454_, new_n11455_, new_n11456_,
    new_n11457_, new_n11458_, new_n11459_, new_n11460_, new_n11461_,
    new_n11462_, new_n11463_, new_n11464_, new_n11465_, new_n11466_,
    new_n11467_, new_n11468_, new_n11469_, new_n11470_, new_n11471_,
    new_n11472_, new_n11473_, new_n11474_, new_n11475_, new_n11476_,
    new_n11477_, new_n11478_, new_n11479_, new_n11480_, new_n11481_,
    new_n11482_, new_n11483_, new_n11484_, new_n11485_, new_n11486_,
    new_n11487_, new_n11488_, new_n11489_, new_n11490_, new_n11491_,
    new_n11492_, new_n11493_, new_n11494_, new_n11495_, new_n11496_,
    new_n11497_, new_n11498_, new_n11499_, new_n11500_, new_n11501_,
    new_n11502_, new_n11503_, new_n11504_, new_n11505_, new_n11506_,
    new_n11507_, new_n11508_, new_n11509_, new_n11510_, new_n11511_,
    new_n11512_, new_n11513_, new_n11514_, new_n11515_, new_n11516_,
    new_n11517_, new_n11518_, new_n11519_, new_n11520_, new_n11521_,
    new_n11522_, new_n11524_, new_n11525_, new_n11526_, new_n11527_,
    new_n11528_, new_n11529_, new_n11530_, new_n11531_, new_n11532_,
    new_n11533_, new_n11534_, new_n11535_, new_n11536_, new_n11537_,
    new_n11538_, new_n11539_, new_n11540_, new_n11541_, new_n11542_,
    new_n11543_, new_n11544_, new_n11545_, new_n11546_, new_n11547_,
    new_n11548_, new_n11549_, new_n11550_, new_n11551_, new_n11552_,
    new_n11553_, new_n11554_, new_n11555_, new_n11556_, new_n11557_,
    new_n11558_, new_n11559_, new_n11560_, new_n11561_, new_n11562_,
    new_n11563_, new_n11564_, new_n11565_, new_n11566_, new_n11567_,
    new_n11568_, new_n11569_, new_n11570_, new_n11571_, new_n11572_,
    new_n11573_, new_n11574_, new_n11575_, new_n11576_, new_n11577_,
    new_n11578_, new_n11579_, new_n11580_, new_n11581_, new_n11582_,
    new_n11583_, new_n11584_, new_n11585_, new_n11586_, new_n11587_,
    new_n11588_, new_n11589_, new_n11590_, new_n11591_, new_n11592_,
    new_n11593_, new_n11594_, new_n11595_, new_n11596_, new_n11597_,
    new_n11598_, new_n11599_, new_n11600_, new_n11601_, new_n11603_,
    new_n11604_, new_n11605_, new_n11606_, new_n11607_, new_n11608_,
    new_n11609_, new_n11610_, new_n11611_, new_n11612_, new_n11613_,
    new_n11614_, new_n11615_, new_n11616_, new_n11617_, new_n11618_,
    new_n11619_, new_n11620_, new_n11621_, new_n11622_, new_n11623_,
    new_n11624_, new_n11625_, new_n11626_, new_n11627_, new_n11628_,
    new_n11629_, new_n11630_, new_n11631_, new_n11632_, new_n11633_,
    new_n11634_, new_n11635_, new_n11636_, new_n11637_, new_n11638_,
    new_n11639_, new_n11640_, new_n11641_, new_n11642_, new_n11643_,
    new_n11644_, new_n11645_, new_n11646_, new_n11647_, new_n11648_,
    new_n11649_, new_n11650_, new_n11651_, new_n11652_, new_n11653_,
    new_n11654_, new_n11655_, new_n11656_, new_n11658_, new_n11659_,
    new_n11660_, new_n11661_, new_n11662_, new_n11663_, new_n11664_,
    new_n11666_, new_n11667_, new_n11668_, new_n11669_, new_n11670_,
    new_n11671_, new_n11672_, new_n11673_, new_n11674_, new_n11675_,
    new_n11676_, new_n11677_, new_n11678_, new_n11679_, new_n11680_,
    new_n11681_, new_n11682_, new_n11683_, new_n11684_, new_n11685_,
    new_n11686_, new_n11687_, new_n11688_, new_n11689_, new_n11690_,
    new_n11691_, new_n11692_, new_n11693_, new_n11694_, new_n11695_,
    new_n11696_, new_n11697_, new_n11698_, new_n11699_, new_n11700_,
    new_n11701_, new_n11702_, new_n11703_, new_n11704_, new_n11705_,
    new_n11706_, new_n11707_, new_n11708_, new_n11709_, new_n11710_,
    new_n11711_, new_n11712_, new_n11713_, new_n11714_, new_n11715_,
    new_n11716_, new_n11717_, new_n11718_, new_n11719_, new_n11720_,
    new_n11721_, new_n11722_, new_n11723_, new_n11724_, new_n11725_,
    new_n11726_, new_n11727_, new_n11728_, new_n11729_, new_n11731_,
    new_n11732_, new_n11733_, new_n11734_, new_n11735_, new_n11736_,
    new_n11737_, new_n11738_, new_n11739_, new_n11740_, new_n11741_,
    new_n11742_, new_n11743_, new_n11744_, new_n11745_, new_n11746_,
    new_n11747_, new_n11748_, new_n11749_, new_n11750_, new_n11751_,
    new_n11752_, new_n11753_, new_n11754_, new_n11755_, new_n11756_,
    new_n11757_, new_n11758_, new_n11759_, new_n11760_, new_n11762_,
    new_n11763_, new_n11764_, new_n11765_, new_n11766_, new_n11767_,
    new_n11768_, new_n11769_, new_n11770_, new_n11771_, new_n11772_,
    new_n11773_, new_n11774_, new_n11775_, new_n11776_, new_n11777_,
    new_n11778_, new_n11779_, new_n11780_, new_n11781_, new_n11782_,
    new_n11783_, new_n11784_, new_n11785_, new_n11786_, new_n11787_,
    new_n11788_, new_n11789_, new_n11790_, new_n11791_, new_n11792_,
    new_n11793_, new_n11794_, new_n11795_, new_n11796_, new_n11797_,
    new_n11798_, new_n11799_, new_n11800_, new_n11801_, new_n11802_,
    new_n11803_, new_n11805_, new_n11806_, new_n11807_, new_n11808_,
    new_n11809_, new_n11810_, new_n11811_, new_n11812_, new_n11813_,
    new_n11814_, new_n11815_, new_n11816_, new_n11817_, new_n11818_,
    new_n11819_, new_n11820_, new_n11821_, new_n11822_, new_n11823_,
    new_n11824_, new_n11825_, new_n11826_, new_n11827_, new_n11828_,
    new_n11829_, new_n11830_, new_n11831_, new_n11832_, new_n11833_,
    new_n11834_, new_n11835_, new_n11836_, new_n11837_, new_n11838_,
    new_n11839_, new_n11840_, new_n11841_, new_n11842_, new_n11843_,
    new_n11844_, new_n11845_, new_n11846_, new_n11847_, new_n11848_,
    new_n11849_, new_n11850_, new_n11851_, new_n11852_, new_n11853_,
    new_n11854_, new_n11855_, new_n11856_, new_n11857_, new_n11858_,
    new_n11859_, new_n11860_, new_n11861_, new_n11862_, new_n11863_,
    new_n11864_, new_n11865_, new_n11866_, new_n11867_, new_n11868_,
    new_n11869_, new_n11870_, new_n11871_, new_n11872_, new_n11873_,
    new_n11874_, new_n11875_, new_n11876_, new_n11877_, new_n11878_,
    new_n11879_, new_n11880_, new_n11881_, new_n11882_, new_n11883_,
    new_n11884_, new_n11885_, new_n11886_, new_n11887_, new_n11888_,
    new_n11889_, new_n11890_, new_n11891_, new_n11892_, new_n11893_,
    new_n11894_, new_n11895_, new_n11896_, new_n11897_, new_n11898_,
    new_n11899_, new_n11900_, new_n11901_, new_n11902_, new_n11903_,
    new_n11904_, new_n11905_, new_n11906_, new_n11907_, new_n11908_,
    new_n11909_, new_n11910_, new_n11911_, new_n11912_, new_n11913_,
    new_n11914_, new_n11915_, new_n11916_, new_n11917_, new_n11918_,
    new_n11919_, new_n11920_, new_n11921_, new_n11922_, new_n11923_,
    new_n11924_, new_n11925_, new_n11926_, new_n11927_, new_n11928_,
    new_n11929_, new_n11930_, new_n11931_, new_n11932_, new_n11933_,
    new_n11934_, new_n11935_, new_n11936_, new_n11937_, new_n11938_,
    new_n11939_, new_n11940_, new_n11941_, new_n11942_, new_n11943_,
    new_n11944_, new_n11945_, new_n11946_, new_n11947_, new_n11948_,
    new_n11949_, new_n11950_, new_n11951_, new_n11952_, new_n11953_,
    new_n11954_, new_n11955_, new_n11956_, new_n11957_, new_n11958_,
    new_n11959_, new_n11960_, new_n11961_, new_n11962_, new_n11963_,
    new_n11964_, new_n11965_, new_n11966_, new_n11967_, new_n11968_,
    new_n11969_, new_n11970_, new_n11971_, new_n11972_, new_n11973_,
    new_n11974_, new_n11975_, new_n11976_, new_n11977_, new_n11978_,
    new_n11979_, new_n11980_, new_n11981_, new_n11982_, new_n11983_,
    new_n11984_, new_n11985_, new_n11986_, new_n11987_, new_n11988_,
    new_n11989_, new_n11990_, new_n11991_, new_n11992_, new_n11993_,
    new_n11994_, new_n11995_, new_n11996_, new_n11997_, new_n11998_,
    new_n11999_, new_n12000_, new_n12001_, new_n12002_, new_n12003_,
    new_n12004_, new_n12005_, new_n12006_, new_n12007_, new_n12008_,
    new_n12009_, new_n12010_, new_n12011_, new_n12012_, new_n12013_,
    new_n12014_, new_n12015_, new_n12016_, new_n12017_, new_n12018_,
    new_n12019_, new_n12020_, new_n12021_, new_n12022_, new_n12023_,
    new_n12024_, new_n12025_, new_n12026_, new_n12027_, new_n12028_,
    new_n12029_, new_n12030_, new_n12031_, new_n12032_, new_n12033_,
    new_n12034_, new_n12035_, new_n12036_, new_n12037_, new_n12038_,
    new_n12039_, new_n12040_, new_n12041_, new_n12042_, new_n12043_,
    new_n12044_, new_n12045_, new_n12046_, new_n12047_, new_n12048_,
    new_n12049_, new_n12050_, new_n12051_, new_n12052_, new_n12053_,
    new_n12054_, new_n12055_, new_n12056_, new_n12057_, new_n12058_,
    new_n12059_, new_n12060_, new_n12061_, new_n12062_, new_n12063_,
    new_n12064_, new_n12065_, new_n12066_, new_n12067_, new_n12068_,
    new_n12069_, new_n12070_, new_n12071_, new_n12072_, new_n12073_,
    new_n12074_, new_n12075_, new_n12076_, new_n12077_, new_n12078_,
    new_n12079_, new_n12080_, new_n12081_, new_n12082_, new_n12083_,
    new_n12084_, new_n12085_, new_n12086_, new_n12087_, new_n12088_,
    new_n12089_, new_n12090_, new_n12091_, new_n12092_, new_n12093_,
    new_n12094_, new_n12095_, new_n12096_, new_n12097_, new_n12098_,
    new_n12099_, new_n12100_, new_n12101_, new_n12102_, new_n12103_,
    new_n12104_, new_n12105_, new_n12106_, new_n12107_, new_n12108_,
    new_n12109_, new_n12110_, new_n12111_, new_n12112_, new_n12113_,
    new_n12114_, new_n12115_, new_n12116_, new_n12117_, new_n12118_,
    new_n12119_, new_n12120_, new_n12121_, new_n12122_, new_n12123_,
    new_n12124_, new_n12125_, new_n12126_, new_n12127_, new_n12128_,
    new_n12129_, new_n12130_, new_n12131_, new_n12132_, new_n12133_,
    new_n12134_, new_n12135_, new_n12136_, new_n12137_, new_n12138_,
    new_n12139_, new_n12140_, new_n12141_, new_n12142_, new_n12143_,
    new_n12144_, new_n12145_, new_n12146_, new_n12147_, new_n12148_,
    new_n12149_, new_n12150_, new_n12151_, new_n12152_, new_n12153_,
    new_n12154_, new_n12155_, new_n12156_, new_n12157_, new_n12158_,
    new_n12159_, new_n12160_, new_n12161_, new_n12162_, new_n12163_,
    new_n12164_, new_n12165_, new_n12166_, new_n12167_, new_n12168_,
    new_n12169_, new_n12170_, new_n12171_, new_n12172_, new_n12173_,
    new_n12174_, new_n12175_, new_n12176_, new_n12177_, new_n12178_,
    new_n12179_, new_n12180_, new_n12181_, new_n12182_, new_n12183_,
    new_n12184_, new_n12185_, new_n12186_, new_n12187_, new_n12188_,
    new_n12189_, new_n12190_, new_n12191_, new_n12192_, new_n12193_,
    new_n12194_, new_n12195_, new_n12196_, new_n12197_, new_n12198_,
    new_n12199_, new_n12200_, new_n12201_, new_n12202_, new_n12203_,
    new_n12204_, new_n12205_, new_n12206_, new_n12207_, new_n12208_,
    new_n12209_, new_n12210_, new_n12211_, new_n12212_, new_n12213_,
    new_n12214_, new_n12215_, new_n12216_, new_n12217_, new_n12218_,
    new_n12219_, new_n12220_, new_n12221_, new_n12222_, new_n12223_,
    new_n12224_, new_n12225_, new_n12226_, new_n12227_, new_n12228_,
    new_n12229_, new_n12230_, new_n12231_, new_n12232_, new_n12233_,
    new_n12234_, new_n12235_, new_n12236_, new_n12237_, new_n12238_,
    new_n12239_, new_n12240_, new_n12241_, new_n12242_, new_n12243_,
    new_n12244_, new_n12245_, new_n12246_, new_n12247_, new_n12248_,
    new_n12249_, new_n12250_, new_n12251_, new_n12252_, new_n12253_,
    new_n12254_, new_n12255_, new_n12256_, new_n12257_, new_n12258_,
    new_n12259_, new_n12260_, new_n12261_, new_n12262_, new_n12263_,
    new_n12264_, new_n12265_, new_n12266_, new_n12267_, new_n12268_,
    new_n12269_, new_n12270_, new_n12271_, new_n12272_, new_n12273_,
    new_n12274_, new_n12275_, new_n12276_, new_n12277_, new_n12278_,
    new_n12279_, new_n12280_, new_n12281_, new_n12282_, new_n12283_,
    new_n12284_, new_n12285_, new_n12286_, new_n12287_, new_n12288_,
    new_n12289_, new_n12290_, new_n12291_, new_n12292_, new_n12293_,
    new_n12294_, new_n12295_, new_n12296_, new_n12297_, new_n12298_,
    new_n12299_, new_n12300_, new_n12301_, new_n12302_, new_n12303_,
    new_n12304_, new_n12305_, new_n12306_, new_n12307_, new_n12308_,
    new_n12309_, new_n12310_, new_n12311_, new_n12312_, new_n12313_,
    new_n12314_, new_n12315_, new_n12316_, new_n12317_, new_n12318_,
    new_n12319_, new_n12320_, new_n12321_, new_n12322_, new_n12323_,
    new_n12324_, new_n12325_, new_n12326_, new_n12327_, new_n12328_,
    new_n12329_, new_n12330_, new_n12331_, new_n12332_, new_n12333_,
    new_n12334_, new_n12335_, new_n12336_, new_n12337_, new_n12338_,
    new_n12339_, new_n12340_, new_n12341_, new_n12342_, new_n12343_,
    new_n12344_, new_n12345_, new_n12346_, new_n12347_, new_n12348_,
    new_n12349_, new_n12350_, new_n12351_, new_n12352_, new_n12353_,
    new_n12354_, new_n12355_, new_n12356_, new_n12357_, new_n12358_,
    new_n12359_, new_n12360_, new_n12361_, new_n12362_, new_n12363_,
    new_n12364_, new_n12365_, new_n12366_, new_n12367_, new_n12368_,
    new_n12369_, new_n12370_, new_n12371_, new_n12372_, new_n12373_,
    new_n12374_, new_n12375_, new_n12376_, new_n12377_, new_n12378_,
    new_n12379_, new_n12380_, new_n12381_, new_n12382_, new_n12383_,
    new_n12384_, new_n12385_, new_n12386_, new_n12387_, new_n12388_,
    new_n12389_, new_n12390_, new_n12391_, new_n12392_, new_n12393_,
    new_n12394_, new_n12395_, new_n12396_, new_n12397_, new_n12398_,
    new_n12399_, new_n12400_, new_n12401_, new_n12402_, new_n12403_,
    new_n12404_, new_n12405_, new_n12406_, new_n12407_, new_n12408_,
    new_n12409_, new_n12410_, new_n12411_, new_n12412_, new_n12413_,
    new_n12414_, new_n12415_, new_n12416_, new_n12417_, new_n12418_,
    new_n12419_, new_n12420_, new_n12421_, new_n12422_, new_n12423_,
    new_n12424_, new_n12425_, new_n12426_, new_n12427_, new_n12428_,
    new_n12429_, new_n12430_, new_n12431_, new_n12432_, new_n12433_,
    new_n12434_, new_n12435_, new_n12436_, new_n12437_, new_n12438_,
    new_n12439_, new_n12440_, new_n12441_, new_n12442_, new_n12443_,
    new_n12444_, new_n12445_, new_n12446_, new_n12447_, new_n12448_,
    new_n12449_, new_n12450_, new_n12451_, new_n12452_, new_n12453_,
    new_n12454_, new_n12455_, new_n12456_, new_n12457_, new_n12458_,
    new_n12459_, new_n12460_, new_n12461_, new_n12462_, new_n12463_,
    new_n12464_, new_n12465_, new_n12466_, new_n12467_, new_n12468_,
    new_n12469_, new_n12470_, new_n12471_, new_n12472_, new_n12473_,
    new_n12474_, new_n12475_, new_n12476_, new_n12477_, new_n12478_,
    new_n12479_, new_n12480_, new_n12481_, new_n12482_, new_n12483_,
    new_n12484_, new_n12485_, new_n12486_, new_n12487_, new_n12488_,
    new_n12489_, new_n12490_, new_n12491_, new_n12492_, new_n12493_,
    new_n12494_, new_n12495_, new_n12496_, new_n12497_, new_n12498_,
    new_n12499_, new_n12500_, new_n12501_, new_n12502_, new_n12503_,
    new_n12504_, new_n12505_, new_n12506_, new_n12507_, new_n12508_,
    new_n12509_, new_n12510_, new_n12511_, new_n12512_, new_n12513_,
    new_n12514_, new_n12515_, new_n12516_, new_n12517_, new_n12518_,
    new_n12519_, new_n12520_, new_n12521_, new_n12522_, new_n12523_,
    new_n12524_, new_n12525_, new_n12526_, new_n12527_, new_n12528_,
    new_n12529_, new_n12530_, new_n12531_, new_n12532_, new_n12533_,
    new_n12534_, new_n12535_, new_n12536_, new_n12537_, new_n12538_,
    new_n12539_, new_n12540_, new_n12541_, new_n12542_, new_n12543_,
    new_n12544_, new_n12545_, new_n12546_, new_n12547_, new_n12548_,
    new_n12549_, new_n12550_, new_n12551_, new_n12552_, new_n12553_,
    new_n12554_, new_n12555_, new_n12556_, new_n12557_, new_n12558_,
    new_n12559_, new_n12560_, new_n12561_, new_n12562_, new_n12563_,
    new_n12564_, new_n12565_, new_n12566_, new_n12567_, new_n12568_,
    new_n12569_, new_n12570_, new_n12571_, new_n12572_, new_n12573_,
    new_n12574_, new_n12575_, new_n12576_, new_n12577_, new_n12578_,
    new_n12579_, new_n12580_, new_n12581_, new_n12582_, new_n12583_,
    new_n12584_, new_n12585_, new_n12586_, new_n12587_, new_n12588_,
    new_n12589_, new_n12590_, new_n12591_, new_n12592_, new_n12593_,
    new_n12594_, new_n12595_, new_n12596_, new_n12597_, new_n12598_,
    new_n12599_, new_n12600_, new_n12601_, new_n12602_, new_n12603_,
    new_n12604_, new_n12605_, new_n12606_, new_n12607_, new_n12608_,
    new_n12609_, new_n12610_, new_n12611_, new_n12612_, new_n12613_,
    new_n12614_, new_n12615_, new_n12616_, new_n12617_, new_n12618_,
    new_n12619_, new_n12620_, new_n12621_, new_n12622_, new_n12623_,
    new_n12624_, new_n12625_, new_n12626_, new_n12627_, new_n12628_,
    new_n12629_, new_n12630_, new_n12631_, new_n12632_, new_n12633_,
    new_n12634_, new_n12635_, new_n12636_, new_n12637_, new_n12638_,
    new_n12639_, new_n12640_, new_n12641_, new_n12642_, new_n12643_,
    new_n12644_, new_n12645_, new_n12646_, new_n12647_, new_n12648_,
    new_n12649_, new_n12650_, new_n12651_, new_n12652_, new_n12653_,
    new_n12654_, new_n12655_, new_n12656_, new_n12657_, new_n12658_,
    new_n12659_, new_n12660_, new_n12661_, new_n12662_, new_n12663_,
    new_n12664_, new_n12665_, new_n12666_, new_n12667_, new_n12668_,
    new_n12669_, new_n12670_, new_n12671_, new_n12672_, new_n12673_,
    new_n12674_, new_n12675_, new_n12676_, new_n12677_, new_n12678_,
    new_n12679_, new_n12680_, new_n12681_, new_n12682_, new_n12683_,
    new_n12684_, new_n12685_, new_n12686_, new_n12687_, new_n12688_,
    new_n12689_, new_n12690_, new_n12691_, new_n12692_, new_n12693_,
    new_n12694_, new_n12695_, new_n12696_, new_n12697_, new_n12698_,
    new_n12699_, new_n12700_, new_n12701_, new_n12702_, new_n12703_,
    new_n12704_, new_n12705_, new_n12706_, new_n12707_, new_n12708_,
    new_n12709_, new_n12710_, new_n12711_, new_n12712_, new_n12713_,
    new_n12714_, new_n12715_, new_n12716_, new_n12717_, new_n12718_,
    new_n12719_, new_n12720_, new_n12721_, new_n12722_, new_n12723_,
    new_n12724_, new_n12725_, new_n12726_, new_n12727_, new_n12728_,
    new_n12729_, new_n12730_, new_n12731_, new_n12732_, new_n12733_,
    new_n12734_, new_n12735_, new_n12736_, new_n12737_, new_n12738_,
    new_n12739_, new_n12740_, new_n12741_, new_n12742_, new_n12743_,
    new_n12744_, new_n12745_, new_n12746_, new_n12747_, new_n12748_,
    new_n12749_, new_n12750_, new_n12751_, new_n12752_, new_n12753_,
    new_n12754_, new_n12755_, new_n12756_, new_n12757_, new_n12758_,
    new_n12759_, new_n12760_, new_n12761_, new_n12762_, new_n12763_,
    new_n12764_, new_n12765_, new_n12766_, new_n12767_, new_n12768_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13086_, new_n13087_, new_n13088_, new_n13089_, new_n13090_,
    new_n13091_, new_n13092_, new_n13093_, new_n13094_, new_n13095_,
    new_n13096_, new_n13097_, new_n13098_, new_n13099_, new_n13100_,
    new_n13101_, new_n13102_, new_n13103_, new_n13104_, new_n13105_,
    new_n13106_, new_n13107_, new_n13108_, new_n13109_, new_n13110_,
    new_n13111_, new_n13112_, new_n13113_, new_n13114_, new_n13115_,
    new_n13116_, new_n13117_, new_n13118_, new_n13119_, new_n13120_,
    new_n13121_, new_n13122_, new_n13123_, new_n13124_, new_n13125_,
    new_n13126_, new_n13127_, new_n13128_, new_n13129_, new_n13130_,
    new_n13131_, new_n13132_, new_n13133_, new_n13134_, new_n13135_,
    new_n13136_, new_n13137_, new_n13138_, new_n13139_, new_n13140_,
    new_n13141_, new_n13142_, new_n13143_, new_n13144_, new_n13145_,
    new_n13146_, new_n13147_, new_n13148_, new_n13149_, new_n13150_,
    new_n13151_, new_n13152_, new_n13153_, new_n13154_, new_n13155_,
    new_n13156_, new_n13157_, new_n13158_, new_n13159_, new_n13160_,
    new_n13161_, new_n13162_, new_n13163_, new_n13164_, new_n13165_,
    new_n13166_, new_n13167_, new_n13168_, new_n13169_, new_n13170_,
    new_n13171_, new_n13172_, new_n13173_, new_n13174_, new_n13175_,
    new_n13176_, new_n13177_, new_n13178_, new_n13179_, new_n13180_,
    new_n13181_, new_n13182_, new_n13183_, new_n13184_, new_n13185_,
    new_n13186_, new_n13187_, new_n13188_, new_n13189_, new_n13190_,
    new_n13191_, new_n13192_, new_n13193_, new_n13194_, new_n13195_,
    new_n13196_, new_n13197_, new_n13198_, new_n13199_, new_n13200_,
    new_n13201_, new_n13202_, new_n13203_, new_n13204_, new_n13205_,
    new_n13206_, new_n13207_, new_n13208_, new_n13209_, new_n13210_,
    new_n13211_, new_n13212_, new_n13213_, new_n13214_, new_n13215_,
    new_n13216_, new_n13217_, new_n13218_, new_n13219_, new_n13220_,
    new_n13221_, new_n13222_, new_n13223_, new_n13224_, new_n13225_,
    new_n13226_, new_n13227_, new_n13228_, new_n13229_, new_n13230_,
    new_n13231_, new_n13232_, new_n13233_, new_n13234_, new_n13235_,
    new_n13236_, new_n13237_, new_n13238_, new_n13239_, new_n13240_,
    new_n13241_, new_n13242_, new_n13243_, new_n13244_, new_n13245_,
    new_n13246_, new_n13247_, new_n13248_, new_n13249_, new_n13250_,
    new_n13251_, new_n13252_, new_n13253_, new_n13254_, new_n13255_,
    new_n13256_, new_n13257_, new_n13258_, new_n13259_, new_n13260_,
    new_n13261_, new_n13262_, new_n13263_, new_n13264_, new_n13265_,
    new_n13266_, new_n13267_, new_n13268_, new_n13269_, new_n13270_,
    new_n13271_, new_n13272_, new_n13273_, new_n13274_, new_n13275_,
    new_n13276_, new_n13277_, new_n13278_, new_n13279_, new_n13280_,
    new_n13281_, new_n13282_, new_n13283_, new_n13284_, new_n13285_,
    new_n13286_, new_n13287_, new_n13288_, new_n13289_, new_n13290_,
    new_n13291_, new_n13292_, new_n13293_, new_n13294_, new_n13295_,
    new_n13296_, new_n13297_, new_n13298_, new_n13299_, new_n13300_,
    new_n13301_, new_n13302_, new_n13303_, new_n13304_, new_n13305_,
    new_n13306_, new_n13307_, new_n13308_, new_n13309_, new_n13310_,
    new_n13311_, new_n13312_, new_n13313_, new_n13314_, new_n13315_,
    new_n13316_, new_n13317_, new_n13318_, new_n13319_, new_n13320_,
    new_n13321_, new_n13322_, new_n13323_, new_n13324_, new_n13325_,
    new_n13326_, new_n13327_, new_n13328_, new_n13329_, new_n13330_,
    new_n13331_, new_n13332_, new_n13333_, new_n13334_, new_n13335_,
    new_n13336_, new_n13337_, new_n13338_, new_n13339_, new_n13340_,
    new_n13341_, new_n13342_, new_n13343_, new_n13344_, new_n13345_,
    new_n13346_, new_n13347_, new_n13348_, new_n13349_, new_n13350_,
    new_n13351_, new_n13352_, new_n13353_, new_n13354_, new_n13355_,
    new_n13356_, new_n13357_, new_n13358_, new_n13359_, new_n13360_,
    new_n13361_, new_n13362_, new_n13363_, new_n13364_, new_n13365_,
    new_n13366_, new_n13367_, new_n13368_, new_n13369_, new_n13370_,
    new_n13371_, new_n13372_, new_n13373_, new_n13374_, new_n13375_,
    new_n13376_, new_n13377_, new_n13378_, new_n13379_, new_n13380_,
    new_n13381_, new_n13382_, new_n13383_, new_n13384_, new_n13385_,
    new_n13386_, new_n13387_, new_n13388_, new_n13389_, new_n13390_,
    new_n13391_, new_n13392_, new_n13393_, new_n13394_, new_n13395_,
    new_n13396_, new_n13397_, new_n13398_, new_n13399_, new_n13400_,
    new_n13401_, new_n13402_, new_n13403_, new_n13404_, new_n13405_,
    new_n13406_, new_n13407_, new_n13408_, new_n13409_, new_n13410_,
    new_n13411_, new_n13412_, new_n13413_, new_n13414_, new_n13415_,
    new_n13416_, new_n13417_, new_n13418_, new_n13419_, new_n13420_,
    new_n13421_, new_n13422_, new_n13423_, new_n13424_, new_n13425_,
    new_n13426_, new_n13427_, new_n13428_, new_n13429_, new_n13430_,
    new_n13431_, new_n13432_, new_n13433_, new_n13434_, new_n13435_,
    new_n13436_, new_n13437_, new_n13438_, new_n13439_, new_n13440_,
    new_n13441_, new_n13442_, new_n13443_, new_n13444_, new_n13445_,
    new_n13446_, new_n13447_, new_n13448_, new_n13449_, new_n13450_,
    new_n13451_, new_n13452_, new_n13453_, new_n13454_, new_n13455_,
    new_n13456_, new_n13457_, new_n13458_, new_n13459_, new_n13460_,
    new_n13461_, new_n13462_, new_n13463_, new_n13464_, new_n13465_,
    new_n13466_, new_n13467_, new_n13468_, new_n13469_, new_n13470_,
    new_n13471_, new_n13472_, new_n13473_, new_n13474_, new_n13475_,
    new_n13476_, new_n13477_, new_n13478_, new_n13479_, new_n13480_,
    new_n13481_, new_n13482_, new_n13483_, new_n13484_, new_n13485_,
    new_n13486_, new_n13487_, new_n13488_, new_n13489_, new_n13490_,
    new_n13491_, new_n13492_, new_n13493_, new_n13494_, new_n13495_,
    new_n13496_, new_n13497_, new_n13498_, new_n13499_, new_n13500_,
    new_n13501_, new_n13502_, new_n13503_, new_n13504_, new_n13505_,
    new_n13506_, new_n13507_, new_n13508_, new_n13509_, new_n13510_,
    new_n13511_, new_n13512_, new_n13513_, new_n13514_, new_n13515_,
    new_n13516_, new_n13517_, new_n13518_, new_n13519_, new_n13520_,
    new_n13521_, new_n13522_, new_n13523_, new_n13524_, new_n13525_,
    new_n13526_, new_n13527_, new_n13528_, new_n13529_, new_n13530_,
    new_n13531_, new_n13532_, new_n13533_, new_n13534_, new_n13535_,
    new_n13536_, new_n13538_, new_n13539_, new_n13540_, new_n13541_,
    new_n13542_, new_n13543_, new_n13544_, new_n13545_, new_n13546_,
    new_n13547_, new_n13548_, new_n13549_, new_n13550_, new_n13551_,
    new_n13552_, new_n13553_, new_n13554_, new_n13555_, new_n13556_,
    new_n13557_, new_n13558_, new_n13559_, new_n13560_, new_n13561_,
    new_n13562_, new_n13563_, new_n13564_, new_n13565_, new_n13566_,
    new_n13567_, new_n13568_, new_n13569_, new_n13570_, new_n13571_,
    new_n13572_, new_n13573_, new_n13574_, new_n13575_, new_n13576_,
    new_n13577_, new_n13578_, new_n13579_, new_n13580_, new_n13581_,
    new_n13582_, new_n13583_, new_n13584_, new_n13585_, new_n13586_,
    new_n13587_, new_n13588_, new_n13589_, new_n13590_, new_n13591_,
    new_n13592_, new_n13593_, new_n13594_, new_n13595_, new_n13596_,
    new_n13597_, new_n13598_, new_n13599_, new_n13600_, new_n13601_,
    new_n13602_, new_n13603_, new_n13604_, new_n13605_, new_n13606_,
    new_n13607_, new_n13608_, new_n13609_, new_n13610_, new_n13611_,
    new_n13612_, new_n13613_, new_n13614_, new_n13615_, new_n13616_,
    new_n13617_, new_n13618_, new_n13619_, new_n13620_, new_n13621_,
    new_n13622_, new_n13623_, new_n13624_, new_n13625_, new_n13626_,
    new_n13627_, new_n13628_, new_n13629_, new_n13630_, new_n13631_,
    new_n13632_, new_n13633_, new_n13634_, new_n13635_, new_n13636_,
    new_n13637_, new_n13638_, new_n13639_, new_n13640_, new_n13641_,
    new_n13642_, new_n13643_, new_n13644_, new_n13645_, new_n13646_,
    new_n13647_, new_n13648_, new_n13649_, new_n13650_, new_n13651_,
    new_n13652_, new_n13653_, new_n13654_, new_n13655_, new_n13656_,
    new_n13657_, new_n13658_, new_n13659_, new_n13660_, new_n13661_,
    new_n13662_, new_n13663_, new_n13664_, new_n13665_, new_n13666_,
    new_n13667_, new_n13668_, new_n13669_, new_n13670_, new_n13671_,
    new_n13672_, new_n13673_, new_n13674_, new_n13675_, new_n13676_,
    new_n13677_, new_n13678_, new_n13679_, new_n13680_, new_n13681_,
    new_n13682_, new_n13683_, new_n13684_, new_n13685_, new_n13686_,
    new_n13687_, new_n13688_, new_n13689_, new_n13690_, new_n13691_,
    new_n13692_, new_n13693_, new_n13694_, new_n13695_, new_n13696_,
    new_n13697_, new_n13698_, new_n13699_, new_n13700_, new_n13701_,
    new_n13702_, new_n13703_, new_n13704_, new_n13705_, new_n13706_,
    new_n13707_, new_n13708_, new_n13709_, new_n13710_, new_n13711_,
    new_n13712_, new_n13713_, new_n13714_, new_n13715_, new_n13716_,
    new_n13717_, new_n13718_, new_n13719_, new_n13720_, new_n13721_,
    new_n13722_, new_n13723_, new_n13724_, new_n13725_, new_n13726_,
    new_n13727_, new_n13728_, new_n13729_, new_n13730_, new_n13731_,
    new_n13732_, new_n13733_, new_n13734_, new_n13735_, new_n13736_,
    new_n13737_, new_n13738_, new_n13739_, new_n13740_, new_n13741_,
    new_n13742_, new_n13743_, new_n13744_, new_n13745_, new_n13746_,
    new_n13747_, new_n13748_, new_n13749_, new_n13750_, new_n13751_,
    new_n13752_, new_n13753_, new_n13754_, new_n13755_, new_n13756_,
    new_n13757_, new_n13758_, new_n13759_, new_n13760_, new_n13761_,
    new_n13762_, new_n13763_, new_n13764_, new_n13765_, new_n13766_,
    new_n13767_, new_n13768_, new_n13769_, new_n13770_, new_n13771_,
    new_n13772_, new_n13773_, new_n13774_, new_n13775_, new_n13776_,
    new_n13777_, new_n13778_, new_n13779_, new_n13780_, new_n13781_,
    new_n13782_, new_n13783_, new_n13784_, new_n13785_, new_n13786_,
    new_n13787_, new_n13788_, new_n13789_, new_n13790_, new_n13791_,
    new_n13792_, new_n13793_, new_n13794_, new_n13795_, new_n13796_,
    new_n13797_, new_n13798_, new_n13799_, new_n13800_, new_n13801_,
    new_n13802_, new_n13803_, new_n13804_, new_n13805_, new_n13806_,
    new_n13807_, new_n13808_, new_n13809_, new_n13810_, new_n13811_,
    new_n13812_, new_n13813_, new_n13814_, new_n13815_, new_n13816_,
    new_n13817_, new_n13818_, new_n13819_, new_n13820_, new_n13821_,
    new_n13822_, new_n13823_, new_n13824_, new_n13825_, new_n13826_,
    new_n13827_, new_n13828_, new_n13829_, new_n13830_, new_n13832_,
    new_n13833_, new_n13834_, new_n13835_, new_n13836_, new_n13837_,
    new_n13838_, new_n13839_, new_n13840_, new_n13841_, new_n13842_,
    new_n13843_, new_n13844_, new_n13845_, new_n13846_, new_n13847_,
    new_n13848_, new_n13849_, new_n13850_, new_n13851_, new_n13852_,
    new_n13853_, new_n13854_, new_n13855_, new_n13856_, new_n13857_,
    new_n13858_, new_n13859_, new_n13860_, new_n13861_, new_n13862_,
    new_n13863_, new_n13864_, new_n13865_, new_n13866_, new_n13867_,
    new_n13868_, new_n13869_, new_n13870_, new_n13871_, new_n13872_,
    new_n13873_, new_n13874_, new_n13875_, new_n13876_, new_n13877_,
    new_n13878_, new_n13879_, new_n13880_, new_n13881_, new_n13882_,
    new_n13883_, new_n13884_, new_n13885_, new_n13886_, new_n13887_,
    new_n13888_, new_n13889_, new_n13890_, new_n13891_, new_n13892_,
    new_n13893_, new_n13894_, new_n13895_, new_n13896_, new_n13897_,
    new_n13898_, new_n13899_, new_n13900_, new_n13901_, new_n13902_,
    new_n13903_, new_n13904_, new_n13905_, new_n13906_, new_n13907_,
    new_n13908_, new_n13909_, new_n13910_, new_n13911_, new_n13912_,
    new_n13913_, new_n13914_, new_n13915_, new_n13916_, new_n13917_,
    new_n13918_, new_n13919_, new_n13920_, new_n13921_, new_n13922_,
    new_n13923_, new_n13924_, new_n13925_, new_n13926_, new_n13927_,
    new_n13928_, new_n13929_, new_n13930_, new_n13931_, new_n13932_,
    new_n13933_, new_n13934_, new_n13935_, new_n13936_, new_n13937_,
    new_n13938_, new_n13939_, new_n13940_, new_n13941_, new_n13942_,
    new_n13943_, new_n13944_, new_n13945_, new_n13946_, new_n13947_,
    new_n13948_, new_n13949_, new_n13950_, new_n13951_, new_n13952_,
    new_n13953_, new_n13954_, new_n13955_, new_n13956_, new_n13957_,
    new_n13958_, new_n13959_, new_n13960_, new_n13961_, new_n13962_,
    new_n13963_, new_n13964_, new_n13965_, new_n13966_, new_n13967_,
    new_n13968_, new_n13969_, new_n13970_, new_n13971_, new_n13972_,
    new_n13973_, new_n13974_, new_n13975_, new_n13976_, new_n13977_,
    new_n13978_, new_n13979_, new_n13980_, new_n13981_, new_n13982_,
    new_n13983_, new_n13984_, new_n13985_, new_n13986_, new_n13987_,
    new_n13988_, new_n13989_, new_n13990_, new_n13991_, new_n13992_,
    new_n13993_, new_n13994_, new_n13995_, new_n13996_, new_n13997_,
    new_n13998_, new_n13999_, new_n14000_, new_n14001_, new_n14002_,
    new_n14003_, new_n14004_, new_n14005_, new_n14006_, new_n14007_,
    new_n14008_, new_n14009_, new_n14010_, new_n14011_, new_n14012_,
    new_n14013_, new_n14014_, new_n14015_, new_n14016_, new_n14017_,
    new_n14018_, new_n14019_, new_n14020_, new_n14021_, new_n14022_,
    new_n14023_, new_n14024_, new_n14025_, new_n14026_, new_n14027_,
    new_n14028_, new_n14029_, new_n14030_, new_n14031_, new_n14032_,
    new_n14033_, new_n14034_, new_n14035_, new_n14036_, new_n14037_,
    new_n14038_, new_n14039_, new_n14040_, new_n14041_, new_n14042_,
    new_n14043_, new_n14044_, new_n14045_, new_n14046_, new_n14047_,
    new_n14048_, new_n14049_, new_n14050_, new_n14051_, new_n14052_,
    new_n14053_, new_n14054_, new_n14055_, new_n14056_, new_n14057_,
    new_n14058_, new_n14059_, new_n14060_, new_n14061_, new_n14062_,
    new_n14063_, new_n14064_, new_n14065_, new_n14066_, new_n14067_,
    new_n14068_, new_n14069_, new_n14070_, new_n14071_, new_n14072_,
    new_n14073_, new_n14074_, new_n14075_, new_n14076_, new_n14077_,
    new_n14078_, new_n14079_, new_n14080_, new_n14081_, new_n14082_,
    new_n14083_, new_n14084_, new_n14085_, new_n14086_, new_n14087_,
    new_n14088_, new_n14089_, new_n14090_, new_n14091_, new_n14092_,
    new_n14093_, new_n14094_, new_n14095_, new_n14096_, new_n14097_,
    new_n14098_, new_n14099_, new_n14100_, new_n14101_, new_n14102_,
    new_n14103_, new_n14104_, new_n14105_, new_n14106_, new_n14107_,
    new_n14108_, new_n14109_, new_n14110_, new_n14111_, new_n14112_,
    new_n14113_, new_n14114_, new_n14115_, new_n14116_, new_n14117_,
    new_n14118_, new_n14119_, new_n14120_, new_n14121_, new_n14122_,
    new_n14123_, new_n14124_, new_n14125_, new_n14126_, new_n14127_,
    new_n14128_, new_n14129_, new_n14130_, new_n14131_, new_n14132_,
    new_n14133_, new_n14134_, new_n14135_, new_n14136_, new_n14137_,
    new_n14138_, new_n14139_, new_n14140_, new_n14141_, new_n14142_,
    new_n14143_, new_n14144_, new_n14145_, new_n14146_, new_n14147_,
    new_n14148_, new_n14149_, new_n14150_, new_n14151_, new_n14152_,
    new_n14153_, new_n14154_, new_n14155_, new_n14157_, new_n14158_,
    new_n14159_, new_n14160_, new_n14161_, new_n14162_, new_n14163_,
    new_n14164_, new_n14165_, new_n14166_, new_n14167_, new_n14168_,
    new_n14169_, new_n14170_, new_n14171_, new_n14172_, new_n14173_,
    new_n14174_, new_n14175_, new_n14176_, new_n14177_, new_n14178_,
    new_n14179_, new_n14180_, new_n14181_, new_n14182_, new_n14183_,
    new_n14184_, new_n14185_, new_n14186_, new_n14187_, new_n14188_,
    new_n14189_, new_n14190_, new_n14191_, new_n14192_, new_n14193_,
    new_n14194_, new_n14195_, new_n14196_, new_n14197_, new_n14198_,
    new_n14199_, new_n14200_, new_n14201_, new_n14202_, new_n14203_,
    new_n14204_, new_n14205_, new_n14206_, new_n14207_, new_n14208_,
    new_n14209_, new_n14210_, new_n14211_, new_n14212_, new_n14213_,
    new_n14214_, new_n14215_, new_n14216_, new_n14217_, new_n14218_,
    new_n14219_, new_n14220_, new_n14221_, new_n14222_, new_n14223_,
    new_n14224_, new_n14225_, new_n14226_, new_n14227_, new_n14228_,
    new_n14229_, new_n14230_, new_n14231_, new_n14232_, new_n14233_,
    new_n14234_, new_n14235_, new_n14236_, new_n14237_, new_n14238_,
    new_n14239_, new_n14240_, new_n14241_, new_n14242_, new_n14243_,
    new_n14244_, new_n14245_, new_n14246_, new_n14247_, new_n14248_,
    new_n14249_, new_n14250_, new_n14251_, new_n14252_, new_n14253_,
    new_n14254_, new_n14255_, new_n14256_, new_n14257_, new_n14258_,
    new_n14259_, new_n14260_, new_n14261_, new_n14262_, new_n14263_,
    new_n14264_, new_n14265_, new_n14266_, new_n14267_, new_n14268_,
    new_n14269_, new_n14270_, new_n14271_, new_n14272_, new_n14273_,
    new_n14274_, new_n14275_, new_n14276_, new_n14277_, new_n14278_,
    new_n14279_, new_n14280_, new_n14281_, new_n14282_, new_n14283_,
    new_n14284_, new_n14285_, new_n14286_, new_n14287_, new_n14288_,
    new_n14289_, new_n14290_, new_n14291_, new_n14292_, new_n14293_,
    new_n14294_, new_n14295_, new_n14296_, new_n14297_, new_n14298_,
    new_n14299_, new_n14300_, new_n14301_, new_n14302_, new_n14303_,
    new_n14304_, new_n14305_, new_n14306_, new_n14307_, new_n14308_,
    new_n14309_, new_n14310_, new_n14311_, new_n14312_, new_n14313_,
    new_n14314_, new_n14315_, new_n14316_, new_n14317_, new_n14318_,
    new_n14319_, new_n14320_, new_n14321_, new_n14322_, new_n14323_,
    new_n14324_, new_n14325_, new_n14326_, new_n14327_, new_n14328_,
    new_n14329_, new_n14330_, new_n14331_, new_n14332_, new_n14333_,
    new_n14334_, new_n14335_, new_n14336_, new_n14337_, new_n14338_,
    new_n14339_, new_n14340_, new_n14341_, new_n14342_, new_n14343_,
    new_n14344_, new_n14345_, new_n14346_, new_n14347_, new_n14348_,
    new_n14349_, new_n14350_, new_n14351_, new_n14352_, new_n14353_,
    new_n14354_, new_n14355_, new_n14356_, new_n14357_, new_n14358_,
    new_n14359_, new_n14360_, new_n14361_, new_n14362_, new_n14363_,
    new_n14364_, new_n14365_, new_n14366_, new_n14367_, new_n14368_,
    new_n14369_, new_n14370_, new_n14371_, new_n14372_, new_n14373_,
    new_n14374_, new_n14375_, new_n14376_, new_n14377_, new_n14378_,
    new_n14379_, new_n14380_, new_n14381_, new_n14382_, new_n14383_,
    new_n14384_, new_n14385_, new_n14386_, new_n14387_, new_n14388_,
    new_n14389_, new_n14390_, new_n14391_, new_n14392_, new_n14393_,
    new_n14394_, new_n14395_, new_n14396_, new_n14397_, new_n14398_,
    new_n14399_, new_n14400_, new_n14401_, new_n14402_, new_n14403_,
    new_n14404_, new_n14405_, new_n14406_, new_n14407_, new_n14408_,
    new_n14409_, new_n14410_, new_n14411_, new_n14412_, new_n14413_,
    new_n14414_, new_n14415_, new_n14416_, new_n14417_, new_n14418_,
    new_n14419_, new_n14420_, new_n14421_, new_n14422_, new_n14423_,
    new_n14424_, new_n14425_, new_n14426_, new_n14427_, new_n14428_,
    new_n14429_, new_n14430_, new_n14431_, new_n14432_, new_n14433_,
    new_n14434_, new_n14435_, new_n14436_, new_n14437_, new_n14438_,
    new_n14439_, new_n14440_, new_n14441_, new_n14442_, new_n14443_,
    new_n14444_, new_n14445_, new_n14446_, new_n14447_, new_n14448_,
    new_n14449_, new_n14450_, new_n14451_, new_n14453_, new_n14454_,
    new_n14455_, new_n14456_, new_n14457_, new_n14458_, new_n14459_,
    new_n14460_, new_n14461_, new_n14462_, new_n14463_, new_n14464_,
    new_n14465_, new_n14466_, new_n14467_, new_n14468_, new_n14469_,
    new_n14470_, new_n14471_, new_n14472_, new_n14473_, new_n14474_,
    new_n14475_, new_n14476_, new_n14477_, new_n14478_, new_n14479_,
    new_n14480_, new_n14481_, new_n14482_, new_n14483_, new_n14484_,
    new_n14485_, new_n14486_, new_n14487_, new_n14488_, new_n14489_,
    new_n14490_, new_n14491_, new_n14492_, new_n14493_, new_n14494_,
    new_n14495_, new_n14496_, new_n14497_, new_n14498_, new_n14500_,
    new_n14501_, new_n14502_, new_n14503_, new_n14504_, new_n14505_,
    new_n14506_, new_n14507_, new_n14508_, new_n14509_, new_n14510_,
    new_n14511_, new_n14512_, new_n14513_, new_n14514_, new_n14515_,
    new_n14516_, new_n14517_, new_n14518_, new_n14519_, new_n14520_,
    new_n14521_, new_n14522_, new_n14523_, new_n14524_, new_n14525_,
    new_n14526_, new_n14527_, new_n14528_, new_n14529_, new_n14530_,
    new_n14531_, new_n14532_, new_n14533_, new_n14534_, new_n14535_,
    new_n14536_, new_n14537_, new_n14538_, new_n14539_, new_n14540_,
    new_n14541_, new_n14542_, new_n14543_, new_n14544_, new_n14545_,
    new_n14546_, new_n14547_, new_n14548_, new_n14549_, new_n14550_,
    new_n14551_, new_n14552_, new_n14553_, new_n14554_, new_n14555_,
    new_n14556_, new_n14557_, new_n14558_, new_n14559_, new_n14560_,
    new_n14561_, new_n14562_, new_n14563_, new_n14564_, new_n14565_,
    new_n14566_, new_n14567_, new_n14568_, new_n14569_, new_n14570_,
    new_n14571_, new_n14572_, new_n14573_, new_n14574_, new_n14575_,
    new_n14576_, new_n14577_, new_n14578_, new_n14579_, new_n14580_,
    new_n14581_, new_n14582_, new_n14583_, new_n14584_, new_n14585_,
    new_n14586_, new_n14587_, new_n14588_, new_n14589_, new_n14590_,
    new_n14591_, new_n14592_, new_n14593_, new_n14594_, new_n14595_,
    new_n14596_, new_n14597_, new_n14599_, new_n14600_, new_n14601_,
    new_n14602_, new_n14603_, new_n14604_, new_n14605_, new_n14606_,
    new_n14607_, new_n14608_, new_n14609_, new_n14610_, new_n14611_,
    new_n14612_, new_n14613_, new_n14614_, new_n14615_, new_n14616_,
    new_n14617_, new_n14618_, new_n14619_, new_n14620_, new_n14621_,
    new_n14622_, new_n14623_, new_n14624_, new_n14625_, new_n14626_,
    new_n14627_, new_n14628_, new_n14629_, new_n14630_, new_n14631_,
    new_n14632_, new_n14633_, new_n14634_, new_n14635_, new_n14636_,
    new_n14637_, new_n14638_, new_n14640_, new_n14641_, new_n14642_,
    new_n14643_, new_n14644_, new_n14645_, new_n14646_, new_n14647_,
    new_n14648_, new_n14649_, new_n14650_, new_n14651_, new_n14652_,
    new_n14653_, new_n14654_, new_n14655_, new_n14656_, new_n14657_,
    new_n14658_, new_n14659_, new_n14660_, new_n14661_, new_n14662_,
    new_n14663_, new_n14664_, new_n14665_, new_n14666_, new_n14667_,
    new_n14668_, new_n14669_, new_n14670_, new_n14671_, new_n14672_,
    new_n14673_, new_n14674_, new_n14675_, new_n14677_, new_n14678_,
    new_n14679_, new_n14680_, new_n14681_, new_n14682_, new_n14683_,
    new_n14684_, new_n14685_, new_n14686_, new_n14687_, new_n14688_,
    new_n14689_, new_n14690_, new_n14691_, new_n14692_, new_n14693_,
    new_n14694_, new_n14695_, new_n14696_, new_n14697_, new_n14698_,
    new_n14699_, new_n14700_, new_n14701_, new_n14702_, new_n14703_,
    new_n14704_, new_n14705_, new_n14706_, new_n14707_, new_n14709_,
    new_n14710_, new_n14711_, new_n14712_, new_n14713_, new_n14714_,
    new_n14715_, new_n14716_, new_n14717_, new_n14718_, new_n14719_,
    new_n14720_, new_n14721_, new_n14722_, new_n14723_, new_n14724_,
    new_n14725_, new_n14726_, new_n14727_, new_n14728_, new_n14729_,
    new_n14730_, new_n14731_, new_n14732_, new_n14733_, new_n14734_,
    new_n14735_, new_n14736_, new_n14737_, new_n14738_, new_n14739_,
    new_n14740_, new_n14741_, new_n14742_, new_n14743_, new_n14744_,
    new_n14745_, new_n14746_, new_n14747_, new_n14748_, new_n14749_,
    new_n14750_, new_n14751_, new_n14752_, new_n14753_, new_n14754_,
    new_n14755_, new_n14756_, new_n14757_, new_n14758_, new_n14759_,
    new_n14760_, new_n14761_, new_n14762_, new_n14763_, new_n14764_,
    new_n14765_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14790_,
    new_n14791_, new_n14792_, new_n14793_, new_n14794_, new_n14795_,
    new_n14796_, new_n14797_, new_n14798_, new_n14799_, new_n14800_,
    new_n14801_, new_n14802_, new_n14803_, new_n14804_, new_n14805_,
    new_n14806_, new_n14807_, new_n14808_, new_n14809_, new_n14810_,
    new_n14811_, new_n14812_, new_n14813_, new_n14814_, new_n14815_,
    new_n14816_, new_n14817_, new_n14818_, new_n14819_, new_n14820_,
    new_n14821_, new_n14822_, new_n14823_, new_n14824_, new_n14825_,
    new_n14826_, new_n14827_, new_n14828_, new_n14829_, new_n14830_,
    new_n14831_, new_n14832_, new_n14833_, new_n14834_, new_n14835_,
    new_n14836_, new_n14837_, new_n14839_, new_n14840_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14846_,
    new_n14847_, new_n14848_, new_n14849_, new_n14850_, new_n14851_,
    new_n14852_, new_n14853_, new_n14854_, new_n14855_, new_n14856_,
    new_n14857_, new_n14858_, new_n14859_, new_n14860_, new_n14861_,
    new_n14862_, new_n14863_, new_n14864_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14871_,
    new_n14872_, new_n14873_, new_n14874_, new_n14875_, new_n14876_,
    new_n14877_, new_n14878_, new_n14879_, new_n14880_, new_n14881_,
    new_n14882_, new_n14883_, new_n14884_, new_n14885_, new_n14886_,
    new_n14887_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14893_, new_n14894_, new_n14895_, new_n14896_, new_n14897_,
    new_n14898_, new_n14899_, new_n14900_, new_n14901_, new_n14902_,
    new_n14903_, new_n14904_, new_n14905_, new_n14906_, new_n14907_,
    new_n14908_, new_n14909_, new_n14910_, new_n14911_, new_n14912_,
    new_n14913_, new_n14914_, new_n14915_, new_n14916_, new_n14917_,
    new_n14918_, new_n14919_, new_n14920_, new_n14921_, new_n14922_,
    new_n14923_, new_n14924_, new_n14925_, new_n14926_, new_n14928_,
    new_n14929_, new_n14930_, new_n14931_, new_n14932_, new_n14933_,
    new_n14934_, new_n14935_, new_n14936_, new_n14937_, new_n14938_,
    new_n14939_, new_n14940_, new_n14941_, new_n14942_, new_n14943_,
    new_n14944_, new_n14945_, new_n14946_, new_n14947_, new_n14948_,
    new_n14949_, new_n14950_, new_n14952_, new_n14953_, new_n14954_,
    new_n14955_, new_n14956_, new_n14957_, new_n14958_, new_n14959_,
    new_n14960_, new_n14961_, new_n14962_, new_n14963_, new_n14964_,
    new_n14965_, new_n14966_, new_n14967_, new_n14968_, new_n14970_,
    new_n14971_, new_n14972_, new_n14973_, new_n14974_, new_n14975_,
    new_n14976_, new_n14977_, new_n14978_, new_n14979_, new_n14980_,
    new_n14981_, new_n14982_, new_n14983_, new_n14984_, new_n14985_,
    new_n14986_, new_n14987_, new_n14988_, new_n14989_, new_n14990_,
    new_n14991_, new_n14992_, new_n14993_, new_n14994_, new_n14995_,
    new_n14996_, new_n14997_, new_n14998_, new_n14999_, new_n15000_,
    new_n15001_, new_n15002_, new_n15003_, new_n15004_, new_n15006_,
    new_n15007_, new_n15008_, new_n15009_, new_n15010_, new_n15011_,
    new_n15012_, new_n15013_, new_n15014_, new_n15015_, new_n15016_,
    new_n15017_, new_n15018_, new_n15019_, new_n15020_, new_n15021_,
    new_n15022_, new_n15023_, new_n15024_, new_n15025_, new_n15026_,
    new_n15027_, new_n15028_, new_n15029_, new_n15030_, new_n15031_,
    new_n15032_, new_n15033_, new_n15034_, new_n15035_, new_n15037_,
    new_n15038_, new_n15039_, new_n15040_, new_n15041_, new_n15042_,
    new_n15043_, new_n15044_, new_n15045_, new_n15046_, new_n15047_,
    new_n15048_, new_n15049_, new_n15050_, new_n15051_, new_n15052_,
    new_n15053_, new_n15054_, new_n15055_, new_n15056_, new_n15057_,
    new_n15058_, new_n15059_, new_n15060_, new_n15061_, new_n15062_,
    new_n15063_, new_n15064_, new_n15065_, new_n15066_, new_n15068_,
    new_n15069_, new_n15070_, new_n15071_, new_n15072_, new_n15073_,
    new_n15074_, new_n15075_, new_n15076_, new_n15077_, new_n15078_,
    new_n15079_, new_n15080_, new_n15081_, new_n15082_, new_n15083_,
    new_n15084_, new_n15085_, new_n15086_, new_n15087_, new_n15088_,
    new_n15089_, new_n15090_, new_n15091_, new_n15092_, new_n15093_,
    new_n15094_, new_n15095_, new_n15096_, new_n15097_, new_n15098_,
    new_n15099_, new_n15100_, new_n15101_, new_n15102_, new_n15104_,
    new_n15105_, new_n15106_, new_n15107_, new_n15108_, new_n15109_,
    new_n15110_, new_n15111_, new_n15112_, new_n15113_, new_n15114_,
    new_n15115_, new_n15116_, new_n15117_, new_n15118_, new_n15119_,
    new_n15120_, new_n15121_, new_n15122_, new_n15123_, new_n15124_,
    new_n15125_, new_n15126_, new_n15127_, new_n15128_, new_n15129_,
    new_n15130_, new_n15131_, new_n15132_, new_n15133_, new_n15134_,
    new_n15135_, new_n15136_, new_n15137_, new_n15138_, new_n15139_,
    new_n15140_, new_n15141_, new_n15142_, new_n15143_, new_n15144_,
    new_n15145_, new_n15146_, new_n15147_, new_n15148_, new_n15149_,
    new_n15150_, new_n15151_, new_n15152_, new_n15153_, new_n15154_,
    new_n15155_, new_n15156_, new_n15157_, new_n15158_, new_n15159_,
    new_n15161_, new_n15162_, new_n15163_, new_n15164_, new_n15165_,
    new_n15166_, new_n15167_, new_n15168_, new_n15169_, new_n15170_,
    new_n15171_, new_n15172_, new_n15173_, new_n15174_, new_n15175_,
    new_n15176_, new_n15177_, new_n15178_, new_n15179_, new_n15180_,
    new_n15181_, new_n15182_, new_n15183_, new_n15184_, new_n15185_,
    new_n15186_, new_n15187_, new_n15188_, new_n15189_, new_n15190_,
    new_n15191_, new_n15193_, new_n15194_, new_n15195_, new_n15196_,
    new_n15197_, new_n15198_, new_n15199_, new_n15200_, new_n15201_,
    new_n15202_, new_n15203_, new_n15204_, new_n15205_, new_n15206_,
    new_n15207_, new_n15208_, new_n15209_, new_n15210_, new_n15211_,
    new_n15212_, new_n15213_, new_n15214_, new_n15215_, new_n15216_,
    new_n15217_, new_n15218_, new_n15219_, new_n15220_, new_n15221_,
    new_n15222_, new_n15223_, new_n15224_, new_n15225_, new_n15226_,
    new_n15227_, new_n15229_, new_n15230_, new_n15231_, new_n15232_,
    new_n15233_, new_n15234_, new_n15235_, new_n15236_, new_n15237_,
    new_n15238_, new_n15239_, new_n15240_, new_n15241_, new_n15242_,
    new_n15243_, new_n15244_, new_n15245_, new_n15246_, new_n15247_,
    new_n15248_, new_n15249_, new_n15250_, new_n15252_, new_n15253_,
    new_n15254_, new_n15255_, new_n15256_, new_n15257_, new_n15258_,
    new_n15259_, new_n15260_, new_n15261_, new_n15262_, new_n15263_,
    new_n15264_, new_n15265_, new_n15266_, new_n15267_, new_n15268_,
    new_n15269_, new_n15270_, new_n15271_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15335_,
    new_n15336_, new_n15337_, new_n15338_, new_n15339_, new_n15340_,
    new_n15341_, new_n15342_, new_n15343_, new_n15344_, new_n15345_,
    new_n15346_, new_n15347_, new_n15348_, new_n15349_, new_n15350_,
    new_n15351_, new_n15352_, new_n15353_, new_n15354_, new_n15355_,
    new_n15356_, new_n15357_, new_n15358_, new_n15360_, new_n15361_,
    new_n15362_, new_n15363_, new_n15364_, new_n15365_, new_n15366_,
    new_n15367_, new_n15368_, new_n15369_, new_n15370_, new_n15371_,
    new_n15372_, new_n15373_, new_n15374_, new_n15375_, new_n15376_,
    new_n15377_, new_n15378_, new_n15379_, new_n15380_, new_n15381_,
    new_n15382_, new_n15383_, new_n15384_, new_n15385_, new_n15386_,
    new_n15387_, new_n15388_, new_n15389_, new_n15390_, new_n15391_,
    new_n15392_, new_n15393_, new_n15394_, new_n15395_, new_n15396_,
    new_n15397_, new_n15398_, new_n15399_, new_n15400_, new_n15401_,
    new_n15402_, new_n15403_, new_n15404_, new_n15405_, new_n15406_,
    new_n15407_, new_n15408_, new_n15409_, new_n15411_, new_n15412_,
    new_n15413_, new_n15414_, new_n15415_, new_n15416_, new_n15417_,
    new_n15418_, new_n15419_, new_n15420_, new_n15421_, new_n15422_,
    new_n15423_, new_n15424_, new_n15425_, new_n15426_, new_n15427_,
    new_n15428_, new_n15429_, new_n15430_, new_n15431_, new_n15432_,
    new_n15433_, new_n15434_, new_n15435_, new_n15436_, new_n15437_,
    new_n15438_, new_n15439_, new_n15440_, new_n15441_, new_n15442_,
    new_n15443_, new_n15444_, new_n15445_, new_n15446_, new_n15447_,
    new_n15448_, new_n15449_, new_n15450_, new_n15451_, new_n15452_,
    new_n15453_, new_n15454_, new_n15455_, new_n15456_, new_n15457_,
    new_n15458_, new_n15459_, new_n15460_, new_n15462_, new_n15463_,
    new_n15464_, new_n15465_, new_n15466_, new_n15467_, new_n15468_,
    new_n15469_, new_n15470_, new_n15471_, new_n15472_, new_n15473_,
    new_n15474_, new_n15475_, new_n15476_, new_n15477_, new_n15478_,
    new_n15479_, new_n15480_, new_n15481_, new_n15482_, new_n15483_,
    new_n15484_, new_n15485_, new_n15486_, new_n15487_, new_n15488_,
    new_n15489_, new_n15490_, new_n15491_, new_n15492_, new_n15493_,
    new_n15494_, new_n15495_, new_n15496_, new_n15497_, new_n15498_,
    new_n15499_, new_n15500_, new_n15501_, new_n15502_, new_n15503_,
    new_n15504_, new_n15505_, new_n15506_, new_n15507_, new_n15508_,
    new_n15509_, new_n15510_, new_n15512_, new_n15513_, new_n15514_,
    new_n15515_, new_n15516_, new_n15517_, new_n15518_, new_n15519_,
    new_n15520_, new_n15521_, new_n15522_, new_n15523_, new_n15524_,
    new_n15525_, new_n15526_, new_n15527_, new_n15528_, new_n15529_,
    new_n15530_, new_n15531_, new_n15532_, new_n15533_, new_n15534_,
    new_n15535_, new_n15536_, new_n15537_, new_n15538_, new_n15539_,
    new_n15540_, new_n15541_, new_n15542_, new_n15543_, new_n15544_,
    new_n15545_, new_n15546_, new_n15547_, new_n15548_, new_n15549_,
    new_n15550_, new_n15551_, new_n15552_, new_n15553_, new_n15554_,
    new_n15555_, new_n15556_, new_n15557_, new_n15558_, new_n15559_,
    new_n15560_, new_n15561_, new_n15563_, new_n15564_, new_n15565_,
    new_n15566_, new_n15567_, new_n15568_, new_n15569_, new_n15570_,
    new_n15571_, new_n15572_, new_n15573_, new_n15574_, new_n15575_,
    new_n15576_, new_n15577_, new_n15578_, new_n15579_, new_n15580_,
    new_n15581_, new_n15582_, new_n15583_, new_n15584_, new_n15585_,
    new_n15586_, new_n15587_, new_n15588_, new_n15589_, new_n15590_,
    new_n15591_, new_n15592_, new_n15593_, new_n15594_, new_n15595_,
    new_n15596_, new_n15597_, new_n15598_, new_n15599_, new_n15600_,
    new_n15601_, new_n15602_, new_n15603_, new_n15604_, new_n15605_,
    new_n15606_, new_n15607_, new_n15608_, new_n15609_, new_n15610_,
    new_n15611_, new_n15612_, new_n15613_, new_n15615_, new_n15616_,
    new_n15617_, new_n15618_, new_n15619_, new_n15620_, new_n15621_,
    new_n15622_, new_n15623_, new_n15624_, new_n15625_, new_n15626_,
    new_n15627_, new_n15628_, new_n15629_, new_n15630_, new_n15631_,
    new_n15632_, new_n15633_, new_n15634_, new_n15635_, new_n15636_,
    new_n15637_, new_n15638_, new_n15639_, new_n15640_, new_n15641_,
    new_n15642_, new_n15643_, new_n15644_, new_n15645_, new_n15646_,
    new_n15647_, new_n15648_, new_n15649_, new_n15650_, new_n15651_,
    new_n15652_, new_n15653_, new_n15654_, new_n15655_, new_n15656_,
    new_n15657_, new_n15658_, new_n15659_, new_n15660_, new_n15661_,
    new_n15662_, new_n15663_, new_n15664_, new_n15665_, new_n15666_,
    new_n15667_, new_n15668_, new_n15669_, new_n15670_, new_n15671_,
    new_n15672_, new_n15673_, new_n15674_, new_n15675_, new_n15676_,
    new_n15677_, new_n15678_, new_n15679_, new_n15680_, new_n15681_,
    new_n15682_, new_n15683_, new_n15684_, new_n15685_, new_n15686_,
    new_n15687_, new_n15688_, new_n15689_, new_n15690_, new_n15691_,
    new_n15692_, new_n15693_, new_n15694_, new_n15695_, new_n15696_,
    new_n15697_, new_n15698_, new_n15699_, new_n15700_, new_n15701_,
    new_n15702_, new_n15703_, new_n15704_, new_n15705_, new_n15706_,
    new_n15707_, new_n15708_, new_n15709_, new_n15710_, new_n15711_,
    new_n15712_, new_n15713_, new_n15714_, new_n15715_, new_n15716_,
    new_n15717_, new_n15718_, new_n15719_, new_n15720_, new_n15721_,
    new_n15722_, new_n15723_, new_n15724_, new_n15725_, new_n15726_,
    new_n15727_, new_n15728_, new_n15729_, new_n15730_, new_n15731_,
    new_n15732_, new_n15733_, new_n15734_, new_n15735_, new_n15736_,
    new_n15737_, new_n15738_, new_n15739_, new_n15740_, new_n15741_,
    new_n15742_, new_n15743_, new_n15744_, new_n15745_, new_n15746_,
    new_n15747_, new_n15748_, new_n15749_, new_n15750_, new_n15751_,
    new_n15752_, new_n15753_, new_n15754_, new_n15755_, new_n15756_,
    new_n15757_, new_n15758_, new_n15759_, new_n15760_, new_n15761_,
    new_n15762_, new_n15763_, new_n15764_, new_n15765_, new_n15766_,
    new_n15767_, new_n15768_, new_n15769_, new_n15770_, new_n15771_,
    new_n15772_, new_n15773_, new_n15774_, new_n15775_, new_n15776_,
    new_n15777_, new_n15778_, new_n15779_, new_n15780_, new_n15781_,
    new_n15782_, new_n15783_, new_n15784_, new_n15785_, new_n15786_,
    new_n15787_, new_n15788_, new_n15789_, new_n15790_, new_n15791_,
    new_n15792_, new_n15793_, new_n15794_, new_n15795_, new_n15796_,
    new_n15797_, new_n15798_, new_n15799_, new_n15800_, new_n15801_,
    new_n15802_, new_n15803_, new_n15804_, new_n15805_, new_n15806_,
    new_n15807_, new_n15808_, new_n15809_, new_n15810_, new_n15811_,
    new_n15812_, new_n15813_, new_n15814_, new_n15815_, new_n15816_,
    new_n15817_, new_n15818_, new_n15819_, new_n15820_, new_n15821_,
    new_n15822_, new_n15823_, new_n15824_, new_n15825_, new_n15826_,
    new_n15827_, new_n15828_, new_n15829_, new_n15830_, new_n15831_,
    new_n15832_, new_n15833_, new_n15834_, new_n15835_, new_n15836_,
    new_n15837_, new_n15838_, new_n15839_, new_n15840_, new_n15841_,
    new_n15842_, new_n15843_, new_n15844_, new_n15845_, new_n15846_,
    new_n15847_, new_n15848_, new_n15849_, new_n15850_, new_n15851_,
    new_n15852_, new_n15853_, new_n15854_, new_n15855_, new_n15856_,
    new_n15857_, new_n15858_, new_n15859_, new_n15860_, new_n15861_,
    new_n15862_, new_n15863_, new_n15864_, new_n15865_, new_n15866_,
    new_n15867_, new_n15868_, new_n15869_, new_n15870_, new_n15871_,
    new_n15872_, new_n15873_, new_n15874_, new_n15875_, new_n15876_,
    new_n15877_, new_n15878_, new_n15879_, new_n15880_, new_n15881_,
    new_n15882_, new_n15883_, new_n15884_, new_n15885_, new_n15886_,
    new_n15887_, new_n15888_, new_n15890_, new_n15891_, new_n15892_,
    new_n15893_, new_n15894_, new_n15895_, new_n15896_, new_n15897_,
    new_n15898_, new_n15899_, new_n15900_, new_n15901_, new_n15902_,
    new_n15903_, new_n15904_, new_n15905_, new_n15906_, new_n15907_,
    new_n15908_, new_n15909_, new_n15910_, new_n15911_, new_n15912_,
    new_n15913_, new_n15914_, new_n15915_, new_n15916_, new_n15917_,
    new_n15918_, new_n15919_, new_n15920_, new_n15921_, new_n15922_,
    new_n15923_, new_n15924_, new_n15925_, new_n15926_, new_n15927_,
    new_n15928_, new_n15929_, new_n15930_, new_n15931_, new_n15932_,
    new_n15933_, new_n15934_, new_n15935_, new_n15936_, new_n15937_,
    new_n15938_, new_n15939_, new_n15940_, new_n15941_, new_n15942_,
    new_n15943_, new_n15944_, new_n15945_, new_n15946_, new_n15947_,
    new_n15948_, new_n15949_, new_n15950_, new_n15951_, new_n15952_,
    new_n15953_, new_n15954_, new_n15955_, new_n15956_, new_n15957_,
    new_n15958_, new_n15959_, new_n15960_, new_n15961_, new_n15962_,
    new_n15963_, new_n15964_, new_n15965_, new_n15966_, new_n15967_,
    new_n15968_, new_n15969_, new_n15970_, new_n15971_, new_n15972_,
    new_n15973_, new_n15974_, new_n15975_, new_n15976_, new_n15977_,
    new_n15978_, new_n15979_, new_n15980_, new_n15981_, new_n15982_,
    new_n15983_, new_n15984_, new_n15985_, new_n15986_, new_n15987_,
    new_n15988_, new_n15989_, new_n15990_, new_n15991_, new_n15992_,
    new_n15993_, new_n15994_, new_n15995_, new_n15996_, new_n15997_,
    new_n15998_, new_n15999_, new_n16000_, new_n16001_, new_n16002_,
    new_n16003_, new_n16004_, new_n16005_, new_n16006_, new_n16007_,
    new_n16008_, new_n16009_, new_n16010_, new_n16011_, new_n16012_,
    new_n16013_, new_n16014_, new_n16015_, new_n16016_, new_n16017_,
    new_n16018_, new_n16019_, new_n16020_, new_n16021_, new_n16022_,
    new_n16023_, new_n16024_, new_n16025_, new_n16026_, new_n16027_,
    new_n16028_, new_n16029_, new_n16030_, new_n16031_, new_n16032_,
    new_n16033_, new_n16034_, new_n16035_, new_n16036_, new_n16037_,
    new_n16038_, new_n16039_, new_n16040_, new_n16041_, new_n16042_,
    new_n16043_, new_n16044_, new_n16045_, new_n16046_, new_n16047_,
    new_n16048_, new_n16049_, new_n16050_, new_n16051_, new_n16052_,
    new_n16053_, new_n16054_, new_n16055_, new_n16056_, new_n16057_,
    new_n16058_, new_n16059_, new_n16060_, new_n16061_, new_n16062_,
    new_n16063_, new_n16064_, new_n16065_, new_n16066_, new_n16067_,
    new_n16068_, new_n16069_, new_n16070_, new_n16071_, new_n16072_,
    new_n16073_, new_n16074_, new_n16075_, new_n16076_, new_n16077_,
    new_n16078_, new_n16079_, new_n16080_, new_n16081_, new_n16082_,
    new_n16083_, new_n16084_, new_n16085_, new_n16086_, new_n16087_,
    new_n16088_, new_n16089_, new_n16090_, new_n16091_, new_n16092_,
    new_n16093_, new_n16094_, new_n16095_, new_n16096_, new_n16097_,
    new_n16098_, new_n16099_, new_n16100_, new_n16101_, new_n16102_,
    new_n16103_, new_n16104_, new_n16105_, new_n16106_, new_n16107_,
    new_n16108_, new_n16109_, new_n16110_, new_n16111_, new_n16112_,
    new_n16113_, new_n16114_, new_n16115_, new_n16116_, new_n16117_,
    new_n16118_, new_n16119_, new_n16120_, new_n16121_, new_n16122_,
    new_n16123_, new_n16124_, new_n16125_, new_n16126_, new_n16127_,
    new_n16128_, new_n16129_, new_n16130_, new_n16131_, new_n16132_,
    new_n16133_, new_n16134_, new_n16135_, new_n16136_, new_n16137_,
    new_n16138_, new_n16139_, new_n16140_, new_n16141_, new_n16142_,
    new_n16143_, new_n16144_, new_n16145_, new_n16146_, new_n16147_,
    new_n16148_, new_n16149_, new_n16150_, new_n16151_, new_n16152_,
    new_n16153_, new_n16154_, new_n16155_, new_n16156_, new_n16157_,
    new_n16158_, new_n16159_, new_n16160_, new_n16161_, new_n16162_,
    new_n16163_, new_n16164_, new_n16165_, new_n16166_, new_n16167_,
    new_n16168_, new_n16169_, new_n16170_, new_n16171_, new_n16172_,
    new_n16173_, new_n16174_, new_n16175_, new_n16177_, new_n16178_,
    new_n16179_, new_n16180_, new_n16181_, new_n16182_, new_n16183_,
    new_n16184_, new_n16185_, new_n16186_, new_n16187_, new_n16188_,
    new_n16189_, new_n16190_, new_n16191_, new_n16192_, new_n16193_,
    new_n16194_, new_n16195_, new_n16196_, new_n16197_, new_n16198_,
    new_n16199_, new_n16200_, new_n16201_, new_n16202_, new_n16203_,
    new_n16204_, new_n16205_, new_n16206_, new_n16207_, new_n16208_,
    new_n16209_, new_n16210_, new_n16211_, new_n16212_, new_n16213_,
    new_n16214_, new_n16215_, new_n16216_, new_n16217_, new_n16218_,
    new_n16219_, new_n16220_, new_n16221_, new_n16222_, new_n16223_,
    new_n16224_, new_n16225_, new_n16226_, new_n16227_, new_n16228_,
    new_n16229_, new_n16230_, new_n16231_, new_n16232_, new_n16233_,
    new_n16234_, new_n16235_, new_n16236_, new_n16237_, new_n16238_,
    new_n16239_, new_n16240_, new_n16241_, new_n16242_, new_n16243_,
    new_n16244_, new_n16245_, new_n16246_, new_n16247_, new_n16248_,
    new_n16249_, new_n16250_, new_n16251_, new_n16252_, new_n16253_,
    new_n16254_, new_n16255_, new_n16256_, new_n16257_, new_n16258_,
    new_n16259_, new_n16260_, new_n16261_, new_n16262_, new_n16263_,
    new_n16264_, new_n16265_, new_n16266_, new_n16267_, new_n16268_,
    new_n16269_, new_n16270_, new_n16271_, new_n16272_, new_n16273_,
    new_n16274_, new_n16275_, new_n16276_, new_n16277_, new_n16278_,
    new_n16279_, new_n16280_, new_n16281_, new_n16282_, new_n16283_,
    new_n16284_, new_n16285_, new_n16286_, new_n16287_, new_n16288_,
    new_n16289_, new_n16290_, new_n16291_, new_n16292_, new_n16293_,
    new_n16294_, new_n16295_, new_n16296_, new_n16297_, new_n16298_,
    new_n16299_, new_n16300_, new_n16301_, new_n16302_, new_n16303_,
    new_n16304_, new_n16305_, new_n16306_, new_n16307_, new_n16308_,
    new_n16309_, new_n16310_, new_n16311_, new_n16312_, new_n16313_,
    new_n16314_, new_n16315_, new_n16316_, new_n16317_, new_n16318_,
    new_n16319_, new_n16320_, new_n16321_, new_n16322_, new_n16323_,
    new_n16324_, new_n16325_, new_n16326_, new_n16327_, new_n16328_,
    new_n16329_, new_n16330_, new_n16331_, new_n16332_, new_n16333_,
    new_n16334_, new_n16335_, new_n16336_, new_n16337_, new_n16338_,
    new_n16339_, new_n16340_, new_n16341_, new_n16342_, new_n16343_,
    new_n16344_, new_n16345_, new_n16346_, new_n16347_, new_n16348_,
    new_n16349_, new_n16350_, new_n16351_, new_n16352_, new_n16353_,
    new_n16354_, new_n16355_, new_n16356_, new_n16357_, new_n16358_,
    new_n16359_, new_n16360_, new_n16361_, new_n16362_, new_n16363_,
    new_n16364_, new_n16365_, new_n16366_, new_n16367_, new_n16368_,
    new_n16369_, new_n16370_, new_n16371_, new_n16372_, new_n16373_,
    new_n16374_, new_n16375_, new_n16376_, new_n16377_, new_n16378_,
    new_n16379_, new_n16380_, new_n16381_, new_n16382_, new_n16383_,
    new_n16384_, new_n16385_, new_n16386_, new_n16387_, new_n16388_,
    new_n16389_, new_n16390_, new_n16391_, new_n16392_, new_n16393_,
    new_n16394_, new_n16395_, new_n16396_, new_n16397_, new_n16398_,
    new_n16399_, new_n16400_, new_n16401_, new_n16402_, new_n16403_,
    new_n16404_, new_n16405_, new_n16406_, new_n16407_, new_n16408_,
    new_n16409_, new_n16410_, new_n16411_, new_n16412_, new_n16413_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16420_, new_n16421_, new_n16422_, new_n16423_,
    new_n16424_, new_n16425_, new_n16426_, new_n16427_, new_n16428_,
    new_n16429_, new_n16430_, new_n16431_, new_n16432_, new_n16433_,
    new_n16434_, new_n16435_, new_n16436_, new_n16437_, new_n16438_,
    new_n16439_, new_n16440_, new_n16441_, new_n16442_, new_n16443_,
    new_n16444_, new_n16445_, new_n16446_, new_n16447_, new_n16448_,
    new_n16449_, new_n16450_, new_n16451_, new_n16452_, new_n16453_,
    new_n16454_, new_n16455_, new_n16456_, new_n16457_, new_n16458_,
    new_n16459_, new_n16460_, new_n16462_, new_n16463_, new_n16464_,
    new_n16465_, new_n16466_, new_n16467_, new_n16468_, new_n16469_,
    new_n16470_, new_n16471_, new_n16472_, new_n16473_, new_n16474_,
    new_n16475_, new_n16476_, new_n16477_, new_n16478_, new_n16479_,
    new_n16480_, new_n16481_, new_n16482_, new_n16483_, new_n16484_,
    new_n16485_, new_n16486_, new_n16487_, new_n16488_, new_n16489_,
    new_n16490_, new_n16491_, new_n16492_, new_n16493_, new_n16494_,
    new_n16495_, new_n16496_, new_n16497_, new_n16498_, new_n16499_,
    new_n16500_, new_n16501_, new_n16502_, new_n16503_, new_n16504_,
    new_n16505_, new_n16506_, new_n16507_, new_n16508_, new_n16509_,
    new_n16510_, new_n16511_, new_n16512_, new_n16513_, new_n16514_,
    new_n16515_, new_n16516_, new_n16517_, new_n16518_, new_n16519_,
    new_n16520_, new_n16521_, new_n16522_, new_n16523_, new_n16524_,
    new_n16525_, new_n16526_, new_n16527_, new_n16528_, new_n16529_,
    new_n16530_, new_n16531_, new_n16532_, new_n16533_, new_n16534_,
    new_n16535_, new_n16536_, new_n16537_, new_n16538_, new_n16539_,
    new_n16540_, new_n16541_, new_n16542_, new_n16543_, new_n16544_,
    new_n16545_, new_n16546_, new_n16547_, new_n16548_, new_n16549_,
    new_n16550_, new_n16551_, new_n16552_, new_n16553_, new_n16554_,
    new_n16555_, new_n16556_, new_n16557_, new_n16558_, new_n16559_,
    new_n16560_, new_n16561_, new_n16562_, new_n16563_, new_n16564_,
    new_n16565_, new_n16566_, new_n16567_, new_n16568_, new_n16569_,
    new_n16570_, new_n16571_, new_n16572_, new_n16573_, new_n16574_,
    new_n16575_, new_n16576_, new_n16577_, new_n16578_, new_n16579_,
    new_n16580_, new_n16581_, new_n16582_, new_n16583_, new_n16584_,
    new_n16585_, new_n16586_, new_n16587_, new_n16588_, new_n16589_,
    new_n16590_, new_n16591_, new_n16592_, new_n16593_, new_n16594_,
    new_n16595_, new_n16596_, new_n16597_, new_n16598_, new_n16599_,
    new_n16600_, new_n16601_, new_n16602_, new_n16603_, new_n16604_,
    new_n16605_, new_n16606_, new_n16607_, new_n16608_, new_n16609_,
    new_n16610_, new_n16611_, new_n16612_, new_n16613_, new_n16614_,
    new_n16615_, new_n16616_, new_n16617_, new_n16618_, new_n16619_,
    new_n16620_, new_n16621_, new_n16622_, new_n16623_, new_n16624_,
    new_n16625_, new_n16626_, new_n16627_, new_n16628_, new_n16629_,
    new_n16630_, new_n16631_, new_n16632_, new_n16633_, new_n16634_,
    new_n16635_, new_n16636_, new_n16637_, new_n16638_, new_n16639_,
    new_n16640_, new_n16641_, new_n16642_, new_n16643_, new_n16644_,
    new_n16645_, new_n16646_, new_n16647_, new_n16648_, new_n16649_,
    new_n16650_, new_n16651_, new_n16652_, new_n16653_, new_n16654_,
    new_n16655_, new_n16656_, new_n16657_, new_n16658_, new_n16659_,
    new_n16660_, new_n16661_, new_n16662_, new_n16663_, new_n16664_,
    new_n16665_, new_n16666_, new_n16667_, new_n16668_, new_n16669_,
    new_n16670_, new_n16671_, new_n16672_, new_n16673_, new_n16674_,
    new_n16675_, new_n16676_, new_n16677_, new_n16678_, new_n16679_,
    new_n16680_, new_n16681_, new_n16682_, new_n16683_, new_n16684_,
    new_n16685_, new_n16686_, new_n16687_, new_n16688_, new_n16689_,
    new_n16690_, new_n16691_, new_n16692_, new_n16693_, new_n16694_,
    new_n16695_, new_n16696_, new_n16697_, new_n16698_, new_n16699_,
    new_n16700_, new_n16701_, new_n16702_, new_n16703_, new_n16704_,
    new_n16705_, new_n16706_, new_n16707_, new_n16708_, new_n16709_,
    new_n16710_, new_n16711_, new_n16712_, new_n16713_, new_n16714_,
    new_n16715_, new_n16716_, new_n16717_, new_n16718_, new_n16719_,
    new_n16720_, new_n16721_, new_n16722_, new_n16723_, new_n16724_,
    new_n16725_, new_n16726_, new_n16728_, new_n16729_, new_n16730_,
    new_n16731_, new_n16732_, new_n16733_, new_n16734_, new_n16735_,
    new_n16736_, new_n16737_, new_n16738_, new_n16739_, new_n16740_,
    new_n16741_, new_n16742_, new_n16743_, new_n16744_, new_n16745_,
    new_n16746_, new_n16747_, new_n16748_, new_n16749_, new_n16750_,
    new_n16751_, new_n16752_, new_n16753_, new_n16754_, new_n16755_,
    new_n16756_, new_n16757_, new_n16758_, new_n16759_, new_n16760_,
    new_n16761_, new_n16762_, new_n16763_, new_n16764_, new_n16765_,
    new_n16766_, new_n16767_, new_n16768_, new_n16769_, new_n16770_,
    new_n16771_, new_n16772_, new_n16773_, new_n16774_, new_n16775_,
    new_n16776_, new_n16777_, new_n16778_, new_n16779_, new_n16780_,
    new_n16781_, new_n16782_, new_n16783_, new_n16784_, new_n16785_,
    new_n16786_, new_n16787_, new_n16788_, new_n16789_, new_n16790_,
    new_n16791_, new_n16792_, new_n16793_, new_n16794_, new_n16795_,
    new_n16796_, new_n16797_, new_n16798_, new_n16799_, new_n16800_,
    new_n16801_, new_n16802_, new_n16803_, new_n16804_, new_n16805_,
    new_n16806_, new_n16807_, new_n16808_, new_n16809_, new_n16810_,
    new_n16811_, new_n16812_, new_n16813_, new_n16814_, new_n16815_,
    new_n16816_, new_n16817_, new_n16818_, new_n16819_, new_n16820_,
    new_n16821_, new_n16822_, new_n16823_, new_n16824_, new_n16825_,
    new_n16826_, new_n16827_, new_n16828_, new_n16829_, new_n16830_,
    new_n16831_, new_n16832_, new_n16833_, new_n16834_, new_n16835_,
    new_n16836_, new_n16837_, new_n16838_, new_n16839_, new_n16840_,
    new_n16841_, new_n16842_, new_n16843_, new_n16844_, new_n16845_,
    new_n16846_, new_n16847_, new_n16848_, new_n16849_, new_n16850_,
    new_n16851_, new_n16852_, new_n16853_, new_n16854_, new_n16855_,
    new_n16856_, new_n16857_, new_n16858_, new_n16859_, new_n16860_,
    new_n16861_, new_n16862_, new_n16863_, new_n16864_, new_n16865_,
    new_n16866_, new_n16867_, new_n16868_, new_n16869_, new_n16870_,
    new_n16871_, new_n16872_, new_n16873_, new_n16874_, new_n16875_,
    new_n16876_, new_n16877_, new_n16878_, new_n16879_, new_n16880_,
    new_n16881_, new_n16882_, new_n16883_, new_n16884_, new_n16885_,
    new_n16886_, new_n16887_, new_n16888_, new_n16889_, new_n16890_,
    new_n16891_, new_n16892_, new_n16893_, new_n16894_, new_n16895_,
    new_n16896_, new_n16897_, new_n16898_, new_n16899_, new_n16900_,
    new_n16901_, new_n16902_, new_n16903_, new_n16904_, new_n16905_,
    new_n16906_, new_n16907_, new_n16908_, new_n16909_, new_n16910_,
    new_n16911_, new_n16912_, new_n16913_, new_n16914_, new_n16915_,
    new_n16916_, new_n16917_, new_n16918_, new_n16919_, new_n16920_,
    new_n16921_, new_n16922_, new_n16923_, new_n16924_, new_n16925_,
    new_n16926_, new_n16927_, new_n16928_, new_n16929_, new_n16930_,
    new_n16931_, new_n16932_, new_n16933_, new_n16934_, new_n16935_,
    new_n16936_, new_n16937_, new_n16938_, new_n16939_, new_n16940_,
    new_n16941_, new_n16942_, new_n16943_, new_n16944_, new_n16945_,
    new_n16946_, new_n16947_, new_n16948_, new_n16949_, new_n16950_,
    new_n16951_, new_n16952_, new_n16953_, new_n16954_, new_n16955_,
    new_n16956_, new_n16957_, new_n16958_, new_n16959_, new_n16960_,
    new_n16961_, new_n16962_, new_n16963_, new_n16964_, new_n16965_,
    new_n16966_, new_n16967_, new_n16968_, new_n16969_, new_n16970_,
    new_n16971_, new_n16972_, new_n16973_, new_n16974_, new_n16975_,
    new_n16976_, new_n16977_, new_n16978_, new_n16979_, new_n16980_,
    new_n16981_, new_n16982_, new_n16983_, new_n16984_, new_n16985_,
    new_n16986_, new_n16987_, new_n16988_, new_n16989_, new_n16990_,
    new_n16991_, new_n16992_, new_n16993_, new_n16994_, new_n16995_,
    new_n16996_, new_n16997_, new_n16998_, new_n16999_, new_n17000_,
    new_n17001_, new_n17002_, new_n17003_, new_n17004_, new_n17005_,
    new_n17006_, new_n17007_, new_n17008_, new_n17009_, new_n17010_,
    new_n17011_, new_n17012_, new_n17013_, new_n17014_, new_n17016_,
    new_n17017_, new_n17018_, new_n17019_, new_n17020_, new_n17021_,
    new_n17022_, new_n17023_, new_n17024_, new_n17025_, new_n17026_,
    new_n17027_, new_n17028_, new_n17029_, new_n17030_, new_n17031_,
    new_n17032_, new_n17033_, new_n17034_, new_n17035_, new_n17036_,
    new_n17037_, new_n17038_, new_n17039_, new_n17040_, new_n17041_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17105_, new_n17106_,
    new_n17107_, new_n17108_, new_n17109_, new_n17110_, new_n17111_,
    new_n17112_, new_n17113_, new_n17114_, new_n17115_, new_n17116_,
    new_n17117_, new_n17118_, new_n17119_, new_n17120_, new_n17121_,
    new_n17122_, new_n17123_, new_n17124_, new_n17125_, new_n17126_,
    new_n17127_, new_n17128_, new_n17129_, new_n17130_, new_n17131_,
    new_n17132_, new_n17133_, new_n17134_, new_n17135_, new_n17136_,
    new_n17137_, new_n17138_, new_n17139_, new_n17140_, new_n17141_,
    new_n17142_, new_n17143_, new_n17144_, new_n17145_, new_n17146_,
    new_n17147_, new_n17148_, new_n17149_, new_n17150_, new_n17151_,
    new_n17152_, new_n17153_, new_n17154_, new_n17155_, new_n17156_,
    new_n17157_, new_n17158_, new_n17159_, new_n17160_, new_n17161_,
    new_n17162_, new_n17163_, new_n17164_, new_n17165_, new_n17166_,
    new_n17167_, new_n17168_, new_n17169_, new_n17170_, new_n17171_,
    new_n17172_, new_n17173_, new_n17174_, new_n17175_, new_n17176_,
    new_n17177_, new_n17178_, new_n17179_, new_n17180_, new_n17181_,
    new_n17182_, new_n17183_, new_n17184_, new_n17185_, new_n17186_,
    new_n17187_, new_n17188_, new_n17189_, new_n17190_, new_n17191_,
    new_n17192_, new_n17193_, new_n17194_, new_n17195_, new_n17196_,
    new_n17197_, new_n17198_, new_n17199_, new_n17200_, new_n17201_,
    new_n17202_, new_n17203_, new_n17204_, new_n17205_, new_n17206_,
    new_n17207_, new_n17208_, new_n17209_, new_n17210_, new_n17211_,
    new_n17212_, new_n17213_, new_n17214_, new_n17215_, new_n17216_,
    new_n17217_, new_n17218_, new_n17219_, new_n17220_, new_n17221_,
    new_n17222_, new_n17223_, new_n17224_, new_n17225_, new_n17226_,
    new_n17227_, new_n17228_, new_n17229_, new_n17230_, new_n17231_,
    new_n17232_, new_n17233_, new_n17234_, new_n17235_, new_n17236_,
    new_n17237_, new_n17238_, new_n17239_, new_n17240_, new_n17241_,
    new_n17242_, new_n17243_, new_n17244_, new_n17245_, new_n17246_,
    new_n17247_, new_n17248_, new_n17249_, new_n17250_, new_n17251_,
    new_n17252_, new_n17253_, new_n17254_, new_n17255_, new_n17256_,
    new_n17257_, new_n17258_, new_n17259_, new_n17260_, new_n17261_,
    new_n17262_, new_n17263_, new_n17264_, new_n17265_, new_n17266_,
    new_n17267_, new_n17268_, new_n17269_, new_n17270_, new_n17271_,
    new_n17272_, new_n17273_, new_n17274_, new_n17275_, new_n17276_,
    new_n17277_, new_n17278_, new_n17279_, new_n17280_, new_n17281_,
    new_n17282_, new_n17284_, new_n17285_, new_n17286_, new_n17287_,
    new_n17288_, new_n17289_, new_n17290_, new_n17291_, new_n17292_,
    new_n17293_, new_n17294_, new_n17295_, new_n17296_, new_n17297_,
    new_n17298_, new_n17299_, new_n17300_, new_n17301_, new_n17302_,
    new_n17303_, new_n17304_, new_n17305_, new_n17306_, new_n17307_,
    new_n17308_, new_n17309_, new_n17310_, new_n17311_, new_n17312_,
    new_n17313_, new_n17314_, new_n17315_, new_n17316_, new_n17317_,
    new_n17318_, new_n17319_, new_n17320_, new_n17321_, new_n17322_,
    new_n17323_, new_n17324_, new_n17325_, new_n17326_, new_n17327_,
    new_n17328_, new_n17329_, new_n17330_, new_n17331_, new_n17332_,
    new_n17333_, new_n17334_, new_n17335_, new_n17336_, new_n17337_,
    new_n17338_, new_n17339_, new_n17340_, new_n17341_, new_n17342_,
    new_n17343_, new_n17344_, new_n17345_, new_n17346_, new_n17347_,
    new_n17348_, new_n17349_, new_n17350_, new_n17351_, new_n17352_,
    new_n17353_, new_n17354_, new_n17355_, new_n17356_, new_n17357_,
    new_n17358_, new_n17359_, new_n17360_, new_n17361_, new_n17362_,
    new_n17363_, new_n17364_, new_n17365_, new_n17366_, new_n17367_,
    new_n17368_, new_n17369_, new_n17370_, new_n17371_, new_n17372_,
    new_n17373_, new_n17374_, new_n17375_, new_n17376_, new_n17377_,
    new_n17378_, new_n17379_, new_n17380_, new_n17381_, new_n17382_,
    new_n17383_, new_n17384_, new_n17385_, new_n17386_, new_n17387_,
    new_n17388_, new_n17389_, new_n17390_, new_n17391_, new_n17392_,
    new_n17393_, new_n17394_, new_n17395_, new_n17396_, new_n17397_,
    new_n17398_, new_n17399_, new_n17400_, new_n17401_, new_n17402_,
    new_n17403_, new_n17404_, new_n17405_, new_n17406_, new_n17407_,
    new_n17408_, new_n17409_, new_n17410_, new_n17411_, new_n17412_,
    new_n17413_, new_n17414_, new_n17415_, new_n17416_, new_n17417_,
    new_n17418_, new_n17419_, new_n17420_, new_n17421_, new_n17422_,
    new_n17423_, new_n17424_, new_n17425_, new_n17426_, new_n17427_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17441_, new_n17442_,
    new_n17443_, new_n17444_, new_n17445_, new_n17446_, new_n17447_,
    new_n17448_, new_n17449_, new_n17450_, new_n17451_, new_n17452_,
    new_n17453_, new_n17454_, new_n17455_, new_n17456_, new_n17457_,
    new_n17458_, new_n17459_, new_n17460_, new_n17461_, new_n17462_,
    new_n17463_, new_n17464_, new_n17465_, new_n17466_, new_n17467_,
    new_n17468_, new_n17469_, new_n17470_, new_n17471_, new_n17472_,
    new_n17473_, new_n17474_, new_n17475_, new_n17476_, new_n17477_,
    new_n17478_, new_n17479_, new_n17480_, new_n17481_, new_n17482_,
    new_n17483_, new_n17484_, new_n17485_, new_n17486_, new_n17487_,
    new_n17488_, new_n17489_, new_n17490_, new_n17491_, new_n17492_,
    new_n17493_, new_n17494_, new_n17495_, new_n17496_, new_n17497_,
    new_n17498_, new_n17499_, new_n17500_, new_n17501_, new_n17502_,
    new_n17503_, new_n17504_, new_n17505_, new_n17506_, new_n17507_,
    new_n17508_, new_n17509_, new_n17510_, new_n17511_, new_n17512_,
    new_n17513_, new_n17514_, new_n17515_, new_n17516_, new_n17517_,
    new_n17518_, new_n17519_, new_n17520_, new_n17521_, new_n17522_,
    new_n17523_, new_n17524_, new_n17525_, new_n17526_, new_n17527_,
    new_n17528_, new_n17529_, new_n17530_, new_n17531_, new_n17532_,
    new_n17533_, new_n17534_, new_n17535_, new_n17536_, new_n17537_,
    new_n17538_, new_n17539_, new_n17540_, new_n17541_, new_n17542_,
    new_n17543_, new_n17544_, new_n17545_, new_n17546_, new_n17547_,
    new_n17548_, new_n17549_, new_n17550_, new_n17551_, new_n17552_,
    new_n17553_, new_n17554_, new_n17555_, new_n17556_, new_n17557_,
    new_n17558_, new_n17559_, new_n17561_, new_n17562_, new_n17563_,
    new_n17564_, new_n17565_, new_n17566_, new_n17567_, new_n17568_,
    new_n17569_, new_n17570_, new_n17571_, new_n17572_, new_n17573_,
    new_n17574_, new_n17575_, new_n17576_, new_n17577_, new_n17578_,
    new_n17579_, new_n17580_, new_n17581_, new_n17582_, new_n17583_,
    new_n17584_, new_n17585_, new_n17586_, new_n17587_, new_n17588_,
    new_n17589_, new_n17590_, new_n17591_, new_n17592_, new_n17593_,
    new_n17594_, new_n17595_, new_n17596_, new_n17597_, new_n17598_,
    new_n17599_, new_n17600_, new_n17601_, new_n17602_, new_n17603_,
    new_n17604_, new_n17605_, new_n17606_, new_n17607_, new_n17608_,
    new_n17609_, new_n17610_, new_n17611_, new_n17612_, new_n17613_,
    new_n17614_, new_n17615_, new_n17616_, new_n17617_, new_n17618_,
    new_n17619_, new_n17620_, new_n17621_, new_n17622_, new_n17623_,
    new_n17624_, new_n17625_, new_n17626_, new_n17627_, new_n17628_,
    new_n17629_, new_n17630_, new_n17631_, new_n17632_, new_n17633_,
    new_n17634_, new_n17635_, new_n17636_, new_n17637_, new_n17638_,
    new_n17639_, new_n17640_, new_n17641_, new_n17642_, new_n17643_,
    new_n17644_, new_n17645_, new_n17646_, new_n17647_, new_n17648_,
    new_n17649_, new_n17650_, new_n17651_, new_n17652_, new_n17653_,
    new_n17654_, new_n17655_, new_n17656_, new_n17657_, new_n17658_,
    new_n17659_, new_n17660_, new_n17661_, new_n17662_, new_n17663_,
    new_n17664_, new_n17665_, new_n17666_, new_n17667_, new_n17668_,
    new_n17669_, new_n17670_, new_n17671_, new_n17672_, new_n17673_,
    new_n17674_, new_n17675_, new_n17676_, new_n17677_, new_n17678_,
    new_n17679_, new_n17680_, new_n17681_, new_n17682_, new_n17683_,
    new_n17684_, new_n17685_, new_n17686_, new_n17687_, new_n17688_,
    new_n17689_, new_n17690_, new_n17691_, new_n17692_, new_n17693_,
    new_n17694_, new_n17695_, new_n17696_, new_n17697_, new_n17698_,
    new_n17699_, new_n17700_, new_n17701_, new_n17702_, new_n17703_,
    new_n17704_, new_n17705_, new_n17706_, new_n17707_, new_n17708_,
    new_n17709_, new_n17710_, new_n17711_, new_n17712_, new_n17713_,
    new_n17714_, new_n17715_, new_n17716_, new_n17717_, new_n17718_,
    new_n17719_, new_n17720_, new_n17721_, new_n17722_, new_n17723_,
    new_n17724_, new_n17725_, new_n17726_, new_n17727_, new_n17728_,
    new_n17729_, new_n17730_, new_n17731_, new_n17732_, new_n17733_,
    new_n17734_, new_n17735_, new_n17736_, new_n17737_, new_n17738_,
    new_n17739_, new_n17740_, new_n17741_, new_n17742_, new_n17743_,
    new_n17744_, new_n17745_, new_n17746_, new_n17747_, new_n17748_,
    new_n17749_, new_n17750_, new_n17751_, new_n17752_, new_n17753_,
    new_n17754_, new_n17755_, new_n17756_, new_n17757_, new_n17758_,
    new_n17759_, new_n17760_, new_n17761_, new_n17762_, new_n17763_,
    new_n17764_, new_n17765_, new_n17766_, new_n17767_, new_n17768_,
    new_n17769_, new_n17770_, new_n17771_, new_n17772_, new_n17773_,
    new_n17774_, new_n17775_, new_n17776_, new_n17777_, new_n17778_,
    new_n17779_, new_n17780_, new_n17781_, new_n17782_, new_n17783_,
    new_n17784_, new_n17785_, new_n17786_, new_n17787_, new_n17788_,
    new_n17789_, new_n17790_, new_n17791_, new_n17792_, new_n17793_,
    new_n17794_, new_n17795_, new_n17796_, new_n17797_, new_n17798_,
    new_n17799_, new_n17800_, new_n17801_, new_n17802_, new_n17803_,
    new_n17804_, new_n17805_, new_n17806_, new_n17807_, new_n17808_,
    new_n17809_, new_n17810_, new_n17811_, new_n17812_, new_n17813_,
    new_n17814_, new_n17815_, new_n17816_, new_n17817_, new_n17818_,
    new_n17819_, new_n17820_, new_n17821_, new_n17822_, new_n17823_,
    new_n17824_, new_n17825_, new_n17826_, new_n17827_, new_n17828_,
    new_n17829_, new_n17830_, new_n17831_, new_n17832_, new_n17833_,
    new_n17835_, new_n17836_, new_n17837_, new_n17838_, new_n17839_,
    new_n17840_, new_n17841_, new_n17842_, new_n17843_, new_n17844_,
    new_n17845_, new_n17846_, new_n17847_, new_n17848_, new_n17849_,
    new_n17850_, new_n17851_, new_n17852_, new_n17853_, new_n17854_,
    new_n17855_, new_n17856_, new_n17857_, new_n17858_, new_n17859_,
    new_n17860_, new_n17861_, new_n17862_, new_n17863_, new_n17864_,
    new_n17865_, new_n17866_, new_n17867_, new_n17868_, new_n17869_,
    new_n17870_, new_n17871_, new_n17872_, new_n17873_, new_n17874_,
    new_n17875_, new_n17876_, new_n17877_, new_n17878_, new_n17879_,
    new_n17880_, new_n17881_, new_n17882_, new_n17883_, new_n17884_,
    new_n17885_, new_n17886_, new_n17887_, new_n17888_, new_n17889_,
    new_n17890_, new_n17891_, new_n17892_, new_n17893_, new_n17894_,
    new_n17895_, new_n17896_, new_n17897_, new_n17898_, new_n17899_,
    new_n17900_, new_n17901_, new_n17902_, new_n17903_, new_n17904_,
    new_n17905_, new_n17906_, new_n17907_, new_n17908_, new_n17909_,
    new_n17910_, new_n17911_, new_n17912_, new_n17913_, new_n17914_,
    new_n17915_, new_n17916_, new_n17917_, new_n17918_, new_n17919_,
    new_n17920_, new_n17921_, new_n17922_, new_n17923_, new_n17924_,
    new_n17925_, new_n17926_, new_n17927_, new_n17928_, new_n17929_,
    new_n17930_, new_n17931_, new_n17932_, new_n17933_, new_n17934_,
    new_n17935_, new_n17936_, new_n17937_, new_n17938_, new_n17939_,
    new_n17940_, new_n17941_, new_n17942_, new_n17943_, new_n17944_,
    new_n17945_, new_n17946_, new_n17947_, new_n17948_, new_n17949_,
    new_n17950_, new_n17951_, new_n17952_, new_n17953_, new_n17954_,
    new_n17955_, new_n17956_, new_n17957_, new_n17958_, new_n17959_,
    new_n17960_, new_n17961_, new_n17962_, new_n17963_, new_n17964_,
    new_n17965_, new_n17966_, new_n17967_, new_n17968_, new_n17969_,
    new_n17970_, new_n17971_, new_n17972_, new_n17973_, new_n17974_,
    new_n17975_, new_n17976_, new_n17977_, new_n17978_, new_n17979_,
    new_n17980_, new_n17981_, new_n17982_, new_n17983_, new_n17984_,
    new_n17985_, new_n17986_, new_n17987_, new_n17988_, new_n17989_,
    new_n17990_, new_n17991_, new_n17992_, new_n17993_, new_n17994_,
    new_n17995_, new_n17996_, new_n17997_, new_n17998_, new_n17999_,
    new_n18000_, new_n18001_, new_n18002_, new_n18003_, new_n18004_,
    new_n18005_, new_n18006_, new_n18007_, new_n18008_, new_n18009_,
    new_n18010_, new_n18011_, new_n18012_, new_n18013_, new_n18014_,
    new_n18015_, new_n18016_, new_n18017_, new_n18018_, new_n18019_,
    new_n18020_, new_n18021_, new_n18022_, new_n18023_, new_n18024_,
    new_n18025_, new_n18026_, new_n18027_, new_n18028_, new_n18029_,
    new_n18030_, new_n18031_, new_n18032_, new_n18033_, new_n18034_,
    new_n18035_, new_n18036_, new_n18037_, new_n18038_, new_n18039_,
    new_n18040_, new_n18041_, new_n18042_, new_n18043_, new_n18044_,
    new_n18045_, new_n18046_, new_n18047_, new_n18048_, new_n18049_,
    new_n18050_, new_n18051_, new_n18052_, new_n18053_, new_n18054_,
    new_n18055_, new_n18056_, new_n18057_, new_n18058_, new_n18059_,
    new_n18060_, new_n18061_, new_n18062_, new_n18063_, new_n18064_,
    new_n18065_, new_n18066_, new_n18067_, new_n18068_, new_n18069_,
    new_n18070_, new_n18071_, new_n18072_, new_n18073_, new_n18074_,
    new_n18075_, new_n18076_, new_n18077_, new_n18078_, new_n18079_,
    new_n18080_, new_n18081_, new_n18082_, new_n18083_, new_n18084_,
    new_n18085_, new_n18086_, new_n18087_, new_n18088_, new_n18089_,
    new_n18090_, new_n18091_, new_n18092_, new_n18093_, new_n18094_,
    new_n18095_, new_n18096_, new_n18097_, new_n18098_, new_n18099_,
    new_n18100_, new_n18101_, new_n18102_, new_n18103_, new_n18104_,
    new_n18105_, new_n18106_, new_n18107_, new_n18109_, new_n18110_,
    new_n18111_, new_n18112_, new_n18113_, new_n18114_, new_n18115_,
    new_n18116_, new_n18117_, new_n18118_, new_n18119_, new_n18120_,
    new_n18121_, new_n18122_, new_n18123_, new_n18124_, new_n18125_,
    new_n18126_, new_n18127_, new_n18128_, new_n18129_, new_n18130_,
    new_n18131_, new_n18132_, new_n18133_, new_n18134_, new_n18135_,
    new_n18136_, new_n18137_, new_n18138_, new_n18139_, new_n18140_,
    new_n18141_, new_n18142_, new_n18143_, new_n18144_, new_n18145_,
    new_n18146_, new_n18147_, new_n18148_, new_n18149_, new_n18150_,
    new_n18151_, new_n18152_, new_n18153_, new_n18154_, new_n18155_,
    new_n18156_, new_n18157_, new_n18158_, new_n18159_, new_n18160_,
    new_n18161_, new_n18162_, new_n18163_, new_n18164_, new_n18165_,
    new_n18166_, new_n18167_, new_n18168_, new_n18169_, new_n18170_,
    new_n18171_, new_n18172_, new_n18173_, new_n18174_, new_n18175_,
    new_n18176_, new_n18177_, new_n18178_, new_n18179_, new_n18180_,
    new_n18181_, new_n18182_, new_n18183_, new_n18184_, new_n18185_,
    new_n18186_, new_n18187_, new_n18188_, new_n18189_, new_n18190_,
    new_n18191_, new_n18192_, new_n18193_, new_n18194_, new_n18195_,
    new_n18196_, new_n18197_, new_n18198_, new_n18199_, new_n18200_,
    new_n18201_, new_n18202_, new_n18203_, new_n18204_, new_n18205_,
    new_n18206_, new_n18207_, new_n18208_, new_n18209_, new_n18210_,
    new_n18211_, new_n18212_, new_n18213_, new_n18214_, new_n18215_,
    new_n18216_, new_n18217_, new_n18218_, new_n18219_, new_n18220_,
    new_n18221_, new_n18222_, new_n18223_, new_n18224_, new_n18225_,
    new_n18226_, new_n18227_, new_n18228_, new_n18229_, new_n18230_,
    new_n18231_, new_n18232_, new_n18233_, new_n18234_, new_n18235_,
    new_n18236_, new_n18237_, new_n18238_, new_n18239_, new_n18240_,
    new_n18241_, new_n18242_, new_n18243_, new_n18244_, new_n18245_,
    new_n18246_, new_n18247_, new_n18248_, new_n18249_, new_n18250_,
    new_n18251_, new_n18252_, new_n18253_, new_n18254_, new_n18255_,
    new_n18256_, new_n18257_, new_n18258_, new_n18259_, new_n18260_,
    new_n18261_, new_n18262_, new_n18263_, new_n18264_, new_n18265_,
    new_n18266_, new_n18267_, new_n18268_, new_n18269_, new_n18270_,
    new_n18271_, new_n18272_, new_n18273_, new_n18274_, new_n18275_,
    new_n18276_, new_n18277_, new_n18278_, new_n18279_, new_n18280_,
    new_n18281_, new_n18282_, new_n18283_, new_n18284_, new_n18285_,
    new_n18286_, new_n18287_, new_n18288_, new_n18289_, new_n18290_,
    new_n18291_, new_n18292_, new_n18293_, new_n18294_, new_n18295_,
    new_n18296_, new_n18297_, new_n18298_, new_n18299_, new_n18300_,
    new_n18301_, new_n18302_, new_n18303_, new_n18304_, new_n18305_,
    new_n18306_, new_n18307_, new_n18308_, new_n18309_, new_n18310_,
    new_n18311_, new_n18312_, new_n18313_, new_n18314_, new_n18315_,
    new_n18316_, new_n18317_, new_n18318_, new_n18319_, new_n18320_,
    new_n18321_, new_n18322_, new_n18323_, new_n18324_, new_n18325_,
    new_n18326_, new_n18327_, new_n18328_, new_n18329_, new_n18330_,
    new_n18331_, new_n18332_, new_n18333_, new_n18334_, new_n18335_,
    new_n18336_, new_n18337_, new_n18338_, new_n18339_, new_n18340_,
    new_n18341_, new_n18342_, new_n18343_, new_n18344_, new_n18345_,
    new_n18346_, new_n18347_, new_n18348_, new_n18349_, new_n18350_,
    new_n18351_, new_n18352_, new_n18353_, new_n18354_, new_n18355_,
    new_n18356_, new_n18357_, new_n18358_, new_n18359_, new_n18360_,
    new_n18361_, new_n18362_, new_n18363_, new_n18364_, new_n18365_,
    new_n18366_, new_n18367_, new_n18368_, new_n18369_, new_n18370_,
    new_n18371_, new_n18372_, new_n18373_, new_n18374_, new_n18375_,
    new_n18377_, new_n18378_, new_n18379_, new_n18380_, new_n18381_,
    new_n18382_, new_n18383_, new_n18384_, new_n18385_, new_n18386_,
    new_n18387_, new_n18388_, new_n18389_, new_n18390_, new_n18391_,
    new_n18392_, new_n18393_, new_n18394_, new_n18395_, new_n18396_,
    new_n18397_, new_n18398_, new_n18399_, new_n18400_, new_n18401_,
    new_n18402_, new_n18403_, new_n18404_, new_n18405_, new_n18406_,
    new_n18407_, new_n18408_, new_n18409_, new_n18410_, new_n18411_,
    new_n18412_, new_n18413_, new_n18414_, new_n18415_, new_n18416_,
    new_n18417_, new_n18418_, new_n18419_, new_n18420_, new_n18421_,
    new_n18422_, new_n18423_, new_n18424_, new_n18425_, new_n18426_,
    new_n18427_, new_n18428_, new_n18429_, new_n18430_, new_n18431_,
    new_n18432_, new_n18433_, new_n18434_, new_n18435_, new_n18436_,
    new_n18437_, new_n18438_, new_n18439_, new_n18440_, new_n18441_,
    new_n18442_, new_n18443_, new_n18444_, new_n18445_, new_n18446_,
    new_n18447_, new_n18448_, new_n18449_, new_n18450_, new_n18451_,
    new_n18452_, new_n18453_, new_n18454_, new_n18455_, new_n18456_,
    new_n18457_, new_n18458_, new_n18459_, new_n18460_, new_n18461_,
    new_n18462_, new_n18463_, new_n18464_, new_n18465_, new_n18466_,
    new_n18467_, new_n18468_, new_n18469_, new_n18470_, new_n18471_,
    new_n18472_, new_n18473_, new_n18474_, new_n18475_, new_n18476_,
    new_n18477_, new_n18478_, new_n18479_, new_n18480_, new_n18481_,
    new_n18482_, new_n18483_, new_n18484_, new_n18485_, new_n18486_,
    new_n18487_, new_n18488_, new_n18489_, new_n18490_, new_n18491_,
    new_n18492_, new_n18493_, new_n18494_, new_n18495_, new_n18496_,
    new_n18497_, new_n18498_, new_n18499_, new_n18500_, new_n18501_,
    new_n18502_, new_n18503_, new_n18504_, new_n18505_, new_n18506_,
    new_n18507_, new_n18508_, new_n18509_, new_n18510_, new_n18511_,
    new_n18512_, new_n18513_, new_n18514_, new_n18515_, new_n18516_,
    new_n18517_, new_n18518_, new_n18519_, new_n18520_, new_n18521_,
    new_n18522_, new_n18523_, new_n18524_, new_n18525_, new_n18526_,
    new_n18527_, new_n18528_, new_n18529_, new_n18530_, new_n18531_,
    new_n18532_, new_n18533_, new_n18534_, new_n18535_, new_n18536_,
    new_n18537_, new_n18538_, new_n18539_, new_n18540_, new_n18541_,
    new_n18542_, new_n18543_, new_n18544_, new_n18545_, new_n18546_,
    new_n18547_, new_n18548_, new_n18549_, new_n18550_, new_n18551_,
    new_n18552_, new_n18553_, new_n18554_, new_n18555_, new_n18556_,
    new_n18557_, new_n18558_, new_n18559_, new_n18560_, new_n18561_,
    new_n18562_, new_n18563_, new_n18564_, new_n18565_, new_n18566_,
    new_n18567_, new_n18568_, new_n18569_, new_n18570_, new_n18571_,
    new_n18572_, new_n18573_, new_n18574_, new_n18575_, new_n18576_,
    new_n18577_, new_n18578_, new_n18579_, new_n18580_, new_n18581_,
    new_n18582_, new_n18583_, new_n18584_, new_n18585_, new_n18586_,
    new_n18587_, new_n18588_, new_n18589_, new_n18590_, new_n18591_,
    new_n18592_, new_n18593_, new_n18594_, new_n18595_, new_n18596_,
    new_n18597_, new_n18598_, new_n18599_, new_n18600_, new_n18601_,
    new_n18602_, new_n18603_, new_n18604_, new_n18605_, new_n18606_,
    new_n18607_, new_n18608_, new_n18609_, new_n18610_, new_n18611_,
    new_n18612_, new_n18613_, new_n18614_, new_n18615_, new_n18616_,
    new_n18617_, new_n18618_, new_n18619_, new_n18620_, new_n18621_,
    new_n18622_, new_n18623_, new_n18624_, new_n18625_, new_n18626_,
    new_n18627_, new_n18628_, new_n18629_, new_n18630_, new_n18631_,
    new_n18632_, new_n18633_, new_n18634_, new_n18635_, new_n18636_,
    new_n18637_, new_n18638_, new_n18639_, new_n18640_, new_n18641_,
    new_n18642_, new_n18643_, new_n18645_, new_n18646_, new_n18647_,
    new_n18648_, new_n18649_, new_n18650_, new_n18651_, new_n18652_,
    new_n18653_, new_n18654_, new_n18655_, new_n18656_, new_n18657_,
    new_n18658_, new_n18659_, new_n18660_, new_n18661_, new_n18662_,
    new_n18663_, new_n18664_, new_n18665_, new_n18666_, new_n18667_,
    new_n18668_, new_n18669_, new_n18670_, new_n18671_, new_n18672_,
    new_n18673_, new_n18674_, new_n18675_, new_n18676_, new_n18677_,
    new_n18678_, new_n18679_, new_n18680_, new_n18681_, new_n18682_,
    new_n18683_, new_n18684_, new_n18685_, new_n18686_, new_n18687_,
    new_n18688_, new_n18689_, new_n18690_, new_n18691_, new_n18692_,
    new_n18693_, new_n18694_, new_n18695_, new_n18696_, new_n18697_,
    new_n18698_, new_n18699_, new_n18700_, new_n18701_, new_n18702_,
    new_n18703_, new_n18704_, new_n18705_, new_n18706_, new_n18707_,
    new_n18708_, new_n18709_, new_n18710_, new_n18711_, new_n18712_,
    new_n18713_, new_n18714_, new_n18715_, new_n18716_, new_n18717_,
    new_n18718_, new_n18719_, new_n18720_, new_n18721_, new_n18722_,
    new_n18723_, new_n18724_, new_n18725_, new_n18726_, new_n18727_,
    new_n18728_, new_n18729_, new_n18730_, new_n18731_, new_n18732_,
    new_n18733_, new_n18734_, new_n18735_, new_n18736_, new_n18737_,
    new_n18738_, new_n18739_, new_n18740_, new_n18741_, new_n18742_,
    new_n18743_, new_n18744_, new_n18745_, new_n18746_, new_n18747_,
    new_n18748_, new_n18749_, new_n18750_, new_n18751_, new_n18752_,
    new_n18753_, new_n18754_, new_n18755_, new_n18756_, new_n18757_,
    new_n18758_, new_n18759_, new_n18760_, new_n18761_, new_n18762_,
    new_n18763_, new_n18764_, new_n18765_, new_n18766_, new_n18767_,
    new_n18768_, new_n18769_, new_n18770_, new_n18771_, new_n18772_,
    new_n18773_, new_n18774_, new_n18775_, new_n18776_, new_n18777_,
    new_n18778_, new_n18779_, new_n18780_, new_n18781_, new_n18782_,
    new_n18783_, new_n18784_, new_n18785_, new_n18786_, new_n18787_,
    new_n18788_, new_n18789_, new_n18790_, new_n18791_, new_n18792_,
    new_n18793_, new_n18794_, new_n18795_, new_n18796_, new_n18797_,
    new_n18798_, new_n18799_, new_n18800_, new_n18801_, new_n18802_,
    new_n18803_, new_n18804_, new_n18805_, new_n18806_, new_n18807_,
    new_n18808_, new_n18809_, new_n18810_, new_n18811_, new_n18812_,
    new_n18813_, new_n18814_, new_n18815_, new_n18816_, new_n18817_,
    new_n18818_, new_n18819_, new_n18820_, new_n18821_, new_n18822_,
    new_n18823_, new_n18824_, new_n18825_, new_n18826_, new_n18827_,
    new_n18828_, new_n18829_, new_n18830_, new_n18831_, new_n18832_,
    new_n18833_, new_n18834_, new_n18835_, new_n18836_, new_n18837_,
    new_n18838_, new_n18839_, new_n18840_, new_n18841_, new_n18842_,
    new_n18843_, new_n18844_, new_n18845_, new_n18846_, new_n18847_,
    new_n18848_, new_n18849_, new_n18850_, new_n18851_, new_n18852_,
    new_n18853_, new_n18854_, new_n18855_, new_n18856_, new_n18857_,
    new_n18858_, new_n18859_, new_n18860_, new_n18861_, new_n18862_,
    new_n18863_, new_n18864_, new_n18865_, new_n18866_, new_n18867_,
    new_n18868_, new_n18869_, new_n18870_, new_n18871_, new_n18872_,
    new_n18873_, new_n18874_, new_n18875_, new_n18876_, new_n18877_,
    new_n18878_, new_n18879_, new_n18880_, new_n18881_, new_n18882_,
    new_n18883_, new_n18884_, new_n18885_, new_n18886_, new_n18887_,
    new_n18888_, new_n18889_, new_n18890_, new_n18891_, new_n18892_,
    new_n18893_, new_n18894_, new_n18895_, new_n18896_, new_n18897_,
    new_n18898_, new_n18899_, new_n18900_, new_n18901_, new_n18902_,
    new_n18903_, new_n18904_, new_n18905_, new_n18906_, new_n18907_,
    new_n18908_, new_n18909_, new_n18910_, new_n18911_, new_n18913_,
    new_n18914_, new_n18915_, new_n18916_, new_n18917_, new_n18918_,
    new_n18919_, new_n18920_, new_n18921_, new_n18922_, new_n18923_,
    new_n18924_, new_n18925_, new_n18926_, new_n18927_, new_n18928_,
    new_n18929_, new_n18930_, new_n18931_, new_n18932_, new_n18933_,
    new_n18934_, new_n18935_, new_n18936_, new_n18937_, new_n18938_,
    new_n18939_, new_n18940_, new_n18941_, new_n18942_, new_n18943_,
    new_n18944_, new_n18945_, new_n18946_, new_n18947_, new_n18948_,
    new_n18949_, new_n18950_, new_n18951_, new_n18952_, new_n18953_,
    new_n18954_, new_n18955_, new_n18956_, new_n18957_, new_n18958_,
    new_n18959_, new_n18960_, new_n18961_, new_n18962_, new_n18963_,
    new_n18964_, new_n18965_, new_n18966_, new_n18967_, new_n18968_,
    new_n18969_, new_n18970_, new_n18971_, new_n18972_, new_n18973_,
    new_n18974_, new_n18975_, new_n18976_, new_n18977_, new_n18978_,
    new_n18979_, new_n18980_, new_n18981_, new_n18982_, new_n18983_,
    new_n18984_, new_n18985_, new_n18986_, new_n18987_, new_n18988_,
    new_n18989_, new_n18990_, new_n18991_, new_n18992_, new_n18993_,
    new_n18994_, new_n18995_, new_n18996_, new_n18997_, new_n18998_,
    new_n18999_, new_n19000_, new_n19001_, new_n19002_, new_n19003_,
    new_n19004_, new_n19005_, new_n19006_, new_n19007_, new_n19008_,
    new_n19009_, new_n19010_, new_n19011_, new_n19012_, new_n19013_,
    new_n19014_, new_n19015_, new_n19016_, new_n19017_, new_n19018_,
    new_n19019_, new_n19020_, new_n19021_, new_n19022_, new_n19023_,
    new_n19024_, new_n19025_, new_n19026_, new_n19027_, new_n19028_,
    new_n19029_, new_n19030_, new_n19031_, new_n19032_, new_n19033_,
    new_n19034_, new_n19035_, new_n19036_, new_n19037_, new_n19038_,
    new_n19039_, new_n19040_, new_n19041_, new_n19042_, new_n19043_,
    new_n19044_, new_n19045_, new_n19046_, new_n19047_, new_n19048_,
    new_n19049_, new_n19050_, new_n19051_, new_n19052_, new_n19053_,
    new_n19054_, new_n19055_, new_n19056_, new_n19057_, new_n19058_,
    new_n19059_, new_n19060_, new_n19061_, new_n19062_, new_n19063_,
    new_n19064_, new_n19065_, new_n19066_, new_n19067_, new_n19068_,
    new_n19069_, new_n19070_, new_n19071_, new_n19072_, new_n19073_,
    new_n19074_, new_n19075_, new_n19076_, new_n19077_, new_n19078_,
    new_n19079_, new_n19080_, new_n19081_, new_n19082_, new_n19083_,
    new_n19084_, new_n19085_, new_n19086_, new_n19087_, new_n19088_,
    new_n19089_, new_n19090_, new_n19091_, new_n19092_, new_n19093_,
    new_n19094_, new_n19095_, new_n19096_, new_n19097_, new_n19098_,
    new_n19099_, new_n19100_, new_n19101_, new_n19102_, new_n19103_,
    new_n19104_, new_n19105_, new_n19106_, new_n19107_, new_n19108_,
    new_n19109_, new_n19110_, new_n19111_, new_n19112_, new_n19113_,
    new_n19114_, new_n19115_, new_n19116_, new_n19117_, new_n19118_,
    new_n19119_, new_n19120_, new_n19121_, new_n19122_, new_n19123_,
    new_n19124_, new_n19125_, new_n19126_, new_n19127_, new_n19128_,
    new_n19129_, new_n19130_, new_n19131_, new_n19132_, new_n19133_,
    new_n19134_, new_n19135_, new_n19136_, new_n19137_, new_n19138_,
    new_n19139_, new_n19140_, new_n19141_, new_n19142_, new_n19143_,
    new_n19144_, new_n19145_, new_n19146_, new_n19147_, new_n19148_,
    new_n19149_, new_n19150_, new_n19151_, new_n19152_, new_n19153_,
    new_n19154_, new_n19155_, new_n19156_, new_n19157_, new_n19158_,
    new_n19159_, new_n19160_, new_n19161_, new_n19162_, new_n19163_,
    new_n19164_, new_n19165_, new_n19166_, new_n19167_, new_n19168_,
    new_n19169_, new_n19170_, new_n19171_, new_n19172_, new_n19173_,
    new_n19174_, new_n19175_, new_n19176_, new_n19177_, new_n19178_,
    new_n19179_, new_n19180_, new_n19181_, new_n19182_, new_n19183_,
    new_n19184_, new_n19185_, new_n19187_, new_n19188_, new_n19189_,
    new_n19190_, new_n19191_, new_n19192_, new_n19193_, new_n19194_,
    new_n19195_, new_n19196_, new_n19197_, new_n19198_, new_n19199_,
    new_n19200_, new_n19201_, new_n19202_, new_n19203_, new_n19204_,
    new_n19205_, new_n19206_, new_n19207_, new_n19208_, new_n19209_,
    new_n19210_, new_n19211_, new_n19212_, new_n19213_, new_n19214_,
    new_n19215_, new_n19216_, new_n19217_, new_n19218_, new_n19219_,
    new_n19220_, new_n19221_, new_n19222_, new_n19223_, new_n19224_,
    new_n19225_, new_n19226_, new_n19227_, new_n19228_, new_n19229_,
    new_n19230_, new_n19231_, new_n19232_, new_n19233_, new_n19234_,
    new_n19235_, new_n19236_, new_n19237_, new_n19238_, new_n19239_,
    new_n19240_, new_n19241_, new_n19242_, new_n19243_, new_n19244_,
    new_n19245_, new_n19246_, new_n19247_, new_n19248_, new_n19249_,
    new_n19250_, new_n19251_, new_n19252_, new_n19253_, new_n19254_,
    new_n19255_, new_n19256_, new_n19257_, new_n19258_, new_n19259_,
    new_n19260_, new_n19261_, new_n19262_, new_n19263_, new_n19264_,
    new_n19265_, new_n19266_, new_n19267_, new_n19268_, new_n19269_,
    new_n19270_, new_n19271_, new_n19272_, new_n19273_, new_n19274_,
    new_n19275_, new_n19276_, new_n19277_, new_n19278_, new_n19279_,
    new_n19280_, new_n19281_, new_n19282_, new_n19283_, new_n19284_,
    new_n19285_, new_n19286_, new_n19287_, new_n19288_, new_n19289_,
    new_n19290_, new_n19291_, new_n19292_, new_n19293_, new_n19294_,
    new_n19295_, new_n19296_, new_n19297_, new_n19298_, new_n19299_,
    new_n19300_, new_n19301_, new_n19302_, new_n19303_, new_n19304_,
    new_n19305_, new_n19306_, new_n19307_, new_n19308_, new_n19309_,
    new_n19310_, new_n19311_, new_n19312_, new_n19313_, new_n19314_,
    new_n19315_, new_n19316_, new_n19317_, new_n19318_, new_n19319_,
    new_n19320_, new_n19321_, new_n19322_, new_n19323_, new_n19324_,
    new_n19325_, new_n19326_, new_n19327_, new_n19328_, new_n19329_,
    new_n19330_, new_n19331_, new_n19332_, new_n19333_, new_n19334_,
    new_n19335_, new_n19336_, new_n19337_, new_n19338_, new_n19339_,
    new_n19340_, new_n19341_, new_n19342_, new_n19343_, new_n19344_,
    new_n19345_, new_n19346_, new_n19347_, new_n19348_, new_n19349_,
    new_n19350_, new_n19351_, new_n19352_, new_n19353_, new_n19354_,
    new_n19355_, new_n19356_, new_n19357_, new_n19358_, new_n19359_,
    new_n19360_, new_n19361_, new_n19362_, new_n19363_, new_n19364_,
    new_n19365_, new_n19366_, new_n19367_, new_n19368_, new_n19369_,
    new_n19370_, new_n19371_, new_n19372_, new_n19373_, new_n19374_,
    new_n19375_, new_n19376_, new_n19377_, new_n19378_, new_n19379_,
    new_n19380_, new_n19381_, new_n19382_, new_n19383_, new_n19384_,
    new_n19385_, new_n19386_, new_n19387_, new_n19388_, new_n19389_,
    new_n19390_, new_n19391_, new_n19392_, new_n19393_, new_n19394_,
    new_n19395_, new_n19396_, new_n19397_, new_n19398_, new_n19399_,
    new_n19400_, new_n19401_, new_n19402_, new_n19403_, new_n19404_,
    new_n19405_, new_n19406_, new_n19407_, new_n19408_, new_n19409_,
    new_n19410_, new_n19411_, new_n19412_, new_n19413_, new_n19414_,
    new_n19415_, new_n19416_, new_n19417_, new_n19418_, new_n19419_,
    new_n19420_, new_n19421_, new_n19422_, new_n19423_, new_n19424_,
    new_n19425_, new_n19426_, new_n19427_, new_n19428_, new_n19429_,
    new_n19430_, new_n19431_, new_n19432_, new_n19433_, new_n19434_,
    new_n19435_, new_n19436_, new_n19437_, new_n19438_, new_n19439_,
    new_n19440_, new_n19441_, new_n19442_, new_n19443_, new_n19444_,
    new_n19445_, new_n19446_, new_n19447_, new_n19448_, new_n19449_,
    new_n19450_, new_n19451_, new_n19452_, new_n19453_, new_n19454_,
    new_n19455_, new_n19457_, new_n19458_, new_n19459_, new_n19460_,
    new_n19461_, new_n19462_, new_n19463_, new_n19464_, new_n19465_,
    new_n19466_, new_n19467_, new_n19468_, new_n19469_, new_n19470_,
    new_n19471_, new_n19472_, new_n19473_, new_n19474_, new_n19475_,
    new_n19476_, new_n19477_, new_n19478_, new_n19479_, new_n19480_,
    new_n19481_, new_n19482_, new_n19483_, new_n19484_, new_n19485_,
    new_n19486_, new_n19487_, new_n19488_, new_n19489_, new_n19490_,
    new_n19491_, new_n19492_, new_n19493_, new_n19494_, new_n19495_,
    new_n19496_, new_n19497_, new_n19498_, new_n19499_, new_n19500_,
    new_n19501_, new_n19502_, new_n19503_, new_n19504_, new_n19505_,
    new_n19506_, new_n19507_, new_n19508_, new_n19509_, new_n19510_,
    new_n19511_, new_n19512_, new_n19513_, new_n19514_, new_n19515_,
    new_n19516_, new_n19517_, new_n19518_, new_n19519_, new_n19520_,
    new_n19521_, new_n19522_, new_n19523_, new_n19524_, new_n19525_,
    new_n19526_, new_n19527_, new_n19528_, new_n19529_, new_n19530_,
    new_n19531_, new_n19532_, new_n19533_, new_n19534_, new_n19535_,
    new_n19536_, new_n19537_, new_n19538_, new_n19539_, new_n19540_,
    new_n19541_, new_n19542_, new_n19543_, new_n19544_, new_n19545_,
    new_n19546_, new_n19547_, new_n19548_, new_n19549_, new_n19550_,
    new_n19551_, new_n19552_, new_n19553_, new_n19554_, new_n19555_,
    new_n19556_, new_n19557_, new_n19558_, new_n19559_, new_n19560_,
    new_n19561_, new_n19562_, new_n19563_, new_n19564_, new_n19565_,
    new_n19566_, new_n19567_, new_n19568_, new_n19569_, new_n19570_,
    new_n19571_, new_n19572_, new_n19573_, new_n19574_, new_n19575_,
    new_n19576_, new_n19577_, new_n19578_, new_n19579_, new_n19580_,
    new_n19581_, new_n19582_, new_n19583_, new_n19584_, new_n19585_,
    new_n19586_, new_n19587_, new_n19588_, new_n19589_, new_n19590_,
    new_n19591_, new_n19592_, new_n19593_, new_n19594_, new_n19595_,
    new_n19596_, new_n19597_, new_n19598_, new_n19599_, new_n19600_,
    new_n19601_, new_n19602_, new_n19603_, new_n19604_, new_n19605_,
    new_n19606_, new_n19607_, new_n19608_, new_n19609_, new_n19610_,
    new_n19611_, new_n19612_, new_n19613_, new_n19614_, new_n19615_,
    new_n19616_, new_n19617_, new_n19618_, new_n19619_, new_n19620_,
    new_n19621_, new_n19622_, new_n19623_, new_n19624_, new_n19625_,
    new_n19626_, new_n19627_, new_n19628_, new_n19629_, new_n19630_,
    new_n19631_, new_n19632_, new_n19633_, new_n19634_, new_n19635_,
    new_n19636_, new_n19637_, new_n19638_, new_n19639_, new_n19640_,
    new_n19641_, new_n19642_, new_n19643_, new_n19644_, new_n19645_,
    new_n19646_, new_n19647_, new_n19648_, new_n19649_, new_n19650_,
    new_n19651_, new_n19652_, new_n19653_, new_n19654_, new_n19655_,
    new_n19656_, new_n19657_, new_n19658_, new_n19659_, new_n19660_,
    new_n19661_, new_n19662_, new_n19663_, new_n19664_, new_n19665_,
    new_n19666_, new_n19667_, new_n19668_, new_n19669_, new_n19670_,
    new_n19671_, new_n19672_, new_n19673_, new_n19674_, new_n19675_,
    new_n19676_, new_n19677_, new_n19678_, new_n19679_, new_n19680_,
    new_n19681_, new_n19682_, new_n19683_, new_n19684_, new_n19685_,
    new_n19686_, new_n19687_, new_n19688_, new_n19689_, new_n19690_,
    new_n19691_, new_n19692_, new_n19693_, new_n19694_, new_n19695_,
    new_n19696_, new_n19697_, new_n19698_, new_n19699_, new_n19700_,
    new_n19701_, new_n19702_, new_n19703_, new_n19704_, new_n19705_,
    new_n19706_, new_n19707_, new_n19708_, new_n19709_, new_n19710_,
    new_n19711_, new_n19712_, new_n19713_, new_n19714_, new_n19715_,
    new_n19716_, new_n19717_, new_n19718_, new_n19719_, new_n19720_,
    new_n19721_, new_n19722_, new_n19723_, new_n19724_, new_n19725_,
    new_n19726_, new_n19727_, new_n19728_, new_n19729_, new_n19730_,
    new_n19731_, new_n19732_, new_n19733_, new_n19734_, new_n19736_,
    new_n19737_, new_n19738_, new_n19739_, new_n19740_, new_n19741_,
    new_n19742_, new_n19743_, new_n19744_, new_n19745_, new_n19746_,
    new_n19747_, new_n19748_, new_n19749_, new_n19750_, new_n19751_,
    new_n19752_, new_n19753_, new_n19754_, new_n19755_, new_n19756_,
    new_n19757_, new_n19758_, new_n19759_, new_n19760_, new_n19761_,
    new_n19762_, new_n19763_, new_n19764_, new_n19765_, new_n19766_,
    new_n19767_, new_n19768_, new_n19769_, new_n19770_, new_n19771_,
    new_n19772_, new_n19773_, new_n19774_, new_n19775_, new_n19776_,
    new_n19777_, new_n19778_, new_n19779_, new_n19780_, new_n19781_,
    new_n19782_, new_n19783_, new_n19784_, new_n19785_, new_n19786_,
    new_n19787_, new_n19788_, new_n19789_, new_n19790_, new_n19791_,
    new_n19792_, new_n19793_, new_n19794_, new_n19795_, new_n19796_,
    new_n19797_, new_n19798_, new_n19799_, new_n19800_, new_n19801_,
    new_n19802_, new_n19803_, new_n19804_, new_n19805_, new_n19806_,
    new_n19807_, new_n19808_, new_n19809_, new_n19810_, new_n19811_,
    new_n19812_, new_n19813_, new_n19814_, new_n19815_, new_n19816_,
    new_n19817_, new_n19818_, new_n19819_, new_n19820_, new_n19821_,
    new_n19822_, new_n19823_, new_n19824_, new_n19825_, new_n19826_,
    new_n19827_, new_n19828_, new_n19829_, new_n19830_, new_n19831_,
    new_n19832_, new_n19833_, new_n19834_, new_n19835_, new_n19836_,
    new_n19837_, new_n19838_, new_n19839_, new_n19840_, new_n19841_,
    new_n19842_, new_n19843_, new_n19844_, new_n19845_, new_n19846_,
    new_n19847_, new_n19848_, new_n19849_, new_n19850_, new_n19851_,
    new_n19852_, new_n19853_, new_n19854_, new_n19855_, new_n19856_,
    new_n19857_, new_n19858_, new_n19859_, new_n19860_, new_n19861_,
    new_n19862_, new_n19863_, new_n19864_, new_n19865_, new_n19866_,
    new_n19867_, new_n19868_, new_n19869_, new_n19870_, new_n19871_,
    new_n19872_, new_n19873_, new_n19874_, new_n19875_, new_n19876_,
    new_n19877_, new_n19878_, new_n19879_, new_n19880_, new_n19881_,
    new_n19882_, new_n19883_, new_n19884_, new_n19885_, new_n19886_,
    new_n19887_, new_n19888_, new_n19889_, new_n19890_, new_n19891_,
    new_n19892_, new_n19893_, new_n19894_, new_n19895_, new_n19896_,
    new_n19897_, new_n19898_, new_n19899_, new_n19900_, new_n19901_,
    new_n19902_, new_n19903_, new_n19904_, new_n19905_, new_n19906_,
    new_n19907_, new_n19908_, new_n19909_, new_n19910_, new_n19911_,
    new_n19912_, new_n19913_, new_n19914_, new_n19915_, new_n19916_,
    new_n19917_, new_n19918_, new_n19919_, new_n19920_, new_n19921_,
    new_n19922_, new_n19923_, new_n19924_, new_n19925_, new_n19926_,
    new_n19927_, new_n19928_, new_n19929_, new_n19930_, new_n19931_,
    new_n19932_, new_n19933_, new_n19934_, new_n19935_, new_n19936_,
    new_n19937_, new_n19938_, new_n19939_, new_n19940_, new_n19941_,
    new_n19942_, new_n19943_, new_n19944_, new_n19945_, new_n19946_,
    new_n19947_, new_n19948_, new_n19949_, new_n19950_, new_n19951_,
    new_n19952_, new_n19953_, new_n19954_, new_n19955_, new_n19956_,
    new_n19957_, new_n19958_, new_n19959_, new_n19960_, new_n19961_,
    new_n19962_, new_n19963_, new_n19964_, new_n19965_, new_n19966_,
    new_n19967_, new_n19968_, new_n19969_, new_n19970_, new_n19971_,
    new_n19972_, new_n19973_, new_n19974_, new_n19975_, new_n19976_,
    new_n19977_, new_n19978_, new_n19979_, new_n19980_, new_n19981_,
    new_n19982_, new_n19983_, new_n19984_, new_n19985_, new_n19986_,
    new_n19987_, new_n19988_, new_n19989_, new_n19990_, new_n19991_,
    new_n19992_, new_n19993_, new_n19994_, new_n19995_, new_n19996_,
    new_n19997_, new_n19998_, new_n19999_, new_n20000_, new_n20001_,
    new_n20002_, new_n20003_, new_n20004_, new_n20005_, new_n20006_,
    new_n20007_, new_n20008_, new_n20009_, new_n20010_, new_n20011_,
    new_n20012_, new_n20013_, new_n20015_, new_n20016_, new_n20017_,
    new_n20018_, new_n20019_, new_n20020_, new_n20021_, new_n20022_,
    new_n20023_, new_n20024_, new_n20025_, new_n20026_, new_n20027_,
    new_n20028_, new_n20029_, new_n20030_, new_n20031_, new_n20032_,
    new_n20033_, new_n20034_, new_n20035_, new_n20036_, new_n20037_,
    new_n20038_, new_n20039_, new_n20040_, new_n20041_, new_n20042_,
    new_n20043_, new_n20044_, new_n20045_, new_n20046_, new_n20047_,
    new_n20048_, new_n20049_, new_n20050_, new_n20051_, new_n20052_,
    new_n20053_, new_n20054_, new_n20055_, new_n20056_, new_n20057_,
    new_n20058_, new_n20059_, new_n20060_, new_n20061_, new_n20062_,
    new_n20063_, new_n20064_, new_n20065_, new_n20066_, new_n20067_,
    new_n20068_, new_n20069_, new_n20070_, new_n20071_, new_n20072_,
    new_n20073_, new_n20074_, new_n20075_, new_n20076_, new_n20077_,
    new_n20078_, new_n20079_, new_n20080_, new_n20081_, new_n20082_,
    new_n20083_, new_n20084_, new_n20085_, new_n20086_, new_n20087_,
    new_n20088_, new_n20089_, new_n20090_, new_n20091_, new_n20092_,
    new_n20093_, new_n20094_, new_n20095_, new_n20096_, new_n20097_,
    new_n20098_, new_n20099_, new_n20100_, new_n20101_, new_n20102_,
    new_n20103_, new_n20104_, new_n20105_, new_n20106_, new_n20107_,
    new_n20108_, new_n20109_, new_n20110_, new_n20111_, new_n20112_,
    new_n20113_, new_n20114_, new_n20115_, new_n20116_, new_n20117_,
    new_n20118_, new_n20119_, new_n20120_, new_n20121_, new_n20122_,
    new_n20123_, new_n20124_, new_n20125_, new_n20126_, new_n20127_,
    new_n20128_, new_n20129_, new_n20130_, new_n20131_, new_n20132_,
    new_n20133_, new_n20134_, new_n20135_, new_n20136_, new_n20137_,
    new_n20138_, new_n20139_, new_n20140_, new_n20141_, new_n20142_,
    new_n20143_, new_n20144_, new_n20145_, new_n20146_, new_n20147_,
    new_n20148_, new_n20149_, new_n20150_, new_n20151_, new_n20152_,
    new_n20153_, new_n20154_, new_n20155_, new_n20156_, new_n20157_,
    new_n20158_, new_n20159_, new_n20160_, new_n20161_, new_n20162_,
    new_n20163_, new_n20164_, new_n20165_, new_n20166_, new_n20167_,
    new_n20168_, new_n20169_, new_n20170_, new_n20171_, new_n20172_,
    new_n20173_, new_n20174_, new_n20175_, new_n20176_, new_n20177_,
    new_n20178_, new_n20179_, new_n20180_, new_n20181_, new_n20182_,
    new_n20183_, new_n20184_, new_n20185_, new_n20186_, new_n20187_,
    new_n20188_, new_n20189_, new_n20190_, new_n20191_, new_n20192_,
    new_n20193_, new_n20194_, new_n20195_, new_n20196_, new_n20197_,
    new_n20198_, new_n20199_, new_n20200_, new_n20201_, new_n20202_,
    new_n20203_, new_n20204_, new_n20205_, new_n20206_, new_n20207_,
    new_n20208_, new_n20209_, new_n20210_, new_n20211_, new_n20212_,
    new_n20213_, new_n20214_, new_n20215_, new_n20216_, new_n20217_,
    new_n20218_, new_n20219_, new_n20220_, new_n20221_, new_n20222_,
    new_n20223_, new_n20224_, new_n20225_, new_n20226_, new_n20227_,
    new_n20228_, new_n20229_, new_n20230_, new_n20231_, new_n20232_,
    new_n20233_, new_n20234_, new_n20235_, new_n20236_, new_n20237_,
    new_n20238_, new_n20239_, new_n20240_, new_n20241_, new_n20242_,
    new_n20243_, new_n20244_, new_n20245_, new_n20246_, new_n20247_,
    new_n20248_, new_n20249_, new_n20250_, new_n20251_, new_n20252_,
    new_n20253_, new_n20254_, new_n20255_, new_n20256_, new_n20257_,
    new_n20258_, new_n20259_, new_n20260_, new_n20261_, new_n20262_,
    new_n20263_, new_n20264_, new_n20265_, new_n20266_, new_n20267_,
    new_n20268_, new_n20269_, new_n20270_, new_n20271_, new_n20272_,
    new_n20273_, new_n20274_, new_n20275_, new_n20276_, new_n20277_,
    new_n20278_, new_n20279_, new_n20280_, new_n20281_, new_n20282_,
    new_n20283_, new_n20284_, new_n20285_, new_n20286_, new_n20287_,
    new_n20288_, new_n20289_, new_n20291_, new_n20292_, new_n20293_,
    new_n20294_, new_n20295_, new_n20296_, new_n20297_, new_n20298_,
    new_n20299_, new_n20300_, new_n20301_, new_n20302_, new_n20303_,
    new_n20304_, new_n20305_, new_n20306_, new_n20307_, new_n20308_,
    new_n20309_, new_n20310_, new_n20311_, new_n20312_, new_n20313_,
    new_n20314_, new_n20315_, new_n20316_, new_n20317_, new_n20318_,
    new_n20319_, new_n20320_, new_n20321_, new_n20322_, new_n20323_,
    new_n20324_, new_n20325_, new_n20326_, new_n20327_, new_n20328_,
    new_n20329_, new_n20330_, new_n20331_, new_n20332_, new_n20333_,
    new_n20334_, new_n20335_, new_n20336_, new_n20337_, new_n20338_,
    new_n20339_, new_n20340_, new_n20341_, new_n20342_, new_n20343_,
    new_n20344_, new_n20345_, new_n20346_, new_n20347_, new_n20348_,
    new_n20349_, new_n20350_, new_n20351_, new_n20352_, new_n20353_,
    new_n20354_, new_n20355_, new_n20356_, new_n20357_, new_n20358_,
    new_n20359_, new_n20360_, new_n20361_, new_n20362_, new_n20363_,
    new_n20364_, new_n20365_, new_n20366_, new_n20367_, new_n20368_,
    new_n20369_, new_n20370_, new_n20371_, new_n20372_, new_n20373_,
    new_n20374_, new_n20375_, new_n20376_, new_n20377_, new_n20378_,
    new_n20379_, new_n20380_, new_n20381_, new_n20382_, new_n20383_,
    new_n20384_, new_n20385_, new_n20386_, new_n20387_, new_n20388_,
    new_n20389_, new_n20390_, new_n20391_, new_n20392_, new_n20393_,
    new_n20394_, new_n20395_, new_n20396_, new_n20397_, new_n20398_,
    new_n20399_, new_n20400_, new_n20401_, new_n20402_, new_n20403_,
    new_n20404_, new_n20405_, new_n20406_, new_n20407_, new_n20408_,
    new_n20409_, new_n20410_, new_n20411_, new_n20412_, new_n20413_,
    new_n20414_, new_n20415_, new_n20416_, new_n20417_, new_n20418_,
    new_n20419_, new_n20420_, new_n20421_, new_n20422_, new_n20423_,
    new_n20424_, new_n20425_, new_n20426_, new_n20427_, new_n20428_,
    new_n20429_, new_n20430_, new_n20431_, new_n20432_, new_n20433_,
    new_n20434_, new_n20435_, new_n20436_, new_n20437_, new_n20438_,
    new_n20439_, new_n20440_, new_n20441_, new_n20442_, new_n20443_,
    new_n20444_, new_n20445_, new_n20446_, new_n20447_, new_n20448_,
    new_n20449_, new_n20450_, new_n20451_, new_n20452_, new_n20453_,
    new_n20454_, new_n20455_, new_n20456_, new_n20457_, new_n20458_,
    new_n20459_, new_n20460_, new_n20461_, new_n20462_, new_n20463_,
    new_n20464_, new_n20465_, new_n20466_, new_n20467_, new_n20468_,
    new_n20469_, new_n20470_, new_n20471_, new_n20472_, new_n20473_,
    new_n20474_, new_n20475_, new_n20476_, new_n20477_, new_n20478_,
    new_n20479_, new_n20480_, new_n20481_, new_n20482_, new_n20483_,
    new_n20484_, new_n20485_, new_n20486_, new_n20487_, new_n20488_,
    new_n20489_, new_n20490_, new_n20491_, new_n20492_, new_n20493_,
    new_n20494_, new_n20495_, new_n20496_, new_n20497_, new_n20498_,
    new_n20499_, new_n20500_, new_n20501_, new_n20502_, new_n20503_,
    new_n20504_, new_n20505_, new_n20506_, new_n20507_, new_n20508_,
    new_n20509_, new_n20510_, new_n20511_, new_n20512_, new_n20513_,
    new_n20514_, new_n20515_, new_n20516_, new_n20517_, new_n20518_,
    new_n20519_, new_n20520_, new_n20521_, new_n20522_, new_n20523_,
    new_n20524_, new_n20525_, new_n20526_, new_n20527_, new_n20528_,
    new_n20529_, new_n20530_, new_n20531_, new_n20532_, new_n20533_,
    new_n20534_, new_n20535_, new_n20536_, new_n20537_, new_n20538_,
    new_n20539_, new_n20540_, new_n20541_, new_n20542_, new_n20543_,
    new_n20544_, new_n20545_, new_n20546_, new_n20547_, new_n20548_,
    new_n20549_, new_n20550_, new_n20551_, new_n20552_, new_n20553_,
    new_n20554_, new_n20555_, new_n20556_, new_n20557_, new_n20558_,
    new_n20559_, new_n20560_, new_n20561_, new_n20562_, new_n20564_,
    new_n20565_, new_n20566_, new_n20567_, new_n20568_, new_n20569_,
    new_n20570_, new_n20571_, new_n20572_, new_n20573_, new_n20574_,
    new_n20575_, new_n20576_, new_n20577_, new_n20578_, new_n20579_,
    new_n20580_, new_n20581_, new_n20582_, new_n20583_, new_n20584_,
    new_n20585_, new_n20586_, new_n20587_, new_n20588_, new_n20589_,
    new_n20590_, new_n20591_, new_n20592_, new_n20593_, new_n20594_,
    new_n20595_, new_n20596_, new_n20597_, new_n20598_, new_n20599_,
    new_n20600_, new_n20601_, new_n20602_, new_n20603_, new_n20604_,
    new_n20605_, new_n20606_, new_n20607_, new_n20608_, new_n20609_,
    new_n20610_, new_n20611_, new_n20612_, new_n20613_, new_n20614_,
    new_n20615_, new_n20616_, new_n20617_, new_n20618_, new_n20619_,
    new_n20620_, new_n20621_, new_n20622_, new_n20623_, new_n20624_,
    new_n20625_, new_n20626_, new_n20627_, new_n20628_, new_n20629_,
    new_n20630_, new_n20631_, new_n20632_, new_n20633_, new_n20634_,
    new_n20635_, new_n20636_, new_n20637_, new_n20638_, new_n20639_,
    new_n20640_, new_n20641_, new_n20642_, new_n20643_, new_n20644_,
    new_n20645_, new_n20646_, new_n20647_, new_n20648_, new_n20649_,
    new_n20650_, new_n20651_, new_n20652_, new_n20653_, new_n20654_,
    new_n20655_, new_n20656_, new_n20657_, new_n20658_, new_n20659_,
    new_n20660_, new_n20661_, new_n20662_, new_n20663_, new_n20664_,
    new_n20665_, new_n20666_, new_n20667_, new_n20668_, new_n20669_,
    new_n20670_, new_n20671_, new_n20672_, new_n20673_, new_n20674_,
    new_n20675_, new_n20676_, new_n20677_, new_n20678_, new_n20679_,
    new_n20680_, new_n20681_, new_n20682_, new_n20683_, new_n20684_,
    new_n20685_, new_n20686_, new_n20687_, new_n20688_, new_n20689_,
    new_n20690_, new_n20691_, new_n20692_, new_n20693_, new_n20694_,
    new_n20695_, new_n20696_, new_n20697_, new_n20698_, new_n20699_,
    new_n20700_, new_n20701_, new_n20702_, new_n20703_, new_n20704_,
    new_n20705_, new_n20706_, new_n20707_, new_n20708_, new_n20709_,
    new_n20710_, new_n20711_, new_n20712_, new_n20713_, new_n20714_,
    new_n20715_, new_n20716_, new_n20717_, new_n20718_, new_n20719_,
    new_n20720_, new_n20721_, new_n20722_, new_n20723_, new_n20724_,
    new_n20725_, new_n20726_, new_n20727_, new_n20728_, new_n20729_,
    new_n20730_, new_n20731_, new_n20732_, new_n20733_, new_n20734_,
    new_n20735_, new_n20736_, new_n20737_, new_n20738_, new_n20739_,
    new_n20740_, new_n20741_, new_n20742_, new_n20743_, new_n20744_,
    new_n20745_, new_n20746_, new_n20747_, new_n20748_, new_n20749_,
    new_n20750_, new_n20751_, new_n20752_, new_n20753_, new_n20754_,
    new_n20755_, new_n20756_, new_n20757_, new_n20758_, new_n20759_,
    new_n20760_, new_n20761_, new_n20762_, new_n20763_, new_n20764_,
    new_n20765_, new_n20766_, new_n20767_, new_n20768_, new_n20769_,
    new_n20770_, new_n20771_, new_n20772_, new_n20773_, new_n20774_,
    new_n20775_, new_n20776_, new_n20777_, new_n20778_, new_n20779_,
    new_n20780_, new_n20781_, new_n20782_, new_n20783_, new_n20784_,
    new_n20785_, new_n20786_, new_n20787_, new_n20788_, new_n20789_,
    new_n20790_, new_n20791_, new_n20792_, new_n20793_, new_n20794_,
    new_n20795_, new_n20796_, new_n20797_, new_n20798_, new_n20799_,
    new_n20800_, new_n20801_, new_n20802_, new_n20803_, new_n20804_,
    new_n20805_, new_n20806_, new_n20807_, new_n20808_, new_n20809_,
    new_n20810_, new_n20811_, new_n20812_, new_n20813_, new_n20814_,
    new_n20815_, new_n20816_, new_n20817_, new_n20818_, new_n20819_,
    new_n20820_, new_n20821_, new_n20822_, new_n20823_, new_n20824_,
    new_n20825_, new_n20826_, new_n20827_, new_n20828_, new_n20829_,
    new_n20830_, new_n20831_, new_n20832_, new_n20833_, new_n20834_,
    new_n20835_, new_n20837_, new_n20838_, new_n20839_, new_n20840_,
    new_n20841_, new_n20842_, new_n20843_, new_n20844_, new_n20845_,
    new_n20846_, new_n20847_, new_n20848_, new_n20849_, new_n20850_,
    new_n20851_, new_n20852_, new_n20853_, new_n20854_, new_n20855_,
    new_n20856_, new_n20857_, new_n20858_, new_n20859_, new_n20860_,
    new_n20861_, new_n20862_, new_n20863_, new_n20864_, new_n20865_,
    new_n20866_, new_n20867_, new_n20868_, new_n20869_, new_n20870_,
    new_n20871_, new_n20872_, new_n20873_, new_n20874_, new_n20875_,
    new_n20876_, new_n20877_, new_n20878_, new_n20879_, new_n20880_,
    new_n20881_, new_n20882_, new_n20883_, new_n20884_, new_n20885_,
    new_n20886_, new_n20887_, new_n20888_, new_n20889_, new_n20890_,
    new_n20891_, new_n20892_, new_n20893_, new_n20894_, new_n20895_,
    new_n20896_, new_n20897_, new_n20898_, new_n20899_, new_n20900_,
    new_n20901_, new_n20902_, new_n20903_, new_n20904_, new_n20905_,
    new_n20906_, new_n20907_, new_n20908_, new_n20909_, new_n20910_,
    new_n20911_, new_n20912_, new_n20913_, new_n20914_, new_n20915_,
    new_n20916_, new_n20917_, new_n20918_, new_n20919_, new_n20920_,
    new_n20921_, new_n20922_, new_n20923_, new_n20924_, new_n20925_,
    new_n20926_, new_n20927_, new_n20928_, new_n20929_, new_n20930_,
    new_n20931_, new_n20932_, new_n20933_, new_n20934_, new_n20935_,
    new_n20936_, new_n20937_, new_n20938_, new_n20939_, new_n20940_,
    new_n20941_, new_n20942_, new_n20943_, new_n20944_, new_n20945_,
    new_n20946_, new_n20947_, new_n20948_, new_n20949_, new_n20950_,
    new_n20951_, new_n20952_, new_n20953_, new_n20954_, new_n20955_,
    new_n20956_, new_n20957_, new_n20958_, new_n20959_, new_n20960_,
    new_n20961_, new_n20962_, new_n20963_, new_n20964_, new_n20965_,
    new_n20966_, new_n20967_, new_n20968_, new_n20969_, new_n20970_,
    new_n20971_, new_n20972_, new_n20973_, new_n20974_, new_n20975_,
    new_n20976_, new_n20977_, new_n20978_, new_n20979_, new_n20980_,
    new_n20981_, new_n20982_, new_n20983_, new_n20984_, new_n20985_,
    new_n20986_, new_n20987_, new_n20988_, new_n20989_, new_n20990_,
    new_n20991_, new_n20992_, new_n20993_, new_n20994_, new_n20995_,
    new_n20996_, new_n20997_, new_n20998_, new_n20999_, new_n21000_,
    new_n21001_, new_n21002_, new_n21003_, new_n21004_, new_n21005_,
    new_n21006_, new_n21007_, new_n21008_, new_n21009_, new_n21010_,
    new_n21011_, new_n21012_, new_n21013_, new_n21014_, new_n21015_,
    new_n21016_, new_n21017_, new_n21018_, new_n21019_, new_n21020_,
    new_n21021_, new_n21022_, new_n21023_, new_n21024_, new_n21025_,
    new_n21026_, new_n21027_, new_n21028_, new_n21029_, new_n21030_,
    new_n21031_, new_n21032_, new_n21033_, new_n21034_, new_n21035_,
    new_n21036_, new_n21037_, new_n21038_, new_n21039_, new_n21040_,
    new_n21041_, new_n21042_, new_n21043_, new_n21044_, new_n21045_,
    new_n21046_, new_n21047_, new_n21048_, new_n21049_, new_n21050_,
    new_n21051_, new_n21052_, new_n21053_, new_n21054_, new_n21055_,
    new_n21056_, new_n21057_, new_n21058_, new_n21059_, new_n21060_,
    new_n21061_, new_n21062_, new_n21063_, new_n21064_, new_n21065_,
    new_n21066_, new_n21067_, new_n21068_, new_n21069_, new_n21070_,
    new_n21071_, new_n21072_, new_n21073_, new_n21074_, new_n21075_,
    new_n21076_, new_n21077_, new_n21078_, new_n21079_, new_n21080_,
    new_n21081_, new_n21082_, new_n21083_, new_n21084_, new_n21085_,
    new_n21086_, new_n21087_, new_n21088_, new_n21089_, new_n21090_,
    new_n21091_, new_n21092_, new_n21093_, new_n21094_, new_n21095_,
    new_n21096_, new_n21097_, new_n21098_, new_n21099_, new_n21100_,
    new_n21101_, new_n21102_, new_n21103_, new_n21104_, new_n21105_,
    new_n21106_, new_n21107_, new_n21108_, new_n21110_, new_n21111_,
    new_n21112_, new_n21113_, new_n21114_, new_n21115_, new_n21116_,
    new_n21117_, new_n21118_, new_n21119_, new_n21120_, new_n21121_,
    new_n21122_, new_n21123_, new_n21124_, new_n21125_, new_n21126_,
    new_n21127_, new_n21128_, new_n21129_, new_n21130_, new_n21131_,
    new_n21132_, new_n21133_, new_n21134_, new_n21135_, new_n21136_,
    new_n21137_, new_n21138_, new_n21139_, new_n21140_, new_n21141_,
    new_n21142_, new_n21143_, new_n21144_, new_n21145_, new_n21146_,
    new_n21147_, new_n21148_, new_n21149_, new_n21150_, new_n21151_,
    new_n21152_, new_n21153_, new_n21154_, new_n21155_, new_n21156_,
    new_n21157_, new_n21158_, new_n21159_, new_n21160_, new_n21161_,
    new_n21162_, new_n21163_, new_n21164_, new_n21165_, new_n21166_,
    new_n21167_, new_n21168_, new_n21169_, new_n21170_, new_n21171_,
    new_n21172_, new_n21173_, new_n21174_, new_n21175_, new_n21176_,
    new_n21177_, new_n21178_, new_n21179_, new_n21180_, new_n21181_,
    new_n21182_, new_n21183_, new_n21184_, new_n21185_, new_n21186_,
    new_n21187_, new_n21188_, new_n21189_, new_n21190_, new_n21191_,
    new_n21192_, new_n21193_, new_n21194_, new_n21195_, new_n21196_,
    new_n21197_, new_n21198_, new_n21199_, new_n21200_, new_n21201_,
    new_n21202_, new_n21203_, new_n21204_, new_n21205_, new_n21206_,
    new_n21207_, new_n21208_, new_n21209_, new_n21210_, new_n21211_,
    new_n21212_, new_n21213_, new_n21214_, new_n21215_, new_n21216_,
    new_n21217_, new_n21218_, new_n21219_, new_n21220_, new_n21221_,
    new_n21222_, new_n21223_, new_n21224_, new_n21225_, new_n21226_,
    new_n21227_, new_n21228_, new_n21229_, new_n21230_, new_n21231_,
    new_n21232_, new_n21233_, new_n21234_, new_n21235_, new_n21236_,
    new_n21237_, new_n21238_, new_n21239_, new_n21240_, new_n21241_,
    new_n21242_, new_n21243_, new_n21244_, new_n21245_, new_n21246_,
    new_n21247_, new_n21248_, new_n21249_, new_n21250_, new_n21251_,
    new_n21252_, new_n21253_, new_n21254_, new_n21255_, new_n21256_,
    new_n21257_, new_n21258_, new_n21259_, new_n21260_, new_n21261_,
    new_n21262_, new_n21263_, new_n21264_, new_n21265_, new_n21266_,
    new_n21267_, new_n21268_, new_n21269_, new_n21270_, new_n21271_,
    new_n21272_, new_n21273_, new_n21274_, new_n21275_, new_n21276_,
    new_n21277_, new_n21278_, new_n21279_, new_n21280_, new_n21281_,
    new_n21282_, new_n21283_, new_n21284_, new_n21285_, new_n21286_,
    new_n21287_, new_n21288_, new_n21289_, new_n21290_, new_n21291_,
    new_n21292_, new_n21293_, new_n21294_, new_n21295_, new_n21296_,
    new_n21297_, new_n21298_, new_n21299_, new_n21300_, new_n21301_,
    new_n21302_, new_n21303_, new_n21304_, new_n21305_, new_n21306_,
    new_n21307_, new_n21308_, new_n21309_, new_n21310_, new_n21311_,
    new_n21312_, new_n21313_, new_n21314_, new_n21315_, new_n21316_,
    new_n21317_, new_n21318_, new_n21319_, new_n21320_, new_n21321_,
    new_n21322_, new_n21323_, new_n21324_, new_n21325_, new_n21326_,
    new_n21327_, new_n21328_, new_n21329_, new_n21330_, new_n21331_,
    new_n21332_, new_n21333_, new_n21334_, new_n21335_, new_n21336_,
    new_n21337_, new_n21338_, new_n21339_, new_n21340_, new_n21341_,
    new_n21342_, new_n21343_, new_n21344_, new_n21345_, new_n21346_,
    new_n21347_, new_n21348_, new_n21349_, new_n21350_, new_n21351_,
    new_n21352_, new_n21353_, new_n21354_, new_n21355_, new_n21356_,
    new_n21357_, new_n21358_, new_n21359_, new_n21360_, new_n21361_,
    new_n21362_, new_n21363_, new_n21364_, new_n21365_, new_n21366_,
    new_n21367_, new_n21368_, new_n21369_, new_n21370_, new_n21371_,
    new_n21372_, new_n21373_, new_n21374_, new_n21375_, new_n21376_,
    new_n21378_, new_n21379_, new_n21380_, new_n21381_, new_n21382_,
    new_n21383_, new_n21384_, new_n21385_, new_n21386_, new_n21387_,
    new_n21388_, new_n21389_, new_n21390_, new_n21391_, new_n21392_,
    new_n21393_, new_n21394_, new_n21395_, new_n21396_, new_n21397_,
    new_n21398_, new_n21399_, new_n21400_, new_n21401_, new_n21402_,
    new_n21403_, new_n21404_, new_n21405_, new_n21406_, new_n21407_,
    new_n21408_, new_n21409_, new_n21410_, new_n21411_, new_n21412_,
    new_n21413_, new_n21414_, new_n21415_, new_n21416_, new_n21417_,
    new_n21418_, new_n21419_, new_n21420_, new_n21421_, new_n21422_,
    new_n21423_, new_n21424_, new_n21425_, new_n21426_, new_n21427_,
    new_n21428_, new_n21429_, new_n21430_, new_n21431_, new_n21432_,
    new_n21433_, new_n21434_, new_n21435_, new_n21436_, new_n21437_,
    new_n21438_, new_n21439_, new_n21440_, new_n21441_, new_n21442_,
    new_n21443_, new_n21444_, new_n21445_, new_n21446_, new_n21447_,
    new_n21448_, new_n21449_, new_n21450_, new_n21451_, new_n21452_,
    new_n21453_, new_n21454_, new_n21455_, new_n21456_, new_n21457_,
    new_n21458_, new_n21459_, new_n21460_, new_n21461_, new_n21462_,
    new_n21463_, new_n21464_, new_n21465_, new_n21466_, new_n21467_,
    new_n21468_, new_n21469_, new_n21470_, new_n21471_, new_n21472_,
    new_n21473_, new_n21474_, new_n21475_, new_n21476_, new_n21477_,
    new_n21478_, new_n21479_, new_n21480_, new_n21481_, new_n21482_,
    new_n21483_, new_n21484_, new_n21485_, new_n21486_, new_n21487_,
    new_n21488_, new_n21489_, new_n21490_, new_n21491_, new_n21492_,
    new_n21493_, new_n21494_, new_n21495_, new_n21496_, new_n21497_,
    new_n21498_, new_n21499_, new_n21500_, new_n21501_, new_n21502_,
    new_n21503_, new_n21504_, new_n21505_, new_n21506_, new_n21507_,
    new_n21508_, new_n21509_, new_n21510_, new_n21511_, new_n21512_,
    new_n21513_, new_n21514_, new_n21515_, new_n21516_, new_n21517_,
    new_n21518_, new_n21519_, new_n21520_, new_n21521_, new_n21522_,
    new_n21523_, new_n21524_, new_n21525_, new_n21526_, new_n21527_,
    new_n21528_, new_n21529_, new_n21530_, new_n21531_, new_n21532_,
    new_n21533_, new_n21534_, new_n21535_, new_n21536_, new_n21537_,
    new_n21538_, new_n21539_, new_n21540_, new_n21541_, new_n21542_,
    new_n21543_, new_n21544_, new_n21545_, new_n21546_, new_n21547_,
    new_n21548_, new_n21549_, new_n21550_, new_n21551_, new_n21552_,
    new_n21553_, new_n21554_, new_n21555_, new_n21556_, new_n21557_,
    new_n21558_, new_n21559_, new_n21560_, new_n21561_, new_n21562_,
    new_n21563_, new_n21564_, new_n21565_, new_n21566_, new_n21567_,
    new_n21568_, new_n21569_, new_n21570_, new_n21571_, new_n21572_,
    new_n21573_, new_n21574_, new_n21575_, new_n21576_, new_n21577_,
    new_n21578_, new_n21579_, new_n21580_, new_n21581_, new_n21582_,
    new_n21583_, new_n21584_, new_n21585_, new_n21586_, new_n21587_,
    new_n21588_, new_n21589_, new_n21590_, new_n21591_, new_n21592_,
    new_n21593_, new_n21594_, new_n21595_, new_n21596_, new_n21597_,
    new_n21598_, new_n21599_, new_n21600_, new_n21601_, new_n21602_,
    new_n21603_, new_n21604_, new_n21605_, new_n21606_, new_n21607_,
    new_n21608_, new_n21609_, new_n21610_, new_n21611_, new_n21612_,
    new_n21613_, new_n21614_, new_n21615_, new_n21616_, new_n21617_,
    new_n21618_, new_n21619_, new_n21620_, new_n21621_, new_n21622_,
    new_n21623_, new_n21624_, new_n21625_, new_n21626_, new_n21627_,
    new_n21628_, new_n21629_, new_n21630_, new_n21631_, new_n21632_,
    new_n21633_, new_n21634_, new_n21635_, new_n21636_, new_n21637_,
    new_n21639_, new_n21640_, new_n21641_, new_n21642_, new_n21643_,
    new_n21644_, new_n21645_, new_n21646_, new_n21647_, new_n21648_,
    new_n21649_, new_n21650_, new_n21651_, new_n21652_, new_n21653_,
    new_n21654_, new_n21655_, new_n21656_, new_n21657_, new_n21658_,
    new_n21659_, new_n21660_, new_n21661_, new_n21662_, new_n21663_,
    new_n21664_, new_n21665_, new_n21667_, new_n21668_, new_n21669_,
    new_n21670_, new_n21671_, new_n21672_, new_n21673_, new_n21674_,
    new_n21675_, new_n21676_, new_n21677_, new_n21678_, new_n21679_,
    new_n21680_, new_n21681_, new_n21682_, new_n21683_, new_n21684_,
    new_n21685_, new_n21686_, new_n21687_, new_n21688_, new_n21689_,
    new_n21690_, new_n21691_, new_n21692_, new_n21693_, new_n21694_,
    new_n21695_, new_n21696_, new_n21697_, new_n21698_, new_n21699_,
    new_n21700_, new_n21701_, new_n21702_, new_n21703_, new_n21704_,
    new_n21705_, new_n21706_, new_n21707_, new_n21708_, new_n21709_,
    new_n21710_, new_n21711_, new_n21712_, new_n21714_, new_n21715_,
    new_n21716_, new_n21717_, new_n21718_, new_n21719_, new_n21720_,
    new_n21721_, new_n21722_, new_n21723_, new_n21724_, new_n21725_,
    new_n21726_, new_n21727_, new_n21728_, new_n21729_, new_n21730_,
    new_n21731_, new_n21732_, new_n21733_, new_n21734_, new_n21735_,
    new_n21736_, new_n21737_, new_n21738_, new_n21739_, new_n21740_,
    new_n21741_, new_n21742_, new_n21743_, new_n21744_, new_n21745_,
    new_n21746_, new_n21747_, new_n21749_, new_n21750_, new_n21751_,
    new_n21752_, new_n21753_, new_n21754_, new_n21755_, new_n21756_,
    new_n21757_, new_n21758_, new_n21759_, new_n21760_, new_n21761_,
    new_n21762_, new_n21763_, new_n21764_, new_n21765_, new_n21766_,
    new_n21767_, new_n21768_, new_n21769_, new_n21770_, new_n21771_,
    new_n21772_, new_n21773_, new_n21774_, new_n21775_, new_n21776_,
    new_n21777_, new_n21778_, new_n21779_, new_n21780_, new_n21781_,
    new_n21782_, new_n21783_, new_n21784_, new_n21785_, new_n21786_,
    new_n21787_, new_n21788_, new_n21789_, new_n21790_, new_n21791_,
    new_n21792_, new_n21793_, new_n21794_, new_n21795_, new_n21796_,
    new_n21797_, new_n21798_, new_n21799_, new_n21800_, new_n21801_,
    new_n21802_, new_n21803_, new_n21804_, new_n21805_, new_n21806_,
    new_n21807_, new_n21808_, new_n21809_, new_n21810_, new_n21811_,
    new_n21812_, new_n21813_, new_n21814_, new_n21815_, new_n21816_,
    new_n21817_, new_n21818_, new_n21819_, new_n21820_, new_n21821_,
    new_n21822_, new_n21823_, new_n21824_, new_n21825_, new_n21826_,
    new_n21827_, new_n21828_, new_n21829_, new_n21830_, new_n21831_,
    new_n21832_, new_n21833_, new_n21834_, new_n21835_, new_n21836_,
    new_n21837_, new_n21838_, new_n21839_, new_n21840_, new_n21841_,
    new_n21842_, new_n21843_, new_n21844_, new_n21845_, new_n21846_,
    new_n21847_, new_n21848_, new_n21849_, new_n21850_, new_n21851_,
    new_n21852_, new_n21853_, new_n21854_, new_n21855_, new_n21856_,
    new_n21857_, new_n21858_, new_n21859_, new_n21860_, new_n21861_,
    new_n21862_, new_n21863_, new_n21864_, new_n21865_, new_n21866_,
    new_n21867_, new_n21868_, new_n21869_, new_n21870_, new_n21871_,
    new_n21872_, new_n21873_, new_n21874_, new_n21875_, new_n21876_,
    new_n21877_, new_n21878_, new_n21879_, new_n21880_, new_n21881_,
    new_n21882_, new_n21883_, new_n21884_, new_n21885_, new_n21886_,
    new_n21887_, new_n21888_, new_n21889_, new_n21890_, new_n21891_,
    new_n21892_, new_n21893_, new_n21894_, new_n21895_, new_n21896_,
    new_n21897_, new_n21898_, new_n21899_, new_n21900_, new_n21901_,
    new_n21902_, new_n21903_, new_n21904_, new_n21905_, new_n21906_,
    new_n21907_, new_n21908_, new_n21909_, new_n21910_, new_n21911_,
    new_n21912_, new_n21913_, new_n21914_, new_n21915_, new_n21916_,
    new_n21917_, new_n21918_, new_n21919_, new_n21920_, new_n21921_,
    new_n21922_, new_n21923_, new_n21924_, new_n21925_, new_n21926_,
    new_n21927_, new_n21928_, new_n21929_, new_n21930_, new_n21931_,
    new_n21932_, new_n21933_, new_n21934_, new_n21935_, new_n21936_,
    new_n21937_, new_n21938_, new_n21939_, new_n21940_, new_n21941_,
    new_n21942_, new_n21943_, new_n21944_, new_n21945_, new_n21946_,
    new_n21947_, new_n21948_, new_n21949_, new_n21950_, new_n21951_,
    new_n21952_, new_n21953_, new_n21954_, new_n21955_, new_n21956_,
    new_n21957_, new_n21958_, new_n21959_, new_n21960_, new_n21961_,
    new_n21962_, new_n21963_, new_n21964_, new_n21965_, new_n21966_,
    new_n21967_, new_n21968_, new_n21969_, new_n21970_, new_n21971_,
    new_n21972_, new_n21973_, new_n21974_, new_n21975_, new_n21976_,
    new_n21977_, new_n21978_, new_n21979_, new_n21980_, new_n21981_,
    new_n21982_, new_n21983_, new_n21984_, new_n21985_, new_n21986_,
    new_n21987_, new_n21988_, new_n21989_, new_n21990_, new_n21991_,
    new_n21992_, new_n21993_, new_n21994_, new_n21995_, new_n21996_,
    new_n21997_, new_n21998_, new_n21999_, new_n22000_, new_n22001_,
    new_n22002_, new_n22003_, new_n22004_, new_n22005_, new_n22006_,
    new_n22007_, new_n22008_, new_n22009_, new_n22010_, new_n22011_,
    new_n22012_, new_n22013_, new_n22014_, new_n22015_, new_n22016_,
    new_n22017_, new_n22018_, new_n22019_, new_n22020_, new_n22021_,
    new_n22022_, new_n22023_, new_n22024_, new_n22025_, new_n22026_,
    new_n22027_, new_n22028_, new_n22029_, new_n22030_, new_n22031_,
    new_n22032_, new_n22033_, new_n22034_, new_n22035_, new_n22036_,
    new_n22037_, new_n22038_, new_n22039_, new_n22040_, new_n22041_,
    new_n22042_, new_n22043_, new_n22044_, new_n22045_, new_n22046_,
    new_n22047_, new_n22048_, new_n22049_, new_n22050_, new_n22051_,
    new_n22052_, new_n22053_, new_n22054_, new_n22055_, new_n22056_,
    new_n22057_, new_n22058_, new_n22059_, new_n22060_, new_n22061_,
    new_n22062_, new_n22063_, new_n22064_, new_n22065_, new_n22066_,
    new_n22067_, new_n22068_, new_n22069_, new_n22070_, new_n22071_,
    new_n22072_, new_n22073_, new_n22074_, new_n22075_, new_n22076_,
    new_n22077_, new_n22078_, new_n22079_, new_n22080_, new_n22081_,
    new_n22082_, new_n22083_, new_n22084_, new_n22085_, new_n22086_,
    new_n22087_, new_n22088_, new_n22089_, new_n22090_, new_n22091_,
    new_n22092_, new_n22093_, new_n22094_, new_n22095_, new_n22096_,
    new_n22097_, new_n22098_, new_n22099_, new_n22100_, new_n22101_,
    new_n22102_, new_n22103_, new_n22104_, new_n22105_, new_n22106_,
    new_n22107_, new_n22108_, new_n22109_, new_n22110_, new_n22111_,
    new_n22112_, new_n22113_, new_n22114_, new_n22115_, new_n22116_,
    new_n22117_, new_n22118_, new_n22119_, new_n22120_, new_n22121_,
    new_n22122_, new_n22123_, new_n22124_, new_n22125_, new_n22126_,
    new_n22127_, new_n22128_, new_n22129_, new_n22130_, new_n22131_,
    new_n22132_, new_n22133_, new_n22134_, new_n22135_, new_n22136_,
    new_n22137_, new_n22139_, new_n22140_, new_n22141_, new_n22142_,
    new_n22143_, new_n22144_, new_n22145_, new_n22146_, new_n22147_,
    new_n22148_, new_n22149_, new_n22150_, new_n22151_, new_n22152_,
    new_n22153_, new_n22154_, new_n22155_, new_n22156_, new_n22157_,
    new_n22158_, new_n22159_, new_n22160_, new_n22161_, new_n22162_,
    new_n22163_, new_n22164_, new_n22165_, new_n22166_, new_n22167_,
    new_n22168_, new_n22169_, new_n22170_, new_n22171_, new_n22172_,
    new_n22173_, new_n22174_, new_n22175_, new_n22176_, new_n22177_,
    new_n22178_, new_n22179_, new_n22180_, new_n22181_, new_n22182_,
    new_n22183_, new_n22184_, new_n22185_, new_n22186_, new_n22187_,
    new_n22188_, new_n22189_, new_n22190_, new_n22191_, new_n22192_,
    new_n22193_, new_n22194_, new_n22195_, new_n22196_, new_n22197_,
    new_n22198_, new_n22199_, new_n22200_, new_n22201_, new_n22202_,
    new_n22203_, new_n22204_, new_n22205_, new_n22206_, new_n22207_,
    new_n22208_, new_n22209_, new_n22210_, new_n22211_, new_n22212_,
    new_n22213_, new_n22214_, new_n22215_, new_n22216_, new_n22217_,
    new_n22218_, new_n22219_, new_n22220_, new_n22221_, new_n22222_,
    new_n22223_, new_n22224_, new_n22225_, new_n22226_, new_n22227_,
    new_n22228_, new_n22229_, new_n22230_, new_n22231_, new_n22232_,
    new_n22233_, new_n22234_, new_n22235_, new_n22236_, new_n22237_,
    new_n22238_, new_n22239_, new_n22240_, new_n22241_, new_n22242_,
    new_n22243_, new_n22244_, new_n22245_, new_n22246_, new_n22247_,
    new_n22248_, new_n22249_, new_n22250_, new_n22251_, new_n22252_,
    new_n22253_, new_n22254_, new_n22255_, new_n22256_, new_n22257_,
    new_n22258_, new_n22259_, new_n22260_, new_n22261_, new_n22262_,
    new_n22263_, new_n22264_, new_n22265_, new_n22266_, new_n22267_,
    new_n22268_, new_n22269_, new_n22270_, new_n22271_, new_n22272_,
    new_n22273_, new_n22274_, new_n22275_, new_n22276_, new_n22277_,
    new_n22278_, new_n22279_, new_n22280_, new_n22281_, new_n22282_,
    new_n22283_, new_n22284_, new_n22285_, new_n22286_, new_n22287_,
    new_n22288_, new_n22289_, new_n22290_, new_n22291_, new_n22292_,
    new_n22293_, new_n22294_, new_n22295_, new_n22297_, new_n22298_,
    new_n22299_, new_n22300_, new_n22301_, new_n22302_, new_n22303_,
    new_n22304_, new_n22305_, new_n22306_, new_n22307_, new_n22308_,
    new_n22309_, new_n22310_, new_n22311_, new_n22312_, new_n22313_,
    new_n22314_, new_n22315_, new_n22316_, new_n22317_, new_n22318_,
    new_n22319_, new_n22320_, new_n22321_, new_n22322_, new_n22323_,
    new_n22324_, new_n22325_, new_n22326_, new_n22327_, new_n22328_,
    new_n22329_, new_n22330_, new_n22331_, new_n22332_, new_n22333_,
    new_n22334_, new_n22335_, new_n22336_, new_n22337_, new_n22338_,
    new_n22339_, new_n22340_, new_n22341_, new_n22342_, new_n22343_,
    new_n22344_, new_n22345_, new_n22346_, new_n22347_, new_n22348_,
    new_n22349_, new_n22350_, new_n22351_, new_n22352_, new_n22353_,
    new_n22354_, new_n22355_, new_n22356_, new_n22357_, new_n22358_,
    new_n22359_, new_n22360_, new_n22361_, new_n22362_, new_n22363_,
    new_n22364_, new_n22365_, new_n22366_, new_n22367_, new_n22368_,
    new_n22369_, new_n22370_, new_n22371_, new_n22372_, new_n22373_,
    new_n22374_, new_n22375_, new_n22376_, new_n22377_, new_n22378_,
    new_n22379_, new_n22380_, new_n22381_, new_n22382_, new_n22383_,
    new_n22384_, new_n22385_, new_n22386_, new_n22387_, new_n22388_,
    new_n22389_, new_n22390_, new_n22391_, new_n22392_, new_n22393_,
    new_n22394_, new_n22395_, new_n22396_, new_n22397_, new_n22398_,
    new_n22399_, new_n22400_, new_n22401_, new_n22402_, new_n22403_,
    new_n22404_, new_n22405_, new_n22406_, new_n22407_, new_n22408_,
    new_n22409_, new_n22410_, new_n22411_, new_n22412_, new_n22413_,
    new_n22414_, new_n22415_, new_n22416_, new_n22417_, new_n22418_,
    new_n22419_, new_n22420_, new_n22421_, new_n22422_, new_n22423_,
    new_n22424_, new_n22425_, new_n22426_, new_n22427_, new_n22428_,
    new_n22429_, new_n22430_, new_n22431_, new_n22432_, new_n22433_,
    new_n22434_, new_n22435_, new_n22436_, new_n22437_, new_n22438_,
    new_n22439_, new_n22440_, new_n22441_, new_n22442_, new_n22443_,
    new_n22444_, new_n22445_, new_n22446_, new_n22447_, new_n22448_,
    new_n22449_, new_n22450_, new_n22451_, new_n22452_, new_n22453_,
    new_n22454_, new_n22455_, new_n22457_, new_n22458_, new_n22459_,
    new_n22460_, new_n22461_, new_n22462_, new_n22463_, new_n22464_,
    new_n22465_, new_n22466_, new_n22467_, new_n22468_, new_n22469_,
    new_n22470_, new_n22471_, new_n22472_, new_n22473_, new_n22474_,
    new_n22475_, new_n22476_, new_n22477_, new_n22478_, new_n22479_,
    new_n22480_, new_n22481_, new_n22482_, new_n22483_, new_n22484_,
    new_n22485_, new_n22486_, new_n22487_, new_n22488_, new_n22489_,
    new_n22490_, new_n22491_, new_n22492_, new_n22493_, new_n22494_,
    new_n22495_, new_n22496_, new_n22497_, new_n22498_, new_n22499_,
    new_n22500_, new_n22501_, new_n22502_, new_n22503_, new_n22504_,
    new_n22505_, new_n22506_, new_n22507_, new_n22508_, new_n22509_,
    new_n22510_, new_n22511_, new_n22512_, new_n22513_, new_n22514_,
    new_n22515_, new_n22516_, new_n22517_, new_n22518_, new_n22519_,
    new_n22520_, new_n22521_, new_n22522_, new_n22523_, new_n22524_,
    new_n22525_, new_n22526_, new_n22527_, new_n22528_, new_n22529_,
    new_n22530_, new_n22531_, new_n22532_, new_n22533_, new_n22534_,
    new_n22535_, new_n22536_, new_n22537_, new_n22538_, new_n22539_,
    new_n22540_, new_n22541_, new_n22542_, new_n22543_, new_n22544_,
    new_n22545_, new_n22546_, new_n22547_, new_n22548_, new_n22549_,
    new_n22550_, new_n22551_, new_n22552_, new_n22553_, new_n22554_,
    new_n22555_, new_n22556_, new_n22557_, new_n22558_, new_n22559_,
    new_n22560_, new_n22561_, new_n22562_, new_n22563_, new_n22564_,
    new_n22565_, new_n22566_, new_n22567_, new_n22568_, new_n22569_,
    new_n22570_, new_n22571_, new_n22572_, new_n22573_, new_n22574_,
    new_n22575_, new_n22576_, new_n22578_, new_n22579_, new_n22580_,
    new_n22581_, new_n22582_, new_n22584_, new_n22585_, new_n22586_,
    new_n22587_, new_n22589_, new_n22590_, new_n22591_, new_n22592_,
    new_n22593_, new_n22594_, new_n22595_, new_n22596_, new_n22597_,
    new_n22598_, new_n22599_, new_n22600_, new_n22601_, new_n22602_,
    new_n22603_, new_n22604_, new_n22605_, new_n22606_, new_n22607_,
    new_n22608_, new_n22609_, new_n22610_, new_n22611_, new_n22612_,
    new_n22613_, new_n22614_, new_n22615_, new_n22616_, new_n22617_,
    new_n22618_, new_n22619_, new_n22620_, new_n22621_, new_n22622_,
    new_n22623_, new_n22624_, new_n22625_, new_n22626_, new_n22627_,
    new_n22628_, new_n22629_, new_n22630_, new_n22631_, new_n22632_,
    new_n22633_, new_n22634_, new_n22635_, new_n22636_, new_n22637_,
    new_n22638_, new_n22639_, new_n22640_, new_n22641_, new_n22642_,
    new_n22643_, new_n22644_, new_n22645_, new_n22646_, new_n22647_,
    new_n22648_, new_n22650_, new_n22651_, new_n22652_, new_n22654_,
    new_n22655_, new_n22656_, new_n22657_, new_n22658_, new_n22660_,
    new_n22661_, new_n22662_, new_n22663_, new_n22664_, new_n22665_,
    new_n22666_, new_n22667_, new_n22668_, new_n22669_, new_n22670_,
    new_n22671_, new_n22672_, new_n22673_, new_n22674_, new_n22675_,
    new_n22676_, new_n22677_, new_n22678_, new_n22679_, new_n22680_,
    new_n22681_, new_n22682_, new_n22683_, new_n22684_, new_n22685_,
    new_n22686_, new_n22687_, new_n22688_, new_n22689_, new_n22690_,
    new_n22691_, new_n22692_, new_n22693_, new_n22694_, new_n22695_,
    new_n22696_, new_n22697_, new_n22698_, new_n22699_, new_n22700_,
    new_n22701_, new_n22702_, new_n22703_, new_n22704_, new_n22705_,
    new_n22706_, new_n22707_, new_n22708_, new_n22709_, new_n22710_,
    new_n22711_, new_n22712_, new_n22713_, new_n22714_, new_n22715_,
    new_n22716_, new_n22717_, new_n22718_, new_n22719_, new_n22720_,
    new_n22721_, new_n22722_, new_n22723_, new_n22724_, new_n22725_,
    new_n22726_, new_n22727_, new_n22728_, new_n22729_, new_n22730_,
    new_n22731_, new_n22732_, new_n22733_, new_n22734_, new_n22735_,
    new_n22736_, new_n22737_, new_n22738_, new_n22739_, new_n22740_,
    new_n22741_, new_n22742_, new_n22743_, new_n22744_, new_n22745_,
    new_n22746_, new_n22747_, new_n22748_, new_n22749_, new_n22750_,
    new_n22751_, new_n22752_, new_n22753_, new_n22754_, new_n22755_,
    new_n22756_, new_n22757_, new_n22758_, new_n22759_, new_n22760_,
    new_n22761_, new_n22762_, new_n22763_, new_n22764_, new_n22765_,
    new_n22766_, new_n22767_, new_n22768_, new_n22769_, new_n22770_,
    new_n22771_, new_n22772_, new_n22773_, new_n22774_, new_n22775_,
    new_n22776_, new_n22777_, new_n22778_, new_n22779_, new_n22780_,
    new_n22781_, new_n22782_, new_n22783_, new_n22784_, new_n22785_,
    new_n22786_, new_n22787_, new_n22788_, new_n22789_, new_n22790_,
    new_n22791_, new_n22792_, new_n22793_, new_n22794_, new_n22795_,
    new_n22796_, new_n22797_, new_n22798_, new_n22799_, new_n22800_,
    new_n22801_, new_n22802_, new_n22803_, new_n22804_, new_n22805_,
    new_n22806_, new_n22807_, new_n22808_, new_n22809_, new_n22810_,
    new_n22811_, new_n22812_, new_n22813_, new_n22814_, new_n22815_,
    new_n22816_, new_n22817_, new_n22818_, new_n22819_, new_n22820_,
    new_n22821_, new_n22822_, new_n22823_, new_n22824_, new_n22825_,
    new_n22826_, new_n22827_, new_n22828_, new_n22829_, new_n22830_,
    new_n22831_, new_n22832_, new_n22833_, new_n22834_, new_n22835_,
    new_n22836_, new_n22837_, new_n22838_, new_n22839_, new_n22840_,
    new_n22841_, new_n22842_, new_n22843_, new_n22844_, new_n22845_,
    new_n22846_, new_n22847_, new_n22848_, new_n22849_, new_n22850_,
    new_n22851_, new_n22852_, new_n22853_, new_n22854_, new_n22855_,
    new_n22856_, new_n22857_, new_n22858_, new_n22859_, new_n22860_,
    new_n22861_, new_n22862_, new_n22863_, new_n22864_, new_n22865_,
    new_n22866_, new_n22867_, new_n22868_, new_n22869_, new_n22870_,
    new_n22871_, new_n22872_, new_n22873_, new_n22874_, new_n22875_,
    new_n22876_, new_n22877_, new_n22878_, new_n22879_, new_n22880_,
    new_n22881_, new_n22882_, new_n22883_, new_n22884_, new_n22885_,
    new_n22886_, new_n22887_, new_n22888_, new_n22889_, new_n22890_,
    new_n22891_, new_n22892_, new_n22893_, new_n22894_, new_n22895_,
    new_n22896_, new_n22897_, new_n22898_, new_n22899_, new_n22900_,
    new_n22901_, new_n22902_, new_n22903_, new_n22904_, new_n22905_,
    new_n22906_, new_n22907_, new_n22908_, new_n22909_, new_n22910_,
    new_n22911_, new_n22912_, new_n22913_, new_n22914_, new_n22915_,
    new_n22916_, new_n22917_, new_n22918_, new_n22919_, new_n22920_,
    new_n22921_, new_n22922_, new_n22923_, new_n22924_, new_n22925_,
    new_n22926_, new_n22927_, new_n22928_, new_n22929_, new_n22930_,
    new_n22931_, new_n22932_, new_n22933_, new_n22934_, new_n22935_,
    new_n22936_, new_n22937_, new_n22938_, new_n22939_, new_n22940_,
    new_n22941_, new_n22942_, new_n22943_, new_n22944_, new_n22945_,
    new_n22946_, new_n22947_, new_n22948_, new_n22949_, new_n22950_,
    new_n22951_, new_n22952_, new_n22953_, new_n22954_, new_n22955_,
    new_n22956_, new_n22957_, new_n22959_, new_n22960_, new_n22961_,
    new_n22962_, new_n22963_, new_n22964_, new_n22965_, new_n22966_,
    new_n22967_, new_n22968_, new_n22969_, new_n22970_, new_n22971_,
    new_n22972_, new_n22973_, new_n22974_, new_n22975_, new_n22976_,
    new_n22977_, new_n22978_, new_n22979_, new_n22980_, new_n22981_,
    new_n22982_, new_n22983_, new_n22984_, new_n22985_, new_n22986_,
    new_n22987_, new_n22988_, new_n22989_, new_n22990_, new_n22991_,
    new_n22992_, new_n22993_, new_n22994_, new_n22995_, new_n22996_,
    new_n22997_, new_n22998_, new_n22999_, new_n23000_, new_n23002_,
    new_n23003_, new_n23004_, new_n23005_, new_n23006_, new_n23007_,
    new_n23008_, new_n23009_, new_n23010_, new_n23011_, new_n23012_,
    new_n23013_, new_n23014_, new_n23015_, new_n23016_, new_n23017_,
    new_n23018_, new_n23019_, new_n23020_, new_n23021_, new_n23022_,
    new_n23023_, new_n23024_, new_n23025_, new_n23026_, new_n23027_,
    new_n23028_, new_n23029_, new_n23030_, new_n23031_, new_n23032_,
    new_n23033_, new_n23034_, new_n23035_, new_n23036_, new_n23037_,
    new_n23038_, new_n23039_, new_n23040_, new_n23041_, new_n23042_,
    new_n23043_, new_n23044_, new_n23045_, new_n23046_, new_n23047_,
    new_n23048_, new_n23049_, new_n23050_, new_n23051_, new_n23052_,
    new_n23053_, new_n23054_, new_n23055_, new_n23056_, new_n23057_,
    new_n23058_, new_n23059_, new_n23060_, new_n23061_, new_n23062_,
    new_n23063_, new_n23064_, new_n23065_, new_n23066_, new_n23067_,
    new_n23068_, new_n23069_, new_n23070_, new_n23071_, new_n23072_,
    new_n23073_, new_n23074_, new_n23075_, new_n23076_, new_n23077_,
    new_n23078_, new_n23079_, new_n23080_, new_n23081_, new_n23082_,
    new_n23083_, new_n23084_, new_n23085_, new_n23086_, new_n23087_,
    new_n23088_, new_n23089_, new_n23090_, new_n23091_, new_n23092_,
    new_n23093_, new_n23094_, new_n23095_, new_n23096_, new_n23097_,
    new_n23099_, new_n23100_, new_n23101_, new_n23102_, new_n23103_,
    new_n23104_, new_n23105_, new_n23106_, new_n23107_, new_n23108_,
    new_n23109_, new_n23110_, new_n23111_, new_n23112_, new_n23113_,
    new_n23114_, new_n23115_, new_n23116_, new_n23117_, new_n23118_,
    new_n23119_, new_n23120_, new_n23121_, new_n23122_, new_n23123_,
    new_n23124_, new_n23125_, new_n23126_, new_n23127_, new_n23128_,
    new_n23129_, new_n23130_, new_n23131_, new_n23132_, new_n23133_,
    new_n23134_, new_n23135_, new_n23136_, new_n23137_, new_n23138_,
    new_n23139_, new_n23140_, new_n23141_, new_n23142_, new_n23143_,
    new_n23144_, new_n23145_, new_n23146_, new_n23147_, new_n23148_,
    new_n23149_, new_n23150_, new_n23151_, new_n23152_, new_n23153_,
    new_n23154_, new_n23155_, new_n23156_, new_n23157_, new_n23158_,
    new_n23159_, new_n23160_, new_n23161_, new_n23162_, new_n23163_,
    new_n23164_, new_n23165_, new_n23166_, new_n23167_, new_n23168_,
    new_n23169_, new_n23170_, new_n23171_, new_n23173_, new_n23174_,
    new_n23175_, new_n23176_, new_n23177_, new_n23178_, new_n23179_,
    new_n23180_, new_n23181_, new_n23182_, new_n23183_, new_n23184_,
    new_n23185_, new_n23186_, new_n23187_, new_n23188_, new_n23189_,
    new_n23191_, new_n23192_, new_n23193_, new_n23194_, new_n23195_,
    new_n23196_, new_n23197_, new_n23198_, new_n23199_, new_n23200_,
    new_n23202_, new_n23203_, new_n23204_, new_n23205_, new_n23206_,
    new_n23207_, new_n23208_, new_n23209_, new_n23210_, new_n23211_,
    new_n23212_, new_n23214_, new_n23215_, new_n23216_, new_n23217_,
    new_n23218_, new_n23219_, new_n23220_, new_n23221_, new_n23222_,
    new_n23223_, new_n23225_, new_n23226_, new_n23227_, new_n23228_,
    new_n23229_, new_n23230_, new_n23231_, new_n23232_, new_n23233_,
    new_n23234_, new_n23235_, new_n23236_, new_n23237_, new_n23238_,
    new_n23239_, new_n23240_, new_n23241_, new_n23242_, new_n23243_,
    new_n23244_, new_n23245_, new_n23246_, new_n23247_, new_n23248_,
    new_n23249_, new_n23250_, new_n23251_, new_n23252_, new_n23253_,
    new_n23254_, new_n23255_, new_n23256_, new_n23257_, new_n23258_,
    new_n23259_, new_n23260_, new_n23261_, new_n23262_, new_n23263_,
    new_n23264_, new_n23265_, new_n23266_, new_n23267_, new_n23268_,
    new_n23269_, new_n23270_, new_n23271_, new_n23272_, new_n23273_,
    new_n23274_, new_n23275_, new_n23276_, new_n23277_, new_n23278_,
    new_n23279_, new_n23280_, new_n23281_, new_n23282_, new_n23283_,
    new_n23284_, new_n23285_, new_n23286_, new_n23287_, new_n23288_,
    new_n23289_, new_n23290_, new_n23291_, new_n23292_, new_n23293_,
    new_n23294_, new_n23295_, new_n23297_, new_n23298_, new_n23299_,
    new_n23300_, new_n23301_, new_n23302_, new_n23303_, new_n23304_,
    new_n23305_, new_n23306_, new_n23307_, new_n23308_, new_n23309_,
    new_n23310_, new_n23311_, new_n23312_, new_n23313_, new_n23314_,
    new_n23315_, new_n23316_, new_n23317_, new_n23318_, new_n23319_,
    new_n23320_, new_n23321_, new_n23322_, new_n23323_, new_n23324_,
    new_n23325_, new_n23326_, new_n23327_, new_n23328_, new_n23329_,
    new_n23330_, new_n23331_, new_n23332_, new_n23333_, new_n23334_,
    new_n23335_, new_n23336_, new_n23337_, new_n23338_, new_n23339_,
    new_n23340_, new_n23341_, new_n23342_, new_n23343_, new_n23344_,
    new_n23345_, new_n23346_, new_n23347_, new_n23348_, new_n23349_,
    new_n23350_, new_n23351_, new_n23352_, new_n23353_, new_n23354_,
    new_n23355_, new_n23356_, new_n23357_, new_n23358_, new_n23359_,
    new_n23360_, new_n23361_, new_n23362_, new_n23363_, new_n23364_,
    new_n23366_, new_n23367_, new_n23368_, new_n23369_, new_n23370_,
    new_n23371_, new_n23372_, new_n23373_, new_n23374_, new_n23375_,
    new_n23376_, new_n23377_, new_n23378_, new_n23379_, new_n23381_,
    new_n23382_, new_n23383_, new_n23385_, new_n23386_, new_n23387_,
    new_n23388_, new_n23389_, new_n23390_, new_n23391_, new_n23392_,
    new_n23393_, new_n23394_, new_n23396_, new_n23397_, new_n23398_,
    new_n23400_, new_n23401_, new_n23402_, new_n23403_, new_n23404_,
    new_n23405_, new_n23406_, new_n23407_, new_n23408_, new_n23409_,
    new_n23410_, new_n23411_, new_n23412_, new_n23413_, new_n23414_,
    new_n23415_, new_n23416_, new_n23417_, new_n23418_, new_n23419_,
    new_n23420_, new_n23421_, new_n23422_, new_n23423_, new_n23424_,
    new_n23425_, new_n23426_, new_n23427_, new_n23428_, new_n23429_,
    new_n23430_, new_n23431_, new_n23432_, new_n23433_, new_n23434_,
    new_n23435_, new_n23436_, new_n23437_, new_n23438_, new_n23439_,
    new_n23440_, new_n23441_, new_n23442_, new_n23443_, new_n23444_,
    new_n23445_, new_n23446_, new_n23447_, new_n23448_, new_n23449_,
    new_n23450_, new_n23451_, new_n23452_, new_n23453_, new_n23454_,
    new_n23455_, new_n23456_, new_n23457_, new_n23458_, new_n23459_,
    new_n23460_, new_n23461_, new_n23462_, new_n23463_, new_n23464_,
    new_n23465_, new_n23466_, new_n23468_, new_n23469_, new_n23470_,
    new_n23471_, new_n23472_, new_n23473_, new_n23474_, new_n23475_,
    new_n23476_, new_n23477_, new_n23478_, new_n23479_, new_n23480_,
    new_n23481_, new_n23482_, new_n23483_, new_n23484_, new_n23485_,
    new_n23486_, new_n23487_, new_n23488_, new_n23489_, new_n23490_,
    new_n23491_, new_n23492_, new_n23493_, new_n23494_, new_n23495_,
    new_n23496_, new_n23497_, new_n23498_, new_n23499_, new_n23500_,
    new_n23501_, new_n23502_, new_n23503_, new_n23504_, new_n23505_,
    new_n23506_, new_n23507_, new_n23508_, new_n23509_, new_n23510_,
    new_n23511_, new_n23512_, new_n23513_, new_n23514_, new_n23515_,
    new_n23516_, new_n23517_, new_n23518_, new_n23519_, new_n23520_,
    new_n23521_, new_n23522_, new_n23523_, new_n23524_, new_n23525_,
    new_n23526_, new_n23527_, new_n23528_, new_n23529_, new_n23530_,
    new_n23531_, new_n23532_, new_n23533_, new_n23534_, new_n23535_,
    new_n23536_, new_n23537_, new_n23538_, new_n23539_, new_n23540_,
    new_n23541_, new_n23542_, new_n23543_, new_n23544_, new_n23545_,
    new_n23546_, new_n23547_, new_n23548_, new_n23549_, new_n23550_,
    new_n23551_, new_n23552_, new_n23553_, new_n23554_, new_n23555_,
    new_n23556_, new_n23557_, new_n23558_, new_n23559_, new_n23560_,
    new_n23561_, new_n23562_, new_n23563_, new_n23564_, new_n23565_,
    new_n23566_, new_n23567_, new_n23568_, new_n23569_, new_n23570_,
    new_n23571_, new_n23572_, new_n23573_, new_n23574_, new_n23575_,
    new_n23576_, new_n23577_, new_n23578_, new_n23579_, new_n23580_,
    new_n23581_, new_n23582_, new_n23583_, new_n23584_, new_n23585_,
    new_n23586_, new_n23587_, new_n23588_, new_n23589_, new_n23590_,
    new_n23591_, new_n23592_, new_n23593_, new_n23594_, new_n23595_,
    new_n23596_, new_n23597_, new_n23598_, new_n23599_, new_n23600_,
    new_n23601_, new_n23602_, new_n23603_, new_n23604_, new_n23605_,
    new_n23606_, new_n23607_, new_n23608_, new_n23609_, new_n23610_,
    new_n23611_, new_n23612_, new_n23613_, new_n23614_, new_n23615_,
    new_n23616_, new_n23617_, new_n23618_, new_n23619_, new_n23620_,
    new_n23621_, new_n23622_, new_n23623_, new_n23624_, new_n23625_,
    new_n23626_, new_n23627_, new_n23628_, new_n23629_, new_n23630_,
    new_n23631_, new_n23632_, new_n23633_, new_n23634_, new_n23635_,
    new_n23636_, new_n23637_, new_n23638_, new_n23639_, new_n23640_,
    new_n23641_, new_n23642_, new_n23643_, new_n23644_, new_n23645_,
    new_n23646_, new_n23647_, new_n23648_, new_n23649_, new_n23650_,
    new_n23651_, new_n23652_, new_n23653_, new_n23654_, new_n23655_,
    new_n23656_, new_n23657_, new_n23658_, new_n23659_, new_n23660_,
    new_n23661_, new_n23662_, new_n23663_, new_n23664_, new_n23665_,
    new_n23666_, new_n23667_, new_n23668_, new_n23669_, new_n23670_,
    new_n23671_, new_n23672_, new_n23673_, new_n23674_, new_n23675_,
    new_n23676_, new_n23677_, new_n23678_, new_n23679_, new_n23680_,
    new_n23681_, new_n23682_, new_n23683_, new_n23684_, new_n23685_,
    new_n23686_, new_n23687_, new_n23688_, new_n23689_, new_n23690_,
    new_n23691_, new_n23692_, new_n23693_, new_n23694_, new_n23695_,
    new_n23696_, new_n23697_, new_n23698_, new_n23699_, new_n23700_,
    new_n23701_, new_n23702_, new_n23703_, new_n23704_, new_n23705_,
    new_n23706_, new_n23707_, new_n23708_, new_n23709_, new_n23710_,
    new_n23711_, new_n23712_, new_n23713_, new_n23714_, new_n23715_,
    new_n23716_, new_n23717_, new_n23718_, new_n23719_, new_n23720_,
    new_n23721_, new_n23722_, new_n23723_, new_n23724_, new_n23725_,
    new_n23726_, new_n23727_, new_n23728_, new_n23729_, new_n23730_,
    new_n23731_, new_n23732_, new_n23733_, new_n23734_, new_n23735_,
    new_n23736_, new_n23737_, new_n23738_, new_n23739_, new_n23740_,
    new_n23741_, new_n23742_, new_n23743_, new_n23744_, new_n23745_,
    new_n23746_, new_n23747_, new_n23748_, new_n23749_, new_n23750_,
    new_n23751_, new_n23752_, new_n23753_, new_n23754_, new_n23755_,
    new_n23756_, new_n23757_, new_n23758_, new_n23759_, new_n23760_,
    new_n23761_, new_n23762_, new_n23763_, new_n23764_, new_n23765_,
    new_n23766_, new_n23767_, new_n23768_, new_n23769_, new_n23770_,
    new_n23771_, new_n23772_, new_n23773_, new_n23774_, new_n23775_,
    new_n23776_, new_n23777_, new_n23778_, new_n23779_, new_n23780_,
    new_n23781_, new_n23782_, new_n23783_, new_n23784_, new_n23785_,
    new_n23786_, new_n23787_, new_n23788_, new_n23789_, new_n23790_,
    new_n23791_, new_n23792_, new_n23793_, new_n23794_, new_n23795_,
    new_n23796_, new_n23797_, new_n23798_, new_n23799_, new_n23800_,
    new_n23801_, new_n23802_, new_n23803_, new_n23804_, new_n23805_,
    new_n23806_, new_n23807_, new_n23808_, new_n23809_, new_n23810_,
    new_n23811_, new_n23812_, new_n23813_, new_n23814_, new_n23815_,
    new_n23816_, new_n23817_, new_n23818_, new_n23819_, new_n23820_,
    new_n23821_, new_n23822_, new_n23823_, new_n23824_, new_n23825_,
    new_n23826_, new_n23827_, new_n23828_, new_n23829_, new_n23830_,
    new_n23831_, new_n23832_, new_n23833_, new_n23834_, new_n23835_,
    new_n23836_, new_n23837_, new_n23838_, new_n23839_, new_n23840_,
    new_n23841_, new_n23842_, new_n23843_, new_n23844_, new_n23845_,
    new_n23846_, new_n23847_, new_n23848_, new_n23849_, new_n23850_,
    new_n23851_, new_n23852_, new_n23853_, new_n23854_, new_n23855_,
    new_n23856_, new_n23857_, new_n23858_, new_n23859_, new_n23860_,
    new_n23861_, new_n23862_, new_n23863_, new_n23864_, new_n23865_,
    new_n23866_, new_n23867_, new_n23868_, new_n23869_, new_n23871_,
    new_n23872_, new_n23873_, new_n23874_, new_n23875_, new_n23876_,
    new_n23877_, new_n23878_, new_n23879_, new_n23880_, new_n23881_,
    new_n23882_, new_n23883_, new_n23884_, new_n23885_, new_n23886_,
    new_n23887_, new_n23888_, new_n23889_, new_n23890_, new_n23891_,
    new_n23892_, new_n23893_, new_n23894_, new_n23895_, new_n23896_,
    new_n23897_, new_n23898_, new_n23899_, new_n23900_, new_n23901_,
    new_n23902_, new_n23903_, new_n23904_, new_n23905_, new_n23906_,
    new_n23907_, new_n23908_, new_n23909_, new_n23910_, new_n23911_,
    new_n23912_, new_n23913_, new_n23914_, new_n23915_, new_n23916_,
    new_n23917_, new_n23918_, new_n23919_, new_n23920_, new_n23921_,
    new_n23922_, new_n23923_, new_n23924_, new_n23925_, new_n23926_,
    new_n23927_, new_n23928_, new_n23929_, new_n23930_, new_n23931_,
    new_n23932_, new_n23933_, new_n23934_, new_n23935_, new_n23936_,
    new_n23937_, new_n23938_, new_n23939_, new_n23940_, new_n23941_,
    new_n23942_, new_n23943_, new_n23944_, new_n23945_, new_n23946_,
    new_n23947_, new_n23948_, new_n23949_, new_n23950_, new_n23951_,
    new_n23952_, new_n23953_, new_n23954_, new_n23955_, new_n23956_,
    new_n23957_, new_n23958_, new_n23959_, new_n23960_, new_n23961_,
    new_n23962_, new_n23963_, new_n23964_, new_n23965_, new_n23966_,
    new_n23967_, new_n23968_, new_n23969_, new_n23970_, new_n23971_,
    new_n23972_, new_n23973_, new_n23974_, new_n23975_, new_n23976_,
    new_n23977_, new_n23978_, new_n23979_, new_n23980_, new_n23981_,
    new_n23982_, new_n23983_, new_n23984_, new_n23985_, new_n23986_,
    new_n23987_, new_n23988_, new_n23989_, new_n23990_, new_n23991_,
    new_n23992_, new_n23993_, new_n23994_, new_n23995_, new_n23996_,
    new_n23997_, new_n23998_, new_n23999_, new_n24000_, new_n24001_,
    new_n24002_, new_n24003_, new_n24004_, new_n24005_, new_n24006_,
    new_n24007_, new_n24008_, new_n24009_, new_n24010_, new_n24011_,
    new_n24012_, new_n24013_, new_n24014_, new_n24015_, new_n24016_,
    new_n24017_, new_n24018_, new_n24019_, new_n24020_, new_n24021_,
    new_n24022_, new_n24023_, new_n24024_, new_n24025_, new_n24026_,
    new_n24027_, new_n24028_, new_n24029_, new_n24030_, new_n24031_,
    new_n24032_, new_n24033_, new_n24034_, new_n24035_, new_n24036_,
    new_n24037_, new_n24038_, new_n24039_, new_n24040_, new_n24041_,
    new_n24042_, new_n24043_, new_n24044_, new_n24045_, new_n24046_,
    new_n24047_, new_n24048_, new_n24049_, new_n24050_, new_n24051_,
    new_n24052_, new_n24053_, new_n24054_, new_n24055_, new_n24056_,
    new_n24057_, new_n24058_, new_n24059_, new_n24060_, new_n24061_,
    new_n24062_, new_n24063_, new_n24064_, new_n24065_, new_n24066_,
    new_n24067_, new_n24068_, new_n24069_, new_n24070_, new_n24071_,
    new_n24072_, new_n24073_, new_n24074_, new_n24075_, new_n24076_,
    new_n24077_, new_n24078_, new_n24079_, new_n24080_, new_n24081_,
    new_n24082_, new_n24083_, new_n24084_, new_n24085_, new_n24086_,
    new_n24087_, new_n24088_, new_n24089_, new_n24090_, new_n24091_,
    new_n24092_, new_n24093_, new_n24094_, new_n24095_, new_n24096_,
    new_n24097_, new_n24098_, new_n24099_, new_n24100_, new_n24101_,
    new_n24102_, new_n24103_, new_n24104_, new_n24105_, new_n24106_,
    new_n24107_, new_n24108_, new_n24109_, new_n24110_, new_n24111_,
    new_n24112_, new_n24113_, new_n24114_, new_n24115_, new_n24116_,
    new_n24117_, new_n24118_, new_n24119_, new_n24120_, new_n24121_,
    new_n24122_, new_n24123_, new_n24124_, new_n24125_, new_n24126_,
    new_n24127_, new_n24128_, new_n24129_, new_n24130_, new_n24131_,
    new_n24132_, new_n24133_, new_n24134_, new_n24135_, new_n24136_,
    new_n24137_, new_n24138_, new_n24139_, new_n24140_, new_n24141_,
    new_n24142_, new_n24143_, new_n24144_, new_n24145_, new_n24146_,
    new_n24147_, new_n24148_, new_n24149_, new_n24150_, new_n24151_,
    new_n24152_, new_n24153_, new_n24154_, new_n24155_, new_n24156_,
    new_n24157_, new_n24158_, new_n24159_, new_n24160_, new_n24161_,
    new_n24162_, new_n24163_, new_n24164_, new_n24165_, new_n24166_,
    new_n24167_, new_n24168_, new_n24169_, new_n24170_, new_n24171_,
    new_n24172_, new_n24173_, new_n24174_, new_n24175_, new_n24176_,
    new_n24177_, new_n24178_, new_n24179_, new_n24180_, new_n24181_,
    new_n24182_, new_n24183_, new_n24184_, new_n24185_, new_n24186_,
    new_n24187_, new_n24188_, new_n24189_, new_n24190_, new_n24191_,
    new_n24192_, new_n24193_, new_n24194_, new_n24195_, new_n24196_,
    new_n24197_, new_n24198_, new_n24199_, new_n24200_, new_n24201_,
    new_n24202_, new_n24203_, new_n24204_, new_n24205_, new_n24206_,
    new_n24207_, new_n24208_, new_n24209_, new_n24210_, new_n24211_,
    new_n24212_, new_n24213_, new_n24214_, new_n24215_, new_n24216_,
    new_n24217_, new_n24218_, new_n24219_, new_n24220_, new_n24221_,
    new_n24222_, new_n24223_, new_n24224_, new_n24225_, new_n24226_,
    new_n24227_, new_n24228_, new_n24229_, new_n24230_, new_n24231_,
    new_n24232_, new_n24233_, new_n24234_, new_n24235_, new_n24236_,
    new_n24237_, new_n24238_, new_n24239_, new_n24241_, new_n24242_,
    new_n24243_, new_n24244_, new_n24245_, new_n24246_, new_n24247_,
    new_n24248_, new_n24249_, new_n24250_, new_n24251_, new_n24252_,
    new_n24253_, new_n24254_, new_n24255_, new_n24256_, new_n24257_,
    new_n24258_, new_n24259_, new_n24260_, new_n24261_, new_n24262_,
    new_n24263_, new_n24264_, new_n24265_, new_n24266_, new_n24267_,
    new_n24268_, new_n24269_, new_n24270_, new_n24271_, new_n24272_,
    new_n24273_, new_n24274_, new_n24275_, new_n24276_, new_n24277_,
    new_n24278_, new_n24279_, new_n24280_, new_n24281_, new_n24282_,
    new_n24283_, new_n24284_, new_n24285_, new_n24286_, new_n24287_,
    new_n24288_, new_n24289_, new_n24290_, new_n24291_, new_n24292_,
    new_n24293_, new_n24294_, new_n24295_, new_n24296_, new_n24297_,
    new_n24298_, new_n24299_, new_n24300_, new_n24301_, new_n24302_,
    new_n24303_, new_n24304_, new_n24305_, new_n24306_, new_n24307_,
    new_n24308_, new_n24309_, new_n24310_, new_n24311_, new_n24312_,
    new_n24313_, new_n24314_, new_n24315_, new_n24316_, new_n24317_,
    new_n24318_, new_n24319_, new_n24320_, new_n24321_, new_n24322_,
    new_n24323_, new_n24324_, new_n24325_, new_n24326_, new_n24327_,
    new_n24328_, new_n24329_, new_n24330_, new_n24331_, new_n24332_,
    new_n24333_, new_n24334_, new_n24335_, new_n24336_, new_n24337_,
    new_n24338_, new_n24339_, new_n24340_, new_n24341_, new_n24342_,
    new_n24343_, new_n24344_, new_n24345_, new_n24346_, new_n24347_,
    new_n24348_, new_n24349_, new_n24350_, new_n24351_, new_n24352_,
    new_n24353_, new_n24354_, new_n24355_, new_n24356_, new_n24357_,
    new_n24358_, new_n24359_, new_n24360_, new_n24361_, new_n24362_,
    new_n24363_, new_n24364_, new_n24365_, new_n24366_, new_n24367_,
    new_n24368_, new_n24369_, new_n24370_, new_n24371_, new_n24372_,
    new_n24373_, new_n24374_, new_n24375_, new_n24376_, new_n24377_,
    new_n24378_, new_n24379_, new_n24380_, new_n24381_, new_n24382_,
    new_n24383_, new_n24384_, new_n24385_, new_n24386_, new_n24387_,
    new_n24388_, new_n24389_, new_n24390_, new_n24391_, new_n24392_,
    new_n24393_, new_n24394_, new_n24395_, new_n24396_, new_n24397_,
    new_n24398_, new_n24399_, new_n24400_, new_n24401_, new_n24402_,
    new_n24403_, new_n24404_, new_n24405_, new_n24406_, new_n24407_,
    new_n24408_, new_n24409_, new_n24410_, new_n24411_, new_n24412_,
    new_n24413_, new_n24414_, new_n24415_, new_n24416_, new_n24417_,
    new_n24418_, new_n24419_, new_n24420_, new_n24421_, new_n24422_,
    new_n24423_, new_n24424_, new_n24425_, new_n24426_, new_n24427_,
    new_n24428_, new_n24429_, new_n24430_, new_n24431_, new_n24432_,
    new_n24433_, new_n24434_, new_n24435_, new_n24436_, new_n24437_,
    new_n24438_, new_n24439_, new_n24440_, new_n24441_, new_n24442_,
    new_n24443_, new_n24444_, new_n24445_, new_n24446_, new_n24447_,
    new_n24448_, new_n24449_, new_n24450_, new_n24451_, new_n24452_,
    new_n24453_, new_n24454_, new_n24455_, new_n24456_, new_n24457_,
    new_n24458_, new_n24459_, new_n24460_, new_n24461_, new_n24462_,
    new_n24463_, new_n24464_, new_n24465_, new_n24466_, new_n24467_,
    new_n24468_, new_n24469_, new_n24470_, new_n24471_, new_n24472_,
    new_n24473_, new_n24474_, new_n24475_, new_n24476_, new_n24477_,
    new_n24478_, new_n24479_, new_n24480_, new_n24481_, new_n24482_,
    new_n24483_, new_n24484_, new_n24485_, new_n24486_, new_n24487_,
    new_n24488_, new_n24489_, new_n24490_, new_n24491_, new_n24492_,
    new_n24493_, new_n24494_, new_n24495_, new_n24496_, new_n24497_,
    new_n24498_, new_n24499_, new_n24500_, new_n24501_, new_n24502_,
    new_n24503_, new_n24504_, new_n24505_, new_n24506_, new_n24507_,
    new_n24508_, new_n24509_, new_n24510_, new_n24511_, new_n24512_,
    new_n24513_, new_n24514_, new_n24515_, new_n24516_, new_n24517_,
    new_n24518_, new_n24519_, new_n24520_, new_n24521_, new_n24522_,
    new_n24523_, new_n24524_, new_n24525_, new_n24526_, new_n24527_,
    new_n24528_, new_n24529_, new_n24530_, new_n24531_, new_n24532_,
    new_n24533_, new_n24534_, new_n24535_, new_n24536_, new_n24537_,
    new_n24538_, new_n24539_, new_n24540_, new_n24541_, new_n24542_,
    new_n24543_, new_n24544_, new_n24545_, new_n24546_, new_n24547_,
    new_n24548_, new_n24549_, new_n24550_, new_n24551_, new_n24552_,
    new_n24553_, new_n24554_, new_n24555_, new_n24556_, new_n24557_,
    new_n24558_, new_n24559_, new_n24560_, new_n24561_, new_n24562_,
    new_n24563_, new_n24564_, new_n24565_, new_n24566_, new_n24567_,
    new_n24568_, new_n24569_, new_n24570_, new_n24571_, new_n24572_,
    new_n24573_, new_n24574_, new_n24575_, new_n24576_, new_n24577_,
    new_n24578_, new_n24579_, new_n24580_, new_n24581_, new_n24582_,
    new_n24583_, new_n24584_, new_n24586_, new_n24587_, new_n24588_,
    new_n24589_, new_n24590_, new_n24591_, new_n24592_, new_n24593_,
    new_n24594_, new_n24595_, new_n24596_, new_n24597_, new_n24598_,
    new_n24599_, new_n24600_, new_n24601_, new_n24602_, new_n24603_,
    new_n24604_, new_n24605_, new_n24606_, new_n24607_, new_n24608_,
    new_n24609_, new_n24610_, new_n24611_, new_n24612_, new_n24613_,
    new_n24614_, new_n24615_, new_n24616_, new_n24617_, new_n24618_,
    new_n24619_, new_n24620_, new_n24621_, new_n24622_, new_n24623_,
    new_n24624_, new_n24625_, new_n24626_, new_n24627_, new_n24628_,
    new_n24629_, new_n24630_, new_n24631_, new_n24632_, new_n24633_,
    new_n24634_, new_n24635_, new_n24636_, new_n24637_, new_n24638_,
    new_n24639_, new_n24640_, new_n24641_, new_n24642_, new_n24643_,
    new_n24644_, new_n24645_, new_n24646_, new_n24647_, new_n24648_,
    new_n24649_, new_n24650_, new_n24651_, new_n24652_, new_n24653_,
    new_n24654_, new_n24655_, new_n24656_, new_n24657_, new_n24658_,
    new_n24659_, new_n24660_, new_n24661_, new_n24663_, new_n24664_,
    new_n24665_, new_n24666_, new_n24667_, new_n24668_, new_n24669_,
    new_n24670_, new_n24671_, new_n24672_, new_n24673_, new_n24674_,
    new_n24675_, new_n24676_, new_n24677_, new_n24678_, new_n24679_,
    new_n24680_, new_n24681_, new_n24682_, new_n24683_, new_n24684_,
    new_n24685_, new_n24686_, new_n24687_, new_n24688_, new_n24689_,
    new_n24690_, new_n24691_, new_n24692_, new_n24694_, new_n24695_,
    new_n24696_, new_n24697_, new_n24698_, new_n24699_, new_n24700_,
    new_n24701_, new_n24702_, new_n24703_, new_n24704_, new_n24705_,
    new_n24706_, new_n24707_, new_n24708_, new_n24709_, new_n24710_,
    new_n24711_, new_n24712_, new_n24713_, new_n24714_, new_n24716_,
    new_n24717_, new_n24718_, new_n24719_, new_n24720_, new_n24721_,
    new_n24723_, new_n24724_, new_n24725_, new_n24726_, new_n24727_,
    new_n24728_, new_n24729_, new_n24730_, new_n24731_, new_n24732_,
    new_n24733_, new_n24734_, new_n24735_, new_n24736_, new_n24737_,
    new_n24738_, new_n24739_, new_n24740_, new_n24741_, new_n24742_,
    new_n24743_, new_n24744_, new_n24745_, new_n24746_, new_n24747_,
    new_n24748_, new_n24749_, new_n24750_, new_n24751_, new_n24752_,
    new_n24753_, new_n24754_, new_n24755_, new_n24756_, new_n24757_,
    new_n24758_, new_n24759_, new_n24760_, new_n24761_, new_n24762_,
    new_n24763_, new_n24764_, new_n24765_, new_n24766_, new_n24767_,
    new_n24768_, new_n24769_, new_n24770_, new_n24771_, new_n24772_,
    new_n24773_, new_n24774_, new_n24775_, new_n24776_, new_n24777_,
    new_n24778_, new_n24780_, new_n24781_, new_n24782_, new_n24783_,
    new_n24784_, new_n24785_, new_n24786_, new_n24787_, new_n24788_,
    new_n24789_, new_n24790_, new_n24791_, new_n24792_, new_n24793_,
    new_n24794_, new_n24795_, new_n24796_, new_n24797_, new_n24798_,
    new_n24800_, new_n24801_, new_n24802_, new_n24803_, new_n24804_,
    new_n24805_, new_n24806_, new_n24807_, new_n24808_, new_n24809_,
    new_n24810_, new_n24811_, new_n24812_, new_n24814_, new_n24815_,
    new_n24816_, new_n24817_, new_n24818_, new_n24819_, new_n24820_,
    new_n24821_, new_n24822_, new_n24823_, new_n24824_, new_n24825_,
    new_n24826_, new_n24827_, new_n24828_, new_n24829_, new_n24830_,
    new_n24831_, new_n24832_, new_n24833_, new_n24834_, new_n24835_,
    new_n24836_, new_n24837_, new_n24838_, new_n24839_, new_n24840_,
    new_n24841_, new_n24842_, new_n24843_, new_n24844_, new_n24845_,
    new_n24846_, new_n24847_, new_n24848_, new_n24849_, new_n24850_,
    new_n24851_, new_n24852_, new_n24853_, new_n24854_, new_n24855_,
    new_n24856_, new_n24857_, new_n24858_, new_n24859_, new_n24860_,
    new_n24861_, new_n24862_, new_n24863_, new_n24864_, new_n24865_,
    new_n24866_, new_n24867_, new_n24868_, new_n24869_, new_n24870_,
    new_n24871_, new_n24872_, new_n24873_, new_n24874_, new_n24875_,
    new_n24876_, new_n24877_, new_n24878_, new_n24879_, new_n24880_,
    new_n24881_, new_n24882_, new_n24883_, new_n24884_, new_n24885_,
    new_n24886_, new_n24887_, new_n24888_, new_n24889_, new_n24890_,
    new_n24891_, new_n24892_, new_n24893_, new_n24894_, new_n24895_,
    new_n24896_, new_n24897_, new_n24898_, new_n24899_, new_n24900_,
    new_n24901_, new_n24902_, new_n24903_, new_n24904_, new_n24905_,
    new_n24906_, new_n24907_, new_n24908_, new_n24909_, new_n24910_,
    new_n24911_, new_n24912_, new_n24913_, new_n24914_, new_n24915_,
    new_n24916_, new_n24917_, new_n24918_, new_n24919_, new_n24920_,
    new_n24921_, new_n24922_, new_n24923_, new_n24924_, new_n24925_,
    new_n24926_, new_n24927_, new_n24928_, new_n24929_, new_n24930_,
    new_n24931_, new_n24932_, new_n24933_, new_n24934_, new_n24935_,
    new_n24936_, new_n24937_, new_n24938_, new_n24939_, new_n24940_,
    new_n24941_, new_n24942_, new_n24943_, new_n24944_, new_n24945_,
    new_n24946_, new_n24947_, new_n24948_, new_n24949_, new_n24950_,
    new_n24951_, new_n24952_, new_n24953_, new_n24954_, new_n24955_,
    new_n24956_, new_n24957_, new_n24958_, new_n24959_, new_n24960_,
    new_n24961_, new_n24962_, new_n24963_, new_n24964_, new_n24965_,
    new_n24966_, new_n24967_, new_n24968_, new_n24969_, new_n24970_,
    new_n24971_, new_n24972_, new_n24973_, new_n24974_, new_n24975_,
    new_n24976_, new_n24977_, new_n24978_, new_n24979_, new_n24980_,
    new_n24981_, new_n24982_, new_n24983_, new_n24984_, new_n24985_,
    new_n24986_, new_n24987_, new_n24988_, new_n24989_, new_n24990_,
    new_n24991_, new_n24992_, new_n24993_, new_n24994_, new_n24995_,
    new_n24996_, new_n24997_, new_n24998_, new_n24999_, new_n25000_,
    new_n25001_, new_n25002_, new_n25003_, new_n25004_, new_n25005_,
    new_n25006_, new_n25007_, new_n25008_, new_n25009_, new_n25010_,
    new_n25011_, new_n25012_, new_n25013_, new_n25014_, new_n25015_,
    new_n25016_, new_n25017_, new_n25018_, new_n25019_, new_n25020_,
    new_n25021_, new_n25022_, new_n25023_, new_n25024_, new_n25025_,
    new_n25026_, new_n25027_, new_n25028_, new_n25029_, new_n25030_,
    new_n25031_, new_n25032_, new_n25033_, new_n25034_, new_n25035_,
    new_n25036_, new_n25037_, new_n25038_, new_n25039_, new_n25040_,
    new_n25041_, new_n25042_, new_n25043_, new_n25044_, new_n25045_,
    new_n25046_, new_n25047_, new_n25048_, new_n25049_, new_n25050_,
    new_n25051_, new_n25052_, new_n25053_, new_n25054_, new_n25055_,
    new_n25056_, new_n25057_, new_n25058_, new_n25059_, new_n25060_,
    new_n25061_, new_n25062_, new_n25063_, new_n25064_, new_n25065_,
    new_n25066_, new_n25067_, new_n25068_, new_n25069_, new_n25070_,
    new_n25071_, new_n25072_, new_n25073_, new_n25074_, new_n25075_,
    new_n25076_, new_n25077_, new_n25078_, new_n25079_, new_n25080_,
    new_n25081_, new_n25082_, new_n25083_, new_n25084_, new_n25085_,
    new_n25086_, new_n25087_, new_n25088_, new_n25089_, new_n25090_,
    new_n25091_, new_n25092_, new_n25093_, new_n25094_, new_n25095_,
    new_n25096_, new_n25097_, new_n25098_, new_n25099_, new_n25100_,
    new_n25101_, new_n25102_, new_n25103_, new_n25104_, new_n25105_,
    new_n25106_, new_n25107_, new_n25109_, new_n25110_, new_n25111_,
    new_n25112_, new_n25113_, new_n25114_, new_n25115_, new_n25116_,
    new_n25117_, new_n25118_, new_n25119_, new_n25120_, new_n25121_,
    new_n25122_, new_n25123_, new_n25124_, new_n25125_, new_n25126_,
    new_n25127_, new_n25128_, new_n25129_, new_n25130_, new_n25131_,
    new_n25132_, new_n25133_, new_n25134_, new_n25135_, new_n25136_,
    new_n25137_, new_n25138_, new_n25139_, new_n25140_, new_n25141_,
    new_n25142_, new_n25143_, new_n25144_, new_n25145_, new_n25146_,
    new_n25147_, new_n25148_, new_n25149_, new_n25150_, new_n25151_,
    new_n25152_, new_n25153_, new_n25154_, new_n25155_, new_n25156_,
    new_n25157_, new_n25158_, new_n25159_, new_n25160_, new_n25161_,
    new_n25162_, new_n25163_, new_n25164_, new_n25165_, new_n25166_,
    new_n25167_, new_n25168_, new_n25169_, new_n25170_, new_n25171_,
    new_n25172_, new_n25173_, new_n25174_, new_n25175_, new_n25176_,
    new_n25177_, new_n25178_, new_n25179_, new_n25180_, new_n25181_,
    new_n25182_, new_n25183_, new_n25184_, new_n25185_, new_n25186_,
    new_n25187_, new_n25188_, new_n25189_, new_n25190_, new_n25191_,
    new_n25192_, new_n25193_, new_n25194_, new_n25195_, new_n25196_,
    new_n25197_, new_n25198_, new_n25199_, new_n25200_, new_n25201_,
    new_n25202_, new_n25203_, new_n25204_, new_n25205_, new_n25206_,
    new_n25207_, new_n25208_, new_n25209_, new_n25210_, new_n25211_,
    new_n25212_, new_n25213_, new_n25214_, new_n25215_, new_n25216_,
    new_n25217_, new_n25218_, new_n25219_, new_n25220_, new_n25221_,
    new_n25222_, new_n25223_, new_n25224_, new_n25225_, new_n25226_,
    new_n25227_, new_n25228_, new_n25229_, new_n25230_, new_n25231_,
    new_n25232_, new_n25233_, new_n25234_, new_n25235_, new_n25236_,
    new_n25237_, new_n25238_, new_n25239_, new_n25240_, new_n25241_,
    new_n25242_, new_n25243_, new_n25244_, new_n25245_, new_n25246_,
    new_n25247_, new_n25248_, new_n25249_, new_n25250_, new_n25251_,
    new_n25252_, new_n25253_, new_n25254_, new_n25255_, new_n25256_,
    new_n25257_, new_n25258_, new_n25259_, new_n25260_, new_n25261_,
    new_n25262_, new_n25263_, new_n25264_, new_n25265_, new_n25266_,
    new_n25267_, new_n25268_, new_n25269_, new_n25270_, new_n25271_,
    new_n25272_, new_n25273_, new_n25274_, new_n25275_, new_n25276_,
    new_n25277_, new_n25278_, new_n25279_, new_n25280_, new_n25281_,
    new_n25282_, new_n25283_, new_n25284_, new_n25285_, new_n25286_,
    new_n25287_, new_n25288_, new_n25289_, new_n25290_, new_n25291_,
    new_n25292_, new_n25293_, new_n25294_, new_n25295_, new_n25296_,
    new_n25297_, new_n25298_, new_n25299_, new_n25300_, new_n25301_,
    new_n25302_, new_n25303_, new_n25304_, new_n25305_, new_n25306_,
    new_n25307_, new_n25308_, new_n25309_, new_n25310_, new_n25311_,
    new_n25312_, new_n25313_, new_n25314_, new_n25315_, new_n25316_,
    new_n25317_, new_n25318_, new_n25319_, new_n25320_, new_n25321_,
    new_n25322_, new_n25323_, new_n25324_, new_n25325_, new_n25326_,
    new_n25327_, new_n25328_, new_n25329_, new_n25330_, new_n25331_,
    new_n25332_, new_n25333_, new_n25334_, new_n25335_, new_n25336_,
    new_n25337_, new_n25338_, new_n25339_, new_n25341_, new_n25342_,
    new_n25343_, new_n25344_, new_n25345_, new_n25346_, new_n25347_,
    new_n25348_, new_n25349_, new_n25350_, new_n25351_, new_n25352_,
    new_n25353_, new_n25354_, new_n25355_, new_n25356_, new_n25357_,
    new_n25358_, new_n25359_, new_n25360_, new_n25361_, new_n25362_,
    new_n25363_, new_n25364_, new_n25365_, new_n25366_, new_n25367_,
    new_n25368_, new_n25369_, new_n25370_, new_n25371_, new_n25372_,
    new_n25373_, new_n25374_, new_n25375_, new_n25376_, new_n25377_,
    new_n25378_, new_n25379_, new_n25380_, new_n25381_, new_n25382_,
    new_n25383_, new_n25384_, new_n25385_, new_n25386_, new_n25387_,
    new_n25388_, new_n25389_, new_n25390_, new_n25391_, new_n25392_,
    new_n25393_, new_n25394_, new_n25395_, new_n25396_, new_n25397_,
    new_n25398_, new_n25399_, new_n25400_, new_n25401_, new_n25402_,
    new_n25403_, new_n25404_, new_n25405_, new_n25406_, new_n25407_,
    new_n25408_, new_n25409_, new_n25410_, new_n25411_, new_n25412_,
    new_n25413_, new_n25414_, new_n25415_, new_n25416_, new_n25417_,
    new_n25418_, new_n25419_, new_n25420_, new_n25421_, new_n25422_,
    new_n25423_, new_n25424_, new_n25425_, new_n25426_, new_n25427_,
    new_n25428_, new_n25429_, new_n25430_, new_n25431_, new_n25432_,
    new_n25433_, new_n25434_, new_n25435_, new_n25436_, new_n25437_,
    new_n25438_, new_n25439_, new_n25440_, new_n25441_, new_n25442_,
    new_n25443_, new_n25444_, new_n25445_, new_n25446_, new_n25447_,
    new_n25448_, new_n25449_, new_n25450_, new_n25451_, new_n25452_,
    new_n25453_, new_n25454_, new_n25455_, new_n25456_, new_n25457_,
    new_n25458_, new_n25459_, new_n25460_, new_n25461_, new_n25462_,
    new_n25463_, new_n25464_, new_n25465_, new_n25466_, new_n25467_,
    new_n25468_, new_n25469_, new_n25470_, new_n25471_, new_n25472_,
    new_n25473_, new_n25474_, new_n25476_, new_n25477_, new_n25478_,
    new_n25479_, new_n25480_, new_n25481_, new_n25483_, new_n25484_,
    new_n25485_, new_n25486_, new_n25487_, new_n25488_, new_n25489_,
    new_n25490_, new_n25491_, new_n25492_, new_n25493_, new_n25494_,
    new_n25495_, new_n25496_, new_n25497_, new_n25498_, new_n25499_,
    new_n25500_, new_n25501_, new_n25502_, new_n25503_, new_n25504_,
    new_n25505_, new_n25506_, new_n25507_, new_n25508_, new_n25509_,
    new_n25510_, new_n25511_, new_n25512_, new_n25513_, new_n25514_,
    new_n25515_, new_n25516_, new_n25517_, new_n25518_, new_n25519_,
    new_n25520_, new_n25521_, new_n25522_, new_n25523_, new_n25524_,
    new_n25525_, new_n25526_, new_n25527_, new_n25528_, new_n25529_,
    new_n25530_, new_n25531_, new_n25532_, new_n25533_, new_n25534_,
    new_n25535_, new_n25536_, new_n25537_, new_n25538_, new_n25539_,
    new_n25540_, new_n25541_, new_n25542_, new_n25543_, new_n25544_,
    new_n25545_, new_n25546_, new_n25547_, new_n25548_, new_n25549_,
    new_n25550_, new_n25551_, new_n25552_, new_n25553_, new_n25554_,
    new_n25555_, new_n25556_, new_n25557_, new_n25558_, new_n25559_,
    new_n25560_, new_n25561_, new_n25562_, new_n25563_, new_n25564_,
    new_n25565_, new_n25566_, new_n25567_, new_n25568_, new_n25569_,
    new_n25570_, new_n25571_, new_n25572_, new_n25573_, new_n25574_,
    new_n25575_, new_n25576_, new_n25577_, new_n25578_, new_n25579_,
    new_n25580_, new_n25581_, new_n25582_, new_n25583_, new_n25584_,
    new_n25585_, new_n25586_, new_n25587_, new_n25588_, new_n25589_,
    new_n25590_, new_n25591_, new_n25592_, new_n25593_, new_n25594_,
    new_n25595_, new_n25596_, new_n25597_, new_n25598_, new_n25599_,
    new_n25600_, new_n25601_, new_n25602_, new_n25603_, new_n25604_,
    new_n25605_, new_n25606_, new_n25607_, new_n25608_, new_n25609_,
    new_n25610_, new_n25611_, new_n25612_, new_n25613_, new_n25614_,
    new_n25615_, new_n25616_, new_n25617_, new_n25618_, new_n25619_,
    new_n25620_, new_n25621_, new_n25622_, new_n25623_, new_n25624_,
    new_n25625_, new_n25626_, new_n25627_, new_n25628_, new_n25629_,
    new_n25630_, new_n25631_, new_n25632_, new_n25633_, new_n25634_,
    new_n25635_, new_n25636_, new_n25637_, new_n25638_, new_n25639_,
    new_n25640_, new_n25641_, new_n25642_, new_n25643_, new_n25644_,
    new_n25645_, new_n25646_, new_n25647_, new_n25648_, new_n25649_,
    new_n25651_, new_n25652_, new_n25653_, new_n25654_, new_n25655_,
    new_n25656_, new_n25657_, new_n25658_, new_n25659_, new_n25660_,
    new_n25661_, new_n25662_, new_n25663_, new_n25664_, new_n25665_,
    new_n25666_, new_n25667_, new_n25668_, new_n25669_, new_n25670_,
    new_n25671_, new_n25672_, new_n25673_, new_n25674_, new_n25675_,
    new_n25676_, new_n25677_, new_n25678_, new_n25679_, new_n25680_,
    new_n25681_, new_n25682_, new_n25683_, new_n25684_, new_n25685_,
    new_n25686_, new_n25687_, new_n25688_, new_n25689_, new_n25690_,
    new_n25691_, new_n25692_, new_n25693_, new_n25694_, new_n25695_,
    new_n25696_, new_n25697_, new_n25698_, new_n25699_, new_n25700_,
    new_n25701_, new_n25702_, new_n25703_, new_n25704_, new_n25705_,
    new_n25706_, new_n25707_, new_n25708_, new_n25709_, new_n25710_,
    new_n25711_, new_n25712_, new_n25713_, new_n25714_, new_n25715_,
    new_n25716_, new_n25717_, new_n25718_, new_n25719_, new_n25720_,
    new_n25721_, new_n25722_, new_n25723_, new_n25724_, new_n25725_,
    new_n25726_, new_n25727_, new_n25728_, new_n25729_, new_n25730_,
    new_n25731_, new_n25732_, new_n25733_, new_n25734_, new_n25735_,
    new_n25736_, new_n25737_, new_n25738_, new_n25739_, new_n25740_,
    new_n25741_, new_n25742_, new_n25743_, new_n25744_, new_n25745_,
    new_n25746_, new_n25747_, new_n25748_, new_n25749_, new_n25750_,
    new_n25751_, new_n25752_, new_n25753_, new_n25754_, new_n25755_,
    new_n25756_, new_n25757_, new_n25758_, new_n25759_, new_n25760_,
    new_n25761_, new_n25762_, new_n25763_, new_n25764_, new_n25765_,
    new_n25766_, new_n25767_, new_n25768_, new_n25769_, new_n25770_,
    new_n25771_, new_n25772_, new_n25773_, new_n25774_, new_n25775_,
    new_n25776_, new_n25777_, new_n25778_, new_n25779_, new_n25780_,
    new_n25781_, new_n25782_, new_n25783_, new_n25784_, new_n25785_,
    new_n25786_, new_n25787_, new_n25788_, new_n25789_, new_n25790_,
    new_n25791_, new_n25792_, new_n25793_, new_n25794_, new_n25795_,
    new_n25796_, new_n25797_, new_n25798_, new_n25799_, new_n25800_,
    new_n25801_, new_n25802_, new_n25803_, new_n25804_, new_n25805_,
    new_n25806_, new_n25807_, new_n25808_, new_n25809_, new_n25810_,
    new_n25811_, new_n25812_, new_n25813_, new_n25814_, new_n25815_,
    new_n25816_, new_n25817_, new_n25818_, new_n25819_, new_n25820_,
    new_n25821_, new_n25822_, new_n25823_, new_n25824_, new_n25825_,
    new_n25826_, new_n25827_, new_n25828_, new_n25829_, new_n25830_,
    new_n25831_, new_n25832_, new_n25833_, new_n25834_, new_n25835_,
    new_n25836_, new_n25837_, new_n25838_, new_n25839_, new_n25840_,
    new_n25841_, new_n25842_, new_n25843_, new_n25844_, new_n25845_,
    new_n25846_, new_n25847_, new_n25848_, new_n25849_, new_n25850_,
    new_n25851_, new_n25852_, new_n25853_, new_n25854_, new_n25855_,
    new_n25856_, new_n25857_, new_n25858_, new_n25859_, new_n25860_,
    new_n25861_, new_n25862_, new_n25863_, new_n25864_, new_n25865_,
    new_n25866_, new_n25867_, new_n25868_, new_n25869_, new_n25870_,
    new_n25871_, new_n25872_, new_n25873_, new_n25874_, new_n25875_,
    new_n25876_, new_n25877_, new_n25878_, new_n25880_, new_n25881_,
    new_n25882_, new_n25883_, new_n25884_, new_n25885_, new_n25886_,
    new_n25887_, new_n25888_, new_n25889_, new_n25890_, new_n25891_,
    new_n25892_, new_n25893_, new_n25894_, new_n25895_, new_n25896_,
    new_n25897_, new_n25898_, new_n25899_, new_n25900_, new_n25901_,
    new_n25902_, new_n25903_, new_n25904_, new_n25905_, new_n25906_,
    new_n25907_, new_n25908_, new_n25909_, new_n25910_, new_n25911_,
    new_n25912_, new_n25913_, new_n25914_, new_n25915_, new_n25916_,
    new_n25917_, new_n25918_, new_n25919_, new_n25920_, new_n25921_,
    new_n25922_, new_n25923_, new_n25924_, new_n25925_, new_n25926_,
    new_n25927_, new_n25928_, new_n25929_, new_n25930_, new_n25931_,
    new_n25932_, new_n25933_, new_n25934_, new_n25935_, new_n25936_,
    new_n25937_, new_n25938_, new_n25939_, new_n25941_, new_n25942_,
    new_n25943_, new_n25944_, new_n25945_, new_n25946_, new_n25947_,
    new_n25948_, new_n25949_, new_n25950_, new_n25951_, new_n25952_,
    new_n25953_, new_n25954_, new_n25955_, new_n25956_, new_n25957_,
    new_n25958_, new_n25959_, new_n25960_, new_n25961_, new_n25962_,
    new_n25963_, new_n25964_, new_n25965_, new_n25966_, new_n25967_,
    new_n25968_, new_n25969_, new_n25970_, new_n25971_, new_n25972_,
    new_n25973_, new_n25974_, new_n25975_, new_n25976_, new_n25977_,
    new_n25978_, new_n25979_, new_n25980_, new_n25981_, new_n25982_,
    new_n25983_, new_n25984_, new_n25985_, new_n25986_, new_n25987_,
    new_n25988_, new_n25989_, new_n25990_, new_n25991_, new_n25992_,
    new_n25993_, new_n25994_, new_n25995_, new_n25996_, new_n25997_,
    new_n25998_, new_n25999_, new_n26000_, new_n26001_, new_n26002_,
    new_n26003_, new_n26004_, new_n26005_, new_n26006_, new_n26007_,
    new_n26008_, new_n26009_, new_n26010_, new_n26011_, new_n26012_,
    new_n26013_, new_n26014_, new_n26015_, new_n26016_, new_n26017_,
    new_n26018_, new_n26019_, new_n26020_, new_n26021_, new_n26022_,
    new_n26023_, new_n26024_, new_n26025_, new_n26026_, new_n26027_,
    new_n26028_, new_n26029_, new_n26030_, new_n26031_, new_n26032_,
    new_n26033_, new_n26034_, new_n26035_, new_n26036_, new_n26037_,
    new_n26038_, new_n26039_, new_n26040_, new_n26041_, new_n26042_,
    new_n26043_, new_n26044_, new_n26045_, new_n26046_, new_n26047_,
    new_n26048_, new_n26049_, new_n26050_, new_n26051_, new_n26052_,
    new_n26053_, new_n26054_, new_n26055_, new_n26056_, new_n26057_,
    new_n26058_, new_n26059_, new_n26060_, new_n26061_, new_n26062_,
    new_n26063_, new_n26064_, new_n26065_, new_n26066_, new_n26067_,
    new_n26068_, new_n26069_, new_n26070_, new_n26071_, new_n26072_,
    new_n26073_, new_n26074_, new_n26075_, new_n26076_, new_n26077_,
    new_n26078_, new_n26079_, new_n26080_, new_n26081_, new_n26082_,
    new_n26083_, new_n26084_, new_n26085_, new_n26086_, new_n26087_,
    new_n26088_, new_n26089_, new_n26090_, new_n26091_, new_n26092_,
    new_n26093_, new_n26094_, new_n26095_, new_n26096_, new_n26097_,
    new_n26098_, new_n26099_, new_n26100_, new_n26101_, new_n26102_,
    new_n26103_, new_n26104_, new_n26105_, new_n26106_, new_n26107_,
    new_n26108_, new_n26109_, new_n26110_, new_n26111_, new_n26112_,
    new_n26113_, new_n26114_, new_n26115_, new_n26116_, new_n26117_,
    new_n26118_, new_n26119_, new_n26120_, new_n26121_, new_n26122_,
    new_n26123_, new_n26124_, new_n26125_, new_n26126_, new_n26127_,
    new_n26128_, new_n26129_, new_n26130_, new_n26131_, new_n26132_,
    new_n26133_, new_n26134_, new_n26135_, new_n26136_, new_n26137_,
    new_n26138_, new_n26139_, new_n26140_, new_n26141_, new_n26142_,
    new_n26143_, new_n26144_, new_n26145_, new_n26146_, new_n26147_,
    new_n26148_, new_n26149_, new_n26150_, new_n26151_, new_n26152_,
    new_n26153_, new_n26154_, new_n26155_, new_n26156_, new_n26157_,
    new_n26158_, new_n26159_, new_n26160_, new_n26161_, new_n26162_,
    new_n26163_, new_n26164_, new_n26165_, new_n26166_, new_n26167_,
    new_n26168_, new_n26169_, new_n26170_, new_n26171_, new_n26172_,
    new_n26173_, new_n26174_, new_n26175_, new_n26176_, new_n26177_,
    new_n26178_, new_n26179_, new_n26180_, new_n26181_, new_n26182_,
    new_n26183_, new_n26184_, new_n26185_, new_n26186_, new_n26187_,
    new_n26188_, new_n26189_, new_n26190_, new_n26191_, new_n26192_,
    new_n26193_, new_n26194_, new_n26195_, new_n26196_, new_n26197_,
    new_n26198_, new_n26199_, new_n26200_, new_n26201_, new_n26202_,
    new_n26203_, new_n26204_, new_n26205_, new_n26206_, new_n26207_,
    new_n26208_, new_n26209_, new_n26210_, new_n26211_, new_n26212_,
    new_n26213_, new_n26214_, new_n26215_, new_n26216_, new_n26217_,
    new_n26218_, new_n26219_, new_n26220_, new_n26221_, new_n26222_,
    new_n26223_, new_n26224_, new_n26225_, new_n26226_, new_n26227_,
    new_n26228_, new_n26229_, new_n26230_, new_n26231_, new_n26232_,
    new_n26233_, new_n26234_, new_n26235_, new_n26236_, new_n26237_,
    new_n26238_, new_n26239_, new_n26240_, new_n26241_, new_n26242_,
    new_n26243_, new_n26244_, new_n26245_, new_n26246_, new_n26247_,
    new_n26248_, new_n26249_, new_n26251_, new_n26252_, new_n26253_,
    new_n26254_, new_n26255_, new_n26256_, new_n26257_, new_n26258_,
    new_n26259_, new_n26260_, new_n26261_, new_n26262_, new_n26263_,
    new_n26264_, new_n26265_, new_n26266_, new_n26267_, new_n26268_,
    new_n26269_, new_n26270_, new_n26271_, new_n26272_, new_n26273_,
    new_n26274_, new_n26275_, new_n26276_, new_n26277_, new_n26278_,
    new_n26279_, new_n26280_, new_n26281_, new_n26282_, new_n26283_,
    new_n26284_, new_n26285_, new_n26286_, new_n26287_, new_n26288_,
    new_n26289_, new_n26290_, new_n26291_, new_n26292_, new_n26293_,
    new_n26294_, new_n26295_, new_n26296_, new_n26297_, new_n26298_,
    new_n26299_, new_n26300_, new_n26301_, new_n26302_, new_n26303_,
    new_n26304_, new_n26305_, new_n26306_, new_n26307_, new_n26308_,
    new_n26309_, new_n26310_, new_n26311_, new_n26312_, new_n26313_,
    new_n26314_, new_n26315_, new_n26316_, new_n26317_, new_n26318_,
    new_n26319_, new_n26320_, new_n26321_, new_n26322_, new_n26323_,
    new_n26324_, new_n26325_, new_n26326_, new_n26327_, new_n26328_,
    new_n26329_, new_n26330_, new_n26331_, new_n26332_, new_n26333_,
    new_n26334_, new_n26335_, new_n26336_, new_n26337_, new_n26338_,
    new_n26339_, new_n26340_, new_n26341_, new_n26342_, new_n26343_,
    new_n26344_, new_n26345_, new_n26346_, new_n26347_, new_n26348_,
    new_n26349_, new_n26350_, new_n26351_, new_n26352_, new_n26353_,
    new_n26354_, new_n26355_, new_n26356_, new_n26357_, new_n26358_,
    new_n26359_, new_n26360_, new_n26361_, new_n26362_, new_n26363_,
    new_n26364_, new_n26365_, new_n26366_, new_n26367_, new_n26368_,
    new_n26369_, new_n26370_, new_n26371_, new_n26372_, new_n26373_,
    new_n26374_, new_n26375_, new_n26376_, new_n26377_, new_n26378_,
    new_n26379_, new_n26380_, new_n26381_, new_n26382_, new_n26383_,
    new_n26384_, new_n26385_, new_n26386_, new_n26387_, new_n26388_,
    new_n26389_, new_n26390_, new_n26391_, new_n26392_, new_n26393_,
    new_n26394_, new_n26395_, new_n26396_, new_n26397_, new_n26398_,
    new_n26399_, new_n26400_, new_n26401_, new_n26402_, new_n26403_,
    new_n26404_, new_n26405_, new_n26406_, new_n26407_, new_n26408_,
    new_n26409_, new_n26410_, new_n26411_, new_n26412_, new_n26413_,
    new_n26414_, new_n26415_, new_n26416_, new_n26417_, new_n26418_,
    new_n26419_, new_n26420_, new_n26421_, new_n26422_, new_n26423_,
    new_n26424_, new_n26425_, new_n26426_, new_n26427_, new_n26428_,
    new_n26429_, new_n26430_, new_n26431_, new_n26432_, new_n26433_,
    new_n26434_, new_n26435_, new_n26436_, new_n26437_, new_n26438_,
    new_n26439_, new_n26440_, new_n26441_, new_n26442_, new_n26443_,
    new_n26444_, new_n26446_, new_n26447_, new_n26448_, new_n26449_,
    new_n26450_, new_n26451_, new_n26452_, new_n26453_, new_n26454_,
    new_n26455_, new_n26456_, new_n26457_, new_n26458_, new_n26459_,
    new_n26460_, new_n26461_, new_n26462_, new_n26463_, new_n26464_,
    new_n26465_, new_n26466_, new_n26467_, new_n26468_, new_n26469_,
    new_n26470_, new_n26471_, new_n26472_, new_n26473_, new_n26474_,
    new_n26475_, new_n26476_, new_n26477_, new_n26478_, new_n26479_,
    new_n26480_, new_n26481_, new_n26482_, new_n26483_, new_n26484_,
    new_n26485_, new_n26486_, new_n26487_, new_n26488_, new_n26489_,
    new_n26490_, new_n26491_, new_n26492_, new_n26493_, new_n26494_,
    new_n26495_, new_n26496_, new_n26497_, new_n26499_, new_n26500_,
    new_n26501_, new_n26502_, new_n26503_, new_n26504_, new_n26505_,
    new_n26506_, new_n26507_, new_n26508_, new_n26509_, new_n26510_,
    new_n26511_, new_n26512_, new_n26513_, new_n26514_, new_n26515_,
    new_n26516_, new_n26517_, new_n26518_, new_n26519_, new_n26520_,
    new_n26521_, new_n26522_, new_n26523_, new_n26524_, new_n26525_,
    new_n26526_, new_n26527_, new_n26528_, new_n26529_, new_n26530_,
    new_n26531_, new_n26532_, new_n26533_, new_n26534_, new_n26535_,
    new_n26536_, new_n26537_, new_n26538_, new_n26539_, new_n26540_,
    new_n26541_, new_n26542_, new_n26543_, new_n26544_, new_n26545_,
    new_n26546_, new_n26547_, new_n26548_, new_n26549_, new_n26550_,
    new_n26551_, new_n26552_, new_n26553_, new_n26554_, new_n26555_,
    new_n26556_, new_n26557_, new_n26558_, new_n26559_, new_n26560_,
    new_n26561_, new_n26562_, new_n26563_, new_n26564_, new_n26565_,
    new_n26566_, new_n26567_, new_n26568_, new_n26569_, new_n26570_,
    new_n26571_, new_n26572_, new_n26573_, new_n26574_, new_n26575_,
    new_n26576_, new_n26577_, new_n26578_, new_n26579_, new_n26580_,
    new_n26581_, new_n26582_, new_n26583_, new_n26584_, new_n26585_,
    new_n26586_, new_n26587_, new_n26588_, new_n26589_, new_n26590_,
    new_n26591_, new_n26592_, new_n26593_, new_n26594_, new_n26595_,
    new_n26596_, new_n26597_, new_n26598_, new_n26599_, new_n26600_,
    new_n26601_, new_n26602_, new_n26603_, new_n26604_, new_n26605_,
    new_n26606_, new_n26607_, new_n26608_, new_n26609_, new_n26610_,
    new_n26611_, new_n26612_, new_n26613_, new_n26614_, new_n26615_,
    new_n26616_, new_n26617_, new_n26618_, new_n26619_, new_n26620_,
    new_n26621_, new_n26622_, new_n26623_, new_n26624_, new_n26625_,
    new_n26626_, new_n26627_, new_n26628_, new_n26629_, new_n26630_,
    new_n26631_, new_n26632_, new_n26633_, new_n26634_, new_n26635_,
    new_n26636_, new_n26637_, new_n26638_, new_n26639_, new_n26640_,
    new_n26641_, new_n26642_, new_n26643_, new_n26644_, new_n26645_,
    new_n26646_, new_n26647_, new_n26648_, new_n26649_, new_n26650_,
    new_n26651_, new_n26652_, new_n26653_, new_n26654_, new_n26655_,
    new_n26656_, new_n26657_, new_n26658_, new_n26659_, new_n26660_,
    new_n26661_, new_n26662_, new_n26663_, new_n26664_, new_n26665_,
    new_n26666_, new_n26667_, new_n26668_, new_n26669_, new_n26670_,
    new_n26671_, new_n26672_, new_n26673_, new_n26674_, new_n26675_,
    new_n26676_, new_n26677_, new_n26678_, new_n26679_, new_n26680_,
    new_n26681_, new_n26682_, new_n26683_, new_n26684_, new_n26685_,
    new_n26686_, new_n26687_, new_n26688_, new_n26689_, new_n26690_,
    new_n26691_, new_n26692_, new_n26693_, new_n26694_, new_n26695_,
    new_n26696_, new_n26697_, new_n26698_, new_n26699_, new_n26700_,
    new_n26701_, new_n26702_, new_n26703_, new_n26704_, new_n26705_,
    new_n26706_, new_n26707_, new_n26708_, new_n26709_, new_n26710_,
    new_n26711_, new_n26712_, new_n26713_, new_n26714_, new_n26715_,
    new_n26716_, new_n26717_, new_n26718_, new_n26719_, new_n26720_,
    new_n26722_, new_n26723_, new_n26724_, new_n26725_, new_n26726_,
    new_n26727_, new_n26728_, new_n26729_, new_n26730_, new_n26731_,
    new_n26732_, new_n26733_, new_n26734_, new_n26735_, new_n26736_,
    new_n26737_, new_n26738_, new_n26739_, new_n26740_, new_n26741_,
    new_n26742_, new_n26743_, new_n26744_, new_n26745_, new_n26746_,
    new_n26747_, new_n26748_, new_n26749_, new_n26750_, new_n26751_,
    new_n26752_, new_n26753_, new_n26754_, new_n26756_, new_n26757_,
    new_n26758_, new_n26759_, new_n26760_, new_n26761_, new_n26762_,
    new_n26763_, new_n26764_, new_n26765_, new_n26766_, new_n26767_,
    new_n26768_, new_n26769_, new_n26770_, new_n26771_, new_n26772_,
    new_n26773_, new_n26774_, new_n26775_, new_n26776_, new_n26777_,
    new_n26778_, new_n26779_, new_n26780_, new_n26781_, new_n26782_,
    new_n26783_, new_n26784_, new_n26785_, new_n26786_, new_n26787_,
    new_n26788_, new_n26789_, new_n26790_, new_n26791_, new_n26792_,
    new_n26793_, new_n26794_, new_n26795_, new_n26796_, new_n26797_,
    new_n26798_, new_n26799_, new_n26800_, new_n26801_, new_n26802_,
    new_n26803_, new_n26804_, new_n26805_, new_n26806_, new_n26807_,
    new_n26808_, new_n26809_, new_n26810_, new_n26811_, new_n26812_,
    new_n26813_, new_n26814_, new_n26815_, new_n26816_, new_n26817_,
    new_n26818_, new_n26819_, new_n26820_, new_n26821_, new_n26822_,
    new_n26823_, new_n26824_, new_n26825_, new_n26826_, new_n26827_,
    new_n26828_, new_n26829_, new_n26830_, new_n26831_, new_n26832_,
    new_n26833_, new_n26834_, new_n26835_, new_n26836_, new_n26837_,
    new_n26838_, new_n26839_, new_n26840_, new_n26841_, new_n26842_,
    new_n26843_, new_n26844_, new_n26845_, new_n26846_, new_n26847_,
    new_n26848_, new_n26849_, new_n26850_, new_n26851_, new_n26852_,
    new_n26853_, new_n26854_, new_n26855_, new_n26856_, new_n26857_,
    new_n26858_, new_n26859_, new_n26860_, new_n26861_, new_n26862_,
    new_n26863_, new_n26864_, new_n26865_, new_n26866_, new_n26867_,
    new_n26868_, new_n26869_, new_n26870_, new_n26871_, new_n26872_,
    new_n26873_, new_n26874_, new_n26875_, new_n26876_, new_n26877_,
    new_n26878_, new_n26879_, new_n26880_, new_n26881_, new_n26882_,
    new_n26883_, new_n26884_, new_n26885_, new_n26886_, new_n26887_,
    new_n26888_, new_n26889_, new_n26890_, new_n26891_, new_n26892_,
    new_n26893_, new_n26894_, new_n26895_, new_n26896_, new_n26897_,
    new_n26898_, new_n26899_, new_n26900_, new_n26901_, new_n26902_,
    new_n26903_, new_n26904_, new_n26905_, new_n26906_, new_n26907_,
    new_n26908_, new_n26909_, new_n26910_, new_n26911_, new_n26912_,
    new_n26913_, new_n26914_, new_n26915_, new_n26916_, new_n26917_,
    new_n26918_, new_n26919_, new_n26920_, new_n26921_, new_n26922_,
    new_n26923_, new_n26925_, new_n26926_, new_n26927_, new_n26928_,
    new_n26929_, new_n26930_, new_n26931_, new_n26932_, new_n26933_,
    new_n26934_, new_n26935_, new_n26936_, new_n26937_, new_n26938_,
    new_n26939_, new_n26940_, new_n26941_, new_n26942_, new_n26943_,
    new_n26944_, new_n26945_, new_n26946_, new_n26947_, new_n26948_,
    new_n26949_, new_n26950_, new_n26951_, new_n26952_, new_n26953_,
    new_n26954_, new_n26955_, new_n26956_, new_n26957_, new_n26958_,
    new_n26959_, new_n26960_, new_n26961_, new_n26962_, new_n26963_,
    new_n26964_, new_n26965_, new_n26966_, new_n26967_, new_n26968_,
    new_n26969_, new_n26970_, new_n26971_, new_n26972_, new_n26973_,
    new_n26974_, new_n26975_, new_n26976_, new_n26977_, new_n26978_,
    new_n26979_, new_n26980_, new_n26981_, new_n26982_, new_n26983_,
    new_n26984_, new_n26985_, new_n26986_, new_n26987_, new_n26988_,
    new_n26989_, new_n26990_, new_n26991_, new_n26992_, new_n26993_,
    new_n26994_, new_n26995_, new_n26996_, new_n26997_, new_n26998_,
    new_n26999_, new_n27000_, new_n27001_, new_n27002_, new_n27003_,
    new_n27004_, new_n27005_, new_n27006_, new_n27007_, new_n27008_,
    new_n27009_, new_n27010_, new_n27011_, new_n27012_, new_n27013_,
    new_n27014_, new_n27015_, new_n27016_, new_n27017_, new_n27018_,
    new_n27019_, new_n27020_, new_n27021_, new_n27022_, new_n27023_,
    new_n27024_, new_n27025_, new_n27026_, new_n27027_, new_n27028_,
    new_n27029_, new_n27030_, new_n27031_, new_n27032_, new_n27033_,
    new_n27034_, new_n27035_, new_n27036_, new_n27037_, new_n27038_,
    new_n27039_, new_n27040_, new_n27041_, new_n27042_, new_n27043_,
    new_n27044_, new_n27045_, new_n27046_, new_n27047_, new_n27048_,
    new_n27049_, new_n27050_, new_n27051_, new_n27052_, new_n27053_,
    new_n27054_, new_n27055_, new_n27056_, new_n27057_, new_n27058_,
    new_n27059_, new_n27060_, new_n27061_, new_n27062_, new_n27063_,
    new_n27064_, new_n27065_, new_n27066_, new_n27067_, new_n27068_,
    new_n27069_, new_n27070_, new_n27071_, new_n27072_, new_n27073_,
    new_n27074_, new_n27075_, new_n27076_, new_n27077_, new_n27078_,
    new_n27079_, new_n27080_, new_n27081_, new_n27082_, new_n27083_,
    new_n27084_, new_n27085_, new_n27086_, new_n27087_, new_n27088_,
    new_n27089_, new_n27090_, new_n27091_, new_n27092_, new_n27093_,
    new_n27094_, new_n27095_, new_n27096_, new_n27098_, new_n27099_,
    new_n27100_, new_n27101_, new_n27102_, new_n27103_, new_n27104_,
    new_n27105_, new_n27106_, new_n27107_, new_n27108_, new_n27109_,
    new_n27110_, new_n27111_, new_n27112_, new_n27113_, new_n27114_,
    new_n27115_, new_n27116_, new_n27117_, new_n27118_, new_n27119_,
    new_n27120_, new_n27121_, new_n27122_, new_n27123_, new_n27124_,
    new_n27125_, new_n27126_, new_n27127_, new_n27128_, new_n27129_,
    new_n27130_, new_n27131_, new_n27132_, new_n27133_, new_n27134_,
    new_n27135_, new_n27136_, new_n27137_, new_n27138_, new_n27139_,
    new_n27140_, new_n27141_, new_n27142_, new_n27143_, new_n27144_,
    new_n27145_, new_n27146_, new_n27147_, new_n27148_, new_n27149_,
    new_n27150_, new_n27151_, new_n27152_, new_n27153_, new_n27154_,
    new_n27155_, new_n27156_, new_n27157_, new_n27158_, new_n27159_,
    new_n27160_, new_n27161_, new_n27162_, new_n27163_, new_n27164_,
    new_n27165_, new_n27166_, new_n27167_, new_n27168_, new_n27169_,
    new_n27170_, new_n27171_, new_n27172_, new_n27173_, new_n27174_,
    new_n27175_, new_n27176_, new_n27177_, new_n27178_, new_n27179_,
    new_n27180_, new_n27181_, new_n27182_, new_n27183_, new_n27184_,
    new_n27185_, new_n27186_, new_n27187_, new_n27188_, new_n27189_,
    new_n27190_, new_n27191_, new_n27192_, new_n27193_, new_n27194_,
    new_n27195_, new_n27196_, new_n27197_, new_n27198_, new_n27199_,
    new_n27200_, new_n27201_, new_n27202_, new_n27203_, new_n27204_,
    new_n27205_, new_n27206_, new_n27207_, new_n27208_, new_n27209_,
    new_n27210_, new_n27211_, new_n27212_, new_n27213_, new_n27214_,
    new_n27215_, new_n27216_, new_n27217_, new_n27218_, new_n27219_,
    new_n27220_, new_n27221_, new_n27222_, new_n27223_, new_n27224_,
    new_n27225_, new_n27226_, new_n27227_, new_n27228_, new_n27229_,
    new_n27230_, new_n27231_, new_n27232_, new_n27233_, new_n27234_,
    new_n27235_, new_n27236_, new_n27237_, new_n27238_, new_n27239_,
    new_n27240_, new_n27241_, new_n27242_, new_n27243_, new_n27244_,
    new_n27245_, new_n27246_, new_n27247_, new_n27248_, new_n27249_,
    new_n27250_, new_n27251_, new_n27252_, new_n27253_, new_n27254_,
    new_n27256_, new_n27257_, new_n27258_, new_n27259_, new_n27260_,
    new_n27261_, new_n27262_, new_n27263_, new_n27264_, new_n27265_,
    new_n27266_, new_n27267_, new_n27268_, new_n27269_, new_n27270_,
    new_n27271_, new_n27272_, new_n27273_, new_n27274_, new_n27275_,
    new_n27276_, new_n27277_, new_n27278_, new_n27279_, new_n27280_,
    new_n27281_, new_n27282_, new_n27283_, new_n27284_, new_n27285_,
    new_n27286_, new_n27287_, new_n27288_, new_n27289_, new_n27290_,
    new_n27291_, new_n27292_, new_n27293_, new_n27294_, new_n27295_,
    new_n27296_, new_n27297_, new_n27298_, new_n27299_, new_n27300_,
    new_n27301_, new_n27302_, new_n27303_, new_n27304_, new_n27305_,
    new_n27306_, new_n27307_, new_n27308_, new_n27309_, new_n27310_,
    new_n27311_, new_n27312_, new_n27313_, new_n27314_, new_n27315_,
    new_n27316_, new_n27317_, new_n27318_, new_n27319_, new_n27320_,
    new_n27321_, new_n27322_, new_n27323_, new_n27324_, new_n27325_,
    new_n27326_, new_n27327_, new_n27328_, new_n27329_, new_n27330_,
    new_n27331_, new_n27332_, new_n27333_, new_n27334_, new_n27335_,
    new_n27336_, new_n27337_, new_n27338_, new_n27339_, new_n27340_,
    new_n27341_, new_n27342_, new_n27343_, new_n27344_, new_n27345_,
    new_n27346_, new_n27347_, new_n27348_, new_n27349_, new_n27350_,
    new_n27351_, new_n27352_, new_n27353_, new_n27354_, new_n27355_,
    new_n27356_, new_n27357_, new_n27358_, new_n27359_, new_n27360_,
    new_n27361_, new_n27362_, new_n27364_, new_n27365_, new_n27366_,
    new_n27367_, new_n27368_, new_n27369_, new_n27370_, new_n27371_,
    new_n27372_, new_n27373_, new_n27374_, new_n27375_, new_n27376_,
    new_n27377_, new_n27378_, new_n27379_, new_n27380_, new_n27381_,
    new_n27382_, new_n27383_, new_n27384_, new_n27385_, new_n27386_,
    new_n27387_, new_n27388_, new_n27389_, new_n27390_, new_n27391_,
    new_n27392_, new_n27393_, new_n27394_, new_n27395_, new_n27396_,
    new_n27397_, new_n27398_, new_n27399_, new_n27400_, new_n27401_,
    new_n27402_, new_n27403_, new_n27404_, new_n27405_, new_n27406_,
    new_n27407_, new_n27408_, new_n27409_, new_n27410_, new_n27411_,
    new_n27412_, new_n27413_, new_n27414_, new_n27415_, new_n27416_,
    new_n27417_, new_n27418_, new_n27419_, new_n27420_, new_n27421_,
    new_n27422_, new_n27423_, new_n27424_, new_n27425_, new_n27426_,
    new_n27427_, new_n27428_, new_n27429_, new_n27430_, new_n27431_,
    new_n27432_, new_n27433_, new_n27434_, new_n27435_, new_n27436_,
    new_n27437_, new_n27438_, new_n27439_, new_n27440_, new_n27441_,
    new_n27442_, new_n27443_, new_n27444_, new_n27445_, new_n27446_,
    new_n27447_, new_n27448_, new_n27449_, new_n27450_, new_n27451_,
    new_n27452_, new_n27453_, new_n27454_, new_n27455_, new_n27456_,
    new_n27457_, new_n27458_, new_n27459_, new_n27460_, new_n27461_,
    new_n27462_, new_n27463_, new_n27464_, new_n27465_, new_n27466_,
    new_n27467_, new_n27468_, new_n27469_, new_n27470_, new_n27471_,
    new_n27472_, new_n27473_, new_n27474_, new_n27475_, new_n27476_,
    new_n27477_, new_n27478_, new_n27480_, new_n27481_, new_n27482_,
    new_n27483_, new_n27485_, new_n27486_, new_n27487_, new_n27488_,
    new_n27489_, new_n27490_, new_n27491_, new_n27493_, new_n27494_,
    new_n27495_, new_n27496_, new_n27497_, new_n27498_, new_n27499_,
    new_n27500_, new_n27501_, new_n27502_, new_n27503_, new_n27504_,
    new_n27505_, new_n27506_, new_n27507_, new_n27508_, new_n27509_,
    new_n27510_, new_n27511_, new_n27512_, new_n27513_, new_n27514_,
    new_n27515_, new_n27516_, new_n27517_, new_n27519_, new_n27520_,
    new_n27521_, new_n27522_, new_n27523_, new_n27524_, new_n27525_,
    new_n27526_, new_n27527_, new_n27528_, new_n27529_, new_n27530_,
    new_n27531_, new_n27532_, new_n27533_, new_n27534_, new_n27535_,
    new_n27536_, new_n27537_, new_n27538_, new_n27539_, new_n27540_,
    new_n27541_, new_n27542_, new_n27543_, new_n27544_, new_n27545_,
    new_n27546_, new_n27547_, new_n27548_, new_n27549_, new_n27550_,
    new_n27551_, new_n27552_, new_n27553_, new_n27554_, new_n27555_,
    new_n27556_, new_n27557_, new_n27558_, new_n27559_, new_n27560_,
    new_n27561_, new_n27562_, new_n27563_, new_n27564_, new_n27565_,
    new_n27566_, new_n27567_, new_n27568_, new_n27569_, new_n27570_,
    new_n27571_, new_n27572_, new_n27573_, new_n27574_, new_n27575_,
    new_n27576_, new_n27577_, new_n27578_, new_n27579_, new_n27580_,
    new_n27581_, new_n27582_, new_n27583_, new_n27584_, new_n27585_,
    new_n27586_, new_n27587_, new_n27588_, new_n27589_, new_n27590_,
    new_n27591_, new_n27592_, new_n27593_, new_n27594_, new_n27595_,
    new_n27596_, new_n27597_, new_n27598_, new_n27599_, new_n27600_,
    new_n27601_, new_n27602_, new_n27603_, new_n27604_, new_n27605_,
    new_n27606_, new_n27607_, new_n27608_, new_n27609_, new_n27610_,
    new_n27611_, new_n27612_, new_n27613_, new_n27614_, new_n27615_,
    new_n27616_, new_n27617_, new_n27618_, new_n27619_, new_n27620_,
    new_n27621_, new_n27622_, new_n27623_, new_n27624_, new_n27625_,
    new_n27626_, new_n27627_, new_n27628_, new_n27629_, new_n27630_,
    new_n27631_, new_n27632_, new_n27633_, new_n27634_, new_n27635_,
    new_n27636_, new_n27637_, new_n27638_, new_n27639_, new_n27640_,
    new_n27641_, new_n27642_, new_n27643_, new_n27644_, new_n27645_,
    new_n27646_, new_n27647_, new_n27648_, new_n27649_, new_n27650_,
    new_n27651_, new_n27652_, new_n27653_, new_n27654_, new_n27655_,
    new_n27656_, new_n27657_, new_n27658_, new_n27659_, new_n27660_,
    new_n27661_, new_n27662_, new_n27663_, new_n27664_, new_n27665_,
    new_n27666_, new_n27667_, new_n27668_, new_n27669_, new_n27670_,
    new_n27671_, new_n27672_, new_n27673_, new_n27674_, new_n27675_,
    new_n27676_, new_n27677_, new_n27678_, new_n27679_, new_n27680_,
    new_n27681_, new_n27682_, new_n27683_, new_n27684_, new_n27685_,
    new_n27686_, new_n27687_, new_n27689_, new_n27690_, new_n27691_,
    new_n27692_, new_n27693_, new_n27694_, new_n27695_, new_n27696_,
    new_n27697_, new_n27698_, new_n27699_, new_n27700_, new_n27701_,
    new_n27702_, new_n27703_, new_n27704_, new_n27705_, new_n27706_,
    new_n27707_, new_n27708_, new_n27709_, new_n27710_, new_n27711_,
    new_n27712_, new_n27713_, new_n27714_, new_n27715_, new_n27716_,
    new_n27717_, new_n27718_, new_n27719_, new_n27720_, new_n27721_,
    new_n27722_, new_n27723_, new_n27724_, new_n27725_, new_n27726_,
    new_n27727_, new_n27728_, new_n27729_, new_n27730_, new_n27731_,
    new_n27732_, new_n27733_, new_n27734_, new_n27735_, new_n27736_,
    new_n27737_, new_n27738_, new_n27739_, new_n27740_, new_n27741_,
    new_n27742_, new_n27743_, new_n27744_, new_n27745_, new_n27746_,
    new_n27747_, new_n27748_, new_n27749_, new_n27750_, new_n27751_,
    new_n27752_, new_n27753_, new_n27754_, new_n27755_, new_n27756_,
    new_n27757_, new_n27758_, new_n27759_, new_n27760_, new_n27761_,
    new_n27762_, new_n27763_, new_n27764_, new_n27765_, new_n27766_,
    new_n27767_, new_n27768_, new_n27769_, new_n27770_, new_n27771_,
    new_n27772_, new_n27773_, new_n27774_, new_n27775_, new_n27776_,
    new_n27777_, new_n27778_, new_n27779_, new_n27780_, new_n27781_,
    new_n27782_, new_n27783_, new_n27784_, new_n27785_, new_n27786_,
    new_n27787_, new_n27788_, new_n27789_, new_n27790_, new_n27791_,
    new_n27792_, new_n27793_, new_n27794_, new_n27795_, new_n27796_,
    new_n27797_, new_n27798_, new_n27799_, new_n27800_, new_n27801_,
    new_n27802_, new_n27803_, new_n27804_, new_n27805_, new_n27806_,
    new_n27807_, new_n27808_, new_n27809_, new_n27810_, new_n27811_,
    new_n27812_, new_n27813_, new_n27814_, new_n27815_, new_n27816_,
    new_n27817_, new_n27818_, new_n27819_, new_n27820_, new_n27821_,
    new_n27822_, new_n27823_, new_n27824_, new_n27825_, new_n27826_,
    new_n27827_, new_n27828_, new_n27829_, new_n27830_, new_n27831_,
    new_n27832_, new_n27833_, new_n27834_, new_n27835_, new_n27836_,
    new_n27837_, new_n27838_, new_n27840_, new_n27842_, new_n27844_,
    new_n27846_, new_n27848_, new_n27850_, new_n27851_, new_n27852_,
    new_n27854_, new_n27855_, new_n27856_, new_n27858_, new_n27859_,
    new_n27860_, new_n27861_, new_n27862_, new_n27863_, new_n27864_,
    new_n27865_, new_n27866_, new_n27867_, new_n27868_, new_n27869_,
    new_n27870_, new_n27871_, new_n27872_, new_n27873_, new_n27874_,
    new_n27875_, new_n27876_, new_n27877_, new_n27878_, new_n27880_,
    new_n27881_, new_n27882_, new_n27883_, new_n27884_, new_n27885_,
    new_n27886_, new_n27887_, new_n27888_, new_n27889_, new_n27890_,
    new_n27891_, new_n27892_, new_n27893_, new_n27894_, new_n27895_,
    new_n27896_, new_n27897_, new_n27898_, new_n27899_, new_n27900_,
    new_n27901_, new_n27902_, new_n27903_, new_n27904_, new_n27905_,
    new_n27906_, new_n27907_, new_n27908_, new_n27909_, new_n27910_,
    new_n27911_, new_n27912_, new_n27913_, new_n27914_, new_n27915_,
    new_n27916_, new_n27917_, new_n27918_, new_n27919_, new_n27920_,
    new_n27921_, new_n27922_, new_n27923_, new_n27924_, new_n27925_,
    new_n27926_, new_n27927_, new_n27928_, new_n27929_, new_n27930_,
    new_n27931_, new_n27932_, new_n27933_, new_n27934_, new_n27935_,
    new_n27936_, new_n27937_, new_n27938_, new_n27939_, new_n27940_,
    new_n27941_, new_n27942_, new_n27943_, new_n27944_, new_n27945_,
    new_n27946_, new_n27947_, new_n27948_, new_n27949_, new_n27950_,
    new_n27951_, new_n27952_, new_n27953_, new_n27954_, new_n27955_,
    new_n27956_, new_n27957_, new_n27958_, new_n27959_, new_n27960_,
    new_n27961_, new_n27962_, new_n27963_, new_n27964_, new_n27965_,
    new_n27966_, new_n27967_, new_n27968_, new_n27969_, new_n27970_,
    new_n27971_, new_n27972_, new_n27973_, new_n27974_, new_n27975_,
    new_n27976_, new_n27977_, new_n27978_, new_n27979_, new_n27980_,
    new_n27981_, new_n27982_, new_n27983_, new_n27984_, new_n27985_,
    new_n27986_, new_n27987_, new_n27988_, new_n27989_, new_n27990_,
    new_n27991_, new_n27992_, new_n27993_, new_n27994_, new_n27995_,
    new_n27996_, new_n27997_, new_n27998_, new_n27999_, new_n28000_,
    new_n28001_, new_n28002_, new_n28003_, new_n28004_, new_n28005_,
    new_n28006_, new_n28007_, new_n28008_, new_n28009_, new_n28010_,
    new_n28011_, new_n28012_, new_n28013_, new_n28014_, new_n28015_,
    new_n28016_, new_n28017_, new_n28018_, new_n28019_, new_n28020_,
    new_n28021_, new_n28022_, new_n28023_, new_n28024_, new_n28025_,
    new_n28026_, new_n28028_, new_n28029_, new_n28030_, new_n28031_,
    new_n28032_, new_n28033_, new_n28034_, new_n28035_, new_n28036_,
    new_n28037_, new_n28038_, new_n28039_, new_n28040_, new_n28041_,
    new_n28042_, new_n28043_, new_n28044_, new_n28045_, new_n28046_,
    new_n28047_, new_n28048_, new_n28049_, new_n28050_, new_n28051_,
    new_n28052_, new_n28053_, new_n28054_, new_n28055_, new_n28057_,
    new_n28058_, new_n28059_, new_n28060_, new_n28061_, new_n28062_,
    new_n28063_, new_n28064_, new_n28065_, new_n28066_, new_n28067_,
    new_n28068_, new_n28069_, new_n28070_, new_n28071_, new_n28072_,
    new_n28073_, new_n28074_, new_n28075_, new_n28076_, new_n28077_,
    new_n28078_, new_n28079_, new_n28080_, new_n28081_, new_n28083_,
    new_n28084_, new_n28085_, new_n28086_, new_n28087_, new_n28088_,
    new_n28089_, new_n28090_, new_n28091_, new_n28092_, new_n28093_,
    new_n28094_, new_n28095_, new_n28096_, new_n28097_, new_n28098_,
    new_n28099_, new_n28100_, new_n28101_, new_n28102_, new_n28103_,
    new_n28104_, new_n28105_, new_n28106_, new_n28107_, new_n28108_,
    new_n28109_, new_n28110_, new_n28111_, new_n28112_, new_n28113_,
    new_n28114_, new_n28115_, new_n28116_, new_n28117_, new_n28118_,
    new_n28119_, new_n28121_, new_n28122_, new_n28123_, new_n28124_,
    new_n28125_, new_n28126_, new_n28127_, new_n28128_, new_n28129_,
    new_n28130_, new_n28131_, new_n28132_, new_n28133_, new_n28134_,
    new_n28135_, new_n28136_, new_n28137_, new_n28138_, new_n28139_,
    new_n28140_, new_n28141_, new_n28142_, new_n28143_, new_n28144_,
    new_n28145_, new_n28146_, new_n28147_, new_n28148_, new_n28149_,
    new_n28150_, new_n28151_, new_n28152_, new_n28153_, new_n28154_,
    new_n28155_, new_n28156_, new_n28157_, new_n28158_, new_n28159_,
    new_n28160_, new_n28161_, new_n28162_, new_n28163_, new_n28164_,
    new_n28165_, new_n28166_, new_n28167_, new_n28168_, new_n28169_,
    new_n28170_, new_n28171_, new_n28172_, new_n28173_, new_n28174_,
    new_n28175_, new_n28176_, new_n28177_, new_n28178_, new_n28179_,
    new_n28180_, new_n28181_, new_n28182_, new_n28183_, new_n28184_,
    new_n28185_, new_n28186_, new_n28187_, new_n28188_, new_n28189_,
    new_n28190_, new_n28191_, new_n28192_, new_n28193_, new_n28194_,
    new_n28195_, new_n28196_, new_n28197_, new_n28198_, new_n28199_,
    new_n28200_, new_n28201_, new_n28202_, new_n28203_, new_n28204_,
    new_n28205_, new_n28206_, new_n28207_, new_n28208_, new_n28209_,
    new_n28210_, new_n28211_, new_n28212_, new_n28213_, new_n28214_,
    new_n28215_, new_n28216_, new_n28217_, new_n28218_, new_n28219_,
    new_n28220_, new_n28221_, new_n28222_, new_n28223_, new_n28224_,
    new_n28225_, new_n28226_, new_n28227_, new_n28228_, new_n28229_,
    new_n28230_, new_n28231_, new_n28232_, new_n28233_, new_n28234_,
    new_n28235_, new_n28236_, new_n28237_, new_n28238_, new_n28239_,
    new_n28240_, new_n28241_, new_n28242_, new_n28243_, new_n28244_,
    new_n28245_, new_n28246_, new_n28247_, new_n28248_, new_n28249_,
    new_n28250_, new_n28251_, new_n28252_, new_n28253_, new_n28254_,
    new_n28255_, new_n28256_, new_n28258_, new_n28259_, new_n28260_,
    new_n28261_, new_n28262_, new_n28263_, new_n28264_, new_n28265_,
    new_n28266_, new_n28267_, new_n28268_, new_n28269_, new_n28270_,
    new_n28271_, new_n28272_, new_n28273_, new_n28274_, new_n28275_,
    new_n28276_, new_n28277_, new_n28278_, new_n28279_, new_n28280_,
    new_n28281_, new_n28282_, new_n28283_, new_n28284_, new_n28285_,
    new_n28286_, new_n28287_, new_n28288_, new_n28289_, new_n28290_,
    new_n28291_, new_n28292_, new_n28293_, new_n28294_, new_n28295_,
    new_n28296_, new_n28297_, new_n28298_, new_n28299_, new_n28300_,
    new_n28301_, new_n28302_, new_n28303_, new_n28304_, new_n28305_,
    new_n28306_, new_n28307_, new_n28308_, new_n28309_, new_n28310_,
    new_n28311_, new_n28312_, new_n28313_, new_n28314_, new_n28315_,
    new_n28316_, new_n28317_, new_n28318_, new_n28319_, new_n28320_,
    new_n28321_, new_n28322_, new_n28323_, new_n28324_, new_n28325_,
    new_n28326_, new_n28327_, new_n28328_, new_n28329_, new_n28330_,
    new_n28331_, new_n28332_, new_n28333_, new_n28334_, new_n28335_,
    new_n28336_, new_n28337_, new_n28338_, new_n28339_, new_n28340_,
    new_n28341_, new_n28342_, new_n28343_, new_n28344_, new_n28345_,
    new_n28346_, new_n28347_, new_n28348_, new_n28349_, new_n28350_,
    new_n28351_, new_n28352_, new_n28353_, new_n28354_, new_n28355_,
    new_n28356_, new_n28357_, new_n28358_, new_n28360_, new_n28361_,
    new_n28362_, new_n28363_, new_n28364_, new_n28365_, new_n28366_,
    new_n28367_, new_n28368_, new_n28369_, new_n28370_, new_n28371_,
    new_n28372_, new_n28373_, new_n28374_, new_n28375_, new_n28376_,
    new_n28377_, new_n28378_, new_n28379_, new_n28380_, new_n28381_,
    new_n28383_, new_n28384_, new_n28385_, new_n28386_, new_n28387_,
    new_n28388_, new_n28389_, new_n28390_, new_n28391_, new_n28392_,
    new_n28393_, new_n28394_, new_n28395_, new_n28396_, new_n28397_,
    new_n28398_, new_n28399_, new_n28400_, new_n28401_, new_n28402_,
    new_n28403_, new_n28404_, new_n28405_, new_n28406_, new_n28407_,
    new_n28408_, new_n28409_, new_n28411_, new_n28412_, new_n28413_,
    new_n28414_, new_n28415_, new_n28416_, new_n28417_, new_n28418_,
    new_n28419_, new_n28420_, new_n28421_, new_n28422_, new_n28423_,
    new_n28424_, new_n28425_, new_n28426_, new_n28427_, new_n28428_,
    new_n28429_, new_n28430_, new_n28431_, new_n28432_, new_n28433_,
    new_n28434_, new_n28435_, new_n28436_, new_n28437_, new_n28438_,
    new_n28440_, new_n28441_, new_n28442_, new_n28443_, new_n28444_,
    new_n28445_, new_n28446_, new_n28447_, new_n28448_, new_n28449_,
    new_n28450_, new_n28451_, new_n28452_, new_n28453_, new_n28454_,
    new_n28455_, new_n28456_, new_n28457_, new_n28458_, new_n28459_,
    new_n28460_, new_n28461_, new_n28462_, new_n28463_, new_n28464_,
    new_n28465_, new_n28466_, new_n28467_, new_n28468_, new_n28469_,
    new_n28470_, new_n28471_, new_n28472_, new_n28473_, new_n28474_,
    new_n28475_, new_n28476_, new_n28477_, new_n28478_, new_n28479_,
    new_n28480_, new_n28481_, new_n28482_, new_n28483_, new_n28484_,
    new_n28485_, new_n28486_, new_n28487_, new_n28488_, new_n28489_,
    new_n28490_, new_n28491_, new_n28492_, new_n28493_, new_n28494_,
    new_n28495_, new_n28496_, new_n28497_, new_n28498_, new_n28499_,
    new_n28500_, new_n28501_, new_n28502_, new_n28503_, new_n28504_,
    new_n28505_, new_n28507_, new_n28508_, new_n28509_, new_n28510_,
    new_n28511_, new_n28512_, new_n28513_, new_n28514_, new_n28515_,
    new_n28516_, new_n28517_, new_n28518_, new_n28519_, new_n28520_,
    new_n28521_, new_n28522_, new_n28523_, new_n28524_, new_n28525_,
    new_n28526_, new_n28527_, new_n28528_, new_n28529_, new_n28530_,
    new_n28531_, new_n28532_, new_n28533_, new_n28534_, new_n28535_,
    new_n28536_, new_n28537_, new_n28538_, new_n28539_, new_n28540_,
    new_n28541_, new_n28542_, new_n28543_, new_n28544_, new_n28546_,
    new_n28547_, new_n28548_, new_n28549_, new_n28550_, new_n28551_,
    new_n28552_, new_n28553_, new_n28554_, new_n28555_, new_n28556_,
    new_n28557_, new_n28558_, new_n28559_, new_n28560_, new_n28561_,
    new_n28562_, new_n28563_, new_n28564_, new_n28565_, new_n28566_,
    new_n28567_, new_n28568_, new_n28569_, new_n28570_, new_n28572_,
    new_n28573_, new_n28574_, new_n28575_, new_n28576_, new_n28577_,
    new_n28578_, new_n28579_, new_n28580_, new_n28581_, new_n28582_,
    new_n28583_, new_n28584_, new_n28585_, new_n28586_, new_n28587_,
    new_n28588_, new_n28589_, new_n28590_, new_n28591_, new_n28592_,
    new_n28593_, new_n28594_, new_n28595_, new_n28596_, new_n28597_,
    new_n28598_, new_n28599_, new_n28600_, new_n28601_, new_n28602_,
    new_n28603_, new_n28604_, new_n28605_, new_n28606_, new_n28607_,
    new_n28608_, new_n28609_, new_n28610_, new_n28611_, new_n28612_,
    new_n28613_, new_n28614_, new_n28615_, new_n28617_, new_n28618_,
    new_n28619_, new_n28620_, new_n28621_, new_n28622_, new_n28623_,
    new_n28624_, new_n28625_, new_n28626_, new_n28627_, new_n28628_,
    new_n28629_, new_n28630_, new_n28631_, new_n28632_, new_n28633_,
    new_n28635_, new_n28636_, new_n28637_, new_n28638_, new_n28639_,
    new_n28640_, new_n28641_, new_n28642_, new_n28643_, new_n28644_,
    new_n28645_, new_n28646_, new_n28647_, new_n28648_, new_n28649_,
    new_n28650_, new_n28651_, new_n28652_, new_n28653_, new_n28654_,
    new_n28655_, new_n28656_, new_n28659_, new_n28660_, new_n28661_,
    new_n28662_, new_n28663_, new_n28664_, new_n28665_, new_n28666_,
    new_n28667_, new_n28668_, new_n28669_, new_n28670_, new_n28671_,
    new_n28672_, new_n28673_, new_n28674_, new_n28675_, new_n28676_,
    new_n28677_, new_n28678_, new_n28679_, new_n28680_, new_n28681_,
    new_n28682_, new_n28683_, new_n28684_, new_n28685_, new_n28686_,
    new_n28687_, new_n28688_, new_n28689_, new_n28690_, new_n28691_,
    new_n28692_, new_n28693_, new_n28694_, new_n28695_, new_n28696_,
    new_n28697_, new_n28699_, new_n28700_, new_n28701_, new_n28702_,
    new_n28703_, new_n28704_, new_n28705_, new_n28706_, new_n28707_,
    new_n28708_, new_n28709_, new_n28710_, new_n28711_, new_n28712_,
    new_n28713_, new_n28714_, new_n28715_, new_n28716_, new_n28717_,
    new_n28718_, new_n28719_, new_n28720_, new_n28721_, new_n28722_,
    new_n28723_, new_n28724_, new_n28725_, new_n28726_, new_n28727_,
    new_n28728_, new_n28729_, new_n28730_, new_n28731_, new_n28732_,
    new_n28733_, new_n28735_, new_n28736_, new_n28737_, new_n28738_,
    new_n28739_, new_n28740_, new_n28741_, new_n28742_, new_n28743_,
    new_n28744_, new_n28745_, new_n28746_, new_n28747_, new_n28748_,
    new_n28749_, new_n28750_, new_n28751_, new_n28752_, new_n28753_,
    new_n28754_, new_n28755_, new_n28756_, new_n28757_, new_n28758_,
    new_n28760_, new_n28761_, new_n28762_, new_n28763_, new_n28764_,
    new_n28765_, new_n28766_, new_n28767_, new_n28768_, new_n28769_,
    new_n28770_, new_n28771_, new_n28772_, new_n28773_, new_n28774_,
    new_n28775_, new_n28776_, new_n28777_, new_n28778_, new_n28779_,
    new_n28781_, new_n28782_, new_n28783_, new_n28784_, new_n28785_,
    new_n28786_, new_n28787_, new_n28788_, new_n28789_, new_n28790_,
    new_n28791_, new_n28792_, new_n28793_, new_n28794_, new_n28795_,
    new_n28796_, new_n28797_, new_n28798_, new_n28799_, new_n28800_,
    new_n28802_, new_n28803_, new_n28804_, new_n28805_, new_n28806_,
    new_n28807_, new_n28808_, new_n28809_, new_n28810_, new_n28811_,
    new_n28812_, new_n28813_, new_n28814_, new_n28815_, new_n28816_,
    new_n28817_, new_n28818_, new_n28819_, new_n28820_, new_n28821_,
    new_n28822_, new_n28823_, new_n28824_, new_n28825_, new_n28826_,
    new_n28827_, new_n28828_, new_n28829_, new_n28830_, new_n28831_,
    new_n28832_, new_n28833_, new_n28834_, new_n28836_, new_n28838_,
    new_n28839_, new_n28840_, new_n28841_, new_n28842_, new_n28843_,
    new_n28844_, new_n28845_, new_n28846_, new_n28847_, new_n28849_,
    new_n28850_, new_n28851_, new_n28852_, new_n28853_, new_n28854_,
    new_n28855_, new_n28856_, new_n28857_, new_n28858_, new_n28859_,
    new_n28860_, new_n28861_, new_n28862_, new_n28863_, new_n28866_,
    new_n28868_, new_n28870_, new_n28871_, new_n28872_, new_n28873_,
    new_n28874_, new_n28875_, new_n28876_, new_n28877_, new_n28878_,
    new_n28879_, new_n28880_, new_n28881_, new_n28882_, new_n28893_,
    new_n28894_, new_n28895_, new_n28896_, new_n28898_, new_n28899_,
    new_n28900_, new_n28901_, new_n28903_, new_n28904_, new_n28905_,
    new_n28906_, new_n28908_, new_n28909_, new_n28910_, new_n28911_,
    new_n28912_, new_n28913_, new_n28914_, new_n28915_, new_n28916_,
    new_n28917_, new_n28918_, new_n28919_, new_n28920_, new_n28921_,
    new_n28930_, new_n28931_, new_n28932_, new_n28933_, new_n28934_,
    new_n28935_, new_n28936_, new_n28937_, new_n28938_, new_n28939_,
    new_n28940_, new_n28941_, new_n28942_, new_n28943_, new_n28944_,
    new_n28946_, new_n28948_, new_n28950_, new_n28952_, new_n28954_,
    new_n28955_, new_n28956_, new_n28957_, new_n28958_, new_n28959_,
    new_n28960_, new_n28962_, new_n28965_, new_n28967_, new_n28980_,
    new_n28981_, new_n28982_, new_n28983_, new_n28984_, new_n28986_,
    new_n28988_, new_n28989_, new_n28990_, new_n28991_, new_n28992_,
    new_n28993_, new_n29002_, new_n29003_, new_n29004_, new_n29006_,
    new_n29080_, new_n29124_, new_n29125_, new_n29126_, new_n29127_,
    new_n29128_, new_n29129_, new_n29130_, new_n29131_, new_n29132_,
    new_n29133_, new_n29134_, new_n29135_, new_n29136_, new_n29137_,
    new_n29138_, new_n29139_, new_n29140_, new_n29141_, new_n29142_,
    new_n29151_, new_n29152_, new_n29153_, new_n29154_, new_n29155_,
    new_n29156_, new_n29157_, new_n29158_, new_n29159_, new_n29160_,
    new_n29161_, new_n29162_, new_n29163_, new_n29165_, new_n29166_,
    new_n29167_, new_n29168_, new_n29169_, new_n29170_, new_n29171_,
    new_n29172_, new_n29173_, new_n29174_, new_n29175_, new_n29177_,
    new_n29178_, new_n29179_, new_n29180_, new_n29181_, new_n29182_,
    new_n29183_, new_n29184_, new_n29185_, new_n29186_, new_n29187_,
    new_n29188_, new_n29189_, new_n29190_, new_n29191_, new_n29192_,
    new_n29194_, new_n29196_, new_n29197_, new_n29198_, new_n29199_,
    new_n29200_, new_n29201_, new_n29202_, new_n29203_, new_n29204_,
    new_n29206_, new_n29207_, new_n29208_, new_n29209_, new_n29210_,
    new_n29211_, new_n29212_, new_n29213_, new_n29214_, new_n29216_,
    new_n29217_, new_n29218_, new_n29219_, new_n29220_, new_n29221_,
    new_n29222_, new_n29223_, new_n29224_, new_n29226_, new_n29227_,
    new_n29228_, new_n29229_, new_n29230_, new_n29231_, new_n29232_,
    new_n29233_, new_n29234_, new_n29236_, new_n29237_, new_n29238_,
    new_n29239_, new_n29240_, new_n29242_, new_n29243_, new_n29244_,
    new_n29245_, new_n29246_, new_n29248_, new_n29249_, new_n29250_,
    new_n29251_, new_n29252_, new_n29254_, new_n29255_, new_n29256_,
    new_n29257_, new_n29258_, new_n29259_, new_n29269_, new_n29276_,
    new_n29280_, new_n29289_, new_n29290_, new_n29291_, new_n29292_,
    new_n29293_, new_n29300_, new_n29301_, new_n29302_, new_n29310_,
    new_n29311_, new_n29312_, new_n29313_, new_n29315_, new_n29320_,
    new_n29321_, new_n29322_, new_n29324_, new_n29335_, new_n29346_,
    new_n29347_, new_n29348_, new_n29355_, new_n29363_, new_n29364_,
    new_n29365_, new_n29376_, new_n29377_, new_n29378_, new_n29379_,
    new_n29380_, new_n29381_, new_n29382_, new_n29383_, new_n29384_,
    new_n29385_, new_n29386_, new_n29387_, new_n29388_, new_n29389_,
    new_n29390_, new_n29391_, new_n29392_, new_n29393_, new_n29394_,
    new_n29395_, new_n29396_, new_n29397_, new_n29398_, new_n29399_,
    new_n29400_, new_n29401_, new_n29402_, new_n29403_, new_n29404_,
    new_n29405_, new_n29406_, new_n29407_, new_n29408_, new_n29409_,
    new_n29410_, new_n29411_, new_n29412_, new_n29413_, new_n29414_,
    new_n29415_, new_n29416_, new_n29417_, new_n29418_, new_n29419_,
    new_n29420_, new_n29421_, new_n29422_, new_n29423_, new_n29424_,
    new_n29425_, new_n29426_, new_n29427_, new_n29428_, new_n29429_,
    new_n29430_, new_n29431_, new_n29432_, new_n29433_, new_n29434_,
    new_n29435_, new_n29436_, new_n29439_, new_n29441_, new_n29442_,
    new_n29443_, new_n29460_, new_n29461_, new_n29463_, new_n29464_,
    new_n29466_, new_n29467_, new_n29468_, new_n29469_, new_n29470_,
    new_n29471_, new_n29472_, new_n29473_, new_n29474_, new_n29475_,
    new_n29477_, new_n29478_, new_n29480_, new_n29482_, new_n29484_,
    new_n29485_, new_n29486_, new_n29487_, new_n29488_, new_n29489_,
    new_n29490_, new_n29491_, new_n29492_, new_n29493_, new_n29494_,
    new_n29495_, new_n29496_, new_n29497_, new_n29498_, new_n29499_,
    new_n29500_, new_n29501_, new_n29502_, new_n29503_, new_n29504_,
    new_n29505_, new_n29506_, new_n29507_, new_n29508_, new_n29509_,
    new_n29510_, new_n29511_, new_n29512_, new_n29513_, new_n29514_,
    new_n29515_, new_n29516_, new_n29517_, new_n29518_, new_n29519_,
    new_n29520_, new_n29521_, new_n29522_, new_n29523_, new_n29524_,
    new_n29525_, new_n29526_, new_n29527_, new_n29528_, new_n29529_,
    new_n29530_, new_n29531_, new_n29532_, new_n29533_, new_n29534_,
    new_n29535_, new_n29536_, new_n29537_, new_n29538_, new_n29539_,
    new_n29540_, new_n29541_, new_n29542_, new_n29543_, new_n29544_,
    new_n29545_, new_n29546_, new_n29547_, new_n29548_, new_n29549_,
    new_n29550_, new_n29551_, new_n29552_, new_n29553_, new_n29554_,
    new_n29555_, new_n29556_, new_n29557_, new_n29558_, new_n29559_,
    new_n29560_, new_n29561_, new_n29562_, new_n29563_, new_n29564_,
    new_n29565_, new_n29566_, new_n29567_, new_n29568_, new_n29569_,
    new_n29570_, new_n29571_, new_n29572_, new_n29573_, new_n29574_,
    new_n29575_, new_n29576_, new_n29577_, new_n29578_, new_n29579_,
    new_n29580_, new_n29581_, new_n29582_, new_n29583_, new_n29584_,
    new_n29585_, new_n29586_, new_n29587_, new_n29588_, new_n29589_,
    new_n29590_, new_n29591_, new_n29592_, new_n29593_, new_n29594_,
    new_n29595_, new_n29596_, new_n29597_, new_n29598_, new_n29599_,
    new_n29600_, new_n29601_, new_n29602_, new_n29603_, new_n29604_,
    new_n29605_, new_n29606_, new_n29607_, new_n29608_, new_n29609_,
    new_n29610_, new_n29611_, new_n29612_, new_n29613_, new_n29614_,
    new_n29615_, new_n29616_, new_n29617_, new_n29618_, new_n29619_,
    new_n29620_, new_n29621_, new_n29622_, new_n29623_, new_n29624_,
    new_n29625_, new_n29626_, new_n29627_, new_n29628_, new_n29629_,
    new_n29630_, new_n29631_, new_n29632_, new_n29633_, new_n29634_,
    new_n29635_, new_n29636_, new_n29637_, new_n29638_, new_n29639_,
    new_n29640_, new_n29641_, new_n29642_, new_n29643_, new_n29644_,
    new_n29645_, new_n29646_, new_n29647_, new_n29648_, new_n29649_,
    new_n29650_, new_n29651_, new_n29652_, new_n29653_, new_n29654_,
    new_n29655_, new_n29656_, new_n29657_, new_n29658_, new_n29659_,
    new_n29660_, new_n29661_, new_n29662_, new_n29663_, new_n29664_,
    new_n29665_, new_n29666_, new_n29667_, new_n29668_, new_n29669_,
    new_n29670_, new_n29671_, new_n29672_, new_n29673_, new_n29674_,
    new_n29675_, new_n29676_, new_n29677_, new_n29678_, new_n29679_,
    new_n29680_, new_n29681_, new_n29682_, new_n29683_, new_n29684_,
    new_n29685_, new_n29686_, new_n29687_, new_n29688_, new_n29689_,
    new_n29690_, new_n29691_, new_n29692_, new_n29693_, new_n29694_,
    new_n29695_, new_n29696_, new_n29697_, new_n29698_, new_n29699_,
    new_n29700_, new_n29701_, new_n29702_, new_n29703_, new_n29704_,
    new_n29705_, new_n29706_, new_n29707_, new_n29708_, new_n29709_,
    new_n29710_, new_n29711_, new_n29712_, new_n29713_, new_n29714_,
    new_n29715_, new_n29716_, new_n29717_, new_n29718_, new_n29719_,
    new_n29720_, new_n29721_, new_n29722_, new_n29723_, new_n29724_,
    new_n29725_, new_n29726_, new_n29727_, new_n29728_, new_n29729_,
    new_n29730_, new_n29731_, new_n29732_, new_n29733_, new_n29734_,
    new_n29735_, new_n29736_, new_n29737_, new_n29738_, new_n29739_,
    new_n29740_, new_n29741_, new_n29742_, new_n29743_, new_n29744_,
    new_n29745_, new_n29746_, new_n29747_, new_n29748_, new_n29749_,
    new_n29750_, new_n29751_, new_n29752_, new_n29753_, new_n29754_,
    new_n29755_, new_n29756_, new_n29757_, new_n29758_, new_n29759_,
    new_n29760_, new_n29761_, new_n29762_, new_n29763_, new_n29764_,
    new_n29765_, new_n29766_, new_n29767_, new_n29768_, new_n29769_,
    new_n29770_, new_n29771_, new_n29772_, new_n29773_, new_n29774_,
    new_n29775_, new_n29776_, new_n29777_, new_n29778_, new_n29779_,
    new_n29780_, new_n29781_, new_n29782_, new_n29783_, new_n29784_,
    new_n29785_, new_n29786_, new_n29787_, new_n29788_, new_n29789_,
    new_n29790_, new_n29791_, new_n29792_, new_n29793_, new_n29794_,
    new_n29795_, new_n29796_, new_n29797_, new_n29798_, new_n29799_,
    new_n29800_, new_n29801_, new_n29802_, new_n29803_, new_n29804_,
    new_n29805_, new_n29806_, new_n29807_, new_n29808_, new_n29809_,
    new_n29810_, new_n29811_, new_n29812_, new_n29813_, new_n29814_,
    new_n29815_, new_n29816_, new_n29817_, new_n29818_, new_n29819_,
    new_n29820_, new_n29821_, new_n29822_, new_n29823_, new_n29824_,
    new_n29825_, new_n29826_, new_n29827_, new_n29828_, new_n29829_,
    new_n29830_, new_n29831_, new_n29832_, new_n29833_, new_n29834_,
    new_n29835_, new_n29836_, new_n29837_, new_n29838_, new_n29839_,
    new_n29840_, new_n29841_, new_n29842_, new_n29843_, new_n29844_,
    new_n29845_, new_n29846_, new_n29847_, new_n29848_, new_n29849_,
    new_n29850_, new_n29851_, new_n29852_, new_n29853_, new_n29854_,
    new_n29855_, new_n29856_, new_n29857_, new_n29858_, new_n29859_,
    new_n29860_, new_n29861_, new_n29862_, new_n29863_, new_n29864_,
    new_n29865_, new_n29866_, new_n29867_, new_n29868_, new_n29869_,
    new_n29870_, new_n29871_, new_n29872_, new_n29873_, new_n29874_,
    new_n29875_, new_n29876_, new_n29877_, new_n29878_, new_n29879_,
    new_n29880_, new_n29881_, new_n29882_, new_n29883_, new_n29884_,
    new_n29885_, new_n29886_, new_n29887_, new_n29888_, new_n29889_,
    new_n29890_, new_n29891_, new_n29892_, new_n29893_, new_n29894_,
    new_n29895_, new_n29896_, new_n29897_, new_n29898_, new_n29899_,
    new_n29900_, new_n29901_, new_n29902_, new_n29903_, new_n29904_,
    new_n29905_, new_n29906_, new_n29907_, new_n29908_, new_n29909_,
    new_n29910_, new_n29911_, new_n29912_, new_n29913_, new_n29914_,
    new_n29915_, new_n29916_, new_n29917_, new_n29918_, new_n29919_,
    new_n29920_, new_n29921_, new_n29922_, new_n29923_, new_n29924_,
    new_n29925_, new_n29926_, new_n29927_, new_n29928_, new_n29929_,
    new_n29930_, new_n29931_, new_n29932_, new_n29933_, new_n29934_,
    new_n29935_, new_n29936_, new_n29937_, new_n29938_, new_n29939_,
    new_n29940_, new_n29941_, new_n29942_, new_n29943_, new_n29944_,
    new_n29945_, new_n29946_, new_n29947_, new_n29948_, new_n29949_,
    new_n29950_, new_n29951_, new_n29952_, new_n29953_, new_n29954_,
    new_n29955_, new_n29956_, new_n29957_, new_n29958_, new_n29959_,
    new_n29960_, new_n29961_, new_n29962_, new_n29963_, new_n29964_,
    new_n29965_, new_n29966_, new_n29967_, new_n29968_, new_n29969_,
    new_n29970_, new_n29971_, new_n29972_, new_n29973_, new_n29974_,
    new_n29975_, new_n29976_, new_n29977_, new_n29978_, new_n29979_,
    new_n29980_, new_n29981_, new_n29982_, new_n29983_, new_n29984_,
    new_n29985_, new_n29986_, new_n29987_, new_n29988_, new_n29989_,
    new_n29990_, new_n29991_, new_n29992_, new_n29993_, new_n29994_,
    new_n29995_, new_n29996_, new_n29997_, new_n29998_, new_n29999_,
    new_n30000_, new_n30001_, new_n30003_, new_n30004_, new_n30005_,
    new_n30006_, new_n30008_, new_n30009_, new_n30010_, new_n30011_,
    new_n30013_, new_n30014_, new_n30015_, new_n30017_, new_n30018_,
    new_n30019_, new_n30021_, new_n30022_, new_n30023_, new_n30025_,
    new_n30026_, new_n30028_, new_n30029_, new_n30030_, new_n30032_,
    new_n30033_, new_n30035_, new_n30036_, new_n30037_, new_n30038_,
    new_n30040_, new_n30041_, new_n30042_, new_n30044_, new_n30045_,
    new_n30046_, new_n30047_, new_n30048_, new_n30050_, new_n30051_,
    new_n30052_, new_n30054_, new_n30055_, new_n30057_, new_n30059_,
    new_n30060_, new_n30061_, new_n30063_, new_n30065_, new_n30067_,
    new_n30068_, new_n30070_, new_n30071_, new_n30073_, new_n30075_,
    new_n30076_, new_n30078_, new_n30079_, new_n30080_, new_n30082_,
    new_n30083_, new_n30085_, new_n30086_, new_n30087_, new_n30089_,
    new_n30091_, new_n30093_, new_n30095_, new_n30096_, new_n30098_,
    new_n30100_, new_n30102_, new_n30104_, new_n30105_, new_n30106_,
    new_n30108_, new_n30109_, new_n30111_, new_n30112_, new_n30113_,
    new_n30115_, new_n30117_, new_n30119_, new_n30121_, new_n30123_,
    new_n30125_, new_n30126_, new_n30127_, new_n30129_, new_n30130_,
    new_n30131_, new_n30133_, new_n30135_, new_n30137_, new_n30138_,
    new_n30139_, new_n30141_, new_n30142_, new_n30143_, new_n30145_,
    new_n30147_, new_n30149_, new_n30151_, new_n30152_, new_n30153_,
    new_n30155_, new_n30157_, new_n30159_, new_n30161_, new_n30163_,
    new_n30164_, new_n30165_, new_n30167_, new_n30168_, new_n30169_,
    new_n30171_, new_n30173_, new_n30175_, new_n30176_, new_n30177_,
    new_n30179_, new_n30180_, new_n30182_, new_n30183_, new_n30184_,
    new_n30186_, new_n30187_, new_n30188_, new_n30190_, new_n30191_,
    new_n30192_, new_n30194_, new_n30195_, new_n30197_, new_n30198_,
    new_n30199_, new_n30201_, new_n30202_, new_n30204_, new_n30205_,
    new_n30207_, new_n30208_, new_n30210_, new_n30211_, new_n30212_,
    new_n30213_, new_n30214_, new_n30215_, new_n30216_, new_n30218_,
    new_n30220_, new_n30222_, new_n30224_, new_n30225_, new_n30226_,
    new_n30227_, new_n30228_, new_n30229_, new_n30230_, new_n30231_,
    new_n30232_, new_n30233_, new_n30234_, new_n30235_, new_n30236_,
    new_n30237_, new_n30238_, new_n30239_, new_n30240_, new_n30241_,
    new_n30242_, new_n30243_, new_n30244_, new_n30245_, new_n30246_,
    new_n30247_, new_n30248_, new_n30249_, new_n30250_, new_n30251_,
    new_n30252_, new_n30253_, new_n30254_, new_n30256_, new_n30257_,
    new_n30258_, new_n30259_, new_n30260_, new_n30261_, new_n30262_,
    new_n30263_, new_n30264_, new_n30265_, new_n30266_, new_n30267_,
    new_n30268_, new_n30269_, new_n30270_, new_n30271_, new_n30272_,
    new_n30273_, new_n30274_, new_n30275_, new_n30276_, new_n30277_,
    new_n30278_, new_n30279_, new_n30280_, new_n30281_, new_n30282_,
    new_n30284_, new_n30286_, new_n30287_, new_n30288_, new_n30289_,
    new_n30290_, new_n30291_, new_n30292_, new_n30293_, new_n30294_,
    new_n30295_, new_n30296_, new_n30297_, new_n30298_, new_n30299_,
    new_n30300_, new_n30301_, new_n30302_, new_n30304_, new_n30305_,
    new_n30306_, new_n30307_, new_n30308_, new_n30309_, new_n30310_,
    new_n30311_, new_n30312_, new_n30313_, new_n30314_, new_n30315_,
    new_n30316_, new_n30317_, new_n30318_, new_n30319_, new_n30320_,
    new_n30321_, new_n30323_, new_n30324_, new_n30325_, new_n30326_,
    new_n30327_, new_n30328_, new_n30329_, new_n30330_, new_n30331_,
    new_n30332_, new_n30333_, new_n30334_, new_n30335_, new_n30336_,
    new_n30337_, new_n30338_, new_n30339_, new_n30340_, new_n30341_,
    new_n30343_, new_n30344_, new_n30346_, new_n30347_, new_n30348_,
    new_n30349_, new_n30350_, new_n30351_, new_n30352_, new_n30353_,
    new_n30354_, new_n30355_, new_n30356_, new_n30357_, new_n30358_,
    new_n30359_, new_n30360_, new_n30361_, new_n30362_, new_n30363_,
    new_n30365_, new_n30366_, new_n30367_, new_n30368_, new_n30369_,
    new_n30370_, new_n30371_, new_n30372_, new_n30373_, new_n30374_,
    new_n30375_, new_n30376_, new_n30377_, new_n30378_, new_n30379_,
    new_n30380_, new_n30381_, new_n30383_, new_n30384_, new_n30385_,
    new_n30386_, new_n30387_, new_n30388_, new_n30389_, new_n30390_,
    new_n30391_, new_n30392_, new_n30393_, new_n30394_, new_n30395_,
    new_n30396_, new_n30397_, new_n30398_, new_n30399_, new_n30400_,
    new_n30401_, new_n30403_, new_n30404_, new_n30405_, new_n30406_,
    new_n30407_, new_n30408_, new_n30409_, new_n30410_, new_n30411_,
    new_n30412_, new_n30413_, new_n30414_, new_n30415_, new_n30416_,
    new_n30417_, new_n30418_, new_n30419_, new_n30421_, new_n30422_,
    new_n30423_, new_n30424_, new_n30425_, new_n30426_, new_n30427_,
    new_n30428_, new_n30429_, new_n30430_, new_n30431_, new_n30432_,
    new_n30433_, new_n30434_, new_n30435_, new_n30436_, new_n30437_,
    new_n30438_, new_n30439_, new_n30440_, new_n30442_, new_n30443_,
    new_n30444_, new_n30445_, new_n30446_, new_n30447_, new_n30448_,
    new_n30449_, new_n30450_, new_n30451_, new_n30452_, new_n30453_,
    new_n30454_, new_n30455_, new_n30456_, new_n30457_, new_n30458_,
    new_n30459_, new_n30460_, new_n30462_, new_n30463_, new_n30464_,
    new_n30465_, new_n30466_, new_n30467_, new_n30468_, new_n30469_,
    new_n30470_, new_n30471_, new_n30472_, new_n30473_, new_n30474_,
    new_n30475_, new_n30476_, new_n30477_, new_n30478_, new_n30479_,
    new_n30481_, new_n30482_, new_n30483_, new_n30484_, new_n30485_,
    new_n30486_, new_n30487_, new_n30488_, new_n30489_, new_n30490_,
    new_n30491_, new_n30492_, new_n30493_, new_n30494_, new_n30495_,
    new_n30496_, new_n30497_, new_n30499_, new_n30500_, new_n30501_,
    new_n30502_, new_n30503_, new_n30504_, new_n30505_, new_n30506_,
    new_n30507_, new_n30508_, new_n30509_, new_n30510_, new_n30511_,
    new_n30512_, new_n30513_, new_n30514_, new_n30515_, new_n30517_,
    new_n30518_, new_n30519_, new_n30520_, new_n30521_, new_n30522_,
    new_n30523_, new_n30524_, new_n30525_, new_n30526_, new_n30527_,
    new_n30528_, new_n30529_, new_n30530_, new_n30531_, new_n30532_,
    new_n30533_, new_n30534_, new_n30535_, new_n30537_, new_n30539_,
    new_n30541_, new_n30542_, new_n30543_, new_n30544_, new_n30545_,
    new_n30546_, new_n30547_, new_n30548_, new_n30549_, new_n30550_,
    new_n30551_, new_n30552_, new_n30553_, new_n30554_, new_n30555_,
    new_n30556_, new_n30557_, new_n30559_, new_n30561_, new_n30562_,
    new_n30564_, new_n30565_, new_n30566_, new_n30567_, new_n30568_,
    new_n30569_, new_n30570_, new_n30571_, new_n30572_, new_n30573_,
    new_n30574_, new_n30575_, new_n30576_, new_n30577_, new_n30578_,
    new_n30579_, new_n30580_, new_n30581_, new_n30582_, new_n30583_,
    new_n30585_, new_n30587_, new_n30588_, new_n30590_, new_n30592_,
    new_n30593_, new_n30594_, new_n30595_, new_n30596_, new_n30597_,
    new_n30598_, new_n30599_, new_n30600_, new_n30601_, new_n30602_,
    new_n30603_, new_n30604_, new_n30605_, new_n30606_, new_n30608_,
    new_n30610_, new_n30612_, new_n30613_, new_n30614_, new_n30615_,
    new_n30616_, new_n30617_, new_n30618_, new_n30619_, new_n30620_,
    new_n30621_, new_n30622_, new_n30623_, new_n30624_, new_n30625_,
    new_n30626_, new_n30627_, new_n30628_, new_n30629_, new_n30630_,
    new_n30631_, new_n30632_, new_n30633_, new_n30635_, new_n30636_,
    new_n30638_, new_n30639_, new_n30641_, new_n30642_, new_n30644_,
    new_n30646_, new_n30647_, new_n30649_, new_n30650_, new_n30652_,
    new_n30654_, new_n30656_, new_n30657_, new_n30659_, new_n30660_,
    new_n30662_, new_n30664_, new_n30666_, new_n30668_, new_n30670_,
    new_n30671_, new_n30672_, new_n30673_, new_n30674_, new_n30675_,
    new_n30676_, new_n30677_, new_n30678_, new_n30679_, new_n30680_,
    new_n30681_, new_n30682_, new_n30683_, new_n30684_, new_n30685_,
    new_n30686_, new_n30687_, new_n30688_, new_n30689_, new_n30690_,
    new_n30692_, new_n30693_, new_n30694_, new_n30695_, new_n30696_,
    new_n30697_, new_n30698_, new_n30699_, new_n30700_, new_n30701_,
    new_n30702_, new_n30703_, new_n30704_, new_n30705_, new_n30706_,
    new_n30707_, new_n30708_, new_n30709_, new_n30710_, new_n30711_,
    new_n30712_, new_n30713_, new_n30715_, new_n30716_, new_n30718_,
    new_n30720_, new_n30721_, new_n30722_, new_n30723_, new_n30724_,
    new_n30725_, new_n30726_, new_n30727_, new_n30728_, new_n30729_,
    new_n30730_, new_n30731_, new_n30732_, new_n30733_, new_n30734_,
    new_n30735_, new_n30736_, new_n30738_, new_n30739_, new_n30740_,
    new_n30741_, new_n30742_, new_n30743_, new_n30744_, new_n30745_,
    new_n30746_, new_n30747_, new_n30748_, new_n30749_, new_n30750_,
    new_n30751_, new_n30752_, new_n30753_, new_n30754_, new_n30755_,
    new_n30756_, new_n30758_, new_n30759_, new_n30760_, new_n30761_,
    new_n30762_, new_n30763_, new_n30764_, new_n30765_, new_n30766_,
    new_n30767_, new_n30768_, new_n30769_, new_n30770_, new_n30771_,
    new_n30772_, new_n30773_, new_n30774_, new_n30776_, new_n30777_,
    new_n30778_, new_n30779_, new_n30780_, new_n30781_, new_n30782_,
    new_n30783_, new_n30784_, new_n30785_, new_n30786_, new_n30787_,
    new_n30788_, new_n30789_, new_n30790_, new_n30792_, new_n30794_,
    new_n30795_, new_n30796_, new_n30797_, new_n30798_, new_n30799_,
    new_n30800_, new_n30801_, new_n30802_, new_n30803_, new_n30804_,
    new_n30805_, new_n30806_, new_n30807_, new_n30808_, new_n30809_,
    new_n30810_, new_n30811_, new_n30812_, new_n30814_, new_n30815_,
    new_n30816_, new_n30817_, new_n30818_, new_n30819_, new_n30820_,
    new_n30821_, new_n30822_, new_n30823_, new_n30824_, new_n30825_,
    new_n30826_, new_n30827_, new_n30828_, new_n30829_, new_n30830_,
    new_n30831_, new_n30833_, new_n30834_, new_n30835_, new_n30836_,
    new_n30837_, new_n30838_, new_n30839_, new_n30840_, new_n30841_,
    new_n30842_, new_n30843_, new_n30844_, new_n30845_, new_n30846_,
    new_n30847_, new_n30848_, new_n30849_, new_n30850_, new_n30851_,
    new_n30853_, new_n30854_, new_n30855_, new_n30856_, new_n30857_,
    new_n30858_, new_n30859_, new_n30860_, new_n30861_, new_n30862_,
    new_n30863_, new_n30864_, new_n30865_, new_n30866_, new_n30867_,
    new_n30868_, new_n30869_, new_n30870_, new_n30872_, new_n30873_,
    new_n30874_, new_n30875_, new_n30876_, new_n30877_, new_n30878_,
    new_n30879_, new_n30880_, new_n30881_, new_n30882_, new_n30883_,
    new_n30884_, new_n30885_, new_n30886_, new_n30887_, new_n30889_,
    new_n30890_, new_n30891_, new_n30892_, new_n30893_, new_n30894_,
    new_n30895_, new_n30896_, new_n30897_, new_n30898_, new_n30899_,
    new_n30900_, new_n30901_, new_n30902_, new_n30903_, new_n30904_,
    new_n30905_, new_n30906_, new_n30907_, new_n30908_, new_n30909_,
    new_n30910_, new_n30911_, new_n30912_, new_n30913_, new_n30914_,
    new_n30915_, new_n30916_, new_n30917_, new_n30918_, new_n30919_,
    new_n30920_, new_n30921_, new_n30922_, new_n30923_, new_n30924_,
    new_n30925_, new_n30927_, new_n30928_, new_n30929_, new_n30930_,
    new_n30931_, new_n30932_, new_n30933_, new_n30934_, new_n30935_,
    new_n30936_, new_n30937_, new_n30938_, new_n30939_, new_n30940_,
    new_n30941_, new_n30942_, new_n30943_, new_n30944_, new_n30945_,
    new_n30947_, new_n30949_, new_n30951_, new_n30952_, new_n30954_,
    new_n30956_, new_n30958_, new_n30959_, new_n30961_, new_n30963_,
    new_n30965_, new_n30966_, new_n30967_, new_n30968_, new_n30969_,
    new_n30970_, new_n30971_, new_n30972_, new_n30973_, new_n30974_,
    new_n30975_, new_n30976_, new_n30977_, new_n30979_, new_n30981_,
    new_n30982_, new_n30983_, new_n30984_, new_n30985_, new_n30986_,
    new_n30987_, new_n30988_, new_n30989_, new_n30990_, new_n30991_,
    new_n30992_, new_n30993_, new_n30994_, new_n30995_, new_n30996_,
    new_n30997_, new_n30998_, new_n30999_, new_n31001_, new_n31002_,
    new_n31004_, new_n31006_, new_n31008_, new_n31009_, new_n31011_,
    new_n31012_, new_n31015_, new_n31016_, new_n31018_, new_n31020_,
    new_n31022_, new_n31023_, new_n31025_, new_n31027_, new_n31029_,
    new_n31030_, new_n31032_, new_n31033_, new_n31034_, new_n31035_,
    new_n31036_, new_n31037_, new_n31038_, new_n31039_, new_n31040_,
    new_n31042_, new_n31043_, new_n31045_, new_n31046_, new_n31048_,
    new_n31050_, new_n31052_, new_n31054_, new_n31056_, new_n31058_,
    new_n31060_, new_n31062_, new_n31064_, new_n31065_, new_n31067_,
    new_n31068_, new_n31070_, new_n31072_, new_n31074_, new_n31076_,
    new_n31077_, new_n31078_, new_n31080_, new_n31081_, new_n31083_,
    new_n31085_, new_n31086_, new_n31087_, new_n31088_, new_n31089_,
    new_n31090_, new_n31091_, new_n31092_, new_n31093_, new_n31094_,
    new_n31095_, new_n31096_, new_n31097_, new_n31098_, new_n31099_,
    new_n31100_, new_n31101_, new_n31102_, new_n31103_, new_n31105_,
    new_n31106_, new_n31108_, new_n31110_, new_n31112_, new_n31113_,
    new_n31114_, new_n31115_, new_n31116_, new_n31117_, new_n31118_,
    new_n31119_, new_n31120_, new_n31121_, new_n31122_, new_n31124_,
    new_n31126_, new_n31127_, new_n31128_, new_n31129_, new_n31130_,
    new_n31131_, new_n31133_, new_n31134_, new_n31136_, new_n31137_,
    new_n31139_, new_n31140_, new_n31141_, new_n31142_, new_n31144_,
    new_n31146_, new_n31147_, new_n31148_, new_n31149_, new_n31150_,
    new_n31151_, new_n31152_, new_n31153_, new_n31154_, new_n31156_,
    new_n31158_, new_n31160_, new_n31161_, new_n31162_, new_n31167_,
    new_n31179_, new_n31180_, new_n31183_, new_n31184_, new_n31185_,
    new_n31188_, new_n31192_, new_n31194_, new_n31197_, new_n31201_,
    new_n31205_, new_n31208_, new_n31215_, new_n31218_, new_n31220_,
    new_n31221_, new_n31222_, new_n31223_, new_n31224_, new_n31225_,
    new_n31226_, new_n31227_, new_n31228_, new_n31229_, new_n31230_,
    new_n31231_, new_n31233_, new_n31234_, new_n31236_, new_n31237_,
    new_n31238_, new_n31239_, new_n31240_, new_n31241_, new_n31242_,
    new_n31243_, new_n31244_, new_n31245_, new_n31247_, new_n31248_,
    new_n31250_, new_n31251_, new_n31252_, new_n31253_, new_n31254_,
    new_n31255_, new_n31256_, new_n31257_, new_n31258_, new_n31259_,
    new_n31261_, new_n31262_, new_n31264_, new_n31265_, new_n31266_,
    new_n31267_, new_n31268_, new_n31269_, new_n31270_, new_n31271_,
    new_n31272_, new_n31273_, new_n31275_, new_n31276_, new_n31278_,
    new_n31309_, new_n31310_, new_n31311_, new_n31320_, new_n31321_,
    new_n31322_, new_n31329_, new_n31330_, new_n31331_, new_n31334_,
    new_n31335_, new_n31336_, new_n31338_, new_n31339_, new_n31340_,
    new_n31342_, new_n31343_, new_n31344_, new_n31390_, new_n31391_,
    new_n31392_, new_n31393_, new_n31394_, new_n31395_, new_n31396_,
    new_n31425_, new_n31450_;
  INVX1    g00000(.A(pi0057), .Y(new_n2436_));
  INVX1    g00001(.A(pi0221), .Y(new_n2437_));
  INVX1    g00002(.A(pi0216), .Y(new_n2438_));
  INVX1    g00003(.A(pi1144), .Y(new_n2439_));
  AOI21X1  g00004(.A0(pi0833), .A1(new_n2438_), .B0(new_n2439_), .Y(new_n2440_));
  AND3X1   g00005(.A(pi0929), .B(pi0833), .C(new_n2438_), .Y(new_n2441_));
  NOR3X1   g00006(.A(new_n2441_), .B(new_n2440_), .C(pi0332), .Y(new_n2442_));
  NOR2X1   g00007(.A(new_n2442_), .B(new_n2437_), .Y(new_n2443_));
  INVX1    g00008(.A(pi0332), .Y(new_n2444_));
  AOI21X1  g00009(.A0(new_n2444_), .A1(pi0265), .B0(new_n2438_), .Y(new_n2445_));
  INVX1    g00010(.A(new_n2445_), .Y(new_n2446_));
  INVX1    g00011(.A(pi0105), .Y(new_n2447_));
  AND2X1   g00012(.A(new_n2444_), .B(pi0153), .Y(new_n2448_));
  INVX1    g00013(.A(new_n2448_), .Y(new_n2449_));
  NOR3X1   g00014(.A(pi0166), .B(pi0161), .C(pi0152), .Y(new_n2450_));
  INVX1    g00015(.A(new_n2450_), .Y(new_n2451_));
  INVX1    g00016(.A(pi0137), .Y(new_n2452_));
  INVX1    g00017(.A(pi0479), .Y(new_n2453_));
  AND2X1   g00018(.A(new_n2453_), .B(pi0095), .Y(new_n2454_));
  INVX1    g00019(.A(pi0032), .Y(new_n2455_));
  NOR2X1   g00020(.A(pi0072), .B(pi0040), .Y(new_n2456_));
  OR4X1    g00021(.A(pi0098), .B(pi0088), .C(pi0077), .D(pi0050), .Y(new_n2457_));
  OR2X1    g00022(.A(new_n2457_), .B(pi0102), .Y(new_n2458_));
  OR2X1    g00023(.A(pi0071), .B(pi0065), .Y(new_n2459_));
  OR2X1    g00024(.A(pi0103), .B(pi0083), .Y(new_n2460_));
  OR2X1    g00025(.A(pi0069), .B(pi0067), .Y(new_n2461_));
  OR2X1    g00026(.A(pi0073), .B(pi0066), .Y(new_n2462_));
  OR4X1    g00027(.A(pi0106), .B(pi0085), .C(pi0076), .D(pi0061), .Y(new_n2463_));
  OR4X1    g00028(.A(new_n2463_), .B(pi0089), .C(pi0049), .D(pi0048), .Y(new_n2464_));
  OR3X1    g00029(.A(pi0111), .B(pi0082), .C(pi0036), .Y(new_n2465_));
  OR3X1    g00030(.A(new_n2465_), .B(pi0084), .C(pi0068), .Y(new_n2466_));
  OR4X1    g00031(.A(new_n2466_), .B(new_n2464_), .C(pi0104), .D(pi0045), .Y(new_n2467_));
  OR4X1    g00032(.A(new_n2467_), .B(new_n2462_), .C(new_n2461_), .D(new_n2460_), .Y(new_n2468_));
  OR2X1    g00033(.A(pi0107), .B(pi0063), .Y(new_n2469_));
  OR4X1    g00034(.A(new_n2469_), .B(new_n2468_), .C(new_n2459_), .D(pi0064), .Y(new_n2470_));
  OR2X1    g00035(.A(new_n2470_), .B(pi0081), .Y(new_n2471_));
  OR3X1    g00036(.A(pi0086), .B(pi0060), .C(pi0053), .Y(new_n2472_));
  OR2X1    g00037(.A(pi0108), .B(pi0097), .Y(new_n2473_));
  OR4X1    g00038(.A(new_n2473_), .B(new_n2472_), .C(pi0094), .D(pi0046), .Y(new_n2474_));
  OR3X1    g00039(.A(pi0091), .B(pi0058), .C(pi0047), .Y(new_n2475_));
  OR3X1    g00040(.A(new_n2475_), .B(pi0110), .C(pi0109), .Y(new_n2476_));
  NOR4X1   g00041(.A(new_n2476_), .B(new_n2474_), .C(new_n2471_), .D(new_n2458_), .Y(new_n2477_));
  OR4X1    g00042(.A(pi0096), .B(pi0070), .C(pi0051), .D(pi0035), .Y(new_n2478_));
  NOR3X1   g00043(.A(new_n2478_), .B(pi0093), .C(pi0090), .Y(new_n2479_));
  AND3X1   g00044(.A(new_n2479_), .B(new_n2477_), .C(new_n2456_), .Y(new_n2480_));
  AOI21X1  g00045(.A0(new_n2480_), .A1(pi0225), .B0(new_n2455_), .Y(new_n2481_));
  NOR2X1   g00046(.A(new_n2481_), .B(pi0095), .Y(new_n2482_));
  NOR2X1   g00047(.A(pi0093), .B(pi0090), .Y(new_n2483_));
  INVX1    g00048(.A(new_n2483_), .Y(new_n2484_));
  INVX1    g00049(.A(pi0053), .Y(new_n2485_));
  INVX1    g00050(.A(pi0060), .Y(new_n2486_));
  OR4X1    g00051(.A(new_n2470_), .B(new_n2458_), .C(pi0081), .D(new_n2486_), .Y(new_n2487_));
  AND2X1   g00052(.A(new_n2487_), .B(new_n2485_), .Y(new_n2488_));
  NOR2X1   g00053(.A(pi0094), .B(pi0086), .Y(new_n2489_));
  INVX1    g00054(.A(new_n2489_), .Y(new_n2490_));
  OR4X1    g00055(.A(new_n2470_), .B(new_n2458_), .C(pi0081), .D(pi0060), .Y(new_n2491_));
  AOI21X1  g00056(.A0(new_n2491_), .A1(pi0053), .B0(new_n2490_), .Y(new_n2492_));
  INVX1    g00057(.A(new_n2492_), .Y(new_n2493_));
  INVX1    g00058(.A(pi0058), .Y(new_n2494_));
  OR3X1    g00059(.A(pi0110), .B(pi0109), .C(pi0046), .Y(new_n2495_));
  NOR4X1   g00060(.A(new_n2495_), .B(new_n2473_), .C(pi0091), .D(pi0047), .Y(new_n2496_));
  AND2X1   g00061(.A(new_n2496_), .B(new_n2494_), .Y(new_n2497_));
  INVX1    g00062(.A(new_n2497_), .Y(new_n2498_));
  NOR4X1   g00063(.A(new_n2498_), .B(new_n2493_), .C(new_n2488_), .D(new_n2484_), .Y(new_n2499_));
  OR2X1    g00064(.A(new_n2499_), .B(pi0035), .Y(new_n2500_));
  NOR2X1   g00065(.A(pi0090), .B(pi0058), .Y(new_n2501_));
  INVX1    g00066(.A(new_n2501_), .Y(new_n2502_));
  OR3X1    g00067(.A(new_n2474_), .B(pi0110), .C(pi0109), .Y(new_n2503_));
  OR3X1    g00068(.A(new_n2503_), .B(pi0091), .C(pi0047), .Y(new_n2504_));
  OR4X1    g00069(.A(new_n2504_), .B(new_n2470_), .C(new_n2458_), .D(pi0081), .Y(new_n2505_));
  OR3X1    g00070(.A(new_n2505_), .B(new_n2502_), .C(pi0093), .Y(new_n2506_));
  AND2X1   g00071(.A(new_n2506_), .B(pi0035), .Y(new_n2507_));
  INVX1    g00072(.A(pi0035), .Y(new_n2508_));
  OR4X1    g00073(.A(new_n2505_), .B(new_n2502_), .C(pi0093), .D(new_n2508_), .Y(new_n2509_));
  NOR2X1   g00074(.A(new_n2509_), .B(pi0225), .Y(new_n2510_));
  NOR4X1   g00075(.A(new_n2510_), .B(new_n2507_), .C(pi0070), .D(pi0051), .Y(new_n2511_));
  AOI21X1  g00076(.A0(new_n2511_), .A1(new_n2500_), .B0(pi0096), .Y(new_n2512_));
  INVX1    g00077(.A(pi0096), .Y(new_n2513_));
  OR4X1    g00078(.A(new_n2474_), .B(pi0110), .C(pi0109), .D(pi0047), .Y(new_n2514_));
  INVX1    g00079(.A(pi0091), .Y(new_n2515_));
  INVX1    g00080(.A(pi0093), .Y(new_n2516_));
  NOR3X1   g00081(.A(pi0070), .B(pi0051), .C(pi0035), .Y(new_n2517_));
  NAND4X1  g00082(.A(new_n2517_), .B(new_n2501_), .C(new_n2516_), .D(new_n2515_), .Y(new_n2518_));
  NOR4X1   g00083(.A(new_n2518_), .B(new_n2514_), .C(new_n2471_), .D(new_n2458_), .Y(new_n2519_));
  OAI21X1  g00084(.A0(new_n2519_), .A1(new_n2513_), .B0(new_n2456_), .Y(new_n2520_));
  OAI21X1  g00085(.A0(new_n2520_), .A1(new_n2512_), .B0(new_n2455_), .Y(new_n2521_));
  AOI21X1  g00086(.A0(new_n2521_), .A1(new_n2482_), .B0(new_n2454_), .Y(new_n2522_));
  INVX1    g00087(.A(pi0095), .Y(new_n2523_));
  NOR2X1   g00088(.A(pi0093), .B(pi0035), .Y(new_n2524_));
  INVX1    g00089(.A(new_n2524_), .Y(new_n2525_));
  OR4X1    g00090(.A(pi0096), .B(pi0072), .C(pi0070), .D(pi0051), .Y(new_n2526_));
  NOR4X1   g00091(.A(new_n2526_), .B(new_n2525_), .C(new_n2505_), .D(new_n2502_), .Y(new_n2527_));
  AOI21X1  g00092(.A0(new_n2527_), .A1(pi0040), .B0(pi0032), .Y(new_n2528_));
  INVX1    g00093(.A(pi0040), .Y(new_n2529_));
  INVX1    g00094(.A(pi0072), .Y(new_n2530_));
  AND2X1   g00095(.A(new_n2479_), .B(new_n2477_), .Y(new_n2531_));
  OR2X1    g00096(.A(new_n2531_), .B(new_n2530_), .Y(new_n2532_));
  AND2X1   g00097(.A(new_n2532_), .B(new_n2529_), .Y(new_n2533_));
  INVX1    g00098(.A(pi0051), .Y(new_n2534_));
  INVX1    g00099(.A(pi0070), .Y(new_n2535_));
  OR4X1    g00100(.A(new_n2525_), .B(new_n2505_), .C(new_n2502_), .D(pi0070), .Y(new_n2536_));
  AOI21X1  g00101(.A0(new_n2536_), .A1(pi0051), .B0(pi0096), .Y(new_n2537_));
  OAI21X1  g00102(.A0(new_n2535_), .A1(pi0051), .B0(new_n2537_), .Y(new_n2538_));
  INVX1    g00103(.A(pi0225), .Y(new_n2539_));
  OAI21X1  g00104(.A0(new_n2506_), .A1(new_n2539_), .B0(pi0035), .Y(new_n2540_));
  OR3X1    g00105(.A(new_n2505_), .B(new_n2502_), .C(new_n2516_), .Y(new_n2541_));
  AND2X1   g00106(.A(new_n2541_), .B(new_n2508_), .Y(new_n2542_));
  INVX1    g00107(.A(new_n2542_), .Y(new_n2543_));
  NOR4X1   g00108(.A(new_n2514_), .B(new_n2470_), .C(new_n2458_), .D(pi0081), .Y(new_n2544_));
  AOI21X1  g00109(.A0(new_n2544_), .A1(pi0091), .B0(new_n2502_), .Y(new_n2545_));
  INVX1    g00110(.A(pi0109), .Y(new_n2546_));
  INVX1    g00111(.A(pi0110), .Y(new_n2547_));
  NOR4X1   g00112(.A(new_n2474_), .B(new_n2470_), .C(new_n2458_), .D(pi0081), .Y(new_n2548_));
  AOI21X1  g00113(.A0(new_n2548_), .A1(new_n2546_), .B0(new_n2547_), .Y(new_n2549_));
  INVX1    g00114(.A(pi0047), .Y(new_n2550_));
  NOR3X1   g00115(.A(new_n2470_), .B(new_n2458_), .C(pi0081), .Y(new_n2551_));
  INVX1    g00116(.A(new_n2503_), .Y(new_n2552_));
  AOI21X1  g00117(.A0(new_n2552_), .A1(new_n2551_), .B0(new_n2550_), .Y(new_n2553_));
  NOR3X1   g00118(.A(new_n2553_), .B(new_n2549_), .C(pi0091), .Y(new_n2554_));
  NOR2X1   g00119(.A(pi0110), .B(pi0047), .Y(new_n2555_));
  INVX1    g00120(.A(new_n2555_), .Y(new_n2556_));
  NOR2X1   g00121(.A(new_n2548_), .B(new_n2546_), .Y(new_n2557_));
  OR2X1    g00122(.A(pi0098), .B(pi0088), .Y(new_n2558_));
  OR4X1    g00123(.A(new_n2470_), .B(new_n2558_), .C(pi0102), .D(pi0081), .Y(new_n2559_));
  NOR4X1   g00124(.A(pi0077), .B(pi0060), .C(pi0053), .D(pi0050), .Y(new_n2560_));
  NAND2X1  g00125(.A(new_n2560_), .B(new_n2489_), .Y(new_n2561_));
  OR3X1    g00126(.A(new_n2561_), .B(new_n2559_), .C(pi0097), .Y(new_n2562_));
  AOI21X1  g00127(.A0(new_n2562_), .A1(pi0108), .B0(pi0046), .Y(new_n2563_));
  OR2X1    g00128(.A(new_n2561_), .B(new_n2559_), .Y(new_n2564_));
  AND2X1   g00129(.A(new_n2564_), .B(pi0097), .Y(new_n2565_));
  INVX1    g00130(.A(pi0086), .Y(new_n2566_));
  OR3X1    g00131(.A(new_n2470_), .B(pi0102), .C(pi0081), .Y(new_n2567_));
  OR3X1    g00132(.A(pi0060), .B(pi0053), .C(pi0050), .Y(new_n2568_));
  NOR4X1   g00133(.A(new_n2568_), .B(new_n2567_), .C(new_n2558_), .D(pi0077), .Y(new_n2569_));
  AND3X1   g00134(.A(new_n2569_), .B(pi0094), .C(new_n2566_), .Y(new_n2570_));
  NOR2X1   g00135(.A(new_n2570_), .B(pi0097), .Y(new_n2571_));
  INVX1    g00136(.A(pi0094), .Y(new_n2572_));
  OAI21X1  g00137(.A0(new_n2569_), .A1(new_n2566_), .B0(new_n2572_), .Y(new_n2573_));
  INVX1    g00138(.A(new_n2573_), .Y(new_n2574_));
  AND2X1   g00139(.A(new_n2491_), .B(pi0053), .Y(new_n2575_));
  INVX1    g00140(.A(pi0077), .Y(new_n2576_));
  NOR2X1   g00141(.A(new_n2559_), .B(new_n2576_), .Y(new_n2577_));
  NOR2X1   g00142(.A(new_n2577_), .B(pi0050), .Y(new_n2578_));
  INVX1    g00143(.A(pi0081), .Y(new_n2579_));
  INVX1    g00144(.A(pi0102), .Y(new_n2580_));
  NOR4X1   g00145(.A(new_n2469_), .B(new_n2468_), .C(new_n2459_), .D(pi0064), .Y(new_n2581_));
  AOI21X1  g00146(.A0(new_n2581_), .A1(new_n2579_), .B0(new_n2580_), .Y(new_n2582_));
  AOI21X1  g00147(.A0(new_n2470_), .A1(pi0081), .B0(new_n2582_), .Y(new_n2583_));
  INVX1    g00148(.A(pi0064), .Y(new_n2584_));
  NOR3X1   g00149(.A(new_n2469_), .B(new_n2468_), .C(new_n2459_), .Y(new_n2585_));
  NOR2X1   g00150(.A(new_n2585_), .B(new_n2584_), .Y(new_n2586_));
  INVX1    g00151(.A(pi0107), .Y(new_n2587_));
  AND2X1   g00152(.A(new_n2468_), .B(pi0071), .Y(new_n2588_));
  OR2X1    g00153(.A(new_n2588_), .B(pi0065), .Y(new_n2589_));
  INVX1    g00154(.A(pi0071), .Y(new_n2590_));
  INVX1    g00155(.A(pi0069), .Y(new_n2591_));
  NOR3X1   g00156(.A(new_n2467_), .B(new_n2462_), .C(pi0067), .Y(new_n2592_));
  NOR2X1   g00157(.A(new_n2592_), .B(new_n2591_), .Y(new_n2593_));
  INVX1    g00158(.A(pi0083), .Y(new_n2594_));
  INVX1    g00159(.A(pi0103), .Y(new_n2595_));
  NOR3X1   g00160(.A(new_n2467_), .B(new_n2462_), .C(new_n2461_), .Y(new_n2596_));
  OAI21X1  g00161(.A0(new_n2596_), .A1(new_n2594_), .B0(new_n2595_), .Y(new_n2597_));
  NOR2X1   g00162(.A(new_n2597_), .B(new_n2593_), .Y(new_n2598_));
  NOR2X1   g00163(.A(pi0083), .B(pi0069), .Y(new_n2599_));
  INVX1    g00164(.A(new_n2599_), .Y(new_n2600_));
  NOR2X1   g00165(.A(pi0111), .B(pi0068), .Y(new_n2601_));
  INVX1    g00166(.A(new_n2601_), .Y(new_n2602_));
  INVX1    g00167(.A(pi0084), .Y(new_n2603_));
  OR4X1    g00168(.A(new_n2464_), .B(new_n2462_), .C(pi0104), .D(pi0045), .Y(new_n2604_));
  AND2X1   g00169(.A(new_n2604_), .B(pi0084), .Y(new_n2605_));
  NOR3X1   g00170(.A(new_n2464_), .B(pi0104), .C(pi0045), .Y(new_n2606_));
  NOR2X1   g00171(.A(new_n2464_), .B(pi0104), .Y(new_n2607_));
  OR3X1    g00172(.A(new_n2463_), .B(pi0089), .C(pi0048), .Y(new_n2608_));
  INVX1    g00173(.A(pi0048), .Y(new_n2609_));
  INVX1    g00174(.A(new_n2463_), .Y(new_n2610_));
  OR2X1    g00175(.A(pi0076), .B(pi0061), .Y(new_n2611_));
  OR2X1    g00176(.A(pi0106), .B(pi0085), .Y(new_n2612_));
  AND2X1   g00177(.A(pi0106), .B(pi0085), .Y(new_n2613_));
  AND2X1   g00178(.A(pi0076), .B(pi0061), .Y(new_n2614_));
  OAI22X1  g00179(.A0(new_n2614_), .A1(new_n2612_), .B0(new_n2613_), .B1(new_n2611_), .Y(new_n2615_));
  AOI21X1  g00180(.A0(new_n2615_), .A1(new_n2609_), .B0(new_n2610_), .Y(new_n2616_));
  INVX1    g00181(.A(pi0049), .Y(new_n2617_));
  OAI21X1  g00182(.A0(new_n2463_), .A1(pi0048), .B0(pi0089), .Y(new_n2618_));
  NAND2X1  g00183(.A(new_n2618_), .B(new_n2617_), .Y(new_n2619_));
  OAI21X1  g00184(.A0(new_n2619_), .A1(new_n2616_), .B0(new_n2608_), .Y(new_n2620_));
  AOI21X1  g00185(.A0(new_n2464_), .A1(pi0104), .B0(pi0045), .Y(new_n2621_));
  AOI21X1  g00186(.A0(new_n2621_), .A1(new_n2620_), .B0(new_n2607_), .Y(new_n2622_));
  NOR2X1   g00187(.A(new_n2622_), .B(new_n2606_), .Y(new_n2623_));
  INVX1    g00188(.A(new_n2606_), .Y(new_n2624_));
  AND2X1   g00189(.A(pi0073), .B(pi0066), .Y(new_n2625_));
  AOI21X1  g00190(.A0(new_n2624_), .A1(new_n2462_), .B0(new_n2625_), .Y(new_n2626_));
  OAI21X1  g00191(.A0(new_n2623_), .A1(new_n2462_), .B0(new_n2626_), .Y(new_n2627_));
  AOI21X1  g00192(.A0(new_n2627_), .A1(new_n2603_), .B0(new_n2605_), .Y(new_n2628_));
  INVX1    g00193(.A(pi0082), .Y(new_n2629_));
  INVX1    g00194(.A(pi0111), .Y(new_n2630_));
  NOR3X1   g00195(.A(new_n2604_), .B(pi0084), .C(pi0068), .Y(new_n2631_));
  OAI21X1  g00196(.A0(new_n2631_), .A1(new_n2630_), .B0(new_n2629_), .Y(new_n2632_));
  OR2X1    g00197(.A(new_n2604_), .B(pi0084), .Y(new_n2633_));
  AND2X1   g00198(.A(new_n2633_), .B(pi0068), .Y(new_n2634_));
  NOR2X1   g00199(.A(new_n2634_), .B(new_n2632_), .Y(new_n2635_));
  OAI21X1  g00200(.A0(new_n2628_), .A1(new_n2602_), .B0(new_n2635_), .Y(new_n2636_));
  OR2X1    g00201(.A(pi0067), .B(pi0036), .Y(new_n2637_));
  NOR4X1   g00202(.A(new_n2604_), .B(new_n2602_), .C(pi0084), .D(new_n2629_), .Y(new_n2638_));
  NOR2X1   g00203(.A(new_n2638_), .B(new_n2637_), .Y(new_n2639_));
  INVX1    g00204(.A(pi0036), .Y(new_n2640_));
  OAI21X1  g00205(.A0(new_n2467_), .A1(new_n2462_), .B0(pi0067), .Y(new_n2641_));
  OR2X1    g00206(.A(pi0111), .B(pi0082), .Y(new_n2642_));
  NOR4X1   g00207(.A(new_n2604_), .B(new_n2642_), .C(pi0084), .D(pi0068), .Y(new_n2643_));
  OAI21X1  g00208(.A0(new_n2643_), .A1(new_n2640_), .B0(new_n2641_), .Y(new_n2644_));
  AOI21X1  g00209(.A0(new_n2639_), .A1(new_n2636_), .B0(new_n2644_), .Y(new_n2645_));
  OAI21X1  g00210(.A0(new_n2645_), .A1(new_n2600_), .B0(new_n2598_), .Y(new_n2646_));
  NAND3X1  g00211(.A(new_n2599_), .B(new_n2592_), .C(pi0103), .Y(new_n2647_));
  AND3X1   g00212(.A(new_n2647_), .B(new_n2646_), .C(new_n2590_), .Y(new_n2648_));
  OAI21X1  g00213(.A0(new_n2648_), .A1(new_n2589_), .B0(new_n2587_), .Y(new_n2649_));
  INVX1    g00214(.A(pi0065), .Y(new_n2650_));
  NOR3X1   g00215(.A(new_n2468_), .B(pi0071), .C(new_n2650_), .Y(new_n2651_));
  OR2X1    g00216(.A(new_n2468_), .B(new_n2459_), .Y(new_n2652_));
  AOI21X1  g00217(.A0(new_n2652_), .A1(pi0107), .B0(pi0063), .Y(new_n2653_));
  OAI21X1  g00218(.A0(new_n2651_), .A1(new_n2649_), .B0(new_n2653_), .Y(new_n2654_));
  AOI21X1  g00219(.A0(new_n2654_), .A1(new_n2584_), .B0(new_n2586_), .Y(new_n2655_));
  INVX1    g00220(.A(pi0063), .Y(new_n2656_));
  OR2X1    g00221(.A(pi0107), .B(new_n2656_), .Y(new_n2657_));
  OAI21X1  g00222(.A0(new_n2657_), .A1(new_n2652_), .B0(new_n2584_), .Y(new_n2658_));
  AOI21X1  g00223(.A0(new_n2653_), .A1(new_n2649_), .B0(new_n2658_), .Y(new_n2659_));
  NOR2X1   g00224(.A(new_n2659_), .B(new_n2586_), .Y(new_n2660_));
  OR4X1    g00225(.A(new_n2660_), .B(new_n2655_), .C(pi0102), .D(pi0081), .Y(new_n2661_));
  AOI21X1  g00226(.A0(new_n2661_), .A1(new_n2583_), .B0(new_n2558_), .Y(new_n2662_));
  INVX1    g00227(.A(pi0088), .Y(new_n2663_));
  NOR4X1   g00228(.A(new_n2470_), .B(pi0102), .C(pi0098), .D(pi0081), .Y(new_n2664_));
  AOI21X1  g00229(.A0(new_n2567_), .A1(pi0098), .B0(pi0077), .Y(new_n2665_));
  OAI21X1  g00230(.A0(new_n2664_), .A1(new_n2663_), .B0(new_n2665_), .Y(new_n2666_));
  OAI21X1  g00231(.A0(new_n2666_), .A1(new_n2662_), .B0(new_n2578_), .Y(new_n2667_));
  NOR3X1   g00232(.A(new_n2567_), .B(new_n2558_), .C(pi0077), .Y(new_n2668_));
  INVX1    g00233(.A(new_n2668_), .Y(new_n2669_));
  AOI21X1  g00234(.A0(new_n2669_), .A1(pi0050), .B0(pi0060), .Y(new_n2670_));
  NAND2X1  g00235(.A(new_n2670_), .B(new_n2667_), .Y(new_n2671_));
  AOI21X1  g00236(.A0(new_n2671_), .A1(new_n2488_), .B0(new_n2575_), .Y(new_n2672_));
  OAI21X1  g00237(.A0(new_n2672_), .A1(pi0086), .B0(new_n2574_), .Y(new_n2673_));
  AOI21X1  g00238(.A0(new_n2673_), .A1(new_n2571_), .B0(new_n2565_), .Y(new_n2674_));
  OAI21X1  g00239(.A0(new_n2674_), .A1(pi0108), .B0(new_n2563_), .Y(new_n2675_));
  INVX1    g00240(.A(pi0046), .Y(new_n2676_));
  NOR4X1   g00241(.A(new_n2561_), .B(new_n2559_), .C(new_n2473_), .D(new_n2676_), .Y(new_n2677_));
  NOR2X1   g00242(.A(new_n2677_), .B(pi0109), .Y(new_n2678_));
  AOI21X1  g00243(.A0(new_n2678_), .A1(new_n2675_), .B0(new_n2557_), .Y(new_n2679_));
  OAI21X1  g00244(.A0(new_n2679_), .A1(new_n2556_), .B0(new_n2554_), .Y(new_n2680_));
  AND2X1   g00245(.A(new_n2505_), .B(pi0058), .Y(new_n2681_));
  INVX1    g00246(.A(pi0090), .Y(new_n2682_));
  NOR2X1   g00247(.A(new_n2477_), .B(new_n2682_), .Y(new_n2683_));
  OR3X1    g00248(.A(new_n2683_), .B(new_n2681_), .C(pi0093), .Y(new_n2684_));
  AOI21X1  g00249(.A0(new_n2680_), .A1(new_n2545_), .B0(new_n2684_), .Y(new_n2685_));
  OAI21X1  g00250(.A0(new_n2685_), .A1(new_n2543_), .B0(new_n2540_), .Y(new_n2686_));
  AOI21X1  g00251(.A0(new_n2686_), .A1(new_n2534_), .B0(new_n2538_), .Y(new_n2687_));
  OAI21X1  g00252(.A0(new_n2687_), .A1(pi0072), .B0(new_n2533_), .Y(new_n2688_));
  OR3X1    g00253(.A(new_n2525_), .B(new_n2505_), .C(new_n2502_), .Y(new_n2689_));
  NAND2X1  g00254(.A(new_n2519_), .B(pi0096), .Y(new_n2690_));
  OR2X1    g00255(.A(pi0072), .B(pi0051), .Y(new_n2691_));
  OR4X1    g00256(.A(new_n2691_), .B(new_n2690_), .C(new_n2689_), .D(pi0040), .Y(new_n2692_));
  AND3X1   g00257(.A(new_n2692_), .B(new_n2688_), .C(new_n2528_), .Y(new_n2693_));
  OAI21X1  g00258(.A0(new_n2693_), .A1(new_n2481_), .B0(new_n2523_), .Y(new_n2694_));
  NOR2X1   g00259(.A(pi0040), .B(pi0032), .Y(new_n2695_));
  AOI21X1  g00260(.A0(new_n2695_), .A1(new_n2527_), .B0(new_n2523_), .Y(new_n2696_));
  AND2X1   g00261(.A(new_n2696_), .B(pi0479), .Y(new_n2697_));
  INVX1    g00262(.A(new_n2697_), .Y(new_n2698_));
  AOI21X1  g00263(.A0(new_n2698_), .A1(new_n2694_), .B0(new_n2452_), .Y(new_n2699_));
  AOI21X1  g00264(.A0(new_n2522_), .A1(new_n2452_), .B0(new_n2699_), .Y(new_n2700_));
  INVX1    g00265(.A(pi0833), .Y(new_n2701_));
  INVX1    g00266(.A(pi1091), .Y(new_n2702_));
  AOI21X1  g00267(.A0(pi0957), .A1(new_n2701_), .B0(new_n2702_), .Y(new_n2703_));
  INVX1    g00268(.A(new_n2703_), .Y(new_n2704_));
  INVX1    g00269(.A(pi0841), .Y(new_n2705_));
  NOR4X1   g00270(.A(new_n2505_), .B(new_n2502_), .C(new_n2705_), .D(pi0093), .Y(new_n2706_));
  OR2X1    g00271(.A(pi0096), .B(pi0070), .Y(new_n2707_));
  NOR4X1   g00272(.A(new_n2707_), .B(new_n2539_), .C(pi0040), .D(pi0035), .Y(new_n2708_));
  NAND4X1  g00273(.A(new_n2708_), .B(new_n2706_), .C(new_n2530_), .D(new_n2534_), .Y(new_n2709_));
  AND2X1   g00274(.A(new_n2709_), .B(pi0032), .Y(new_n2710_));
  OAI21X1  g00275(.A0(new_n2710_), .A1(new_n2693_), .B0(new_n2523_), .Y(new_n2711_));
  AOI21X1  g00276(.A0(new_n2711_), .A1(new_n2698_), .B0(new_n2452_), .Y(new_n2712_));
  AND2X1   g00277(.A(pi0479), .B(pi0095), .Y(new_n2713_));
  INVX1    g00278(.A(new_n2710_), .Y(new_n2714_));
  AOI21X1  g00279(.A0(new_n2714_), .A1(new_n2521_), .B0(pi0095), .Y(new_n2715_));
  NOR2X1   g00280(.A(new_n2715_), .B(new_n2713_), .Y(new_n2716_));
  NOR2X1   g00281(.A(new_n2716_), .B(pi0137), .Y(new_n2717_));
  NOR2X1   g00282(.A(new_n2717_), .B(new_n2712_), .Y(new_n2718_));
  AND2X1   g00283(.A(pi0950), .B(pi0829), .Y(new_n2719_));
  AND2X1   g00284(.A(pi1093), .B(pi1092), .Y(new_n2720_));
  AND2X1   g00285(.A(new_n2720_), .B(new_n2719_), .Y(new_n2721_));
  NOR3X1   g00286(.A(new_n2721_), .B(new_n2715_), .C(new_n2713_), .Y(new_n2722_));
  INVX1    g00287(.A(new_n2722_), .Y(new_n2723_));
  INVX1    g00288(.A(new_n2719_), .Y(new_n2724_));
  INVX1    g00289(.A(new_n2720_), .Y(new_n2725_));
  INVX1    g00290(.A(new_n2511_), .Y(new_n2726_));
  NOR3X1   g00291(.A(new_n2565_), .B(pi0110), .C(pi0108), .Y(new_n2727_));
  OR3X1    g00292(.A(pi0093), .B(pi0090), .C(pi0058), .Y(new_n2728_));
  INVX1    g00293(.A(new_n2488_), .Y(new_n2729_));
  AOI21X1  g00294(.A0(new_n2492_), .A1(new_n2729_), .B0(pi0097), .Y(new_n2730_));
  NOR4X1   g00295(.A(pi0109), .B(pi0091), .C(pi0047), .D(pi0046), .Y(new_n2731_));
  INVX1    g00296(.A(new_n2731_), .Y(new_n2732_));
  NOR3X1   g00297(.A(new_n2732_), .B(new_n2730_), .C(new_n2728_), .Y(new_n2733_));
  AOI21X1  g00298(.A0(new_n2733_), .A1(new_n2727_), .B0(pi0035), .Y(new_n2734_));
  OR2X1    g00299(.A(new_n2734_), .B(new_n2726_), .Y(new_n2735_));
  AND2X1   g00300(.A(new_n2735_), .B(new_n2513_), .Y(new_n2736_));
  OAI21X1  g00301(.A0(new_n2736_), .A1(new_n2520_), .B0(new_n2455_), .Y(new_n2737_));
  AOI21X1  g00302(.A0(new_n2737_), .A1(new_n2714_), .B0(pi0095), .Y(new_n2738_));
  OR4X1    g00303(.A(new_n2738_), .B(new_n2725_), .C(new_n2724_), .D(new_n2713_), .Y(new_n2739_));
  AND3X1   g00304(.A(new_n2739_), .B(new_n2723_), .C(new_n2452_), .Y(new_n2740_));
  NOR3X1   g00305(.A(new_n2740_), .B(new_n2712_), .C(new_n2704_), .Y(new_n2741_));
  AOI21X1  g00306(.A0(new_n2718_), .A1(new_n2704_), .B0(new_n2741_), .Y(new_n2742_));
  INVX1    g00307(.A(new_n2742_), .Y(new_n2743_));
  MX2X1    g00308(.A(new_n2743_), .B(new_n2700_), .S0(pi0210), .Y(new_n2744_));
  NOR2X1   g00309(.A(new_n2499_), .B(pi0035), .Y(new_n2745_));
  NOR3X1   g00310(.A(pi0096), .B(pi0072), .C(pi0040), .Y(new_n2746_));
  INVX1    g00311(.A(new_n2746_), .Y(new_n2747_));
  NOR3X1   g00312(.A(new_n2747_), .B(new_n2726_), .C(new_n2745_), .Y(new_n2748_));
  OAI21X1  g00313(.A0(new_n2748_), .A1(pi0032), .B0(new_n2482_), .Y(new_n2749_));
  AND2X1   g00314(.A(new_n2749_), .B(new_n2452_), .Y(new_n2750_));
  NOR2X1   g00315(.A(new_n2696_), .B(new_n2454_), .Y(new_n2751_));
  AND2X1   g00316(.A(new_n2688_), .B(new_n2528_), .Y(new_n2752_));
  OAI21X1  g00317(.A0(new_n2752_), .A1(new_n2481_), .B0(new_n2523_), .Y(new_n2753_));
  AOI21X1  g00318(.A0(new_n2753_), .A1(new_n2751_), .B0(new_n2452_), .Y(new_n2754_));
  OAI21X1  g00319(.A0(new_n2754_), .A1(new_n2750_), .B0(pi0210), .Y(new_n2755_));
  OR2X1    g00320(.A(new_n2710_), .B(pi0095), .Y(new_n2756_));
  AND2X1   g00321(.A(new_n2721_), .B(new_n2703_), .Y(new_n2757_));
  INVX1    g00322(.A(pi0957), .Y(new_n2758_));
  AND2X1   g00323(.A(pi1093), .B(pi1091), .Y(new_n2759_));
  OAI21X1  g00324(.A0(new_n2758_), .A1(pi0833), .B0(new_n2759_), .Y(new_n2760_));
  AND3X1   g00325(.A(pi1092), .B(pi0950), .C(pi0829), .Y(new_n2761_));
  INVX1    g00326(.A(new_n2761_), .Y(new_n2762_));
  OR2X1    g00327(.A(new_n2762_), .B(new_n2760_), .Y(new_n2763_));
  OAI22X1  g00328(.A0(new_n2763_), .A1(new_n2734_), .B0(new_n2757_), .B1(new_n2745_), .Y(new_n2764_));
  AND2X1   g00329(.A(new_n2746_), .B(new_n2511_), .Y(new_n2765_));
  AOI21X1  g00330(.A0(new_n2765_), .A1(new_n2764_), .B0(pi0032), .Y(new_n2766_));
  OR2X1    g00331(.A(new_n2766_), .B(new_n2756_), .Y(new_n2767_));
  OAI21X1  g00332(.A0(new_n2710_), .A1(new_n2752_), .B0(new_n2523_), .Y(new_n2768_));
  AOI21X1  g00333(.A0(new_n2768_), .A1(new_n2751_), .B0(new_n2452_), .Y(new_n2769_));
  AOI21X1  g00334(.A0(new_n2767_), .A1(new_n2452_), .B0(new_n2769_), .Y(new_n2770_));
  OAI21X1  g00335(.A0(new_n2770_), .A1(pi0210), .B0(new_n2755_), .Y(new_n2771_));
  OAI21X1  g00336(.A0(new_n2771_), .A1(pi0234), .B0(new_n2444_), .Y(new_n2772_));
  AOI21X1  g00337(.A0(new_n2744_), .A1(pi0234), .B0(new_n2772_), .Y(new_n2773_));
  AND2X1   g00338(.A(new_n2444_), .B(pi0234), .Y(new_n2774_));
  NOR2X1   g00339(.A(new_n2718_), .B(pi0210), .Y(new_n2775_));
  INVX1    g00340(.A(pi0146), .Y(new_n2776_));
  INVX1    g00341(.A(pi0210), .Y(new_n2777_));
  OAI21X1  g00342(.A0(new_n2700_), .A1(new_n2777_), .B0(new_n2776_), .Y(new_n2778_));
  OAI21X1  g00343(.A0(new_n2778_), .A1(new_n2775_), .B0(new_n2774_), .Y(new_n2779_));
  AOI21X1  g00344(.A0(new_n2744_), .A1(pi0146), .B0(new_n2779_), .Y(new_n2780_));
  NOR2X1   g00345(.A(new_n2771_), .B(new_n2776_), .Y(new_n2781_));
  NOR2X1   g00346(.A(new_n2748_), .B(pi0032), .Y(new_n2782_));
  NOR2X1   g00347(.A(new_n2756_), .B(new_n2782_), .Y(new_n2783_));
  NOR2X1   g00348(.A(new_n2783_), .B(pi0137), .Y(new_n2784_));
  OR2X1    g00349(.A(new_n2784_), .B(new_n2769_), .Y(new_n2785_));
  AND2X1   g00350(.A(new_n2785_), .B(new_n2777_), .Y(new_n2786_));
  NAND2X1  g00351(.A(new_n2755_), .B(new_n2776_), .Y(new_n2787_));
  NOR2X1   g00352(.A(pi0332), .B(pi0234), .Y(new_n2788_));
  OAI21X1  g00353(.A0(new_n2787_), .A1(new_n2786_), .B0(new_n2788_), .Y(new_n2789_));
  OAI21X1  g00354(.A0(new_n2789_), .A1(new_n2781_), .B0(new_n2451_), .Y(new_n2790_));
  OAI22X1  g00355(.A0(new_n2790_), .A1(new_n2780_), .B0(new_n2773_), .B1(new_n2451_), .Y(new_n2791_));
  MX2X1    g00356(.A(new_n2791_), .B(new_n2449_), .S0(new_n2447_), .Y(new_n2792_));
  INVX1    g00357(.A(pi0228), .Y(new_n2793_));
  INVX1    g00358(.A(new_n2696_), .Y(new_n2794_));
  INVX1    g00359(.A(new_n2528_), .Y(new_n2795_));
  AOI21X1  g00360(.A0(new_n2675_), .A1(new_n2546_), .B0(new_n2557_), .Y(new_n2796_));
  OAI21X1  g00361(.A0(new_n2796_), .A1(new_n2556_), .B0(new_n2554_), .Y(new_n2797_));
  AOI21X1  g00362(.A0(new_n2797_), .A1(new_n2545_), .B0(new_n2684_), .Y(new_n2798_));
  OR2X1    g00363(.A(new_n2798_), .B(new_n2543_), .Y(new_n2799_));
  AOI21X1  g00364(.A0(new_n2799_), .A1(new_n2540_), .B0(pi0051), .Y(new_n2800_));
  OAI21X1  g00365(.A0(new_n2800_), .A1(new_n2538_), .B0(new_n2530_), .Y(new_n2801_));
  AOI21X1  g00366(.A0(new_n2801_), .A1(new_n2533_), .B0(new_n2795_), .Y(new_n2802_));
  AND2X1   g00367(.A(new_n2802_), .B(new_n2692_), .Y(new_n2803_));
  OAI21X1  g00368(.A0(new_n2803_), .A1(new_n2710_), .B0(new_n2523_), .Y(new_n2804_));
  AOI21X1  g00369(.A0(new_n2804_), .A1(new_n2794_), .B0(new_n2452_), .Y(new_n2805_));
  OAI21X1  g00370(.A0(new_n2450_), .A1(pi0146), .B0(new_n2703_), .Y(new_n2806_));
  NOR3X1   g00371(.A(new_n2715_), .B(new_n2713_), .C(new_n2696_), .Y(new_n2807_));
  OAI21X1  g00372(.A0(new_n2806_), .A1(new_n2722_), .B0(new_n2807_), .Y(new_n2808_));
  OR3X1    g00373(.A(new_n2806_), .B(new_n2739_), .C(new_n2696_), .Y(new_n2809_));
  AND3X1   g00374(.A(new_n2809_), .B(new_n2808_), .C(new_n2452_), .Y(new_n2810_));
  OAI21X1  g00375(.A0(new_n2810_), .A1(new_n2805_), .B0(new_n2777_), .Y(new_n2811_));
  OAI21X1  g00376(.A0(new_n2802_), .A1(new_n2710_), .B0(new_n2523_), .Y(new_n2812_));
  AOI21X1  g00377(.A0(new_n2812_), .A1(new_n2751_), .B0(new_n2452_), .Y(new_n2813_));
  OAI21X1  g00378(.A0(new_n2766_), .A1(new_n2756_), .B0(new_n2452_), .Y(new_n2814_));
  NOR2X1   g00379(.A(new_n2450_), .B(pi0146), .Y(new_n2815_));
  OR2X1    g00380(.A(pi0234), .B(pi0210), .Y(new_n2816_));
  AOI21X1  g00381(.A0(new_n2815_), .A1(new_n2784_), .B0(new_n2816_), .Y(new_n2817_));
  OAI21X1  g00382(.A0(new_n2815_), .A1(new_n2814_), .B0(new_n2817_), .Y(new_n2818_));
  OAI21X1  g00383(.A0(new_n2802_), .A1(new_n2481_), .B0(new_n2523_), .Y(new_n2819_));
  AOI21X1  g00384(.A0(new_n2819_), .A1(new_n2751_), .B0(new_n2452_), .Y(new_n2820_));
  OR2X1    g00385(.A(new_n2750_), .B(new_n2777_), .Y(new_n2821_));
  OAI22X1  g00386(.A0(new_n2821_), .A1(new_n2820_), .B0(new_n2818_), .B1(new_n2813_), .Y(new_n2822_));
  AOI21X1  g00387(.A0(new_n2811_), .A1(pi0234), .B0(new_n2822_), .Y(new_n2823_));
  OAI21X1  g00388(.A0(new_n2803_), .A1(new_n2481_), .B0(new_n2523_), .Y(new_n2824_));
  NOR2X1   g00389(.A(new_n2696_), .B(new_n2452_), .Y(new_n2825_));
  OR2X1    g00390(.A(new_n2696_), .B(pi0137), .Y(new_n2826_));
  AND2X1   g00391(.A(pi0234), .B(pi0210), .Y(new_n2827_));
  OAI21X1  g00392(.A0(new_n2826_), .A1(new_n2522_), .B0(new_n2827_), .Y(new_n2828_));
  AOI21X1  g00393(.A0(new_n2825_), .A1(new_n2824_), .B0(new_n2828_), .Y(new_n2829_));
  OAI21X1  g00394(.A0(new_n2829_), .A1(new_n2823_), .B0(new_n2448_), .Y(new_n2830_));
  INVX1    g00395(.A(new_n2757_), .Y(new_n2831_));
  NOR3X1   g00396(.A(new_n2510_), .B(pi0070), .C(pi0051), .Y(new_n2832_));
  OR2X1    g00397(.A(new_n2505_), .B(new_n2502_), .Y(new_n2833_));
  AOI21X1  g00398(.A0(new_n2833_), .A1(pi0093), .B0(pi0035), .Y(new_n2834_));
  NOR2X1   g00399(.A(new_n2683_), .B(new_n2681_), .Y(new_n2835_));
  INVX1    g00400(.A(new_n2835_), .Y(new_n2836_));
  INVX1    g00401(.A(pi0108), .Y(new_n2837_));
  INVX1    g00402(.A(new_n2571_), .Y(new_n2838_));
  OAI21X1  g00403(.A0(new_n2671_), .A1(pi0053), .B0(new_n2566_), .Y(new_n2839_));
  AOI21X1  g00404(.A0(new_n2839_), .A1(new_n2574_), .B0(new_n2838_), .Y(new_n2840_));
  OAI21X1  g00405(.A0(new_n2840_), .A1(new_n2565_), .B0(new_n2837_), .Y(new_n2841_));
  AOI21X1  g00406(.A0(new_n2841_), .A1(new_n2563_), .B0(pi0109), .Y(new_n2842_));
  NOR2X1   g00407(.A(new_n2842_), .B(new_n2557_), .Y(new_n2843_));
  OAI21X1  g00408(.A0(new_n2843_), .A1(new_n2556_), .B0(new_n2554_), .Y(new_n2844_));
  AOI21X1  g00409(.A0(new_n2844_), .A1(new_n2545_), .B0(new_n2836_), .Y(new_n2845_));
  OAI21X1  g00410(.A0(new_n2845_), .A1(pi0093), .B0(new_n2834_), .Y(new_n2846_));
  AND2X1   g00411(.A(new_n2536_), .B(pi0051), .Y(new_n2847_));
  AND2X1   g00412(.A(new_n2689_), .B(pi0070), .Y(new_n2848_));
  NOR3X1   g00413(.A(new_n2848_), .B(new_n2847_), .C(pi0096), .Y(new_n2849_));
  INVX1    g00414(.A(new_n2849_), .Y(new_n2850_));
  AOI21X1  g00415(.A0(new_n2846_), .A1(new_n2832_), .B0(new_n2850_), .Y(new_n2851_));
  AOI21X1  g00416(.A0(new_n2519_), .A1(pi0096), .B0(pi0072), .Y(new_n2852_));
  INVX1    g00417(.A(new_n2852_), .Y(new_n2853_));
  OR2X1    g00418(.A(new_n2853_), .B(new_n2851_), .Y(new_n2854_));
  AOI21X1  g00419(.A0(new_n2854_), .A1(new_n2533_), .B0(new_n2795_), .Y(new_n2855_));
  NAND2X1  g00420(.A(new_n2855_), .B(new_n2831_), .Y(new_n2856_));
  INVX1    g00421(.A(new_n2480_), .Y(new_n2857_));
  AND2X1   g00422(.A(pi0841), .B(pi0225), .Y(new_n2858_));
  OAI21X1  g00423(.A0(new_n2858_), .A1(new_n2857_), .B0(pi0032), .Y(new_n2859_));
  INVX1    g00424(.A(new_n2859_), .Y(new_n2860_));
  AND2X1   g00425(.A(new_n2757_), .B(new_n2528_), .Y(new_n2861_));
  OAI21X1  g00426(.A0(new_n2840_), .A1(pi0097), .B0(new_n2837_), .Y(new_n2862_));
  AOI21X1  g00427(.A0(new_n2862_), .A1(new_n2563_), .B0(pi0109), .Y(new_n2863_));
  NOR2X1   g00428(.A(new_n2863_), .B(new_n2557_), .Y(new_n2864_));
  OAI21X1  g00429(.A0(new_n2864_), .A1(new_n2556_), .B0(new_n2554_), .Y(new_n2865_));
  AOI21X1  g00430(.A0(new_n2865_), .A1(new_n2545_), .B0(new_n2836_), .Y(new_n2866_));
  OAI21X1  g00431(.A0(new_n2866_), .A1(pi0093), .B0(new_n2834_), .Y(new_n2867_));
  AOI21X1  g00432(.A0(new_n2867_), .A1(new_n2832_), .B0(new_n2850_), .Y(new_n2868_));
  OAI21X1  g00433(.A0(new_n2868_), .A1(new_n2853_), .B0(new_n2533_), .Y(new_n2869_));
  AOI21X1  g00434(.A0(new_n2869_), .A1(new_n2861_), .B0(new_n2860_), .Y(new_n2870_));
  AOI21X1  g00435(.A0(new_n2870_), .A1(new_n2856_), .B0(pi0095), .Y(new_n2871_));
  OAI21X1  g00436(.A0(new_n2871_), .A1(new_n2696_), .B0(new_n2452_), .Y(new_n2872_));
  OAI21X1  g00437(.A0(new_n2509_), .A1(pi0225), .B0(new_n2535_), .Y(new_n2873_));
  NOR3X1   g00438(.A(new_n2848_), .B(pi0096), .C(pi0051), .Y(new_n2874_));
  AND3X1   g00439(.A(new_n2874_), .B(new_n2873_), .C(new_n2456_), .Y(new_n2875_));
  INVX1    g00440(.A(new_n2695_), .Y(new_n2876_));
  NOR3X1   g00441(.A(new_n2876_), .B(new_n2690_), .C(pi0072), .Y(new_n2877_));
  NOR3X1   g00442(.A(new_n2877_), .B(new_n2875_), .C(pi0032), .Y(new_n2878_));
  NOR3X1   g00443(.A(new_n2878_), .B(new_n2860_), .C(pi0095), .Y(new_n2879_));
  AND3X1   g00444(.A(new_n2695_), .B(new_n2527_), .C(new_n2454_), .Y(new_n2880_));
  OR3X1    g00445(.A(new_n2880_), .B(new_n2879_), .C(new_n2452_), .Y(new_n2881_));
  AOI21X1  g00446(.A0(new_n2881_), .A1(new_n2872_), .B0(pi0210), .Y(new_n2882_));
  NAND2X1  g00447(.A(new_n2882_), .B(pi0146), .Y(new_n2883_));
  AND2X1   g00448(.A(new_n2854_), .B(new_n2533_), .Y(new_n2884_));
  OAI21X1  g00449(.A0(new_n2857_), .A1(pi0225), .B0(pi0032), .Y(new_n2885_));
  OAI21X1  g00450(.A0(new_n2884_), .A1(new_n2795_), .B0(new_n2885_), .Y(new_n2886_));
  AOI21X1  g00451(.A0(new_n2886_), .A1(new_n2523_), .B0(new_n2826_), .Y(new_n2887_));
  INVX1    g00452(.A(new_n2878_), .Y(new_n2888_));
  AND2X1   g00453(.A(new_n2885_), .B(new_n2523_), .Y(new_n2889_));
  AOI21X1  g00454(.A0(new_n2889_), .A1(new_n2888_), .B0(new_n2880_), .Y(new_n2890_));
  OAI21X1  g00455(.A0(new_n2890_), .A1(new_n2452_), .B0(pi0210), .Y(new_n2891_));
  OAI21X1  g00456(.A0(new_n2891_), .A1(new_n2887_), .B0(new_n2788_), .Y(new_n2892_));
  NOR2X1   g00457(.A(pi0210), .B(pi0146), .Y(new_n2893_));
  OAI21X1  g00458(.A0(new_n2860_), .A1(new_n2855_), .B0(new_n2523_), .Y(new_n2894_));
  AND2X1   g00459(.A(new_n2894_), .B(new_n2794_), .Y(new_n2895_));
  OAI21X1  g00460(.A0(new_n2895_), .A1(pi0137), .B0(new_n2881_), .Y(new_n2896_));
  AOI21X1  g00461(.A0(new_n2896_), .A1(new_n2893_), .B0(new_n2892_), .Y(new_n2897_));
  NAND2X1  g00462(.A(new_n2897_), .B(new_n2883_), .Y(new_n2898_));
  AND2X1   g00463(.A(new_n2859_), .B(new_n2523_), .Y(new_n2899_));
  OAI21X1  g00464(.A0(new_n2875_), .A1(pi0032), .B0(new_n2899_), .Y(new_n2900_));
  OAI21X1  g00465(.A0(new_n2851_), .A1(pi0072), .B0(new_n2533_), .Y(new_n2901_));
  NAND3X1  g00466(.A(new_n2901_), .B(new_n2831_), .C(new_n2528_), .Y(new_n2902_));
  OAI21X1  g00467(.A0(new_n2868_), .A1(pi0072), .B0(new_n2533_), .Y(new_n2903_));
  NAND2X1  g00468(.A(new_n2903_), .B(new_n2861_), .Y(new_n2904_));
  AND3X1   g00469(.A(new_n2904_), .B(new_n2902_), .C(new_n2859_), .Y(new_n2905_));
  OAI21X1  g00470(.A0(new_n2905_), .A1(pi0095), .B0(new_n2751_), .Y(new_n2906_));
  MX2X1    g00471(.A(new_n2906_), .B(new_n2900_), .S0(pi0137), .Y(new_n2907_));
  NAND2X1  g00472(.A(new_n2907_), .B(new_n2777_), .Y(new_n2908_));
  NAND2X1  g00473(.A(new_n2901_), .B(new_n2528_), .Y(new_n2909_));
  AOI21X1  g00474(.A0(new_n2909_), .A1(new_n2885_), .B0(pi0095), .Y(new_n2910_));
  NOR3X1   g00475(.A(new_n2696_), .B(new_n2454_), .C(pi0137), .Y(new_n2911_));
  INVX1    g00476(.A(new_n2911_), .Y(new_n2912_));
  AND3X1   g00477(.A(new_n2885_), .B(pi0137), .C(new_n2523_), .Y(new_n2913_));
  OAI21X1  g00478(.A0(new_n2875_), .A1(pi0032), .B0(new_n2913_), .Y(new_n2914_));
  AND2X1   g00479(.A(new_n2914_), .B(pi0210), .Y(new_n2915_));
  OAI21X1  g00480(.A0(new_n2912_), .A1(new_n2910_), .B0(new_n2915_), .Y(new_n2916_));
  NAND2X1  g00481(.A(new_n2916_), .B(new_n2774_), .Y(new_n2917_));
  AOI21X1  g00482(.A0(new_n2901_), .A1(new_n2528_), .B0(new_n2860_), .Y(new_n2918_));
  OAI21X1  g00483(.A0(new_n2918_), .A1(pi0095), .B0(new_n2751_), .Y(new_n2919_));
  MX2X1    g00484(.A(new_n2919_), .B(new_n2900_), .S0(pi0137), .Y(new_n2920_));
  AOI21X1  g00485(.A0(new_n2920_), .A1(new_n2893_), .B0(new_n2917_), .Y(new_n2921_));
  OAI21X1  g00486(.A0(new_n2908_), .A1(new_n2776_), .B0(new_n2921_), .Y(new_n2922_));
  AND3X1   g00487(.A(new_n2922_), .B(new_n2898_), .C(new_n2451_), .Y(new_n2923_));
  INVX1    g00488(.A(pi0153), .Y(new_n2924_));
  AOI21X1  g00489(.A0(new_n2907_), .A1(new_n2777_), .B0(new_n2917_), .Y(new_n2925_));
  OAI21X1  g00490(.A0(new_n2892_), .A1(new_n2882_), .B0(new_n2450_), .Y(new_n2926_));
  OAI21X1  g00491(.A0(new_n2926_), .A1(new_n2925_), .B0(new_n2924_), .Y(new_n2927_));
  OR2X1    g00492(.A(new_n2927_), .B(new_n2923_), .Y(new_n2928_));
  AND3X1   g00493(.A(new_n2928_), .B(new_n2830_), .C(new_n2793_), .Y(new_n2929_));
  AOI21X1  g00494(.A0(new_n2792_), .A1(pi0228), .B0(new_n2929_), .Y(new_n2930_));
  OAI21X1  g00495(.A0(new_n2930_), .A1(pi0216), .B0(new_n2446_), .Y(new_n2931_));
  AOI21X1  g00496(.A0(new_n2931_), .A1(new_n2437_), .B0(new_n2443_), .Y(new_n2932_));
  INVX1    g00497(.A(pi0299), .Y(new_n2933_));
  INVX1    g00498(.A(pi0215), .Y(new_n2934_));
  NOR2X1   g00499(.A(pi1144), .B(pi0332), .Y(new_n2935_));
  NOR2X1   g00500(.A(new_n2935_), .B(new_n2934_), .Y(new_n2936_));
  NOR2X1   g00501(.A(new_n2936_), .B(new_n2933_), .Y(new_n2937_));
  OAI21X1  g00502(.A0(new_n2932_), .A1(pi0215), .B0(new_n2937_), .Y(new_n2938_));
  INVX1    g00503(.A(pi0039), .Y(new_n2939_));
  INVX1    g00504(.A(pi0223), .Y(new_n2940_));
  INVX1    g00505(.A(pi0222), .Y(new_n2941_));
  INVX1    g00506(.A(pi0224), .Y(new_n2942_));
  AOI21X1  g00507(.A0(pi0833), .A1(new_n2942_), .B0(new_n2941_), .Y(new_n2943_));
  NOR2X1   g00508(.A(new_n2943_), .B(pi0223), .Y(new_n2944_));
  NOR3X1   g00509(.A(new_n2944_), .B(pi1144), .C(pi0332), .Y(new_n2945_));
  AOI21X1  g00510(.A0(new_n2444_), .A1(pi0265), .B0(new_n2942_), .Y(new_n2946_));
  OR4X1    g00511(.A(pi0929), .B(new_n2701_), .C(pi0332), .D(pi0224), .Y(new_n2947_));
  OAI21X1  g00512(.A0(new_n2946_), .A1(pi0222), .B0(new_n2947_), .Y(new_n2948_));
  AOI21X1  g00513(.A0(new_n2948_), .A1(new_n2940_), .B0(new_n2945_), .Y(new_n2949_));
  NOR2X1   g00514(.A(new_n2949_), .B(pi0299), .Y(new_n2950_));
  NOR2X1   g00515(.A(pi0224), .B(pi0222), .Y(new_n2951_));
  INVX1    g00516(.A(new_n2951_), .Y(new_n2952_));
  INVX1    g00517(.A(pi0142), .Y(new_n2953_));
  INVX1    g00518(.A(pi0198), .Y(new_n2954_));
  OR2X1    g00519(.A(new_n2700_), .B(new_n2954_), .Y(new_n2955_));
  OAI21X1  g00520(.A0(new_n2743_), .A1(pi0198), .B0(new_n2955_), .Y(new_n2956_));
  OAI21X1  g00521(.A0(new_n2717_), .A1(new_n2712_), .B0(new_n2954_), .Y(new_n2957_));
  NAND3X1  g00522(.A(new_n2957_), .B(new_n2955_), .C(new_n2953_), .Y(new_n2958_));
  AND2X1   g00523(.A(new_n2958_), .B(new_n2774_), .Y(new_n2959_));
  OAI21X1  g00524(.A0(new_n2956_), .A1(new_n2953_), .B0(new_n2959_), .Y(new_n2960_));
  NOR3X1   g00525(.A(pi0189), .B(pi0174), .C(pi0144), .Y(new_n2961_));
  NOR2X1   g00526(.A(new_n2961_), .B(pi0223), .Y(new_n2962_));
  INVX1    g00527(.A(new_n2962_), .Y(new_n2963_));
  NOR2X1   g00528(.A(new_n2754_), .B(new_n2750_), .Y(new_n2964_));
  MX2X1    g00529(.A(new_n2770_), .B(new_n2964_), .S0(pi0198), .Y(new_n2965_));
  NAND2X1  g00530(.A(new_n2965_), .B(pi0142), .Y(new_n2966_));
  INVX1    g00531(.A(new_n2788_), .Y(new_n2967_));
  OAI21X1  g00532(.A0(new_n2754_), .A1(new_n2750_), .B0(pi0198), .Y(new_n2968_));
  AOI21X1  g00533(.A0(new_n2785_), .A1(new_n2954_), .B0(pi0142), .Y(new_n2969_));
  AOI21X1  g00534(.A0(new_n2969_), .A1(new_n2968_), .B0(new_n2967_), .Y(new_n2970_));
  AOI21X1  g00535(.A0(new_n2970_), .A1(new_n2966_), .B0(new_n2963_), .Y(new_n2971_));
  NOR4X1   g00536(.A(pi0223), .B(pi0189), .C(pi0174), .D(pi0144), .Y(new_n2972_));
  INVX1    g00537(.A(pi0234), .Y(new_n2973_));
  AOI21X1  g00538(.A0(new_n2965_), .A1(new_n2973_), .B0(pi0332), .Y(new_n2974_));
  OAI21X1  g00539(.A0(new_n2956_), .A1(new_n2973_), .B0(new_n2974_), .Y(new_n2975_));
  AOI22X1  g00540(.A0(new_n2975_), .A1(new_n2972_), .B0(new_n2971_), .B1(new_n2960_), .Y(new_n2976_));
  OAI21X1  g00541(.A0(new_n2976_), .A1(new_n2952_), .B0(new_n2950_), .Y(new_n2977_));
  AND2X1   g00542(.A(new_n2977_), .B(new_n2939_), .Y(new_n2978_));
  INVX1    g00543(.A(pi0038), .Y(new_n2979_));
  AOI21X1  g00544(.A0(new_n2454_), .A1(pi0234), .B0(pi0332), .Y(new_n2980_));
  INVX1    g00545(.A(new_n2980_), .Y(new_n2981_));
  AND3X1   g00546(.A(new_n2695_), .B(new_n2527_), .C(new_n2523_), .Y(new_n2982_));
  OR2X1    g00547(.A(new_n2982_), .B(new_n2454_), .Y(new_n2983_));
  NOR4X1   g00548(.A(pi0095), .B(pi0072), .C(pi0040), .D(pi0032), .Y(new_n2984_));
  NAND3X1  g00549(.A(new_n2984_), .B(new_n2513_), .C(new_n2534_), .Y(new_n2985_));
  OR2X1    g00550(.A(new_n2985_), .B(new_n2536_), .Y(new_n2986_));
  INVX1    g00551(.A(new_n2986_), .Y(new_n2987_));
  MX2X1    g00552(.A(new_n2987_), .B(new_n2983_), .S0(pi0234), .Y(new_n2988_));
  AOI21X1  g00553(.A0(new_n2988_), .A1(pi0137), .B0(new_n2981_), .Y(new_n2989_));
  NOR3X1   g00554(.A(pi0224), .B(pi0223), .C(pi0222), .Y(new_n2990_));
  INVX1    g00555(.A(new_n2990_), .Y(new_n2991_));
  NOR2X1   g00556(.A(new_n2991_), .B(new_n2989_), .Y(new_n2992_));
  NOR2X1   g00557(.A(new_n2992_), .B(new_n2949_), .Y(new_n2993_));
  INVX1    g00558(.A(new_n2443_), .Y(new_n2994_));
  MX2X1    g00559(.A(new_n2989_), .B(new_n2448_), .S0(new_n2447_), .Y(new_n2995_));
  INVX1    g00560(.A(new_n2982_), .Y(new_n2996_));
  NOR4X1   g00561(.A(new_n2996_), .B(pi0332), .C(pi0153), .D(pi0137), .Y(new_n2997_));
  NOR3X1   g00562(.A(new_n2985_), .B(new_n2536_), .C(new_n2452_), .Y(new_n2998_));
  OAI21X1  g00563(.A0(new_n2998_), .A1(new_n2449_), .B0(new_n2793_), .Y(new_n2999_));
  OAI22X1  g00564(.A0(new_n2999_), .A1(new_n2997_), .B0(new_n2995_), .B1(new_n2793_), .Y(new_n3000_));
  AOI21X1  g00565(.A0(new_n3000_), .A1(new_n2438_), .B0(new_n2445_), .Y(new_n3001_));
  OAI21X1  g00566(.A0(new_n3001_), .A1(pi0221), .B0(new_n2994_), .Y(new_n3002_));
  AOI21X1  g00567(.A0(new_n3002_), .A1(new_n2934_), .B0(new_n2936_), .Y(new_n3003_));
  MX2X1    g00568(.A(new_n3003_), .B(new_n2993_), .S0(new_n2933_), .Y(new_n3004_));
  OAI21X1  g00569(.A0(new_n3004_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n3005_));
  AOI21X1  g00570(.A0(new_n2978_), .A1(new_n2938_), .B0(new_n3005_), .Y(new_n3006_));
  INVX1    g00571(.A(pi0100), .Y(new_n3007_));
  OAI21X1  g00572(.A0(new_n2992_), .A1(new_n2949_), .B0(new_n2933_), .Y(new_n3008_));
  AND2X1   g00573(.A(pi0228), .B(pi0105), .Y(new_n3009_));
  AND2X1   g00574(.A(new_n3009_), .B(new_n2980_), .Y(new_n3010_));
  INVX1    g00575(.A(new_n3009_), .Y(new_n3011_));
  AOI21X1  g00576(.A0(new_n3011_), .A1(new_n2448_), .B0(pi0216), .Y(new_n3012_));
  INVX1    g00577(.A(new_n3012_), .Y(new_n3013_));
  OAI21X1  g00578(.A0(new_n3013_), .A1(new_n3010_), .B0(new_n2446_), .Y(new_n3014_));
  AOI21X1  g00579(.A0(new_n3014_), .A1(new_n2437_), .B0(new_n2443_), .Y(new_n3015_));
  MX2X1    g00580(.A(new_n3015_), .B(new_n2935_), .S0(pi0215), .Y(new_n3016_));
  INVX1    g00581(.A(new_n3016_), .Y(new_n3017_));
  NOR2X1   g00582(.A(pi0221), .B(pi0215), .Y(new_n3018_));
  INVX1    g00583(.A(new_n3018_), .Y(new_n3019_));
  NOR3X1   g00584(.A(new_n3019_), .B(new_n3013_), .C(new_n2989_), .Y(new_n3020_));
  OAI21X1  g00585(.A0(new_n3020_), .A1(new_n3017_), .B0(pi0299), .Y(new_n3021_));
  AOI21X1  g00586(.A0(new_n3021_), .A1(new_n3008_), .B0(pi0039), .Y(new_n3022_));
  NOR2X1   g00587(.A(new_n2991_), .B(new_n2980_), .Y(new_n3023_));
  NOR3X1   g00588(.A(new_n3023_), .B(new_n2949_), .C(pi0299), .Y(new_n3024_));
  AOI21X1  g00589(.A0(new_n3016_), .A1(pi0299), .B0(new_n3024_), .Y(new_n3025_));
  INVX1    g00590(.A(new_n3025_), .Y(new_n3026_));
  OAI21X1  g00591(.A0(new_n3026_), .A1(new_n2939_), .B0(pi0038), .Y(new_n3027_));
  OAI21X1  g00592(.A0(new_n3027_), .A1(new_n3022_), .B0(new_n3007_), .Y(new_n3028_));
  AOI21X1  g00593(.A0(new_n2449_), .A1(new_n2447_), .B0(new_n2793_), .Y(new_n3029_));
  AOI21X1  g00594(.A0(pi0234), .A1(pi0095), .B0(pi0137), .Y(new_n3030_));
  OAI21X1  g00595(.A0(new_n2815_), .A1(pi0210), .B0(new_n3030_), .Y(new_n3031_));
  AOI21X1  g00596(.A0(new_n3031_), .A1(new_n2988_), .B0(pi0332), .Y(new_n3032_));
  OAI21X1  g00597(.A0(new_n3032_), .A1(new_n2447_), .B0(new_n3029_), .Y(new_n3033_));
  INVX1    g00598(.A(new_n2997_), .Y(new_n3034_));
  INVX1    g00599(.A(pi0252), .Y(new_n3035_));
  OAI21X1  g00600(.A0(new_n2777_), .A1(pi0137), .B0(new_n3035_), .Y(new_n3036_));
  NOR4X1   g00601(.A(new_n3036_), .B(new_n2996_), .C(new_n2815_), .D(pi0332), .Y(new_n3037_));
  INVX1    g00602(.A(new_n2815_), .Y(new_n3038_));
  NOR4X1   g00603(.A(new_n2985_), .B(new_n3038_), .C(new_n2536_), .D(new_n2452_), .Y(new_n3039_));
  OR2X1    g00604(.A(new_n3039_), .B(new_n2449_), .Y(new_n3040_));
  AOI21X1  g00605(.A0(new_n3035_), .A1(pi0210), .B0(new_n2815_), .Y(new_n3041_));
  OAI22X1  g00606(.A0(new_n3041_), .A1(new_n3034_), .B0(new_n3040_), .B1(new_n3037_), .Y(new_n3042_));
  AOI21X1  g00607(.A0(new_n3042_), .A1(new_n2793_), .B0(pi0216), .Y(new_n3043_));
  AOI21X1  g00608(.A0(new_n3043_), .A1(new_n3033_), .B0(new_n2445_), .Y(new_n3044_));
  OAI21X1  g00609(.A0(new_n3044_), .A1(pi0221), .B0(new_n2994_), .Y(new_n3045_));
  AOI21X1  g00610(.A0(new_n3045_), .A1(new_n2934_), .B0(new_n2936_), .Y(new_n3046_));
  NOR2X1   g00611(.A(pi0039), .B(pi0038), .Y(new_n3047_));
  OAI21X1  g00612(.A0(pi0198), .A1(new_n2953_), .B0(new_n2452_), .Y(new_n3048_));
  AOI21X1  g00613(.A0(new_n3048_), .A1(new_n2988_), .B0(new_n2981_), .Y(new_n3049_));
  INVX1    g00614(.A(new_n2774_), .Y(new_n3050_));
  OR3X1    g00615(.A(new_n2954_), .B(pi0137), .C(pi0095), .Y(new_n3051_));
  AOI21X1  g00616(.A0(new_n3051_), .A1(new_n2983_), .B0(new_n3050_), .Y(new_n3052_));
  AOI21X1  g00617(.A0(pi0198), .A1(new_n2452_), .B0(new_n2986_), .Y(new_n3053_));
  OAI21X1  g00618(.A0(new_n3053_), .A1(new_n2967_), .B0(new_n2972_), .Y(new_n3054_));
  OAI22X1  g00619(.A0(new_n3054_), .A1(new_n3052_), .B0(new_n3049_), .B1(new_n2963_), .Y(new_n3055_));
  AOI21X1  g00620(.A0(new_n3055_), .A1(new_n2951_), .B0(new_n2949_), .Y(new_n3056_));
  OR2X1    g00621(.A(new_n3056_), .B(pi0299), .Y(new_n3057_));
  AND2X1   g00622(.A(new_n3057_), .B(new_n3047_), .Y(new_n3058_));
  OAI21X1  g00623(.A0(new_n3046_), .A1(new_n2933_), .B0(new_n3058_), .Y(new_n3059_));
  INVX1    g00624(.A(new_n3047_), .Y(new_n3060_));
  AOI21X1  g00625(.A0(new_n3060_), .A1(new_n3026_), .B0(new_n3007_), .Y(new_n3061_));
  AOI21X1  g00626(.A0(new_n3061_), .A1(new_n3059_), .B0(pi0087), .Y(new_n3062_));
  OAI21X1  g00627(.A0(new_n3028_), .A1(new_n3006_), .B0(new_n3062_), .Y(new_n3063_));
  NOR3X1   g00628(.A(pi0100), .B(pi0039), .C(pi0038), .Y(new_n3064_));
  MX2X1    g00629(.A(new_n3026_), .B(new_n3004_), .S0(new_n3064_), .Y(new_n3065_));
  AOI21X1  g00630(.A0(new_n3065_), .A1(pi0087), .B0(pi0075), .Y(new_n3066_));
  AOI21X1  g00631(.A0(new_n3033_), .A1(new_n3012_), .B0(new_n2445_), .Y(new_n3067_));
  OAI21X1  g00632(.A0(new_n3067_), .A1(pi0221), .B0(new_n2994_), .Y(new_n3068_));
  AOI21X1  g00633(.A0(new_n3068_), .A1(new_n2934_), .B0(new_n2936_), .Y(new_n3069_));
  NOR4X1   g00634(.A(pi0100), .B(pi0087), .C(pi0039), .D(pi0038), .Y(new_n3070_));
  AND2X1   g00635(.A(new_n3070_), .B(new_n3057_), .Y(new_n3071_));
  OAI21X1  g00636(.A0(new_n3069_), .A1(new_n2933_), .B0(new_n3071_), .Y(new_n3072_));
  INVX1    g00637(.A(pi0075), .Y(new_n3073_));
  INVX1    g00638(.A(new_n3070_), .Y(new_n3074_));
  AOI21X1  g00639(.A0(new_n3074_), .A1(new_n3026_), .B0(new_n3073_), .Y(new_n3075_));
  AOI22X1  g00640(.A0(new_n3075_), .A1(new_n3072_), .B0(new_n3066_), .B1(new_n3063_), .Y(new_n3076_));
  NOR2X1   g00641(.A(pi0087), .B(pi0075), .Y(new_n3077_));
  NAND2X1  g00642(.A(new_n3077_), .B(new_n3065_), .Y(new_n3078_));
  INVX1    g00643(.A(pi0092), .Y(new_n3079_));
  INVX1    g00644(.A(new_n3077_), .Y(new_n3080_));
  AOI21X1  g00645(.A0(new_n3080_), .A1(new_n3026_), .B0(new_n3079_), .Y(new_n3081_));
  AOI21X1  g00646(.A0(new_n3081_), .A1(new_n3078_), .B0(pi0054), .Y(new_n3082_));
  OAI21X1  g00647(.A0(new_n3076_), .A1(pi0092), .B0(new_n3082_), .Y(new_n3083_));
  NOR2X1   g00648(.A(pi0092), .B(pi0075), .Y(new_n3084_));
  AND2X1   g00649(.A(new_n3084_), .B(new_n3070_), .Y(new_n3085_));
  INVX1    g00650(.A(new_n3085_), .Y(new_n3086_));
  NOR3X1   g00651(.A(pi0100), .B(pi0087), .C(pi0038), .Y(new_n3087_));
  AND2X1   g00652(.A(new_n3087_), .B(new_n3084_), .Y(new_n3088_));
  AOI22X1  g00653(.A0(new_n3088_), .A1(new_n3022_), .B0(new_n3086_), .B1(new_n3025_), .Y(new_n3089_));
  AOI21X1  g00654(.A0(new_n3089_), .A1(pi0054), .B0(pi0074), .Y(new_n3090_));
  INVX1    g00655(.A(pi0054), .Y(new_n3091_));
  OAI21X1  g00656(.A0(new_n3025_), .A1(new_n3091_), .B0(pi0074), .Y(new_n3092_));
  AOI21X1  g00657(.A0(new_n3089_), .A1(new_n3091_), .B0(new_n3092_), .Y(new_n3093_));
  AOI21X1  g00658(.A0(new_n3090_), .A1(new_n3083_), .B0(new_n3093_), .Y(new_n3094_));
  OAI21X1  g00659(.A0(new_n2988_), .A1(pi0332), .B0(pi0105), .Y(new_n3095_));
  AND3X1   g00660(.A(new_n2986_), .B(new_n2448_), .C(new_n2793_), .Y(new_n3096_));
  OR2X1    g00661(.A(new_n3096_), .B(pi0216), .Y(new_n3097_));
  AOI21X1  g00662(.A0(new_n3095_), .A1(new_n3029_), .B0(new_n3097_), .Y(new_n3098_));
  OAI21X1  g00663(.A0(new_n3098_), .A1(new_n2445_), .B0(new_n2437_), .Y(new_n3099_));
  AOI21X1  g00664(.A0(new_n3099_), .A1(new_n2994_), .B0(pi0215), .Y(new_n3100_));
  NOR2X1   g00665(.A(pi0100), .B(pi0087), .Y(new_n3101_));
  NOR2X1   g00666(.A(pi0074), .B(pi0054), .Y(new_n3102_));
  AND3X1   g00667(.A(new_n3102_), .B(new_n3101_), .C(new_n3084_), .Y(new_n3103_));
  AND2X1   g00668(.A(new_n3103_), .B(new_n3047_), .Y(new_n3104_));
  INVX1    g00669(.A(new_n3104_), .Y(new_n3105_));
  OR3X1    g00670(.A(new_n3105_), .B(new_n3100_), .C(new_n2936_), .Y(new_n3106_));
  INVX1    g00671(.A(pi0055), .Y(new_n3107_));
  AOI21X1  g00672(.A0(new_n3105_), .A1(new_n3016_), .B0(new_n3107_), .Y(new_n3108_));
  AOI21X1  g00673(.A0(new_n3108_), .A1(new_n3106_), .B0(pi0056), .Y(new_n3109_));
  OAI21X1  g00674(.A0(new_n3094_), .A1(pi0055), .B0(new_n3109_), .Y(new_n3110_));
  NOR3X1   g00675(.A(pi0100), .B(pi0039), .C(pi0038), .Y(new_n3111_));
  OR3X1    g00676(.A(pi0092), .B(pi0087), .C(pi0075), .Y(new_n3112_));
  NOR4X1   g00677(.A(new_n3112_), .B(pi0074), .C(pi0055), .D(pi0054), .Y(new_n3113_));
  AND2X1   g00678(.A(new_n3113_), .B(new_n3111_), .Y(new_n3114_));
  INVX1    g00679(.A(new_n3114_), .Y(new_n3115_));
  MX2X1    g00680(.A(new_n3003_), .B(new_n3016_), .S0(new_n3115_), .Y(new_n3116_));
  AOI21X1  g00681(.A0(new_n3116_), .A1(pi0056), .B0(pi0062), .Y(new_n3117_));
  INVX1    g00682(.A(pi0056), .Y(new_n3118_));
  OAI21X1  g00683(.A0(new_n3017_), .A1(new_n3118_), .B0(pi0062), .Y(new_n3119_));
  AOI21X1  g00684(.A0(new_n3116_), .A1(new_n3118_), .B0(new_n3119_), .Y(new_n3120_));
  OR2X1    g00685(.A(new_n3120_), .B(pi0059), .Y(new_n3121_));
  AOI21X1  g00686(.A0(new_n3117_), .A1(new_n3110_), .B0(new_n3121_), .Y(new_n3122_));
  NOR2X1   g00687(.A(pi0062), .B(pi0056), .Y(new_n3123_));
  AND3X1   g00688(.A(new_n3123_), .B(new_n3114_), .C(new_n3020_), .Y(new_n3124_));
  NAND2X1  g00689(.A(new_n3016_), .B(pi0059), .Y(new_n3125_));
  OAI21X1  g00690(.A0(new_n3125_), .A1(new_n3124_), .B0(new_n2436_), .Y(new_n3126_));
  INVX1    g00691(.A(pi0059), .Y(new_n3127_));
  AOI21X1  g00692(.A0(new_n3124_), .A1(new_n3127_), .B0(new_n3017_), .Y(new_n3128_));
  OAI22X1  g00693(.A0(new_n3128_), .A1(new_n2436_), .B0(new_n3126_), .B1(new_n3122_), .Y(po0153));
  INVX1    g00694(.A(new_n3102_), .Y(new_n3130_));
  INVX1    g00695(.A(pi0087), .Y(new_n3131_));
  INVX1    g00696(.A(new_n3064_), .Y(new_n3132_));
  INVX1    g00697(.A(pi0154), .Y(new_n3133_));
  AND2X1   g00698(.A(pi0833), .B(new_n2942_), .Y(new_n3134_));
  INVX1    g00699(.A(pi0939), .Y(new_n3135_));
  AOI21X1  g00700(.A0(new_n3134_), .A1(new_n3135_), .B0(new_n2941_), .Y(new_n3136_));
  OAI21X1  g00701(.A0(new_n3134_), .A1(pi1146), .B0(new_n3136_), .Y(new_n3137_));
  AND2X1   g00702(.A(pi0224), .B(new_n2941_), .Y(new_n3138_));
  AOI21X1  g00703(.A0(new_n3138_), .A1(pi0276), .B0(pi0223), .Y(new_n3139_));
  INVX1    g00704(.A(pi1146), .Y(new_n3140_));
  AOI21X1  g00705(.A0(new_n3140_), .A1(pi0223), .B0(pi0299), .Y(new_n3141_));
  INVX1    g00706(.A(new_n3141_), .Y(new_n3142_));
  AOI21X1  g00707(.A0(new_n3139_), .A1(new_n3137_), .B0(new_n3142_), .Y(new_n3143_));
  INVX1    g00708(.A(new_n3143_), .Y(new_n3144_));
  AND2X1   g00709(.A(pi0833), .B(new_n2438_), .Y(new_n3145_));
  AOI21X1  g00710(.A0(new_n3145_), .A1(new_n3135_), .B0(new_n2437_), .Y(new_n3146_));
  OAI21X1  g00711(.A0(new_n3145_), .A1(pi1146), .B0(new_n3146_), .Y(new_n3147_));
  OAI21X1  g00712(.A0(new_n3140_), .A1(new_n2934_), .B0(new_n3147_), .Y(new_n3148_));
  NOR4X1   g00713(.A(new_n3148_), .B(new_n2986_), .C(pi0228), .D(pi0216), .Y(new_n3149_));
  OAI21X1  g00714(.A0(new_n2701_), .A1(pi0216), .B0(new_n3140_), .Y(new_n3150_));
  INVX1    g00715(.A(pi0276), .Y(new_n3151_));
  AND2X1   g00716(.A(new_n2437_), .B(pi0216), .Y(new_n3152_));
  INVX1    g00717(.A(new_n3152_), .Y(new_n3153_));
  OAI22X1  g00718(.A0(new_n3153_), .A1(new_n3151_), .B0(new_n3009_), .B1(pi0216), .Y(new_n3154_));
  AOI22X1  g00719(.A0(new_n3154_), .A1(new_n2437_), .B0(new_n3146_), .B1(new_n3150_), .Y(new_n3155_));
  MX2X1    g00720(.A(new_n3155_), .B(new_n3140_), .S0(pi0215), .Y(new_n3156_));
  OR2X1    g00721(.A(new_n3156_), .B(new_n2933_), .Y(new_n3157_));
  OAI21X1  g00722(.A0(new_n3157_), .A1(new_n3149_), .B0(new_n3144_), .Y(new_n3158_));
  OAI21X1  g00723(.A0(new_n3153_), .A1(new_n3151_), .B0(new_n3147_), .Y(new_n3159_));
  MX2X1    g00724(.A(new_n3159_), .B(pi1146), .S0(pi0215), .Y(new_n3160_));
  AOI21X1  g00725(.A0(new_n3160_), .A1(pi0299), .B0(new_n3143_), .Y(new_n3161_));
  OAI21X1  g00726(.A0(new_n3161_), .A1(new_n3133_), .B0(new_n3064_), .Y(new_n3162_));
  AOI21X1  g00727(.A0(new_n3158_), .A1(new_n3133_), .B0(new_n3162_), .Y(new_n3163_));
  INVX1    g00728(.A(new_n3160_), .Y(new_n3164_));
  MX2X1    g00729(.A(new_n3164_), .B(new_n3156_), .S0(new_n3133_), .Y(new_n3165_));
  INVX1    g00730(.A(new_n3165_), .Y(new_n3166_));
  AOI21X1  g00731(.A0(new_n3166_), .A1(pi0299), .B0(new_n3143_), .Y(new_n3167_));
  AOI21X1  g00732(.A0(new_n3167_), .A1(new_n3132_), .B0(new_n3163_), .Y(new_n3168_));
  AND2X1   g00733(.A(new_n2986_), .B(pi0039), .Y(new_n3169_));
  INVX1    g00734(.A(new_n2537_), .Y(new_n3170_));
  AOI22X1  g00735(.A0(new_n2689_), .A1(pi0070), .B0(new_n2506_), .B1(pi0035), .Y(new_n3171_));
  OAI21X1  g00736(.A0(new_n2799_), .A1(pi0070), .B0(new_n3171_), .Y(new_n3172_));
  AOI21X1  g00737(.A0(new_n3172_), .A1(new_n2534_), .B0(new_n3170_), .Y(new_n3173_));
  OAI21X1  g00738(.A0(new_n3173_), .A1(new_n2853_), .B0(new_n2532_), .Y(new_n3174_));
  OR2X1    g00739(.A(new_n2527_), .B(new_n2529_), .Y(new_n3175_));
  OR2X1    g00740(.A(new_n2480_), .B(new_n2455_), .Y(new_n3176_));
  AND2X1   g00741(.A(new_n3176_), .B(new_n3175_), .Y(new_n3177_));
  INVX1    g00742(.A(new_n3177_), .Y(new_n3178_));
  AOI21X1  g00743(.A0(new_n3174_), .A1(new_n2695_), .B0(new_n3178_), .Y(new_n3179_));
  OAI21X1  g00744(.A0(new_n3179_), .A1(pi0095), .B0(new_n2794_), .Y(new_n3180_));
  AOI21X1  g00745(.A0(new_n3180_), .A1(new_n2939_), .B0(new_n3169_), .Y(new_n3181_));
  NOR3X1   g00746(.A(new_n3148_), .B(pi0228), .C(pi0216), .Y(new_n3182_));
  AOI21X1  g00747(.A0(new_n3182_), .A1(new_n3181_), .B0(new_n3157_), .Y(new_n3183_));
  OAI21X1  g00748(.A0(new_n3183_), .A1(new_n3143_), .B0(new_n3133_), .Y(new_n3184_));
  OR2X1    g00749(.A(new_n3161_), .B(new_n3133_), .Y(new_n3185_));
  AND2X1   g00750(.A(new_n3185_), .B(new_n2979_), .Y(new_n3186_));
  INVX1    g00751(.A(new_n3167_), .Y(new_n3187_));
  OAI21X1  g00752(.A0(new_n3187_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3188_));
  AOI21X1  g00753(.A0(new_n3186_), .A1(new_n3184_), .B0(new_n3188_), .Y(new_n3189_));
  AOI21X1  g00754(.A0(pi0252), .A1(pi0146), .B0(new_n2986_), .Y(new_n3190_));
  INVX1    g00755(.A(new_n3190_), .Y(new_n3191_));
  OR2X1    g00756(.A(pi0166), .B(pi0161), .Y(new_n3192_));
  INVX1    g00757(.A(pi0152), .Y(new_n3193_));
  NOR3X1   g00758(.A(new_n2985_), .B(new_n2536_), .C(pi0252), .Y(new_n3194_));
  INVX1    g00759(.A(new_n3194_), .Y(new_n3195_));
  OAI21X1  g00760(.A0(new_n3192_), .A1(new_n3195_), .B0(new_n3193_), .Y(new_n3196_));
  AOI21X1  g00761(.A0(new_n3192_), .A1(new_n3190_), .B0(new_n3196_), .Y(new_n3197_));
  AOI21X1  g00762(.A0(new_n3191_), .A1(pi0152), .B0(new_n3197_), .Y(new_n3198_));
  INVX1    g00763(.A(new_n3198_), .Y(new_n3199_));
  OR3X1    g00764(.A(pi0228), .B(pi0216), .C(pi0038), .Y(new_n3200_));
  OR4X1    g00765(.A(new_n3200_), .B(new_n2933_), .C(pi0154), .D(pi0039), .Y(new_n3201_));
  NOR3X1   g00766(.A(new_n3201_), .B(new_n3199_), .C(new_n3148_), .Y(new_n3202_));
  OR2X1    g00767(.A(new_n3167_), .B(new_n3007_), .Y(new_n3203_));
  OAI21X1  g00768(.A0(new_n3203_), .A1(new_n3202_), .B0(new_n3131_), .Y(new_n3204_));
  OAI22X1  g00769(.A0(new_n3204_), .A1(new_n3189_), .B0(new_n3168_), .B1(new_n3131_), .Y(new_n3205_));
  OAI21X1  g00770(.A0(new_n3187_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3206_));
  AOI21X1  g00771(.A0(new_n3205_), .A1(new_n3073_), .B0(new_n3206_), .Y(new_n3207_));
  AND2X1   g00772(.A(new_n3111_), .B(new_n3077_), .Y(new_n3208_));
  OAI21X1  g00773(.A0(new_n3208_), .A1(new_n3187_), .B0(pi0092), .Y(new_n3209_));
  AOI21X1  g00774(.A0(new_n3163_), .A1(new_n3077_), .B0(new_n3209_), .Y(new_n3210_));
  NOR3X1   g00775(.A(new_n3210_), .B(new_n3207_), .C(new_n3130_), .Y(new_n3211_));
  OAI21X1  g00776(.A0(new_n3187_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n3212_));
  OAI21X1  g00777(.A0(new_n3164_), .A1(new_n3133_), .B0(new_n3149_), .Y(new_n3213_));
  NOR2X1   g00778(.A(new_n3165_), .B(new_n3107_), .Y(new_n3214_));
  OAI21X1  g00779(.A0(new_n3213_), .A1(new_n3105_), .B0(new_n3214_), .Y(new_n3215_));
  AND2X1   g00780(.A(new_n3215_), .B(new_n3118_), .Y(new_n3216_));
  OAI21X1  g00781(.A0(new_n3212_), .A1(new_n3211_), .B0(new_n3216_), .Y(new_n3217_));
  NOR3X1   g00782(.A(new_n3165_), .B(new_n3105_), .C(pi0055), .Y(new_n3218_));
  NAND2X1  g00783(.A(new_n3218_), .B(new_n3213_), .Y(new_n3219_));
  AOI21X1  g00784(.A0(new_n3166_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n3220_));
  AOI21X1  g00785(.A0(new_n3220_), .A1(new_n3219_), .B0(pi0062), .Y(new_n3221_));
  INVX1    g00786(.A(pi0062), .Y(new_n3222_));
  NOR2X1   g00787(.A(pi0059), .B(pi0057), .Y(new_n3223_));
  AND3X1   g00788(.A(new_n3113_), .B(new_n3111_), .C(new_n3118_), .Y(new_n3224_));
  INVX1    g00789(.A(new_n3224_), .Y(new_n3225_));
  AOI22X1  g00790(.A0(new_n3225_), .A1(new_n3166_), .B0(new_n3218_), .B1(new_n3213_), .Y(new_n3226_));
  OAI21X1  g00791(.A0(new_n3226_), .A1(new_n3222_), .B0(new_n3223_), .Y(new_n3227_));
  AOI21X1  g00792(.A0(new_n3221_), .A1(new_n3217_), .B0(new_n3227_), .Y(new_n3228_));
  INVX1    g00793(.A(pi0239), .Y(new_n3229_));
  OAI21X1  g00794(.A0(new_n3223_), .A1(new_n3166_), .B0(new_n3229_), .Y(new_n3230_));
  AND3X1   g00795(.A(new_n2984_), .B(new_n2519_), .C(pi0096), .Y(new_n3231_));
  NOR2X1   g00796(.A(new_n3231_), .B(new_n2454_), .Y(new_n3232_));
  OAI21X1  g00797(.A0(pi0276), .A1(new_n2942_), .B0(new_n2941_), .Y(new_n3233_));
  AOI21X1  g00798(.A0(new_n3232_), .A1(new_n2942_), .B0(new_n3233_), .Y(new_n3234_));
  NAND2X1  g00799(.A(new_n3137_), .B(new_n2940_), .Y(new_n3235_));
  OAI22X1  g00800(.A0(new_n3235_), .A1(new_n3234_), .B0(pi1146), .B1(new_n2940_), .Y(new_n3236_));
  INVX1    g00801(.A(new_n2751_), .Y(new_n3237_));
  MX2X1    g00802(.A(new_n3173_), .B(new_n2531_), .S0(pi0072), .Y(new_n3238_));
  OAI21X1  g00803(.A0(new_n3238_), .A1(new_n2876_), .B0(new_n3177_), .Y(new_n3239_));
  AOI21X1  g00804(.A0(new_n3239_), .A1(new_n2523_), .B0(new_n3237_), .Y(new_n3240_));
  AOI22X1  g00805(.A0(new_n3240_), .A1(new_n2793_), .B0(new_n3232_), .B1(new_n3009_), .Y(new_n3241_));
  NOR3X1   g00806(.A(pi0221), .B(pi0216), .C(pi0215), .Y(new_n3242_));
  NOR2X1   g00807(.A(new_n3232_), .B(new_n2447_), .Y(new_n3243_));
  NOR2X1   g00808(.A(new_n3232_), .B(new_n2696_), .Y(new_n3244_));
  MX2X1    g00809(.A(new_n3244_), .B(new_n3243_), .S0(pi0228), .Y(new_n3245_));
  OR2X1    g00810(.A(new_n3245_), .B(new_n3133_), .Y(new_n3246_));
  AND2X1   g00811(.A(new_n3246_), .B(new_n3242_), .Y(new_n3247_));
  OAI21X1  g00812(.A0(new_n3241_), .A1(pi0154), .B0(new_n3247_), .Y(new_n3248_));
  NOR2X1   g00813(.A(new_n3160_), .B(new_n2933_), .Y(new_n3249_));
  AOI22X1  g00814(.A0(new_n3249_), .A1(new_n3248_), .B0(new_n3236_), .B1(new_n2933_), .Y(new_n3250_));
  NOR2X1   g00815(.A(pi0100), .B(pi0038), .Y(new_n3251_));
  INVX1    g00816(.A(new_n3251_), .Y(new_n3252_));
  OR2X1    g00817(.A(new_n3156_), .B(pi0154), .Y(new_n3253_));
  AND3X1   g00818(.A(new_n3009_), .B(new_n2453_), .C(pi0095), .Y(new_n3254_));
  AND2X1   g00819(.A(new_n3254_), .B(new_n3242_), .Y(new_n3255_));
  OAI21X1  g00820(.A0(new_n3255_), .A1(new_n3160_), .B0(new_n2934_), .Y(new_n3256_));
  INVX1    g00821(.A(new_n3255_), .Y(new_n3257_));
  AOI21X1  g00822(.A0(new_n3257_), .A1(new_n3164_), .B0(new_n3133_), .Y(new_n3258_));
  INVX1    g00823(.A(new_n3258_), .Y(new_n3259_));
  AND3X1   g00824(.A(new_n3259_), .B(new_n3256_), .C(new_n3253_), .Y(new_n3260_));
  OR4X1    g00825(.A(pi0299), .B(pi0224), .C(pi0223), .D(pi0222), .Y(new_n3261_));
  NOR3X1   g00826(.A(new_n3261_), .B(pi0479), .C(new_n2523_), .Y(new_n3262_));
  NOR2X1   g00827(.A(new_n3262_), .B(new_n3143_), .Y(new_n3263_));
  OAI21X1  g00828(.A0(new_n3260_), .A1(new_n2933_), .B0(new_n3263_), .Y(new_n3264_));
  AND2X1   g00829(.A(new_n3259_), .B(new_n3149_), .Y(new_n3265_));
  OAI21X1  g00830(.A0(new_n3265_), .A1(new_n3260_), .B0(pi0299), .Y(new_n3266_));
  AOI21X1  g00831(.A0(new_n3266_), .A1(new_n3264_), .B0(new_n2939_), .Y(new_n3267_));
  NOR2X1   g00832(.A(new_n3267_), .B(new_n3252_), .Y(new_n3268_));
  OAI21X1  g00833(.A0(new_n3250_), .A1(pi0039), .B0(new_n3268_), .Y(new_n3269_));
  INVX1    g00834(.A(new_n3264_), .Y(new_n3270_));
  NOR4X1   g00835(.A(new_n3201_), .B(new_n3199_), .C(new_n3148_), .D(new_n3007_), .Y(new_n3271_));
  OR3X1    g00836(.A(new_n3271_), .B(new_n3270_), .C(new_n3251_), .Y(new_n3272_));
  AOI21X1  g00837(.A0(new_n3272_), .A1(new_n3269_), .B0(pi0087), .Y(new_n3273_));
  NOR2X1   g00838(.A(new_n3266_), .B(new_n3132_), .Y(new_n3274_));
  NAND2X1  g00839(.A(new_n3264_), .B(pi0087), .Y(new_n3275_));
  OAI21X1  g00840(.A0(new_n3275_), .A1(new_n3274_), .B0(new_n3073_), .Y(new_n3276_));
  AOI21X1  g00841(.A0(new_n3270_), .A1(pi0075), .B0(pi0092), .Y(new_n3277_));
  OAI21X1  g00842(.A0(new_n3276_), .A1(new_n3273_), .B0(new_n3277_), .Y(new_n3278_));
  INVX1    g00843(.A(new_n3208_), .Y(new_n3279_));
  OR2X1    g00844(.A(new_n3266_), .B(new_n3279_), .Y(new_n3280_));
  AND2X1   g00845(.A(new_n3264_), .B(pi0092), .Y(new_n3281_));
  AOI21X1  g00846(.A0(new_n3281_), .A1(new_n3280_), .B0(new_n3130_), .Y(new_n3282_));
  OAI21X1  g00847(.A0(new_n3264_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n3283_));
  AOI21X1  g00848(.A0(new_n3282_), .A1(new_n3278_), .B0(new_n3283_), .Y(new_n3284_));
  AND3X1   g00849(.A(new_n3259_), .B(new_n3149_), .C(new_n3104_), .Y(new_n3285_));
  NOR3X1   g00850(.A(new_n3285_), .B(new_n3260_), .C(new_n3107_), .Y(new_n3286_));
  OR3X1    g00851(.A(new_n3286_), .B(new_n3284_), .C(pi0056), .Y(new_n3287_));
  NOR4X1   g00852(.A(new_n3265_), .B(new_n3260_), .C(new_n3105_), .D(pi0055), .Y(new_n3288_));
  INVX1    g00853(.A(new_n3288_), .Y(new_n3289_));
  INVX1    g00854(.A(new_n3260_), .Y(new_n3290_));
  AOI21X1  g00855(.A0(new_n3290_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n3291_));
  AOI21X1  g00856(.A0(new_n3291_), .A1(new_n3289_), .B0(pi0062), .Y(new_n3292_));
  AOI22X1  g00857(.A0(new_n3288_), .A1(new_n3118_), .B0(new_n3290_), .B1(new_n3225_), .Y(new_n3293_));
  OAI21X1  g00858(.A0(new_n3293_), .A1(new_n3222_), .B0(new_n3223_), .Y(new_n3294_));
  AOI21X1  g00859(.A0(new_n3292_), .A1(new_n3287_), .B0(new_n3294_), .Y(new_n3295_));
  OAI21X1  g00860(.A0(new_n3290_), .A1(new_n3223_), .B0(pi0239), .Y(new_n3296_));
  OAI22X1  g00861(.A0(new_n3296_), .A1(new_n3295_), .B0(new_n3230_), .B1(new_n3228_), .Y(po0154));
  AOI21X1  g00862(.A0(pi0833), .A1(new_n2438_), .B0(pi1145), .Y(new_n3298_));
  INVX1    g00863(.A(new_n3145_), .Y(new_n3299_));
  OAI21X1  g00864(.A0(new_n3299_), .A1(pi0927), .B0(pi0221), .Y(new_n3300_));
  NOR2X1   g00865(.A(new_n3300_), .B(new_n3298_), .Y(new_n3301_));
  AOI21X1  g00866(.A0(pi0274), .A1(pi0216), .B0(pi0221), .Y(new_n3302_));
  INVX1    g00867(.A(new_n3241_), .Y(new_n3303_));
  AOI21X1  g00868(.A0(new_n3245_), .A1(pi0151), .B0(pi0216), .Y(new_n3304_));
  OAI21X1  g00869(.A0(new_n3303_), .A1(pi0151), .B0(new_n3304_), .Y(new_n3305_));
  AOI21X1  g00870(.A0(new_n3305_), .A1(new_n3302_), .B0(new_n3301_), .Y(new_n3306_));
  AOI21X1  g00871(.A0(pi1145), .A1(pi0215), .B0(new_n2933_), .Y(new_n3307_));
  OAI21X1  g00872(.A0(new_n3306_), .A1(pi0215), .B0(new_n3307_), .Y(new_n3308_));
  INVX1    g00873(.A(pi1145), .Y(new_n3309_));
  INVX1    g00874(.A(new_n3134_), .Y(new_n3310_));
  OAI21X1  g00875(.A0(new_n3310_), .A1(pi0927), .B0(pi0222), .Y(new_n3311_));
  AOI21X1  g00876(.A0(new_n3310_), .A1(new_n3309_), .B0(new_n3311_), .Y(new_n3312_));
  INVX1    g00877(.A(pi0274), .Y(new_n3313_));
  OAI21X1  g00878(.A0(new_n3313_), .A1(new_n2942_), .B0(new_n2941_), .Y(new_n3314_));
  AOI21X1  g00879(.A0(new_n3232_), .A1(new_n2942_), .B0(new_n3314_), .Y(new_n3315_));
  OAI21X1  g00880(.A0(new_n3315_), .A1(new_n3312_), .B0(new_n2940_), .Y(new_n3316_));
  AOI21X1  g00881(.A0(pi1145), .A1(pi0223), .B0(pi0299), .Y(new_n3317_));
  AOI21X1  g00882(.A0(new_n3317_), .A1(new_n3316_), .B0(pi0039), .Y(new_n3318_));
  NAND2X1  g00883(.A(pi1145), .B(pi0223), .Y(new_n3319_));
  AND3X1   g00884(.A(new_n3313_), .B(pi0224), .C(new_n2941_), .Y(new_n3320_));
  OAI21X1  g00885(.A0(new_n3320_), .A1(new_n3312_), .B0(new_n2940_), .Y(new_n3321_));
  AOI21X1  g00886(.A0(new_n3321_), .A1(new_n3319_), .B0(pi0299), .Y(new_n3322_));
  NOR2X1   g00887(.A(new_n3322_), .B(new_n3262_), .Y(new_n3323_));
  INVX1    g00888(.A(new_n3323_), .Y(new_n3324_));
  AOI21X1  g00889(.A0(pi0228), .A1(pi0105), .B0(pi0151), .Y(new_n3325_));
  NOR2X1   g00890(.A(new_n3325_), .B(new_n3254_), .Y(new_n3326_));
  NOR4X1   g00891(.A(new_n2985_), .B(new_n2536_), .C(pi0228), .D(pi0151), .Y(new_n3327_));
  OAI21X1  g00892(.A0(new_n3327_), .A1(new_n3326_), .B0(new_n2438_), .Y(new_n3328_));
  AOI21X1  g00893(.A0(new_n3328_), .A1(new_n3302_), .B0(new_n3301_), .Y(new_n3329_));
  MX2X1    g00894(.A(new_n3329_), .B(new_n3309_), .S0(pi0215), .Y(new_n3330_));
  INVX1    g00895(.A(new_n3330_), .Y(new_n3331_));
  AOI21X1  g00896(.A0(new_n3331_), .A1(pi0299), .B0(new_n3324_), .Y(new_n3332_));
  OAI21X1  g00897(.A0(new_n3332_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n3333_));
  AOI21X1  g00898(.A0(new_n3318_), .A1(new_n3308_), .B0(new_n3333_), .Y(new_n3334_));
  OAI21X1  g00899(.A0(new_n3325_), .A1(pi0216), .B0(new_n3302_), .Y(new_n3335_));
  OAI21X1  g00900(.A0(new_n3300_), .A1(new_n3298_), .B0(new_n3335_), .Y(new_n3336_));
  MX2X1    g00901(.A(new_n3336_), .B(pi1145), .S0(pi0215), .Y(new_n3337_));
  INVX1    g00902(.A(new_n3337_), .Y(new_n3338_));
  AND2X1   g00903(.A(new_n3254_), .B(new_n3018_), .Y(new_n3339_));
  OAI21X1  g00904(.A0(new_n3313_), .A1(new_n2438_), .B0(new_n3339_), .Y(new_n3340_));
  AND2X1   g00905(.A(new_n3340_), .B(new_n3338_), .Y(new_n3341_));
  INVX1    g00906(.A(new_n3341_), .Y(new_n3342_));
  AOI21X1  g00907(.A0(new_n3342_), .A1(pi0299), .B0(new_n3324_), .Y(new_n3343_));
  INVX1    g00908(.A(new_n3343_), .Y(new_n3344_));
  OAI21X1  g00909(.A0(new_n3344_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3345_));
  INVX1    g00910(.A(new_n3302_), .Y(new_n3346_));
  INVX1    g00911(.A(pi0151), .Y(new_n3347_));
  INVX1    g00912(.A(new_n2454_), .Y(new_n3348_));
  AOI22X1  g00913(.A0(new_n3198_), .A1(new_n2793_), .B0(new_n3009_), .B1(new_n3348_), .Y(new_n3349_));
  AOI21X1  g00914(.A0(new_n3349_), .A1(new_n3347_), .B0(new_n3328_), .Y(new_n3350_));
  OAI22X1  g00915(.A0(new_n3350_), .A1(new_n3346_), .B0(new_n3300_), .B1(new_n3298_), .Y(new_n3351_));
  MX2X1    g00916(.A(new_n3351_), .B(pi1145), .S0(pi0215), .Y(new_n3352_));
  OR3X1    g00917(.A(new_n3322_), .B(new_n3262_), .C(new_n3060_), .Y(new_n3353_));
  AOI21X1  g00918(.A0(new_n3352_), .A1(pi0299), .B0(new_n3353_), .Y(new_n3354_));
  OAI21X1  g00919(.A0(new_n3344_), .A1(new_n3047_), .B0(pi0100), .Y(new_n3355_));
  OAI22X1  g00920(.A0(new_n3355_), .A1(new_n3354_), .B0(new_n3345_), .B1(new_n3334_), .Y(new_n3356_));
  MX2X1    g00921(.A(new_n3343_), .B(new_n3332_), .S0(new_n3064_), .Y(new_n3357_));
  OAI21X1  g00922(.A0(new_n3357_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n3358_));
  AOI21X1  g00923(.A0(new_n3356_), .A1(new_n3131_), .B0(new_n3358_), .Y(new_n3359_));
  OAI21X1  g00924(.A0(new_n3344_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3360_));
  NAND2X1  g00925(.A(new_n3357_), .B(new_n3077_), .Y(new_n3361_));
  AOI21X1  g00926(.A0(new_n3343_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n3362_));
  AOI21X1  g00927(.A0(new_n3362_), .A1(new_n3361_), .B0(new_n3130_), .Y(new_n3363_));
  OAI21X1  g00928(.A0(new_n3360_), .A1(new_n3359_), .B0(new_n3363_), .Y(new_n3364_));
  AOI21X1  g00929(.A0(new_n3343_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3365_));
  OAI21X1  g00930(.A0(new_n3342_), .A1(new_n3104_), .B0(pi0055), .Y(new_n3366_));
  AOI21X1  g00931(.A0(new_n3330_), .A1(new_n3104_), .B0(new_n3366_), .Y(new_n3367_));
  OR2X1    g00932(.A(new_n3367_), .B(pi0056), .Y(new_n3368_));
  AOI21X1  g00933(.A0(new_n3365_), .A1(new_n3364_), .B0(new_n3368_), .Y(new_n3369_));
  OAI21X1  g00934(.A0(new_n3341_), .A1(new_n3114_), .B0(pi0056), .Y(new_n3370_));
  AOI21X1  g00935(.A0(new_n3331_), .A1(new_n3114_), .B0(new_n3370_), .Y(new_n3371_));
  OR3X1    g00936(.A(new_n3371_), .B(new_n3369_), .C(pi0062), .Y(new_n3372_));
  INVX1    g00937(.A(pi0235), .Y(new_n3373_));
  INVX1    g00938(.A(new_n3223_), .Y(new_n3374_));
  OAI21X1  g00939(.A0(new_n3342_), .A1(new_n3224_), .B0(pi0062), .Y(new_n3375_));
  AOI21X1  g00940(.A0(new_n3330_), .A1(new_n3224_), .B0(new_n3375_), .Y(new_n3376_));
  NOR3X1   g00941(.A(new_n3376_), .B(new_n3374_), .C(new_n3373_), .Y(new_n3377_));
  INVX1    g00942(.A(new_n3111_), .Y(new_n3378_));
  OAI22X1  g00943(.A0(new_n3300_), .A1(new_n3298_), .B0(new_n3309_), .B1(new_n2934_), .Y(new_n3379_));
  NOR4X1   g00944(.A(new_n3379_), .B(new_n2986_), .C(pi0228), .D(pi0216), .Y(new_n3380_));
  AND2X1   g00945(.A(new_n3337_), .B(pi0299), .Y(new_n3381_));
  INVX1    g00946(.A(new_n3381_), .Y(new_n3382_));
  NOR2X1   g00947(.A(new_n3382_), .B(new_n3380_), .Y(new_n3383_));
  NOR3X1   g00948(.A(new_n3383_), .B(new_n3322_), .C(new_n3378_), .Y(new_n3384_));
  NOR3X1   g00949(.A(new_n3381_), .B(new_n3322_), .C(new_n3064_), .Y(new_n3385_));
  OAI21X1  g00950(.A0(new_n3385_), .A1(new_n3384_), .B0(pi0087), .Y(new_n3386_));
  INVX1    g00951(.A(new_n3181_), .Y(new_n3387_));
  AND2X1   g00952(.A(pi0100), .B(new_n2939_), .Y(new_n3388_));
  NAND2X1  g00953(.A(new_n3388_), .B(new_n3198_), .Y(new_n3389_));
  OAI21X1  g00954(.A0(new_n3387_), .A1(pi0100), .B0(new_n3389_), .Y(new_n3390_));
  NOR2X1   g00955(.A(new_n3379_), .B(new_n3200_), .Y(new_n3391_));
  AOI21X1  g00956(.A0(new_n3391_), .A1(new_n3390_), .B0(new_n3382_), .Y(new_n3392_));
  OR2X1    g00957(.A(new_n3322_), .B(pi0087), .Y(new_n3393_));
  OAI21X1  g00958(.A0(new_n3393_), .A1(new_n3392_), .B0(new_n3386_), .Y(new_n3394_));
  NOR2X1   g00959(.A(new_n3381_), .B(new_n3322_), .Y(new_n3395_));
  INVX1    g00960(.A(new_n3395_), .Y(new_n3396_));
  OAI21X1  g00961(.A0(new_n3396_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3397_));
  AOI21X1  g00962(.A0(new_n3394_), .A1(new_n3073_), .B0(new_n3397_), .Y(new_n3398_));
  NOR4X1   g00963(.A(new_n3383_), .B(new_n3322_), .C(new_n3378_), .D(new_n3080_), .Y(new_n3399_));
  OAI21X1  g00964(.A0(new_n3396_), .A1(new_n3208_), .B0(pi0092), .Y(new_n3400_));
  OAI21X1  g00965(.A0(new_n3400_), .A1(new_n3399_), .B0(new_n3102_), .Y(new_n3401_));
  AOI21X1  g00966(.A0(new_n3395_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3402_));
  OAI21X1  g00967(.A0(new_n3401_), .A1(new_n3398_), .B0(new_n3402_), .Y(new_n3403_));
  NAND2X1  g00968(.A(new_n3380_), .B(new_n3104_), .Y(new_n3404_));
  AND2X1   g00969(.A(new_n3337_), .B(pi0055), .Y(new_n3405_));
  AOI21X1  g00970(.A0(new_n3405_), .A1(new_n3404_), .B0(pi0056), .Y(new_n3406_));
  AOI21X1  g00971(.A0(new_n3380_), .A1(new_n3114_), .B0(new_n3338_), .Y(new_n3407_));
  OAI21X1  g00972(.A0(new_n3407_), .A1(new_n3118_), .B0(new_n3222_), .Y(new_n3408_));
  AOI21X1  g00973(.A0(new_n3406_), .A1(new_n3403_), .B0(new_n3408_), .Y(new_n3409_));
  AND3X1   g00974(.A(new_n3380_), .B(new_n3114_), .C(new_n3118_), .Y(new_n3410_));
  NAND2X1  g00975(.A(new_n3337_), .B(pi0062), .Y(new_n3411_));
  NOR3X1   g00976(.A(pi0235), .B(pi0059), .C(pi0057), .Y(new_n3412_));
  OAI21X1  g00977(.A0(new_n3411_), .A1(new_n3410_), .B0(new_n3412_), .Y(new_n3413_));
  OAI21X1  g00978(.A0(new_n3340_), .A1(new_n3373_), .B0(new_n3374_), .Y(new_n3414_));
  OAI22X1  g00979(.A0(new_n3414_), .A1(new_n3337_), .B0(new_n3413_), .B1(new_n3409_), .Y(new_n3415_));
  AOI21X1  g00980(.A0(new_n3377_), .A1(new_n3372_), .B0(new_n3415_), .Y(po0155));
  AND2X1   g00981(.A(pi1143), .B(pi0215), .Y(new_n3417_));
  NOR2X1   g00982(.A(new_n3417_), .B(new_n2933_), .Y(new_n3418_));
  INVX1    g00983(.A(pi0944), .Y(new_n3419_));
  AOI21X1  g00984(.A0(new_n3145_), .A1(new_n3419_), .B0(new_n2437_), .Y(new_n3420_));
  OAI21X1  g00985(.A0(new_n3145_), .A1(pi1143), .B0(new_n3420_), .Y(new_n3421_));
  AOI21X1  g00986(.A0(pi0264), .A1(pi0216), .B0(pi0221), .Y(new_n3422_));
  AOI21X1  g00987(.A0(new_n3244_), .A1(pi0146), .B0(pi0284), .Y(new_n3423_));
  AND3X1   g00988(.A(new_n3180_), .B(pi0284), .C(pi0146), .Y(new_n3424_));
  OAI22X1  g00989(.A0(new_n3424_), .A1(new_n3423_), .B0(new_n3240_), .B1(pi0146), .Y(new_n3425_));
  INVX1    g00990(.A(pi0284), .Y(new_n3426_));
  AOI21X1  g00991(.A0(new_n2453_), .A1(pi0095), .B0(new_n3426_), .Y(new_n3427_));
  AOI21X1  g00992(.A0(pi0146), .A1(new_n2447_), .B0(new_n2793_), .Y(new_n3428_));
  OAI21X1  g00993(.A0(new_n3427_), .A1(new_n2447_), .B0(new_n3428_), .Y(new_n3429_));
  OAI21X1  g00994(.A0(new_n3232_), .A1(new_n3011_), .B0(new_n3429_), .Y(new_n3430_));
  AOI21X1  g00995(.A0(new_n3425_), .A1(new_n2793_), .B0(new_n3430_), .Y(new_n3431_));
  OAI21X1  g00996(.A0(new_n3431_), .A1(pi0216), .B0(new_n3422_), .Y(new_n3432_));
  AND2X1   g00997(.A(new_n3432_), .B(new_n3421_), .Y(new_n3433_));
  OAI21X1  g00998(.A0(new_n3433_), .A1(pi0215), .B0(new_n3418_), .Y(new_n3434_));
  AOI21X1  g00999(.A0(pi1143), .A1(pi0223), .B0(pi0299), .Y(new_n3435_));
  AOI21X1  g01000(.A0(new_n3134_), .A1(new_n3419_), .B0(new_n2941_), .Y(new_n3436_));
  OAI21X1  g01001(.A0(new_n3134_), .A1(pi1143), .B0(new_n3436_), .Y(new_n3437_));
  AOI21X1  g01002(.A0(pi0264), .A1(pi0224), .B0(pi0222), .Y(new_n3438_));
  INVX1    g01003(.A(new_n3438_), .Y(new_n3439_));
  AOI21X1  g01004(.A0(new_n3232_), .A1(new_n3426_), .B0(pi0224), .Y(new_n3440_));
  OAI21X1  g01005(.A0(new_n3440_), .A1(new_n3439_), .B0(new_n3437_), .Y(new_n3441_));
  NOR2X1   g01006(.A(new_n3439_), .B(new_n3232_), .Y(new_n3442_));
  OAI21X1  g01007(.A0(new_n3442_), .A1(new_n3441_), .B0(new_n2940_), .Y(new_n3443_));
  AOI21X1  g01008(.A0(new_n3443_), .A1(new_n3435_), .B0(pi0039), .Y(new_n3444_));
  AND2X1   g01009(.A(pi1143), .B(pi0223), .Y(new_n3445_));
  OR3X1    g01010(.A(new_n3441_), .B(new_n3445_), .C(pi0299), .Y(new_n3446_));
  AND2X1   g01011(.A(new_n3446_), .B(new_n3444_), .Y(new_n3447_));
  AOI21X1  g01012(.A0(new_n3427_), .A1(new_n2942_), .B0(new_n3439_), .Y(new_n3448_));
  INVX1    g01013(.A(new_n3448_), .Y(new_n3449_));
  AOI21X1  g01014(.A0(new_n3449_), .A1(new_n3437_), .B0(pi0223), .Y(new_n3450_));
  OAI21X1  g01015(.A0(new_n3450_), .A1(new_n3445_), .B0(new_n2933_), .Y(new_n3451_));
  AOI21X1  g01016(.A0(new_n2990_), .A1(new_n2454_), .B0(new_n3451_), .Y(new_n3452_));
  INVX1    g01017(.A(new_n3421_), .Y(new_n3453_));
  INVX1    g01018(.A(new_n3422_), .Y(new_n3454_));
  MX2X1    g01019(.A(new_n3426_), .B(pi0146), .S0(new_n2986_), .Y(new_n3455_));
  INVX1    g01020(.A(new_n3254_), .Y(new_n3456_));
  AND2X1   g01021(.A(new_n3429_), .B(new_n3456_), .Y(new_n3457_));
  OAI21X1  g01022(.A0(new_n3455_), .A1(pi0228), .B0(new_n3457_), .Y(new_n3458_));
  AOI21X1  g01023(.A0(new_n3458_), .A1(new_n2438_), .B0(new_n3454_), .Y(new_n3459_));
  OR2X1    g01024(.A(new_n3459_), .B(new_n3453_), .Y(new_n3460_));
  AOI21X1  g01025(.A0(new_n3460_), .A1(new_n2934_), .B0(new_n3417_), .Y(new_n3461_));
  NOR2X1   g01026(.A(new_n3461_), .B(new_n2933_), .Y(new_n3462_));
  NOR2X1   g01027(.A(new_n3462_), .B(new_n3452_), .Y(new_n3463_));
  OAI21X1  g01028(.A0(new_n3463_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n3464_));
  AOI21X1  g01029(.A0(new_n3447_), .A1(new_n3434_), .B0(new_n3464_), .Y(new_n3465_));
  OR2X1    g01030(.A(pi0228), .B(pi0146), .Y(new_n3466_));
  AND3X1   g01031(.A(new_n3466_), .B(new_n3429_), .C(new_n3456_), .Y(new_n3467_));
  OAI21X1  g01032(.A0(new_n3467_), .A1(pi0216), .B0(new_n3422_), .Y(new_n3468_));
  AOI21X1  g01033(.A0(new_n3468_), .A1(new_n3421_), .B0(pi0215), .Y(new_n3469_));
  NOR2X1   g01034(.A(new_n3469_), .B(new_n3417_), .Y(new_n3470_));
  INVX1    g01035(.A(new_n3470_), .Y(new_n3471_));
  AOI21X1  g01036(.A0(new_n3471_), .A1(pi0299), .B0(new_n3452_), .Y(new_n3472_));
  INVX1    g01037(.A(new_n3472_), .Y(new_n3473_));
  OAI21X1  g01038(.A0(new_n3473_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3474_));
  AOI21X1  g01039(.A0(new_n2450_), .A1(pi0252), .B0(pi0284), .Y(new_n3475_));
  AOI21X1  g01040(.A0(new_n3475_), .A1(new_n2987_), .B0(pi0228), .Y(new_n3476_));
  OAI21X1  g01041(.A0(new_n3194_), .A1(new_n2776_), .B0(new_n3476_), .Y(new_n3477_));
  AOI21X1  g01042(.A0(new_n3477_), .A1(new_n3457_), .B0(pi0216), .Y(new_n3478_));
  OAI21X1  g01043(.A0(new_n3478_), .A1(new_n3454_), .B0(new_n3421_), .Y(new_n3479_));
  MX2X1    g01044(.A(new_n3479_), .B(pi1143), .S0(pi0215), .Y(new_n3480_));
  OR2X1    g01045(.A(new_n3452_), .B(new_n3060_), .Y(new_n3481_));
  AOI21X1  g01046(.A0(new_n3480_), .A1(pi0299), .B0(new_n3481_), .Y(new_n3482_));
  OAI21X1  g01047(.A0(new_n3473_), .A1(new_n3047_), .B0(pi0100), .Y(new_n3483_));
  OAI22X1  g01048(.A0(new_n3483_), .A1(new_n3482_), .B0(new_n3474_), .B1(new_n3465_), .Y(new_n3484_));
  MX2X1    g01049(.A(new_n3472_), .B(new_n3463_), .S0(new_n3064_), .Y(new_n3485_));
  OAI21X1  g01050(.A0(new_n3485_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n3486_));
  AOI21X1  g01051(.A0(new_n3484_), .A1(new_n3131_), .B0(new_n3486_), .Y(new_n3487_));
  OAI21X1  g01052(.A0(new_n3473_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3488_));
  NAND2X1  g01053(.A(new_n3485_), .B(new_n3077_), .Y(new_n3489_));
  AOI21X1  g01054(.A0(new_n3472_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n3490_));
  AOI21X1  g01055(.A0(new_n3490_), .A1(new_n3489_), .B0(new_n3130_), .Y(new_n3491_));
  OAI21X1  g01056(.A0(new_n3488_), .A1(new_n3487_), .B0(new_n3491_), .Y(new_n3492_));
  AOI21X1  g01057(.A0(new_n3472_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3493_));
  OAI21X1  g01058(.A0(new_n3471_), .A1(new_n3104_), .B0(pi0055), .Y(new_n3494_));
  AOI21X1  g01059(.A0(new_n3461_), .A1(new_n3104_), .B0(new_n3494_), .Y(new_n3495_));
  OR2X1    g01060(.A(new_n3495_), .B(pi0056), .Y(new_n3496_));
  AOI21X1  g01061(.A0(new_n3493_), .A1(new_n3492_), .B0(new_n3496_), .Y(new_n3497_));
  AOI21X1  g01062(.A0(new_n3471_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n3498_));
  OAI21X1  g01063(.A0(new_n3461_), .A1(new_n3115_), .B0(new_n3498_), .Y(new_n3499_));
  NAND2X1  g01064(.A(new_n3499_), .B(new_n3222_), .Y(new_n3500_));
  OAI21X1  g01065(.A0(new_n3471_), .A1(new_n3224_), .B0(pi0062), .Y(new_n3501_));
  AOI21X1  g01066(.A0(new_n3461_), .A1(new_n3224_), .B0(new_n3501_), .Y(new_n3502_));
  NOR3X1   g01067(.A(new_n3502_), .B(new_n3374_), .C(pi0238), .Y(new_n3503_));
  OAI21X1  g01068(.A0(new_n3500_), .A1(new_n3497_), .B0(new_n3503_), .Y(new_n3504_));
  NOR2X1   g01069(.A(new_n3429_), .B(new_n3243_), .Y(new_n3505_));
  AOI21X1  g01070(.A0(new_n3244_), .A1(new_n2776_), .B0(new_n3426_), .Y(new_n3506_));
  OAI21X1  g01071(.A0(new_n3240_), .A1(new_n2776_), .B0(new_n3506_), .Y(new_n3507_));
  NAND3X1  g01072(.A(new_n3180_), .B(new_n3426_), .C(new_n2776_), .Y(new_n3508_));
  AOI21X1  g01073(.A0(new_n3508_), .A1(new_n3507_), .B0(pi0228), .Y(new_n3509_));
  OAI21X1  g01074(.A0(new_n3509_), .A1(new_n3505_), .B0(new_n2438_), .Y(new_n3510_));
  AOI21X1  g01075(.A0(new_n3510_), .A1(new_n3422_), .B0(new_n3453_), .Y(new_n3511_));
  OAI21X1  g01076(.A0(new_n3511_), .A1(pi0215), .B0(new_n3418_), .Y(new_n3512_));
  NOR2X1   g01077(.A(new_n3450_), .B(new_n3445_), .Y(new_n3513_));
  OAI21X1  g01078(.A0(new_n3455_), .A1(pi0228), .B0(new_n3429_), .Y(new_n3514_));
  AOI21X1  g01079(.A0(new_n3514_), .A1(new_n2438_), .B0(new_n3454_), .Y(new_n3515_));
  OR2X1    g01080(.A(new_n3515_), .B(new_n3453_), .Y(new_n3516_));
  AOI21X1  g01081(.A0(new_n3516_), .A1(new_n2934_), .B0(new_n3417_), .Y(new_n3517_));
  MX2X1    g01082(.A(new_n3517_), .B(new_n3513_), .S0(new_n2933_), .Y(new_n3518_));
  OAI21X1  g01083(.A0(new_n3518_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n3519_));
  AOI21X1  g01084(.A0(new_n3512_), .A1(new_n3444_), .B0(new_n3519_), .Y(new_n3520_));
  INVX1    g01085(.A(pi0264), .Y(new_n3521_));
  OAI21X1  g01086(.A0(new_n3521_), .A1(new_n2438_), .B0(new_n3339_), .Y(new_n3522_));
  AND2X1   g01087(.A(new_n3522_), .B(new_n3470_), .Y(new_n3523_));
  MX2X1    g01088(.A(new_n3523_), .B(new_n3513_), .S0(new_n2933_), .Y(new_n3524_));
  INVX1    g01089(.A(new_n3524_), .Y(new_n3525_));
  OAI21X1  g01090(.A0(new_n3525_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3526_));
  AOI21X1  g01091(.A0(new_n3477_), .A1(new_n3429_), .B0(pi0216), .Y(new_n3527_));
  OAI21X1  g01092(.A0(new_n3527_), .A1(new_n3454_), .B0(new_n3421_), .Y(new_n3528_));
  MX2X1    g01093(.A(new_n3528_), .B(pi1143), .S0(pi0215), .Y(new_n3529_));
  NAND2X1  g01094(.A(new_n3451_), .B(new_n3047_), .Y(new_n3530_));
  AOI21X1  g01095(.A0(new_n3529_), .A1(pi0299), .B0(new_n3530_), .Y(new_n3531_));
  OAI21X1  g01096(.A0(new_n3525_), .A1(new_n3047_), .B0(pi0100), .Y(new_n3532_));
  OAI22X1  g01097(.A0(new_n3532_), .A1(new_n3531_), .B0(new_n3526_), .B1(new_n3520_), .Y(new_n3533_));
  MX2X1    g01098(.A(new_n3524_), .B(new_n3518_), .S0(new_n3064_), .Y(new_n3534_));
  OAI21X1  g01099(.A0(new_n3534_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n3535_));
  AOI21X1  g01100(.A0(new_n3533_), .A1(new_n3131_), .B0(new_n3535_), .Y(new_n3536_));
  OAI21X1  g01101(.A0(new_n3525_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3537_));
  NAND2X1  g01102(.A(new_n3534_), .B(new_n3077_), .Y(new_n3538_));
  AOI21X1  g01103(.A0(new_n3524_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n3539_));
  AOI21X1  g01104(.A0(new_n3539_), .A1(new_n3538_), .B0(new_n3130_), .Y(new_n3540_));
  OAI21X1  g01105(.A0(new_n3537_), .A1(new_n3536_), .B0(new_n3540_), .Y(new_n3541_));
  AOI21X1  g01106(.A0(new_n3524_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3542_));
  INVX1    g01107(.A(new_n3523_), .Y(new_n3543_));
  OAI21X1  g01108(.A0(new_n3543_), .A1(new_n3104_), .B0(pi0055), .Y(new_n3544_));
  AOI21X1  g01109(.A0(new_n3517_), .A1(new_n3104_), .B0(new_n3544_), .Y(new_n3545_));
  OR2X1    g01110(.A(new_n3545_), .B(pi0056), .Y(new_n3546_));
  AOI21X1  g01111(.A0(new_n3542_), .A1(new_n3541_), .B0(new_n3546_), .Y(new_n3547_));
  AOI21X1  g01112(.A0(new_n3543_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n3548_));
  OAI21X1  g01113(.A0(new_n3517_), .A1(new_n3115_), .B0(new_n3548_), .Y(new_n3549_));
  NAND2X1  g01114(.A(new_n3549_), .B(new_n3222_), .Y(new_n3550_));
  INVX1    g01115(.A(pi0238), .Y(new_n3551_));
  OAI21X1  g01116(.A0(new_n3543_), .A1(new_n3224_), .B0(pi0062), .Y(new_n3552_));
  AOI21X1  g01117(.A0(new_n3517_), .A1(new_n3224_), .B0(new_n3552_), .Y(new_n3553_));
  NOR3X1   g01118(.A(new_n3553_), .B(new_n3374_), .C(new_n3551_), .Y(new_n3554_));
  OAI21X1  g01119(.A0(new_n3550_), .A1(new_n3547_), .B0(new_n3554_), .Y(new_n3555_));
  OAI21X1  g01120(.A0(new_n3522_), .A1(new_n3551_), .B0(new_n3374_), .Y(new_n3556_));
  OR3X1    g01121(.A(new_n3556_), .B(new_n3469_), .C(new_n3417_), .Y(new_n3557_));
  AND3X1   g01122(.A(new_n3557_), .B(new_n3555_), .C(new_n3504_), .Y(po0156));
  AND2X1   g01123(.A(pi1142), .B(pi0215), .Y(new_n3559_));
  OR2X1    g01124(.A(new_n3559_), .B(new_n2933_), .Y(new_n3560_));
  INVX1    g01125(.A(pi0932), .Y(new_n3561_));
  AOI21X1  g01126(.A0(new_n3145_), .A1(new_n3561_), .B0(new_n2437_), .Y(new_n3562_));
  OAI21X1  g01127(.A0(new_n3145_), .A1(pi1142), .B0(new_n3562_), .Y(new_n3563_));
  AOI21X1  g01128(.A0(pi0277), .A1(pi0216), .B0(pi0221), .Y(new_n3564_));
  INVX1    g01129(.A(new_n3564_), .Y(new_n3565_));
  INVX1    g01130(.A(pi0262), .Y(new_n3566_));
  AOI21X1  g01131(.A0(new_n3244_), .A1(new_n3566_), .B0(pi0172), .Y(new_n3567_));
  AND3X1   g01132(.A(new_n3240_), .B(new_n3566_), .C(pi0172), .Y(new_n3568_));
  OR2X1    g01133(.A(new_n3568_), .B(new_n3567_), .Y(new_n3569_));
  INVX1    g01134(.A(new_n3180_), .Y(new_n3570_));
  AOI21X1  g01135(.A0(new_n3570_), .A1(pi0262), .B0(pi0228), .Y(new_n3571_));
  AOI21X1  g01136(.A0(new_n2453_), .A1(pi0095), .B0(new_n3566_), .Y(new_n3572_));
  AND2X1   g01137(.A(new_n3572_), .B(pi0105), .Y(new_n3573_));
  INVX1    g01138(.A(new_n3573_), .Y(new_n3574_));
  AOI21X1  g01139(.A0(pi0172), .A1(new_n2447_), .B0(new_n2793_), .Y(new_n3575_));
  OAI21X1  g01140(.A0(new_n3574_), .A1(new_n3231_), .B0(new_n3575_), .Y(new_n3576_));
  OAI21X1  g01141(.A0(new_n3576_), .A1(new_n3243_), .B0(new_n2438_), .Y(new_n3577_));
  AOI21X1  g01142(.A0(new_n3571_), .A1(new_n3569_), .B0(new_n3577_), .Y(new_n3578_));
  OAI21X1  g01143(.A0(new_n3578_), .A1(new_n3565_), .B0(new_n3563_), .Y(new_n3579_));
  AOI21X1  g01144(.A0(new_n3579_), .A1(new_n2934_), .B0(new_n3560_), .Y(new_n3580_));
  AOI21X1  g01145(.A0(pi1142), .A1(pi0223), .B0(pi0299), .Y(new_n3581_));
  AOI21X1  g01146(.A0(new_n3134_), .A1(new_n3561_), .B0(new_n2941_), .Y(new_n3582_));
  OAI21X1  g01147(.A0(new_n3134_), .A1(pi1142), .B0(new_n3582_), .Y(new_n3583_));
  AOI21X1  g01148(.A0(pi0277), .A1(pi0224), .B0(pi0222), .Y(new_n3584_));
  NOR3X1   g01149(.A(new_n3231_), .B(new_n2454_), .C(pi0262), .Y(new_n3585_));
  OAI21X1  g01150(.A0(new_n3585_), .A1(pi0224), .B0(new_n3584_), .Y(new_n3586_));
  AND3X1   g01151(.A(new_n3586_), .B(new_n3583_), .C(new_n3581_), .Y(new_n3587_));
  INVX1    g01152(.A(new_n3581_), .Y(new_n3588_));
  OAI21X1  g01153(.A0(new_n3231_), .A1(new_n2454_), .B0(new_n3584_), .Y(new_n3589_));
  NAND3X1  g01154(.A(new_n3589_), .B(new_n3586_), .C(new_n3583_), .Y(new_n3590_));
  AOI21X1  g01155(.A0(new_n3590_), .A1(new_n2940_), .B0(new_n3588_), .Y(new_n3591_));
  OR2X1    g01156(.A(new_n3591_), .B(pi0039), .Y(new_n3592_));
  OR3X1    g01157(.A(new_n3592_), .B(new_n3587_), .C(new_n3580_), .Y(new_n3593_));
  NAND3X1  g01158(.A(new_n2990_), .B(new_n2453_), .C(pi0095), .Y(new_n3594_));
  AND2X1   g01159(.A(pi1142), .B(pi0223), .Y(new_n3595_));
  INVX1    g01160(.A(new_n3595_), .Y(new_n3596_));
  INVX1    g01161(.A(new_n3583_), .Y(new_n3597_));
  INVX1    g01162(.A(new_n3584_), .Y(new_n3598_));
  AOI21X1  g01163(.A0(new_n3572_), .A1(new_n2942_), .B0(new_n3598_), .Y(new_n3599_));
  OAI21X1  g01164(.A0(new_n3599_), .A1(new_n3597_), .B0(new_n2940_), .Y(new_n3600_));
  AOI21X1  g01165(.A0(new_n3600_), .A1(new_n3596_), .B0(pi0299), .Y(new_n3601_));
  AND2X1   g01166(.A(new_n3601_), .B(new_n3594_), .Y(new_n3602_));
  NOR3X1   g01167(.A(new_n2985_), .B(new_n2536_), .C(pi0228), .Y(new_n3603_));
  INVX1    g01168(.A(new_n3603_), .Y(new_n3604_));
  AND2X1   g01169(.A(new_n2793_), .B(pi0172), .Y(new_n3605_));
  INVX1    g01170(.A(new_n3605_), .Y(new_n3606_));
  AOI22X1  g01171(.A0(new_n3606_), .A1(new_n3604_), .B0(new_n2987_), .B1(new_n3566_), .Y(new_n3607_));
  INVX1    g01172(.A(new_n3607_), .Y(new_n3608_));
  AND2X1   g01173(.A(pi0172), .B(new_n2447_), .Y(new_n3609_));
  OAI21X1  g01174(.A0(new_n3609_), .A1(new_n3573_), .B0(pi0228), .Y(new_n3610_));
  AND2X1   g01175(.A(new_n3610_), .B(new_n3456_), .Y(new_n3611_));
  AOI21X1  g01176(.A0(new_n3611_), .A1(new_n3608_), .B0(pi0216), .Y(new_n3612_));
  OAI21X1  g01177(.A0(new_n3612_), .A1(new_n3565_), .B0(new_n3563_), .Y(new_n3613_));
  AOI21X1  g01178(.A0(new_n3613_), .A1(new_n2934_), .B0(new_n3559_), .Y(new_n3614_));
  INVX1    g01179(.A(new_n3614_), .Y(new_n3615_));
  AOI21X1  g01180(.A0(new_n3615_), .A1(pi0299), .B0(new_n3602_), .Y(new_n3616_));
  INVX1    g01181(.A(new_n3616_), .Y(new_n3617_));
  AOI21X1  g01182(.A0(new_n3617_), .A1(pi0039), .B0(pi0038), .Y(new_n3618_));
  AOI21X1  g01183(.A0(new_n3610_), .A1(new_n3606_), .B0(pi0216), .Y(new_n3619_));
  OAI21X1  g01184(.A0(new_n3619_), .A1(new_n3565_), .B0(new_n3563_), .Y(new_n3620_));
  AOI21X1  g01185(.A0(new_n3620_), .A1(new_n2934_), .B0(new_n3559_), .Y(new_n3621_));
  NOR3X1   g01186(.A(new_n3621_), .B(new_n3255_), .C(new_n2933_), .Y(new_n3622_));
  NOR2X1   g01187(.A(new_n3622_), .B(new_n3602_), .Y(new_n3623_));
  INVX1    g01188(.A(new_n3623_), .Y(new_n3624_));
  OAI21X1  g01189(.A0(new_n3624_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3625_));
  AOI21X1  g01190(.A0(new_n3618_), .A1(new_n3593_), .B0(new_n3625_), .Y(new_n3626_));
  AND2X1   g01191(.A(new_n3198_), .B(new_n2793_), .Y(new_n3627_));
  OAI22X1  g01192(.A0(new_n3605_), .A1(new_n3627_), .B0(new_n3199_), .B1(pi0262), .Y(new_n3628_));
  AOI21X1  g01193(.A0(new_n3628_), .A1(new_n3611_), .B0(pi0216), .Y(new_n3629_));
  OAI21X1  g01194(.A0(new_n3629_), .A1(new_n3565_), .B0(new_n3563_), .Y(new_n3630_));
  AOI21X1  g01195(.A0(new_n3630_), .A1(new_n2934_), .B0(new_n3559_), .Y(new_n3631_));
  AOI21X1  g01196(.A0(new_n3601_), .A1(new_n3594_), .B0(new_n3060_), .Y(new_n3632_));
  OAI21X1  g01197(.A0(new_n3631_), .A1(new_n2933_), .B0(new_n3632_), .Y(new_n3633_));
  AOI21X1  g01198(.A0(new_n3623_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n3634_));
  AND2X1   g01199(.A(new_n3634_), .B(new_n3633_), .Y(new_n3635_));
  OAI21X1  g01200(.A0(new_n3635_), .A1(new_n3626_), .B0(new_n3131_), .Y(new_n3636_));
  MX2X1    g01201(.A(new_n3624_), .B(new_n3617_), .S0(new_n3064_), .Y(new_n3637_));
  AOI21X1  g01202(.A0(new_n3637_), .A1(pi0087), .B0(pi0075), .Y(new_n3638_));
  OAI21X1  g01203(.A0(new_n3624_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3639_));
  AOI21X1  g01204(.A0(new_n3638_), .A1(new_n3636_), .B0(new_n3639_), .Y(new_n3640_));
  NOR2X1   g01205(.A(new_n3637_), .B(new_n3080_), .Y(new_n3641_));
  OAI21X1  g01206(.A0(new_n3624_), .A1(new_n3077_), .B0(pi0092), .Y(new_n3642_));
  OAI21X1  g01207(.A0(new_n3642_), .A1(new_n3641_), .B0(new_n3102_), .Y(new_n3643_));
  AOI21X1  g01208(.A0(new_n3623_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3644_));
  OAI21X1  g01209(.A0(new_n3643_), .A1(new_n3640_), .B0(new_n3644_), .Y(new_n3645_));
  NAND2X1  g01210(.A(new_n3614_), .B(new_n3104_), .Y(new_n3646_));
  NOR2X1   g01211(.A(new_n3621_), .B(new_n3255_), .Y(new_n3647_));
  INVX1    g01212(.A(new_n3647_), .Y(new_n3648_));
  AOI21X1  g01213(.A0(new_n3648_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n3649_));
  AOI21X1  g01214(.A0(new_n3649_), .A1(new_n3646_), .B0(pi0056), .Y(new_n3650_));
  AOI21X1  g01215(.A0(new_n3647_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n3651_));
  OAI21X1  g01216(.A0(new_n3614_), .A1(new_n3115_), .B0(new_n3651_), .Y(new_n3652_));
  NAND2X1  g01217(.A(new_n3652_), .B(new_n3222_), .Y(new_n3653_));
  AOI21X1  g01218(.A0(new_n3650_), .A1(new_n3645_), .B0(new_n3653_), .Y(new_n3654_));
  OAI21X1  g01219(.A0(new_n3647_), .A1(new_n3224_), .B0(pi0062), .Y(new_n3655_));
  AOI21X1  g01220(.A0(new_n3614_), .A1(new_n3224_), .B0(new_n3655_), .Y(new_n3656_));
  OR2X1    g01221(.A(new_n3656_), .B(new_n3374_), .Y(new_n3657_));
  AOI21X1  g01222(.A0(new_n3648_), .A1(new_n3374_), .B0(pi0249), .Y(new_n3658_));
  OAI21X1  g01223(.A0(new_n3657_), .A1(new_n3654_), .B0(new_n3658_), .Y(new_n3659_));
  AOI21X1  g01224(.A0(new_n3240_), .A1(pi0262), .B0(pi0172), .Y(new_n3660_));
  OAI21X1  g01225(.A0(new_n3244_), .A1(new_n3566_), .B0(pi0172), .Y(new_n3661_));
  AOI21X1  g01226(.A0(new_n3180_), .A1(new_n3566_), .B0(new_n3661_), .Y(new_n3662_));
  OAI21X1  g01227(.A0(new_n3662_), .A1(new_n3660_), .B0(new_n2793_), .Y(new_n3663_));
  AND3X1   g01228(.A(new_n3663_), .B(new_n3576_), .C(new_n2438_), .Y(new_n3664_));
  OAI21X1  g01229(.A0(new_n3664_), .A1(new_n3565_), .B0(new_n3563_), .Y(new_n3665_));
  AOI21X1  g01230(.A0(new_n3665_), .A1(new_n2934_), .B0(new_n3560_), .Y(new_n3666_));
  AND2X1   g01231(.A(new_n3600_), .B(new_n3596_), .Y(new_n3667_));
  AOI21X1  g01232(.A0(new_n3610_), .A1(new_n3608_), .B0(pi0216), .Y(new_n3668_));
  OAI21X1  g01233(.A0(new_n3668_), .A1(new_n3565_), .B0(new_n3563_), .Y(new_n3669_));
  AOI21X1  g01234(.A0(new_n3669_), .A1(new_n2934_), .B0(new_n3559_), .Y(new_n3670_));
  MX2X1    g01235(.A(new_n3670_), .B(new_n3667_), .S0(new_n2933_), .Y(new_n3671_));
  INVX1    g01236(.A(new_n3671_), .Y(new_n3672_));
  AOI21X1  g01237(.A0(new_n3672_), .A1(pi0039), .B0(pi0038), .Y(new_n3673_));
  OAI21X1  g01238(.A0(new_n3666_), .A1(new_n3592_), .B0(new_n3673_), .Y(new_n3674_));
  MX2X1    g01239(.A(new_n3621_), .B(new_n3667_), .S0(new_n2933_), .Y(new_n3675_));
  AOI21X1  g01240(.A0(new_n3675_), .A1(pi0038), .B0(pi0100), .Y(new_n3676_));
  AOI21X1  g01241(.A0(new_n3628_), .A1(new_n3610_), .B0(pi0216), .Y(new_n3677_));
  OAI21X1  g01242(.A0(new_n3677_), .A1(new_n3565_), .B0(new_n3563_), .Y(new_n3678_));
  AOI21X1  g01243(.A0(new_n3678_), .A1(new_n2934_), .B0(new_n3559_), .Y(new_n3679_));
  NOR2X1   g01244(.A(new_n3601_), .B(new_n3060_), .Y(new_n3680_));
  OAI21X1  g01245(.A0(new_n3679_), .A1(new_n2933_), .B0(new_n3680_), .Y(new_n3681_));
  AOI21X1  g01246(.A0(new_n3675_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n3682_));
  AOI22X1  g01247(.A0(new_n3682_), .A1(new_n3681_), .B0(new_n3676_), .B1(new_n3674_), .Y(new_n3683_));
  INVX1    g01248(.A(new_n3675_), .Y(new_n3684_));
  MX2X1    g01249(.A(new_n3684_), .B(new_n3672_), .S0(new_n3064_), .Y(new_n3685_));
  AOI21X1  g01250(.A0(new_n3685_), .A1(pi0087), .B0(pi0075), .Y(new_n3686_));
  OAI21X1  g01251(.A0(new_n3683_), .A1(pi0087), .B0(new_n3686_), .Y(new_n3687_));
  AOI21X1  g01252(.A0(new_n3675_), .A1(pi0075), .B0(pi0092), .Y(new_n3688_));
  NOR2X1   g01253(.A(new_n3685_), .B(new_n3080_), .Y(new_n3689_));
  OAI21X1  g01254(.A0(new_n3684_), .A1(new_n3077_), .B0(pi0092), .Y(new_n3690_));
  OAI21X1  g01255(.A0(new_n3690_), .A1(new_n3689_), .B0(new_n3102_), .Y(new_n3691_));
  AOI21X1  g01256(.A0(new_n3688_), .A1(new_n3687_), .B0(new_n3691_), .Y(new_n3692_));
  OAI21X1  g01257(.A0(new_n3684_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n3693_));
  NAND2X1  g01258(.A(new_n3670_), .B(new_n3104_), .Y(new_n3694_));
  AOI21X1  g01259(.A0(new_n3621_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n3695_));
  AOI21X1  g01260(.A0(new_n3695_), .A1(new_n3694_), .B0(pi0056), .Y(new_n3696_));
  OAI21X1  g01261(.A0(new_n3693_), .A1(new_n3692_), .B0(new_n3696_), .Y(new_n3697_));
  INVX1    g01262(.A(new_n3621_), .Y(new_n3698_));
  AOI21X1  g01263(.A0(new_n3698_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n3699_));
  OAI21X1  g01264(.A0(new_n3670_), .A1(new_n3115_), .B0(new_n3699_), .Y(new_n3700_));
  AND2X1   g01265(.A(new_n3700_), .B(new_n3222_), .Y(new_n3701_));
  OAI21X1  g01266(.A0(new_n3698_), .A1(new_n3224_), .B0(pi0062), .Y(new_n3702_));
  AOI21X1  g01267(.A0(new_n3670_), .A1(new_n3224_), .B0(new_n3702_), .Y(new_n3703_));
  OR2X1    g01268(.A(new_n3703_), .B(new_n3374_), .Y(new_n3704_));
  AOI21X1  g01269(.A0(new_n3701_), .A1(new_n3697_), .B0(new_n3704_), .Y(new_n3705_));
  OAI21X1  g01270(.A0(new_n3698_), .A1(new_n3223_), .B0(pi0249), .Y(new_n3706_));
  OAI21X1  g01271(.A0(new_n3706_), .A1(new_n3705_), .B0(new_n3659_), .Y(po0157));
  AND2X1   g01272(.A(pi1141), .B(pi0215), .Y(new_n3708_));
  NOR2X1   g01273(.A(new_n3708_), .B(new_n2933_), .Y(new_n3709_));
  INVX1    g01274(.A(pi0935), .Y(new_n3710_));
  AOI21X1  g01275(.A0(new_n3145_), .A1(new_n3710_), .B0(new_n2437_), .Y(new_n3711_));
  OAI21X1  g01276(.A0(new_n3145_), .A1(pi1141), .B0(new_n3711_), .Y(new_n3712_));
  INVX1    g01277(.A(new_n3712_), .Y(new_n3713_));
  AOI21X1  g01278(.A0(pi0270), .A1(pi0216), .B0(pi0221), .Y(new_n3714_));
  INVX1    g01279(.A(pi0171), .Y(new_n3715_));
  INVX1    g01280(.A(pi0861), .Y(new_n3716_));
  OR3X1    g01281(.A(new_n3232_), .B(new_n2696_), .C(new_n3716_), .Y(new_n3717_));
  AND2X1   g01282(.A(new_n3717_), .B(new_n3715_), .Y(new_n3718_));
  MX2X1    g01283(.A(new_n3717_), .B(new_n3240_), .S0(pi0171), .Y(new_n3719_));
  AOI22X1  g01284(.A0(new_n3719_), .A1(pi0861), .B0(new_n3718_), .B1(new_n3180_), .Y(new_n3720_));
  INVX1    g01285(.A(new_n3243_), .Y(new_n3721_));
  AOI21X1  g01286(.A0(new_n2453_), .A1(pi0095), .B0(new_n3716_), .Y(new_n3722_));
  INVX1    g01287(.A(new_n3722_), .Y(new_n3723_));
  OAI21X1  g01288(.A0(new_n3715_), .A1(pi0105), .B0(pi0228), .Y(new_n3724_));
  AOI21X1  g01289(.A0(new_n3723_), .A1(pi0105), .B0(new_n3724_), .Y(new_n3725_));
  AOI21X1  g01290(.A0(new_n3725_), .A1(new_n3721_), .B0(pi0216), .Y(new_n3726_));
  OAI21X1  g01291(.A0(new_n3720_), .A1(pi0228), .B0(new_n3726_), .Y(new_n3727_));
  AOI21X1  g01292(.A0(new_n3727_), .A1(new_n3714_), .B0(new_n3713_), .Y(new_n3728_));
  OAI21X1  g01293(.A0(new_n3728_), .A1(pi0215), .B0(new_n3709_), .Y(new_n3729_));
  AND2X1   g01294(.A(pi1141), .B(pi0223), .Y(new_n3730_));
  AOI21X1  g01295(.A0(new_n3134_), .A1(new_n3710_), .B0(new_n2941_), .Y(new_n3731_));
  OAI21X1  g01296(.A0(new_n3134_), .A1(pi1141), .B0(new_n3731_), .Y(new_n3732_));
  AOI21X1  g01297(.A0(pi0270), .A1(pi0224), .B0(pi0222), .Y(new_n3733_));
  INVX1    g01298(.A(new_n3733_), .Y(new_n3734_));
  AOI21X1  g01299(.A0(new_n3232_), .A1(pi0861), .B0(pi0224), .Y(new_n3735_));
  OAI21X1  g01300(.A0(new_n3735_), .A1(new_n3734_), .B0(new_n3732_), .Y(new_n3736_));
  OR3X1    g01301(.A(new_n3736_), .B(new_n3730_), .C(pi0299), .Y(new_n3737_));
  AOI21X1  g01302(.A0(pi1141), .A1(pi0223), .B0(pi0299), .Y(new_n3738_));
  NOR2X1   g01303(.A(new_n3734_), .B(new_n3232_), .Y(new_n3739_));
  OAI21X1  g01304(.A0(new_n3739_), .A1(new_n3736_), .B0(new_n2940_), .Y(new_n3740_));
  AOI21X1  g01305(.A0(new_n3740_), .A1(new_n3738_), .B0(pi0039), .Y(new_n3741_));
  AND2X1   g01306(.A(new_n3741_), .B(new_n3737_), .Y(new_n3742_));
  AOI21X1  g01307(.A0(new_n3723_), .A1(new_n2942_), .B0(new_n3734_), .Y(new_n3743_));
  INVX1    g01308(.A(new_n3743_), .Y(new_n3744_));
  AOI21X1  g01309(.A0(new_n3744_), .A1(new_n3732_), .B0(pi0223), .Y(new_n3745_));
  OAI21X1  g01310(.A0(new_n3745_), .A1(new_n3730_), .B0(new_n2933_), .Y(new_n3746_));
  INVX1    g01311(.A(new_n3746_), .Y(new_n3747_));
  INVX1    g01312(.A(new_n3708_), .Y(new_n3748_));
  INVX1    g01313(.A(new_n3714_), .Y(new_n3749_));
  NOR2X1   g01314(.A(new_n3725_), .B(pi0216), .Y(new_n3750_));
  AOI21X1  g01315(.A0(new_n2986_), .A1(pi0171), .B0(pi0228), .Y(new_n3751_));
  OAI21X1  g01316(.A0(new_n2986_), .A1(pi0861), .B0(new_n3751_), .Y(new_n3752_));
  AOI21X1  g01317(.A0(new_n3752_), .A1(new_n3750_), .B0(new_n3749_), .Y(new_n3753_));
  OAI21X1  g01318(.A0(new_n3753_), .A1(new_n3713_), .B0(new_n2934_), .Y(new_n3754_));
  AOI21X1  g01319(.A0(new_n3754_), .A1(new_n3748_), .B0(new_n2933_), .Y(new_n3755_));
  NOR2X1   g01320(.A(new_n3755_), .B(new_n3747_), .Y(new_n3756_));
  OAI21X1  g01321(.A0(new_n3756_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n3757_));
  AOI21X1  g01322(.A0(new_n3742_), .A1(new_n3729_), .B0(new_n3757_), .Y(new_n3758_));
  INVX1    g01323(.A(pi1141), .Y(new_n3759_));
  OAI21X1  g01324(.A0(pi0228), .A1(pi0171), .B0(new_n3750_), .Y(new_n3760_));
  AOI21X1  g01325(.A0(new_n3760_), .A1(new_n3714_), .B0(new_n3713_), .Y(new_n3761_));
  MX2X1    g01326(.A(new_n3761_), .B(new_n3759_), .S0(pi0215), .Y(new_n3762_));
  INVX1    g01327(.A(new_n3762_), .Y(new_n3763_));
  AOI21X1  g01328(.A0(new_n3763_), .A1(pi0299), .B0(new_n3747_), .Y(new_n3764_));
  INVX1    g01329(.A(new_n3764_), .Y(new_n3765_));
  OAI21X1  g01330(.A0(new_n3765_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3766_));
  AOI21X1  g01331(.A0(new_n3199_), .A1(pi0171), .B0(pi0228), .Y(new_n3767_));
  OAI21X1  g01332(.A0(new_n3199_), .A1(pi0861), .B0(new_n3767_), .Y(new_n3768_));
  AOI21X1  g01333(.A0(new_n3768_), .A1(new_n3750_), .B0(new_n3749_), .Y(new_n3769_));
  OAI21X1  g01334(.A0(new_n3769_), .A1(new_n3713_), .B0(new_n2934_), .Y(new_n3770_));
  AOI21X1  g01335(.A0(new_n3770_), .A1(new_n3748_), .B0(new_n2933_), .Y(new_n3771_));
  NOR3X1   g01336(.A(new_n3771_), .B(new_n3747_), .C(new_n3060_), .Y(new_n3772_));
  OAI21X1  g01337(.A0(new_n3765_), .A1(new_n3047_), .B0(pi0100), .Y(new_n3773_));
  OAI22X1  g01338(.A0(new_n3773_), .A1(new_n3772_), .B0(new_n3766_), .B1(new_n3758_), .Y(new_n3774_));
  MX2X1    g01339(.A(new_n3764_), .B(new_n3756_), .S0(new_n3064_), .Y(new_n3775_));
  OAI21X1  g01340(.A0(new_n3775_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n3776_));
  AOI21X1  g01341(.A0(new_n3774_), .A1(new_n3131_), .B0(new_n3776_), .Y(new_n3777_));
  OAI21X1  g01342(.A0(new_n3765_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3778_));
  NAND2X1  g01343(.A(new_n3775_), .B(new_n3077_), .Y(new_n3779_));
  AOI21X1  g01344(.A0(new_n3764_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n3780_));
  AOI21X1  g01345(.A0(new_n3780_), .A1(new_n3779_), .B0(new_n3130_), .Y(new_n3781_));
  OAI21X1  g01346(.A0(new_n3778_), .A1(new_n3777_), .B0(new_n3781_), .Y(new_n3782_));
  AOI21X1  g01347(.A0(new_n3764_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3783_));
  AND3X1   g01348(.A(new_n3754_), .B(new_n3748_), .C(new_n3104_), .Y(new_n3784_));
  OAI21X1  g01349(.A0(new_n3763_), .A1(new_n3104_), .B0(pi0055), .Y(new_n3785_));
  OAI21X1  g01350(.A0(new_n3785_), .A1(new_n3784_), .B0(new_n3118_), .Y(new_n3786_));
  AOI21X1  g01351(.A0(new_n3783_), .A1(new_n3782_), .B0(new_n3786_), .Y(new_n3787_));
  AOI21X1  g01352(.A0(new_n3754_), .A1(new_n3748_), .B0(new_n3115_), .Y(new_n3788_));
  OAI21X1  g01353(.A0(new_n3762_), .A1(new_n3114_), .B0(pi0056), .Y(new_n3789_));
  OAI21X1  g01354(.A0(new_n3789_), .A1(new_n3788_), .B0(new_n3222_), .Y(new_n3790_));
  NAND3X1  g01355(.A(new_n3754_), .B(new_n3748_), .C(new_n3224_), .Y(new_n3791_));
  AOI21X1  g01356(.A0(new_n3762_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n3792_));
  OR3X1    g01357(.A(pi0241), .B(pi0059), .C(pi0057), .Y(new_n3793_));
  AOI21X1  g01358(.A0(new_n3792_), .A1(new_n3791_), .B0(new_n3793_), .Y(new_n3794_));
  OAI21X1  g01359(.A0(new_n3790_), .A1(new_n3787_), .B0(new_n3794_), .Y(new_n3795_));
  INVX1    g01360(.A(new_n3709_), .Y(new_n3796_));
  INVX1    g01361(.A(new_n3240_), .Y(new_n3797_));
  OAI21X1  g01362(.A0(new_n3797_), .A1(pi0861), .B0(new_n3715_), .Y(new_n3798_));
  INVX1    g01363(.A(new_n3244_), .Y(new_n3799_));
  AOI21X1  g01364(.A0(new_n3799_), .A1(new_n3716_), .B0(new_n3715_), .Y(new_n3800_));
  OAI21X1  g01365(.A0(new_n3570_), .A1(new_n3716_), .B0(new_n3800_), .Y(new_n3801_));
  AOI21X1  g01366(.A0(new_n3801_), .A1(new_n3798_), .B0(pi0228), .Y(new_n3802_));
  OAI21X1  g01367(.A0(new_n3232_), .A1(new_n3011_), .B0(new_n3750_), .Y(new_n3803_));
  OAI21X1  g01368(.A0(new_n3803_), .A1(new_n3802_), .B0(new_n3714_), .Y(new_n3804_));
  AOI21X1  g01369(.A0(new_n3804_), .A1(new_n3712_), .B0(pi0215), .Y(new_n3805_));
  OAI21X1  g01370(.A0(new_n3805_), .A1(new_n3796_), .B0(new_n3741_), .Y(new_n3806_));
  INVX1    g01371(.A(new_n3262_), .Y(new_n3807_));
  AND2X1   g01372(.A(new_n3746_), .B(new_n3807_), .Y(new_n3808_));
  INVX1    g01373(.A(new_n3808_), .Y(new_n3809_));
  NOR3X1   g01374(.A(new_n3725_), .B(new_n3254_), .C(pi0216), .Y(new_n3810_));
  AOI21X1  g01375(.A0(new_n3810_), .A1(new_n3752_), .B0(new_n3749_), .Y(new_n3811_));
  OAI21X1  g01376(.A0(new_n3811_), .A1(new_n3713_), .B0(new_n2934_), .Y(new_n3812_));
  AOI21X1  g01377(.A0(new_n3812_), .A1(new_n3748_), .B0(new_n2933_), .Y(new_n3813_));
  NOR2X1   g01378(.A(new_n3813_), .B(new_n3809_), .Y(new_n3814_));
  INVX1    g01379(.A(new_n3814_), .Y(new_n3815_));
  AOI21X1  g01380(.A0(new_n3815_), .A1(pi0039), .B0(pi0038), .Y(new_n3816_));
  INVX1    g01381(.A(pi0270), .Y(new_n3817_));
  OAI21X1  g01382(.A0(new_n3817_), .A1(new_n2438_), .B0(new_n3339_), .Y(new_n3818_));
  AND2X1   g01383(.A(new_n3818_), .B(new_n3762_), .Y(new_n3819_));
  INVX1    g01384(.A(new_n3819_), .Y(new_n3820_));
  AOI21X1  g01385(.A0(new_n3820_), .A1(pi0299), .B0(new_n3809_), .Y(new_n3821_));
  INVX1    g01386(.A(new_n3821_), .Y(new_n3822_));
  OAI21X1  g01387(.A0(new_n3822_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3823_));
  AOI21X1  g01388(.A0(new_n3816_), .A1(new_n3806_), .B0(new_n3823_), .Y(new_n3824_));
  AND2X1   g01389(.A(new_n3810_), .B(new_n3768_), .Y(new_n3825_));
  OAI21X1  g01390(.A0(new_n3825_), .A1(new_n3749_), .B0(new_n3712_), .Y(new_n3826_));
  AOI21X1  g01391(.A0(new_n3826_), .A1(new_n2934_), .B0(new_n3708_), .Y(new_n3827_));
  AND3X1   g01392(.A(new_n3746_), .B(new_n3807_), .C(new_n3047_), .Y(new_n3828_));
  OAI21X1  g01393(.A0(new_n3827_), .A1(new_n2933_), .B0(new_n3828_), .Y(new_n3829_));
  AOI21X1  g01394(.A0(new_n3821_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n3830_));
  AND2X1   g01395(.A(new_n3830_), .B(new_n3829_), .Y(new_n3831_));
  OAI21X1  g01396(.A0(new_n3831_), .A1(new_n3824_), .B0(new_n3131_), .Y(new_n3832_));
  MX2X1    g01397(.A(new_n3822_), .B(new_n3815_), .S0(new_n3064_), .Y(new_n3833_));
  AOI21X1  g01398(.A0(new_n3833_), .A1(pi0087), .B0(pi0075), .Y(new_n3834_));
  OAI21X1  g01399(.A0(new_n3822_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3835_));
  AOI21X1  g01400(.A0(new_n3834_), .A1(new_n3832_), .B0(new_n3835_), .Y(new_n3836_));
  AOI21X1  g01401(.A0(new_n3821_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n3837_));
  OAI21X1  g01402(.A0(new_n3833_), .A1(new_n3080_), .B0(new_n3837_), .Y(new_n3838_));
  NAND2X1  g01403(.A(new_n3838_), .B(new_n3102_), .Y(new_n3839_));
  OR2X1    g01404(.A(new_n3839_), .B(new_n3836_), .Y(new_n3840_));
  AOI21X1  g01405(.A0(new_n3821_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3841_));
  AND3X1   g01406(.A(new_n3812_), .B(new_n3748_), .C(new_n3104_), .Y(new_n3842_));
  OAI21X1  g01407(.A0(new_n3820_), .A1(new_n3104_), .B0(pi0055), .Y(new_n3843_));
  OAI21X1  g01408(.A0(new_n3843_), .A1(new_n3842_), .B0(new_n3118_), .Y(new_n3844_));
  AOI21X1  g01409(.A0(new_n3841_), .A1(new_n3840_), .B0(new_n3844_), .Y(new_n3845_));
  AOI21X1  g01410(.A0(new_n3812_), .A1(new_n3748_), .B0(new_n3115_), .Y(new_n3846_));
  OAI21X1  g01411(.A0(new_n3819_), .A1(new_n3114_), .B0(pi0056), .Y(new_n3847_));
  OAI21X1  g01412(.A0(new_n3847_), .A1(new_n3846_), .B0(new_n3222_), .Y(new_n3848_));
  NAND3X1  g01413(.A(new_n3812_), .B(new_n3748_), .C(new_n3224_), .Y(new_n3849_));
  AOI21X1  g01414(.A0(new_n3819_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n3850_));
  NAND2X1  g01415(.A(new_n3223_), .B(pi0241), .Y(new_n3851_));
  AOI21X1  g01416(.A0(new_n3850_), .A1(new_n3849_), .B0(new_n3851_), .Y(new_n3852_));
  OAI21X1  g01417(.A0(new_n3848_), .A1(new_n3845_), .B0(new_n3852_), .Y(new_n3853_));
  INVX1    g01418(.A(pi0241), .Y(new_n3854_));
  OR2X1    g01419(.A(new_n3818_), .B(new_n3854_), .Y(new_n3855_));
  NAND3X1  g01420(.A(new_n3855_), .B(new_n3762_), .C(new_n3374_), .Y(new_n3856_));
  AND3X1   g01421(.A(new_n3856_), .B(new_n3853_), .C(new_n3795_), .Y(po0158));
  AND2X1   g01422(.A(pi1140), .B(pi0215), .Y(new_n3858_));
  NOR2X1   g01423(.A(new_n3858_), .B(new_n2933_), .Y(new_n3859_));
  INVX1    g01424(.A(pi0921), .Y(new_n3860_));
  AOI21X1  g01425(.A0(new_n3145_), .A1(new_n3860_), .B0(new_n2437_), .Y(new_n3861_));
  OAI21X1  g01426(.A0(new_n3145_), .A1(pi1140), .B0(new_n3861_), .Y(new_n3862_));
  INVX1    g01427(.A(new_n3862_), .Y(new_n3863_));
  AOI21X1  g01428(.A0(pi0282), .A1(pi0216), .B0(pi0221), .Y(new_n3864_));
  INVX1    g01429(.A(pi0170), .Y(new_n3865_));
  INVX1    g01430(.A(pi0869), .Y(new_n3866_));
  OR3X1    g01431(.A(new_n3232_), .B(new_n2696_), .C(new_n3866_), .Y(new_n3867_));
  AND2X1   g01432(.A(new_n3867_), .B(new_n3865_), .Y(new_n3868_));
  MX2X1    g01433(.A(new_n3867_), .B(new_n3240_), .S0(pi0170), .Y(new_n3869_));
  AOI22X1  g01434(.A0(new_n3869_), .A1(pi0869), .B0(new_n3868_), .B1(new_n3180_), .Y(new_n3870_));
  AOI21X1  g01435(.A0(new_n2453_), .A1(pi0095), .B0(new_n3866_), .Y(new_n3871_));
  INVX1    g01436(.A(new_n3871_), .Y(new_n3872_));
  OAI21X1  g01437(.A0(new_n3865_), .A1(pi0105), .B0(pi0228), .Y(new_n3873_));
  AOI21X1  g01438(.A0(new_n3872_), .A1(pi0105), .B0(new_n3873_), .Y(new_n3874_));
  AOI21X1  g01439(.A0(new_n3874_), .A1(new_n3721_), .B0(pi0216), .Y(new_n3875_));
  OAI21X1  g01440(.A0(new_n3870_), .A1(pi0228), .B0(new_n3875_), .Y(new_n3876_));
  AOI21X1  g01441(.A0(new_n3876_), .A1(new_n3864_), .B0(new_n3863_), .Y(new_n3877_));
  OAI21X1  g01442(.A0(new_n3877_), .A1(pi0215), .B0(new_n3859_), .Y(new_n3878_));
  AND2X1   g01443(.A(pi1140), .B(pi0223), .Y(new_n3879_));
  AOI21X1  g01444(.A0(new_n3134_), .A1(new_n3860_), .B0(new_n2941_), .Y(new_n3880_));
  OAI21X1  g01445(.A0(new_n3134_), .A1(pi1140), .B0(new_n3880_), .Y(new_n3881_));
  AOI21X1  g01446(.A0(pi0282), .A1(pi0224), .B0(pi0222), .Y(new_n3882_));
  INVX1    g01447(.A(new_n3882_), .Y(new_n3883_));
  AOI21X1  g01448(.A0(new_n3232_), .A1(pi0869), .B0(pi0224), .Y(new_n3884_));
  OAI21X1  g01449(.A0(new_n3884_), .A1(new_n3883_), .B0(new_n3881_), .Y(new_n3885_));
  OR3X1    g01450(.A(new_n3885_), .B(new_n3879_), .C(pi0299), .Y(new_n3886_));
  AOI21X1  g01451(.A0(pi1140), .A1(pi0223), .B0(pi0299), .Y(new_n3887_));
  NOR2X1   g01452(.A(new_n3883_), .B(new_n3232_), .Y(new_n3888_));
  OAI21X1  g01453(.A0(new_n3888_), .A1(new_n3885_), .B0(new_n2940_), .Y(new_n3889_));
  AOI21X1  g01454(.A0(new_n3889_), .A1(new_n3887_), .B0(pi0039), .Y(new_n3890_));
  AND2X1   g01455(.A(new_n3890_), .B(new_n3886_), .Y(new_n3891_));
  AOI21X1  g01456(.A0(new_n3872_), .A1(new_n2942_), .B0(new_n3883_), .Y(new_n3892_));
  INVX1    g01457(.A(new_n3892_), .Y(new_n3893_));
  AOI21X1  g01458(.A0(new_n3893_), .A1(new_n3881_), .B0(pi0223), .Y(new_n3894_));
  OAI21X1  g01459(.A0(new_n3894_), .A1(new_n3879_), .B0(new_n2933_), .Y(new_n3895_));
  INVX1    g01460(.A(new_n3895_), .Y(new_n3896_));
  INVX1    g01461(.A(new_n3858_), .Y(new_n3897_));
  INVX1    g01462(.A(new_n3864_), .Y(new_n3898_));
  NOR2X1   g01463(.A(new_n3874_), .B(pi0216), .Y(new_n3899_));
  AOI21X1  g01464(.A0(new_n2986_), .A1(pi0170), .B0(pi0228), .Y(new_n3900_));
  OAI21X1  g01465(.A0(new_n2986_), .A1(pi0869), .B0(new_n3900_), .Y(new_n3901_));
  AOI21X1  g01466(.A0(new_n3901_), .A1(new_n3899_), .B0(new_n3898_), .Y(new_n3902_));
  OAI21X1  g01467(.A0(new_n3902_), .A1(new_n3863_), .B0(new_n2934_), .Y(new_n3903_));
  AOI21X1  g01468(.A0(new_n3903_), .A1(new_n3897_), .B0(new_n2933_), .Y(new_n3904_));
  NOR2X1   g01469(.A(new_n3904_), .B(new_n3896_), .Y(new_n3905_));
  OAI21X1  g01470(.A0(new_n3905_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n3906_));
  AOI21X1  g01471(.A0(new_n3891_), .A1(new_n3878_), .B0(new_n3906_), .Y(new_n3907_));
  INVX1    g01472(.A(pi1140), .Y(new_n3908_));
  OAI21X1  g01473(.A0(pi0228), .A1(pi0170), .B0(new_n3899_), .Y(new_n3909_));
  AOI21X1  g01474(.A0(new_n3909_), .A1(new_n3864_), .B0(new_n3863_), .Y(new_n3910_));
  MX2X1    g01475(.A(new_n3910_), .B(new_n3908_), .S0(pi0215), .Y(new_n3911_));
  INVX1    g01476(.A(new_n3911_), .Y(new_n3912_));
  AOI21X1  g01477(.A0(new_n3912_), .A1(pi0299), .B0(new_n3896_), .Y(new_n3913_));
  INVX1    g01478(.A(new_n3913_), .Y(new_n3914_));
  OAI21X1  g01479(.A0(new_n3914_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3915_));
  AOI21X1  g01480(.A0(new_n3199_), .A1(pi0170), .B0(pi0228), .Y(new_n3916_));
  OAI21X1  g01481(.A0(new_n3199_), .A1(pi0869), .B0(new_n3916_), .Y(new_n3917_));
  AOI21X1  g01482(.A0(new_n3917_), .A1(new_n3899_), .B0(new_n3898_), .Y(new_n3918_));
  OAI21X1  g01483(.A0(new_n3918_), .A1(new_n3863_), .B0(new_n2934_), .Y(new_n3919_));
  AOI21X1  g01484(.A0(new_n3919_), .A1(new_n3897_), .B0(new_n2933_), .Y(new_n3920_));
  NOR3X1   g01485(.A(new_n3920_), .B(new_n3896_), .C(new_n3060_), .Y(new_n3921_));
  OAI21X1  g01486(.A0(new_n3914_), .A1(new_n3047_), .B0(pi0100), .Y(new_n3922_));
  OAI22X1  g01487(.A0(new_n3922_), .A1(new_n3921_), .B0(new_n3915_), .B1(new_n3907_), .Y(new_n3923_));
  MX2X1    g01488(.A(new_n3913_), .B(new_n3905_), .S0(new_n3064_), .Y(new_n3924_));
  OAI21X1  g01489(.A0(new_n3924_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n3925_));
  AOI21X1  g01490(.A0(new_n3923_), .A1(new_n3131_), .B0(new_n3925_), .Y(new_n3926_));
  OAI21X1  g01491(.A0(new_n3914_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3927_));
  NAND2X1  g01492(.A(new_n3924_), .B(new_n3077_), .Y(new_n3928_));
  AOI21X1  g01493(.A0(new_n3913_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n3929_));
  AOI21X1  g01494(.A0(new_n3929_), .A1(new_n3928_), .B0(new_n3130_), .Y(new_n3930_));
  OAI21X1  g01495(.A0(new_n3927_), .A1(new_n3926_), .B0(new_n3930_), .Y(new_n3931_));
  AOI21X1  g01496(.A0(new_n3913_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3932_));
  AND3X1   g01497(.A(new_n3903_), .B(new_n3897_), .C(new_n3104_), .Y(new_n3933_));
  OAI21X1  g01498(.A0(new_n3912_), .A1(new_n3104_), .B0(pi0055), .Y(new_n3934_));
  OAI21X1  g01499(.A0(new_n3934_), .A1(new_n3933_), .B0(new_n3118_), .Y(new_n3935_));
  AOI21X1  g01500(.A0(new_n3932_), .A1(new_n3931_), .B0(new_n3935_), .Y(new_n3936_));
  AOI21X1  g01501(.A0(new_n3903_), .A1(new_n3897_), .B0(new_n3115_), .Y(new_n3937_));
  OAI21X1  g01502(.A0(new_n3911_), .A1(new_n3114_), .B0(pi0056), .Y(new_n3938_));
  OAI21X1  g01503(.A0(new_n3938_), .A1(new_n3937_), .B0(new_n3222_), .Y(new_n3939_));
  NAND3X1  g01504(.A(new_n3903_), .B(new_n3897_), .C(new_n3224_), .Y(new_n3940_));
  AOI21X1  g01505(.A0(new_n3911_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n3941_));
  OR3X1    g01506(.A(pi0248), .B(pi0059), .C(pi0057), .Y(new_n3942_));
  AOI21X1  g01507(.A0(new_n3941_), .A1(new_n3940_), .B0(new_n3942_), .Y(new_n3943_));
  OAI21X1  g01508(.A0(new_n3939_), .A1(new_n3936_), .B0(new_n3943_), .Y(new_n3944_));
  INVX1    g01509(.A(new_n3859_), .Y(new_n3945_));
  OAI21X1  g01510(.A0(new_n3797_), .A1(pi0869), .B0(new_n3865_), .Y(new_n3946_));
  AOI21X1  g01511(.A0(new_n3799_), .A1(new_n3866_), .B0(new_n3865_), .Y(new_n3947_));
  OAI21X1  g01512(.A0(new_n3570_), .A1(new_n3866_), .B0(new_n3947_), .Y(new_n3948_));
  AOI21X1  g01513(.A0(new_n3948_), .A1(new_n3946_), .B0(pi0228), .Y(new_n3949_));
  OAI21X1  g01514(.A0(new_n3232_), .A1(new_n3011_), .B0(new_n3899_), .Y(new_n3950_));
  OAI21X1  g01515(.A0(new_n3950_), .A1(new_n3949_), .B0(new_n3864_), .Y(new_n3951_));
  AOI21X1  g01516(.A0(new_n3951_), .A1(new_n3862_), .B0(pi0215), .Y(new_n3952_));
  OAI21X1  g01517(.A0(new_n3952_), .A1(new_n3945_), .B0(new_n3890_), .Y(new_n3953_));
  AND2X1   g01518(.A(new_n3895_), .B(new_n3807_), .Y(new_n3954_));
  INVX1    g01519(.A(new_n3954_), .Y(new_n3955_));
  NOR3X1   g01520(.A(new_n3874_), .B(new_n3254_), .C(pi0216), .Y(new_n3956_));
  AOI21X1  g01521(.A0(new_n3956_), .A1(new_n3901_), .B0(new_n3898_), .Y(new_n3957_));
  OAI21X1  g01522(.A0(new_n3957_), .A1(new_n3863_), .B0(new_n2934_), .Y(new_n3958_));
  AOI21X1  g01523(.A0(new_n3958_), .A1(new_n3897_), .B0(new_n2933_), .Y(new_n3959_));
  NOR2X1   g01524(.A(new_n3959_), .B(new_n3955_), .Y(new_n3960_));
  INVX1    g01525(.A(new_n3960_), .Y(new_n3961_));
  AOI21X1  g01526(.A0(new_n3961_), .A1(pi0039), .B0(pi0038), .Y(new_n3962_));
  INVX1    g01527(.A(pi0282), .Y(new_n3963_));
  OAI21X1  g01528(.A0(new_n3963_), .A1(new_n2438_), .B0(new_n3339_), .Y(new_n3964_));
  AND2X1   g01529(.A(new_n3964_), .B(new_n3911_), .Y(new_n3965_));
  INVX1    g01530(.A(new_n3965_), .Y(new_n3966_));
  AOI21X1  g01531(.A0(new_n3966_), .A1(pi0299), .B0(new_n3955_), .Y(new_n3967_));
  INVX1    g01532(.A(new_n3967_), .Y(new_n3968_));
  OAI21X1  g01533(.A0(new_n3968_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n3969_));
  AOI21X1  g01534(.A0(new_n3962_), .A1(new_n3953_), .B0(new_n3969_), .Y(new_n3970_));
  AND2X1   g01535(.A(new_n3956_), .B(new_n3917_), .Y(new_n3971_));
  OAI21X1  g01536(.A0(new_n3971_), .A1(new_n3898_), .B0(new_n3862_), .Y(new_n3972_));
  AOI21X1  g01537(.A0(new_n3972_), .A1(new_n2934_), .B0(new_n3858_), .Y(new_n3973_));
  AND3X1   g01538(.A(new_n3895_), .B(new_n3807_), .C(new_n3047_), .Y(new_n3974_));
  OAI21X1  g01539(.A0(new_n3973_), .A1(new_n2933_), .B0(new_n3974_), .Y(new_n3975_));
  AOI21X1  g01540(.A0(new_n3967_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n3976_));
  AND2X1   g01541(.A(new_n3976_), .B(new_n3975_), .Y(new_n3977_));
  OAI21X1  g01542(.A0(new_n3977_), .A1(new_n3970_), .B0(new_n3131_), .Y(new_n3978_));
  MX2X1    g01543(.A(new_n3968_), .B(new_n3961_), .S0(new_n3064_), .Y(new_n3979_));
  AOI21X1  g01544(.A0(new_n3979_), .A1(pi0087), .B0(pi0075), .Y(new_n3980_));
  OAI21X1  g01545(.A0(new_n3968_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n3981_));
  AOI21X1  g01546(.A0(new_n3980_), .A1(new_n3978_), .B0(new_n3981_), .Y(new_n3982_));
  AOI21X1  g01547(.A0(new_n3967_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n3983_));
  OAI21X1  g01548(.A0(new_n3979_), .A1(new_n3080_), .B0(new_n3983_), .Y(new_n3984_));
  NAND2X1  g01549(.A(new_n3984_), .B(new_n3102_), .Y(new_n3985_));
  OR2X1    g01550(.A(new_n3985_), .B(new_n3982_), .Y(new_n3986_));
  AOI21X1  g01551(.A0(new_n3967_), .A1(new_n3130_), .B0(pi0055), .Y(new_n3987_));
  AND3X1   g01552(.A(new_n3958_), .B(new_n3897_), .C(new_n3104_), .Y(new_n3988_));
  OAI21X1  g01553(.A0(new_n3966_), .A1(new_n3104_), .B0(pi0055), .Y(new_n3989_));
  OAI21X1  g01554(.A0(new_n3989_), .A1(new_n3988_), .B0(new_n3118_), .Y(new_n3990_));
  AOI21X1  g01555(.A0(new_n3987_), .A1(new_n3986_), .B0(new_n3990_), .Y(new_n3991_));
  AOI21X1  g01556(.A0(new_n3958_), .A1(new_n3897_), .B0(new_n3115_), .Y(new_n3992_));
  OAI21X1  g01557(.A0(new_n3965_), .A1(new_n3114_), .B0(pi0056), .Y(new_n3993_));
  OAI21X1  g01558(.A0(new_n3993_), .A1(new_n3992_), .B0(new_n3222_), .Y(new_n3994_));
  NAND3X1  g01559(.A(new_n3958_), .B(new_n3897_), .C(new_n3224_), .Y(new_n3995_));
  AOI21X1  g01560(.A0(new_n3965_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n3996_));
  NAND2X1  g01561(.A(new_n3223_), .B(pi0248), .Y(new_n3997_));
  AOI21X1  g01562(.A0(new_n3996_), .A1(new_n3995_), .B0(new_n3997_), .Y(new_n3998_));
  OAI21X1  g01563(.A0(new_n3994_), .A1(new_n3991_), .B0(new_n3998_), .Y(new_n3999_));
  INVX1    g01564(.A(pi0248), .Y(new_n4000_));
  OR2X1    g01565(.A(new_n3964_), .B(new_n4000_), .Y(new_n4001_));
  NAND3X1  g01566(.A(new_n4001_), .B(new_n3911_), .C(new_n3374_), .Y(new_n4002_));
  AND3X1   g01567(.A(new_n4002_), .B(new_n3999_), .C(new_n3944_), .Y(po0159));
  NOR2X1   g01568(.A(pi0215), .B(pi0148), .Y(new_n4004_));
  INVX1    g01569(.A(new_n4004_), .Y(new_n4005_));
  AND2X1   g01570(.A(pi0920), .B(pi0833), .Y(new_n4006_));
  INVX1    g01571(.A(new_n4006_), .Y(new_n4007_));
  AOI21X1  g01572(.A0(pi1139), .A1(new_n2701_), .B0(pi0216), .Y(new_n4008_));
  AOI21X1  g01573(.A0(new_n4008_), .A1(new_n4007_), .B0(new_n2437_), .Y(new_n4009_));
  OAI21X1  g01574(.A0(pi1139), .A1(new_n2438_), .B0(new_n4009_), .Y(new_n4010_));
  INVX1    g01575(.A(new_n4010_), .Y(new_n4011_));
  AOI21X1  g01576(.A0(pi0281), .A1(pi0216), .B0(pi0221), .Y(new_n4012_));
  AOI21X1  g01577(.A0(new_n3456_), .A1(pi0862), .B0(pi0216), .Y(new_n4013_));
  OAI21X1  g01578(.A0(new_n3603_), .A1(new_n3009_), .B0(new_n4013_), .Y(new_n4014_));
  AOI21X1  g01579(.A0(new_n4014_), .A1(new_n4012_), .B0(new_n4011_), .Y(new_n4015_));
  INVX1    g01580(.A(new_n4012_), .Y(new_n4016_));
  OR3X1    g01581(.A(new_n4016_), .B(new_n3627_), .C(new_n3009_), .Y(new_n4017_));
  AOI21X1  g01582(.A0(new_n4017_), .A1(new_n4015_), .B0(new_n4005_), .Y(new_n4018_));
  INVX1    g01583(.A(pi1139), .Y(new_n4019_));
  AOI21X1  g01584(.A0(new_n3009_), .A1(new_n3348_), .B0(new_n3603_), .Y(new_n4020_));
  NOR3X1   g01585(.A(new_n4020_), .B(pi0862), .C(pi0216), .Y(new_n4021_));
  OAI21X1  g01586(.A0(new_n4021_), .A1(new_n4016_), .B0(new_n4010_), .Y(new_n4022_));
  AOI21X1  g01587(.A0(new_n4012_), .A1(new_n3349_), .B0(new_n4022_), .Y(new_n4023_));
  AND2X1   g01588(.A(new_n2934_), .B(pi0148), .Y(new_n4024_));
  INVX1    g01589(.A(new_n4024_), .Y(new_n4025_));
  NOR2X1   g01590(.A(new_n4009_), .B(pi0216), .Y(new_n4026_));
  AND2X1   g01591(.A(new_n4026_), .B(new_n3349_), .Y(new_n4027_));
  OR3X1    g01592(.A(new_n4027_), .B(new_n4025_), .C(new_n4023_), .Y(new_n4028_));
  OAI21X1  g01593(.A0(new_n4019_), .A1(new_n2934_), .B0(new_n4028_), .Y(new_n4029_));
  OAI21X1  g01594(.A0(new_n4029_), .A1(new_n4018_), .B0(pi0299), .Y(new_n4030_));
  OAI21X1  g01595(.A0(new_n3310_), .A1(pi0920), .B0(pi0222), .Y(new_n4031_));
  AOI21X1  g01596(.A0(new_n3310_), .A1(new_n4019_), .B0(new_n4031_), .Y(new_n4032_));
  AND2X1   g01597(.A(pi1139), .B(pi0223), .Y(new_n4033_));
  NOR3X1   g01598(.A(new_n4033_), .B(new_n4032_), .C(pi0224), .Y(new_n4034_));
  INVX1    g01599(.A(new_n4034_), .Y(new_n4035_));
  NOR4X1   g01600(.A(new_n4033_), .B(new_n4032_), .C(pi0862), .D(pi0224), .Y(new_n4036_));
  AOI21X1  g01601(.A0(pi0281), .A1(pi0224), .B0(pi0222), .Y(new_n4037_));
  NOR2X1   g01602(.A(new_n4037_), .B(new_n4032_), .Y(new_n4038_));
  MX2X1    g01603(.A(new_n4038_), .B(new_n4019_), .S0(pi0223), .Y(new_n4039_));
  NOR3X1   g01604(.A(new_n4039_), .B(new_n4036_), .C(pi0299), .Y(new_n4040_));
  OAI21X1  g01605(.A0(new_n4035_), .A1(new_n3348_), .B0(new_n4040_), .Y(new_n4041_));
  AND2X1   g01606(.A(new_n4041_), .B(new_n3047_), .Y(new_n4042_));
  INVX1    g01607(.A(new_n4041_), .Y(new_n4043_));
  NOR4X1   g01608(.A(new_n3011_), .B(new_n2454_), .C(pi0862), .D(pi0216), .Y(new_n4044_));
  OAI21X1  g01609(.A0(new_n4044_), .A1(new_n4016_), .B0(new_n4010_), .Y(new_n4045_));
  INVX1    g01610(.A(pi0148), .Y(new_n4046_));
  OR4X1    g01611(.A(new_n4009_), .B(new_n3009_), .C(pi0216), .D(new_n4046_), .Y(new_n4047_));
  AND2X1   g01612(.A(new_n4047_), .B(new_n2934_), .Y(new_n4048_));
  AOI22X1  g01613(.A0(new_n4048_), .A1(new_n4045_), .B0(pi1139), .B1(pi0215), .Y(new_n4049_));
  NOR2X1   g01614(.A(new_n4049_), .B(new_n3255_), .Y(new_n4050_));
  AOI21X1  g01615(.A0(new_n4050_), .A1(pi0299), .B0(new_n4043_), .Y(new_n4051_));
  INVX1    g01616(.A(new_n4051_), .Y(new_n4052_));
  OAI21X1  g01617(.A0(new_n4052_), .A1(new_n3047_), .B0(pi0100), .Y(new_n4053_));
  AOI21X1  g01618(.A0(new_n4042_), .A1(new_n4030_), .B0(new_n4053_), .Y(new_n4054_));
  INVX1    g01619(.A(pi0862), .Y(new_n4055_));
  MX2X1    g01620(.A(new_n3180_), .B(new_n2447_), .S0(pi0228), .Y(new_n4056_));
  OAI21X1  g01621(.A0(new_n3245_), .A1(new_n4055_), .B0(new_n2438_), .Y(new_n4057_));
  AOI21X1  g01622(.A0(new_n4056_), .A1(new_n4055_), .B0(new_n4057_), .Y(new_n4058_));
  OAI21X1  g01623(.A0(new_n4058_), .A1(new_n4016_), .B0(new_n4010_), .Y(new_n4059_));
  AND2X1   g01624(.A(new_n4059_), .B(new_n4004_), .Y(new_n4060_));
  NOR3X1   g01625(.A(new_n3241_), .B(pi0862), .C(pi0216), .Y(new_n4061_));
  OAI21X1  g01626(.A0(new_n4061_), .A1(new_n4016_), .B0(new_n4010_), .Y(new_n4062_));
  INVX1    g01627(.A(new_n4062_), .Y(new_n4063_));
  AND2X1   g01628(.A(new_n4026_), .B(new_n3241_), .Y(new_n4064_));
  OR2X1    g01629(.A(new_n4064_), .B(new_n4025_), .Y(new_n4065_));
  AOI21X1  g01630(.A0(pi1139), .A1(pi0215), .B0(new_n2933_), .Y(new_n4066_));
  OAI21X1  g01631(.A0(new_n4065_), .A1(new_n4063_), .B0(new_n4066_), .Y(new_n4067_));
  NOR2X1   g01632(.A(new_n4039_), .B(new_n4036_), .Y(new_n4068_));
  OAI21X1  g01633(.A0(new_n4035_), .A1(new_n3232_), .B0(new_n4068_), .Y(new_n4069_));
  AOI21X1  g01634(.A0(new_n4069_), .A1(new_n2933_), .B0(pi0039), .Y(new_n4070_));
  OAI21X1  g01635(.A0(new_n4067_), .A1(new_n4060_), .B0(new_n4070_), .Y(new_n4071_));
  AOI21X1  g01636(.A0(new_n4026_), .A1(new_n4020_), .B0(new_n4025_), .Y(new_n4072_));
  AOI22X1  g01637(.A0(new_n4072_), .A1(new_n4022_), .B0(pi1139), .B1(pi0215), .Y(new_n4073_));
  OAI21X1  g01638(.A0(new_n4015_), .A1(new_n4005_), .B0(new_n4073_), .Y(new_n4074_));
  AOI21X1  g01639(.A0(new_n4074_), .A1(pi0299), .B0(new_n4043_), .Y(new_n4075_));
  INVX1    g01640(.A(new_n4075_), .Y(new_n4076_));
  AOI21X1  g01641(.A0(new_n4076_), .A1(pi0039), .B0(pi0038), .Y(new_n4077_));
  OAI21X1  g01642(.A0(new_n4052_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4078_));
  AOI21X1  g01643(.A0(new_n4077_), .A1(new_n4071_), .B0(new_n4078_), .Y(new_n4079_));
  OAI21X1  g01644(.A0(new_n4079_), .A1(new_n4054_), .B0(new_n3131_), .Y(new_n4080_));
  MX2X1    g01645(.A(new_n4052_), .B(new_n4076_), .S0(new_n3064_), .Y(new_n4081_));
  AOI21X1  g01646(.A0(new_n4081_), .A1(pi0087), .B0(pi0075), .Y(new_n4082_));
  OAI21X1  g01647(.A0(new_n4052_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4083_));
  AOI21X1  g01648(.A0(new_n4082_), .A1(new_n4080_), .B0(new_n4083_), .Y(new_n4084_));
  OR2X1    g01649(.A(new_n4081_), .B(new_n3080_), .Y(new_n4085_));
  AOI21X1  g01650(.A0(new_n4051_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4086_));
  AND2X1   g01651(.A(new_n4086_), .B(new_n4085_), .Y(new_n4087_));
  NOR3X1   g01652(.A(new_n4087_), .B(new_n4084_), .C(new_n3130_), .Y(new_n4088_));
  OAI21X1  g01653(.A0(new_n4052_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4089_));
  OAI21X1  g01654(.A0(new_n4049_), .A1(new_n3255_), .B0(new_n3105_), .Y(new_n4090_));
  AND2X1   g01655(.A(new_n4090_), .B(pi0055), .Y(new_n4091_));
  OAI21X1  g01656(.A0(new_n4074_), .A1(new_n3105_), .B0(new_n4091_), .Y(new_n4092_));
  AND2X1   g01657(.A(new_n4092_), .B(new_n3118_), .Y(new_n4093_));
  OAI21X1  g01658(.A0(new_n4089_), .A1(new_n4088_), .B0(new_n4093_), .Y(new_n4094_));
  NAND2X1  g01659(.A(new_n4074_), .B(new_n3114_), .Y(new_n4095_));
  AOI21X1  g01660(.A0(new_n4050_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4096_));
  AOI21X1  g01661(.A0(new_n4096_), .A1(new_n4095_), .B0(pi0062), .Y(new_n4097_));
  NOR2X1   g01662(.A(new_n4074_), .B(new_n3225_), .Y(new_n4098_));
  OAI21X1  g01663(.A0(new_n4050_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4099_));
  OAI21X1  g01664(.A0(new_n4099_), .A1(new_n4098_), .B0(new_n3223_), .Y(new_n4100_));
  AOI21X1  g01665(.A0(new_n4097_), .A1(new_n4094_), .B0(new_n4100_), .Y(new_n4101_));
  INVX1    g01666(.A(pi0247), .Y(new_n4102_));
  OAI21X1  g01667(.A0(new_n4050_), .A1(new_n3223_), .B0(new_n4102_), .Y(new_n4103_));
  NOR2X1   g01668(.A(new_n4023_), .B(new_n4005_), .Y(new_n4104_));
  NOR4X1   g01669(.A(new_n4011_), .B(new_n3627_), .C(new_n3009_), .D(pi0216), .Y(new_n4105_));
  NAND2X1  g01670(.A(new_n4024_), .B(new_n4022_), .Y(new_n4106_));
  OAI22X1  g01671(.A0(new_n4106_), .A1(new_n4105_), .B0(new_n4019_), .B1(new_n2934_), .Y(new_n4107_));
  OAI21X1  g01672(.A0(new_n4107_), .A1(new_n4104_), .B0(pi0299), .Y(new_n4108_));
  NOR3X1   g01673(.A(new_n4040_), .B(new_n3262_), .C(new_n3060_), .Y(new_n4109_));
  INVX1    g01674(.A(new_n4049_), .Y(new_n4110_));
  NOR2X1   g01675(.A(new_n4040_), .B(new_n3262_), .Y(new_n4111_));
  INVX1    g01676(.A(new_n4111_), .Y(new_n4112_));
  AOI21X1  g01677(.A0(new_n4110_), .A1(pi0299), .B0(new_n4112_), .Y(new_n4113_));
  INVX1    g01678(.A(new_n4113_), .Y(new_n4114_));
  OAI21X1  g01679(.A0(new_n4114_), .A1(new_n3047_), .B0(pi0100), .Y(new_n4115_));
  AOI21X1  g01680(.A0(new_n4109_), .A1(new_n4108_), .B0(new_n4115_), .Y(new_n4116_));
  OR2X1    g01681(.A(new_n4039_), .B(pi0299), .Y(new_n4117_));
  AOI21X1  g01682(.A0(new_n4036_), .A1(new_n3232_), .B0(new_n4117_), .Y(new_n4118_));
  AOI21X1  g01683(.A0(new_n3245_), .A1(new_n4055_), .B0(pi0216), .Y(new_n4119_));
  OAI21X1  g01684(.A0(new_n4056_), .A1(new_n4055_), .B0(new_n4119_), .Y(new_n4120_));
  AOI21X1  g01685(.A0(new_n4120_), .A1(new_n4012_), .B0(new_n4011_), .Y(new_n4121_));
  OR2X1    g01686(.A(new_n4121_), .B(new_n4025_), .Y(new_n4122_));
  AOI22X1  g01687(.A0(new_n4062_), .A1(new_n4004_), .B0(pi1139), .B1(pi0215), .Y(new_n4123_));
  AOI21X1  g01688(.A0(new_n4123_), .A1(new_n4122_), .B0(new_n2933_), .Y(new_n4124_));
  OAI21X1  g01689(.A0(new_n4124_), .A1(new_n4118_), .B0(new_n2939_), .Y(new_n4125_));
  NAND2X1  g01690(.A(new_n4048_), .B(new_n4022_), .Y(new_n4126_));
  AND2X1   g01691(.A(new_n4126_), .B(new_n4073_), .Y(new_n4127_));
  OAI21X1  g01692(.A0(new_n4127_), .A1(new_n2933_), .B0(new_n4111_), .Y(new_n4128_));
  AOI21X1  g01693(.A0(new_n4128_), .A1(pi0039), .B0(pi0038), .Y(new_n4129_));
  OAI21X1  g01694(.A0(new_n4114_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4130_));
  AOI21X1  g01695(.A0(new_n4129_), .A1(new_n4125_), .B0(new_n4130_), .Y(new_n4131_));
  OAI21X1  g01696(.A0(new_n4131_), .A1(new_n4116_), .B0(new_n3131_), .Y(new_n4132_));
  MX2X1    g01697(.A(new_n4114_), .B(new_n4128_), .S0(new_n3064_), .Y(new_n4133_));
  AOI21X1  g01698(.A0(new_n4133_), .A1(pi0087), .B0(pi0075), .Y(new_n4134_));
  OAI21X1  g01699(.A0(new_n4114_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4135_));
  AOI21X1  g01700(.A0(new_n4134_), .A1(new_n4132_), .B0(new_n4135_), .Y(new_n4136_));
  OR2X1    g01701(.A(new_n4133_), .B(new_n3080_), .Y(new_n4137_));
  AOI21X1  g01702(.A0(new_n4113_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4138_));
  AND2X1   g01703(.A(new_n4138_), .B(new_n4137_), .Y(new_n4139_));
  NOR3X1   g01704(.A(new_n4139_), .B(new_n4136_), .C(new_n3130_), .Y(new_n4140_));
  OAI21X1  g01705(.A0(new_n4114_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4141_));
  NAND3X1  g01706(.A(new_n4126_), .B(new_n4073_), .C(new_n3104_), .Y(new_n4142_));
  AOI21X1  g01707(.A0(new_n4049_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n4143_));
  AOI21X1  g01708(.A0(new_n4143_), .A1(new_n4142_), .B0(pi0056), .Y(new_n4144_));
  OAI21X1  g01709(.A0(new_n4141_), .A1(new_n4140_), .B0(new_n4144_), .Y(new_n4145_));
  AOI21X1  g01710(.A0(new_n4110_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4146_));
  OAI21X1  g01711(.A0(new_n4127_), .A1(new_n3115_), .B0(new_n4146_), .Y(new_n4147_));
  AND2X1   g01712(.A(new_n4147_), .B(new_n3222_), .Y(new_n4148_));
  AND3X1   g01713(.A(new_n4126_), .B(new_n4073_), .C(new_n3224_), .Y(new_n4149_));
  OAI21X1  g01714(.A0(new_n4110_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4150_));
  OAI21X1  g01715(.A0(new_n4150_), .A1(new_n4149_), .B0(new_n3223_), .Y(new_n4151_));
  AOI21X1  g01716(.A0(new_n4148_), .A1(new_n4145_), .B0(new_n4151_), .Y(new_n4152_));
  OAI21X1  g01717(.A0(new_n4110_), .A1(new_n3223_), .B0(pi0247), .Y(new_n4153_));
  OAI22X1  g01718(.A0(new_n4153_), .A1(new_n4152_), .B0(new_n4103_), .B1(new_n4101_), .Y(po0160));
  AND2X1   g01719(.A(pi1138), .B(pi0215), .Y(new_n4155_));
  NOR2X1   g01720(.A(new_n4155_), .B(new_n2933_), .Y(new_n4156_));
  INVX1    g01721(.A(pi0940), .Y(new_n4157_));
  AOI21X1  g01722(.A0(new_n3145_), .A1(new_n4157_), .B0(new_n2437_), .Y(new_n4158_));
  OAI21X1  g01723(.A0(new_n3145_), .A1(pi1138), .B0(new_n4158_), .Y(new_n4159_));
  INVX1    g01724(.A(new_n4159_), .Y(new_n4160_));
  AOI21X1  g01725(.A0(pi0269), .A1(pi0216), .B0(pi0221), .Y(new_n4161_));
  INVX1    g01726(.A(pi0169), .Y(new_n4162_));
  INVX1    g01727(.A(pi0877), .Y(new_n4163_));
  OR3X1    g01728(.A(new_n3232_), .B(new_n2696_), .C(new_n4163_), .Y(new_n4164_));
  AND2X1   g01729(.A(new_n4164_), .B(new_n4162_), .Y(new_n4165_));
  MX2X1    g01730(.A(new_n4164_), .B(new_n3240_), .S0(pi0169), .Y(new_n4166_));
  AOI22X1  g01731(.A0(new_n4166_), .A1(pi0877), .B0(new_n4165_), .B1(new_n3180_), .Y(new_n4167_));
  AOI21X1  g01732(.A0(new_n2453_), .A1(pi0095), .B0(new_n4163_), .Y(new_n4168_));
  INVX1    g01733(.A(new_n4168_), .Y(new_n4169_));
  OAI21X1  g01734(.A0(new_n4162_), .A1(pi0105), .B0(pi0228), .Y(new_n4170_));
  AOI21X1  g01735(.A0(new_n4169_), .A1(pi0105), .B0(new_n4170_), .Y(new_n4171_));
  AOI21X1  g01736(.A0(new_n4171_), .A1(new_n3721_), .B0(pi0216), .Y(new_n4172_));
  OAI21X1  g01737(.A0(new_n4167_), .A1(pi0228), .B0(new_n4172_), .Y(new_n4173_));
  AOI21X1  g01738(.A0(new_n4173_), .A1(new_n4161_), .B0(new_n4160_), .Y(new_n4174_));
  OAI21X1  g01739(.A0(new_n4174_), .A1(pi0215), .B0(new_n4156_), .Y(new_n4175_));
  AND2X1   g01740(.A(pi1138), .B(pi0223), .Y(new_n4176_));
  AOI21X1  g01741(.A0(new_n3134_), .A1(new_n4157_), .B0(new_n2941_), .Y(new_n4177_));
  OAI21X1  g01742(.A0(new_n3134_), .A1(pi1138), .B0(new_n4177_), .Y(new_n4178_));
  AOI21X1  g01743(.A0(pi0269), .A1(pi0224), .B0(pi0222), .Y(new_n4179_));
  INVX1    g01744(.A(new_n4179_), .Y(new_n4180_));
  AOI21X1  g01745(.A0(new_n3232_), .A1(pi0877), .B0(pi0224), .Y(new_n4181_));
  OAI21X1  g01746(.A0(new_n4181_), .A1(new_n4180_), .B0(new_n4178_), .Y(new_n4182_));
  OR3X1    g01747(.A(new_n4182_), .B(new_n4176_), .C(pi0299), .Y(new_n4183_));
  AOI21X1  g01748(.A0(pi1138), .A1(pi0223), .B0(pi0299), .Y(new_n4184_));
  NOR2X1   g01749(.A(new_n4180_), .B(new_n3232_), .Y(new_n4185_));
  OAI21X1  g01750(.A0(new_n4185_), .A1(new_n4182_), .B0(new_n2940_), .Y(new_n4186_));
  AOI21X1  g01751(.A0(new_n4186_), .A1(new_n4184_), .B0(pi0039), .Y(new_n4187_));
  AND2X1   g01752(.A(new_n4187_), .B(new_n4183_), .Y(new_n4188_));
  AOI21X1  g01753(.A0(new_n4169_), .A1(new_n2942_), .B0(new_n4180_), .Y(new_n4189_));
  INVX1    g01754(.A(new_n4189_), .Y(new_n4190_));
  AOI21X1  g01755(.A0(new_n4190_), .A1(new_n4178_), .B0(pi0223), .Y(new_n4191_));
  OAI21X1  g01756(.A0(new_n4191_), .A1(new_n4176_), .B0(new_n2933_), .Y(new_n4192_));
  INVX1    g01757(.A(new_n4192_), .Y(new_n4193_));
  INVX1    g01758(.A(new_n4155_), .Y(new_n4194_));
  INVX1    g01759(.A(new_n4161_), .Y(new_n4195_));
  NOR2X1   g01760(.A(new_n4171_), .B(pi0216), .Y(new_n4196_));
  AOI21X1  g01761(.A0(new_n2986_), .A1(pi0169), .B0(pi0228), .Y(new_n4197_));
  OAI21X1  g01762(.A0(new_n2986_), .A1(pi0877), .B0(new_n4197_), .Y(new_n4198_));
  AOI21X1  g01763(.A0(new_n4198_), .A1(new_n4196_), .B0(new_n4195_), .Y(new_n4199_));
  OAI21X1  g01764(.A0(new_n4199_), .A1(new_n4160_), .B0(new_n2934_), .Y(new_n4200_));
  AOI21X1  g01765(.A0(new_n4200_), .A1(new_n4194_), .B0(new_n2933_), .Y(new_n4201_));
  NOR2X1   g01766(.A(new_n4201_), .B(new_n4193_), .Y(new_n4202_));
  OAI21X1  g01767(.A0(new_n4202_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n4203_));
  AOI21X1  g01768(.A0(new_n4188_), .A1(new_n4175_), .B0(new_n4203_), .Y(new_n4204_));
  INVX1    g01769(.A(pi1138), .Y(new_n4205_));
  OAI21X1  g01770(.A0(pi0228), .A1(pi0169), .B0(new_n4196_), .Y(new_n4206_));
  AOI21X1  g01771(.A0(new_n4206_), .A1(new_n4161_), .B0(new_n4160_), .Y(new_n4207_));
  MX2X1    g01772(.A(new_n4207_), .B(new_n4205_), .S0(pi0215), .Y(new_n4208_));
  INVX1    g01773(.A(new_n4208_), .Y(new_n4209_));
  AOI21X1  g01774(.A0(new_n4209_), .A1(pi0299), .B0(new_n4193_), .Y(new_n4210_));
  INVX1    g01775(.A(new_n4210_), .Y(new_n4211_));
  OAI21X1  g01776(.A0(new_n4211_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4212_));
  AOI21X1  g01777(.A0(new_n3199_), .A1(pi0169), .B0(pi0228), .Y(new_n4213_));
  OAI21X1  g01778(.A0(new_n3199_), .A1(pi0877), .B0(new_n4213_), .Y(new_n4214_));
  AOI21X1  g01779(.A0(new_n4214_), .A1(new_n4196_), .B0(new_n4195_), .Y(new_n4215_));
  OAI21X1  g01780(.A0(new_n4215_), .A1(new_n4160_), .B0(new_n2934_), .Y(new_n4216_));
  AOI21X1  g01781(.A0(new_n4216_), .A1(new_n4194_), .B0(new_n2933_), .Y(new_n4217_));
  NOR3X1   g01782(.A(new_n4217_), .B(new_n4193_), .C(new_n3060_), .Y(new_n4218_));
  OAI21X1  g01783(.A0(new_n4211_), .A1(new_n3047_), .B0(pi0100), .Y(new_n4219_));
  OAI22X1  g01784(.A0(new_n4219_), .A1(new_n4218_), .B0(new_n4212_), .B1(new_n4204_), .Y(new_n4220_));
  MX2X1    g01785(.A(new_n4210_), .B(new_n4202_), .S0(new_n3064_), .Y(new_n4221_));
  OAI21X1  g01786(.A0(new_n4221_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n4222_));
  AOI21X1  g01787(.A0(new_n4220_), .A1(new_n3131_), .B0(new_n4222_), .Y(new_n4223_));
  OAI21X1  g01788(.A0(new_n4211_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4224_));
  NAND2X1  g01789(.A(new_n4221_), .B(new_n3077_), .Y(new_n4225_));
  AOI21X1  g01790(.A0(new_n4210_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4226_));
  AOI21X1  g01791(.A0(new_n4226_), .A1(new_n4225_), .B0(new_n3130_), .Y(new_n4227_));
  OAI21X1  g01792(.A0(new_n4224_), .A1(new_n4223_), .B0(new_n4227_), .Y(new_n4228_));
  AOI21X1  g01793(.A0(new_n4210_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4229_));
  AND3X1   g01794(.A(new_n4200_), .B(new_n4194_), .C(new_n3104_), .Y(new_n4230_));
  OAI21X1  g01795(.A0(new_n4209_), .A1(new_n3104_), .B0(pi0055), .Y(new_n4231_));
  OAI21X1  g01796(.A0(new_n4231_), .A1(new_n4230_), .B0(new_n3118_), .Y(new_n4232_));
  AOI21X1  g01797(.A0(new_n4229_), .A1(new_n4228_), .B0(new_n4232_), .Y(new_n4233_));
  AOI21X1  g01798(.A0(new_n4200_), .A1(new_n4194_), .B0(new_n3115_), .Y(new_n4234_));
  OAI21X1  g01799(.A0(new_n4208_), .A1(new_n3114_), .B0(pi0056), .Y(new_n4235_));
  OAI21X1  g01800(.A0(new_n4235_), .A1(new_n4234_), .B0(new_n3222_), .Y(new_n4236_));
  NAND3X1  g01801(.A(new_n4200_), .B(new_n4194_), .C(new_n3224_), .Y(new_n4237_));
  AOI21X1  g01802(.A0(new_n4208_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n4238_));
  OR3X1    g01803(.A(pi0246), .B(pi0059), .C(pi0057), .Y(new_n4239_));
  AOI21X1  g01804(.A0(new_n4238_), .A1(new_n4237_), .B0(new_n4239_), .Y(new_n4240_));
  OAI21X1  g01805(.A0(new_n4236_), .A1(new_n4233_), .B0(new_n4240_), .Y(new_n4241_));
  INVX1    g01806(.A(new_n4156_), .Y(new_n4242_));
  OAI21X1  g01807(.A0(new_n3797_), .A1(pi0877), .B0(new_n4162_), .Y(new_n4243_));
  AOI21X1  g01808(.A0(new_n3799_), .A1(new_n4163_), .B0(new_n4162_), .Y(new_n4244_));
  OAI21X1  g01809(.A0(new_n3570_), .A1(new_n4163_), .B0(new_n4244_), .Y(new_n4245_));
  AOI21X1  g01810(.A0(new_n4245_), .A1(new_n4243_), .B0(pi0228), .Y(new_n4246_));
  OAI21X1  g01811(.A0(new_n3232_), .A1(new_n3011_), .B0(new_n4196_), .Y(new_n4247_));
  OAI21X1  g01812(.A0(new_n4247_), .A1(new_n4246_), .B0(new_n4161_), .Y(new_n4248_));
  AOI21X1  g01813(.A0(new_n4248_), .A1(new_n4159_), .B0(pi0215), .Y(new_n4249_));
  OAI21X1  g01814(.A0(new_n4249_), .A1(new_n4242_), .B0(new_n4187_), .Y(new_n4250_));
  AND2X1   g01815(.A(new_n4192_), .B(new_n3807_), .Y(new_n4251_));
  INVX1    g01816(.A(new_n4251_), .Y(new_n4252_));
  NOR3X1   g01817(.A(new_n4171_), .B(new_n3254_), .C(pi0216), .Y(new_n4253_));
  AOI21X1  g01818(.A0(new_n4253_), .A1(new_n4198_), .B0(new_n4195_), .Y(new_n4254_));
  OAI21X1  g01819(.A0(new_n4254_), .A1(new_n4160_), .B0(new_n2934_), .Y(new_n4255_));
  AOI21X1  g01820(.A0(new_n4255_), .A1(new_n4194_), .B0(new_n2933_), .Y(new_n4256_));
  NOR2X1   g01821(.A(new_n4256_), .B(new_n4252_), .Y(new_n4257_));
  INVX1    g01822(.A(new_n4257_), .Y(new_n4258_));
  AOI21X1  g01823(.A0(new_n4258_), .A1(pi0039), .B0(pi0038), .Y(new_n4259_));
  INVX1    g01824(.A(pi0269), .Y(new_n4260_));
  OAI21X1  g01825(.A0(new_n4260_), .A1(new_n2438_), .B0(new_n3339_), .Y(new_n4261_));
  AND2X1   g01826(.A(new_n4261_), .B(new_n4208_), .Y(new_n4262_));
  INVX1    g01827(.A(new_n4262_), .Y(new_n4263_));
  AOI21X1  g01828(.A0(new_n4263_), .A1(pi0299), .B0(new_n4252_), .Y(new_n4264_));
  INVX1    g01829(.A(new_n4264_), .Y(new_n4265_));
  OAI21X1  g01830(.A0(new_n4265_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4266_));
  AOI21X1  g01831(.A0(new_n4259_), .A1(new_n4250_), .B0(new_n4266_), .Y(new_n4267_));
  AND2X1   g01832(.A(new_n4253_), .B(new_n4214_), .Y(new_n4268_));
  OAI21X1  g01833(.A0(new_n4268_), .A1(new_n4195_), .B0(new_n4159_), .Y(new_n4269_));
  AOI21X1  g01834(.A0(new_n4269_), .A1(new_n2934_), .B0(new_n4155_), .Y(new_n4270_));
  AND3X1   g01835(.A(new_n4192_), .B(new_n3807_), .C(new_n3047_), .Y(new_n4271_));
  OAI21X1  g01836(.A0(new_n4270_), .A1(new_n2933_), .B0(new_n4271_), .Y(new_n4272_));
  AOI21X1  g01837(.A0(new_n4264_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4273_));
  AND2X1   g01838(.A(new_n4273_), .B(new_n4272_), .Y(new_n4274_));
  OAI21X1  g01839(.A0(new_n4274_), .A1(new_n4267_), .B0(new_n3131_), .Y(new_n4275_));
  MX2X1    g01840(.A(new_n4265_), .B(new_n4258_), .S0(new_n3064_), .Y(new_n4276_));
  AOI21X1  g01841(.A0(new_n4276_), .A1(pi0087), .B0(pi0075), .Y(new_n4277_));
  OAI21X1  g01842(.A0(new_n4265_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4278_));
  AOI21X1  g01843(.A0(new_n4277_), .A1(new_n4275_), .B0(new_n4278_), .Y(new_n4279_));
  AOI21X1  g01844(.A0(new_n4264_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4280_));
  OAI21X1  g01845(.A0(new_n4276_), .A1(new_n3080_), .B0(new_n4280_), .Y(new_n4281_));
  NAND2X1  g01846(.A(new_n4281_), .B(new_n3102_), .Y(new_n4282_));
  OR2X1    g01847(.A(new_n4282_), .B(new_n4279_), .Y(new_n4283_));
  AOI21X1  g01848(.A0(new_n4264_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4284_));
  AND3X1   g01849(.A(new_n4255_), .B(new_n4194_), .C(new_n3104_), .Y(new_n4285_));
  OAI21X1  g01850(.A0(new_n4263_), .A1(new_n3104_), .B0(pi0055), .Y(new_n4286_));
  OAI21X1  g01851(.A0(new_n4286_), .A1(new_n4285_), .B0(new_n3118_), .Y(new_n4287_));
  AOI21X1  g01852(.A0(new_n4284_), .A1(new_n4283_), .B0(new_n4287_), .Y(new_n4288_));
  AOI21X1  g01853(.A0(new_n4255_), .A1(new_n4194_), .B0(new_n3115_), .Y(new_n4289_));
  OAI21X1  g01854(.A0(new_n4262_), .A1(new_n3114_), .B0(pi0056), .Y(new_n4290_));
  OAI21X1  g01855(.A0(new_n4290_), .A1(new_n4289_), .B0(new_n3222_), .Y(new_n4291_));
  NAND3X1  g01856(.A(new_n4255_), .B(new_n4194_), .C(new_n3224_), .Y(new_n4292_));
  AOI21X1  g01857(.A0(new_n4262_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n4293_));
  NAND2X1  g01858(.A(new_n3223_), .B(pi0246), .Y(new_n4294_));
  AOI21X1  g01859(.A0(new_n4293_), .A1(new_n4292_), .B0(new_n4294_), .Y(new_n4295_));
  OAI21X1  g01860(.A0(new_n4291_), .A1(new_n4288_), .B0(new_n4295_), .Y(new_n4296_));
  NAND2X1  g01861(.A(pi0269), .B(pi0216), .Y(new_n4297_));
  NAND4X1  g01862(.A(new_n4297_), .B(new_n3254_), .C(new_n3018_), .D(pi0246), .Y(new_n4298_));
  NAND3X1  g01863(.A(new_n4298_), .B(new_n4208_), .C(new_n3374_), .Y(new_n4299_));
  AND3X1   g01864(.A(new_n4299_), .B(new_n4296_), .C(new_n4241_), .Y(po0161));
  AND2X1   g01865(.A(pi1137), .B(pi0215), .Y(new_n4301_));
  NOR2X1   g01866(.A(new_n4301_), .B(new_n2933_), .Y(new_n4302_));
  INVX1    g01867(.A(pi0933), .Y(new_n4303_));
  AOI21X1  g01868(.A0(new_n3145_), .A1(new_n4303_), .B0(new_n2437_), .Y(new_n4304_));
  OAI21X1  g01869(.A0(new_n3145_), .A1(pi1137), .B0(new_n4304_), .Y(new_n4305_));
  INVX1    g01870(.A(new_n4305_), .Y(new_n4306_));
  AOI21X1  g01871(.A0(pi0280), .A1(pi0216), .B0(pi0221), .Y(new_n4307_));
  INVX1    g01872(.A(pi0168), .Y(new_n4308_));
  INVX1    g01873(.A(pi0878), .Y(new_n4309_));
  OR3X1    g01874(.A(new_n3232_), .B(new_n2696_), .C(new_n4309_), .Y(new_n4310_));
  AND2X1   g01875(.A(new_n4310_), .B(new_n4308_), .Y(new_n4311_));
  MX2X1    g01876(.A(new_n4310_), .B(new_n3240_), .S0(pi0168), .Y(new_n4312_));
  AOI22X1  g01877(.A0(new_n4312_), .A1(pi0878), .B0(new_n4311_), .B1(new_n3180_), .Y(new_n4313_));
  AOI21X1  g01878(.A0(new_n2453_), .A1(pi0095), .B0(new_n4309_), .Y(new_n4314_));
  INVX1    g01879(.A(new_n4314_), .Y(new_n4315_));
  OAI21X1  g01880(.A0(new_n4308_), .A1(pi0105), .B0(pi0228), .Y(new_n4316_));
  AOI21X1  g01881(.A0(new_n4315_), .A1(pi0105), .B0(new_n4316_), .Y(new_n4317_));
  AOI21X1  g01882(.A0(new_n4317_), .A1(new_n3721_), .B0(pi0216), .Y(new_n4318_));
  OAI21X1  g01883(.A0(new_n4313_), .A1(pi0228), .B0(new_n4318_), .Y(new_n4319_));
  AOI21X1  g01884(.A0(new_n4319_), .A1(new_n4307_), .B0(new_n4306_), .Y(new_n4320_));
  OAI21X1  g01885(.A0(new_n4320_), .A1(pi0215), .B0(new_n4302_), .Y(new_n4321_));
  AND2X1   g01886(.A(pi1137), .B(pi0223), .Y(new_n4322_));
  AOI21X1  g01887(.A0(new_n3134_), .A1(new_n4303_), .B0(new_n2941_), .Y(new_n4323_));
  OAI21X1  g01888(.A0(new_n3134_), .A1(pi1137), .B0(new_n4323_), .Y(new_n4324_));
  AOI21X1  g01889(.A0(pi0280), .A1(pi0224), .B0(pi0222), .Y(new_n4325_));
  INVX1    g01890(.A(new_n4325_), .Y(new_n4326_));
  AOI21X1  g01891(.A0(new_n3232_), .A1(pi0878), .B0(pi0224), .Y(new_n4327_));
  OAI21X1  g01892(.A0(new_n4327_), .A1(new_n4326_), .B0(new_n4324_), .Y(new_n4328_));
  OR3X1    g01893(.A(new_n4328_), .B(new_n4322_), .C(pi0299), .Y(new_n4329_));
  AOI21X1  g01894(.A0(pi1137), .A1(pi0223), .B0(pi0299), .Y(new_n4330_));
  NOR2X1   g01895(.A(new_n4326_), .B(new_n3232_), .Y(new_n4331_));
  OAI21X1  g01896(.A0(new_n4331_), .A1(new_n4328_), .B0(new_n2940_), .Y(new_n4332_));
  AOI21X1  g01897(.A0(new_n4332_), .A1(new_n4330_), .B0(pi0039), .Y(new_n4333_));
  AND2X1   g01898(.A(new_n4333_), .B(new_n4329_), .Y(new_n4334_));
  AOI21X1  g01899(.A0(new_n4315_), .A1(new_n2942_), .B0(new_n4326_), .Y(new_n4335_));
  INVX1    g01900(.A(new_n4335_), .Y(new_n4336_));
  AOI21X1  g01901(.A0(new_n4336_), .A1(new_n4324_), .B0(pi0223), .Y(new_n4337_));
  OAI21X1  g01902(.A0(new_n4337_), .A1(new_n4322_), .B0(new_n2933_), .Y(new_n4338_));
  INVX1    g01903(.A(new_n4338_), .Y(new_n4339_));
  INVX1    g01904(.A(new_n4301_), .Y(new_n4340_));
  INVX1    g01905(.A(new_n4307_), .Y(new_n4341_));
  NOR2X1   g01906(.A(new_n4317_), .B(pi0216), .Y(new_n4342_));
  AOI21X1  g01907(.A0(new_n2986_), .A1(pi0168), .B0(pi0228), .Y(new_n4343_));
  OAI21X1  g01908(.A0(new_n2986_), .A1(pi0878), .B0(new_n4343_), .Y(new_n4344_));
  AOI21X1  g01909(.A0(new_n4344_), .A1(new_n4342_), .B0(new_n4341_), .Y(new_n4345_));
  OAI21X1  g01910(.A0(new_n4345_), .A1(new_n4306_), .B0(new_n2934_), .Y(new_n4346_));
  AOI21X1  g01911(.A0(new_n4346_), .A1(new_n4340_), .B0(new_n2933_), .Y(new_n4347_));
  NOR2X1   g01912(.A(new_n4347_), .B(new_n4339_), .Y(new_n4348_));
  OAI21X1  g01913(.A0(new_n4348_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n4349_));
  AOI21X1  g01914(.A0(new_n4334_), .A1(new_n4321_), .B0(new_n4349_), .Y(new_n4350_));
  INVX1    g01915(.A(pi1137), .Y(new_n4351_));
  OAI21X1  g01916(.A0(pi0228), .A1(pi0168), .B0(new_n4342_), .Y(new_n4352_));
  AOI21X1  g01917(.A0(new_n4352_), .A1(new_n4307_), .B0(new_n4306_), .Y(new_n4353_));
  MX2X1    g01918(.A(new_n4353_), .B(new_n4351_), .S0(pi0215), .Y(new_n4354_));
  INVX1    g01919(.A(new_n4354_), .Y(new_n4355_));
  AOI21X1  g01920(.A0(new_n4355_), .A1(pi0299), .B0(new_n4339_), .Y(new_n4356_));
  INVX1    g01921(.A(new_n4356_), .Y(new_n4357_));
  OAI21X1  g01922(.A0(new_n4357_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4358_));
  AOI21X1  g01923(.A0(new_n3199_), .A1(pi0168), .B0(pi0228), .Y(new_n4359_));
  OAI21X1  g01924(.A0(new_n3199_), .A1(pi0878), .B0(new_n4359_), .Y(new_n4360_));
  AOI21X1  g01925(.A0(new_n4360_), .A1(new_n4342_), .B0(new_n4341_), .Y(new_n4361_));
  OAI21X1  g01926(.A0(new_n4361_), .A1(new_n4306_), .B0(new_n2934_), .Y(new_n4362_));
  AOI21X1  g01927(.A0(new_n4362_), .A1(new_n4340_), .B0(new_n2933_), .Y(new_n4363_));
  NOR3X1   g01928(.A(new_n4363_), .B(new_n4339_), .C(new_n3060_), .Y(new_n4364_));
  OAI21X1  g01929(.A0(new_n4357_), .A1(new_n3047_), .B0(pi0100), .Y(new_n4365_));
  OAI22X1  g01930(.A0(new_n4365_), .A1(new_n4364_), .B0(new_n4358_), .B1(new_n4350_), .Y(new_n4366_));
  MX2X1    g01931(.A(new_n4356_), .B(new_n4348_), .S0(new_n3064_), .Y(new_n4367_));
  OAI21X1  g01932(.A0(new_n4367_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n4368_));
  AOI21X1  g01933(.A0(new_n4366_), .A1(new_n3131_), .B0(new_n4368_), .Y(new_n4369_));
  OAI21X1  g01934(.A0(new_n4357_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4370_));
  NAND2X1  g01935(.A(new_n4367_), .B(new_n3077_), .Y(new_n4371_));
  AOI21X1  g01936(.A0(new_n4356_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4372_));
  AOI21X1  g01937(.A0(new_n4372_), .A1(new_n4371_), .B0(new_n3130_), .Y(new_n4373_));
  OAI21X1  g01938(.A0(new_n4370_), .A1(new_n4369_), .B0(new_n4373_), .Y(new_n4374_));
  AOI21X1  g01939(.A0(new_n4356_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4375_));
  AND3X1   g01940(.A(new_n4346_), .B(new_n4340_), .C(new_n3104_), .Y(new_n4376_));
  OAI21X1  g01941(.A0(new_n4355_), .A1(new_n3104_), .B0(pi0055), .Y(new_n4377_));
  OAI21X1  g01942(.A0(new_n4377_), .A1(new_n4376_), .B0(new_n3118_), .Y(new_n4378_));
  AOI21X1  g01943(.A0(new_n4375_), .A1(new_n4374_), .B0(new_n4378_), .Y(new_n4379_));
  AOI21X1  g01944(.A0(new_n4346_), .A1(new_n4340_), .B0(new_n3115_), .Y(new_n4380_));
  OAI21X1  g01945(.A0(new_n4354_), .A1(new_n3114_), .B0(pi0056), .Y(new_n4381_));
  OAI21X1  g01946(.A0(new_n4381_), .A1(new_n4380_), .B0(new_n3222_), .Y(new_n4382_));
  NAND3X1  g01947(.A(new_n4346_), .B(new_n4340_), .C(new_n3224_), .Y(new_n4383_));
  AOI21X1  g01948(.A0(new_n4354_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n4384_));
  OR3X1    g01949(.A(pi0240), .B(pi0059), .C(pi0057), .Y(new_n4385_));
  AOI21X1  g01950(.A0(new_n4384_), .A1(new_n4383_), .B0(new_n4385_), .Y(new_n4386_));
  OAI21X1  g01951(.A0(new_n4382_), .A1(new_n4379_), .B0(new_n4386_), .Y(new_n4387_));
  INVX1    g01952(.A(new_n4302_), .Y(new_n4388_));
  OAI21X1  g01953(.A0(new_n3797_), .A1(pi0878), .B0(new_n4308_), .Y(new_n4389_));
  AOI21X1  g01954(.A0(new_n3799_), .A1(new_n4309_), .B0(new_n4308_), .Y(new_n4390_));
  OAI21X1  g01955(.A0(new_n3570_), .A1(new_n4309_), .B0(new_n4390_), .Y(new_n4391_));
  AOI21X1  g01956(.A0(new_n4391_), .A1(new_n4389_), .B0(pi0228), .Y(new_n4392_));
  OAI21X1  g01957(.A0(new_n3232_), .A1(new_n3011_), .B0(new_n4342_), .Y(new_n4393_));
  OAI21X1  g01958(.A0(new_n4393_), .A1(new_n4392_), .B0(new_n4307_), .Y(new_n4394_));
  AOI21X1  g01959(.A0(new_n4394_), .A1(new_n4305_), .B0(pi0215), .Y(new_n4395_));
  OAI21X1  g01960(.A0(new_n4395_), .A1(new_n4388_), .B0(new_n4333_), .Y(new_n4396_));
  AND2X1   g01961(.A(new_n4338_), .B(new_n3807_), .Y(new_n4397_));
  INVX1    g01962(.A(new_n4397_), .Y(new_n4398_));
  NOR3X1   g01963(.A(new_n4317_), .B(new_n3254_), .C(pi0216), .Y(new_n4399_));
  AOI21X1  g01964(.A0(new_n4399_), .A1(new_n4344_), .B0(new_n4341_), .Y(new_n4400_));
  OAI21X1  g01965(.A0(new_n4400_), .A1(new_n4306_), .B0(new_n2934_), .Y(new_n4401_));
  AOI21X1  g01966(.A0(new_n4401_), .A1(new_n4340_), .B0(new_n2933_), .Y(new_n4402_));
  NOR2X1   g01967(.A(new_n4402_), .B(new_n4398_), .Y(new_n4403_));
  INVX1    g01968(.A(new_n4403_), .Y(new_n4404_));
  AOI21X1  g01969(.A0(new_n4404_), .A1(pi0039), .B0(pi0038), .Y(new_n4405_));
  INVX1    g01970(.A(pi0280), .Y(new_n4406_));
  OAI21X1  g01971(.A0(new_n4406_), .A1(new_n2438_), .B0(new_n3339_), .Y(new_n4407_));
  AND2X1   g01972(.A(new_n4407_), .B(new_n4354_), .Y(new_n4408_));
  INVX1    g01973(.A(new_n4408_), .Y(new_n4409_));
  AOI21X1  g01974(.A0(new_n4409_), .A1(pi0299), .B0(new_n4398_), .Y(new_n4410_));
  INVX1    g01975(.A(new_n4410_), .Y(new_n4411_));
  OAI21X1  g01976(.A0(new_n4411_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4412_));
  AOI21X1  g01977(.A0(new_n4405_), .A1(new_n4396_), .B0(new_n4412_), .Y(new_n4413_));
  AND2X1   g01978(.A(new_n4399_), .B(new_n4360_), .Y(new_n4414_));
  OAI21X1  g01979(.A0(new_n4414_), .A1(new_n4341_), .B0(new_n4305_), .Y(new_n4415_));
  AOI21X1  g01980(.A0(new_n4415_), .A1(new_n2934_), .B0(new_n4301_), .Y(new_n4416_));
  AND3X1   g01981(.A(new_n4338_), .B(new_n3807_), .C(new_n3047_), .Y(new_n4417_));
  OAI21X1  g01982(.A0(new_n4416_), .A1(new_n2933_), .B0(new_n4417_), .Y(new_n4418_));
  AOI21X1  g01983(.A0(new_n4410_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4419_));
  AND2X1   g01984(.A(new_n4419_), .B(new_n4418_), .Y(new_n4420_));
  OAI21X1  g01985(.A0(new_n4420_), .A1(new_n4413_), .B0(new_n3131_), .Y(new_n4421_));
  MX2X1    g01986(.A(new_n4411_), .B(new_n4404_), .S0(new_n3064_), .Y(new_n4422_));
  AOI21X1  g01987(.A0(new_n4422_), .A1(pi0087), .B0(pi0075), .Y(new_n4423_));
  OAI21X1  g01988(.A0(new_n4411_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4424_));
  AOI21X1  g01989(.A0(new_n4423_), .A1(new_n4421_), .B0(new_n4424_), .Y(new_n4425_));
  AOI21X1  g01990(.A0(new_n4410_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4426_));
  OAI21X1  g01991(.A0(new_n4422_), .A1(new_n3080_), .B0(new_n4426_), .Y(new_n4427_));
  NAND2X1  g01992(.A(new_n4427_), .B(new_n3102_), .Y(new_n4428_));
  OR2X1    g01993(.A(new_n4428_), .B(new_n4425_), .Y(new_n4429_));
  AOI21X1  g01994(.A0(new_n4410_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4430_));
  AND3X1   g01995(.A(new_n4401_), .B(new_n4340_), .C(new_n3104_), .Y(new_n4431_));
  OAI21X1  g01996(.A0(new_n4409_), .A1(new_n3104_), .B0(pi0055), .Y(new_n4432_));
  OAI21X1  g01997(.A0(new_n4432_), .A1(new_n4431_), .B0(new_n3118_), .Y(new_n4433_));
  AOI21X1  g01998(.A0(new_n4430_), .A1(new_n4429_), .B0(new_n4433_), .Y(new_n4434_));
  AOI21X1  g01999(.A0(new_n4401_), .A1(new_n4340_), .B0(new_n3115_), .Y(new_n4435_));
  OAI21X1  g02000(.A0(new_n4408_), .A1(new_n3114_), .B0(pi0056), .Y(new_n4436_));
  OAI21X1  g02001(.A0(new_n4436_), .A1(new_n4435_), .B0(new_n3222_), .Y(new_n4437_));
  NAND3X1  g02002(.A(new_n4401_), .B(new_n4340_), .C(new_n3224_), .Y(new_n4438_));
  AOI21X1  g02003(.A0(new_n4408_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n4439_));
  NAND2X1  g02004(.A(new_n3223_), .B(pi0240), .Y(new_n4440_));
  AOI21X1  g02005(.A0(new_n4439_), .A1(new_n4438_), .B0(new_n4440_), .Y(new_n4441_));
  OAI21X1  g02006(.A0(new_n4437_), .A1(new_n4434_), .B0(new_n4441_), .Y(new_n4442_));
  INVX1    g02007(.A(pi0240), .Y(new_n4443_));
  OR2X1    g02008(.A(new_n4407_), .B(new_n4443_), .Y(new_n4444_));
  NAND3X1  g02009(.A(new_n4444_), .B(new_n4354_), .C(new_n3374_), .Y(new_n4445_));
  AND3X1   g02010(.A(new_n4445_), .B(new_n4442_), .C(new_n4387_), .Y(po0162));
  INVX1    g02011(.A(pi0928), .Y(new_n4447_));
  AOI21X1  g02012(.A0(new_n3145_), .A1(new_n4447_), .B0(new_n2437_), .Y(new_n4448_));
  OAI21X1  g02013(.A0(new_n3145_), .A1(pi1136), .B0(new_n4448_), .Y(new_n4449_));
  AND2X1   g02014(.A(pi0266), .B(pi0216), .Y(new_n4450_));
  NOR2X1   g02015(.A(new_n3243_), .B(new_n2793_), .Y(new_n4451_));
  INVX1    g02016(.A(new_n4451_), .Y(new_n4452_));
  INVX1    g02017(.A(pi0875), .Y(new_n4453_));
  AOI21X1  g02018(.A0(new_n2453_), .A1(pi0095), .B0(new_n4453_), .Y(new_n4454_));
  MX2X1    g02019(.A(new_n4454_), .B(pi0166), .S0(new_n2447_), .Y(new_n4455_));
  INVX1    g02020(.A(new_n4455_), .Y(new_n4456_));
  AOI21X1  g02021(.A0(new_n4456_), .A1(new_n4451_), .B0(pi0216), .Y(new_n4457_));
  INVX1    g02022(.A(new_n4457_), .Y(new_n4458_));
  INVX1    g02023(.A(pi0166), .Y(new_n4459_));
  OAI21X1  g02024(.A0(new_n3799_), .A1(new_n4459_), .B0(pi0875), .Y(new_n4460_));
  AOI21X1  g02025(.A0(new_n3797_), .A1(new_n4459_), .B0(new_n4460_), .Y(new_n4461_));
  AND3X1   g02026(.A(new_n3180_), .B(new_n4453_), .C(pi0166), .Y(new_n4462_));
  OAI21X1  g02027(.A0(new_n4462_), .A1(new_n4461_), .B0(new_n2793_), .Y(new_n4463_));
  AOI21X1  g02028(.A0(new_n4463_), .A1(new_n4452_), .B0(new_n4458_), .Y(new_n4464_));
  OAI21X1  g02029(.A0(new_n4464_), .A1(new_n4450_), .B0(new_n2437_), .Y(new_n4465_));
  AOI21X1  g02030(.A0(new_n4465_), .A1(new_n4449_), .B0(pi0215), .Y(new_n4466_));
  AND2X1   g02031(.A(pi1136), .B(pi0215), .Y(new_n4467_));
  OR2X1    g02032(.A(new_n4467_), .B(new_n2933_), .Y(new_n4468_));
  OR3X1    g02033(.A(new_n2454_), .B(pi0875), .C(pi0224), .Y(new_n4469_));
  INVX1    g02034(.A(pi0266), .Y(new_n4470_));
  AOI21X1  g02035(.A0(new_n4470_), .A1(pi0224), .B0(pi0222), .Y(new_n4471_));
  AND2X1   g02036(.A(new_n4471_), .B(new_n4469_), .Y(new_n4472_));
  OAI21X1  g02037(.A0(new_n3231_), .A1(new_n2454_), .B0(new_n2951_), .Y(new_n4473_));
  NAND2X1  g02038(.A(new_n4473_), .B(new_n4472_), .Y(new_n4474_));
  AOI21X1  g02039(.A0(new_n3134_), .A1(new_n4447_), .B0(new_n2941_), .Y(new_n4475_));
  OAI21X1  g02040(.A0(new_n3134_), .A1(pi1136), .B0(new_n4475_), .Y(new_n4476_));
  AOI21X1  g02041(.A0(pi1136), .A1(pi0223), .B0(pi0299), .Y(new_n4477_));
  AND2X1   g02042(.A(new_n4477_), .B(new_n4476_), .Y(new_n4478_));
  INVX1    g02043(.A(new_n4477_), .Y(new_n4479_));
  INVX1    g02044(.A(new_n4472_), .Y(new_n4480_));
  AND2X1   g02045(.A(new_n4476_), .B(new_n4480_), .Y(new_n4481_));
  AOI21X1  g02046(.A0(new_n4481_), .A1(new_n4473_), .B0(pi0223), .Y(new_n4482_));
  OAI21X1  g02047(.A0(new_n4482_), .A1(new_n4479_), .B0(new_n2939_), .Y(new_n4483_));
  AOI21X1  g02048(.A0(new_n4478_), .A1(new_n4474_), .B0(new_n4483_), .Y(new_n4484_));
  OAI21X1  g02049(.A0(new_n4468_), .A1(new_n4466_), .B0(new_n4484_), .Y(new_n4485_));
  AND2X1   g02050(.A(pi1136), .B(pi0223), .Y(new_n4486_));
  AOI21X1  g02051(.A0(new_n4476_), .A1(new_n4480_), .B0(pi0223), .Y(new_n4487_));
  OAI21X1  g02052(.A0(new_n4487_), .A1(new_n4486_), .B0(new_n2933_), .Y(new_n4488_));
  INVX1    g02053(.A(new_n4488_), .Y(new_n4489_));
  OAI21X1  g02054(.A0(new_n4454_), .A1(new_n2991_), .B0(new_n4489_), .Y(new_n4490_));
  AND2X1   g02055(.A(new_n4455_), .B(pi0228), .Y(new_n4491_));
  INVX1    g02056(.A(new_n4491_), .Y(new_n4492_));
  AOI21X1  g02057(.A0(new_n2987_), .A1(new_n4453_), .B0(pi0228), .Y(new_n4493_));
  OAI21X1  g02058(.A0(new_n2987_), .A1(pi0166), .B0(new_n4493_), .Y(new_n4494_));
  AOI21X1  g02059(.A0(new_n4494_), .A1(new_n4492_), .B0(pi0216), .Y(new_n4495_));
  OAI21X1  g02060(.A0(new_n4495_), .A1(new_n4450_), .B0(new_n2437_), .Y(new_n4496_));
  AOI21X1  g02061(.A0(new_n4496_), .A1(new_n4449_), .B0(pi0215), .Y(new_n4497_));
  OAI21X1  g02062(.A0(new_n4497_), .A1(new_n4467_), .B0(pi0299), .Y(new_n4498_));
  NAND2X1  g02063(.A(new_n4498_), .B(new_n4490_), .Y(new_n4499_));
  AOI21X1  g02064(.A0(new_n4499_), .A1(pi0039), .B0(pi0038), .Y(new_n4500_));
  AOI21X1  g02065(.A0(new_n2793_), .A1(pi0166), .B0(new_n4491_), .Y(new_n4501_));
  MX2X1    g02066(.A(new_n4501_), .B(new_n4470_), .S0(pi0216), .Y(new_n4502_));
  OAI21X1  g02067(.A0(new_n4502_), .A1(pi0221), .B0(new_n4449_), .Y(new_n4503_));
  AOI21X1  g02068(.A0(new_n4503_), .A1(new_n2934_), .B0(new_n4467_), .Y(new_n4504_));
  OAI21X1  g02069(.A0(new_n4504_), .A1(new_n2933_), .B0(new_n4490_), .Y(new_n4505_));
  OAI21X1  g02070(.A0(new_n4505_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4506_));
  AOI21X1  g02071(.A0(new_n4500_), .A1(new_n4485_), .B0(new_n4506_), .Y(new_n4507_));
  AOI21X1  g02072(.A0(new_n3190_), .A1(new_n4453_), .B0(new_n4459_), .Y(new_n4508_));
  INVX1    g02073(.A(new_n4508_), .Y(new_n4509_));
  NOR2X1   g02074(.A(pi0161), .B(pi0152), .Y(new_n4510_));
  AOI21X1  g02075(.A0(new_n3195_), .A1(new_n4510_), .B0(new_n4453_), .Y(new_n4511_));
  OAI21X1  g02076(.A0(new_n3190_), .A1(new_n4510_), .B0(new_n4511_), .Y(new_n4512_));
  AOI21X1  g02077(.A0(new_n4512_), .A1(new_n4509_), .B0(pi0228), .Y(new_n4513_));
  OR2X1    g02078(.A(new_n4513_), .B(new_n4491_), .Y(new_n4514_));
  AOI21X1  g02079(.A0(new_n4514_), .A1(new_n2438_), .B0(new_n4450_), .Y(new_n4515_));
  OAI21X1  g02080(.A0(new_n4515_), .A1(pi0221), .B0(new_n4449_), .Y(new_n4516_));
  AOI21X1  g02081(.A0(new_n4516_), .A1(new_n2934_), .B0(new_n4467_), .Y(new_n4517_));
  AND2X1   g02082(.A(new_n4490_), .B(new_n3047_), .Y(new_n4518_));
  OAI21X1  g02083(.A0(new_n4517_), .A1(new_n2933_), .B0(new_n4518_), .Y(new_n4519_));
  INVX1    g02084(.A(new_n4505_), .Y(new_n4520_));
  AOI21X1  g02085(.A0(new_n4520_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4521_));
  AND2X1   g02086(.A(new_n4521_), .B(new_n4519_), .Y(new_n4522_));
  OAI21X1  g02087(.A0(new_n4522_), .A1(new_n4507_), .B0(new_n3131_), .Y(new_n4523_));
  MX2X1    g02088(.A(new_n4505_), .B(new_n4499_), .S0(new_n3064_), .Y(new_n4524_));
  AOI21X1  g02089(.A0(new_n4524_), .A1(pi0087), .B0(pi0075), .Y(new_n4525_));
  OAI21X1  g02090(.A0(new_n4505_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4526_));
  AOI21X1  g02091(.A0(new_n4525_), .A1(new_n4523_), .B0(new_n4526_), .Y(new_n4527_));
  OR2X1    g02092(.A(new_n4524_), .B(new_n3080_), .Y(new_n4528_));
  AOI21X1  g02093(.A0(new_n4520_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4529_));
  AND2X1   g02094(.A(new_n4529_), .B(new_n4528_), .Y(new_n4530_));
  NOR3X1   g02095(.A(new_n4530_), .B(new_n4527_), .C(new_n3130_), .Y(new_n4531_));
  OAI21X1  g02096(.A0(new_n4505_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4532_));
  OR3X1    g02097(.A(new_n4497_), .B(new_n4467_), .C(new_n3105_), .Y(new_n4533_));
  AOI21X1  g02098(.A0(new_n4504_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n4534_));
  AOI21X1  g02099(.A0(new_n4534_), .A1(new_n4533_), .B0(pi0056), .Y(new_n4535_));
  OAI21X1  g02100(.A0(new_n4532_), .A1(new_n4531_), .B0(new_n4535_), .Y(new_n4536_));
  OAI21X1  g02101(.A0(new_n4497_), .A1(new_n4467_), .B0(new_n3114_), .Y(new_n4537_));
  INVX1    g02102(.A(new_n4504_), .Y(new_n4538_));
  AOI21X1  g02103(.A0(new_n4538_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4539_));
  AOI21X1  g02104(.A0(new_n4539_), .A1(new_n4537_), .B0(pi0062), .Y(new_n4540_));
  NOR3X1   g02105(.A(new_n4497_), .B(new_n4467_), .C(new_n3225_), .Y(new_n4541_));
  OAI21X1  g02106(.A0(new_n4538_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4542_));
  OAI21X1  g02107(.A0(new_n4542_), .A1(new_n4541_), .B0(new_n3223_), .Y(new_n4543_));
  AOI21X1  g02108(.A0(new_n4540_), .A1(new_n4536_), .B0(new_n4543_), .Y(new_n4544_));
  INVX1    g02109(.A(pi0245), .Y(new_n4545_));
  OAI21X1  g02110(.A0(new_n4538_), .A1(new_n3223_), .B0(new_n4545_), .Y(new_n4546_));
  OAI21X1  g02111(.A0(new_n3244_), .A1(pi0166), .B0(new_n4453_), .Y(new_n4547_));
  AOI21X1  g02112(.A0(new_n3240_), .A1(pi0166), .B0(new_n4547_), .Y(new_n4548_));
  AOI21X1  g02113(.A0(new_n3180_), .A1(new_n4459_), .B0(new_n4453_), .Y(new_n4549_));
  OR3X1    g02114(.A(new_n4549_), .B(new_n4548_), .C(pi0228), .Y(new_n4550_));
  AOI21X1  g02115(.A0(new_n4550_), .A1(new_n4457_), .B0(new_n4450_), .Y(new_n4551_));
  OAI21X1  g02116(.A0(new_n4551_), .A1(pi0221), .B0(new_n4449_), .Y(new_n4552_));
  AOI21X1  g02117(.A0(new_n4552_), .A1(new_n2934_), .B0(new_n4468_), .Y(new_n4553_));
  INVX1    g02118(.A(pi1136), .Y(new_n4554_));
  INVX1    g02119(.A(new_n4449_), .Y(new_n4555_));
  INVX1    g02120(.A(new_n4450_), .Y(new_n4556_));
  AND3X1   g02121(.A(new_n4494_), .B(new_n4492_), .C(new_n3456_), .Y(new_n4557_));
  OAI21X1  g02122(.A0(new_n4557_), .A1(pi0216), .B0(new_n4556_), .Y(new_n4558_));
  AOI21X1  g02123(.A0(new_n4558_), .A1(new_n2437_), .B0(new_n4555_), .Y(new_n4559_));
  MX2X1    g02124(.A(new_n4559_), .B(new_n4554_), .S0(pi0215), .Y(new_n4560_));
  OAI21X1  g02125(.A0(new_n4560_), .A1(new_n2933_), .B0(new_n4488_), .Y(new_n4561_));
  AOI21X1  g02126(.A0(new_n4561_), .A1(pi0039), .B0(pi0038), .Y(new_n4562_));
  OAI21X1  g02127(.A0(new_n4553_), .A1(new_n4483_), .B0(new_n4562_), .Y(new_n4563_));
  AND2X1   g02128(.A(new_n4504_), .B(new_n3257_), .Y(new_n4564_));
  INVX1    g02129(.A(new_n4564_), .Y(new_n4565_));
  AOI21X1  g02130(.A0(new_n4565_), .A1(pi0299), .B0(new_n4489_), .Y(new_n4566_));
  AOI21X1  g02131(.A0(new_n4566_), .A1(pi0038), .B0(pi0100), .Y(new_n4567_));
  INVX1    g02132(.A(new_n4467_), .Y(new_n4568_));
  OR2X1    g02133(.A(new_n4491_), .B(new_n3254_), .Y(new_n4569_));
  OAI21X1  g02134(.A0(new_n4569_), .A1(new_n4513_), .B0(new_n2438_), .Y(new_n4570_));
  AOI21X1  g02135(.A0(new_n4570_), .A1(new_n4556_), .B0(pi0221), .Y(new_n4571_));
  OAI21X1  g02136(.A0(new_n4571_), .A1(new_n4555_), .B0(new_n2934_), .Y(new_n4572_));
  AOI21X1  g02137(.A0(new_n4572_), .A1(new_n4568_), .B0(new_n2933_), .Y(new_n4573_));
  OR3X1    g02138(.A(new_n4573_), .B(new_n4489_), .C(new_n3060_), .Y(new_n4574_));
  AOI21X1  g02139(.A0(new_n4566_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4575_));
  AOI22X1  g02140(.A0(new_n4575_), .A1(new_n4574_), .B0(new_n4567_), .B1(new_n4563_), .Y(new_n4576_));
  INVX1    g02141(.A(new_n4566_), .Y(new_n4577_));
  MX2X1    g02142(.A(new_n4577_), .B(new_n4561_), .S0(new_n3064_), .Y(new_n4578_));
  AOI21X1  g02143(.A0(new_n4578_), .A1(pi0087), .B0(pi0075), .Y(new_n4579_));
  OAI21X1  g02144(.A0(new_n4576_), .A1(pi0087), .B0(new_n4579_), .Y(new_n4580_));
  AOI21X1  g02145(.A0(new_n4566_), .A1(pi0075), .B0(pi0092), .Y(new_n4581_));
  NOR2X1   g02146(.A(new_n4578_), .B(new_n3080_), .Y(new_n4582_));
  OAI21X1  g02147(.A0(new_n4577_), .A1(new_n3077_), .B0(pi0092), .Y(new_n4583_));
  OAI21X1  g02148(.A0(new_n4583_), .A1(new_n4582_), .B0(new_n3102_), .Y(new_n4584_));
  AOI21X1  g02149(.A0(new_n4581_), .A1(new_n4580_), .B0(new_n4584_), .Y(new_n4585_));
  OAI21X1  g02150(.A0(new_n4577_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4586_));
  NAND2X1  g02151(.A(new_n4560_), .B(new_n3104_), .Y(new_n4587_));
  AOI21X1  g02152(.A0(new_n4564_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n4588_));
  AOI21X1  g02153(.A0(new_n4588_), .A1(new_n4587_), .B0(pi0056), .Y(new_n4589_));
  OAI21X1  g02154(.A0(new_n4586_), .A1(new_n4585_), .B0(new_n4589_), .Y(new_n4590_));
  AOI21X1  g02155(.A0(new_n4565_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4591_));
  OAI21X1  g02156(.A0(new_n4560_), .A1(new_n3115_), .B0(new_n4591_), .Y(new_n4592_));
  AND3X1   g02157(.A(new_n4592_), .B(new_n4590_), .C(new_n3222_), .Y(new_n4593_));
  OAI21X1  g02158(.A0(new_n4565_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4594_));
  AOI21X1  g02159(.A0(new_n4560_), .A1(new_n3224_), .B0(new_n4594_), .Y(new_n4595_));
  OR2X1    g02160(.A(new_n4595_), .B(new_n3374_), .Y(new_n4596_));
  AOI21X1  g02161(.A0(new_n4564_), .A1(new_n3374_), .B0(new_n4545_), .Y(new_n4597_));
  OAI21X1  g02162(.A0(new_n4596_), .A1(new_n4593_), .B0(new_n4597_), .Y(new_n4598_));
  OAI21X1  g02163(.A0(new_n4546_), .A1(new_n4544_), .B0(new_n4598_), .Y(po0163));
  AOI21X1  g02164(.A0(pi0833), .A1(new_n2438_), .B0(pi1135), .Y(new_n4600_));
  OAI21X1  g02165(.A0(new_n3299_), .A1(pi0938), .B0(pi0221), .Y(new_n4601_));
  NOR2X1   g02166(.A(new_n4601_), .B(new_n4600_), .Y(new_n4602_));
  INVX1    g02167(.A(new_n4602_), .Y(new_n4603_));
  AND2X1   g02168(.A(pi0279), .B(pi0216), .Y(new_n4604_));
  INVX1    g02169(.A(pi0879), .Y(new_n4605_));
  AOI21X1  g02170(.A0(new_n2453_), .A1(pi0095), .B0(new_n4605_), .Y(new_n4606_));
  MX2X1    g02171(.A(new_n4606_), .B(pi0161), .S0(new_n2447_), .Y(new_n4607_));
  INVX1    g02172(.A(new_n4607_), .Y(new_n4608_));
  AOI21X1  g02173(.A0(new_n4608_), .A1(new_n4451_), .B0(pi0216), .Y(new_n4609_));
  INVX1    g02174(.A(new_n4609_), .Y(new_n4610_));
  INVX1    g02175(.A(pi0161), .Y(new_n4611_));
  OAI21X1  g02176(.A0(new_n3799_), .A1(new_n4611_), .B0(pi0879), .Y(new_n4612_));
  AOI21X1  g02177(.A0(new_n3797_), .A1(new_n4611_), .B0(new_n4612_), .Y(new_n4613_));
  AND3X1   g02178(.A(new_n3180_), .B(new_n4605_), .C(pi0161), .Y(new_n4614_));
  OAI21X1  g02179(.A0(new_n4614_), .A1(new_n4613_), .B0(new_n2793_), .Y(new_n4615_));
  AOI21X1  g02180(.A0(new_n4615_), .A1(new_n4452_), .B0(new_n4610_), .Y(new_n4616_));
  OAI21X1  g02181(.A0(new_n4616_), .A1(new_n4604_), .B0(new_n2437_), .Y(new_n4617_));
  AOI21X1  g02182(.A0(new_n4617_), .A1(new_n4603_), .B0(pi0215), .Y(new_n4618_));
  AND2X1   g02183(.A(pi1135), .B(pi0215), .Y(new_n4619_));
  OR2X1    g02184(.A(new_n4619_), .B(new_n2933_), .Y(new_n4620_));
  AOI21X1  g02185(.A0(pi1135), .A1(pi0223), .B0(pi0299), .Y(new_n4621_));
  INVX1    g02186(.A(pi1135), .Y(new_n4622_));
  OAI21X1  g02187(.A0(new_n3310_), .A1(pi0938), .B0(pi0222), .Y(new_n4623_));
  AOI21X1  g02188(.A0(new_n3310_), .A1(new_n4622_), .B0(new_n4623_), .Y(new_n4624_));
  OR3X1    g02189(.A(new_n2454_), .B(pi0879), .C(pi0224), .Y(new_n4625_));
  INVX1    g02190(.A(pi0279), .Y(new_n4626_));
  AOI21X1  g02191(.A0(new_n4626_), .A1(pi0224), .B0(pi0222), .Y(new_n4627_));
  AOI21X1  g02192(.A0(new_n4627_), .A1(new_n4625_), .B0(new_n4624_), .Y(new_n4628_));
  NOR2X1   g02193(.A(new_n4628_), .B(pi0223), .Y(new_n4629_));
  OAI21X1  g02194(.A0(new_n4624_), .A1(new_n4473_), .B0(new_n4629_), .Y(new_n4630_));
  AOI21X1  g02195(.A0(new_n4630_), .A1(new_n4621_), .B0(pi0039), .Y(new_n4631_));
  OAI21X1  g02196(.A0(new_n4620_), .A1(new_n4618_), .B0(new_n4631_), .Y(new_n4632_));
  AND2X1   g02197(.A(pi1135), .B(pi0223), .Y(new_n4633_));
  OAI21X1  g02198(.A0(new_n4629_), .A1(new_n4633_), .B0(new_n2933_), .Y(new_n4634_));
  INVX1    g02199(.A(new_n4634_), .Y(new_n4635_));
  OAI21X1  g02200(.A0(new_n4606_), .A1(new_n2991_), .B0(new_n4635_), .Y(new_n4636_));
  AND2X1   g02201(.A(new_n4607_), .B(pi0228), .Y(new_n4637_));
  INVX1    g02202(.A(new_n4637_), .Y(new_n4638_));
  AND2X1   g02203(.A(new_n2793_), .B(pi0161), .Y(new_n4639_));
  OAI22X1  g02204(.A0(new_n4639_), .A1(new_n3603_), .B0(new_n2986_), .B1(pi0879), .Y(new_n4640_));
  AOI21X1  g02205(.A0(new_n4640_), .A1(new_n4638_), .B0(pi0216), .Y(new_n4641_));
  OAI21X1  g02206(.A0(new_n4641_), .A1(new_n4604_), .B0(new_n2437_), .Y(new_n4642_));
  AOI21X1  g02207(.A0(new_n4642_), .A1(new_n4603_), .B0(pi0215), .Y(new_n4643_));
  OAI21X1  g02208(.A0(new_n4643_), .A1(new_n4619_), .B0(pi0299), .Y(new_n4644_));
  NAND2X1  g02209(.A(new_n4644_), .B(new_n4636_), .Y(new_n4645_));
  AOI21X1  g02210(.A0(new_n4645_), .A1(pi0039), .B0(pi0038), .Y(new_n4646_));
  AOI21X1  g02211(.A0(new_n4607_), .A1(pi0228), .B0(new_n4639_), .Y(new_n4647_));
  MX2X1    g02212(.A(new_n4647_), .B(new_n4626_), .S0(pi0216), .Y(new_n4648_));
  OAI22X1  g02213(.A0(new_n4648_), .A1(pi0221), .B0(new_n4601_), .B1(new_n4600_), .Y(new_n4649_));
  AOI21X1  g02214(.A0(new_n4649_), .A1(new_n2934_), .B0(new_n4619_), .Y(new_n4650_));
  OAI21X1  g02215(.A0(new_n4650_), .A1(new_n2933_), .B0(new_n4636_), .Y(new_n4651_));
  OAI21X1  g02216(.A0(new_n4651_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4652_));
  AOI21X1  g02217(.A0(new_n4646_), .A1(new_n4632_), .B0(new_n4652_), .Y(new_n4653_));
  AOI21X1  g02218(.A0(new_n3190_), .A1(new_n4605_), .B0(new_n4611_), .Y(new_n4654_));
  INVX1    g02219(.A(new_n4654_), .Y(new_n4655_));
  NOR2X1   g02220(.A(pi0166), .B(pi0152), .Y(new_n4656_));
  AOI21X1  g02221(.A0(new_n4656_), .A1(new_n3195_), .B0(new_n4605_), .Y(new_n4657_));
  OAI21X1  g02222(.A0(new_n4656_), .A1(new_n3190_), .B0(new_n4657_), .Y(new_n4658_));
  AOI21X1  g02223(.A0(new_n4658_), .A1(new_n4655_), .B0(pi0228), .Y(new_n4659_));
  OR2X1    g02224(.A(new_n4659_), .B(new_n4637_), .Y(new_n4660_));
  AOI21X1  g02225(.A0(new_n4660_), .A1(new_n2438_), .B0(new_n4604_), .Y(new_n4661_));
  OAI21X1  g02226(.A0(new_n4661_), .A1(pi0221), .B0(new_n4603_), .Y(new_n4662_));
  AOI21X1  g02227(.A0(new_n4662_), .A1(new_n2934_), .B0(new_n4619_), .Y(new_n4663_));
  AND2X1   g02228(.A(new_n4636_), .B(new_n3047_), .Y(new_n4664_));
  OAI21X1  g02229(.A0(new_n4663_), .A1(new_n2933_), .B0(new_n4664_), .Y(new_n4665_));
  INVX1    g02230(.A(new_n4651_), .Y(new_n4666_));
  AOI21X1  g02231(.A0(new_n4666_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4667_));
  AND2X1   g02232(.A(new_n4667_), .B(new_n4665_), .Y(new_n4668_));
  OAI21X1  g02233(.A0(new_n4668_), .A1(new_n4653_), .B0(new_n3131_), .Y(new_n4669_));
  MX2X1    g02234(.A(new_n4651_), .B(new_n4645_), .S0(new_n3064_), .Y(new_n4670_));
  AOI21X1  g02235(.A0(new_n4670_), .A1(pi0087), .B0(pi0075), .Y(new_n4671_));
  OAI21X1  g02236(.A0(new_n4651_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4672_));
  AOI21X1  g02237(.A0(new_n4671_), .A1(new_n4669_), .B0(new_n4672_), .Y(new_n4673_));
  OR2X1    g02238(.A(new_n4670_), .B(new_n3080_), .Y(new_n4674_));
  AOI21X1  g02239(.A0(new_n4666_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4675_));
  AND2X1   g02240(.A(new_n4675_), .B(new_n4674_), .Y(new_n4676_));
  NOR3X1   g02241(.A(new_n4676_), .B(new_n4673_), .C(new_n3130_), .Y(new_n4677_));
  OAI21X1  g02242(.A0(new_n4651_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4678_));
  OR3X1    g02243(.A(new_n4643_), .B(new_n4619_), .C(new_n3105_), .Y(new_n4679_));
  AOI21X1  g02244(.A0(new_n4650_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n4680_));
  AOI21X1  g02245(.A0(new_n4680_), .A1(new_n4679_), .B0(pi0056), .Y(new_n4681_));
  OAI21X1  g02246(.A0(new_n4678_), .A1(new_n4677_), .B0(new_n4681_), .Y(new_n4682_));
  OAI21X1  g02247(.A0(new_n4643_), .A1(new_n4619_), .B0(new_n3114_), .Y(new_n4683_));
  INVX1    g02248(.A(new_n4650_), .Y(new_n4684_));
  AOI21X1  g02249(.A0(new_n4684_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4685_));
  AOI21X1  g02250(.A0(new_n4685_), .A1(new_n4683_), .B0(pi0062), .Y(new_n4686_));
  NOR3X1   g02251(.A(new_n4643_), .B(new_n4619_), .C(new_n3225_), .Y(new_n4687_));
  OAI21X1  g02252(.A0(new_n4684_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4688_));
  OAI21X1  g02253(.A0(new_n4688_), .A1(new_n4687_), .B0(new_n3223_), .Y(new_n4689_));
  AOI21X1  g02254(.A0(new_n4686_), .A1(new_n4682_), .B0(new_n4689_), .Y(new_n4690_));
  INVX1    g02255(.A(pi0244), .Y(new_n4691_));
  OAI21X1  g02256(.A0(new_n4684_), .A1(new_n3223_), .B0(new_n4691_), .Y(new_n4692_));
  OAI21X1  g02257(.A0(new_n3244_), .A1(pi0161), .B0(new_n4605_), .Y(new_n4693_));
  AOI21X1  g02258(.A0(new_n3240_), .A1(pi0161), .B0(new_n4693_), .Y(new_n4694_));
  AOI21X1  g02259(.A0(new_n3180_), .A1(new_n4611_), .B0(new_n4605_), .Y(new_n4695_));
  OR3X1    g02260(.A(new_n4695_), .B(new_n4694_), .C(pi0228), .Y(new_n4696_));
  AOI21X1  g02261(.A0(new_n4696_), .A1(new_n4609_), .B0(new_n4604_), .Y(new_n4697_));
  OAI21X1  g02262(.A0(new_n4697_), .A1(pi0221), .B0(new_n4603_), .Y(new_n4698_));
  AOI21X1  g02263(.A0(new_n4698_), .A1(new_n2934_), .B0(new_n4620_), .Y(new_n4699_));
  INVX1    g02264(.A(new_n4621_), .Y(new_n4700_));
  AOI21X1  g02265(.A0(new_n4628_), .A1(new_n4473_), .B0(pi0223), .Y(new_n4701_));
  OAI21X1  g02266(.A0(new_n4701_), .A1(new_n4700_), .B0(new_n2939_), .Y(new_n4702_));
  INVX1    g02267(.A(new_n4604_), .Y(new_n4703_));
  AND3X1   g02268(.A(new_n4640_), .B(new_n4638_), .C(new_n3456_), .Y(new_n4704_));
  OAI21X1  g02269(.A0(new_n4704_), .A1(pi0216), .B0(new_n4703_), .Y(new_n4705_));
  AOI21X1  g02270(.A0(new_n4705_), .A1(new_n2437_), .B0(new_n4602_), .Y(new_n4706_));
  MX2X1    g02271(.A(new_n4706_), .B(new_n4622_), .S0(pi0215), .Y(new_n4707_));
  OAI21X1  g02272(.A0(new_n4707_), .A1(new_n2933_), .B0(new_n4634_), .Y(new_n4708_));
  AOI21X1  g02273(.A0(new_n4708_), .A1(pi0039), .B0(pi0038), .Y(new_n4709_));
  OAI21X1  g02274(.A0(new_n4702_), .A1(new_n4699_), .B0(new_n4709_), .Y(new_n4710_));
  AND2X1   g02275(.A(new_n4650_), .B(new_n3257_), .Y(new_n4711_));
  INVX1    g02276(.A(new_n4711_), .Y(new_n4712_));
  AOI21X1  g02277(.A0(new_n4712_), .A1(pi0299), .B0(new_n4635_), .Y(new_n4713_));
  AOI21X1  g02278(.A0(new_n4713_), .A1(pi0038), .B0(pi0100), .Y(new_n4714_));
  INVX1    g02279(.A(new_n4619_), .Y(new_n4715_));
  OR2X1    g02280(.A(new_n4637_), .B(new_n3254_), .Y(new_n4716_));
  OAI21X1  g02281(.A0(new_n4716_), .A1(new_n4659_), .B0(new_n2438_), .Y(new_n4717_));
  AOI21X1  g02282(.A0(new_n4717_), .A1(new_n4703_), .B0(pi0221), .Y(new_n4718_));
  OAI21X1  g02283(.A0(new_n4718_), .A1(new_n4602_), .B0(new_n2934_), .Y(new_n4719_));
  AOI21X1  g02284(.A0(new_n4719_), .A1(new_n4715_), .B0(new_n2933_), .Y(new_n4720_));
  OR3X1    g02285(.A(new_n4720_), .B(new_n4635_), .C(new_n3060_), .Y(new_n4721_));
  AOI21X1  g02286(.A0(new_n4713_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4722_));
  AOI22X1  g02287(.A0(new_n4722_), .A1(new_n4721_), .B0(new_n4714_), .B1(new_n4710_), .Y(new_n4723_));
  INVX1    g02288(.A(new_n4713_), .Y(new_n4724_));
  MX2X1    g02289(.A(new_n4724_), .B(new_n4708_), .S0(new_n3064_), .Y(new_n4725_));
  AOI21X1  g02290(.A0(new_n4725_), .A1(pi0087), .B0(pi0075), .Y(new_n4726_));
  OAI21X1  g02291(.A0(new_n4723_), .A1(pi0087), .B0(new_n4726_), .Y(new_n4727_));
  AOI21X1  g02292(.A0(new_n4713_), .A1(pi0075), .B0(pi0092), .Y(new_n4728_));
  NOR2X1   g02293(.A(new_n4725_), .B(new_n3080_), .Y(new_n4729_));
  OAI21X1  g02294(.A0(new_n4724_), .A1(new_n3077_), .B0(pi0092), .Y(new_n4730_));
  OAI21X1  g02295(.A0(new_n4730_), .A1(new_n4729_), .B0(new_n3102_), .Y(new_n4731_));
  AOI21X1  g02296(.A0(new_n4728_), .A1(new_n4727_), .B0(new_n4731_), .Y(new_n4732_));
  OAI21X1  g02297(.A0(new_n4724_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4733_));
  NAND2X1  g02298(.A(new_n4707_), .B(new_n3104_), .Y(new_n4734_));
  AOI21X1  g02299(.A0(new_n4711_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n4735_));
  AOI21X1  g02300(.A0(new_n4735_), .A1(new_n4734_), .B0(pi0056), .Y(new_n4736_));
  OAI21X1  g02301(.A0(new_n4733_), .A1(new_n4732_), .B0(new_n4736_), .Y(new_n4737_));
  AOI21X1  g02302(.A0(new_n4712_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4738_));
  OAI21X1  g02303(.A0(new_n4707_), .A1(new_n3115_), .B0(new_n4738_), .Y(new_n4739_));
  AND3X1   g02304(.A(new_n4739_), .B(new_n4737_), .C(new_n3222_), .Y(new_n4740_));
  OAI21X1  g02305(.A0(new_n4712_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4741_));
  AOI21X1  g02306(.A0(new_n4707_), .A1(new_n3224_), .B0(new_n4741_), .Y(new_n4742_));
  OR2X1    g02307(.A(new_n4742_), .B(new_n3374_), .Y(new_n4743_));
  AOI21X1  g02308(.A0(new_n4711_), .A1(new_n3374_), .B0(new_n4691_), .Y(new_n4744_));
  OAI21X1  g02309(.A0(new_n4743_), .A1(new_n4740_), .B0(new_n4744_), .Y(new_n4745_));
  OAI21X1  g02310(.A0(new_n4692_), .A1(new_n4690_), .B0(new_n4745_), .Y(po0164));
  INVX1    g02311(.A(pi1134), .Y(new_n4747_));
  NOR4X1   g02312(.A(pi0930), .B(new_n2701_), .C(new_n2437_), .D(pi0216), .Y(new_n4748_));
  INVX1    g02313(.A(new_n4748_), .Y(new_n4749_));
  AOI21X1  g02314(.A0(pi0278), .A1(pi0216), .B0(pi0221), .Y(new_n4750_));
  AOI21X1  g02315(.A0(pi0152), .A1(new_n2447_), .B0(new_n2793_), .Y(new_n4751_));
  INVX1    g02316(.A(new_n4751_), .Y(new_n4752_));
  INVX1    g02317(.A(pi0846), .Y(new_n4753_));
  AOI21X1  g02318(.A0(new_n3232_), .A1(new_n4753_), .B0(new_n2447_), .Y(new_n4754_));
  OAI21X1  g02319(.A0(new_n4754_), .A1(new_n4752_), .B0(new_n2438_), .Y(new_n4755_));
  AOI21X1  g02320(.A0(new_n3244_), .A1(new_n3193_), .B0(pi0846), .Y(new_n4756_));
  OAI21X1  g02321(.A0(new_n3240_), .A1(new_n3193_), .B0(new_n4756_), .Y(new_n4757_));
  NAND3X1  g02322(.A(new_n3180_), .B(pi0846), .C(new_n3193_), .Y(new_n4758_));
  AOI21X1  g02323(.A0(new_n4758_), .A1(new_n4757_), .B0(pi0228), .Y(new_n4759_));
  OAI21X1  g02324(.A0(new_n4759_), .A1(new_n4755_), .B0(new_n4750_), .Y(new_n4760_));
  AOI21X1  g02325(.A0(pi0833), .A1(new_n2438_), .B0(new_n2437_), .Y(new_n4761_));
  NOR3X1   g02326(.A(new_n4761_), .B(new_n2933_), .C(pi0215), .Y(new_n4762_));
  AND3X1   g02327(.A(new_n4762_), .B(new_n4760_), .C(new_n4749_), .Y(new_n4763_));
  NOR4X1   g02328(.A(pi0930), .B(new_n2701_), .C(pi0224), .D(new_n2941_), .Y(new_n4764_));
  INVX1    g02329(.A(new_n4764_), .Y(new_n4765_));
  NOR3X1   g02330(.A(new_n3231_), .B(new_n2454_), .C(pi0846), .Y(new_n4766_));
  AOI21X1  g02331(.A0(pi0278), .A1(pi0224), .B0(pi0222), .Y(new_n4767_));
  OAI21X1  g02332(.A0(new_n4766_), .A1(pi0224), .B0(new_n4767_), .Y(new_n4768_));
  NOR2X1   g02333(.A(pi0299), .B(pi0223), .Y(new_n4769_));
  INVX1    g02334(.A(new_n4769_), .Y(new_n4770_));
  NOR2X1   g02335(.A(new_n4770_), .B(new_n2943_), .Y(new_n4771_));
  AND3X1   g02336(.A(new_n4771_), .B(new_n4768_), .C(new_n4765_), .Y(new_n4772_));
  OR2X1    g02337(.A(new_n4772_), .B(pi0039), .Y(new_n4773_));
  INVX1    g02338(.A(new_n4767_), .Y(new_n4774_));
  AOI21X1  g02339(.A0(new_n2453_), .A1(pi0095), .B0(new_n4753_), .Y(new_n4775_));
  AOI21X1  g02340(.A0(new_n4775_), .A1(new_n2942_), .B0(new_n4774_), .Y(new_n4776_));
  NOR4X1   g02341(.A(new_n4776_), .B(new_n4764_), .C(new_n2943_), .D(pi0223), .Y(new_n4777_));
  NOR2X1   g02342(.A(new_n4777_), .B(pi0299), .Y(new_n4778_));
  AND2X1   g02343(.A(new_n4778_), .B(new_n3594_), .Y(new_n4779_));
  NOR3X1   g02344(.A(new_n4761_), .B(new_n4748_), .C(pi0215), .Y(new_n4780_));
  MX2X1    g02345(.A(new_n4775_), .B(pi0152), .S0(new_n2447_), .Y(new_n4781_));
  AND2X1   g02346(.A(new_n4781_), .B(pi0228), .Y(new_n4782_));
  INVX1    g02347(.A(new_n4782_), .Y(new_n4783_));
  AOI21X1  g02348(.A0(new_n2987_), .A1(new_n4753_), .B0(pi0228), .Y(new_n4784_));
  OAI21X1  g02349(.A0(new_n2987_), .A1(pi0152), .B0(new_n4784_), .Y(new_n4785_));
  AND3X1   g02350(.A(new_n4785_), .B(new_n4783_), .C(new_n3456_), .Y(new_n4786_));
  OAI21X1  g02351(.A0(new_n4786_), .A1(pi0216), .B0(new_n4750_), .Y(new_n4787_));
  AOI21X1  g02352(.A0(new_n4787_), .A1(new_n4780_), .B0(new_n2933_), .Y(new_n4788_));
  OR2X1    g02353(.A(new_n4788_), .B(new_n4779_), .Y(new_n4789_));
  AOI21X1  g02354(.A0(new_n4789_), .A1(pi0039), .B0(pi0038), .Y(new_n4790_));
  OAI21X1  g02355(.A0(new_n4773_), .A1(new_n4763_), .B0(new_n4790_), .Y(new_n4791_));
  AOI21X1  g02356(.A0(new_n2793_), .A1(pi0152), .B0(new_n4782_), .Y(new_n4792_));
  OAI21X1  g02357(.A0(new_n4792_), .A1(pi0216), .B0(new_n4750_), .Y(new_n4793_));
  AOI21X1  g02358(.A0(new_n4793_), .A1(new_n4780_), .B0(new_n3255_), .Y(new_n4794_));
  AOI21X1  g02359(.A0(new_n4794_), .A1(pi0299), .B0(new_n4779_), .Y(new_n4795_));
  AOI21X1  g02360(.A0(new_n4795_), .A1(pi0038), .B0(pi0100), .Y(new_n4796_));
  OR2X1    g02361(.A(new_n4782_), .B(new_n3254_), .Y(new_n4797_));
  OAI22X1  g02362(.A0(new_n3197_), .A1(new_n4753_), .B0(new_n3190_), .B1(new_n3193_), .Y(new_n4798_));
  AOI21X1  g02363(.A0(new_n4798_), .A1(new_n2793_), .B0(new_n4797_), .Y(new_n4799_));
  OAI21X1  g02364(.A0(new_n4799_), .A1(pi0216), .B0(new_n4750_), .Y(new_n4800_));
  AOI21X1  g02365(.A0(new_n4800_), .A1(new_n4780_), .B0(new_n2933_), .Y(new_n4801_));
  OR3X1    g02366(.A(new_n4801_), .B(new_n4779_), .C(new_n3060_), .Y(new_n4802_));
  AOI21X1  g02367(.A0(new_n4795_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4803_));
  AOI22X1  g02368(.A0(new_n4803_), .A1(new_n4802_), .B0(new_n4796_), .B1(new_n4791_), .Y(new_n4804_));
  INVX1    g02369(.A(new_n4795_), .Y(new_n4805_));
  MX2X1    g02370(.A(new_n4805_), .B(new_n4789_), .S0(new_n3064_), .Y(new_n4806_));
  AOI21X1  g02371(.A0(new_n4806_), .A1(pi0087), .B0(pi0075), .Y(new_n4807_));
  OAI21X1  g02372(.A0(new_n4804_), .A1(pi0087), .B0(new_n4807_), .Y(new_n4808_));
  AOI21X1  g02373(.A0(new_n4795_), .A1(pi0075), .B0(pi0092), .Y(new_n4809_));
  NOR2X1   g02374(.A(new_n4806_), .B(new_n3080_), .Y(new_n4810_));
  OAI21X1  g02375(.A0(new_n4805_), .A1(new_n3077_), .B0(pi0092), .Y(new_n4811_));
  OAI21X1  g02376(.A0(new_n4811_), .A1(new_n4810_), .B0(new_n3102_), .Y(new_n4812_));
  AOI21X1  g02377(.A0(new_n4809_), .A1(new_n4808_), .B0(new_n4812_), .Y(new_n4813_));
  OAI21X1  g02378(.A0(new_n4805_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4814_));
  NAND3X1  g02379(.A(new_n4787_), .B(new_n4780_), .C(new_n3104_), .Y(new_n4815_));
  OR2X1    g02380(.A(new_n4794_), .B(new_n3104_), .Y(new_n4816_));
  AND2X1   g02381(.A(new_n4816_), .B(pi0055), .Y(new_n4817_));
  AOI21X1  g02382(.A0(new_n4817_), .A1(new_n4815_), .B0(pi0056), .Y(new_n4818_));
  OAI21X1  g02383(.A0(new_n4814_), .A1(new_n4813_), .B0(new_n4818_), .Y(new_n4819_));
  AND2X1   g02384(.A(new_n4787_), .B(new_n4780_), .Y(new_n4820_));
  AOI21X1  g02385(.A0(new_n4794_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4821_));
  OAI21X1  g02386(.A0(new_n4820_), .A1(new_n3115_), .B0(new_n4821_), .Y(new_n4822_));
  AND2X1   g02387(.A(new_n4822_), .B(new_n3222_), .Y(new_n4823_));
  AND3X1   g02388(.A(new_n4787_), .B(new_n4780_), .C(new_n3224_), .Y(new_n4824_));
  OAI21X1  g02389(.A0(new_n4794_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4825_));
  OAI21X1  g02390(.A0(new_n4825_), .A1(new_n4824_), .B0(new_n3223_), .Y(new_n4826_));
  AOI21X1  g02391(.A0(new_n4823_), .A1(new_n4819_), .B0(new_n4826_), .Y(new_n4827_));
  OAI21X1  g02392(.A0(new_n4794_), .A1(new_n3223_), .B0(pi0242), .Y(new_n4828_));
  INVX1    g02393(.A(new_n4762_), .Y(new_n4829_));
  INVX1    g02394(.A(new_n4750_), .Y(new_n4830_));
  AOI21X1  g02395(.A0(new_n3244_), .A1(pi0152), .B0(new_n4753_), .Y(new_n4831_));
  OAI21X1  g02396(.A0(new_n3240_), .A1(pi0152), .B0(new_n4831_), .Y(new_n4832_));
  AND2X1   g02397(.A(new_n4753_), .B(pi0152), .Y(new_n4833_));
  AOI21X1  g02398(.A0(new_n4833_), .A1(new_n3180_), .B0(pi0228), .Y(new_n4834_));
  AND2X1   g02399(.A(new_n4834_), .B(new_n4832_), .Y(new_n4835_));
  NOR2X1   g02400(.A(new_n4752_), .B(new_n3232_), .Y(new_n4836_));
  NOR3X1   g02401(.A(new_n4836_), .B(new_n4835_), .C(new_n4755_), .Y(new_n4837_));
  OAI21X1  g02402(.A0(new_n4837_), .A1(new_n4830_), .B0(new_n4749_), .Y(new_n4838_));
  OR4X1    g02403(.A(new_n3231_), .B(new_n2454_), .C(new_n4753_), .D(pi0224), .Y(new_n4839_));
  AND2X1   g02404(.A(new_n4839_), .B(new_n4767_), .Y(new_n4840_));
  OR4X1    g02405(.A(new_n4840_), .B(new_n4764_), .C(new_n4770_), .D(new_n2943_), .Y(new_n4841_));
  AND2X1   g02406(.A(new_n4841_), .B(new_n2939_), .Y(new_n4842_));
  OAI21X1  g02407(.A0(new_n4838_), .A1(new_n4829_), .B0(new_n4842_), .Y(new_n4843_));
  NOR2X1   g02408(.A(new_n4761_), .B(pi0215), .Y(new_n4844_));
  INVX1    g02409(.A(new_n4844_), .Y(new_n4845_));
  AOI21X1  g02410(.A0(new_n4785_), .A1(new_n4783_), .B0(pi0216), .Y(new_n4846_));
  NOR2X1   g02411(.A(new_n4846_), .B(new_n4830_), .Y(new_n4847_));
  NOR3X1   g02412(.A(new_n4847_), .B(new_n4845_), .C(new_n4748_), .Y(new_n4848_));
  MX2X1    g02413(.A(new_n4848_), .B(new_n4777_), .S0(new_n2933_), .Y(new_n4849_));
  INVX1    g02414(.A(new_n4849_), .Y(new_n4850_));
  AOI21X1  g02415(.A0(new_n4850_), .A1(pi0039), .B0(pi0038), .Y(new_n4851_));
  AND2X1   g02416(.A(new_n4793_), .B(new_n4780_), .Y(new_n4852_));
  MX2X1    g02417(.A(new_n4852_), .B(new_n4777_), .S0(new_n2933_), .Y(new_n4853_));
  INVX1    g02418(.A(new_n4853_), .Y(new_n4854_));
  OAI21X1  g02419(.A0(new_n4854_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4855_));
  AOI21X1  g02420(.A0(new_n4851_), .A1(new_n4843_), .B0(new_n4855_), .Y(new_n4856_));
  AOI21X1  g02421(.A0(new_n4798_), .A1(new_n2793_), .B0(new_n4782_), .Y(new_n4857_));
  OAI21X1  g02422(.A0(new_n4857_), .A1(pi0216), .B0(new_n4750_), .Y(new_n4858_));
  AOI21X1  g02423(.A0(new_n4858_), .A1(new_n4780_), .B0(new_n2933_), .Y(new_n4859_));
  OR3X1    g02424(.A(new_n4859_), .B(new_n4778_), .C(new_n3060_), .Y(new_n4860_));
  AOI21X1  g02425(.A0(new_n4853_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4861_));
  AOI21X1  g02426(.A0(new_n4861_), .A1(new_n4860_), .B0(new_n4856_), .Y(new_n4862_));
  MX2X1    g02427(.A(new_n4854_), .B(new_n4850_), .S0(new_n3064_), .Y(new_n4863_));
  AOI21X1  g02428(.A0(new_n4863_), .A1(pi0087), .B0(pi0075), .Y(new_n4864_));
  OAI21X1  g02429(.A0(new_n4862_), .A1(pi0087), .B0(new_n4864_), .Y(new_n4865_));
  AOI21X1  g02430(.A0(new_n4853_), .A1(pi0075), .B0(pi0092), .Y(new_n4866_));
  NOR2X1   g02431(.A(new_n4863_), .B(new_n3080_), .Y(new_n4867_));
  OAI21X1  g02432(.A0(new_n4854_), .A1(new_n3077_), .B0(pi0092), .Y(new_n4868_));
  OAI21X1  g02433(.A0(new_n4868_), .A1(new_n4867_), .B0(new_n3102_), .Y(new_n4869_));
  AOI21X1  g02434(.A0(new_n4866_), .A1(new_n4865_), .B0(new_n4869_), .Y(new_n4870_));
  OAI21X1  g02435(.A0(new_n4854_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4871_));
  OR4X1    g02436(.A(new_n4847_), .B(new_n4845_), .C(new_n4748_), .D(new_n3105_), .Y(new_n4872_));
  AOI21X1  g02437(.A0(new_n4852_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n4873_));
  AOI21X1  g02438(.A0(new_n4873_), .A1(new_n4872_), .B0(pi0056), .Y(new_n4874_));
  OAI21X1  g02439(.A0(new_n4871_), .A1(new_n4870_), .B0(new_n4874_), .Y(new_n4875_));
  INVX1    g02440(.A(new_n4852_), .Y(new_n4876_));
  AOI21X1  g02441(.A0(new_n4876_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4877_));
  OAI21X1  g02442(.A0(new_n4848_), .A1(new_n3115_), .B0(new_n4877_), .Y(new_n4878_));
  AND2X1   g02443(.A(new_n4878_), .B(new_n3222_), .Y(new_n4879_));
  NOR4X1   g02444(.A(new_n4847_), .B(new_n4845_), .C(new_n4748_), .D(new_n3225_), .Y(new_n4880_));
  OAI21X1  g02445(.A0(new_n4876_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4881_));
  OAI21X1  g02446(.A0(new_n4881_), .A1(new_n4880_), .B0(new_n3223_), .Y(new_n4882_));
  AOI21X1  g02447(.A0(new_n4879_), .A1(new_n4875_), .B0(new_n4882_), .Y(new_n4883_));
  INVX1    g02448(.A(pi0242), .Y(new_n4884_));
  OAI21X1  g02449(.A0(new_n4876_), .A1(new_n3223_), .B0(new_n4884_), .Y(new_n4885_));
  OAI22X1  g02450(.A0(new_n4885_), .A1(new_n4883_), .B0(new_n4828_), .B1(new_n4827_), .Y(new_n4886_));
  AOI21X1  g02451(.A0(new_n4768_), .A1(new_n4765_), .B0(new_n4770_), .Y(new_n4887_));
  OR2X1    g02452(.A(new_n4887_), .B(pi0039), .Y(new_n4888_));
  AND2X1   g02453(.A(pi0299), .B(new_n2934_), .Y(new_n4889_));
  INVX1    g02454(.A(new_n4889_), .Y(new_n4890_));
  AOI21X1  g02455(.A0(new_n4760_), .A1(new_n4749_), .B0(new_n4890_), .Y(new_n4891_));
  AOI21X1  g02456(.A0(new_n4779_), .A1(new_n2944_), .B0(pi0299), .Y(new_n4892_));
  INVX1    g02457(.A(new_n4892_), .Y(new_n4893_));
  AOI21X1  g02458(.A0(new_n4787_), .A1(new_n4749_), .B0(pi0215), .Y(new_n4894_));
  OAI21X1  g02459(.A0(new_n4894_), .A1(new_n2933_), .B0(new_n4893_), .Y(new_n4895_));
  AOI21X1  g02460(.A0(new_n4895_), .A1(pi0039), .B0(pi0038), .Y(new_n4896_));
  OAI21X1  g02461(.A0(new_n4891_), .A1(new_n4888_), .B0(new_n4896_), .Y(new_n4897_));
  AOI21X1  g02462(.A0(new_n4793_), .A1(new_n4749_), .B0(pi0215), .Y(new_n4898_));
  AND2X1   g02463(.A(new_n4898_), .B(new_n3257_), .Y(new_n4899_));
  INVX1    g02464(.A(new_n4899_), .Y(new_n4900_));
  AOI21X1  g02465(.A0(new_n4900_), .A1(pi0299), .B0(new_n4892_), .Y(new_n4901_));
  AOI21X1  g02466(.A0(new_n4901_), .A1(pi0038), .B0(pi0100), .Y(new_n4902_));
  AOI21X1  g02467(.A0(new_n4800_), .A1(new_n4749_), .B0(pi0215), .Y(new_n4903_));
  NOR2X1   g02468(.A(new_n4892_), .B(new_n3060_), .Y(new_n4904_));
  OAI21X1  g02469(.A0(new_n4903_), .A1(new_n2933_), .B0(new_n4904_), .Y(new_n4905_));
  AOI21X1  g02470(.A0(new_n4901_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4906_));
  AOI22X1  g02471(.A0(new_n4906_), .A1(new_n4905_), .B0(new_n4902_), .B1(new_n4897_), .Y(new_n4907_));
  INVX1    g02472(.A(new_n4901_), .Y(new_n4908_));
  MX2X1    g02473(.A(new_n4908_), .B(new_n4895_), .S0(new_n3064_), .Y(new_n4909_));
  AOI21X1  g02474(.A0(new_n4909_), .A1(pi0087), .B0(pi0075), .Y(new_n4910_));
  OAI21X1  g02475(.A0(new_n4907_), .A1(pi0087), .B0(new_n4910_), .Y(new_n4911_));
  AOI21X1  g02476(.A0(new_n4901_), .A1(pi0075), .B0(pi0092), .Y(new_n4912_));
  NOR2X1   g02477(.A(new_n4909_), .B(new_n3080_), .Y(new_n4913_));
  OAI21X1  g02478(.A0(new_n4908_), .A1(new_n3077_), .B0(pi0092), .Y(new_n4914_));
  OAI21X1  g02479(.A0(new_n4914_), .A1(new_n4913_), .B0(new_n3102_), .Y(new_n4915_));
  AOI21X1  g02480(.A0(new_n4912_), .A1(new_n4911_), .B0(new_n4915_), .Y(new_n4916_));
  OAI21X1  g02481(.A0(new_n4908_), .A1(new_n3102_), .B0(new_n3107_), .Y(new_n4917_));
  NAND2X1  g02482(.A(new_n4894_), .B(new_n3104_), .Y(new_n4918_));
  AOI21X1  g02483(.A0(new_n4899_), .A1(new_n3105_), .B0(new_n3107_), .Y(new_n4919_));
  AOI21X1  g02484(.A0(new_n4919_), .A1(new_n4918_), .B0(pi0056), .Y(new_n4920_));
  OAI21X1  g02485(.A0(new_n4917_), .A1(new_n4916_), .B0(new_n4920_), .Y(new_n4921_));
  AOI21X1  g02486(.A0(new_n4900_), .A1(new_n3115_), .B0(new_n3118_), .Y(new_n4922_));
  OAI21X1  g02487(.A0(new_n4894_), .A1(new_n3115_), .B0(new_n4922_), .Y(new_n4923_));
  AND3X1   g02488(.A(new_n4923_), .B(new_n4921_), .C(new_n3222_), .Y(new_n4924_));
  OAI21X1  g02489(.A0(new_n4900_), .A1(new_n3224_), .B0(pi0062), .Y(new_n4925_));
  AOI21X1  g02490(.A0(new_n4894_), .A1(new_n3224_), .B0(new_n4925_), .Y(new_n4926_));
  OR2X1    g02491(.A(new_n4926_), .B(new_n3374_), .Y(new_n4927_));
  AOI21X1  g02492(.A0(new_n4899_), .A1(new_n3374_), .B0(new_n4884_), .Y(new_n4928_));
  OAI21X1  g02493(.A0(new_n4927_), .A1(new_n4924_), .B0(new_n4928_), .Y(new_n4929_));
  NAND2X1  g02494(.A(new_n4838_), .B(new_n4889_), .Y(new_n4930_));
  AOI21X1  g02495(.A0(new_n4840_), .A1(new_n4769_), .B0(new_n4888_), .Y(new_n4931_));
  NAND2X1  g02496(.A(new_n4931_), .B(new_n4930_), .Y(new_n4932_));
  NAND2X1  g02497(.A(new_n4776_), .B(new_n2940_), .Y(new_n4933_));
  OAI21X1  g02498(.A0(new_n4847_), .A1(new_n4748_), .B0(new_n2934_), .Y(new_n4934_));
  AOI22X1  g02499(.A0(new_n4934_), .A1(pi0299), .B0(new_n4933_), .B1(new_n4892_), .Y(new_n4935_));
  INVX1    g02500(.A(new_n4935_), .Y(new_n4936_));
  AOI21X1  g02501(.A0(new_n4936_), .A1(pi0039), .B0(pi0038), .Y(new_n4937_));
  INVX1    g02502(.A(new_n4898_), .Y(new_n4938_));
  AOI22X1  g02503(.A0(new_n4933_), .A1(new_n4892_), .B0(new_n4938_), .B1(pi0299), .Y(new_n4939_));
  INVX1    g02504(.A(new_n4939_), .Y(new_n4940_));
  OAI21X1  g02505(.A0(new_n4940_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n4941_));
  AOI21X1  g02506(.A0(new_n4937_), .A1(new_n4932_), .B0(new_n4941_), .Y(new_n4942_));
  AOI21X1  g02507(.A0(new_n4858_), .A1(new_n4749_), .B0(pi0215), .Y(new_n4943_));
  AOI21X1  g02508(.A0(new_n4933_), .A1(new_n4892_), .B0(new_n3060_), .Y(new_n4944_));
  OAI21X1  g02509(.A0(new_n4943_), .A1(new_n2933_), .B0(new_n4944_), .Y(new_n4945_));
  AOI21X1  g02510(.A0(new_n4939_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n4946_));
  AND2X1   g02511(.A(new_n4946_), .B(new_n4945_), .Y(new_n4947_));
  OAI21X1  g02512(.A0(new_n4947_), .A1(new_n4942_), .B0(new_n3131_), .Y(new_n4948_));
  MX2X1    g02513(.A(new_n4940_), .B(new_n4936_), .S0(new_n3064_), .Y(new_n4949_));
  AOI21X1  g02514(.A0(new_n4949_), .A1(pi0087), .B0(pi0075), .Y(new_n4950_));
  OAI21X1  g02515(.A0(new_n4940_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n4951_));
  AOI21X1  g02516(.A0(new_n4950_), .A1(new_n4948_), .B0(new_n4951_), .Y(new_n4952_));
  AOI21X1  g02517(.A0(new_n4939_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n4953_));
  OAI21X1  g02518(.A0(new_n4949_), .A1(new_n3080_), .B0(new_n4953_), .Y(new_n4954_));
  NAND2X1  g02519(.A(new_n4954_), .B(new_n3102_), .Y(new_n4955_));
  OR2X1    g02520(.A(new_n4955_), .B(new_n4952_), .Y(new_n4956_));
  AOI21X1  g02521(.A0(new_n4939_), .A1(new_n3130_), .B0(pi0055), .Y(new_n4957_));
  NOR2X1   g02522(.A(new_n4934_), .B(new_n3105_), .Y(new_n4958_));
  OAI21X1  g02523(.A0(new_n4938_), .A1(new_n3104_), .B0(pi0055), .Y(new_n4959_));
  OAI21X1  g02524(.A0(new_n4959_), .A1(new_n4958_), .B0(new_n3118_), .Y(new_n4960_));
  AOI21X1  g02525(.A0(new_n4957_), .A1(new_n4956_), .B0(new_n4960_), .Y(new_n4961_));
  OAI21X1  g02526(.A0(new_n4898_), .A1(new_n3114_), .B0(pi0056), .Y(new_n4962_));
  AOI21X1  g02527(.A0(new_n4934_), .A1(new_n3114_), .B0(new_n4962_), .Y(new_n4963_));
  OR2X1    g02528(.A(new_n4963_), .B(pi0062), .Y(new_n4964_));
  AOI21X1  g02529(.A0(new_n4898_), .A1(new_n3225_), .B0(new_n3222_), .Y(new_n4965_));
  OAI21X1  g02530(.A0(new_n4934_), .A1(new_n3225_), .B0(new_n4965_), .Y(new_n4966_));
  AND2X1   g02531(.A(new_n4966_), .B(new_n3223_), .Y(new_n4967_));
  OAI21X1  g02532(.A0(new_n4964_), .A1(new_n4961_), .B0(new_n4967_), .Y(new_n4968_));
  AOI21X1  g02533(.A0(new_n4898_), .A1(new_n3374_), .B0(pi0242), .Y(new_n4969_));
  AOI21X1  g02534(.A0(new_n4969_), .A1(new_n4968_), .B0(new_n4747_), .Y(new_n4970_));
  AOI22X1  g02535(.A0(new_n4970_), .A1(new_n4929_), .B0(new_n4886_), .B1(new_n4747_), .Y(po0165));
  AND2X1   g02536(.A(pi0059), .B(pi0057), .Y(new_n4973_));
  INVX1    g02537(.A(new_n4973_), .Y(new_n4974_));
  INVX1    g02538(.A(new_n3123_), .Y(new_n4975_));
  NOR4X1   g02539(.A(new_n4975_), .B(new_n3115_), .C(new_n2985_), .D(new_n2536_), .Y(new_n4976_));
  OAI21X1  g02540(.A0(new_n4976_), .A1(new_n3223_), .B0(new_n4974_), .Y(new_n4977_));
  INVX1    g02541(.A(new_n4977_), .Y(new_n4978_));
  AND2X1   g02542(.A(new_n3064_), .B(new_n2982_), .Y(new_n4979_));
  AOI21X1  g02543(.A0(new_n4979_), .A1(new_n3113_), .B0(new_n3118_), .Y(new_n4980_));
  INVX1    g02544(.A(new_n4980_), .Y(new_n4981_));
  INVX1    g02545(.A(pi0074), .Y(new_n4982_));
  NOR4X1   g02546(.A(pi0092), .B(pi0087), .C(pi0075), .D(pi0054), .Y(new_n4983_));
  AOI21X1  g02547(.A0(new_n4983_), .A1(new_n4979_), .B0(new_n4982_), .Y(new_n4984_));
  OR2X1    g02548(.A(new_n4984_), .B(pi0055), .Y(new_n4985_));
  AND2X1   g02549(.A(new_n2982_), .B(new_n2939_), .Y(new_n4986_));
  INVX1    g02550(.A(new_n4986_), .Y(new_n4987_));
  AOI21X1  g02551(.A0(new_n4987_), .A1(pi0038), .B0(pi0100), .Y(new_n4988_));
  INVX1    g02552(.A(new_n4988_), .Y(new_n4989_));
  INVX1    g02553(.A(new_n2533_), .Y(new_n4990_));
  OR2X1    g02554(.A(new_n2505_), .B(new_n2494_), .Y(new_n4991_));
  AND2X1   g02555(.A(new_n4991_), .B(new_n2682_), .Y(new_n4992_));
  OR4X1    g02556(.A(new_n2666_), .B(new_n2662_), .C(new_n2568_), .D(new_n2490_), .Y(new_n4993_));
  AOI21X1  g02557(.A0(new_n4993_), .A1(new_n2571_), .B0(new_n2565_), .Y(new_n4994_));
  OAI21X1  g02558(.A0(new_n4994_), .A1(pi0108), .B0(new_n2563_), .Y(new_n4995_));
  NOR3X1   g02559(.A(new_n2677_), .B(pi0110), .C(pi0109), .Y(new_n4996_));
  OR2X1    g02560(.A(new_n2557_), .B(new_n2549_), .Y(new_n4997_));
  AOI21X1  g02561(.A0(new_n4996_), .A1(new_n4995_), .B0(new_n4997_), .Y(new_n4998_));
  OR2X1    g02562(.A(pi0091), .B(pi0058), .Y(new_n4999_));
  NOR2X1   g02563(.A(new_n2553_), .B(new_n4999_), .Y(new_n5000_));
  OAI21X1  g02564(.A0(new_n4998_), .A1(pi0047), .B0(new_n5000_), .Y(new_n5001_));
  AOI21X1  g02565(.A0(new_n5001_), .A1(new_n4992_), .B0(new_n2683_), .Y(new_n5002_));
  OAI21X1  g02566(.A0(new_n2833_), .A1(pi0841), .B0(pi0093), .Y(new_n5003_));
  OAI21X1  g02567(.A0(new_n5002_), .A1(pi0093), .B0(new_n5003_), .Y(new_n5004_));
  OR2X1    g02568(.A(new_n2507_), .B(pi0070), .Y(new_n5005_));
  AOI21X1  g02569(.A0(new_n5004_), .A1(new_n2508_), .B0(new_n5005_), .Y(new_n5006_));
  OAI21X1  g02570(.A0(new_n5006_), .A1(pi0051), .B0(new_n2537_), .Y(new_n5007_));
  AOI21X1  g02571(.A0(new_n5007_), .A1(new_n2852_), .B0(new_n4990_), .Y(new_n5008_));
  MX2X1    g02572(.A(pi0198), .B(pi0210), .S0(pi0299), .Y(new_n5009_));
  NOR2X1   g02573(.A(new_n2526_), .B(pi0035), .Y(new_n5010_));
  AND3X1   g02574(.A(new_n5010_), .B(new_n2706_), .C(new_n2529_), .Y(new_n5011_));
  OR2X1    g02575(.A(new_n5011_), .B(new_n2455_), .Y(new_n5012_));
  MX2X1    g02576(.A(new_n5012_), .B(new_n3176_), .S0(new_n5009_), .Y(new_n5013_));
  OAI21X1  g02577(.A0(new_n5008_), .A1(new_n2795_), .B0(new_n5013_), .Y(new_n5014_));
  AOI21X1  g02578(.A0(new_n5014_), .A1(new_n2523_), .B0(new_n2696_), .Y(new_n5015_));
  INVX1    g02579(.A(pi0642), .Y(new_n5016_));
  NOR2X1   g02580(.A(pi0616), .B(pi0614), .Y(new_n5017_));
  AND3X1   g02581(.A(new_n5017_), .B(new_n5016_), .C(pi0603), .Y(new_n5018_));
  INVX1    g02582(.A(pi0680), .Y(new_n5019_));
  NOR4X1   g02583(.A(pi0681), .B(new_n5019_), .C(pi0662), .D(pi0661), .Y(new_n5020_));
  NOR2X1   g02584(.A(new_n5020_), .B(new_n5018_), .Y(new_n5021_));
  INVX1    g02585(.A(new_n5021_), .Y(po1101));
  NOR2X1   g02586(.A(pi0468), .B(pi0332), .Y(new_n5023_));
  INVX1    g02587(.A(pi1092), .Y(new_n5024_));
  AND2X1   g02588(.A(pi0984), .B(pi0835), .Y(new_n5025_));
  INVX1    g02589(.A(pi0979), .Y(new_n5026_));
  OR2X1    g02590(.A(pi1001), .B(pi0252), .Y(new_n5027_));
  NAND2X1  g02591(.A(new_n5027_), .B(new_n5026_), .Y(new_n5028_));
  NAND2X1  g02592(.A(pi0950), .B(pi0835), .Y(new_n5029_));
  OR4X1    g02593(.A(new_n5029_), .B(new_n5028_), .C(new_n5025_), .D(pi0287), .Y(new_n5030_));
  NOR2X1   g02594(.A(pi0829), .B(pi0824), .Y(new_n5031_));
  INVX1    g02595(.A(pi1093), .Y(new_n5032_));
  AND2X1   g02596(.A(new_n2702_), .B(pi0824), .Y(new_n5033_));
  NOR3X1   g02597(.A(new_n5033_), .B(new_n2703_), .C(new_n5032_), .Y(new_n5034_));
  NOR4X1   g02598(.A(new_n5034_), .B(new_n5031_), .C(new_n5030_), .D(new_n5024_), .Y(new_n5035_));
  OAI21X1  g02599(.A0(new_n5035_), .A1(new_n5023_), .B0(po1101), .Y(new_n5036_));
  AND2X1   g02600(.A(new_n5023_), .B(new_n2982_), .Y(new_n5037_));
  AOI22X1  g02601(.A0(new_n5037_), .A1(po1101), .B0(new_n5036_), .B1(new_n2987_), .Y(new_n5038_));
  NOR4X1   g02602(.A(pi0977), .B(pi0974), .C(pi0971), .D(pi0969), .Y(new_n5039_));
  NOR4X1   g02603(.A(pi0967), .B(pi0961), .C(pi0602), .D(pi0587), .Y(new_n5040_));
  AND2X1   g02604(.A(new_n5040_), .B(new_n5039_), .Y(new_n5041_));
  INVX1    g02605(.A(new_n5041_), .Y(new_n5042_));
  NOR3X1   g02606(.A(new_n5023_), .B(new_n5020_), .C(new_n5018_), .Y(new_n5043_));
  INVX1    g02607(.A(new_n5043_), .Y(new_n5044_));
  AOI21X1  g02608(.A0(new_n5044_), .A1(new_n5035_), .B0(new_n2986_), .Y(new_n5045_));
  AOI21X1  g02609(.A0(new_n5045_), .A1(new_n5042_), .B0(new_n2940_), .Y(new_n5046_));
  OAI21X1  g02610(.A0(new_n5042_), .A1(new_n5038_), .B0(new_n5046_), .Y(new_n5047_));
  INVX1    g02611(.A(new_n5023_), .Y(new_n5048_));
  MX2X1    g02612(.A(new_n5041_), .B(new_n5021_), .S0(new_n5048_), .Y(new_n5049_));
  NOR4X1   g02613(.A(new_n5030_), .B(new_n2725_), .C(new_n2724_), .D(new_n2704_), .Y(new_n5050_));
  INVX1    g02614(.A(new_n5050_), .Y(new_n5051_));
  NOR4X1   g02615(.A(new_n5051_), .B(new_n5049_), .C(new_n2942_), .D(new_n2941_), .Y(new_n5052_));
  OAI21X1  g02616(.A0(new_n5052_), .A1(new_n2986_), .B0(new_n2940_), .Y(new_n5053_));
  AND3X1   g02617(.A(new_n5053_), .B(new_n5047_), .C(new_n2933_), .Y(new_n5054_));
  NOR2X1   g02618(.A(pi0947), .B(pi0907), .Y(new_n5055_));
  OR4X1    g02619(.A(pi0978), .B(pi0975), .C(pi0972), .D(pi0970), .Y(new_n5056_));
  NOR3X1   g02620(.A(new_n5056_), .B(pi0963), .C(pi0960), .Y(new_n5057_));
  AND2X1   g02621(.A(new_n5057_), .B(new_n5055_), .Y(new_n5058_));
  INVX1    g02622(.A(new_n5058_), .Y(new_n5059_));
  AOI21X1  g02623(.A0(new_n5059_), .A1(new_n5045_), .B0(new_n2934_), .Y(new_n5060_));
  OAI21X1  g02624(.A0(new_n5059_), .A1(new_n5038_), .B0(new_n5060_), .Y(new_n5061_));
  MX2X1    g02625(.A(new_n5058_), .B(new_n5021_), .S0(new_n5048_), .Y(new_n5062_));
  NOR4X1   g02626(.A(new_n5062_), .B(new_n5051_), .C(new_n2437_), .D(new_n2438_), .Y(new_n5063_));
  OAI21X1  g02627(.A0(new_n5063_), .A1(new_n2986_), .B0(new_n2934_), .Y(new_n5064_));
  AND3X1   g02628(.A(new_n5064_), .B(new_n5061_), .C(pi0299), .Y(new_n5065_));
  OR3X1    g02629(.A(new_n5065_), .B(new_n5054_), .C(new_n2939_), .Y(new_n5066_));
  OAI21X1  g02630(.A0(new_n5015_), .A1(pi0039), .B0(new_n5066_), .Y(new_n5067_));
  AOI21X1  g02631(.A0(new_n5067_), .A1(new_n2979_), .B0(new_n4989_), .Y(new_n5068_));
  NOR2X1   g02632(.A(new_n2961_), .B(pi0142), .Y(new_n5069_));
  INVX1    g02633(.A(new_n5069_), .Y(new_n5070_));
  MX2X1    g02634(.A(new_n5070_), .B(new_n3038_), .S0(pi0299), .Y(new_n5071_));
  INVX1    g02635(.A(new_n5071_), .Y(new_n5072_));
  NOR2X1   g02636(.A(new_n5072_), .B(new_n3194_), .Y(new_n5073_));
  AND2X1   g02637(.A(pi0100), .B(new_n2979_), .Y(new_n5074_));
  INVX1    g02638(.A(new_n5074_), .Y(new_n5075_));
  NOR4X1   g02639(.A(new_n5075_), .B(new_n2985_), .C(new_n2536_), .D(pi0039), .Y(new_n5076_));
  INVX1    g02640(.A(pi0683), .Y(new_n5077_));
  INVX1    g02641(.A(pi0044), .Y(new_n5078_));
  NOR3X1   g02642(.A(pi0101), .B(pi0099), .C(pi0041), .Y(new_n5079_));
  OR4X1    g02643(.A(pi0116), .B(pi0115), .C(pi0114), .D(pi0113), .Y(new_n5080_));
  NOR4X1   g02644(.A(new_n5080_), .B(pi0052), .C(pi0043), .D(pi0042), .Y(new_n5081_));
  AND3X1   g02645(.A(new_n5081_), .B(new_n5079_), .C(new_n5078_), .Y(new_n5082_));
  INVX1    g02646(.A(pi0129), .Y(new_n5083_));
  INVX1    g02647(.A(pi0950), .Y(new_n5084_));
  NOR4X1   g02648(.A(new_n5031_), .B(pi1093), .C(new_n5024_), .D(new_n5084_), .Y(po0740));
  MX2X1    g02649(.A(po0740), .B(new_n5083_), .S0(pi0250), .Y(new_n5086_));
  OR4X1    g02650(.A(new_n5086_), .B(new_n5082_), .C(new_n5071_), .D(new_n5077_), .Y(new_n5087_));
  NAND2X1  g02651(.A(new_n5087_), .B(new_n5076_), .Y(new_n5088_));
  OAI21X1  g02652(.A0(new_n5088_), .A1(new_n5073_), .B0(new_n3131_), .Y(new_n5089_));
  OR2X1    g02653(.A(new_n4979_), .B(new_n3131_), .Y(new_n5090_));
  AND2X1   g02654(.A(new_n5090_), .B(new_n3073_), .Y(new_n5091_));
  AND3X1   g02655(.A(new_n5091_), .B(new_n3079_), .C(new_n3091_), .Y(new_n5092_));
  OAI21X1  g02656(.A0(new_n5089_), .A1(new_n5068_), .B0(new_n5092_), .Y(new_n5093_));
  AOI21X1  g02657(.A0(new_n5093_), .A1(new_n4982_), .B0(new_n4985_), .Y(new_n5094_));
  OAI21X1  g02658(.A0(new_n5094_), .A1(pi0056), .B0(new_n4981_), .Y(new_n5095_));
  AND2X1   g02659(.A(new_n3113_), .B(new_n3118_), .Y(new_n5096_));
  AOI21X1  g02660(.A0(new_n4979_), .A1(new_n5096_), .B0(new_n3222_), .Y(new_n5097_));
  OR2X1    g02661(.A(new_n5097_), .B(pi0059), .Y(new_n5098_));
  AOI21X1  g02662(.A0(new_n5095_), .A1(new_n3222_), .B0(new_n5098_), .Y(new_n5099_));
  MX2X1    g02663(.A(new_n5099_), .B(new_n4978_), .S0(pi0057), .Y(po0167));
  INVX1    g02664(.A(pi1090), .Y(po0170));
  NOR4X1   g02665(.A(pi0062), .B(pi0059), .C(pi0056), .D(pi0055), .Y(new_n5102_));
  INVX1    g02666(.A(new_n5102_), .Y(new_n5103_));
  AOI21X1  g02667(.A0(new_n5103_), .A1(new_n2793_), .B0(new_n2436_), .Y(new_n5104_));
  MX2X1    g02668(.A(pi0907), .B(new_n5020_), .S0(new_n5048_), .Y(new_n5105_));
  AND2X1   g02669(.A(pi0228), .B(pi0030), .Y(new_n5106_));
  NOR2X1   g02670(.A(new_n5106_), .B(new_n3603_), .Y(new_n5107_));
  AOI21X1  g02671(.A0(new_n3105_), .A1(new_n2793_), .B0(new_n5107_), .Y(new_n5108_));
  AND2X1   g02672(.A(new_n5108_), .B(new_n5105_), .Y(new_n5109_));
  AND2X1   g02673(.A(new_n5106_), .B(new_n5105_), .Y(new_n5110_));
  OR2X1    g02674(.A(new_n5110_), .B(new_n2933_), .Y(new_n5111_));
  INVX1    g02675(.A(new_n5105_), .Y(new_n5112_));
  AND2X1   g02676(.A(pi0159), .B(pi0158), .Y(new_n5113_));
  AND3X1   g02677(.A(new_n5113_), .B(pi0197), .C(pi0160), .Y(new_n5114_));
  INVX1    g02678(.A(new_n2880_), .Y(new_n5115_));
  INVX1    g02679(.A(new_n2683_), .Y(new_n5116_));
  INVX1    g02680(.A(pi0314), .Y(new_n5117_));
  INVX1    g02681(.A(new_n2678_), .Y(new_n5118_));
  NOR2X1   g02682(.A(new_n2557_), .B(new_n2556_), .Y(new_n5119_));
  INVX1    g02683(.A(new_n2575_), .Y(new_n5120_));
  INVX1    g02684(.A(new_n2670_), .Y(new_n5121_));
  INVX1    g02685(.A(new_n2642_), .Y(new_n5122_));
  NOR2X1   g02686(.A(pi0084), .B(pi0068), .Y(new_n5123_));
  INVX1    g02687(.A(pi0085), .Y(new_n5124_));
  NOR3X1   g02688(.A(new_n2622_), .B(new_n2606_), .C(new_n5124_), .Y(new_n5125_));
  OAI21X1  g02689(.A0(new_n5125_), .A1(new_n2462_), .B0(new_n2626_), .Y(new_n5126_));
  OR2X1    g02690(.A(new_n2634_), .B(new_n2605_), .Y(new_n5127_));
  AOI21X1  g02691(.A0(new_n5126_), .A1(new_n5123_), .B0(new_n5127_), .Y(new_n5128_));
  AOI21X1  g02692(.A0(new_n5128_), .A1(new_n5122_), .B0(new_n2638_), .Y(new_n5129_));
  OR2X1    g02693(.A(new_n2467_), .B(new_n2462_), .Y(new_n5130_));
  INVX1    g02694(.A(new_n5130_), .Y(new_n5131_));
  AOI21X1  g02695(.A0(new_n5131_), .A1(pi0067), .B0(new_n2600_), .Y(new_n5132_));
  OAI21X1  g02696(.A0(new_n5129_), .A1(new_n2637_), .B0(new_n5132_), .Y(new_n5133_));
  AOI21X1  g02697(.A0(new_n5133_), .A1(new_n2598_), .B0(pi0071), .Y(new_n5134_));
  OR3X1    g02698(.A(pi0107), .B(pi0064), .C(pi0063), .Y(po1049));
  OR3X1    g02699(.A(po1049), .B(new_n2588_), .C(pi0065), .Y(new_n5136_));
  OAI21X1  g02700(.A0(new_n5136_), .A1(new_n5134_), .B0(new_n2579_), .Y(new_n5137_));
  NOR4X1   g02701(.A(po1049), .B(new_n2647_), .C(new_n2588_), .D(pi0065), .Y(new_n5138_));
  INVX1    g02702(.A(new_n2558_), .Y(new_n5139_));
  AOI21X1  g02703(.A0(new_n2470_), .A1(pi0081), .B0(pi0102), .Y(new_n5140_));
  AND3X1   g02704(.A(new_n5140_), .B(new_n5139_), .C(new_n2576_), .Y(new_n5141_));
  OAI21X1  g02705(.A0(new_n5138_), .A1(new_n5137_), .B0(new_n5141_), .Y(new_n5142_));
  AOI21X1  g02706(.A0(new_n5142_), .A1(new_n2578_), .B0(new_n5121_), .Y(new_n5143_));
  OAI21X1  g02707(.A0(new_n5143_), .A1(new_n2729_), .B0(new_n5120_), .Y(new_n5144_));
  OR3X1    g02708(.A(new_n2573_), .B(new_n2473_), .C(pi0046), .Y(new_n5145_));
  AOI21X1  g02709(.A0(new_n5144_), .A1(new_n2566_), .B0(new_n5145_), .Y(new_n5146_));
  OAI21X1  g02710(.A0(new_n5146_), .A1(new_n5118_), .B0(new_n5119_), .Y(new_n5147_));
  AND3X1   g02711(.A(new_n5147_), .B(new_n5117_), .C(new_n2515_), .Y(new_n5148_));
  INVX1    g02712(.A(new_n2544_), .Y(new_n5149_));
  AOI21X1  g02713(.A0(new_n5149_), .A1(pi0091), .B0(pi0058), .Y(new_n5150_));
  AND2X1   g02714(.A(pi0314), .B(new_n2515_), .Y(new_n5151_));
  INVX1    g02715(.A(new_n5151_), .Y(new_n5152_));
  INVX1    g02716(.A(new_n5119_), .Y(new_n5153_));
  INVX1    g02717(.A(new_n2578_), .Y(new_n5154_));
  AOI21X1  g02718(.A0(new_n5141_), .A1(new_n5137_), .B0(new_n5154_), .Y(new_n5155_));
  OAI21X1  g02719(.A0(new_n5155_), .A1(new_n5121_), .B0(new_n2488_), .Y(new_n5156_));
  AOI21X1  g02720(.A0(new_n5156_), .A1(new_n5120_), .B0(pi0086), .Y(new_n5157_));
  NOR2X1   g02721(.A(new_n5157_), .B(new_n5145_), .Y(new_n5158_));
  INVX1    g02722(.A(new_n5158_), .Y(new_n5159_));
  AOI21X1  g02723(.A0(new_n5159_), .A1(new_n2678_), .B0(new_n5153_), .Y(new_n5160_));
  OAI21X1  g02724(.A0(new_n5160_), .A1(new_n5152_), .B0(new_n5150_), .Y(new_n5161_));
  OAI21X1  g02725(.A0(new_n5161_), .A1(new_n5148_), .B0(new_n2682_), .Y(new_n5162_));
  AOI21X1  g02726(.A0(new_n5162_), .A1(new_n5116_), .B0(pi0093), .Y(new_n5163_));
  NOR3X1   g02727(.A(new_n2505_), .B(new_n2502_), .C(new_n2705_), .Y(new_n5164_));
  OAI21X1  g02728(.A0(new_n5164_), .A1(new_n2516_), .B0(new_n2508_), .Y(new_n5165_));
  OAI21X1  g02729(.A0(new_n5165_), .A1(new_n5163_), .B0(new_n2535_), .Y(new_n5166_));
  AOI21X1  g02730(.A0(new_n5166_), .A1(new_n2874_), .B0(pi0072), .Y(new_n5167_));
  NOR3X1   g02731(.A(pi0095), .B(pi0040), .C(pi0032), .Y(new_n5168_));
  AND2X1   g02732(.A(new_n5168_), .B(new_n2532_), .Y(new_n5169_));
  INVX1    g02733(.A(new_n5169_), .Y(new_n5170_));
  OAI21X1  g02734(.A0(new_n5170_), .A1(new_n5167_), .B0(new_n5115_), .Y(new_n5171_));
  INVX1    g02735(.A(new_n2517_), .Y(new_n5172_));
  OR4X1    g02736(.A(new_n2505_), .B(new_n2502_), .C(pi0841), .D(pi0093), .Y(new_n5173_));
  OR4X1    g02737(.A(new_n5173_), .B(new_n2747_), .C(new_n5172_), .D(new_n2455_), .Y(new_n5174_));
  NOR3X1   g02738(.A(new_n5174_), .B(pi0210), .C(pi0095), .Y(new_n5175_));
  OR2X1    g02739(.A(new_n5175_), .B(new_n5171_), .Y(new_n5176_));
  NOR3X1   g02740(.A(pi0110), .B(pi0109), .C(pi0047), .Y(new_n5177_));
  OAI21X1  g02741(.A0(new_n5146_), .A1(new_n2677_), .B0(new_n5177_), .Y(new_n5178_));
  AND3X1   g02742(.A(new_n5178_), .B(new_n5117_), .C(new_n2515_), .Y(new_n5179_));
  INVX1    g02743(.A(new_n2677_), .Y(new_n5180_));
  INVX1    g02744(.A(new_n5177_), .Y(new_n5181_));
  AOI21X1  g02745(.A0(new_n5159_), .A1(new_n5180_), .B0(new_n5181_), .Y(new_n5182_));
  OAI21X1  g02746(.A0(new_n5182_), .A1(new_n5152_), .B0(new_n5150_), .Y(new_n5183_));
  OAI21X1  g02747(.A0(new_n5183_), .A1(new_n5179_), .B0(new_n2682_), .Y(new_n5184_));
  AOI21X1  g02748(.A0(new_n5184_), .A1(new_n5116_), .B0(pi0093), .Y(new_n5185_));
  OAI21X1  g02749(.A0(new_n5185_), .A1(new_n5165_), .B0(new_n2535_), .Y(new_n5186_));
  AOI21X1  g02750(.A0(new_n5186_), .A1(new_n2874_), .B0(pi0072), .Y(new_n5187_));
  OAI21X1  g02751(.A0(new_n5187_), .A1(new_n5170_), .B0(new_n5115_), .Y(new_n5188_));
  OR2X1    g02752(.A(new_n5188_), .B(new_n5175_), .Y(new_n5189_));
  AND2X1   g02753(.A(new_n5189_), .B(new_n5023_), .Y(new_n5190_));
  AOI21X1  g02754(.A0(new_n5176_), .A1(new_n5048_), .B0(new_n5190_), .Y(new_n5191_));
  OAI21X1  g02755(.A0(new_n5191_), .A1(new_n5112_), .B0(new_n5114_), .Y(new_n5192_));
  INVX1    g02756(.A(new_n5114_), .Y(new_n5193_));
  OAI21X1  g02757(.A0(new_n5175_), .A1(new_n5171_), .B0(new_n5105_), .Y(new_n5194_));
  AOI21X1  g02758(.A0(new_n5194_), .A1(new_n5193_), .B0(pi0228), .Y(new_n5195_));
  AOI21X1  g02759(.A0(new_n5195_), .A1(new_n5192_), .B0(new_n5111_), .Y(new_n5196_));
  MX2X1    g02760(.A(pi0602), .B(new_n5020_), .S0(new_n5048_), .Y(new_n5197_));
  NOR3X1   g02761(.A(new_n5174_), .B(pi0198), .C(pi0095), .Y(new_n5198_));
  OR2X1    g02762(.A(new_n5198_), .B(new_n5171_), .Y(new_n5199_));
  MX2X1    g02763(.A(new_n5199_), .B(pi0030), .S0(pi0228), .Y(new_n5200_));
  AOI21X1  g02764(.A0(new_n5200_), .A1(new_n5197_), .B0(pi0299), .Y(new_n5201_));
  INVX1    g02765(.A(pi0145), .Y(new_n5202_));
  INVX1    g02766(.A(pi0180), .Y(new_n5203_));
  INVX1    g02767(.A(pi0181), .Y(new_n5204_));
  INVX1    g02768(.A(pi0182), .Y(new_n5205_));
  NOR4X1   g02769(.A(new_n5205_), .B(new_n5204_), .C(new_n5203_), .D(new_n5202_), .Y(new_n5206_));
  AOI21X1  g02770(.A0(new_n5206_), .A1(new_n2933_), .B0(new_n5201_), .Y(new_n5207_));
  INVX1    g02771(.A(new_n5206_), .Y(new_n5208_));
  NAND2X1  g02772(.A(new_n5197_), .B(new_n5106_), .Y(new_n5209_));
  OR2X1    g02773(.A(new_n5198_), .B(new_n5188_), .Y(new_n5210_));
  MX2X1    g02774(.A(new_n5210_), .B(new_n5199_), .S0(new_n5048_), .Y(new_n5211_));
  NAND3X1  g02775(.A(new_n5211_), .B(new_n5197_), .C(new_n2793_), .Y(new_n5212_));
  AOI21X1  g02776(.A0(new_n5212_), .A1(new_n5209_), .B0(new_n5208_), .Y(new_n5213_));
  OAI21X1  g02777(.A0(new_n5213_), .A1(new_n5207_), .B0(pi0232), .Y(new_n5214_));
  INVX1    g02778(.A(pi0232), .Y(new_n5215_));
  NOR2X1   g02779(.A(new_n5194_), .B(pi0228), .Y(new_n5216_));
  OAI21X1  g02780(.A0(new_n5216_), .A1(new_n5111_), .B0(new_n5215_), .Y(new_n5217_));
  OAI22X1  g02781(.A0(new_n5217_), .A1(new_n5201_), .B0(new_n5214_), .B1(new_n5196_), .Y(new_n5218_));
  INVX1    g02782(.A(new_n5106_), .Y(new_n5219_));
  AND2X1   g02783(.A(pi0221), .B(new_n2934_), .Y(new_n5220_));
  INVX1    g02784(.A(new_n5220_), .Y(new_n5221_));
  INVX1    g02785(.A(pi0984), .Y(new_n5222_));
  NAND4X1  g02786(.A(new_n5027_), .B(new_n5222_), .C(new_n5026_), .D(pi0835), .Y(new_n5223_));
  OR4X1    g02787(.A(new_n5223_), .B(new_n2985_), .C(new_n2536_), .D(pi0287), .Y(new_n5224_));
  AND2X1   g02788(.A(pi1092), .B(pi0950), .Y(new_n5225_));
  AND2X1   g02789(.A(pi1093), .B(pi0824), .Y(new_n5226_));
  AND2X1   g02790(.A(new_n5226_), .B(new_n5225_), .Y(new_n5227_));
  INVX1    g02791(.A(new_n5227_), .Y(new_n5228_));
  NOR3X1   g02792(.A(new_n5228_), .B(new_n5224_), .C(pi1091), .Y(new_n5229_));
  INVX1    g02793(.A(new_n5225_), .Y(new_n5230_));
  INVX1    g02794(.A(new_n5226_), .Y(new_n5231_));
  AND3X1   g02795(.A(pi1091), .B(pi0957), .C(new_n2701_), .Y(new_n5232_));
  OR3X1    g02796(.A(new_n5232_), .B(new_n5231_), .C(new_n5230_), .Y(new_n5233_));
  AND2X1   g02797(.A(new_n5233_), .B(new_n2831_), .Y(new_n5234_));
  NOR3X1   g02798(.A(new_n5234_), .B(new_n5224_), .C(new_n2702_), .Y(new_n5235_));
  NOR2X1   g02799(.A(new_n5235_), .B(new_n5229_), .Y(new_n5236_));
  INVX1    g02800(.A(pi0829), .Y(new_n5237_));
  OAI21X1  g02801(.A0(new_n2758_), .A1(pi0833), .B0(new_n5237_), .Y(new_n5238_));
  AND2X1   g02802(.A(new_n5238_), .B(pi1091), .Y(new_n5239_));
  NOR3X1   g02803(.A(new_n5239_), .B(new_n5228_), .C(new_n5224_), .Y(new_n5240_));
  INVX1    g02804(.A(new_n5240_), .Y(new_n5241_));
  MX2X1    g02805(.A(new_n5241_), .B(new_n5236_), .S0(pi0216), .Y(new_n5242_));
  OR2X1    g02806(.A(new_n5242_), .B(pi0228), .Y(new_n5243_));
  OAI21X1  g02807(.A0(new_n5243_), .A1(new_n5221_), .B0(new_n5219_), .Y(new_n5244_));
  AOI21X1  g02808(.A0(new_n5244_), .A1(new_n5105_), .B0(new_n2933_), .Y(new_n5245_));
  NOR3X1   g02809(.A(new_n5235_), .B(new_n5229_), .C(new_n2942_), .Y(new_n5246_));
  AND2X1   g02810(.A(new_n2940_), .B(pi0222), .Y(new_n5247_));
  INVX1    g02811(.A(new_n5247_), .Y(new_n5248_));
  NOR2X1   g02812(.A(new_n5240_), .B(pi0224), .Y(new_n5249_));
  OR3X1    g02813(.A(new_n5249_), .B(new_n5248_), .C(new_n5246_), .Y(new_n5250_));
  OAI21X1  g02814(.A0(new_n5250_), .A1(pi0228), .B0(new_n5219_), .Y(new_n5251_));
  AOI21X1  g02815(.A0(new_n5251_), .A1(new_n5197_), .B0(pi0299), .Y(new_n5252_));
  OR2X1    g02816(.A(new_n5252_), .B(new_n2939_), .Y(new_n5253_));
  OAI21X1  g02817(.A0(new_n5253_), .A1(new_n5245_), .B0(new_n2979_), .Y(new_n5254_));
  AOI21X1  g02818(.A0(new_n5218_), .A1(new_n2939_), .B0(new_n5254_), .Y(new_n5255_));
  INVX1    g02819(.A(new_n5197_), .Y(new_n5256_));
  MX2X1    g02820(.A(new_n5256_), .B(new_n5112_), .S0(pi0299), .Y(new_n5257_));
  NOR3X1   g02821(.A(new_n5257_), .B(new_n5107_), .C(pi0039), .Y(new_n5258_));
  NOR2X1   g02822(.A(new_n5257_), .B(new_n5219_), .Y(new_n5259_));
  NOR3X1   g02823(.A(new_n5259_), .B(new_n5258_), .C(new_n2979_), .Y(new_n5260_));
  OAI21X1  g02824(.A0(new_n5260_), .A1(new_n5255_), .B0(new_n3007_), .Y(new_n5261_));
  INVX1    g02825(.A(new_n5020_), .Y(new_n5262_));
  NOR4X1   g02826(.A(new_n5086_), .B(new_n5082_), .C(new_n2986_), .D(new_n5077_), .Y(new_n5263_));
  INVX1    g02827(.A(new_n5263_), .Y(new_n5264_));
  AOI21X1  g02828(.A0(new_n5048_), .A1(new_n5262_), .B0(new_n5264_), .Y(new_n5265_));
  NAND2X1  g02829(.A(new_n5265_), .B(new_n5069_), .Y(new_n5266_));
  NOR2X1   g02830(.A(new_n5069_), .B(new_n3035_), .Y(new_n5267_));
  INVX1    g02831(.A(new_n5267_), .Y(new_n5268_));
  AND3X1   g02832(.A(new_n5023_), .B(new_n2982_), .C(pi0252), .Y(new_n5269_));
  NOR4X1   g02833(.A(new_n5262_), .B(new_n2985_), .C(new_n2536_), .D(new_n3035_), .Y(new_n5270_));
  AOI21X1  g02834(.A0(new_n5269_), .A1(new_n5262_), .B0(new_n5270_), .Y(new_n5271_));
  OAI21X1  g02835(.A0(new_n5271_), .A1(new_n5268_), .B0(new_n5266_), .Y(new_n5272_));
  INVX1    g02836(.A(pi0602), .Y(new_n5273_));
  AOI21X1  g02837(.A0(new_n5023_), .A1(new_n5273_), .B0(pi0228), .Y(new_n5274_));
  NAND2X1  g02838(.A(new_n5209_), .B(new_n2933_), .Y(new_n5275_));
  AOI21X1  g02839(.A0(new_n5274_), .A1(new_n5272_), .B0(new_n5275_), .Y(new_n5276_));
  INVX1    g02840(.A(pi0907), .Y(new_n5277_));
  AOI21X1  g02841(.A0(new_n5023_), .A1(new_n5277_), .B0(pi0228), .Y(new_n5278_));
  OAI21X1  g02842(.A0(new_n5265_), .A1(new_n3038_), .B0(new_n5278_), .Y(new_n5279_));
  AOI21X1  g02843(.A0(new_n5271_), .A1(new_n3038_), .B0(new_n5279_), .Y(new_n5280_));
  OAI21X1  g02844(.A0(new_n5280_), .A1(new_n5111_), .B0(new_n3047_), .Y(new_n5281_));
  AOI21X1  g02845(.A0(new_n5259_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n5282_));
  OAI21X1  g02846(.A0(new_n5281_), .A1(new_n5276_), .B0(new_n5282_), .Y(new_n5283_));
  AND2X1   g02847(.A(new_n5283_), .B(new_n3131_), .Y(new_n5284_));
  INVX1    g02848(.A(new_n5259_), .Y(new_n5285_));
  OAI21X1  g02849(.A0(new_n5285_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n5286_));
  AOI21X1  g02850(.A0(new_n5284_), .A1(new_n5261_), .B0(new_n5286_), .Y(new_n5287_));
  AOI22X1  g02851(.A0(new_n5259_), .A1(new_n3074_), .B0(new_n5258_), .B1(new_n3087_), .Y(new_n5288_));
  AND2X1   g02852(.A(new_n5288_), .B(pi0075), .Y(new_n5289_));
  OR2X1    g02853(.A(new_n5289_), .B(pi0092), .Y(new_n5290_));
  NAND2X1  g02854(.A(new_n5288_), .B(new_n3073_), .Y(new_n5291_));
  AOI21X1  g02855(.A0(new_n5285_), .A1(pi0075), .B0(new_n3079_), .Y(new_n5292_));
  AOI21X1  g02856(.A0(new_n5292_), .A1(new_n5291_), .B0(pi0054), .Y(new_n5293_));
  OAI21X1  g02857(.A0(new_n5290_), .A1(new_n5287_), .B0(new_n5293_), .Y(new_n5294_));
  INVX1    g02858(.A(new_n3084_), .Y(new_n5295_));
  MX2X1    g02859(.A(new_n5288_), .B(new_n5285_), .S0(new_n5295_), .Y(new_n5296_));
  AOI21X1  g02860(.A0(new_n5296_), .A1(pi0054), .B0(pi0074), .Y(new_n5297_));
  AND3X1   g02861(.A(new_n5288_), .B(new_n3084_), .C(new_n3091_), .Y(new_n5298_));
  NOR3X1   g02862(.A(pi0092), .B(pi0075), .C(pi0054), .Y(new_n5299_));
  OAI21X1  g02863(.A0(new_n5299_), .A1(new_n5259_), .B0(pi0074), .Y(new_n5300_));
  OAI21X1  g02864(.A0(new_n5300_), .A1(new_n5298_), .B0(new_n3107_), .Y(new_n5301_));
  AOI21X1  g02865(.A0(new_n5297_), .A1(new_n5294_), .B0(new_n5301_), .Y(new_n5302_));
  OAI21X1  g02866(.A0(new_n5109_), .A1(new_n3107_), .B0(new_n3123_), .Y(new_n5303_));
  AOI21X1  g02867(.A0(new_n5110_), .A1(new_n4975_), .B0(pi0059), .Y(new_n5304_));
  OAI21X1  g02868(.A0(new_n5303_), .A1(new_n5302_), .B0(new_n5304_), .Y(new_n5305_));
  NOR3X1   g02869(.A(pi0062), .B(pi0056), .C(pi0055), .Y(new_n5306_));
  OAI21X1  g02870(.A0(new_n5306_), .A1(pi0228), .B0(new_n5109_), .Y(new_n5307_));
  AOI21X1  g02871(.A0(new_n5307_), .A1(pi0059), .B0(pi0057), .Y(new_n5308_));
  AOI22X1  g02872(.A0(new_n5308_), .A1(new_n5305_), .B0(new_n5109_), .B1(new_n5104_), .Y(po0171));
  MX2X1    g02873(.A(new_n5018_), .B(pi0947), .S0(new_n5023_), .Y(new_n5310_));
  AND2X1   g02874(.A(new_n5310_), .B(new_n5108_), .Y(new_n5311_));
  AOI21X1  g02875(.A0(new_n5310_), .A1(new_n5106_), .B0(new_n2933_), .Y(new_n5312_));
  INVX1    g02876(.A(new_n5312_), .Y(new_n5313_));
  INVX1    g02877(.A(new_n5310_), .Y(new_n5314_));
  OAI21X1  g02878(.A0(new_n5314_), .A1(new_n5191_), .B0(new_n5114_), .Y(new_n5315_));
  OAI21X1  g02879(.A0(new_n5175_), .A1(new_n5171_), .B0(new_n5310_), .Y(new_n5316_));
  AOI21X1  g02880(.A0(new_n5316_), .A1(new_n5193_), .B0(pi0228), .Y(new_n5317_));
  AOI21X1  g02881(.A0(new_n5317_), .A1(new_n5315_), .B0(new_n5313_), .Y(new_n5318_));
  MX2X1    g02882(.A(new_n5018_), .B(pi0587), .S0(new_n5023_), .Y(new_n5319_));
  NAND2X1  g02883(.A(new_n5319_), .B(new_n5106_), .Y(new_n5320_));
  NAND3X1  g02884(.A(new_n5319_), .B(new_n5211_), .C(new_n2793_), .Y(new_n5321_));
  AOI21X1  g02885(.A0(new_n5321_), .A1(new_n5320_), .B0(new_n5208_), .Y(new_n5322_));
  AND3X1   g02886(.A(new_n5319_), .B(new_n5208_), .C(new_n5200_), .Y(new_n5323_));
  OR2X1    g02887(.A(new_n5323_), .B(pi0299), .Y(new_n5324_));
  OAI21X1  g02888(.A0(new_n5324_), .A1(new_n5322_), .B0(pi0232), .Y(new_n5325_));
  AOI21X1  g02889(.A0(new_n5319_), .A1(new_n5200_), .B0(pi0299), .Y(new_n5326_));
  OAI21X1  g02890(.A0(new_n5316_), .A1(pi0228), .B0(new_n5312_), .Y(new_n5327_));
  NAND2X1  g02891(.A(new_n5327_), .B(new_n5215_), .Y(new_n5328_));
  OAI22X1  g02892(.A0(new_n5328_), .A1(new_n5326_), .B0(new_n5325_), .B1(new_n5318_), .Y(new_n5329_));
  AOI21X1  g02893(.A0(new_n5243_), .A1(new_n5219_), .B0(new_n5221_), .Y(new_n5330_));
  AND3X1   g02894(.A(pi0299), .B(pi0221), .C(new_n2934_), .Y(new_n5331_));
  NOR2X1   g02895(.A(new_n5331_), .B(new_n5312_), .Y(new_n5332_));
  AOI21X1  g02896(.A0(new_n5310_), .A1(new_n5330_), .B0(new_n5332_), .Y(new_n5333_));
  AOI21X1  g02897(.A0(new_n5319_), .A1(new_n5251_), .B0(pi0299), .Y(new_n5334_));
  OR2X1    g02898(.A(new_n5334_), .B(new_n2939_), .Y(new_n5335_));
  OAI21X1  g02899(.A0(new_n5335_), .A1(new_n5333_), .B0(new_n2979_), .Y(new_n5336_));
  AOI21X1  g02900(.A0(new_n5329_), .A1(new_n2939_), .B0(new_n5336_), .Y(new_n5337_));
  NOR2X1   g02901(.A(new_n5310_), .B(new_n2933_), .Y(new_n5338_));
  NOR2X1   g02902(.A(new_n5319_), .B(pi0299), .Y(new_n5339_));
  OR2X1    g02903(.A(new_n5339_), .B(new_n5338_), .Y(new_n5340_));
  NOR3X1   g02904(.A(new_n5340_), .B(new_n5107_), .C(pi0039), .Y(new_n5341_));
  NOR3X1   g02905(.A(new_n5339_), .B(new_n5338_), .C(new_n5219_), .Y(new_n5342_));
  NOR3X1   g02906(.A(new_n5342_), .B(new_n5341_), .C(new_n2979_), .Y(new_n5343_));
  OAI21X1  g02907(.A0(new_n5343_), .A1(new_n5337_), .B0(new_n3007_), .Y(new_n5344_));
  NOR3X1   g02908(.A(pi0587), .B(pi0468), .C(pi0332), .Y(new_n5345_));
  INVX1    g02909(.A(new_n5345_), .Y(new_n5346_));
  OR4X1    g02910(.A(pi0228), .B(pi0189), .C(pi0174), .D(pi0144), .Y(new_n5347_));
  INVX1    g02911(.A(new_n5018_), .Y(new_n5348_));
  NOR3X1   g02912(.A(new_n2985_), .B(new_n2536_), .C(new_n3035_), .Y(new_n5349_));
  MX2X1    g02913(.A(new_n5349_), .B(new_n5269_), .S0(new_n5348_), .Y(new_n5350_));
  AOI21X1  g02914(.A0(new_n5350_), .A1(new_n5346_), .B0(new_n5347_), .Y(new_n5351_));
  NOR2X1   g02915(.A(new_n5023_), .B(new_n5018_), .Y(new_n5352_));
  OAI21X1  g02916(.A0(new_n5264_), .A1(new_n5352_), .B0(new_n2953_), .Y(new_n5353_));
  INVX1    g02917(.A(pi0587), .Y(new_n5354_));
  OAI21X1  g02918(.A0(new_n5023_), .A1(new_n5348_), .B0(new_n5354_), .Y(new_n5355_));
  AND3X1   g02919(.A(new_n5355_), .B(new_n5353_), .C(new_n2793_), .Y(new_n5356_));
  OAI21X1  g02920(.A0(new_n5350_), .A1(new_n2953_), .B0(new_n5356_), .Y(new_n5357_));
  AOI22X1  g02921(.A0(new_n5319_), .A1(new_n5106_), .B0(new_n2961_), .B1(new_n2793_), .Y(new_n5358_));
  AOI21X1  g02922(.A0(new_n5358_), .A1(new_n5357_), .B0(new_n5351_), .Y(new_n5359_));
  NOR3X1   g02923(.A(pi0947), .B(pi0468), .C(pi0332), .Y(new_n5360_));
  NOR4X1   g02924(.A(new_n5360_), .B(new_n5264_), .C(new_n5352_), .D(new_n3038_), .Y(new_n5361_));
  INVX1    g02925(.A(pi0947), .Y(new_n5362_));
  OAI21X1  g02926(.A0(new_n5023_), .A1(new_n5348_), .B0(new_n5362_), .Y(new_n5363_));
  AND3X1   g02927(.A(new_n5363_), .B(new_n5350_), .C(new_n3038_), .Y(new_n5364_));
  OAI21X1  g02928(.A0(new_n5364_), .A1(new_n5361_), .B0(new_n2793_), .Y(new_n5365_));
  AOI21X1  g02929(.A0(new_n5365_), .A1(new_n5312_), .B0(new_n3060_), .Y(new_n5366_));
  OAI21X1  g02930(.A0(new_n5359_), .A1(pi0299), .B0(new_n5366_), .Y(new_n5367_));
  AOI21X1  g02931(.A0(new_n5342_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n5368_));
  AOI21X1  g02932(.A0(new_n5368_), .A1(new_n5367_), .B0(pi0087), .Y(new_n5369_));
  INVX1    g02933(.A(new_n5342_), .Y(new_n5370_));
  OAI21X1  g02934(.A0(new_n5370_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n5371_));
  AOI21X1  g02935(.A0(new_n5369_), .A1(new_n5344_), .B0(new_n5371_), .Y(new_n5372_));
  AOI22X1  g02936(.A0(new_n5342_), .A1(new_n3074_), .B0(new_n5341_), .B1(new_n3087_), .Y(new_n5373_));
  AND2X1   g02937(.A(new_n5373_), .B(pi0075), .Y(new_n5374_));
  OR2X1    g02938(.A(new_n5374_), .B(pi0092), .Y(new_n5375_));
  NAND2X1  g02939(.A(new_n5373_), .B(new_n3073_), .Y(new_n5376_));
  AOI21X1  g02940(.A0(new_n5370_), .A1(pi0075), .B0(new_n3079_), .Y(new_n5377_));
  AOI21X1  g02941(.A0(new_n5377_), .A1(new_n5376_), .B0(pi0054), .Y(new_n5378_));
  OAI21X1  g02942(.A0(new_n5375_), .A1(new_n5372_), .B0(new_n5378_), .Y(new_n5379_));
  MX2X1    g02943(.A(new_n5373_), .B(new_n5370_), .S0(new_n5295_), .Y(new_n5380_));
  AOI21X1  g02944(.A0(new_n5380_), .A1(pi0054), .B0(pi0074), .Y(new_n5381_));
  AND3X1   g02945(.A(new_n5373_), .B(new_n3084_), .C(new_n3091_), .Y(new_n5382_));
  OAI21X1  g02946(.A0(new_n5342_), .A1(new_n5299_), .B0(pi0074), .Y(new_n5383_));
  OAI21X1  g02947(.A0(new_n5383_), .A1(new_n5382_), .B0(new_n3107_), .Y(new_n5384_));
  AOI21X1  g02948(.A0(new_n5381_), .A1(new_n5379_), .B0(new_n5384_), .Y(new_n5385_));
  OAI21X1  g02949(.A0(new_n5311_), .A1(new_n3107_), .B0(new_n3123_), .Y(new_n5386_));
  NAND3X1  g02950(.A(new_n5310_), .B(new_n5106_), .C(new_n4975_), .Y(new_n5387_));
  AND2X1   g02951(.A(new_n5387_), .B(new_n3127_), .Y(new_n5388_));
  OAI21X1  g02952(.A0(new_n5386_), .A1(new_n5385_), .B0(new_n5388_), .Y(new_n5389_));
  OAI21X1  g02953(.A0(new_n5306_), .A1(pi0228), .B0(new_n5311_), .Y(new_n5390_));
  AOI21X1  g02954(.A0(new_n5390_), .A1(pi0059), .B0(pi0057), .Y(new_n5391_));
  AOI22X1  g02955(.A0(new_n5391_), .A1(new_n5389_), .B0(new_n5311_), .B1(new_n5104_), .Y(po0172));
  INVX1    g02956(.A(pi0970), .Y(new_n5393_));
  AND3X1   g02957(.A(new_n5023_), .B(pi0228), .C(pi0030), .Y(new_n5394_));
  INVX1    g02958(.A(new_n5394_), .Y(new_n5395_));
  AND2X1   g02959(.A(pi0970), .B(new_n2793_), .Y(new_n5396_));
  NAND4X1  g02960(.A(new_n5396_), .B(new_n5102_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5397_));
  OAI21X1  g02961(.A0(new_n5395_), .A1(new_n5393_), .B0(new_n5397_), .Y(new_n5398_));
  AOI21X1  g02962(.A0(new_n5394_), .A1(pi0970), .B0(new_n2933_), .Y(new_n5399_));
  INVX1    g02963(.A(new_n5399_), .Y(new_n5400_));
  AND2X1   g02964(.A(new_n5176_), .B(new_n5023_), .Y(new_n5401_));
  AOI21X1  g02965(.A0(new_n5401_), .A1(new_n5396_), .B0(new_n5400_), .Y(new_n5402_));
  AOI21X1  g02966(.A0(new_n5113_), .A1(pi0299), .B0(new_n5402_), .Y(new_n5403_));
  AND2X1   g02967(.A(new_n5394_), .B(pi0970), .Y(new_n5404_));
  NAND2X1  g02968(.A(pi0197), .B(pi0160), .Y(new_n5405_));
  MX2X1    g02969(.A(new_n5190_), .B(new_n5176_), .S0(new_n5405_), .Y(new_n5406_));
  AND3X1   g02970(.A(new_n5406_), .B(new_n5396_), .C(new_n5023_), .Y(new_n5407_));
  OR2X1    g02971(.A(new_n5407_), .B(new_n5404_), .Y(new_n5408_));
  AOI21X1  g02972(.A0(new_n5408_), .A1(new_n5113_), .B0(new_n5403_), .Y(new_n5409_));
  AOI21X1  g02973(.A0(new_n5200_), .A1(new_n5023_), .B0(new_n5206_), .Y(new_n5410_));
  NAND3X1  g02974(.A(new_n5210_), .B(new_n5023_), .C(new_n2793_), .Y(new_n5411_));
  OAI21X1  g02975(.A0(new_n5198_), .A1(new_n5171_), .B0(new_n5208_), .Y(new_n5412_));
  AND2X1   g02976(.A(new_n5412_), .B(new_n5395_), .Y(new_n5413_));
  AOI21X1  g02977(.A0(new_n5413_), .A1(new_n5411_), .B0(new_n5410_), .Y(new_n5414_));
  AOI21X1  g02978(.A0(new_n5414_), .A1(pi0967), .B0(pi0299), .Y(new_n5415_));
  OR2X1    g02979(.A(new_n5415_), .B(new_n5215_), .Y(new_n5416_));
  AND2X1   g02980(.A(new_n5200_), .B(new_n5023_), .Y(new_n5417_));
  AOI21X1  g02981(.A0(new_n5417_), .A1(pi0967), .B0(pi0299), .Y(new_n5418_));
  OR3X1    g02982(.A(new_n5418_), .B(new_n5402_), .C(pi0232), .Y(new_n5419_));
  OAI21X1  g02983(.A0(new_n5416_), .A1(new_n5409_), .B0(new_n5419_), .Y(new_n5420_));
  AND2X1   g02984(.A(pi0970), .B(pi0299), .Y(new_n5421_));
  NOR3X1   g02985(.A(new_n5242_), .B(new_n5221_), .C(new_n5048_), .Y(new_n5422_));
  OR2X1    g02986(.A(new_n5422_), .B(pi0228), .Y(new_n5423_));
  AND2X1   g02987(.A(pi0967), .B(new_n2933_), .Y(new_n5424_));
  OAI21X1  g02988(.A0(new_n5250_), .A1(new_n5048_), .B0(new_n2793_), .Y(new_n5425_));
  AOI22X1  g02989(.A0(new_n5425_), .A1(new_n5424_), .B0(new_n5423_), .B1(new_n5421_), .Y(new_n5426_));
  AOI21X1  g02990(.A0(new_n5023_), .A1(pi0030), .B0(new_n2793_), .Y(new_n5427_));
  OR2X1    g02991(.A(new_n5427_), .B(new_n2939_), .Y(new_n5428_));
  OAI21X1  g02992(.A0(new_n5428_), .A1(new_n5426_), .B0(new_n2979_), .Y(new_n5429_));
  AOI21X1  g02993(.A0(new_n5420_), .A1(new_n2939_), .B0(new_n5429_), .Y(new_n5430_));
  INVX1    g02994(.A(new_n5037_), .Y(new_n5431_));
  AOI21X1  g02995(.A0(new_n5431_), .A1(new_n2793_), .B0(new_n5427_), .Y(new_n5432_));
  AOI21X1  g02996(.A0(new_n5432_), .A1(pi0967), .B0(pi0299), .Y(new_n5433_));
  AOI21X1  g02997(.A0(new_n5396_), .A1(new_n5037_), .B0(new_n5400_), .Y(new_n5434_));
  NOR3X1   g02998(.A(new_n5434_), .B(new_n5433_), .C(pi0039), .Y(new_n5435_));
  OAI21X1  g02999(.A0(new_n5424_), .A1(new_n5421_), .B0(new_n5394_), .Y(new_n5436_));
  OAI21X1  g03000(.A0(new_n5436_), .A1(new_n2939_), .B0(pi0038), .Y(new_n5437_));
  NOR2X1   g03001(.A(new_n5437_), .B(new_n5435_), .Y(new_n5438_));
  OAI21X1  g03002(.A0(new_n5438_), .A1(new_n5430_), .B0(new_n3007_), .Y(new_n5439_));
  AND2X1   g03003(.A(new_n5269_), .B(new_n5070_), .Y(new_n5440_));
  AND3X1   g03004(.A(new_n5263_), .B(new_n5069_), .C(new_n5023_), .Y(new_n5441_));
  NOR3X1   g03005(.A(new_n5441_), .B(new_n5440_), .C(pi0228), .Y(new_n5442_));
  NOR2X1   g03006(.A(new_n5442_), .B(new_n5427_), .Y(new_n5443_));
  AOI21X1  g03007(.A0(new_n5443_), .A1(pi0967), .B0(pi0299), .Y(new_n5444_));
  NOR2X1   g03008(.A(new_n5269_), .B(new_n2815_), .Y(new_n5445_));
  AOI21X1  g03009(.A0(new_n5263_), .A1(new_n5023_), .B0(new_n3038_), .Y(new_n5446_));
  NOR4X1   g03010(.A(new_n5446_), .B(new_n5445_), .C(new_n5393_), .D(pi0228), .Y(new_n5447_));
  OAI21X1  g03011(.A0(new_n5447_), .A1(new_n5400_), .B0(new_n3047_), .Y(new_n5448_));
  INVX1    g03012(.A(new_n5436_), .Y(new_n5449_));
  AOI21X1  g03013(.A0(new_n5449_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n5450_));
  OAI21X1  g03014(.A0(new_n5448_), .A1(new_n5444_), .B0(new_n5450_), .Y(new_n5451_));
  AND2X1   g03015(.A(new_n5451_), .B(new_n3131_), .Y(new_n5452_));
  OAI21X1  g03016(.A0(new_n5436_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n5453_));
  AOI21X1  g03017(.A0(new_n5452_), .A1(new_n5439_), .B0(new_n5453_), .Y(new_n5454_));
  AOI22X1  g03018(.A0(new_n5449_), .A1(new_n3074_), .B0(new_n5435_), .B1(new_n3087_), .Y(new_n5455_));
  AND2X1   g03019(.A(new_n5455_), .B(pi0075), .Y(new_n5456_));
  OR2X1    g03020(.A(new_n5456_), .B(pi0092), .Y(new_n5457_));
  NAND2X1  g03021(.A(new_n5455_), .B(new_n3073_), .Y(new_n5458_));
  AOI21X1  g03022(.A0(new_n5436_), .A1(pi0075), .B0(new_n3079_), .Y(new_n5459_));
  AOI21X1  g03023(.A0(new_n5459_), .A1(new_n5458_), .B0(pi0054), .Y(new_n5460_));
  OAI21X1  g03024(.A0(new_n5457_), .A1(new_n5454_), .B0(new_n5460_), .Y(new_n5461_));
  MX2X1    g03025(.A(new_n5455_), .B(new_n5436_), .S0(new_n5295_), .Y(new_n5462_));
  AOI21X1  g03026(.A0(new_n5462_), .A1(pi0054), .B0(pi0074), .Y(new_n5463_));
  AND3X1   g03027(.A(new_n5455_), .B(new_n3084_), .C(new_n3091_), .Y(new_n5464_));
  OAI21X1  g03028(.A0(new_n5449_), .A1(new_n5299_), .B0(pi0074), .Y(new_n5465_));
  OAI21X1  g03029(.A0(new_n5465_), .A1(new_n5464_), .B0(new_n3107_), .Y(new_n5466_));
  AOI21X1  g03030(.A0(new_n5463_), .A1(new_n5461_), .B0(new_n5466_), .Y(new_n5467_));
  AND3X1   g03031(.A(new_n5396_), .B(new_n5037_), .C(new_n3104_), .Y(new_n5468_));
  OR2X1    g03032(.A(new_n5404_), .B(new_n3107_), .Y(new_n5469_));
  OAI21X1  g03033(.A0(new_n5469_), .A1(new_n5468_), .B0(new_n3123_), .Y(new_n5470_));
  AOI21X1  g03034(.A0(new_n5404_), .A1(new_n4975_), .B0(pi0059), .Y(new_n5471_));
  OAI21X1  g03035(.A0(new_n5470_), .A1(new_n5467_), .B0(new_n5471_), .Y(new_n5472_));
  NAND4X1  g03036(.A(new_n5396_), .B(new_n5306_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5473_));
  AOI21X1  g03037(.A0(new_n5394_), .A1(pi0970), .B0(new_n3127_), .Y(new_n5474_));
  AOI21X1  g03038(.A0(new_n5474_), .A1(new_n5473_), .B0(pi0057), .Y(new_n5475_));
  AOI22X1  g03039(.A0(new_n5475_), .A1(new_n5472_), .B0(new_n5398_), .B1(pi0057), .Y(po0173));
  INVX1    g03040(.A(pi0972), .Y(new_n5477_));
  AND2X1   g03041(.A(pi0972), .B(new_n2793_), .Y(new_n5478_));
  NAND4X1  g03042(.A(new_n5478_), .B(new_n5102_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5479_));
  OAI21X1  g03043(.A0(new_n5395_), .A1(new_n5477_), .B0(new_n5479_), .Y(new_n5480_));
  AOI21X1  g03044(.A0(new_n5394_), .A1(pi0972), .B0(new_n2933_), .Y(new_n5481_));
  INVX1    g03045(.A(new_n5481_), .Y(new_n5482_));
  AOI21X1  g03046(.A0(new_n5478_), .A1(new_n5401_), .B0(new_n5482_), .Y(new_n5483_));
  AOI21X1  g03047(.A0(new_n5113_), .A1(pi0299), .B0(new_n5483_), .Y(new_n5484_));
  AND2X1   g03048(.A(new_n5394_), .B(pi0972), .Y(new_n5485_));
  AND3X1   g03049(.A(new_n5478_), .B(new_n5406_), .C(new_n5023_), .Y(new_n5486_));
  OR2X1    g03050(.A(new_n5486_), .B(new_n5485_), .Y(new_n5487_));
  AOI21X1  g03051(.A0(new_n5487_), .A1(new_n5113_), .B0(new_n5484_), .Y(new_n5488_));
  AOI21X1  g03052(.A0(new_n5414_), .A1(pi0961), .B0(pi0299), .Y(new_n5489_));
  OR2X1    g03053(.A(new_n5489_), .B(new_n5215_), .Y(new_n5490_));
  AOI21X1  g03054(.A0(new_n5417_), .A1(pi0961), .B0(pi0299), .Y(new_n5491_));
  OR3X1    g03055(.A(new_n5491_), .B(new_n5483_), .C(pi0232), .Y(new_n5492_));
  OAI21X1  g03056(.A0(new_n5490_), .A1(new_n5488_), .B0(new_n5492_), .Y(new_n5493_));
  AND2X1   g03057(.A(pi0961), .B(new_n2933_), .Y(new_n5494_));
  AND2X1   g03058(.A(pi0972), .B(pi0299), .Y(new_n5495_));
  AOI22X1  g03059(.A0(new_n5495_), .A1(new_n5423_), .B0(new_n5494_), .B1(new_n5425_), .Y(new_n5496_));
  OAI21X1  g03060(.A0(new_n5496_), .A1(new_n5428_), .B0(new_n2979_), .Y(new_n5497_));
  AOI21X1  g03061(.A0(new_n5493_), .A1(new_n2939_), .B0(new_n5497_), .Y(new_n5498_));
  AOI21X1  g03062(.A0(new_n5432_), .A1(pi0961), .B0(pi0299), .Y(new_n5499_));
  AOI21X1  g03063(.A0(new_n5478_), .A1(new_n5037_), .B0(new_n5482_), .Y(new_n5500_));
  NOR3X1   g03064(.A(new_n5500_), .B(new_n5499_), .C(pi0039), .Y(new_n5501_));
  OAI21X1  g03065(.A0(new_n5495_), .A1(new_n5494_), .B0(new_n5394_), .Y(new_n5502_));
  OAI21X1  g03066(.A0(new_n5502_), .A1(new_n2939_), .B0(pi0038), .Y(new_n5503_));
  NOR2X1   g03067(.A(new_n5503_), .B(new_n5501_), .Y(new_n5504_));
  OAI21X1  g03068(.A0(new_n5504_), .A1(new_n5498_), .B0(new_n3007_), .Y(new_n5505_));
  AOI21X1  g03069(.A0(new_n5443_), .A1(pi0961), .B0(pi0299), .Y(new_n5506_));
  NOR4X1   g03070(.A(new_n5446_), .B(new_n5445_), .C(new_n5477_), .D(pi0228), .Y(new_n5507_));
  OAI21X1  g03071(.A0(new_n5507_), .A1(new_n5482_), .B0(new_n3047_), .Y(new_n5508_));
  INVX1    g03072(.A(new_n5502_), .Y(new_n5509_));
  AOI21X1  g03073(.A0(new_n5509_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n5510_));
  OAI21X1  g03074(.A0(new_n5508_), .A1(new_n5506_), .B0(new_n5510_), .Y(new_n5511_));
  AND2X1   g03075(.A(new_n5511_), .B(new_n3131_), .Y(new_n5512_));
  OAI21X1  g03076(.A0(new_n5502_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n5513_));
  AOI21X1  g03077(.A0(new_n5512_), .A1(new_n5505_), .B0(new_n5513_), .Y(new_n5514_));
  AOI22X1  g03078(.A0(new_n5509_), .A1(new_n3074_), .B0(new_n5501_), .B1(new_n3087_), .Y(new_n5515_));
  AND2X1   g03079(.A(new_n5515_), .B(pi0075), .Y(new_n5516_));
  OR2X1    g03080(.A(new_n5516_), .B(pi0092), .Y(new_n5517_));
  NAND2X1  g03081(.A(new_n5515_), .B(new_n3073_), .Y(new_n5518_));
  AOI21X1  g03082(.A0(new_n5502_), .A1(pi0075), .B0(new_n3079_), .Y(new_n5519_));
  AOI21X1  g03083(.A0(new_n5519_), .A1(new_n5518_), .B0(pi0054), .Y(new_n5520_));
  OAI21X1  g03084(.A0(new_n5517_), .A1(new_n5514_), .B0(new_n5520_), .Y(new_n5521_));
  MX2X1    g03085(.A(new_n5515_), .B(new_n5502_), .S0(new_n5295_), .Y(new_n5522_));
  AOI21X1  g03086(.A0(new_n5522_), .A1(pi0054), .B0(pi0074), .Y(new_n5523_));
  AND3X1   g03087(.A(new_n5515_), .B(new_n3084_), .C(new_n3091_), .Y(new_n5524_));
  OAI21X1  g03088(.A0(new_n5509_), .A1(new_n5299_), .B0(pi0074), .Y(new_n5525_));
  OAI21X1  g03089(.A0(new_n5525_), .A1(new_n5524_), .B0(new_n3107_), .Y(new_n5526_));
  AOI21X1  g03090(.A0(new_n5523_), .A1(new_n5521_), .B0(new_n5526_), .Y(new_n5527_));
  AND3X1   g03091(.A(new_n5478_), .B(new_n5037_), .C(new_n3104_), .Y(new_n5528_));
  OR2X1    g03092(.A(new_n5485_), .B(new_n3107_), .Y(new_n5529_));
  OAI21X1  g03093(.A0(new_n5529_), .A1(new_n5528_), .B0(new_n3123_), .Y(new_n5530_));
  AOI21X1  g03094(.A0(new_n5485_), .A1(new_n4975_), .B0(pi0059), .Y(new_n5531_));
  OAI21X1  g03095(.A0(new_n5530_), .A1(new_n5527_), .B0(new_n5531_), .Y(new_n5532_));
  NAND4X1  g03096(.A(new_n5478_), .B(new_n5306_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5533_));
  AOI21X1  g03097(.A0(new_n5394_), .A1(pi0972), .B0(new_n3127_), .Y(new_n5534_));
  AOI21X1  g03098(.A0(new_n5534_), .A1(new_n5533_), .B0(pi0057), .Y(new_n5535_));
  AOI22X1  g03099(.A0(new_n5535_), .A1(new_n5532_), .B0(new_n5480_), .B1(pi0057), .Y(po0174));
  INVX1    g03100(.A(pi0960), .Y(new_n5537_));
  AND2X1   g03101(.A(pi0960), .B(new_n2793_), .Y(new_n5538_));
  NAND4X1  g03102(.A(new_n5538_), .B(new_n5102_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5539_));
  OAI21X1  g03103(.A0(new_n5395_), .A1(new_n5537_), .B0(new_n5539_), .Y(new_n5540_));
  AOI21X1  g03104(.A0(new_n5394_), .A1(pi0960), .B0(new_n2933_), .Y(new_n5541_));
  INVX1    g03105(.A(new_n5541_), .Y(new_n5542_));
  AOI21X1  g03106(.A0(new_n5538_), .A1(new_n5401_), .B0(new_n5542_), .Y(new_n5543_));
  AOI21X1  g03107(.A0(new_n5113_), .A1(pi0299), .B0(new_n5543_), .Y(new_n5544_));
  AND2X1   g03108(.A(new_n5394_), .B(pi0960), .Y(new_n5545_));
  AND3X1   g03109(.A(new_n5538_), .B(new_n5406_), .C(new_n5023_), .Y(new_n5546_));
  OR2X1    g03110(.A(new_n5546_), .B(new_n5545_), .Y(new_n5547_));
  AOI21X1  g03111(.A0(new_n5547_), .A1(new_n5113_), .B0(new_n5544_), .Y(new_n5548_));
  AOI21X1  g03112(.A0(new_n5414_), .A1(pi0977), .B0(pi0299), .Y(new_n5549_));
  OR2X1    g03113(.A(new_n5549_), .B(new_n5215_), .Y(new_n5550_));
  AOI21X1  g03114(.A0(new_n5417_), .A1(pi0977), .B0(pi0299), .Y(new_n5551_));
  OR3X1    g03115(.A(new_n5551_), .B(new_n5543_), .C(pi0232), .Y(new_n5552_));
  OAI21X1  g03116(.A0(new_n5550_), .A1(new_n5548_), .B0(new_n5552_), .Y(new_n5553_));
  AND2X1   g03117(.A(pi0977), .B(new_n2933_), .Y(new_n5554_));
  AND2X1   g03118(.A(pi0960), .B(pi0299), .Y(new_n5555_));
  AOI22X1  g03119(.A0(new_n5555_), .A1(new_n5423_), .B0(new_n5554_), .B1(new_n5425_), .Y(new_n5556_));
  OAI21X1  g03120(.A0(new_n5556_), .A1(new_n5428_), .B0(new_n2979_), .Y(new_n5557_));
  AOI21X1  g03121(.A0(new_n5553_), .A1(new_n2939_), .B0(new_n5557_), .Y(new_n5558_));
  AOI21X1  g03122(.A0(new_n5432_), .A1(pi0977), .B0(pi0299), .Y(new_n5559_));
  AOI21X1  g03123(.A0(new_n5538_), .A1(new_n5037_), .B0(new_n5542_), .Y(new_n5560_));
  NOR3X1   g03124(.A(new_n5560_), .B(new_n5559_), .C(pi0039), .Y(new_n5561_));
  OAI21X1  g03125(.A0(new_n5555_), .A1(new_n5554_), .B0(new_n5394_), .Y(new_n5562_));
  OAI21X1  g03126(.A0(new_n5562_), .A1(new_n2939_), .B0(pi0038), .Y(new_n5563_));
  NOR2X1   g03127(.A(new_n5563_), .B(new_n5561_), .Y(new_n5564_));
  OAI21X1  g03128(.A0(new_n5564_), .A1(new_n5558_), .B0(new_n3007_), .Y(new_n5565_));
  AOI21X1  g03129(.A0(new_n5443_), .A1(pi0977), .B0(pi0299), .Y(new_n5566_));
  NOR4X1   g03130(.A(new_n5446_), .B(new_n5445_), .C(new_n5537_), .D(pi0228), .Y(new_n5567_));
  OAI21X1  g03131(.A0(new_n5567_), .A1(new_n5542_), .B0(new_n3047_), .Y(new_n5568_));
  INVX1    g03132(.A(new_n5562_), .Y(new_n5569_));
  AOI21X1  g03133(.A0(new_n5569_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n5570_));
  OAI21X1  g03134(.A0(new_n5568_), .A1(new_n5566_), .B0(new_n5570_), .Y(new_n5571_));
  AND2X1   g03135(.A(new_n5571_), .B(new_n3131_), .Y(new_n5572_));
  OAI21X1  g03136(.A0(new_n5562_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n5573_));
  AOI21X1  g03137(.A0(new_n5572_), .A1(new_n5565_), .B0(new_n5573_), .Y(new_n5574_));
  AOI22X1  g03138(.A0(new_n5569_), .A1(new_n3074_), .B0(new_n5561_), .B1(new_n3087_), .Y(new_n5575_));
  AND2X1   g03139(.A(new_n5575_), .B(pi0075), .Y(new_n5576_));
  OR2X1    g03140(.A(new_n5576_), .B(pi0092), .Y(new_n5577_));
  NAND2X1  g03141(.A(new_n5575_), .B(new_n3073_), .Y(new_n5578_));
  AOI21X1  g03142(.A0(new_n5562_), .A1(pi0075), .B0(new_n3079_), .Y(new_n5579_));
  AOI21X1  g03143(.A0(new_n5579_), .A1(new_n5578_), .B0(pi0054), .Y(new_n5580_));
  OAI21X1  g03144(.A0(new_n5577_), .A1(new_n5574_), .B0(new_n5580_), .Y(new_n5581_));
  MX2X1    g03145(.A(new_n5575_), .B(new_n5562_), .S0(new_n5295_), .Y(new_n5582_));
  AOI21X1  g03146(.A0(new_n5582_), .A1(pi0054), .B0(pi0074), .Y(new_n5583_));
  AND3X1   g03147(.A(new_n5575_), .B(new_n3084_), .C(new_n3091_), .Y(new_n5584_));
  OAI21X1  g03148(.A0(new_n5569_), .A1(new_n5299_), .B0(pi0074), .Y(new_n5585_));
  OAI21X1  g03149(.A0(new_n5585_), .A1(new_n5584_), .B0(new_n3107_), .Y(new_n5586_));
  AOI21X1  g03150(.A0(new_n5583_), .A1(new_n5581_), .B0(new_n5586_), .Y(new_n5587_));
  AND3X1   g03151(.A(new_n5538_), .B(new_n5037_), .C(new_n3104_), .Y(new_n5588_));
  OR2X1    g03152(.A(new_n5545_), .B(new_n3107_), .Y(new_n5589_));
  OAI21X1  g03153(.A0(new_n5589_), .A1(new_n5588_), .B0(new_n3123_), .Y(new_n5590_));
  AOI21X1  g03154(.A0(new_n5545_), .A1(new_n4975_), .B0(pi0059), .Y(new_n5591_));
  OAI21X1  g03155(.A0(new_n5590_), .A1(new_n5587_), .B0(new_n5591_), .Y(new_n5592_));
  NAND4X1  g03156(.A(new_n5538_), .B(new_n5306_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5593_));
  AOI21X1  g03157(.A0(new_n5394_), .A1(pi0960), .B0(new_n3127_), .Y(new_n5594_));
  AOI21X1  g03158(.A0(new_n5594_), .A1(new_n5593_), .B0(pi0057), .Y(new_n5595_));
  AOI22X1  g03159(.A0(new_n5595_), .A1(new_n5592_), .B0(new_n5540_), .B1(pi0057), .Y(po0175));
  INVX1    g03160(.A(pi0963), .Y(new_n5597_));
  AND2X1   g03161(.A(pi0963), .B(new_n2793_), .Y(new_n5598_));
  NAND4X1  g03162(.A(new_n5598_), .B(new_n5102_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5599_));
  OAI21X1  g03163(.A0(new_n5395_), .A1(new_n5597_), .B0(new_n5599_), .Y(new_n5600_));
  AOI21X1  g03164(.A0(new_n5394_), .A1(pi0963), .B0(new_n2933_), .Y(new_n5601_));
  INVX1    g03165(.A(new_n5601_), .Y(new_n5602_));
  AOI21X1  g03166(.A0(new_n5598_), .A1(new_n5401_), .B0(new_n5602_), .Y(new_n5603_));
  AOI21X1  g03167(.A0(new_n5113_), .A1(pi0299), .B0(new_n5603_), .Y(new_n5604_));
  AND2X1   g03168(.A(new_n5394_), .B(pi0963), .Y(new_n5605_));
  AND3X1   g03169(.A(new_n5598_), .B(new_n5406_), .C(new_n5023_), .Y(new_n5606_));
  OR2X1    g03170(.A(new_n5606_), .B(new_n5605_), .Y(new_n5607_));
  AOI21X1  g03171(.A0(new_n5607_), .A1(new_n5113_), .B0(new_n5604_), .Y(new_n5608_));
  AOI21X1  g03172(.A0(new_n5414_), .A1(pi0969), .B0(pi0299), .Y(new_n5609_));
  OR2X1    g03173(.A(new_n5609_), .B(new_n5215_), .Y(new_n5610_));
  AOI21X1  g03174(.A0(new_n5417_), .A1(pi0969), .B0(pi0299), .Y(new_n5611_));
  OR3X1    g03175(.A(new_n5611_), .B(new_n5603_), .C(pi0232), .Y(new_n5612_));
  OAI21X1  g03176(.A0(new_n5610_), .A1(new_n5608_), .B0(new_n5612_), .Y(new_n5613_));
  AND2X1   g03177(.A(pi0969), .B(new_n2933_), .Y(new_n5614_));
  AND2X1   g03178(.A(pi0963), .B(pi0299), .Y(new_n5615_));
  AOI22X1  g03179(.A0(new_n5615_), .A1(new_n5423_), .B0(new_n5614_), .B1(new_n5425_), .Y(new_n5616_));
  OAI21X1  g03180(.A0(new_n5616_), .A1(new_n5428_), .B0(new_n2979_), .Y(new_n5617_));
  AOI21X1  g03181(.A0(new_n5613_), .A1(new_n2939_), .B0(new_n5617_), .Y(new_n5618_));
  AOI21X1  g03182(.A0(new_n5432_), .A1(pi0969), .B0(pi0299), .Y(new_n5619_));
  AOI21X1  g03183(.A0(new_n5598_), .A1(new_n5037_), .B0(new_n5602_), .Y(new_n5620_));
  NOR3X1   g03184(.A(new_n5620_), .B(new_n5619_), .C(pi0039), .Y(new_n5621_));
  OAI21X1  g03185(.A0(new_n5615_), .A1(new_n5614_), .B0(new_n5394_), .Y(new_n5622_));
  OAI21X1  g03186(.A0(new_n5622_), .A1(new_n2939_), .B0(pi0038), .Y(new_n5623_));
  NOR2X1   g03187(.A(new_n5623_), .B(new_n5621_), .Y(new_n5624_));
  OAI21X1  g03188(.A0(new_n5624_), .A1(new_n5618_), .B0(new_n3007_), .Y(new_n5625_));
  AOI21X1  g03189(.A0(new_n5443_), .A1(pi0969), .B0(pi0299), .Y(new_n5626_));
  NOR4X1   g03190(.A(new_n5446_), .B(new_n5445_), .C(new_n5597_), .D(pi0228), .Y(new_n5627_));
  OAI21X1  g03191(.A0(new_n5627_), .A1(new_n5602_), .B0(new_n3047_), .Y(new_n5628_));
  INVX1    g03192(.A(new_n5622_), .Y(new_n5629_));
  AOI21X1  g03193(.A0(new_n5629_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n5630_));
  OAI21X1  g03194(.A0(new_n5628_), .A1(new_n5626_), .B0(new_n5630_), .Y(new_n5631_));
  AND2X1   g03195(.A(new_n5631_), .B(new_n3131_), .Y(new_n5632_));
  OAI21X1  g03196(.A0(new_n5622_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n5633_));
  AOI21X1  g03197(.A0(new_n5632_), .A1(new_n5625_), .B0(new_n5633_), .Y(new_n5634_));
  AOI22X1  g03198(.A0(new_n5629_), .A1(new_n3074_), .B0(new_n5621_), .B1(new_n3087_), .Y(new_n5635_));
  AND2X1   g03199(.A(new_n5635_), .B(pi0075), .Y(new_n5636_));
  OR2X1    g03200(.A(new_n5636_), .B(pi0092), .Y(new_n5637_));
  NAND2X1  g03201(.A(new_n5635_), .B(new_n3073_), .Y(new_n5638_));
  AOI21X1  g03202(.A0(new_n5622_), .A1(pi0075), .B0(new_n3079_), .Y(new_n5639_));
  AOI21X1  g03203(.A0(new_n5639_), .A1(new_n5638_), .B0(pi0054), .Y(new_n5640_));
  OAI21X1  g03204(.A0(new_n5637_), .A1(new_n5634_), .B0(new_n5640_), .Y(new_n5641_));
  MX2X1    g03205(.A(new_n5635_), .B(new_n5622_), .S0(new_n5295_), .Y(new_n5642_));
  AOI21X1  g03206(.A0(new_n5642_), .A1(pi0054), .B0(pi0074), .Y(new_n5643_));
  AND3X1   g03207(.A(new_n5635_), .B(new_n3084_), .C(new_n3091_), .Y(new_n5644_));
  OAI21X1  g03208(.A0(new_n5629_), .A1(new_n5299_), .B0(pi0074), .Y(new_n5645_));
  OAI21X1  g03209(.A0(new_n5645_), .A1(new_n5644_), .B0(new_n3107_), .Y(new_n5646_));
  AOI21X1  g03210(.A0(new_n5643_), .A1(new_n5641_), .B0(new_n5646_), .Y(new_n5647_));
  AND3X1   g03211(.A(new_n5598_), .B(new_n5037_), .C(new_n3104_), .Y(new_n5648_));
  OR2X1    g03212(.A(new_n5605_), .B(new_n3107_), .Y(new_n5649_));
  OAI21X1  g03213(.A0(new_n5649_), .A1(new_n5648_), .B0(new_n3123_), .Y(new_n5650_));
  AOI21X1  g03214(.A0(new_n5605_), .A1(new_n4975_), .B0(pi0059), .Y(new_n5651_));
  OAI21X1  g03215(.A0(new_n5650_), .A1(new_n5647_), .B0(new_n5651_), .Y(new_n5652_));
  NAND4X1  g03216(.A(new_n5598_), .B(new_n5306_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5653_));
  AOI21X1  g03217(.A0(new_n5394_), .A1(pi0963), .B0(new_n3127_), .Y(new_n5654_));
  AOI21X1  g03218(.A0(new_n5654_), .A1(new_n5653_), .B0(pi0057), .Y(new_n5655_));
  AOI22X1  g03219(.A0(new_n5655_), .A1(new_n5652_), .B0(new_n5600_), .B1(pi0057), .Y(po0176));
  INVX1    g03220(.A(pi0975), .Y(new_n5657_));
  AND2X1   g03221(.A(pi0975), .B(new_n2793_), .Y(new_n5658_));
  NAND4X1  g03222(.A(new_n5658_), .B(new_n5102_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5659_));
  OAI21X1  g03223(.A0(new_n5395_), .A1(new_n5657_), .B0(new_n5659_), .Y(new_n5660_));
  AOI21X1  g03224(.A0(new_n5394_), .A1(pi0975), .B0(new_n2933_), .Y(new_n5661_));
  INVX1    g03225(.A(new_n5661_), .Y(new_n5662_));
  AOI21X1  g03226(.A0(new_n5658_), .A1(new_n5401_), .B0(new_n5662_), .Y(new_n5663_));
  AOI21X1  g03227(.A0(new_n5113_), .A1(pi0299), .B0(new_n5663_), .Y(new_n5664_));
  AND2X1   g03228(.A(new_n5394_), .B(pi0975), .Y(new_n5665_));
  AND3X1   g03229(.A(new_n5658_), .B(new_n5406_), .C(new_n5023_), .Y(new_n5666_));
  OR2X1    g03230(.A(new_n5666_), .B(new_n5665_), .Y(new_n5667_));
  AOI21X1  g03231(.A0(new_n5667_), .A1(new_n5113_), .B0(new_n5664_), .Y(new_n5668_));
  AOI21X1  g03232(.A0(new_n5414_), .A1(pi0971), .B0(pi0299), .Y(new_n5669_));
  OR2X1    g03233(.A(new_n5669_), .B(new_n5215_), .Y(new_n5670_));
  AOI21X1  g03234(.A0(new_n5417_), .A1(pi0971), .B0(pi0299), .Y(new_n5671_));
  OR3X1    g03235(.A(new_n5671_), .B(new_n5663_), .C(pi0232), .Y(new_n5672_));
  OAI21X1  g03236(.A0(new_n5670_), .A1(new_n5668_), .B0(new_n5672_), .Y(new_n5673_));
  AND2X1   g03237(.A(pi0971), .B(new_n2933_), .Y(new_n5674_));
  AND2X1   g03238(.A(pi0975), .B(pi0299), .Y(new_n5675_));
  AOI22X1  g03239(.A0(new_n5675_), .A1(new_n5423_), .B0(new_n5674_), .B1(new_n5425_), .Y(new_n5676_));
  OAI21X1  g03240(.A0(new_n5676_), .A1(new_n5428_), .B0(new_n2979_), .Y(new_n5677_));
  AOI21X1  g03241(.A0(new_n5673_), .A1(new_n2939_), .B0(new_n5677_), .Y(new_n5678_));
  AOI21X1  g03242(.A0(new_n5432_), .A1(pi0971), .B0(pi0299), .Y(new_n5679_));
  AOI21X1  g03243(.A0(new_n5658_), .A1(new_n5037_), .B0(new_n5662_), .Y(new_n5680_));
  NOR3X1   g03244(.A(new_n5680_), .B(new_n5679_), .C(pi0039), .Y(new_n5681_));
  OAI21X1  g03245(.A0(new_n5675_), .A1(new_n5674_), .B0(new_n5394_), .Y(new_n5682_));
  OAI21X1  g03246(.A0(new_n5682_), .A1(new_n2939_), .B0(pi0038), .Y(new_n5683_));
  NOR2X1   g03247(.A(new_n5683_), .B(new_n5681_), .Y(new_n5684_));
  OAI21X1  g03248(.A0(new_n5684_), .A1(new_n5678_), .B0(new_n3007_), .Y(new_n5685_));
  AOI21X1  g03249(.A0(new_n5443_), .A1(pi0971), .B0(pi0299), .Y(new_n5686_));
  NOR4X1   g03250(.A(new_n5446_), .B(new_n5445_), .C(new_n5657_), .D(pi0228), .Y(new_n5687_));
  OAI21X1  g03251(.A0(new_n5687_), .A1(new_n5662_), .B0(new_n3047_), .Y(new_n5688_));
  INVX1    g03252(.A(new_n5682_), .Y(new_n5689_));
  AOI21X1  g03253(.A0(new_n5689_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n5690_));
  OAI21X1  g03254(.A0(new_n5688_), .A1(new_n5686_), .B0(new_n5690_), .Y(new_n5691_));
  AND2X1   g03255(.A(new_n5691_), .B(new_n3131_), .Y(new_n5692_));
  OAI21X1  g03256(.A0(new_n5682_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n5693_));
  AOI21X1  g03257(.A0(new_n5692_), .A1(new_n5685_), .B0(new_n5693_), .Y(new_n5694_));
  AOI22X1  g03258(.A0(new_n5689_), .A1(new_n3074_), .B0(new_n5681_), .B1(new_n3087_), .Y(new_n5695_));
  AND2X1   g03259(.A(new_n5695_), .B(pi0075), .Y(new_n5696_));
  OR2X1    g03260(.A(new_n5696_), .B(pi0092), .Y(new_n5697_));
  NAND2X1  g03261(.A(new_n5695_), .B(new_n3073_), .Y(new_n5698_));
  AOI21X1  g03262(.A0(new_n5682_), .A1(pi0075), .B0(new_n3079_), .Y(new_n5699_));
  AOI21X1  g03263(.A0(new_n5699_), .A1(new_n5698_), .B0(pi0054), .Y(new_n5700_));
  OAI21X1  g03264(.A0(new_n5697_), .A1(new_n5694_), .B0(new_n5700_), .Y(new_n5701_));
  MX2X1    g03265(.A(new_n5695_), .B(new_n5682_), .S0(new_n5295_), .Y(new_n5702_));
  AOI21X1  g03266(.A0(new_n5702_), .A1(pi0054), .B0(pi0074), .Y(new_n5703_));
  AND3X1   g03267(.A(new_n5695_), .B(new_n3084_), .C(new_n3091_), .Y(new_n5704_));
  OAI21X1  g03268(.A0(new_n5689_), .A1(new_n5299_), .B0(pi0074), .Y(new_n5705_));
  OAI21X1  g03269(.A0(new_n5705_), .A1(new_n5704_), .B0(new_n3107_), .Y(new_n5706_));
  AOI21X1  g03270(.A0(new_n5703_), .A1(new_n5701_), .B0(new_n5706_), .Y(new_n5707_));
  AND3X1   g03271(.A(new_n5658_), .B(new_n5037_), .C(new_n3104_), .Y(new_n5708_));
  OR2X1    g03272(.A(new_n5665_), .B(new_n3107_), .Y(new_n5709_));
  OAI21X1  g03273(.A0(new_n5709_), .A1(new_n5708_), .B0(new_n3123_), .Y(new_n5710_));
  AOI21X1  g03274(.A0(new_n5665_), .A1(new_n4975_), .B0(pi0059), .Y(new_n5711_));
  OAI21X1  g03275(.A0(new_n5710_), .A1(new_n5707_), .B0(new_n5711_), .Y(new_n5712_));
  NAND4X1  g03276(.A(new_n5658_), .B(new_n5306_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5713_));
  AOI21X1  g03277(.A0(new_n5394_), .A1(pi0975), .B0(new_n3127_), .Y(new_n5714_));
  AOI21X1  g03278(.A0(new_n5714_), .A1(new_n5713_), .B0(pi0057), .Y(new_n5715_));
  AOI22X1  g03279(.A0(new_n5715_), .A1(new_n5712_), .B0(new_n5660_), .B1(pi0057), .Y(po0177));
  INVX1    g03280(.A(pi0978), .Y(new_n5717_));
  AND2X1   g03281(.A(pi0978), .B(new_n2793_), .Y(new_n5718_));
  NAND4X1  g03282(.A(new_n5718_), .B(new_n5102_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5719_));
  OAI21X1  g03283(.A0(new_n5395_), .A1(new_n5717_), .B0(new_n5719_), .Y(new_n5720_));
  AND2X1   g03284(.A(pi0978), .B(pi0299), .Y(new_n5721_));
  AOI21X1  g03285(.A0(pi0974), .A1(new_n2933_), .B0(new_n5721_), .Y(new_n5722_));
  INVX1    g03286(.A(new_n5722_), .Y(new_n5723_));
  AND2X1   g03287(.A(new_n5723_), .B(new_n5432_), .Y(new_n5724_));
  AND2X1   g03288(.A(new_n5723_), .B(new_n5394_), .Y(new_n5725_));
  INVX1    g03289(.A(new_n5725_), .Y(new_n5726_));
  OAI21X1  g03290(.A0(new_n5726_), .A1(new_n2939_), .B0(pi0038), .Y(new_n5727_));
  AOI21X1  g03291(.A0(new_n5724_), .A1(new_n2939_), .B0(new_n5727_), .Y(new_n5728_));
  AOI21X1  g03292(.A0(new_n5394_), .A1(pi0978), .B0(new_n2933_), .Y(new_n5729_));
  INVX1    g03293(.A(new_n5729_), .Y(new_n5730_));
  AOI21X1  g03294(.A0(new_n5718_), .A1(new_n5401_), .B0(new_n5730_), .Y(new_n5731_));
  AOI21X1  g03295(.A0(new_n5113_), .A1(pi0299), .B0(new_n5731_), .Y(new_n5732_));
  AND2X1   g03296(.A(new_n5394_), .B(pi0978), .Y(new_n5733_));
  AND3X1   g03297(.A(new_n5718_), .B(new_n5406_), .C(new_n5023_), .Y(new_n5734_));
  OR2X1    g03298(.A(new_n5734_), .B(new_n5733_), .Y(new_n5735_));
  AOI21X1  g03299(.A0(new_n5735_), .A1(new_n5113_), .B0(new_n5732_), .Y(new_n5736_));
  AOI21X1  g03300(.A0(new_n5414_), .A1(pi0974), .B0(pi0299), .Y(new_n5737_));
  OR2X1    g03301(.A(new_n5737_), .B(new_n5215_), .Y(new_n5738_));
  AOI21X1  g03302(.A0(new_n5417_), .A1(pi0974), .B0(pi0299), .Y(new_n5739_));
  OR3X1    g03303(.A(new_n5739_), .B(new_n5731_), .C(pi0232), .Y(new_n5740_));
  OAI21X1  g03304(.A0(new_n5738_), .A1(new_n5736_), .B0(new_n5740_), .Y(new_n5741_));
  AND2X1   g03305(.A(pi0974), .B(new_n2933_), .Y(new_n5742_));
  AOI22X1  g03306(.A0(new_n5721_), .A1(new_n5423_), .B0(new_n5742_), .B1(new_n5425_), .Y(new_n5743_));
  OAI21X1  g03307(.A0(new_n5743_), .A1(new_n5428_), .B0(new_n2979_), .Y(new_n5744_));
  AOI21X1  g03308(.A0(new_n5741_), .A1(new_n2939_), .B0(new_n5744_), .Y(new_n5745_));
  OAI21X1  g03309(.A0(new_n5745_), .A1(new_n5728_), .B0(new_n3007_), .Y(new_n5746_));
  AOI21X1  g03310(.A0(new_n5443_), .A1(pi0974), .B0(pi0299), .Y(new_n5747_));
  NOR4X1   g03311(.A(new_n5446_), .B(new_n5445_), .C(new_n5717_), .D(pi0228), .Y(new_n5748_));
  OAI21X1  g03312(.A0(new_n5748_), .A1(new_n5730_), .B0(new_n3047_), .Y(new_n5749_));
  AOI21X1  g03313(.A0(new_n5725_), .A1(new_n3060_), .B0(new_n3007_), .Y(new_n5750_));
  OAI21X1  g03314(.A0(new_n5749_), .A1(new_n5747_), .B0(new_n5750_), .Y(new_n5751_));
  AND2X1   g03315(.A(new_n5751_), .B(new_n3131_), .Y(new_n5752_));
  OAI21X1  g03316(.A0(new_n5726_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n5753_));
  AOI21X1  g03317(.A0(new_n5752_), .A1(new_n5746_), .B0(new_n5753_), .Y(new_n5754_));
  OAI21X1  g03318(.A0(new_n3070_), .A1(pi0228), .B0(new_n5724_), .Y(new_n5755_));
  AND2X1   g03319(.A(new_n5755_), .B(pi0075), .Y(new_n5756_));
  OR2X1    g03320(.A(new_n5756_), .B(pi0092), .Y(new_n5757_));
  OAI21X1  g03321(.A0(new_n5725_), .A1(new_n3073_), .B0(pi0092), .Y(new_n5758_));
  AOI21X1  g03322(.A0(new_n5755_), .A1(new_n3073_), .B0(new_n5758_), .Y(new_n5759_));
  NOR2X1   g03323(.A(new_n5759_), .B(pi0054), .Y(new_n5760_));
  OAI21X1  g03324(.A0(new_n5757_), .A1(new_n5754_), .B0(new_n5760_), .Y(new_n5761_));
  MX2X1    g03325(.A(new_n5755_), .B(new_n5726_), .S0(new_n5295_), .Y(new_n5762_));
  AOI21X1  g03326(.A0(new_n5762_), .A1(pi0054), .B0(pi0074), .Y(new_n5763_));
  AND3X1   g03327(.A(new_n5755_), .B(new_n3084_), .C(new_n3091_), .Y(new_n5764_));
  OAI21X1  g03328(.A0(new_n5725_), .A1(new_n5299_), .B0(pi0074), .Y(new_n5765_));
  OAI21X1  g03329(.A0(new_n5765_), .A1(new_n5764_), .B0(new_n3107_), .Y(new_n5766_));
  AOI21X1  g03330(.A0(new_n5763_), .A1(new_n5761_), .B0(new_n5766_), .Y(new_n5767_));
  AND3X1   g03331(.A(new_n5718_), .B(new_n5037_), .C(new_n3104_), .Y(new_n5768_));
  OR2X1    g03332(.A(new_n5733_), .B(new_n3107_), .Y(new_n5769_));
  OAI21X1  g03333(.A0(new_n5769_), .A1(new_n5768_), .B0(new_n3123_), .Y(new_n5770_));
  AOI21X1  g03334(.A0(new_n5733_), .A1(new_n4975_), .B0(pi0059), .Y(new_n5771_));
  OAI21X1  g03335(.A0(new_n5770_), .A1(new_n5767_), .B0(new_n5771_), .Y(new_n5772_));
  NAND4X1  g03336(.A(new_n5718_), .B(new_n5306_), .C(new_n5037_), .D(new_n3104_), .Y(new_n5773_));
  AOI21X1  g03337(.A0(new_n5394_), .A1(pi0978), .B0(new_n3127_), .Y(new_n5774_));
  AOI21X1  g03338(.A0(new_n5774_), .A1(new_n5773_), .B0(pi0057), .Y(new_n5775_));
  AOI22X1  g03339(.A0(new_n5775_), .A1(new_n5772_), .B0(new_n5720_), .B1(pi0057), .Y(po0178));
  INVX1    g03340(.A(pi0024), .Y(new_n5777_));
  INVX1    g03341(.A(new_n3087_), .Y(new_n5778_));
  NOR4X1   g03342(.A(new_n5778_), .B(new_n2985_), .C(new_n2536_), .D(pi0039), .Y(new_n5779_));
  NOR2X1   g03343(.A(new_n5779_), .B(new_n3073_), .Y(new_n5780_));
  INVX1    g03344(.A(new_n5780_), .Y(new_n5781_));
  NOR3X1   g03345(.A(new_n2985_), .B(new_n2536_), .C(pi0039), .Y(new_n5782_));
  AND3X1   g03346(.A(new_n5782_), .B(new_n3077_), .C(new_n3251_), .Y(new_n5783_));
  OR2X1    g03347(.A(new_n5783_), .B(new_n3079_), .Y(new_n5784_));
  AND2X1   g03348(.A(new_n5784_), .B(new_n5781_), .Y(new_n5785_));
  NOR4X1   g03349(.A(new_n5242_), .B(new_n5221_), .C(new_n5062_), .D(new_n2933_), .Y(new_n5786_));
  OR2X1    g03350(.A(new_n5049_), .B(pi0299), .Y(new_n5787_));
  OAI21X1  g03351(.A0(new_n5787_), .A1(new_n5250_), .B0(pi0039), .Y(new_n5788_));
  NAND3X1  g03352(.A(new_n5210_), .B(new_n5206_), .C(new_n5023_), .Y(new_n5789_));
  AOI21X1  g03353(.A0(new_n5199_), .A1(new_n5048_), .B0(pi0299), .Y(new_n5790_));
  AND3X1   g03354(.A(new_n5790_), .B(new_n5789_), .C(new_n5412_), .Y(new_n5791_));
  OAI21X1  g03355(.A0(new_n5175_), .A1(new_n5171_), .B0(new_n5048_), .Y(new_n5792_));
  NAND3X1  g03356(.A(new_n5792_), .B(new_n5113_), .C(pi0299), .Y(new_n5793_));
  OR4X1    g03357(.A(new_n5175_), .B(new_n5171_), .C(new_n5113_), .D(new_n2933_), .Y(new_n5794_));
  AND2X1   g03358(.A(new_n5794_), .B(pi0232), .Y(new_n5795_));
  OAI21X1  g03359(.A0(new_n5793_), .A1(new_n5406_), .B0(new_n5795_), .Y(new_n5796_));
  OR3X1    g03360(.A(new_n5198_), .B(new_n5171_), .C(pi0299), .Y(new_n5797_));
  NOR3X1   g03361(.A(new_n5175_), .B(new_n5171_), .C(new_n2933_), .Y(new_n5798_));
  NOR2X1   g03362(.A(new_n5798_), .B(pi0232), .Y(new_n5799_));
  AOI21X1  g03363(.A0(new_n5799_), .A1(new_n5797_), .B0(pi0039), .Y(new_n5800_));
  OAI21X1  g03364(.A0(new_n5796_), .A1(new_n5791_), .B0(new_n5800_), .Y(new_n5801_));
  OAI21X1  g03365(.A0(new_n5788_), .A1(new_n5786_), .B0(new_n5801_), .Y(new_n5802_));
  MX2X1    g03366(.A(new_n5802_), .B(new_n4987_), .S0(pi0038), .Y(new_n5803_));
  NOR4X1   g03367(.A(new_n2985_), .B(new_n2536_), .C(pi0039), .D(pi0038), .Y(new_n5804_));
  NOR2X1   g03368(.A(new_n5804_), .B(new_n3007_), .Y(new_n5805_));
  OR2X1    g03369(.A(new_n5805_), .B(new_n5089_), .Y(new_n5806_));
  AOI21X1  g03370(.A0(new_n5803_), .A1(new_n3007_), .B0(new_n5806_), .Y(new_n5807_));
  OAI21X1  g03371(.A0(new_n5807_), .A1(new_n5295_), .B0(new_n5785_), .Y(new_n5808_));
  AND2X1   g03372(.A(new_n5783_), .B(new_n3079_), .Y(new_n5809_));
  INVX1    g03373(.A(new_n5809_), .Y(new_n5810_));
  MX2X1    g03374(.A(new_n5810_), .B(new_n5808_), .S0(new_n3091_), .Y(new_n5811_));
  AOI21X1  g03375(.A0(new_n5811_), .A1(new_n4982_), .B0(new_n4984_), .Y(new_n5812_));
  AND3X1   g03376(.A(new_n3102_), .B(new_n3077_), .C(new_n3079_), .Y(new_n5813_));
  AOI21X1  g03377(.A0(new_n4979_), .A1(new_n5813_), .B0(new_n3107_), .Y(new_n5814_));
  NOR3X1   g03378(.A(new_n5814_), .B(pi0062), .C(pi0056), .Y(new_n5815_));
  OAI21X1  g03379(.A0(new_n5812_), .A1(pi0055), .B0(new_n5815_), .Y(new_n5816_));
  AOI21X1  g03380(.A0(new_n5816_), .A1(new_n3223_), .B0(new_n4977_), .Y(po0195));
  MX2X1    g03381(.A(po0195), .B(new_n5777_), .S0(pi0954), .Y(po0182));
  NOR4X1   g03382(.A(new_n3378_), .B(new_n2985_), .C(new_n2536_), .D(pi0228), .Y(new_n5819_));
  AND2X1   g03383(.A(new_n5819_), .B(new_n5096_), .Y(new_n5820_));
  OAI21X1  g03384(.A0(new_n5820_), .A1(new_n3009_), .B0(pi0062), .Y(new_n5821_));
  OR3X1    g03385(.A(new_n3180_), .B(pi0228), .C(pi0100), .Y(new_n5822_));
  NOR3X1   g03386(.A(new_n5267_), .B(new_n2985_), .C(new_n2536_), .Y(new_n5823_));
  MX2X1    g03387(.A(new_n5823_), .B(new_n3198_), .S0(pi0299), .Y(new_n5824_));
  NAND3X1  g03388(.A(new_n5824_), .B(new_n3603_), .C(pi0100), .Y(new_n5825_));
  AND3X1   g03389(.A(new_n5825_), .B(new_n5822_), .C(new_n2939_), .Y(new_n5826_));
  NOR4X1   g03390(.A(new_n2985_), .B(new_n2536_), .C(pi0228), .D(pi0100), .Y(new_n5827_));
  OAI21X1  g03391(.A0(new_n5827_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n5828_));
  OAI21X1  g03392(.A0(new_n5828_), .A1(new_n5826_), .B0(new_n3011_), .Y(new_n5829_));
  OAI21X1  g03393(.A0(new_n5819_), .A1(new_n3009_), .B0(pi0087), .Y(new_n5830_));
  NAND2X1  g03394(.A(new_n5830_), .B(new_n3073_), .Y(new_n5831_));
  AOI21X1  g03395(.A0(new_n5829_), .A1(new_n3131_), .B0(new_n5831_), .Y(new_n5832_));
  OAI21X1  g03396(.A0(new_n3009_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n5833_));
  NOR4X1   g03397(.A(new_n3279_), .B(new_n2985_), .C(new_n2536_), .D(pi0228), .Y(new_n5834_));
  OAI21X1  g03398(.A0(new_n5834_), .A1(new_n3009_), .B0(pi0092), .Y(new_n5835_));
  AND2X1   g03399(.A(new_n5835_), .B(new_n3102_), .Y(new_n5836_));
  OAI21X1  g03400(.A0(new_n5833_), .A1(new_n5832_), .B0(new_n5836_), .Y(new_n5837_));
  AOI21X1  g03401(.A0(new_n3130_), .A1(new_n3011_), .B0(pi0055), .Y(new_n5838_));
  AND2X1   g03402(.A(new_n4983_), .B(new_n3111_), .Y(new_n5839_));
  INVX1    g03403(.A(new_n5839_), .Y(new_n5840_));
  NOR4X1   g03404(.A(new_n5840_), .B(new_n2985_), .C(new_n2536_), .D(pi0228), .Y(new_n5841_));
  AOI21X1  g03405(.A0(new_n5841_), .A1(new_n4982_), .B0(new_n3009_), .Y(new_n5842_));
  OAI21X1  g03406(.A0(new_n5842_), .A1(new_n3107_), .B0(new_n3118_), .Y(new_n5843_));
  AOI21X1  g03407(.A0(new_n5838_), .A1(new_n5837_), .B0(new_n5843_), .Y(new_n5844_));
  NOR4X1   g03408(.A(new_n3115_), .B(new_n2985_), .C(new_n2536_), .D(pi0228), .Y(new_n5845_));
  OR2X1    g03409(.A(new_n3009_), .B(new_n3118_), .Y(new_n5846_));
  OAI21X1  g03410(.A0(new_n5846_), .A1(new_n5845_), .B0(new_n3222_), .Y(new_n5847_));
  OAI21X1  g03411(.A0(new_n5847_), .A1(new_n5844_), .B0(new_n5821_), .Y(new_n5848_));
  MX2X1    g03412(.A(new_n5848_), .B(new_n3009_), .S0(new_n3374_), .Y(po0183));
  AND2X1   g03413(.A(pi1056), .B(pi0119), .Y(new_n5850_));
  AOI21X1  g03414(.A0(pi0252), .A1(new_n2793_), .B0(pi0119), .Y(new_n5851_));
  OR3X1    g03415(.A(new_n5851_), .B(new_n5850_), .C(pi0468), .Y(po0184));
  AND2X1   g03416(.A(pi1077), .B(pi0119), .Y(new_n5853_));
  OR3X1    g03417(.A(new_n5853_), .B(new_n5851_), .C(pi0468), .Y(po0185));
  AND2X1   g03418(.A(pi1073), .B(pi0119), .Y(new_n5855_));
  OR3X1    g03419(.A(new_n5855_), .B(new_n5851_), .C(pi0468), .Y(po0186));
  AND2X1   g03420(.A(pi1041), .B(pi0119), .Y(new_n5857_));
  OR3X1    g03421(.A(new_n5857_), .B(new_n5851_), .C(pi0468), .Y(po0187));
  XOR2X1   g03422(.A(pi0462), .B(pi0360), .Y(new_n5859_));
  INVX1    g03423(.A(pi0352), .Y(new_n5860_));
  XOR2X1   g03424(.A(pi0353), .B(new_n5860_), .Y(new_n5861_));
  XOR2X1   g03425(.A(new_n5861_), .B(new_n5859_), .Y(new_n5862_));
  XOR2X1   g03426(.A(new_n5862_), .B(pi0354), .Y(new_n5863_));
  INVX1    g03427(.A(pi0356), .Y(new_n5864_));
  INVX1    g03428(.A(pi0357), .Y(new_n5865_));
  INVX1    g03429(.A(pi0461), .Y(new_n5866_));
  XOR2X1   g03430(.A(pi0346), .B(pi0345), .Y(new_n5867_));
  XOR2X1   g03431(.A(new_n5867_), .B(pi0323), .Y(new_n5868_));
  INVX1    g03432(.A(pi0358), .Y(new_n5869_));
  XOR2X1   g03433(.A(pi0450), .B(new_n5869_), .Y(new_n5870_));
  XOR2X1   g03434(.A(new_n5870_), .B(new_n5868_), .Y(new_n5871_));
  XOR2X1   g03435(.A(pi0362), .B(pi0327), .Y(new_n5872_));
  XOR2X1   g03436(.A(pi0344), .B(pi0343), .Y(new_n5873_));
  XOR2X1   g03437(.A(new_n5873_), .B(new_n5872_), .Y(new_n5874_));
  INVX1    g03438(.A(new_n5874_), .Y(new_n5875_));
  INVX1    g03439(.A(pi1197), .Y(new_n5876_));
  AOI21X1  g03440(.A0(new_n5875_), .A1(new_n5871_), .B0(new_n5876_), .Y(new_n5877_));
  OAI21X1  g03441(.A0(new_n5875_), .A1(new_n5871_), .B0(new_n5877_), .Y(new_n5878_));
  INVX1    g03442(.A(new_n5878_), .Y(new_n5879_));
  NOR3X1   g03443(.A(pi0092), .B(pi0074), .C(pi0054), .Y(new_n5880_));
  INVX1    g03444(.A(new_n2984_), .Y(new_n5881_));
  NOR3X1   g03445(.A(new_n5031_), .B(new_n5024_), .C(new_n5084_), .Y(new_n5882_));
  INVX1    g03446(.A(new_n5882_), .Y(new_n5883_));
  INVX1    g03447(.A(new_n2847_), .Y(new_n5884_));
  AND3X1   g03448(.A(new_n5003_), .B(new_n2535_), .C(new_n2508_), .Y(new_n5885_));
  AND3X1   g03449(.A(new_n2477_), .B(new_n2705_), .C(pi0090), .Y(new_n5886_));
  NOR2X1   g03450(.A(new_n5886_), .B(pi0093), .Y(new_n5887_));
  INVX1    g03451(.A(new_n5887_), .Y(new_n5888_));
  AOI21X1  g03452(.A0(new_n5888_), .A1(new_n5885_), .B0(pi0051), .Y(new_n5889_));
  INVX1    g03453(.A(new_n5889_), .Y(new_n5890_));
  NOR2X1   g03454(.A(pi0077), .B(pi0050), .Y(new_n5891_));
  INVX1    g03455(.A(new_n5891_), .Y(new_n5892_));
  INVX1    g03456(.A(pi0098), .Y(new_n5893_));
  OR3X1    g03457(.A(new_n2472_), .B(new_n5893_), .C(pi0088), .Y(new_n5894_));
  NOR4X1   g03458(.A(new_n5894_), .B(new_n5892_), .C(new_n2567_), .D(pi0094), .Y(new_n5895_));
  NOR2X1   g03459(.A(new_n5895_), .B(pi0097), .Y(new_n5896_));
  NOR3X1   g03460(.A(pi0093), .B(pi0090), .C(pi0035), .Y(new_n5897_));
  INVX1    g03461(.A(new_n5897_), .Y(new_n5898_));
  NOR4X1   g03462(.A(new_n5898_), .B(new_n5896_), .C(new_n2498_), .D(pi0070), .Y(new_n5899_));
  OAI21X1  g03463(.A0(new_n5899_), .A1(new_n5890_), .B0(new_n5884_), .Y(new_n5900_));
  NOR4X1   g03464(.A(new_n5900_), .B(new_n5883_), .C(new_n5881_), .D(pi0096), .Y(new_n5901_));
  OAI21X1  g03465(.A0(new_n5237_), .A1(pi0122), .B0(new_n5901_), .Y(new_n5902_));
  AND2X1   g03466(.A(new_n5900_), .B(new_n2513_), .Y(new_n5903_));
  OR2X1    g03467(.A(new_n5173_), .B(new_n5172_), .Y(new_n5904_));
  AND2X1   g03468(.A(new_n5904_), .B(pi0096), .Y(new_n5905_));
  INVX1    g03469(.A(pi0122), .Y(new_n5906_));
  AND3X1   g03470(.A(new_n5225_), .B(pi0829), .C(new_n5906_), .Y(new_n5907_));
  INVX1    g03471(.A(new_n5907_), .Y(new_n5908_));
  OR4X1    g03472(.A(new_n5908_), .B(new_n5905_), .C(new_n5903_), .D(new_n5881_), .Y(new_n5909_));
  AOI21X1  g03473(.A0(new_n5909_), .A1(new_n5902_), .B0(pi1093), .Y(new_n5910_));
  INVX1    g03474(.A(new_n5910_), .Y(new_n5911_));
  INVX1    g03475(.A(po0740), .Y(new_n5912_));
  NOR3X1   g03476(.A(new_n5912_), .B(new_n2985_), .C(new_n2536_), .Y(new_n5913_));
  NOR4X1   g03477(.A(pi0100), .B(pi0075), .C(pi0039), .D(pi0038), .Y(new_n5914_));
  OAI21X1  g03478(.A0(new_n5913_), .A1(new_n3131_), .B0(new_n5914_), .Y(new_n5915_));
  AOI21X1  g03479(.A0(new_n5911_), .A1(new_n3131_), .B0(new_n5915_), .Y(new_n5916_));
  OAI21X1  g03480(.A0(new_n5916_), .A1(pi0567), .B0(new_n5880_), .Y(new_n5917_));
  NOR2X1   g03481(.A(new_n2961_), .B(pi0299), .Y(new_n5918_));
  NOR2X1   g03482(.A(new_n2450_), .B(new_n2933_), .Y(new_n5919_));
  NOR4X1   g03483(.A(new_n5919_), .B(new_n5918_), .C(new_n5048_), .D(new_n5215_), .Y(new_n5920_));
  NOR2X1   g03484(.A(new_n5920_), .B(new_n3074_), .Y(new_n5921_));
  AND2X1   g03485(.A(pi0957), .B(new_n2701_), .Y(new_n5922_));
  OR4X1    g03486(.A(new_n5908_), .B(new_n5082_), .C(new_n5922_), .D(new_n2702_), .Y(new_n5923_));
  NOR4X1   g03487(.A(new_n5923_), .B(new_n2986_), .C(new_n3035_), .D(pi0024), .Y(new_n5924_));
  AND3X1   g03488(.A(new_n5924_), .B(new_n5921_), .C(pi1093), .Y(new_n5925_));
  AOI21X1  g03489(.A0(pi0957), .A1(new_n2701_), .B0(new_n5032_), .Y(new_n5926_));
  AND3X1   g03490(.A(pi1092), .B(pi0950), .C(pi0824), .Y(new_n5927_));
  INVX1    g03491(.A(new_n5927_), .Y(new_n5928_));
  OR4X1    g03492(.A(new_n5889_), .B(new_n5881_), .C(new_n2847_), .D(pi0096), .Y(new_n5929_));
  OR3X1    g03493(.A(new_n5929_), .B(new_n5928_), .C(pi0829), .Y(new_n5930_));
  NAND3X1  g03494(.A(new_n2544_), .B(pi0091), .C(new_n5777_), .Y(new_n5931_));
  NAND4X1  g03495(.A(new_n5177_), .B(new_n2837_), .C(pi0097), .D(new_n2676_), .Y(new_n5932_));
  OR4X1    g03496(.A(new_n5932_), .B(new_n2561_), .C(new_n2559_), .D(pi0091), .Y(new_n5933_));
  NAND2X1  g03497(.A(new_n5933_), .B(new_n5931_), .Y(new_n5934_));
  NAND3X1  g03498(.A(new_n5934_), .B(new_n5885_), .C(new_n2501_), .Y(new_n5935_));
  AOI21X1  g03499(.A0(new_n5935_), .A1(new_n5889_), .B0(new_n2847_), .Y(new_n5936_));
  NOR3X1   g03500(.A(new_n5905_), .B(new_n5881_), .C(new_n2762_), .Y(new_n5937_));
  OAI21X1  g03501(.A0(new_n5936_), .A1(pi0096), .B0(new_n5937_), .Y(new_n5938_));
  AOI21X1  g03502(.A0(new_n5938_), .A1(new_n5930_), .B0(pi0122), .Y(new_n5939_));
  NOR3X1   g03503(.A(new_n5929_), .B(new_n5883_), .C(new_n5906_), .Y(new_n5940_));
  OAI21X1  g03504(.A0(new_n5940_), .A1(new_n5939_), .B0(new_n5926_), .Y(new_n5941_));
  AND2X1   g03505(.A(new_n5941_), .B(pi1091), .Y(new_n5942_));
  AND2X1   g03506(.A(new_n5942_), .B(new_n5911_), .Y(new_n5943_));
  NOR2X1   g03507(.A(new_n5910_), .B(pi1091), .Y(new_n5944_));
  OR2X1    g03508(.A(new_n5944_), .B(new_n5943_), .Y(new_n5945_));
  INVX1    g03509(.A(new_n5062_), .Y(new_n5946_));
  NOR4X1   g03510(.A(new_n5224_), .B(new_n2725_), .C(new_n2724_), .D(new_n5922_), .Y(new_n5947_));
  AND3X1   g03511(.A(new_n5947_), .B(new_n5946_), .C(pi1091), .Y(new_n5948_));
  AND3X1   g03512(.A(new_n5948_), .B(new_n5331_), .C(new_n2438_), .Y(new_n5949_));
  INVX1    g03513(.A(new_n5049_), .Y(new_n5950_));
  NOR4X1   g03514(.A(pi0299), .B(pi0224), .C(pi0223), .D(new_n2941_), .Y(new_n5951_));
  NAND4X1  g03515(.A(new_n5951_), .B(new_n5947_), .C(new_n5950_), .D(pi1091), .Y(new_n5952_));
  NAND2X1  g03516(.A(new_n5952_), .B(pi0039), .Y(new_n5953_));
  OAI21X1  g03517(.A0(new_n5953_), .A1(new_n5949_), .B0(new_n2979_), .Y(new_n5954_));
  AOI21X1  g03518(.A0(new_n5945_), .A1(new_n2939_), .B0(new_n5954_), .Y(new_n5955_));
  OR2X1    g03519(.A(new_n5955_), .B(pi0100), .Y(new_n5956_));
  NOR4X1   g03520(.A(new_n5954_), .B(new_n5942_), .C(new_n5929_), .D(new_n5228_), .Y(new_n5957_));
  NOR4X1   g03521(.A(new_n5908_), .B(new_n5082_), .C(new_n5922_), .D(new_n5032_), .Y(new_n5958_));
  INVX1    g03522(.A(new_n5958_), .Y(new_n5959_));
  NOR4X1   g03523(.A(new_n5959_), .B(new_n2985_), .C(new_n2536_), .D(new_n2702_), .Y(new_n5960_));
  NAND2X1  g03524(.A(new_n5960_), .B(pi0228), .Y(new_n5961_));
  NOR3X1   g03525(.A(new_n5961_), .B(new_n5920_), .C(new_n3060_), .Y(new_n5962_));
  NOR2X1   g03526(.A(new_n5962_), .B(new_n3007_), .Y(new_n5963_));
  INVX1    g03527(.A(new_n5963_), .Y(new_n5964_));
  OAI21X1  g03528(.A0(new_n5957_), .A1(new_n5956_), .B0(new_n5964_), .Y(new_n5965_));
  NOR3X1   g03529(.A(new_n5928_), .B(new_n2985_), .C(new_n2536_), .Y(new_n5966_));
  AND2X1   g03530(.A(pi1093), .B(new_n2702_), .Y(new_n5967_));
  INVX1    g03531(.A(new_n5967_), .Y(new_n5968_));
  NOR2X1   g03532(.A(new_n5968_), .B(new_n5966_), .Y(new_n5969_));
  AND3X1   g03533(.A(pi1093), .B(pi0957), .C(new_n2701_), .Y(new_n5970_));
  NOR4X1   g03534(.A(new_n5970_), .B(new_n5883_), .C(new_n2985_), .D(new_n2536_), .Y(new_n5971_));
  NOR2X1   g03535(.A(new_n5971_), .B(new_n5967_), .Y(new_n5972_));
  NOR3X1   g03536(.A(new_n5972_), .B(new_n5969_), .C(new_n3132_), .Y(new_n5973_));
  NOR2X1   g03537(.A(new_n5973_), .B(new_n3131_), .Y(new_n5974_));
  AOI21X1  g03538(.A0(new_n5965_), .A1(new_n3131_), .B0(new_n5974_), .Y(new_n5975_));
  MX2X1    g03539(.A(new_n5975_), .B(new_n5925_), .S0(pi0075), .Y(new_n5976_));
  INVX1    g03540(.A(new_n5976_), .Y(new_n5977_));
  AOI21X1  g03541(.A0(new_n5977_), .A1(pi0567), .B0(new_n5917_), .Y(new_n5978_));
  INVX1    g03542(.A(pi0567), .Y(new_n5979_));
  INVX1    g03543(.A(new_n5917_), .Y(new_n5980_));
  NOR2X1   g03544(.A(new_n5925_), .B(new_n3073_), .Y(new_n5981_));
  NOR2X1   g03545(.A(new_n5963_), .B(pi0087), .Y(new_n5982_));
  AND2X1   g03546(.A(new_n5982_), .B(new_n5956_), .Y(new_n5983_));
  NOR2X1   g03547(.A(new_n5971_), .B(new_n2702_), .Y(new_n5984_));
  NOR2X1   g03548(.A(new_n5913_), .B(pi1091), .Y(new_n5985_));
  NAND3X1  g03549(.A(new_n3047_), .B(new_n3007_), .C(pi0087), .Y(new_n5986_));
  NOR3X1   g03550(.A(new_n5986_), .B(new_n5985_), .C(new_n5984_), .Y(new_n5987_));
  NOR3X1   g03551(.A(new_n5987_), .B(new_n5983_), .C(pi0075), .Y(new_n5988_));
  NOR2X1   g03552(.A(new_n5988_), .B(new_n5981_), .Y(new_n5989_));
  OAI21X1  g03553(.A0(new_n5989_), .A1(new_n5979_), .B0(new_n5980_), .Y(new_n5990_));
  INVX1    g03554(.A(new_n5990_), .Y(new_n5991_));
  MX2X1    g03555(.A(new_n5991_), .B(new_n5978_), .S0(pi0592), .Y(new_n5992_));
  INVX1    g03556(.A(new_n5992_), .Y(new_n5993_));
  INVX1    g03557(.A(new_n5978_), .Y(new_n5994_));
  OR2X1    g03558(.A(pi0592), .B(pi0350), .Y(new_n5995_));
  INVX1    g03559(.A(pi0321), .Y(new_n5996_));
  XOR2X1   g03560(.A(pi0347), .B(new_n5996_), .Y(new_n5997_));
  XOR2X1   g03561(.A(pi0349), .B(pi0316), .Y(new_n5998_));
  XOR2X1   g03562(.A(new_n5998_), .B(pi0348), .Y(new_n5999_));
  INVX1    g03563(.A(pi0322), .Y(new_n6000_));
  XOR2X1   g03564(.A(pi0359), .B(pi0315), .Y(new_n6001_));
  XOR2X1   g03565(.A(new_n6001_), .B(new_n6000_), .Y(new_n6002_));
  XOR2X1   g03566(.A(new_n6002_), .B(new_n5999_), .Y(new_n6003_));
  XOR2X1   g03567(.A(new_n6003_), .B(new_n5997_), .Y(new_n6004_));
  OAI21X1  g03568(.A0(new_n5991_), .A1(new_n5995_), .B0(new_n6004_), .Y(new_n6005_));
  AOI21X1  g03569(.A0(new_n5995_), .A1(new_n5994_), .B0(new_n6005_), .Y(new_n6006_));
  INVX1    g03570(.A(pi0350), .Y(new_n6007_));
  OR2X1    g03571(.A(pi0592), .B(new_n6007_), .Y(new_n6008_));
  INVX1    g03572(.A(pi0592), .Y(new_n6009_));
  AND3X1   g03573(.A(new_n5990_), .B(new_n6009_), .C(pi0350), .Y(new_n6010_));
  OR2X1    g03574(.A(new_n6010_), .B(new_n6004_), .Y(new_n6011_));
  AOI21X1  g03575(.A0(new_n6008_), .A1(new_n5994_), .B0(new_n6011_), .Y(new_n6012_));
  INVX1    g03576(.A(pi0355), .Y(new_n6013_));
  XOR2X1   g03577(.A(pi0455), .B(pi0452), .Y(new_n6014_));
  XOR2X1   g03578(.A(new_n6014_), .B(new_n6013_), .Y(new_n6015_));
  XOR2X1   g03579(.A(pi0460), .B(pi0320), .Y(new_n6016_));
  XOR2X1   g03580(.A(new_n6016_), .B(pi0342), .Y(new_n6017_));
  INVX1    g03581(.A(pi0361), .Y(new_n6018_));
  XOR2X1   g03582(.A(pi0441), .B(new_n6018_), .Y(new_n6019_));
  XOR2X1   g03583(.A(new_n6019_), .B(new_n6017_), .Y(new_n6020_));
  XOR2X1   g03584(.A(new_n6020_), .B(pi0458), .Y(new_n6021_));
  XOR2X1   g03585(.A(new_n6021_), .B(new_n6015_), .Y(new_n6022_));
  AND2X1   g03586(.A(new_n6022_), .B(pi1196), .Y(new_n6023_));
  OR2X1    g03587(.A(new_n6023_), .B(new_n6012_), .Y(new_n6024_));
  INVX1    g03588(.A(pi1198), .Y(new_n6025_));
  AOI21X1  g03589(.A0(new_n5993_), .A1(new_n6023_), .B0(new_n6025_), .Y(new_n6026_));
  OAI21X1  g03590(.A0(new_n6024_), .A1(new_n6006_), .B0(new_n6026_), .Y(new_n6027_));
  INVX1    g03591(.A(new_n6020_), .Y(new_n6028_));
  INVX1    g03592(.A(pi0458), .Y(new_n6029_));
  INVX1    g03593(.A(pi0452), .Y(new_n6030_));
  MX2X1    g03594(.A(new_n5992_), .B(new_n5978_), .S0(pi0455), .Y(new_n6031_));
  INVX1    g03595(.A(pi0455), .Y(new_n6032_));
  MX2X1    g03596(.A(new_n5992_), .B(new_n5978_), .S0(new_n6032_), .Y(new_n6033_));
  MX2X1    g03597(.A(new_n6033_), .B(new_n6031_), .S0(new_n6030_), .Y(new_n6034_));
  MX2X1    g03598(.A(new_n6033_), .B(new_n6031_), .S0(pi0452), .Y(new_n6035_));
  MX2X1    g03599(.A(new_n6035_), .B(new_n6034_), .S0(new_n6013_), .Y(new_n6036_));
  NOR2X1   g03600(.A(new_n6036_), .B(new_n6029_), .Y(new_n6037_));
  MX2X1    g03601(.A(new_n6035_), .B(new_n6034_), .S0(pi0355), .Y(new_n6038_));
  NOR2X1   g03602(.A(new_n6038_), .B(pi0458), .Y(new_n6039_));
  OR3X1    g03603(.A(new_n6039_), .B(new_n6037_), .C(new_n6028_), .Y(new_n6040_));
  INVX1    g03604(.A(new_n6040_), .Y(new_n6041_));
  NOR2X1   g03605(.A(new_n6038_), .B(new_n6029_), .Y(new_n6042_));
  OAI21X1  g03606(.A0(new_n6036_), .A1(pi0458), .B0(new_n6028_), .Y(new_n6043_));
  OAI21X1  g03607(.A0(new_n6043_), .A1(new_n6042_), .B0(pi1196), .Y(new_n6044_));
  INVX1    g03608(.A(pi1196), .Y(new_n6045_));
  AOI21X1  g03609(.A0(new_n5994_), .A1(new_n6045_), .B0(pi1198), .Y(new_n6046_));
  OAI21X1  g03610(.A0(new_n6044_), .A1(new_n6041_), .B0(new_n6046_), .Y(new_n6047_));
  AND2X1   g03611(.A(new_n6047_), .B(new_n6027_), .Y(new_n6048_));
  MX2X1    g03612(.A(new_n6048_), .B(new_n5993_), .S0(new_n5879_), .Y(new_n6049_));
  INVX1    g03613(.A(pi0351), .Y(new_n6050_));
  AND2X1   g03614(.A(pi1199), .B(new_n6050_), .Y(new_n6051_));
  INVX1    g03615(.A(new_n6051_), .Y(new_n6052_));
  INVX1    g03616(.A(pi1199), .Y(new_n6053_));
  NOR3X1   g03617(.A(new_n5992_), .B(new_n6053_), .C(pi0351), .Y(new_n6054_));
  AOI21X1  g03618(.A0(new_n6052_), .A1(new_n6049_), .B0(new_n6054_), .Y(new_n6055_));
  AND2X1   g03619(.A(pi1199), .B(pi0351), .Y(new_n6056_));
  INVX1    g03620(.A(new_n6056_), .Y(new_n6057_));
  NOR3X1   g03621(.A(new_n5992_), .B(new_n6053_), .C(new_n6050_), .Y(new_n6058_));
  AOI21X1  g03622(.A0(new_n6057_), .A1(new_n6049_), .B0(new_n6058_), .Y(new_n6059_));
  MX2X1    g03623(.A(new_n6059_), .B(new_n6055_), .S0(new_n5866_), .Y(new_n6060_));
  MX2X1    g03624(.A(new_n6059_), .B(new_n6055_), .S0(pi0461), .Y(new_n6061_));
  MX2X1    g03625(.A(new_n6061_), .B(new_n6060_), .S0(new_n5865_), .Y(new_n6062_));
  MX2X1    g03626(.A(new_n6061_), .B(new_n6060_), .S0(pi0357), .Y(new_n6063_));
  MX2X1    g03627(.A(new_n6063_), .B(new_n6062_), .S0(new_n5864_), .Y(new_n6064_));
  OR2X1    g03628(.A(new_n6064_), .B(new_n5863_), .Y(new_n6065_));
  OR2X1    g03629(.A(new_n6063_), .B(pi0356), .Y(new_n6066_));
  OAI21X1  g03630(.A0(new_n6062_), .A1(new_n5864_), .B0(new_n6066_), .Y(new_n6067_));
  AOI21X1  g03631(.A0(new_n6067_), .A1(new_n5863_), .B0(pi0591), .Y(new_n6068_));
  INVX1    g03632(.A(pi0591), .Y(new_n6069_));
  OAI21X1  g03633(.A0(new_n5994_), .A1(new_n6069_), .B0(pi0590), .Y(new_n6070_));
  AOI21X1  g03634(.A0(new_n6068_), .A1(new_n6065_), .B0(new_n6070_), .Y(new_n6071_));
  NOR4X1   g03635(.A(pi0289), .B(pi0288), .C(pi0286), .D(pi0285), .Y(new_n6072_));
  INVX1    g03636(.A(new_n6072_), .Y(new_n6073_));
  INVX1    g03637(.A(pi0375), .Y(new_n6074_));
  INVX1    g03638(.A(pi0373), .Y(new_n6075_));
  INVX1    g03639(.A(pi0371), .Y(new_n6076_));
  INVX1    g03640(.A(pi0370), .Y(new_n6077_));
  INVX1    g03641(.A(pi0369), .Y(new_n6078_));
  INVX1    g03642(.A(pi0374), .Y(new_n6079_));
  XOR2X1   g03643(.A(pi0372), .B(pi0363), .Y(new_n6080_));
  XOR2X1   g03644(.A(new_n6080_), .B(pi0386), .Y(new_n6081_));
  XOR2X1   g03645(.A(pi0388), .B(pi0338), .Y(new_n6082_));
  XOR2X1   g03646(.A(pi0339), .B(pi0337), .Y(new_n6083_));
  XOR2X1   g03647(.A(new_n6083_), .B(pi0387), .Y(new_n6084_));
  XOR2X1   g03648(.A(new_n6084_), .B(pi0380), .Y(new_n6085_));
  XOR2X1   g03649(.A(new_n6085_), .B(new_n6082_), .Y(new_n6086_));
  XOR2X1   g03650(.A(new_n6086_), .B(new_n6081_), .Y(new_n6087_));
  AND2X1   g03651(.A(new_n6087_), .B(pi1196), .Y(new_n6088_));
  XOR2X1   g03652(.A(pi0389), .B(pi0368), .Y(new_n6089_));
  INVX1    g03653(.A(pi0367), .Y(new_n6090_));
  XOR2X1   g03654(.A(pi0447), .B(pi0365), .Y(new_n6091_));
  INVX1    g03655(.A(new_n6091_), .Y(new_n6092_));
  XOR2X1   g03656(.A(pi0383), .B(pi0336), .Y(new_n6093_));
  XOR2X1   g03657(.A(pi0366), .B(pi0364), .Y(new_n6094_));
  XOR2X1   g03658(.A(new_n6094_), .B(new_n6093_), .Y(new_n6095_));
  XOR2X1   g03659(.A(new_n6095_), .B(new_n6092_), .Y(new_n6096_));
  XOR2X1   g03660(.A(new_n6096_), .B(new_n6090_), .Y(new_n6097_));
  OAI21X1  g03661(.A0(new_n6097_), .A1(new_n6089_), .B0(pi1197), .Y(new_n6098_));
  AOI21X1  g03662(.A0(new_n6097_), .A1(new_n6089_), .B0(new_n6098_), .Y(new_n6099_));
  NOR2X1   g03663(.A(new_n6099_), .B(new_n6088_), .Y(new_n6100_));
  AND2X1   g03664(.A(pi0592), .B(pi0377), .Y(new_n6101_));
  XOR2X1   g03665(.A(pi0382), .B(pi0379), .Y(new_n6102_));
  XOR2X1   g03666(.A(pi0439), .B(pi0376), .Y(new_n6103_));
  XOR2X1   g03667(.A(new_n6103_), .B(pi0381), .Y(new_n6104_));
  INVX1    g03668(.A(pi0378), .Y(new_n6105_));
  XOR2X1   g03669(.A(pi0385), .B(pi0317), .Y(new_n6106_));
  XOR2X1   g03670(.A(new_n6106_), .B(new_n6105_), .Y(new_n6107_));
  XOR2X1   g03671(.A(new_n6107_), .B(new_n6104_), .Y(new_n6108_));
  XOR2X1   g03672(.A(new_n6108_), .B(new_n6102_), .Y(new_n6109_));
  INVX1    g03673(.A(new_n6109_), .Y(new_n6110_));
  AOI21X1  g03674(.A0(new_n6101_), .A1(new_n5990_), .B0(new_n6110_), .Y(new_n6111_));
  OAI21X1  g03675(.A0(new_n6101_), .A1(new_n5978_), .B0(new_n6111_), .Y(new_n6112_));
  INVX1    g03676(.A(pi0377), .Y(new_n6113_));
  AND2X1   g03677(.A(pi0592), .B(new_n6113_), .Y(new_n6114_));
  AOI21X1  g03678(.A0(new_n6114_), .A1(new_n5990_), .B0(new_n6109_), .Y(new_n6115_));
  OAI21X1  g03679(.A0(new_n6114_), .A1(new_n5978_), .B0(new_n6115_), .Y(new_n6116_));
  NAND2X1  g03680(.A(new_n6116_), .B(new_n6112_), .Y(new_n6117_));
  MX2X1    g03681(.A(new_n5991_), .B(new_n5978_), .S0(new_n6009_), .Y(new_n6118_));
  MX2X1    g03682(.A(new_n6118_), .B(new_n6117_), .S0(new_n6100_), .Y(new_n6119_));
  NOR2X1   g03683(.A(new_n6119_), .B(new_n6053_), .Y(new_n6120_));
  INVX1    g03684(.A(new_n6087_), .Y(new_n6121_));
  MX2X1    g03685(.A(new_n5978_), .B(new_n6118_), .S0(new_n6099_), .Y(new_n6122_));
  AND2X1   g03686(.A(new_n6122_), .B(new_n6121_), .Y(new_n6123_));
  OAI21X1  g03687(.A0(new_n6099_), .A1(pi1196), .B0(new_n6118_), .Y(new_n6124_));
  OR3X1    g03688(.A(new_n6099_), .B(new_n5994_), .C(pi1196), .Y(new_n6125_));
  AOI21X1  g03689(.A0(new_n6125_), .A1(new_n6124_), .B0(new_n6121_), .Y(new_n6126_));
  NOR3X1   g03690(.A(new_n6126_), .B(new_n6123_), .C(pi1199), .Y(new_n6127_));
  OAI21X1  g03691(.A0(new_n6127_), .A1(new_n6120_), .B0(new_n6079_), .Y(new_n6128_));
  AND2X1   g03692(.A(pi1199), .B(new_n6025_), .Y(new_n6129_));
  INVX1    g03693(.A(new_n6129_), .Y(new_n6130_));
  OAI22X1  g03694(.A0(new_n6130_), .A1(new_n6119_), .B0(new_n6118_), .B1(new_n6025_), .Y(new_n6131_));
  AOI21X1  g03695(.A0(new_n6127_), .A1(new_n6025_), .B0(new_n6131_), .Y(new_n6132_));
  OAI21X1  g03696(.A0(new_n6132_), .A1(new_n6079_), .B0(new_n6128_), .Y(new_n6133_));
  AND2X1   g03697(.A(new_n6133_), .B(pi0369), .Y(new_n6134_));
  OAI21X1  g03698(.A0(new_n6127_), .A1(new_n6120_), .B0(pi0374), .Y(new_n6135_));
  OAI21X1  g03699(.A0(new_n6132_), .A1(pi0374), .B0(new_n6135_), .Y(new_n6136_));
  AOI21X1  g03700(.A0(new_n6136_), .A1(new_n6078_), .B0(new_n6134_), .Y(new_n6137_));
  OR2X1    g03701(.A(new_n6137_), .B(pi0370), .Y(new_n6138_));
  AND2X1   g03702(.A(new_n6133_), .B(new_n6078_), .Y(new_n6139_));
  AOI21X1  g03703(.A0(new_n6136_), .A1(pi0369), .B0(new_n6139_), .Y(new_n6140_));
  OAI21X1  g03704(.A0(new_n6140_), .A1(new_n6077_), .B0(new_n6138_), .Y(new_n6141_));
  AND2X1   g03705(.A(new_n6141_), .B(new_n6076_), .Y(new_n6142_));
  OR2X1    g03706(.A(new_n6140_), .B(pi0370), .Y(new_n6143_));
  OAI21X1  g03707(.A0(new_n6137_), .A1(new_n6077_), .B0(new_n6143_), .Y(new_n6144_));
  AOI21X1  g03708(.A0(new_n6144_), .A1(pi0371), .B0(new_n6142_), .Y(new_n6145_));
  AND2X1   g03709(.A(new_n6144_), .B(new_n6076_), .Y(new_n6146_));
  AOI21X1  g03710(.A0(new_n6141_), .A1(pi0371), .B0(new_n6146_), .Y(new_n6147_));
  MX2X1    g03711(.A(new_n6147_), .B(new_n6145_), .S0(new_n6075_), .Y(new_n6148_));
  NAND2X1  g03712(.A(new_n6148_), .B(new_n6074_), .Y(new_n6149_));
  XOR2X1   g03713(.A(pi0442), .B(pi0384), .Y(new_n6150_));
  XOR2X1   g03714(.A(new_n6150_), .B(pi0440), .Y(new_n6151_));
  INVX1    g03715(.A(new_n6151_), .Y(new_n6152_));
  MX2X1    g03716(.A(new_n6147_), .B(new_n6145_), .S0(pi0373), .Y(new_n6153_));
  AOI21X1  g03717(.A0(new_n6153_), .A1(pi0375), .B0(new_n6152_), .Y(new_n6154_));
  NAND2X1  g03718(.A(new_n6154_), .B(new_n6149_), .Y(new_n6155_));
  NAND2X1  g03719(.A(new_n6148_), .B(pi0375), .Y(new_n6156_));
  AOI21X1  g03720(.A0(new_n6153_), .A1(new_n6074_), .B0(new_n6151_), .Y(new_n6157_));
  AOI21X1  g03721(.A0(new_n6157_), .A1(new_n6156_), .B0(pi0591), .Y(new_n6158_));
  INVX1    g03722(.A(pi0334), .Y(new_n6159_));
  INVX1    g03723(.A(pi0393), .Y(new_n6160_));
  INVX1    g03724(.A(pi0392), .Y(new_n6161_));
  INVX1    g03725(.A(pi0333), .Y(new_n6162_));
  INVX1    g03726(.A(pi0328), .Y(new_n6163_));
  XOR2X1   g03727(.A(pi0408), .B(new_n6163_), .Y(new_n6164_));
  XOR2X1   g03728(.A(pi0396), .B(pi0394), .Y(new_n6165_));
  XOR2X1   g03729(.A(new_n6165_), .B(new_n6164_), .Y(new_n6166_));
  INVX1    g03730(.A(pi0395), .Y(new_n6167_));
  XOR2X1   g03731(.A(pi0399), .B(pi0398), .Y(new_n6168_));
  XOR2X1   g03732(.A(new_n6168_), .B(new_n6167_), .Y(new_n6169_));
  XOR2X1   g03733(.A(new_n6169_), .B(pi0329), .Y(new_n6170_));
  XOR2X1   g03734(.A(new_n6170_), .B(pi0400), .Y(new_n6171_));
  XOR2X1   g03735(.A(new_n6171_), .B(new_n6166_), .Y(new_n6172_));
  AND2X1   g03736(.A(new_n6172_), .B(pi1198), .Y(new_n6173_));
  INVX1    g03737(.A(pi0411), .Y(new_n6174_));
  XOR2X1   g03738(.A(pi0410), .B(pi0390), .Y(new_n6175_));
  XOR2X1   g03739(.A(pi0412), .B(pi0397), .Y(new_n6176_));
  XOR2X1   g03740(.A(new_n6176_), .B(pi0404), .Y(new_n6177_));
  XOR2X1   g03741(.A(pi0324), .B(pi0319), .Y(new_n6178_));
  XOR2X1   g03742(.A(new_n6178_), .B(pi0456), .Y(new_n6179_));
  XOR2X1   g03743(.A(new_n6179_), .B(new_n6177_), .Y(new_n6180_));
  XOR2X1   g03744(.A(new_n6180_), .B(new_n6175_), .Y(new_n6181_));
  XOR2X1   g03745(.A(new_n6181_), .B(new_n6174_), .Y(new_n6182_));
  AOI21X1  g03746(.A0(new_n6182_), .A1(new_n5957_), .B0(new_n5956_), .Y(new_n6183_));
  NOR3X1   g03747(.A(new_n6183_), .B(new_n5963_), .C(pi0087), .Y(new_n6184_));
  AOI21X1  g03748(.A0(new_n6182_), .A1(new_n5966_), .B0(new_n5968_), .Y(new_n6185_));
  NOR3X1   g03749(.A(new_n6185_), .B(new_n5986_), .C(new_n5972_), .Y(new_n6186_));
  NOR2X1   g03750(.A(pi0592), .B(pi0075), .Y(new_n6187_));
  INVX1    g03751(.A(new_n6187_), .Y(new_n6188_));
  OR3X1    g03752(.A(new_n6188_), .B(new_n6186_), .C(new_n6045_), .Y(new_n6189_));
  OR2X1    g03753(.A(new_n6189_), .B(new_n6184_), .Y(new_n6190_));
  OR3X1    g03754(.A(new_n5975_), .B(pi1196), .C(pi0075), .Y(new_n6191_));
  AOI21X1  g03755(.A0(new_n6191_), .A1(new_n6190_), .B0(pi1199), .Y(new_n6192_));
  INVX1    g03756(.A(new_n6192_), .Y(new_n6193_));
  XOR2X1   g03757(.A(pi0409), .B(pi0318), .Y(new_n6194_));
  INVX1    g03758(.A(pi0406), .Y(new_n6195_));
  XOR2X1   g03759(.A(pi0402), .B(pi0401), .Y(new_n6196_));
  XOR2X1   g03760(.A(new_n6196_), .B(new_n6195_), .Y(new_n6197_));
  XOR2X1   g03761(.A(pi0405), .B(pi0403), .Y(new_n6198_));
  XOR2X1   g03762(.A(pi0326), .B(pi0325), .Y(new_n6199_));
  XOR2X1   g03763(.A(new_n6199_), .B(new_n6198_), .Y(new_n6200_));
  XOR2X1   g03764(.A(new_n6200_), .B(new_n6197_), .Y(new_n6201_));
  XOR2X1   g03765(.A(new_n6201_), .B(new_n6194_), .Y(new_n6202_));
  OR3X1    g03766(.A(new_n6182_), .B(new_n6045_), .C(pi0075), .Y(new_n6203_));
  AND3X1   g03767(.A(new_n6203_), .B(new_n6202_), .C(new_n5957_), .Y(new_n6204_));
  OAI21X1  g03768(.A0(new_n6204_), .A1(new_n5956_), .B0(new_n5982_), .Y(new_n6205_));
  AOI21X1  g03769(.A0(new_n6202_), .A1(new_n5966_), .B0(new_n5968_), .Y(new_n6206_));
  NOR4X1   g03770(.A(new_n6206_), .B(new_n5986_), .C(new_n5972_), .D(pi1196), .Y(new_n6207_));
  NOR4X1   g03771(.A(new_n6206_), .B(new_n6185_), .C(new_n5986_), .D(new_n5972_), .Y(new_n6208_));
  NOR4X1   g03772(.A(new_n6208_), .B(new_n6207_), .C(new_n6188_), .D(new_n6053_), .Y(new_n6209_));
  AOI22X1  g03773(.A0(new_n6209_), .A1(new_n6205_), .B0(new_n6188_), .B1(new_n5977_), .Y(new_n6210_));
  AOI21X1  g03774(.A0(new_n6210_), .A1(new_n6193_), .B0(new_n5979_), .Y(new_n6211_));
  NOR3X1   g03775(.A(new_n6211_), .B(new_n6173_), .C(new_n5917_), .Y(new_n6212_));
  AOI21X1  g03776(.A0(new_n6173_), .A1(new_n5992_), .B0(new_n6212_), .Y(new_n6213_));
  INVX1    g03777(.A(new_n6213_), .Y(new_n6214_));
  MX2X1    g03778(.A(new_n6214_), .B(new_n5992_), .S0(pi1197), .Y(new_n6215_));
  MX2X1    g03779(.A(new_n6215_), .B(new_n6214_), .S0(new_n6162_), .Y(new_n6216_));
  MX2X1    g03780(.A(new_n6215_), .B(new_n6214_), .S0(pi0333), .Y(new_n6217_));
  MX2X1    g03781(.A(new_n6217_), .B(new_n6216_), .S0(pi0391), .Y(new_n6218_));
  INVX1    g03782(.A(pi0391), .Y(new_n6219_));
  MX2X1    g03783(.A(new_n6217_), .B(new_n6216_), .S0(new_n6219_), .Y(new_n6220_));
  MX2X1    g03784(.A(new_n6220_), .B(new_n6218_), .S0(new_n6161_), .Y(new_n6221_));
  MX2X1    g03785(.A(new_n6220_), .B(new_n6218_), .S0(pi0392), .Y(new_n6222_));
  MX2X1    g03786(.A(new_n6222_), .B(new_n6221_), .S0(new_n6160_), .Y(new_n6223_));
  NAND2X1  g03787(.A(new_n6223_), .B(new_n6159_), .Y(new_n6224_));
  XOR2X1   g03788(.A(pi0463), .B(pi0407), .Y(new_n6225_));
  XOR2X1   g03789(.A(pi0413), .B(pi0335), .Y(new_n6226_));
  XOR2X1   g03790(.A(new_n6226_), .B(new_n6225_), .Y(new_n6227_));
  MX2X1    g03791(.A(new_n6222_), .B(new_n6221_), .S0(pi0393), .Y(new_n6228_));
  NAND2X1  g03792(.A(new_n6228_), .B(pi0334), .Y(new_n6229_));
  AND3X1   g03793(.A(new_n6229_), .B(new_n6227_), .C(new_n6224_), .Y(new_n6230_));
  AND2X1   g03794(.A(new_n6228_), .B(new_n6159_), .Y(new_n6231_));
  AND2X1   g03795(.A(new_n6223_), .B(pi0334), .Y(new_n6232_));
  NOR3X1   g03796(.A(new_n6232_), .B(new_n6231_), .C(new_n6227_), .Y(new_n6233_));
  NOR3X1   g03797(.A(new_n6233_), .B(new_n6230_), .C(new_n6069_), .Y(new_n6234_));
  OR2X1    g03798(.A(new_n6234_), .B(pi0590), .Y(new_n6235_));
  AOI21X1  g03799(.A0(new_n6158_), .A1(new_n6155_), .B0(new_n6235_), .Y(new_n6236_));
  OR2X1    g03800(.A(new_n6236_), .B(new_n6073_), .Y(new_n6237_));
  INVX1    g03801(.A(new_n5921_), .Y(new_n6238_));
  NOR4X1   g03802(.A(new_n2985_), .B(new_n2536_), .C(new_n3035_), .D(pi0024), .Y(new_n6239_));
  AOI21X1  g03803(.A0(new_n5958_), .A1(new_n6239_), .B0(new_n2702_), .Y(new_n6240_));
  NOR2X1   g03804(.A(new_n6240_), .B(new_n6238_), .Y(new_n6241_));
  INVX1    g03805(.A(new_n6241_), .Y(new_n6242_));
  AND2X1   g03806(.A(pi1093), .B(new_n5906_), .Y(new_n6243_));
  AND2X1   g03807(.A(new_n5927_), .B(new_n5893_), .Y(new_n6244_));
  AOI21X1  g03808(.A0(new_n6244_), .A1(new_n6243_), .B0(pi1091), .Y(new_n6245_));
  AND3X1   g03809(.A(new_n5927_), .B(pi1093), .C(new_n5906_), .Y(new_n6246_));
  AND3X1   g03810(.A(new_n6246_), .B(new_n2702_), .C(new_n5893_), .Y(new_n6247_));
  AOI21X1  g03811(.A0(new_n6247_), .A1(new_n6238_), .B0(new_n3073_), .Y(new_n6248_));
  OAI21X1  g03812(.A0(new_n6245_), .A1(new_n6242_), .B0(new_n6248_), .Y(new_n6249_));
  OR2X1    g03813(.A(new_n5943_), .B(pi0039), .Y(new_n6250_));
  AND3X1   g03814(.A(new_n5927_), .B(new_n5906_), .C(new_n5893_), .Y(new_n6251_));
  NOR3X1   g03815(.A(new_n5929_), .B(new_n5928_), .C(new_n5906_), .Y(new_n6252_));
  OAI21X1  g03816(.A0(new_n6252_), .A1(new_n6251_), .B0(pi1093), .Y(new_n6253_));
  AOI21X1  g03817(.A0(new_n6253_), .A1(new_n5944_), .B0(new_n6250_), .Y(new_n6254_));
  NOR2X1   g03818(.A(new_n5023_), .B(new_n5021_), .Y(new_n6255_));
  INVX1    g03819(.A(new_n6255_), .Y(new_n6256_));
  INVX1    g03820(.A(new_n6247_), .Y(new_n6257_));
  AND2X1   g03821(.A(new_n6244_), .B(new_n6243_), .Y(new_n6258_));
  OR2X1    g03822(.A(new_n6258_), .B(pi1091), .Y(new_n6259_));
  OAI21X1  g03823(.A0(new_n5947_), .A1(new_n2702_), .B0(new_n6259_), .Y(new_n6260_));
  MX2X1    g03824(.A(new_n6260_), .B(new_n6257_), .S0(new_n6256_), .Y(new_n6261_));
  NAND2X1  g03825(.A(new_n6261_), .B(new_n5041_), .Y(new_n6262_));
  MX2X1    g03826(.A(new_n6260_), .B(new_n6257_), .S0(new_n5043_), .Y(new_n6263_));
  AND3X1   g03827(.A(new_n2942_), .B(new_n2940_), .C(pi0222), .Y(new_n6264_));
  INVX1    g03828(.A(new_n6264_), .Y(new_n6265_));
  AOI21X1  g03829(.A0(new_n6263_), .A1(new_n5042_), .B0(new_n6265_), .Y(new_n6266_));
  OAI21X1  g03830(.A0(new_n6264_), .A1(new_n6257_), .B0(new_n2933_), .Y(new_n6267_));
  AOI21X1  g03831(.A0(new_n6266_), .A1(new_n6262_), .B0(new_n6267_), .Y(new_n6268_));
  NAND2X1  g03832(.A(new_n6261_), .B(new_n5058_), .Y(new_n6269_));
  AND3X1   g03833(.A(pi0221), .B(new_n2438_), .C(new_n2934_), .Y(new_n6270_));
  INVX1    g03834(.A(new_n6270_), .Y(new_n6271_));
  AOI21X1  g03835(.A0(new_n6263_), .A1(new_n5059_), .B0(new_n6271_), .Y(new_n6272_));
  OAI21X1  g03836(.A0(new_n6270_), .A1(new_n6257_), .B0(pi0299), .Y(new_n6273_));
  AOI21X1  g03837(.A0(new_n6272_), .A1(new_n6269_), .B0(new_n6273_), .Y(new_n6274_));
  NOR3X1   g03838(.A(new_n6274_), .B(new_n6268_), .C(new_n2939_), .Y(new_n6275_));
  OAI21X1  g03839(.A0(new_n6275_), .A1(new_n6254_), .B0(new_n2979_), .Y(new_n6276_));
  AOI21X1  g03840(.A0(new_n6247_), .A1(pi0038), .B0(pi0100), .Y(new_n6277_));
  NOR2X1   g03841(.A(new_n5920_), .B(new_n2793_), .Y(new_n6278_));
  OR3X1    g03842(.A(new_n5959_), .B(new_n2985_), .C(new_n2536_), .Y(new_n6279_));
  INVX1    g03843(.A(new_n6258_), .Y(new_n6280_));
  MX2X1    g03844(.A(new_n6280_), .B(new_n6279_), .S0(pi1091), .Y(new_n6281_));
  OAI21X1  g03845(.A0(new_n6278_), .A1(new_n6247_), .B0(new_n3047_), .Y(new_n6282_));
  AOI21X1  g03846(.A0(new_n6281_), .A1(new_n6278_), .B0(new_n6282_), .Y(new_n6283_));
  OAI21X1  g03847(.A0(new_n6257_), .A1(new_n3047_), .B0(pi0100), .Y(new_n6284_));
  OAI21X1  g03848(.A0(new_n6284_), .A1(new_n6283_), .B0(new_n3131_), .Y(new_n6285_));
  AOI21X1  g03849(.A0(new_n6277_), .A1(new_n6276_), .B0(new_n6285_), .Y(new_n6286_));
  NOR4X1   g03850(.A(new_n5928_), .B(new_n2985_), .C(new_n2536_), .D(new_n5906_), .Y(new_n6287_));
  OAI21X1  g03851(.A0(new_n6287_), .A1(new_n6251_), .B0(pi1093), .Y(new_n6288_));
  OAI21X1  g03852(.A0(new_n5971_), .A1(new_n2702_), .B0(new_n3064_), .Y(new_n6289_));
  AOI21X1  g03853(.A0(new_n6288_), .A1(new_n5985_), .B0(new_n6289_), .Y(new_n6290_));
  OAI21X1  g03854(.A0(new_n6290_), .A1(new_n6247_), .B0(pi0087), .Y(new_n6291_));
  NAND2X1  g03855(.A(new_n6291_), .B(new_n3073_), .Y(new_n6292_));
  OAI21X1  g03856(.A0(new_n6292_), .A1(new_n6286_), .B0(new_n6249_), .Y(new_n6293_));
  AOI21X1  g03857(.A0(new_n6293_), .A1(pi0567), .B0(new_n5917_), .Y(new_n6294_));
  INVX1    g03858(.A(new_n5880_), .Y(new_n6295_));
  AND3X1   g03859(.A(new_n6247_), .B(new_n6295_), .C(pi0567), .Y(new_n6296_));
  NOR3X1   g03860(.A(new_n6296_), .B(new_n6294_), .C(new_n6009_), .Y(new_n6297_));
  AOI21X1  g03861(.A0(new_n5990_), .A1(new_n6009_), .B0(new_n6297_), .Y(new_n6298_));
  NOR2X1   g03862(.A(new_n6296_), .B(new_n6294_), .Y(new_n6299_));
  INVX1    g03863(.A(new_n6298_), .Y(new_n6300_));
  MX2X1    g03864(.A(new_n6300_), .B(new_n6299_), .S0(new_n6032_), .Y(new_n6301_));
  AND2X1   g03865(.A(new_n6301_), .B(new_n6030_), .Y(new_n6302_));
  XOR2X1   g03866(.A(new_n6021_), .B(new_n6013_), .Y(new_n6303_));
  INVX1    g03867(.A(new_n6303_), .Y(new_n6304_));
  INVX1    g03868(.A(new_n6299_), .Y(new_n6305_));
  MX2X1    g03869(.A(new_n6298_), .B(new_n6305_), .S0(pi0455), .Y(new_n6306_));
  OAI21X1  g03870(.A0(new_n6306_), .A1(new_n6030_), .B0(new_n6304_), .Y(new_n6307_));
  OR2X1    g03871(.A(new_n6307_), .B(new_n6302_), .Y(new_n6308_));
  AOI21X1  g03872(.A0(new_n6301_), .A1(pi0452), .B0(new_n6304_), .Y(new_n6309_));
  OAI21X1  g03873(.A0(new_n6306_), .A1(pi0452), .B0(new_n6309_), .Y(new_n6310_));
  AND3X1   g03874(.A(new_n6310_), .B(new_n6308_), .C(pi1196), .Y(new_n6311_));
  NOR3X1   g03875(.A(new_n6296_), .B(new_n6294_), .C(pi1196), .Y(new_n6312_));
  OR2X1    g03876(.A(new_n6312_), .B(pi1198), .Y(new_n6313_));
  AOI21X1  g03877(.A0(new_n6299_), .A1(new_n6008_), .B0(new_n6011_), .Y(new_n6314_));
  AOI21X1  g03878(.A0(new_n6299_), .A1(new_n5995_), .B0(new_n6005_), .Y(new_n6315_));
  OR3X1    g03879(.A(new_n6315_), .B(new_n6314_), .C(new_n6023_), .Y(new_n6316_));
  AOI21X1  g03880(.A0(new_n6300_), .A1(new_n6023_), .B0(new_n6025_), .Y(new_n6317_));
  AOI21X1  g03881(.A0(new_n6317_), .A1(new_n6316_), .B0(new_n5879_), .Y(new_n6318_));
  OAI21X1  g03882(.A0(new_n6313_), .A1(new_n6311_), .B0(new_n6318_), .Y(new_n6319_));
  OAI21X1  g03883(.A0(new_n6298_), .A1(new_n5878_), .B0(new_n6319_), .Y(new_n6320_));
  NOR3X1   g03884(.A(new_n6298_), .B(new_n6053_), .C(pi0351), .Y(new_n6321_));
  AOI21X1  g03885(.A0(new_n6320_), .A1(new_n6052_), .B0(new_n6321_), .Y(new_n6322_));
  NOR3X1   g03886(.A(new_n6298_), .B(new_n6053_), .C(new_n6050_), .Y(new_n6323_));
  AOI21X1  g03887(.A0(new_n6320_), .A1(new_n6057_), .B0(new_n6323_), .Y(new_n6324_));
  MX2X1    g03888(.A(new_n6324_), .B(new_n6322_), .S0(new_n5866_), .Y(new_n6325_));
  MX2X1    g03889(.A(new_n6324_), .B(new_n6322_), .S0(pi0461), .Y(new_n6326_));
  MX2X1    g03890(.A(new_n6326_), .B(new_n6325_), .S0(new_n5865_), .Y(new_n6327_));
  MX2X1    g03891(.A(new_n6326_), .B(new_n6325_), .S0(pi0357), .Y(new_n6328_));
  MX2X1    g03892(.A(new_n6328_), .B(new_n6327_), .S0(new_n5864_), .Y(new_n6329_));
  NOR2X1   g03893(.A(new_n6329_), .B(new_n5863_), .Y(new_n6330_));
  INVX1    g03894(.A(new_n5863_), .Y(new_n6331_));
  MX2X1    g03895(.A(new_n6328_), .B(new_n6327_), .S0(pi0356), .Y(new_n6332_));
  OAI21X1  g03896(.A0(new_n6332_), .A1(new_n6331_), .B0(new_n6069_), .Y(new_n6333_));
  INVX1    g03897(.A(pi0590), .Y(new_n6334_));
  AOI21X1  g03898(.A0(new_n6305_), .A1(pi0591), .B0(new_n6334_), .Y(new_n6335_));
  OAI21X1  g03899(.A0(new_n6333_), .A1(new_n6330_), .B0(new_n6335_), .Y(new_n6336_));
  XOR2X1   g03900(.A(new_n6151_), .B(pi0375), .Y(new_n6337_));
  XOR2X1   g03901(.A(new_n6337_), .B(new_n6075_), .Y(new_n6338_));
  INVX1    g03902(.A(new_n6100_), .Y(new_n6339_));
  MX2X1    g03903(.A(new_n6305_), .B(new_n5991_), .S0(pi0592), .Y(new_n6340_));
  AND2X1   g03904(.A(new_n6340_), .B(new_n6339_), .Y(new_n6341_));
  NOR2X1   g03905(.A(new_n6299_), .B(new_n6339_), .Y(new_n6342_));
  OR3X1    g03906(.A(new_n6342_), .B(new_n6341_), .C(pi1199), .Y(new_n6343_));
  OAI21X1  g03907(.A0(new_n6305_), .A1(new_n6114_), .B0(new_n6115_), .Y(new_n6344_));
  OAI21X1  g03908(.A0(new_n6305_), .A1(new_n6101_), .B0(new_n6111_), .Y(new_n6345_));
  AOI21X1  g03909(.A0(new_n6345_), .A1(new_n6344_), .B0(new_n6339_), .Y(new_n6346_));
  OR3X1    g03910(.A(new_n6346_), .B(new_n6341_), .C(new_n6053_), .Y(new_n6347_));
  AND2X1   g03911(.A(new_n6347_), .B(new_n6343_), .Y(new_n6348_));
  MX2X1    g03912(.A(new_n6348_), .B(new_n6340_), .S0(pi1198), .Y(new_n6349_));
  MX2X1    g03913(.A(new_n6349_), .B(new_n6348_), .S0(new_n6079_), .Y(new_n6350_));
  MX2X1    g03914(.A(new_n6349_), .B(new_n6348_), .S0(pi0374), .Y(new_n6351_));
  MX2X1    g03915(.A(new_n6351_), .B(new_n6350_), .S0(pi0369), .Y(new_n6352_));
  MX2X1    g03916(.A(new_n6351_), .B(new_n6350_), .S0(new_n6078_), .Y(new_n6353_));
  MX2X1    g03917(.A(new_n6353_), .B(new_n6352_), .S0(new_n6077_), .Y(new_n6354_));
  MX2X1    g03918(.A(new_n6353_), .B(new_n6352_), .S0(pi0370), .Y(new_n6355_));
  MX2X1    g03919(.A(new_n6355_), .B(new_n6354_), .S0(new_n6076_), .Y(new_n6356_));
  OR2X1    g03920(.A(new_n6355_), .B(pi0371), .Y(new_n6357_));
  OAI21X1  g03921(.A0(new_n6354_), .A1(new_n6076_), .B0(new_n6357_), .Y(new_n6358_));
  AOI21X1  g03922(.A0(new_n6358_), .A1(new_n6338_), .B0(pi0591), .Y(new_n6359_));
  OAI21X1  g03923(.A0(new_n6356_), .A1(new_n6338_), .B0(new_n6359_), .Y(new_n6360_));
  XOR2X1   g03924(.A(new_n6227_), .B(new_n6159_), .Y(new_n6361_));
  XOR2X1   g03925(.A(new_n6361_), .B(pi0393), .Y(new_n6362_));
  AND2X1   g03926(.A(pi1196), .B(new_n6009_), .Y(new_n6363_));
  INVX1    g03927(.A(new_n6363_), .Y(new_n6364_));
  AND3X1   g03928(.A(new_n6258_), .B(new_n6182_), .C(new_n2702_), .Y(new_n6365_));
  AND3X1   g03929(.A(new_n6365_), .B(new_n6295_), .C(pi0567), .Y(new_n6366_));
  AND2X1   g03930(.A(new_n6244_), .B(new_n6202_), .Y(new_n6367_));
  AOI21X1  g03931(.A0(new_n6367_), .A1(new_n6366_), .B0(new_n6364_), .Y(new_n6368_));
  INVX1    g03932(.A(new_n6365_), .Y(new_n6369_));
  OAI21X1  g03933(.A0(new_n6369_), .A1(new_n6270_), .B0(pi0299), .Y(new_n6370_));
  AND3X1   g03934(.A(new_n6258_), .B(new_n6202_), .C(new_n2702_), .Y(new_n6371_));
  INVX1    g03935(.A(new_n6371_), .Y(new_n6372_));
  OAI21X1  g03936(.A0(new_n6372_), .A1(new_n6270_), .B0(pi0299), .Y(new_n6373_));
  AND2X1   g03937(.A(new_n6365_), .B(new_n6202_), .Y(new_n6374_));
  AND3X1   g03938(.A(new_n5947_), .B(new_n6255_), .C(pi1091), .Y(new_n6375_));
  OR3X1    g03939(.A(new_n6375_), .B(new_n6374_), .C(new_n5059_), .Y(new_n6376_));
  AND3X1   g03940(.A(new_n5947_), .B(new_n5044_), .C(pi1091), .Y(new_n6377_));
  NOR2X1   g03941(.A(new_n6377_), .B(new_n6374_), .Y(new_n6378_));
  AOI21X1  g03942(.A0(new_n6378_), .A1(new_n5059_), .B0(new_n6271_), .Y(new_n6379_));
  AOI22X1  g03943(.A0(new_n6379_), .A1(new_n6376_), .B0(new_n6373_), .B1(new_n6370_), .Y(new_n6380_));
  OAI21X1  g03944(.A0(new_n6369_), .A1(new_n6264_), .B0(new_n2933_), .Y(new_n6381_));
  OAI21X1  g03945(.A0(new_n6372_), .A1(new_n6264_), .B0(new_n2933_), .Y(new_n6382_));
  OR3X1    g03946(.A(new_n6375_), .B(new_n6374_), .C(new_n5042_), .Y(new_n6383_));
  AOI21X1  g03947(.A0(new_n6378_), .A1(new_n5042_), .B0(new_n6265_), .Y(new_n6384_));
  AOI22X1  g03948(.A0(new_n6384_), .A1(new_n6383_), .B0(new_n6382_), .B1(new_n6381_), .Y(new_n6385_));
  OR3X1    g03949(.A(new_n6385_), .B(new_n6380_), .C(new_n2939_), .Y(new_n6386_));
  OR3X1    g03950(.A(new_n6182_), .B(new_n5910_), .C(pi1091), .Y(new_n6387_));
  NAND2X1  g03951(.A(new_n6387_), .B(new_n6254_), .Y(new_n6388_));
  INVX1    g03952(.A(new_n6202_), .Y(new_n6389_));
  NOR3X1   g03953(.A(new_n6389_), .B(new_n5929_), .C(new_n5928_), .Y(new_n6390_));
  AOI21X1  g03954(.A0(new_n6244_), .A1(new_n6202_), .B0(pi0122), .Y(new_n6391_));
  NOR2X1   g03955(.A(new_n6391_), .B(new_n5032_), .Y(new_n6392_));
  OAI21X1  g03956(.A0(new_n6390_), .A1(new_n5906_), .B0(new_n6392_), .Y(new_n6393_));
  AND2X1   g03957(.A(new_n6393_), .B(new_n5944_), .Y(new_n6394_));
  OAI21X1  g03958(.A0(new_n6394_), .A1(new_n6388_), .B0(new_n6386_), .Y(new_n6395_));
  OAI21X1  g03959(.A0(new_n6369_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n6396_));
  OAI21X1  g03960(.A0(new_n6372_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n6397_));
  AOI22X1  g03961(.A0(new_n6397_), .A1(new_n6396_), .B0(new_n6395_), .B1(new_n2979_), .Y(new_n6398_));
  NAND2X1  g03962(.A(new_n6279_), .B(pi1091), .Y(new_n6399_));
  INVX1    g03963(.A(new_n6374_), .Y(new_n6400_));
  OAI22X1  g03964(.A0(new_n5919_), .A1(new_n5048_), .B0(new_n2961_), .B1(pi0299), .Y(new_n6401_));
  AOI21X1  g03965(.A0(new_n6400_), .A1(new_n2702_), .B0(new_n6401_), .Y(new_n6402_));
  AOI22X1  g03966(.A0(new_n6402_), .A1(new_n6399_), .B0(new_n5960_), .B1(new_n5918_), .Y(new_n6403_));
  OR2X1    g03967(.A(new_n6401_), .B(new_n2793_), .Y(new_n6404_));
  AOI21X1  g03968(.A0(new_n6404_), .A1(new_n6374_), .B0(new_n5215_), .Y(new_n6405_));
  OAI21X1  g03969(.A0(new_n6403_), .A1(new_n2793_), .B0(new_n6405_), .Y(new_n6406_));
  AOI21X1  g03970(.A0(new_n6365_), .A1(new_n6202_), .B0(pi0232), .Y(new_n6407_));
  AOI21X1  g03971(.A0(new_n6407_), .A1(new_n5961_), .B0(new_n3060_), .Y(new_n6408_));
  OAI21X1  g03972(.A0(new_n6400_), .A1(new_n3047_), .B0(pi0100), .Y(new_n6409_));
  AOI21X1  g03973(.A0(new_n6408_), .A1(new_n6406_), .B0(new_n6409_), .Y(new_n6410_));
  OAI21X1  g03974(.A0(new_n6410_), .A1(new_n6398_), .B0(new_n3131_), .Y(new_n6411_));
  AOI21X1  g03975(.A0(new_n6365_), .A1(new_n3132_), .B0(new_n3131_), .Y(new_n6412_));
  AOI21X1  g03976(.A0(new_n6371_), .A1(new_n3132_), .B0(new_n3131_), .Y(new_n6413_));
  NOR3X1   g03977(.A(new_n6182_), .B(new_n5913_), .C(pi1091), .Y(new_n6414_));
  INVX1    g03978(.A(new_n5985_), .Y(new_n6415_));
  OAI21X1  g03979(.A0(new_n6202_), .A1(new_n6415_), .B0(new_n6290_), .Y(new_n6416_));
  OAI22X1  g03980(.A0(new_n6416_), .A1(new_n6414_), .B0(new_n6413_), .B1(new_n6412_), .Y(new_n6417_));
  AOI21X1  g03981(.A0(new_n6417_), .A1(new_n6411_), .B0(pi0075), .Y(new_n6418_));
  OR2X1    g03982(.A(new_n6374_), .B(pi1091), .Y(new_n6419_));
  AOI21X1  g03983(.A0(new_n6365_), .A1(new_n6238_), .B0(new_n3073_), .Y(new_n6420_));
  INVX1    g03984(.A(new_n6420_), .Y(new_n6421_));
  OAI21X1  g03985(.A0(new_n6372_), .A1(new_n5921_), .B0(pi0075), .Y(new_n6422_));
  AOI22X1  g03986(.A0(new_n6422_), .A1(new_n6421_), .B0(new_n6419_), .B1(new_n6241_), .Y(new_n6423_));
  OAI21X1  g03987(.A0(new_n6423_), .A1(new_n6418_), .B0(new_n6368_), .Y(new_n6424_));
  AND3X1   g03988(.A(new_n6371_), .B(new_n6295_), .C(pi0567), .Y(new_n6425_));
  NOR2X1   g03989(.A(pi1196), .B(pi0592), .Y(new_n6426_));
  INVX1    g03990(.A(new_n6426_), .Y(new_n6427_));
  NOR2X1   g03991(.A(new_n6427_), .B(new_n6425_), .Y(new_n6428_));
  NAND2X1  g03992(.A(new_n6416_), .B(new_n6413_), .Y(new_n6429_));
  NOR3X1   g03993(.A(new_n6371_), .B(new_n5962_), .C(new_n3007_), .Y(new_n6430_));
  OR3X1    g03994(.A(new_n6377_), .B(new_n6371_), .C(new_n5058_), .Y(new_n6431_));
  OR3X1    g03995(.A(new_n6375_), .B(new_n6371_), .C(new_n5059_), .Y(new_n6432_));
  AND3X1   g03996(.A(new_n6432_), .B(new_n6431_), .C(new_n6270_), .Y(new_n6433_));
  NOR2X1   g03997(.A(new_n6433_), .B(new_n6373_), .Y(new_n6434_));
  OR3X1    g03998(.A(new_n6377_), .B(new_n6371_), .C(new_n5041_), .Y(new_n6435_));
  OR3X1    g03999(.A(new_n6375_), .B(new_n6371_), .C(new_n5042_), .Y(new_n6436_));
  AND3X1   g04000(.A(new_n6436_), .B(new_n6435_), .C(new_n6264_), .Y(new_n6437_));
  OAI21X1  g04001(.A0(new_n6437_), .A1(new_n6382_), .B0(pi0039), .Y(new_n6438_));
  OAI22X1  g04002(.A0(new_n6438_), .A1(new_n6434_), .B0(new_n6394_), .B1(new_n6250_), .Y(new_n6439_));
  AOI21X1  g04003(.A0(new_n6439_), .A1(new_n2979_), .B0(new_n6397_), .Y(new_n6440_));
  OAI21X1  g04004(.A0(new_n6440_), .A1(new_n6430_), .B0(new_n3131_), .Y(new_n6441_));
  AOI21X1  g04005(.A0(new_n6441_), .A1(new_n6429_), .B0(pi0075), .Y(new_n6442_));
  OAI21X1  g04006(.A0(new_n6280_), .A1(new_n6389_), .B0(new_n2702_), .Y(new_n6443_));
  AOI21X1  g04007(.A0(new_n6443_), .A1(new_n6241_), .B0(new_n6422_), .Y(new_n6444_));
  OAI21X1  g04008(.A0(new_n6444_), .A1(new_n6442_), .B0(new_n6428_), .Y(new_n6445_));
  AOI21X1  g04009(.A0(new_n6445_), .A1(new_n6424_), .B0(new_n5979_), .Y(new_n6446_));
  OR2X1    g04010(.A(new_n6428_), .B(new_n6368_), .Y(new_n6447_));
  AND2X1   g04011(.A(new_n6447_), .B(new_n5917_), .Y(new_n6448_));
  NOR3X1   g04012(.A(new_n6448_), .B(new_n6446_), .C(new_n6053_), .Y(new_n6449_));
  INVX1    g04013(.A(new_n6449_), .Y(new_n6450_));
  INVX1    g04014(.A(new_n6173_), .Y(new_n6451_));
  OR3X1    g04015(.A(new_n6377_), .B(new_n6365_), .C(new_n5058_), .Y(new_n6452_));
  NOR2X1   g04016(.A(new_n6375_), .B(new_n6365_), .Y(new_n6453_));
  AOI21X1  g04017(.A0(new_n6453_), .A1(new_n5058_), .B0(new_n6271_), .Y(new_n6454_));
  AOI21X1  g04018(.A0(new_n6454_), .A1(new_n6452_), .B0(new_n6370_), .Y(new_n6455_));
  OR3X1    g04019(.A(new_n6377_), .B(new_n6365_), .C(new_n5041_), .Y(new_n6456_));
  AOI21X1  g04020(.A0(new_n6453_), .A1(new_n5041_), .B0(new_n6265_), .Y(new_n6457_));
  AOI21X1  g04021(.A0(new_n6457_), .A1(new_n6456_), .B0(new_n6381_), .Y(new_n6458_));
  OR3X1    g04022(.A(new_n6458_), .B(new_n6455_), .C(new_n2939_), .Y(new_n6459_));
  AOI21X1  g04023(.A0(new_n6459_), .A1(new_n6388_), .B0(pi0038), .Y(new_n6460_));
  OAI22X1  g04024(.A0(new_n6460_), .A1(new_n6396_), .B0(new_n6365_), .B1(new_n5964_), .Y(new_n6461_));
  OAI21X1  g04025(.A0(new_n6182_), .A1(new_n6415_), .B0(new_n6290_), .Y(new_n6462_));
  AOI22X1  g04026(.A0(new_n6462_), .A1(new_n6412_), .B0(new_n6461_), .B1(new_n3131_), .Y(new_n6463_));
  AOI21X1  g04027(.A0(new_n6258_), .A1(new_n6182_), .B0(pi1091), .Y(new_n6464_));
  OAI21X1  g04028(.A0(new_n6464_), .A1(new_n6242_), .B0(new_n6420_), .Y(new_n6465_));
  OAI21X1  g04029(.A0(new_n6463_), .A1(pi0075), .B0(new_n6465_), .Y(new_n6466_));
  AOI21X1  g04030(.A0(new_n6466_), .A1(pi0567), .B0(new_n5917_), .Y(new_n6467_));
  NOR3X1   g04031(.A(new_n6467_), .B(new_n6366_), .C(new_n6364_), .Y(new_n6468_));
  OR3X1    g04032(.A(new_n6468_), .B(new_n6312_), .C(pi1199), .Y(new_n6469_));
  AND2X1   g04033(.A(new_n6469_), .B(new_n6451_), .Y(new_n6470_));
  AND2X1   g04034(.A(new_n5990_), .B(new_n6009_), .Y(new_n6471_));
  AOI21X1  g04035(.A0(new_n6173_), .A1(new_n6471_), .B0(new_n6297_), .Y(new_n6472_));
  INVX1    g04036(.A(new_n6472_), .Y(new_n6473_));
  AOI21X1  g04037(.A0(new_n6470_), .A1(new_n6450_), .B0(new_n6473_), .Y(new_n6474_));
  MX2X1    g04038(.A(new_n6474_), .B(new_n6298_), .S0(pi1197), .Y(new_n6475_));
  MX2X1    g04039(.A(new_n6475_), .B(new_n6474_), .S0(pi0333), .Y(new_n6476_));
  MX2X1    g04040(.A(new_n6475_), .B(new_n6474_), .S0(new_n6162_), .Y(new_n6477_));
  MX2X1    g04041(.A(new_n6477_), .B(new_n6476_), .S0(new_n6219_), .Y(new_n6478_));
  MX2X1    g04042(.A(new_n6477_), .B(new_n6476_), .S0(pi0391), .Y(new_n6479_));
  MX2X1    g04043(.A(new_n6479_), .B(new_n6478_), .S0(new_n6161_), .Y(new_n6480_));
  OR2X1    g04044(.A(new_n6480_), .B(new_n6362_), .Y(new_n6481_));
  OR2X1    g04045(.A(new_n6479_), .B(pi0392), .Y(new_n6482_));
  OAI21X1  g04046(.A0(new_n6478_), .A1(new_n6161_), .B0(new_n6482_), .Y(new_n6483_));
  AOI21X1  g04047(.A0(new_n6483_), .A1(new_n6362_), .B0(new_n6069_), .Y(new_n6484_));
  AOI21X1  g04048(.A0(new_n6484_), .A1(new_n6481_), .B0(pi0590), .Y(new_n6485_));
  AOI21X1  g04049(.A0(new_n6485_), .A1(new_n6360_), .B0(new_n6072_), .Y(new_n6486_));
  AOI21X1  g04050(.A0(new_n6486_), .A1(new_n6336_), .B0(pi0588), .Y(new_n6487_));
  OAI21X1  g04051(.A0(new_n6237_), .A1(new_n6071_), .B0(new_n6487_), .Y(new_n6488_));
  AND2X1   g04052(.A(new_n5102_), .B(new_n2436_), .Y(new_n6489_));
  INVX1    g04053(.A(new_n6489_), .Y(po1038));
  INVX1    g04054(.A(pi0448), .Y(new_n6491_));
  INVX1    g04055(.A(pi0449), .Y(new_n6492_));
  XOR2X1   g04056(.A(pi0451), .B(pi0433), .Y(new_n6493_));
  XOR2X1   g04057(.A(new_n6493_), .B(new_n6492_), .Y(new_n6494_));
  XOR2X1   g04058(.A(new_n6494_), .B(new_n6491_), .Y(new_n6495_));
  INVX1    g04059(.A(pi0427), .Y(new_n6496_));
  INVX1    g04060(.A(pi0428), .Y(new_n6497_));
  XOR2X1   g04061(.A(pi0418), .B(pi0417), .Y(new_n6498_));
  XOR2X1   g04062(.A(new_n6498_), .B(pi0437), .Y(new_n6499_));
  INVX1    g04063(.A(pi0453), .Y(new_n6500_));
  XOR2X1   g04064(.A(pi0464), .B(new_n6500_), .Y(new_n6501_));
  XOR2X1   g04065(.A(new_n6501_), .B(new_n6499_), .Y(new_n6502_));
  XOR2X1   g04066(.A(pi0431), .B(pi0415), .Y(new_n6503_));
  INVX1    g04067(.A(pi0416), .Y(new_n6504_));
  XOR2X1   g04068(.A(pi0438), .B(new_n6504_), .Y(new_n6505_));
  XOR2X1   g04069(.A(new_n6505_), .B(new_n6503_), .Y(new_n6506_));
  AND2X1   g04070(.A(new_n6506_), .B(new_n6502_), .Y(new_n6507_));
  OAI21X1  g04071(.A0(new_n6506_), .A1(new_n6502_), .B0(pi1197), .Y(new_n6508_));
  XOR2X1   g04072(.A(pi0454), .B(pi0421), .Y(new_n6509_));
  XOR2X1   g04073(.A(pi0459), .B(pi0432), .Y(new_n6510_));
  XOR2X1   g04074(.A(new_n6510_), .B(new_n6509_), .Y(new_n6511_));
  XOR2X1   g04075(.A(pi0420), .B(pi0419), .Y(new_n6512_));
  XOR2X1   g04076(.A(pi0424), .B(pi0423), .Y(new_n6513_));
  XOR2X1   g04077(.A(new_n6513_), .B(new_n6512_), .Y(new_n6514_));
  XOR2X1   g04078(.A(new_n6514_), .B(new_n6511_), .Y(new_n6515_));
  AND2X1   g04079(.A(new_n6515_), .B(pi0425), .Y(new_n6516_));
  OAI21X1  g04080(.A0(new_n6515_), .A1(pi0425), .B0(pi1198), .Y(new_n6517_));
  OAI22X1  g04081(.A0(new_n6517_), .A1(new_n6516_), .B0(new_n6508_), .B1(new_n6507_), .Y(new_n6518_));
  NOR2X1   g04082(.A(new_n5978_), .B(pi1196), .Y(new_n6519_));
  INVX1    g04083(.A(pi0444), .Y(new_n6520_));
  NOR2X1   g04084(.A(pi0592), .B(pi0443), .Y(new_n6521_));
  MX2X1    g04085(.A(new_n5978_), .B(new_n5991_), .S0(new_n6521_), .Y(new_n6522_));
  AND2X1   g04086(.A(new_n6009_), .B(pi0443), .Y(new_n6523_));
  MX2X1    g04087(.A(new_n5978_), .B(new_n5991_), .S0(new_n6523_), .Y(new_n6524_));
  MX2X1    g04088(.A(new_n6524_), .B(new_n6522_), .S0(new_n6520_), .Y(new_n6525_));
  NOR2X1   g04089(.A(new_n6525_), .B(pi0436), .Y(new_n6526_));
  INVX1    g04090(.A(pi0436), .Y(new_n6527_));
  XOR2X1   g04091(.A(pi0435), .B(pi0429), .Y(new_n6528_));
  XOR2X1   g04092(.A(pi0446), .B(pi0434), .Y(new_n6529_));
  INVX1    g04093(.A(pi0414), .Y(new_n6530_));
  XOR2X1   g04094(.A(pi0422), .B(new_n6530_), .Y(new_n6531_));
  XOR2X1   g04095(.A(new_n6531_), .B(new_n6529_), .Y(new_n6532_));
  INVX1    g04096(.A(new_n6532_), .Y(new_n6533_));
  XOR2X1   g04097(.A(new_n6533_), .B(new_n6528_), .Y(new_n6534_));
  MX2X1    g04098(.A(new_n6524_), .B(new_n6522_), .S0(pi0444), .Y(new_n6535_));
  OAI21X1  g04099(.A0(new_n6535_), .A1(new_n6527_), .B0(new_n6534_), .Y(new_n6536_));
  NOR2X1   g04100(.A(new_n6536_), .B(new_n6526_), .Y(new_n6537_));
  INVX1    g04101(.A(new_n6534_), .Y(new_n6538_));
  OR2X1    g04102(.A(new_n6535_), .B(pi0436), .Y(new_n6539_));
  OR2X1    g04103(.A(new_n6525_), .B(new_n6527_), .Y(new_n6540_));
  AND3X1   g04104(.A(new_n6540_), .B(new_n6539_), .C(new_n6538_), .Y(new_n6541_));
  NOR3X1   g04105(.A(new_n6541_), .B(new_n6537_), .C(new_n6045_), .Y(new_n6542_));
  NOR3X1   g04106(.A(new_n6542_), .B(new_n6518_), .C(new_n6519_), .Y(new_n6543_));
  AOI21X1  g04107(.A0(new_n6518_), .A1(new_n5992_), .B0(new_n6543_), .Y(new_n6544_));
  MX2X1    g04108(.A(new_n6544_), .B(new_n5993_), .S0(new_n6497_), .Y(new_n6545_));
  MX2X1    g04109(.A(new_n6544_), .B(new_n5993_), .S0(pi0428), .Y(new_n6546_));
  MX2X1    g04110(.A(new_n6546_), .B(new_n6545_), .S0(new_n6496_), .Y(new_n6547_));
  MX2X1    g04111(.A(new_n6546_), .B(new_n6545_), .S0(pi0427), .Y(new_n6548_));
  MX2X1    g04112(.A(new_n6548_), .B(new_n6547_), .S0(pi0430), .Y(new_n6549_));
  INVX1    g04113(.A(pi0430), .Y(new_n6550_));
  MX2X1    g04114(.A(new_n6548_), .B(new_n6547_), .S0(new_n6550_), .Y(new_n6551_));
  MX2X1    g04115(.A(new_n6551_), .B(new_n6549_), .S0(pi0426), .Y(new_n6552_));
  INVX1    g04116(.A(pi0426), .Y(new_n6553_));
  MX2X1    g04117(.A(new_n6551_), .B(new_n6549_), .S0(new_n6553_), .Y(new_n6554_));
  MX2X1    g04118(.A(new_n6554_), .B(new_n6552_), .S0(pi0445), .Y(new_n6555_));
  OR2X1    g04119(.A(new_n6555_), .B(new_n6495_), .Y(new_n6556_));
  INVX1    g04120(.A(pi0445), .Y(new_n6557_));
  OR2X1    g04121(.A(new_n6554_), .B(new_n6557_), .Y(new_n6558_));
  OAI21X1  g04122(.A0(new_n6552_), .A1(pi0445), .B0(new_n6558_), .Y(new_n6559_));
  AOI21X1  g04123(.A0(new_n6559_), .A1(new_n6495_), .B0(new_n6053_), .Y(new_n6560_));
  NOR2X1   g04124(.A(pi0591), .B(pi0590), .Y(new_n6561_));
  INVX1    g04125(.A(new_n6561_), .Y(new_n6562_));
  AND2X1   g04126(.A(new_n6544_), .B(new_n6053_), .Y(new_n6563_));
  OR2X1    g04127(.A(new_n6563_), .B(new_n6562_), .Y(new_n6564_));
  AOI21X1  g04128(.A0(new_n6560_), .A1(new_n6556_), .B0(new_n6564_), .Y(new_n6565_));
  OAI21X1  g04129(.A0(new_n6561_), .A1(new_n5994_), .B0(new_n6072_), .Y(new_n6566_));
  XOR2X1   g04130(.A(pi0444), .B(new_n6527_), .Y(new_n6567_));
  XOR2X1   g04131(.A(new_n6567_), .B(new_n6538_), .Y(new_n6568_));
  INVX1    g04132(.A(new_n6568_), .Y(new_n6569_));
  AOI21X1  g04133(.A0(new_n6521_), .A1(new_n5990_), .B0(new_n6569_), .Y(new_n6570_));
  OAI21X1  g04134(.A0(new_n6521_), .A1(new_n6305_), .B0(new_n6570_), .Y(new_n6571_));
  OR3X1    g04135(.A(new_n6523_), .B(new_n6296_), .C(new_n6294_), .Y(new_n6572_));
  AOI21X1  g04136(.A0(new_n6523_), .A1(new_n5990_), .B0(new_n6568_), .Y(new_n6573_));
  AOI21X1  g04137(.A0(new_n6573_), .A1(new_n6572_), .B0(new_n6045_), .Y(new_n6574_));
  AOI21X1  g04138(.A0(new_n6574_), .A1(new_n6571_), .B0(new_n6312_), .Y(new_n6575_));
  MX2X1    g04139(.A(new_n6575_), .B(new_n6298_), .S0(new_n6518_), .Y(new_n6576_));
  OAI21X1  g04140(.A0(new_n6300_), .A1(pi0428), .B0(pi0427), .Y(new_n6577_));
  AOI21X1  g04141(.A0(new_n6576_), .A1(pi0428), .B0(new_n6577_), .Y(new_n6578_));
  OAI21X1  g04142(.A0(new_n6300_), .A1(new_n6497_), .B0(new_n6496_), .Y(new_n6579_));
  AOI21X1  g04143(.A0(new_n6576_), .A1(new_n6497_), .B0(new_n6579_), .Y(new_n6580_));
  OAI21X1  g04144(.A0(new_n6580_), .A1(new_n6578_), .B0(new_n6550_), .Y(new_n6581_));
  XOR2X1   g04145(.A(pi0428), .B(new_n6496_), .Y(new_n6582_));
  MX2X1    g04146(.A(new_n6576_), .B(new_n6298_), .S0(new_n6582_), .Y(new_n6583_));
  OAI21X1  g04147(.A0(new_n6583_), .A1(new_n6550_), .B0(new_n6581_), .Y(new_n6584_));
  OAI21X1  g04148(.A0(new_n6580_), .A1(new_n6578_), .B0(pi0430), .Y(new_n6585_));
  OAI21X1  g04149(.A0(new_n6583_), .A1(pi0430), .B0(new_n6585_), .Y(new_n6586_));
  MX2X1    g04150(.A(new_n6586_), .B(new_n6584_), .S0(new_n6553_), .Y(new_n6587_));
  AND2X1   g04151(.A(new_n6587_), .B(new_n6557_), .Y(new_n6588_));
  MX2X1    g04152(.A(new_n6586_), .B(new_n6584_), .S0(pi0426), .Y(new_n6589_));
  AOI21X1  g04153(.A0(new_n6589_), .A1(pi0445), .B0(new_n6588_), .Y(new_n6590_));
  INVX1    g04154(.A(new_n6494_), .Y(new_n6591_));
  MX2X1    g04155(.A(new_n6589_), .B(new_n6587_), .S0(pi0445), .Y(new_n6592_));
  OAI21X1  g04156(.A0(new_n6592_), .A1(pi0448), .B0(new_n6591_), .Y(new_n6593_));
  AOI21X1  g04157(.A0(new_n6590_), .A1(pi0448), .B0(new_n6593_), .Y(new_n6594_));
  OAI21X1  g04158(.A0(new_n6592_), .A1(new_n6491_), .B0(new_n6494_), .Y(new_n6595_));
  AOI21X1  g04159(.A0(new_n6590_), .A1(new_n6491_), .B0(new_n6595_), .Y(new_n6596_));
  OR2X1    g04160(.A(new_n6596_), .B(new_n6594_), .Y(new_n6597_));
  OAI21X1  g04161(.A0(new_n6576_), .A1(pi1199), .B0(new_n6561_), .Y(new_n6598_));
  AOI21X1  g04162(.A0(new_n6597_), .A1(pi1199), .B0(new_n6598_), .Y(new_n6599_));
  OAI21X1  g04163(.A0(new_n6561_), .A1(new_n6299_), .B0(new_n6073_), .Y(new_n6600_));
  OAI22X1  g04164(.A0(new_n6600_), .A1(new_n6599_), .B0(new_n6566_), .B1(new_n6565_), .Y(new_n6601_));
  AOI21X1  g04165(.A0(new_n6601_), .A1(pi0588), .B0(po1038), .Y(new_n6602_));
  INVX1    g04166(.A(pi0588), .Y(new_n6603_));
  AND2X1   g04167(.A(new_n6247_), .B(pi0567), .Y(new_n6604_));
  INVX1    g04168(.A(new_n6604_), .Y(new_n6605_));
  AND2X1   g04169(.A(new_n6022_), .B(new_n6009_), .Y(new_n6606_));
  NOR3X1   g04170(.A(new_n6606_), .B(new_n6605_), .C(new_n6017_), .Y(new_n6607_));
  INVX1    g04171(.A(new_n6607_), .Y(new_n6608_));
  INVX1    g04172(.A(pi0441), .Y(new_n6609_));
  XOR2X1   g04173(.A(pi0458), .B(new_n6018_), .Y(new_n6610_));
  XOR2X1   g04174(.A(new_n6610_), .B(new_n6015_), .Y(new_n6611_));
  AND2X1   g04175(.A(new_n6611_), .B(new_n6609_), .Y(new_n6612_));
  NOR2X1   g04176(.A(new_n6611_), .B(new_n6609_), .Y(new_n6613_));
  OR3X1    g04177(.A(new_n6613_), .B(new_n6612_), .C(pi0592), .Y(new_n6614_));
  AND3X1   g04178(.A(new_n6247_), .B(new_n6017_), .C(pi0567), .Y(new_n6615_));
  AOI21X1  g04179(.A0(new_n6615_), .A1(new_n6614_), .B0(new_n6045_), .Y(new_n6616_));
  AOI21X1  g04180(.A0(new_n6616_), .A1(new_n6608_), .B0(pi1198), .Y(new_n6617_));
  INVX1    g04181(.A(new_n6617_), .Y(new_n6618_));
  XOR2X1   g04182(.A(new_n6004_), .B(new_n6007_), .Y(new_n6619_));
  INVX1    g04183(.A(new_n6619_), .Y(new_n6620_));
  NAND3X1  g04184(.A(new_n6247_), .B(new_n6009_), .C(pi0567), .Y(new_n6621_));
  OR4X1    g04185(.A(new_n6621_), .B(new_n6620_), .C(new_n6023_), .D(new_n6025_), .Y(new_n6622_));
  AOI21X1  g04186(.A0(new_n6622_), .A1(new_n6618_), .B0(new_n5879_), .Y(new_n6623_));
  INVX1    g04187(.A(new_n6623_), .Y(new_n6624_));
  AOI21X1  g04188(.A0(new_n6624_), .A1(new_n6009_), .B0(new_n6605_), .Y(new_n6625_));
  INVX1    g04189(.A(new_n6625_), .Y(new_n6626_));
  AND3X1   g04190(.A(new_n6247_), .B(pi0592), .C(pi0567), .Y(new_n6627_));
  NOR2X1   g04191(.A(new_n6627_), .B(new_n6053_), .Y(new_n6628_));
  AOI22X1  g04192(.A0(new_n6628_), .A1(pi0351), .B0(new_n6626_), .B1(new_n6057_), .Y(new_n6629_));
  AOI22X1  g04193(.A0(new_n6628_), .A1(new_n6050_), .B0(new_n6626_), .B1(new_n6052_), .Y(new_n6630_));
  MX2X1    g04194(.A(new_n6630_), .B(new_n6629_), .S0(new_n5866_), .Y(new_n6631_));
  MX2X1    g04195(.A(new_n6630_), .B(new_n6629_), .S0(pi0461), .Y(new_n6632_));
  MX2X1    g04196(.A(new_n6632_), .B(new_n6631_), .S0(new_n5865_), .Y(new_n6633_));
  OR2X1    g04197(.A(new_n6633_), .B(pi0356), .Y(new_n6634_));
  MX2X1    g04198(.A(new_n6632_), .B(new_n6631_), .S0(pi0357), .Y(new_n6635_));
  OR2X1    g04199(.A(new_n6635_), .B(new_n5864_), .Y(new_n6636_));
  NAND3X1  g04200(.A(new_n6636_), .B(new_n6634_), .C(new_n5863_), .Y(new_n6637_));
  OR2X1    g04201(.A(new_n6635_), .B(pi0356), .Y(new_n6638_));
  OR2X1    g04202(.A(new_n6633_), .B(new_n5864_), .Y(new_n6639_));
  NAND3X1  g04203(.A(new_n6639_), .B(new_n6638_), .C(new_n6331_), .Y(new_n6640_));
  AOI21X1  g04204(.A0(new_n6640_), .A1(new_n6637_), .B0(new_n6334_), .Y(new_n6641_));
  XOR2X1   g04205(.A(new_n6109_), .B(new_n6113_), .Y(new_n6642_));
  NOR3X1   g04206(.A(new_n6642_), .B(new_n6099_), .C(new_n6088_), .Y(new_n6643_));
  OAI21X1  g04207(.A0(new_n6643_), .A1(new_n6009_), .B0(new_n6604_), .Y(new_n6644_));
  AOI22X1  g04208(.A0(new_n6644_), .A1(pi1199), .B0(new_n6339_), .B1(pi0592), .Y(new_n6645_));
  NAND3X1  g04209(.A(new_n6645_), .B(new_n6627_), .C(new_n6025_), .Y(new_n6646_));
  XOR2X1   g04210(.A(pi0374), .B(pi0369), .Y(new_n6647_));
  XOR2X1   g04211(.A(new_n6647_), .B(pi0370), .Y(new_n6648_));
  XOR2X1   g04212(.A(new_n6648_), .B(pi0371), .Y(new_n6649_));
  XOR2X1   g04213(.A(new_n6649_), .B(pi0373), .Y(new_n6650_));
  XOR2X1   g04214(.A(new_n6650_), .B(new_n6074_), .Y(new_n6651_));
  XOR2X1   g04215(.A(new_n6651_), .B(new_n6151_), .Y(new_n6652_));
  NAND3X1  g04216(.A(new_n6652_), .B(new_n6645_), .C(new_n6627_), .Y(new_n6653_));
  AND3X1   g04217(.A(new_n6653_), .B(new_n6646_), .C(new_n6621_), .Y(new_n6654_));
  OAI21X1  g04218(.A0(new_n6654_), .A1(pi0590), .B0(new_n6069_), .Y(new_n6655_));
  OAI21X1  g04219(.A0(new_n6182_), .A1(new_n6045_), .B0(new_n6009_), .Y(new_n6656_));
  NOR3X1   g04220(.A(new_n6656_), .B(new_n6372_), .C(new_n5979_), .Y(new_n6657_));
  OR3X1    g04221(.A(new_n6657_), .B(new_n6627_), .C(new_n6053_), .Y(new_n6658_));
  NAND4X1  g04222(.A(new_n6258_), .B(new_n6182_), .C(new_n2702_), .D(pi0567), .Y(new_n6659_));
  AOI21X1  g04223(.A0(new_n6364_), .A1(new_n6604_), .B0(pi1199), .Y(new_n6660_));
  OAI21X1  g04224(.A0(new_n6659_), .A1(new_n6364_), .B0(new_n6660_), .Y(new_n6661_));
  AND2X1   g04225(.A(new_n6661_), .B(new_n6658_), .Y(new_n6662_));
  MX2X1    g04226(.A(new_n6662_), .B(new_n6627_), .S0(pi1197), .Y(new_n6663_));
  INVX1    g04227(.A(new_n6662_), .Y(new_n6664_));
  NOR2X1   g04228(.A(new_n6627_), .B(new_n6025_), .Y(new_n6665_));
  INVX1    g04229(.A(new_n6665_), .Y(new_n6666_));
  NAND3X1  g04230(.A(new_n6666_), .B(new_n6661_), .C(new_n6658_), .Y(new_n6667_));
  AND2X1   g04231(.A(new_n6667_), .B(new_n6172_), .Y(new_n6668_));
  AOI21X1  g04232(.A0(new_n6664_), .A1(new_n6162_), .B0(new_n6668_), .Y(new_n6669_));
  OAI21X1  g04233(.A0(new_n6663_), .A1(new_n6162_), .B0(new_n6669_), .Y(new_n6670_));
  NOR2X1   g04234(.A(new_n6663_), .B(pi0333), .Y(new_n6671_));
  OR3X1    g04235(.A(new_n6671_), .B(new_n6668_), .C(new_n6664_), .Y(new_n6672_));
  MX2X1    g04236(.A(new_n6672_), .B(new_n6670_), .S0(new_n6219_), .Y(new_n6673_));
  MX2X1    g04237(.A(new_n6672_), .B(new_n6670_), .S0(pi0391), .Y(new_n6674_));
  MX2X1    g04238(.A(new_n6674_), .B(new_n6673_), .S0(new_n6161_), .Y(new_n6675_));
  NAND2X1  g04239(.A(new_n6675_), .B(new_n6160_), .Y(new_n6676_));
  INVX1    g04240(.A(new_n6361_), .Y(new_n6677_));
  MX2X1    g04241(.A(new_n6674_), .B(new_n6673_), .S0(pi0392), .Y(new_n6678_));
  AOI21X1  g04242(.A0(new_n6678_), .A1(pi0393), .B0(new_n6677_), .Y(new_n6679_));
  NAND2X1  g04243(.A(new_n6678_), .B(new_n6160_), .Y(new_n6680_));
  AOI21X1  g04244(.A0(new_n6675_), .A1(pi0393), .B0(new_n6361_), .Y(new_n6681_));
  AOI22X1  g04245(.A0(new_n6681_), .A1(new_n6680_), .B0(new_n6679_), .B1(new_n6676_), .Y(new_n6682_));
  AOI21X1  g04246(.A0(new_n6604_), .A1(pi0590), .B0(new_n6069_), .Y(new_n6683_));
  OAI21X1  g04247(.A0(new_n6682_), .A1(pi0590), .B0(new_n6683_), .Y(new_n6684_));
  OAI21X1  g04248(.A0(new_n6655_), .A1(new_n6641_), .B0(new_n6684_), .Y(new_n6685_));
  AOI21X1  g04249(.A0(new_n5102_), .A1(new_n2436_), .B0(new_n6072_), .Y(new_n6686_));
  XOR2X1   g04250(.A(pi0443), .B(pi0436), .Y(new_n6687_));
  XOR2X1   g04251(.A(new_n6687_), .B(new_n6520_), .Y(new_n6688_));
  OAI21X1  g04252(.A0(new_n6688_), .A1(new_n6538_), .B0(new_n6363_), .Y(new_n6689_));
  AOI21X1  g04253(.A0(new_n6688_), .A1(new_n6538_), .B0(new_n6689_), .Y(new_n6690_));
  NOR3X1   g04254(.A(new_n6690_), .B(new_n6621_), .C(new_n6518_), .Y(new_n6691_));
  XOR2X1   g04255(.A(new_n6582_), .B(new_n6550_), .Y(new_n6692_));
  XOR2X1   g04256(.A(new_n6692_), .B(pi0426), .Y(new_n6693_));
  XOR2X1   g04257(.A(new_n6693_), .B(pi0445), .Y(new_n6694_));
  XOR2X1   g04258(.A(new_n6694_), .B(new_n6491_), .Y(new_n6695_));
  AOI21X1  g04259(.A0(new_n6695_), .A1(new_n6691_), .B0(new_n6627_), .Y(new_n6696_));
  OR2X1    g04260(.A(new_n6696_), .B(new_n6591_), .Y(new_n6697_));
  NOR4X1   g04261(.A(new_n6695_), .B(new_n6690_), .C(new_n6621_), .D(new_n6518_), .Y(new_n6698_));
  OAI21X1  g04262(.A0(new_n6698_), .A1(new_n6627_), .B0(new_n6591_), .Y(new_n6699_));
  AND2X1   g04263(.A(new_n6699_), .B(pi1199), .Y(new_n6700_));
  OR2X1    g04264(.A(new_n6627_), .B(pi1199), .Y(new_n6701_));
  OAI21X1  g04265(.A0(new_n6701_), .A1(new_n6691_), .B0(new_n6561_), .Y(new_n6702_));
  AOI21X1  g04266(.A0(new_n6700_), .A1(new_n6697_), .B0(new_n6702_), .Y(new_n6703_));
  OAI21X1  g04267(.A0(new_n6561_), .A1(new_n6605_), .B0(pi0588), .Y(new_n6704_));
  OAI21X1  g04268(.A0(new_n6704_), .A1(new_n6703_), .B0(new_n6686_), .Y(new_n6705_));
  AOI21X1  g04269(.A0(new_n6685_), .A1(new_n6603_), .B0(new_n6705_), .Y(new_n6706_));
  OR2X1    g04270(.A(new_n6706_), .B(pi0217), .Y(new_n6707_));
  AOI21X1  g04271(.A0(new_n6602_), .A1(new_n6488_), .B0(new_n6707_), .Y(new_n6708_));
  OAI21X1  g04272(.A0(new_n6305_), .A1(new_n6072_), .B0(new_n6489_), .Y(new_n6709_));
  AOI21X1  g04273(.A0(new_n6072_), .A1(new_n5994_), .B0(new_n6709_), .Y(new_n6710_));
  INVX1    g04274(.A(new_n6686_), .Y(new_n6711_));
  OAI21X1  g04275(.A0(new_n6711_), .A1(new_n6605_), .B0(pi0217), .Y(new_n6712_));
  NOR3X1   g04276(.A(pi1163), .B(pi1162), .C(pi1161), .Y(new_n6713_));
  OAI21X1  g04277(.A0(new_n6712_), .A1(new_n6710_), .B0(new_n6713_), .Y(new_n6714_));
  INVX1    g04278(.A(pi1162), .Y(new_n6715_));
  INVX1    g04279(.A(pi1163), .Y(new_n6716_));
  NAND3X1  g04280(.A(new_n2720_), .B(new_n6716_), .C(pi1161), .Y(new_n6717_));
  OR3X1    g04281(.A(new_n6717_), .B(new_n6715_), .C(pi0031), .Y(new_n6718_));
  OAI21X1  g04282(.A0(new_n6714_), .A1(new_n6708_), .B0(new_n6718_), .Y(po0189));
  NOR4X1   g04283(.A(pi0062), .B(pi0059), .C(pi0057), .D(pi0056), .Y(new_n6720_));
  AND3X1   g04284(.A(new_n6720_), .B(new_n4982_), .C(new_n3107_), .Y(new_n6721_));
  AND3X1   g04285(.A(new_n6721_), .B(new_n3079_), .C(new_n3091_), .Y(new_n6722_));
  AND2X1   g04286(.A(new_n3047_), .B(pi0100), .Y(new_n6723_));
  INVX1    g04287(.A(new_n5082_), .Y(po1057));
  OR4X1    g04288(.A(new_n5086_), .B(po1057), .C(new_n5071_), .D(new_n2986_), .Y(new_n6725_));
  NOR3X1   g04289(.A(new_n2985_), .B(new_n2536_), .C(new_n5083_), .Y(new_n6726_));
  INVX1    g04290(.A(new_n6726_), .Y(new_n6727_));
  NOR2X1   g04291(.A(new_n5920_), .B(new_n5082_), .Y(new_n6728_));
  OR4X1    g04292(.A(new_n6728_), .B(new_n5072_), .C(new_n3035_), .D(pi0137), .Y(new_n6729_));
  OAI22X1  g04293(.A0(new_n6729_), .A1(new_n6727_), .B0(new_n6725_), .B1(pi0137), .Y(new_n6730_));
  OR2X1    g04294(.A(pi0090), .B(pi0024), .Y(new_n6731_));
  OR4X1    g04295(.A(new_n6731_), .B(new_n2526_), .C(pi0040), .D(pi0035), .Y(new_n6732_));
  NOR2X1   g04296(.A(pi0060), .B(pi0053), .Y(new_n6733_));
  INVX1    g04297(.A(pi0050), .Y(new_n6734_));
  NOR4X1   g04298(.A(new_n2567_), .B(new_n2558_), .C(pi0077), .D(new_n6734_), .Y(new_n6735_));
  NAND3X1  g04299(.A(new_n6735_), .B(new_n6733_), .C(new_n2566_), .Y(new_n6736_));
  NOR4X1   g04300(.A(new_n2495_), .B(new_n2475_), .C(new_n2473_), .D(pi0094), .Y(new_n6737_));
  INVX1    g04301(.A(new_n6737_), .Y(new_n6738_));
  OR4X1    g04302(.A(new_n6738_), .B(new_n6736_), .C(new_n6732_), .D(pi0093), .Y(new_n6739_));
  AND3X1   g04303(.A(new_n5225_), .B(new_n5032_), .C(pi0829), .Y(new_n6740_));
  AOI21X1  g04304(.A0(new_n2721_), .A1(new_n2703_), .B0(new_n6740_), .Y(new_n6741_));
  AOI21X1  g04305(.A0(new_n6741_), .A1(new_n6073_), .B0(pi0137), .Y(new_n6742_));
  NOR4X1   g04306(.A(pi0073), .B(pi0068), .C(pi0066), .D(pi0049), .Y(new_n6743_));
  NAND4X1  g04307(.A(new_n6743_), .B(new_n5122_), .C(new_n2603_), .D(pi0076), .Y(new_n6744_));
  OR4X1    g04308(.A(pi0102), .B(pi0089), .C(pi0077), .D(pi0050), .Y(new_n6745_));
  OR4X1    g04309(.A(pi0107), .B(pi0081), .C(pi0064), .D(pi0063), .Y(new_n6746_));
  OR2X1    g04310(.A(new_n6746_), .B(new_n6745_), .Y(new_n6747_));
  OR4X1    g04311(.A(pi0098), .B(pi0088), .C(pi0067), .D(pi0036), .Y(new_n6748_));
  OR3X1    g04312(.A(new_n6748_), .B(new_n2612_), .C(pi0103), .Y(new_n6749_));
  OR4X1    g04313(.A(pi0083), .B(pi0071), .C(pi0069), .D(pi0065), .Y(new_n6750_));
  OR2X1    g04314(.A(pi0048), .B(pi0045), .Y(new_n6751_));
  OR4X1    g04315(.A(new_n6751_), .B(new_n6750_), .C(pi0104), .D(pi0061), .Y(new_n6752_));
  NOR4X1   g04316(.A(new_n6752_), .B(new_n6749_), .C(new_n6747_), .D(new_n6744_), .Y(new_n6753_));
  NOR2X1   g04317(.A(new_n2476_), .B(new_n2474_), .Y(new_n6754_));
  OAI21X1  g04318(.A0(new_n6753_), .A1(new_n6735_), .B0(new_n6754_), .Y(new_n6755_));
  AND2X1   g04319(.A(new_n6755_), .B(new_n5777_), .Y(new_n6756_));
  OR4X1    g04320(.A(new_n6752_), .B(new_n6749_), .C(new_n6747_), .D(new_n6744_), .Y(new_n6757_));
  NOR3X1   g04321(.A(new_n6757_), .B(new_n6738_), .C(new_n2472_), .Y(new_n6758_));
  AND3X1   g04322(.A(new_n2746_), .B(new_n2535_), .C(new_n2534_), .Y(new_n6759_));
  NAND3X1  g04323(.A(new_n6759_), .B(new_n5897_), .C(new_n2452_), .Y(new_n6760_));
  AOI21X1  g04324(.A0(new_n6741_), .A1(new_n6073_), .B0(new_n6760_), .Y(new_n6761_));
  OAI21X1  g04325(.A0(new_n6758_), .A1(new_n5777_), .B0(new_n6761_), .Y(new_n6762_));
  OAI22X1  g04326(.A0(new_n6762_), .A1(new_n6756_), .B0(new_n6742_), .B1(new_n6739_), .Y(new_n6763_));
  AOI21X1  g04327(.A0(new_n2705_), .A1(new_n5777_), .B0(new_n2455_), .Y(new_n6764_));
  AOI22X1  g04328(.A0(new_n6764_), .A1(new_n2480_), .B0(new_n6763_), .B1(new_n2455_), .Y(new_n6765_));
  AND2X1   g04329(.A(new_n6739_), .B(new_n2455_), .Y(new_n6766_));
  OAI21X1  g04330(.A0(new_n5011_), .A1(new_n2455_), .B0(new_n5009_), .Y(new_n6767_));
  OAI22X1  g04331(.A0(new_n6767_), .A1(new_n6766_), .B0(new_n6765_), .B1(new_n5009_), .Y(new_n6768_));
  NOR4X1   g04332(.A(pi0100), .B(pi0095), .C(pi0039), .D(pi0038), .Y(new_n6769_));
  AOI22X1  g04333(.A0(new_n6769_), .A1(new_n6768_), .B0(new_n6730_), .B1(new_n6723_), .Y(new_n6770_));
  INVX1    g04334(.A(new_n6741_), .Y(po0840));
  OR4X1    g04335(.A(new_n2525_), .B(new_n2505_), .C(new_n2502_), .D(pi0024), .Y(new_n6772_));
  NAND3X1  g04336(.A(new_n2984_), .B(new_n2513_), .C(new_n2535_), .Y(new_n6773_));
  OR4X1    g04337(.A(new_n6773_), .B(new_n6772_), .C(po0840), .D(pi0051), .Y(new_n6774_));
  NOR2X1   g04338(.A(new_n5082_), .B(new_n5071_), .Y(new_n6775_));
  NOR2X1   g04339(.A(new_n6728_), .B(new_n3035_), .Y(new_n6776_));
  NOR3X1   g04340(.A(pi0087), .B(pi0039), .C(pi0038), .Y(new_n6777_));
  AND3X1   g04341(.A(new_n6777_), .B(new_n3007_), .C(pi0075), .Y(new_n6778_));
  INVX1    g04342(.A(new_n6778_), .Y(new_n6779_));
  OR4X1    g04343(.A(new_n6779_), .B(new_n6776_), .C(new_n6775_), .D(pi0137), .Y(new_n6780_));
  OAI22X1  g04344(.A0(new_n6780_), .A1(new_n6774_), .B0(new_n6770_), .B1(new_n3080_), .Y(new_n6781_));
  AND2X1   g04345(.A(new_n6781_), .B(new_n6722_), .Y(po0190));
  INVX1    g04346(.A(pi0034), .Y(new_n6783_));
  INVX1    g04347(.A(pi0079), .Y(new_n6784_));
  INVX1    g04348(.A(pi0118), .Y(new_n6785_));
  NOR4X1   g04349(.A(pi0196), .B(pi0195), .C(pi0139), .D(pi0138), .Y(new_n6786_));
  AND3X1   g04350(.A(new_n6786_), .B(new_n6785_), .C(new_n6784_), .Y(new_n6787_));
  AND2X1   g04351(.A(new_n6787_), .B(new_n6783_), .Y(new_n6788_));
  NOR2X1   g04352(.A(pi0157), .B(pi0149), .Y(new_n6789_));
  NOR3X1   g04353(.A(new_n6789_), .B(pi0468), .C(pi0332), .Y(new_n6790_));
  INVX1    g04354(.A(new_n6790_), .Y(new_n6791_));
  AOI21X1  g04355(.A0(pi0157), .A1(pi0149), .B0(new_n6791_), .Y(new_n6792_));
  AOI22X1  g04356(.A0(new_n6792_), .A1(pi0232), .B0(new_n3007_), .B1(new_n3073_), .Y(new_n6793_));
  NOR2X1   g04357(.A(pi0100), .B(pi0075), .Y(new_n6794_));
  AND3X1   g04358(.A(new_n6794_), .B(new_n5023_), .C(pi0232), .Y(new_n6795_));
  AOI21X1  g04359(.A0(new_n6795_), .A1(pi0164), .B0(new_n6793_), .Y(new_n6796_));
  OR2X1    g04360(.A(new_n6796_), .B(pi0074), .Y(new_n6797_));
  AND2X1   g04361(.A(new_n6795_), .B(pi0169), .Y(new_n6798_));
  OAI21X1  g04362(.A0(new_n6798_), .A1(new_n6793_), .B0(pi0074), .Y(new_n6799_));
  NAND3X1  g04363(.A(new_n6799_), .B(new_n6797_), .C(new_n3374_), .Y(new_n6800_));
  INVX1    g04364(.A(pi0178), .Y(new_n6801_));
  INVX1    g04365(.A(pi0183), .Y(new_n6802_));
  OR2X1    g04366(.A(pi0183), .B(pi0178), .Y(new_n6803_));
  AND2X1   g04367(.A(new_n6803_), .B(new_n5023_), .Y(new_n6804_));
  OAI21X1  g04368(.A0(new_n6802_), .A1(new_n6801_), .B0(new_n6804_), .Y(new_n6805_));
  AOI21X1  g04369(.A0(new_n6805_), .A1(new_n2933_), .B0(new_n5215_), .Y(new_n6806_));
  OAI21X1  g04370(.A0(new_n6792_), .A1(new_n2933_), .B0(new_n6806_), .Y(new_n6807_));
  OAI21X1  g04371(.A0(pi0100), .A1(pi0075), .B0(new_n6807_), .Y(new_n6808_));
  INVX1    g04372(.A(new_n6794_), .Y(new_n6809_));
  INVX1    g04373(.A(pi0191), .Y(new_n6810_));
  MX2X1    g04374(.A(new_n6810_), .B(new_n4162_), .S0(pi0299), .Y(new_n6811_));
  OR4X1    g04375(.A(new_n6811_), .B(new_n6809_), .C(new_n5048_), .D(new_n5215_), .Y(new_n6812_));
  AOI21X1  g04376(.A0(new_n6812_), .A1(new_n6808_), .B0(new_n4982_), .Y(new_n6813_));
  NOR2X1   g04377(.A(new_n6813_), .B(pi0055), .Y(new_n6814_));
  MX2X1    g04378(.A(pi0186), .B(pi0164), .S0(pi0299), .Y(new_n6815_));
  NAND4X1  g04379(.A(new_n6815_), .B(new_n6794_), .C(new_n5023_), .D(pi0232), .Y(new_n6816_));
  AOI21X1  g04380(.A0(new_n6816_), .A1(new_n6808_), .B0(new_n3091_), .Y(new_n6817_));
  INVX1    g04381(.A(pi0186), .Y(new_n6818_));
  AND2X1   g04382(.A(new_n5023_), .B(pi0232), .Y(new_n6819_));
  INVX1    g04383(.A(new_n6819_), .Y(new_n6820_));
  NOR3X1   g04384(.A(new_n6820_), .B(new_n4986_), .C(new_n2933_), .Y(new_n6821_));
  INVX1    g04385(.A(new_n6821_), .Y(new_n6822_));
  NOR2X1   g04386(.A(new_n6820_), .B(new_n5782_), .Y(new_n6823_));
  OAI21X1  g04387(.A0(new_n6823_), .A1(new_n6818_), .B0(pi0164), .Y(new_n6824_));
  AOI21X1  g04388(.A0(new_n6822_), .A1(new_n6818_), .B0(new_n6824_), .Y(new_n6825_));
  INVX1    g04389(.A(pi0164), .Y(new_n6826_));
  AND3X1   g04390(.A(new_n5023_), .B(new_n2933_), .C(pi0232), .Y(new_n6827_));
  INVX1    g04391(.A(new_n6827_), .Y(new_n6828_));
  AOI21X1  g04392(.A0(new_n2982_), .A1(new_n2939_), .B0(new_n6828_), .Y(new_n6829_));
  AND3X1   g04393(.A(new_n6829_), .B(pi0186), .C(new_n6826_), .Y(new_n6830_));
  OAI21X1  g04394(.A0(new_n6830_), .A1(new_n6825_), .B0(pi0038), .Y(new_n6831_));
  INVX1    g04395(.A(pi0176), .Y(new_n6832_));
  AND2X1   g04396(.A(pi0232), .B(new_n6832_), .Y(new_n6833_));
  NOR3X1   g04397(.A(pi0107), .B(pi0063), .C(pi0040), .Y(new_n6834_));
  INVX1    g04398(.A(new_n6834_), .Y(new_n6835_));
  OR3X1    g04399(.A(pi0102), .B(pi0081), .C(pi0064), .Y(new_n6836_));
  OR3X1    g04400(.A(new_n6836_), .B(new_n2459_), .C(new_n2457_), .Y(new_n6837_));
  OR2X1    g04401(.A(new_n6837_), .B(new_n2468_), .Y(new_n6838_));
  NAND2X1  g04402(.A(new_n2496_), .B(new_n2489_), .Y(new_n6839_));
  NOR4X1   g04403(.A(new_n6839_), .B(new_n6838_), .C(pi0060), .D(pi0053), .Y(new_n6840_));
  AND3X1   g04404(.A(new_n6840_), .B(new_n5897_), .C(new_n2494_), .Y(new_n6841_));
  INVX1    g04405(.A(new_n6841_), .Y(new_n6842_));
  NOR4X1   g04406(.A(new_n6842_), .B(new_n2526_), .C(pi0095), .D(pi0032), .Y(new_n6843_));
  NOR4X1   g04407(.A(new_n5239_), .B(new_n5231_), .C(new_n5030_), .D(new_n5024_), .Y(new_n6844_));
  OR2X1    g04408(.A(new_n6844_), .B(new_n5050_), .Y(new_n6845_));
  AND2X1   g04409(.A(new_n6845_), .B(new_n6843_), .Y(new_n6846_));
  AOI21X1  g04410(.A0(new_n6846_), .A1(new_n6255_), .B0(new_n6835_), .Y(new_n6847_));
  AND3X1   g04411(.A(pi0224), .B(new_n2940_), .C(pi0222), .Y(new_n6848_));
  NOR2X1   g04412(.A(new_n6848_), .B(new_n6835_), .Y(new_n6849_));
  NOR2X1   g04413(.A(new_n6849_), .B(new_n6847_), .Y(new_n6850_));
  INVX1    g04414(.A(pi0174), .Y(new_n6851_));
  AND3X1   g04415(.A(new_n6844_), .B(new_n6843_), .C(new_n5023_), .Y(new_n6852_));
  OAI21X1  g04416(.A0(new_n6852_), .A1(new_n6835_), .B0(new_n5042_), .Y(new_n6853_));
  NOR3X1   g04417(.A(new_n6853_), .B(new_n6849_), .C(new_n6851_), .Y(new_n6854_));
  OAI21X1  g04418(.A0(new_n6854_), .A1(new_n6850_), .B0(new_n2933_), .Y(new_n6855_));
  AND3X1   g04419(.A(pi0221), .B(pi0216), .C(new_n2934_), .Y(new_n6856_));
  OR2X1    g04420(.A(new_n6856_), .B(new_n6835_), .Y(new_n6857_));
  AND2X1   g04421(.A(new_n6857_), .B(pi0299), .Y(new_n6858_));
  AOI21X1  g04422(.A0(new_n6846_), .A1(new_n5023_), .B0(new_n6835_), .Y(new_n6859_));
  OAI21X1  g04423(.A0(new_n6859_), .A1(new_n5058_), .B0(new_n6847_), .Y(new_n6860_));
  AND3X1   g04424(.A(new_n6843_), .B(new_n5050_), .C(new_n5044_), .Y(new_n6861_));
  OR4X1    g04425(.A(new_n6861_), .B(new_n6835_), .C(new_n5048_), .D(pi0152), .Y(new_n6862_));
  AND3X1   g04426(.A(new_n6862_), .B(new_n6860_), .C(new_n3133_), .Y(new_n6863_));
  INVX1    g04427(.A(new_n6847_), .Y(new_n6864_));
  OR2X1    g04428(.A(new_n5058_), .B(new_n5048_), .Y(new_n6865_));
  AND2X1   g04429(.A(new_n6844_), .B(new_n6843_), .Y(new_n6866_));
  INVX1    g04430(.A(new_n6866_), .Y(new_n6867_));
  AOI21X1  g04431(.A0(new_n6867_), .A1(new_n6834_), .B0(new_n6865_), .Y(new_n6868_));
  AOI21X1  g04432(.A0(new_n6868_), .A1(pi0152), .B0(new_n6864_), .Y(new_n6869_));
  OAI21X1  g04433(.A0(new_n6869_), .A1(new_n3133_), .B0(new_n6856_), .Y(new_n6870_));
  OAI21X1  g04434(.A0(new_n6870_), .A1(new_n6863_), .B0(new_n6858_), .Y(new_n6871_));
  NAND2X1  g04435(.A(new_n6871_), .B(new_n6855_), .Y(new_n6872_));
  NAND4X1  g04436(.A(new_n6843_), .B(new_n5050_), .C(new_n5042_), .D(new_n5023_), .Y(new_n6873_));
  NAND3X1  g04437(.A(new_n6873_), .B(new_n6848_), .C(new_n6834_), .Y(new_n6874_));
  OAI21X1  g04438(.A0(new_n6848_), .A1(new_n6835_), .B0(new_n6874_), .Y(new_n6875_));
  NOR2X1   g04439(.A(new_n6875_), .B(pi0299), .Y(new_n6876_));
  OAI21X1  g04440(.A0(new_n6876_), .A1(new_n6872_), .B0(new_n6833_), .Y(new_n6877_));
  AND2X1   g04441(.A(pi0232), .B(pi0176), .Y(new_n6878_));
  OR2X1    g04442(.A(new_n6859_), .B(new_n5041_), .Y(new_n6879_));
  AOI21X1  g04443(.A0(new_n6879_), .A1(new_n6847_), .B0(new_n6849_), .Y(new_n6880_));
  AOI22X1  g04444(.A0(new_n6880_), .A1(new_n2933_), .B0(new_n6860_), .B1(new_n6858_), .Y(new_n6881_));
  OAI21X1  g04445(.A0(new_n6881_), .A1(pi0232), .B0(pi0039), .Y(new_n6882_));
  AOI21X1  g04446(.A0(new_n6878_), .A1(new_n6872_), .B0(new_n6882_), .Y(new_n6883_));
  AND2X1   g04447(.A(new_n6883_), .B(new_n6877_), .Y(new_n6884_));
  INVX1    g04448(.A(pi0193), .Y(new_n6885_));
  NOR2X1   g04449(.A(new_n6834_), .B(new_n2523_), .Y(new_n6886_));
  INVX1    g04450(.A(new_n6886_), .Y(new_n6887_));
  NOR2X1   g04451(.A(pi0479), .B(pi0040), .Y(new_n6888_));
  NOR3X1   g04452(.A(new_n6842_), .B(new_n2526_), .C(pi0032), .Y(new_n6889_));
  NOR2X1   g04453(.A(new_n6889_), .B(new_n2469_), .Y(new_n6890_));
  AOI22X1  g04454(.A0(new_n6890_), .A1(new_n6888_), .B0(new_n6887_), .B1(new_n3348_), .Y(new_n6891_));
  INVX1    g04455(.A(new_n6891_), .Y(new_n6892_));
  NOR2X1   g04456(.A(new_n6834_), .B(new_n2455_), .Y(new_n6893_));
  NOR2X1   g04457(.A(pi0096), .B(pi0072), .Y(new_n6894_));
  INVX1    g04458(.A(new_n2469_), .Y(new_n6895_));
  AOI21X1  g04459(.A0(new_n6842_), .A1(new_n6895_), .B0(new_n2535_), .Y(new_n6896_));
  INVX1    g04460(.A(new_n6896_), .Y(new_n6897_));
  INVX1    g04461(.A(new_n6840_), .Y(new_n6898_));
  AOI21X1  g04462(.A0(new_n6898_), .A1(new_n6895_), .B0(new_n2494_), .Y(new_n6899_));
  INVX1    g04463(.A(new_n6899_), .Y(new_n6900_));
  NOR3X1   g04464(.A(new_n6837_), .B(new_n2468_), .C(pi0060), .Y(new_n6901_));
  AOI21X1  g04465(.A0(new_n6735_), .A1(new_n2486_), .B0(new_n2729_), .Y(new_n6902_));
  INVX1    g04466(.A(new_n6902_), .Y(new_n6903_));
  OAI21X1  g04467(.A0(new_n6901_), .A1(new_n2485_), .B0(new_n6903_), .Y(new_n6904_));
  OR3X1    g04468(.A(pi0069), .B(pi0068), .C(pi0067), .Y(new_n6905_));
  OR4X1    g04469(.A(new_n6905_), .B(new_n2460_), .C(pi0111), .D(pi0036), .Y(new_n6906_));
  INVX1    g04470(.A(pi0066), .Y(new_n6907_));
  NAND4X1  g04471(.A(new_n2603_), .B(new_n2629_), .C(pi0073), .D(new_n6907_), .Y(new_n6908_));
  OR3X1    g04472(.A(new_n6908_), .B(new_n6906_), .C(new_n6837_), .Y(new_n6909_));
  NOR4X1   g04473(.A(new_n6909_), .B(new_n2464_), .C(pi0104), .D(pi0045), .Y(new_n6910_));
  AOI21X1  g04474(.A0(new_n6910_), .A1(new_n6733_), .B0(new_n2469_), .Y(new_n6911_));
  AOI21X1  g04475(.A0(new_n6911_), .A1(new_n6904_), .B0(new_n2490_), .Y(new_n6912_));
  OAI21X1  g04476(.A0(new_n2489_), .A1(new_n6895_), .B0(new_n2496_), .Y(new_n6913_));
  INVX1    g04477(.A(new_n2496_), .Y(new_n6914_));
  AOI21X1  g04478(.A0(new_n6914_), .A1(new_n6895_), .B0(pi0058), .Y(new_n6915_));
  OAI21X1  g04479(.A0(new_n6913_), .A1(new_n6912_), .B0(new_n6915_), .Y(new_n6916_));
  AOI21X1  g04480(.A0(new_n6916_), .A1(new_n6900_), .B0(pi0090), .Y(new_n6917_));
  AND3X1   g04481(.A(new_n6840_), .B(new_n2705_), .C(new_n2494_), .Y(new_n6918_));
  OAI21X1  g04482(.A0(new_n6918_), .A1(new_n2469_), .B0(pi0090), .Y(new_n6919_));
  NAND2X1  g04483(.A(new_n6919_), .B(new_n2524_), .Y(new_n6920_));
  AOI21X1  g04484(.A0(new_n2525_), .A1(new_n6895_), .B0(pi0070), .Y(new_n6921_));
  OAI21X1  g04485(.A0(new_n6920_), .A1(new_n6917_), .B0(new_n6921_), .Y(new_n6922_));
  AOI21X1  g04486(.A0(new_n6922_), .A1(new_n6897_), .B0(pi0051), .Y(new_n6923_));
  INVX1    g04487(.A(new_n6894_), .Y(new_n6924_));
  AOI21X1  g04488(.A0(new_n2469_), .A1(pi0051), .B0(new_n6924_), .Y(new_n6925_));
  INVX1    g04489(.A(new_n6925_), .Y(new_n6926_));
  OAI22X1  g04490(.A0(new_n6926_), .A1(new_n6923_), .B0(new_n6894_), .B1(new_n2469_), .Y(new_n6927_));
  AOI21X1  g04491(.A0(new_n6927_), .A1(new_n2529_), .B0(pi0032), .Y(new_n6928_));
  OAI21X1  g04492(.A0(new_n6928_), .A1(new_n6893_), .B0(new_n2523_), .Y(new_n6929_));
  AND2X1   g04493(.A(new_n6929_), .B(new_n6892_), .Y(new_n6930_));
  INVX1    g04494(.A(new_n6930_), .Y(new_n6931_));
  OR2X1    g04495(.A(pi0093), .B(pi0072), .Y(new_n6932_));
  NOR3X1   g04496(.A(new_n6932_), .B(new_n2478_), .C(pi0090), .Y(new_n6933_));
  NAND4X1  g04497(.A(new_n6933_), .B(new_n6840_), .C(new_n2705_), .D(new_n2494_), .Y(new_n6934_));
  AOI21X1  g04498(.A0(new_n6934_), .A1(new_n6834_), .B0(new_n2455_), .Y(new_n6935_));
  OAI21X1  g04499(.A0(new_n6935_), .A1(new_n6928_), .B0(new_n2523_), .Y(new_n6936_));
  NOR2X1   g04500(.A(new_n6936_), .B(pi0198), .Y(new_n6937_));
  NOR3X1   g04501(.A(new_n6937_), .B(new_n6931_), .C(new_n5023_), .Y(new_n6938_));
  AND2X1   g04502(.A(new_n6919_), .B(new_n2524_), .Y(new_n6939_));
  OAI21X1  g04503(.A0(new_n6904_), .A1(new_n6839_), .B0(new_n6895_), .Y(new_n6940_));
  AOI21X1  g04504(.A0(new_n6940_), .A1(new_n2494_), .B0(new_n6899_), .Y(new_n6941_));
  OAI21X1  g04505(.A0(new_n6941_), .A1(pi0090), .B0(new_n6939_), .Y(new_n6942_));
  AOI21X1  g04506(.A0(new_n6942_), .A1(new_n6921_), .B0(new_n6896_), .Y(new_n6943_));
  OAI21X1  g04507(.A0(new_n6943_), .A1(pi0051), .B0(new_n6925_), .Y(new_n6944_));
  OAI21X1  g04508(.A0(new_n6894_), .A1(new_n2469_), .B0(new_n6944_), .Y(new_n6945_));
  AOI21X1  g04509(.A0(new_n6945_), .A1(new_n2529_), .B0(pi0032), .Y(new_n6946_));
  OAI21X1  g04510(.A0(new_n6946_), .A1(new_n6935_), .B0(new_n2523_), .Y(new_n6947_));
  OR2X1    g04511(.A(new_n6947_), .B(pi0198), .Y(new_n6948_));
  OAI21X1  g04512(.A0(new_n6946_), .A1(new_n6893_), .B0(new_n2523_), .Y(new_n6949_));
  AND3X1   g04513(.A(new_n6949_), .B(new_n6887_), .C(new_n5023_), .Y(new_n6950_));
  AOI21X1  g04514(.A0(new_n6950_), .A1(new_n6948_), .B0(new_n6938_), .Y(new_n6951_));
  AOI21X1  g04515(.A0(new_n2469_), .A1(pi0032), .B0(pi0040), .Y(new_n6952_));
  INVX1    g04516(.A(new_n6952_), .Y(new_n6953_));
  INVX1    g04517(.A(new_n5010_), .Y(new_n6954_));
  AOI21X1  g04518(.A0(new_n6954_), .A1(new_n6895_), .B0(pi0032), .Y(new_n6955_));
  AOI21X1  g04519(.A0(new_n2469_), .A1(pi0093), .B0(new_n6954_), .Y(new_n6956_));
  OAI21X1  g04520(.A0(new_n6899_), .A1(new_n2469_), .B0(new_n2682_), .Y(new_n6957_));
  AND2X1   g04521(.A(new_n6957_), .B(new_n6919_), .Y(new_n6958_));
  OAI21X1  g04522(.A0(new_n6958_), .A1(pi0093), .B0(new_n6956_), .Y(new_n6959_));
  AOI21X1  g04523(.A0(new_n6959_), .A1(new_n6955_), .B0(new_n6953_), .Y(new_n6960_));
  NOR2X1   g04524(.A(new_n6960_), .B(pi0095), .Y(new_n6961_));
  NOR3X1   g04525(.A(new_n6961_), .B(new_n6886_), .C(new_n5048_), .Y(new_n6962_));
  NOR2X1   g04526(.A(new_n6962_), .B(new_n6938_), .Y(new_n6963_));
  MX2X1    g04527(.A(new_n6963_), .B(new_n6951_), .S0(new_n6802_), .Y(new_n6964_));
  OR2X1    g04528(.A(new_n6891_), .B(pi0174), .Y(new_n6965_));
  AOI21X1  g04529(.A0(new_n6964_), .A1(new_n2523_), .B0(new_n6965_), .Y(new_n6966_));
  NOR2X1   g04530(.A(new_n6937_), .B(new_n6931_), .Y(new_n6967_));
  AND2X1   g04531(.A(new_n5023_), .B(pi0183), .Y(new_n6968_));
  NOR2X1   g04532(.A(new_n6968_), .B(new_n6967_), .Y(new_n6969_));
  NAND3X1  g04533(.A(new_n6910_), .B(new_n6754_), .C(new_n2682_), .Y(new_n6970_));
  AND3X1   g04534(.A(new_n6970_), .B(new_n6957_), .C(new_n6919_), .Y(new_n6971_));
  OAI21X1  g04535(.A0(new_n6971_), .A1(pi0093), .B0(new_n6956_), .Y(new_n6972_));
  AOI21X1  g04536(.A0(new_n6972_), .A1(new_n6955_), .B0(new_n6953_), .Y(new_n6973_));
  NOR2X1   g04537(.A(new_n6973_), .B(pi0095), .Y(new_n6974_));
  OAI21X1  g04538(.A0(new_n6974_), .A1(new_n6891_), .B0(new_n5023_), .Y(new_n6975_));
  OAI21X1  g04539(.A0(new_n6975_), .A1(new_n6802_), .B0(pi0174), .Y(new_n6976_));
  OAI21X1  g04540(.A0(new_n6976_), .A1(new_n6969_), .B0(new_n5203_), .Y(new_n6977_));
  NOR2X1   g04541(.A(new_n6964_), .B(pi0174), .Y(new_n6978_));
  NOR3X1   g04542(.A(new_n6974_), .B(new_n6886_), .C(new_n5048_), .Y(new_n6979_));
  NOR2X1   g04543(.A(new_n6979_), .B(new_n6938_), .Y(new_n6980_));
  NOR3X1   g04544(.A(pi0468), .B(pi0332), .C(pi0040), .Y(new_n6981_));
  INVX1    g04545(.A(new_n6981_), .Y(new_n6982_));
  NAND2X1  g04546(.A(new_n6929_), .B(new_n6887_), .Y(new_n6983_));
  NOR3X1   g04547(.A(new_n6983_), .B(new_n6982_), .C(new_n6937_), .Y(new_n6984_));
  NOR2X1   g04548(.A(new_n6984_), .B(new_n6938_), .Y(new_n6985_));
  MX2X1    g04549(.A(new_n6985_), .B(new_n6980_), .S0(pi0183), .Y(new_n6986_));
  OAI21X1  g04550(.A0(new_n6986_), .A1(new_n6851_), .B0(pi0180), .Y(new_n6987_));
  OAI22X1  g04551(.A0(new_n6987_), .A1(new_n6978_), .B0(new_n6977_), .B1(new_n6966_), .Y(new_n6988_));
  INVX1    g04552(.A(new_n6938_), .Y(new_n6989_));
  AOI21X1  g04553(.A0(new_n2469_), .A1(new_n2529_), .B0(new_n2455_), .Y(new_n6990_));
  NOR4X1   g04554(.A(pi0093), .B(pi0090), .C(pi0058), .D(pi0035), .Y(new_n6991_));
  OAI22X1  g04555(.A0(new_n6991_), .A1(new_n6895_), .B0(new_n6916_), .B1(new_n5898_), .Y(new_n6992_));
  AOI21X1  g04556(.A0(new_n6992_), .A1(new_n2535_), .B0(new_n6896_), .Y(new_n6993_));
  OAI21X1  g04557(.A0(new_n6993_), .A1(pi0051), .B0(new_n6925_), .Y(new_n6994_));
  AOI21X1  g04558(.A0(new_n6924_), .A1(new_n6895_), .B0(pi0040), .Y(new_n6995_));
  AOI21X1  g04559(.A0(new_n6995_), .A1(new_n6994_), .B0(pi0032), .Y(new_n6996_));
  OAI22X1  g04560(.A0(new_n6996_), .A1(new_n6990_), .B0(new_n6834_), .B1(new_n2746_), .Y(new_n6997_));
  AOI21X1  g04561(.A0(new_n6997_), .A1(new_n2523_), .B0(new_n6891_), .Y(new_n6998_));
  NOR3X1   g04562(.A(new_n6834_), .B(pi0468), .C(pi0332), .Y(new_n6999_));
  MX2X1    g04563(.A(new_n6997_), .B(new_n6835_), .S0(pi0095), .Y(new_n7000_));
  AOI21X1  g04564(.A0(new_n2469_), .A1(new_n2529_), .B0(new_n2523_), .Y(new_n7001_));
  INVX1    g04565(.A(new_n7001_), .Y(new_n7002_));
  AND2X1   g04566(.A(new_n6934_), .B(new_n6834_), .Y(new_n7003_));
  OAI21X1  g04567(.A0(new_n7003_), .A1(pi0040), .B0(pi0032), .Y(new_n7004_));
  INVX1    g04568(.A(new_n7004_), .Y(new_n7005_));
  OAI21X1  g04569(.A0(new_n7005_), .A1(new_n6996_), .B0(new_n2523_), .Y(new_n7006_));
  AOI21X1  g04570(.A0(new_n7006_), .A1(new_n7002_), .B0(new_n7000_), .Y(new_n7007_));
  INVX1    g04571(.A(new_n7007_), .Y(new_n7008_));
  AOI21X1  g04572(.A0(new_n7008_), .A1(new_n2954_), .B0(new_n5048_), .Y(new_n7009_));
  OAI21X1  g04573(.A0(new_n7009_), .A1(new_n6999_), .B0(new_n6998_), .Y(new_n7010_));
  AOI21X1  g04574(.A0(new_n7010_), .A1(new_n6989_), .B0(pi0183), .Y(new_n7011_));
  NAND4X1  g04575(.A(new_n6754_), .B(new_n5010_), .C(new_n2483_), .D(new_n2455_), .Y(new_n7012_));
  NOR3X1   g04576(.A(new_n7012_), .B(new_n6909_), .C(new_n2624_), .Y(new_n7013_));
  OR2X1    g04577(.A(new_n7013_), .B(new_n6835_), .Y(new_n7014_));
  AND2X1   g04578(.A(new_n7014_), .B(new_n2523_), .Y(new_n7015_));
  NOR3X1   g04579(.A(new_n7015_), .B(new_n6891_), .C(new_n5048_), .Y(new_n7016_));
  OAI21X1  g04580(.A0(new_n7016_), .A1(new_n6938_), .B0(pi0183), .Y(new_n7017_));
  NAND2X1  g04581(.A(new_n7017_), .B(pi0174), .Y(new_n7018_));
  OAI21X1  g04582(.A0(new_n6937_), .A1(new_n6931_), .B0(new_n5048_), .Y(new_n7019_));
  AOI21X1  g04583(.A0(new_n2587_), .A1(new_n2656_), .B0(new_n6991_), .Y(new_n7020_));
  AND3X1   g04584(.A(new_n6940_), .B(new_n5897_), .C(new_n2494_), .Y(new_n7021_));
  OAI21X1  g04585(.A0(new_n7021_), .A1(new_n7020_), .B0(new_n2535_), .Y(new_n7022_));
  AOI21X1  g04586(.A0(new_n7022_), .A1(new_n6897_), .B0(pi0051), .Y(new_n7023_));
  OAI22X1  g04587(.A0(new_n7023_), .A1(new_n6926_), .B0(new_n6894_), .B1(new_n2469_), .Y(new_n7024_));
  AOI21X1  g04588(.A0(new_n7024_), .A1(new_n2529_), .B0(pi0032), .Y(new_n7025_));
  OR2X1    g04589(.A(new_n7025_), .B(new_n6893_), .Y(new_n7026_));
  AOI21X1  g04590(.A0(new_n7026_), .A1(new_n2523_), .B0(new_n6891_), .Y(new_n7027_));
  OAI21X1  g04591(.A0(new_n7025_), .A1(new_n6935_), .B0(new_n2523_), .Y(new_n7028_));
  OR2X1    g04592(.A(new_n7028_), .B(pi0198), .Y(new_n7029_));
  AND2X1   g04593(.A(new_n7029_), .B(new_n7027_), .Y(new_n7030_));
  OAI21X1  g04594(.A0(new_n7030_), .A1(new_n5048_), .B0(new_n7019_), .Y(new_n7031_));
  OR2X1    g04595(.A(new_n7031_), .B(pi0183), .Y(new_n7032_));
  AOI21X1  g04596(.A0(new_n6835_), .A1(new_n2523_), .B0(new_n6891_), .Y(new_n7033_));
  MX2X1    g04597(.A(new_n7033_), .B(new_n6967_), .S0(new_n5048_), .Y(new_n7034_));
  AOI21X1  g04598(.A0(new_n7034_), .A1(pi0183), .B0(pi0174), .Y(new_n7035_));
  AOI21X1  g04599(.A0(new_n7035_), .A1(new_n7032_), .B0(pi0180), .Y(new_n7036_));
  OAI21X1  g04600(.A0(new_n7018_), .A1(new_n7011_), .B0(new_n7036_), .Y(new_n7037_));
  INVX1    g04601(.A(new_n7009_), .Y(new_n7038_));
  OAI21X1  g04602(.A0(new_n7038_), .A1(new_n7000_), .B0(new_n6989_), .Y(new_n7039_));
  AND2X1   g04603(.A(new_n7039_), .B(new_n6802_), .Y(new_n7040_));
  OR3X1    g04604(.A(new_n7015_), .B(new_n6886_), .C(new_n5048_), .Y(new_n7041_));
  AOI21X1  g04605(.A0(new_n7041_), .A1(new_n6989_), .B0(new_n6802_), .Y(new_n7042_));
  OR3X1    g04606(.A(new_n7042_), .B(new_n7040_), .C(new_n6851_), .Y(new_n7043_));
  INVX1    g04607(.A(new_n6999_), .Y(new_n7044_));
  NAND3X1  g04608(.A(new_n7019_), .B(new_n7044_), .C(pi0183), .Y(new_n7045_));
  AND2X1   g04609(.A(new_n2469_), .B(new_n2529_), .Y(new_n7046_));
  INVX1    g04610(.A(new_n6990_), .Y(new_n7047_));
  OAI21X1  g04611(.A0(new_n7024_), .A1(pi0040), .B0(new_n2455_), .Y(new_n7048_));
  AND2X1   g04612(.A(new_n7048_), .B(new_n7047_), .Y(new_n7049_));
  MX2X1    g04613(.A(new_n7049_), .B(new_n7046_), .S0(pi0095), .Y(new_n7050_));
  AOI21X1  g04614(.A0(new_n7048_), .A1(new_n7004_), .B0(pi0095), .Y(new_n7051_));
  NOR2X1   g04615(.A(new_n7051_), .B(new_n7001_), .Y(new_n7052_));
  MX2X1    g04616(.A(new_n7052_), .B(new_n7050_), .S0(pi0198), .Y(new_n7053_));
  OAI21X1  g04617(.A0(new_n7053_), .A1(new_n6982_), .B0(new_n6989_), .Y(new_n7054_));
  AOI21X1  g04618(.A0(new_n7054_), .A1(new_n6802_), .B0(pi0174), .Y(new_n7055_));
  AOI21X1  g04619(.A0(new_n7055_), .A1(new_n7045_), .B0(new_n5203_), .Y(new_n7056_));
  AOI21X1  g04620(.A0(new_n7056_), .A1(new_n7043_), .B0(new_n6885_), .Y(new_n7057_));
  AOI22X1  g04621(.A0(new_n7057_), .A1(new_n7037_), .B0(new_n6988_), .B1(new_n6885_), .Y(new_n7058_));
  AND2X1   g04622(.A(pi0299), .B(pi0158), .Y(new_n7059_));
  INVX1    g04623(.A(new_n7059_), .Y(new_n7060_));
  NOR2X1   g04624(.A(new_n6936_), .B(pi0210), .Y(new_n7061_));
  NOR3X1   g04625(.A(new_n7061_), .B(new_n6931_), .C(new_n5023_), .Y(new_n7062_));
  OR2X1    g04626(.A(new_n6947_), .B(pi0210), .Y(new_n7063_));
  AOI21X1  g04627(.A0(new_n7063_), .A1(new_n6950_), .B0(new_n7062_), .Y(new_n7064_));
  OR2X1    g04628(.A(new_n7064_), .B(pi0152), .Y(new_n7065_));
  NOR2X1   g04629(.A(new_n7061_), .B(new_n6931_), .Y(new_n7066_));
  NOR2X1   g04630(.A(new_n7061_), .B(new_n6983_), .Y(new_n7067_));
  MX2X1    g04631(.A(new_n7067_), .B(new_n7066_), .S0(new_n5048_), .Y(new_n7068_));
  AOI21X1  g04632(.A0(new_n7068_), .A1(pi0152), .B0(pi0172), .Y(new_n7069_));
  INVX1    g04633(.A(new_n7062_), .Y(new_n7070_));
  AOI21X1  g04634(.A0(new_n7008_), .A1(new_n2777_), .B0(new_n5048_), .Y(new_n7071_));
  INVX1    g04635(.A(new_n7071_), .Y(new_n7072_));
  OAI21X1  g04636(.A0(new_n7072_), .A1(new_n7000_), .B0(new_n7070_), .Y(new_n7073_));
  NAND2X1  g04637(.A(new_n7073_), .B(pi0152), .Y(new_n7074_));
  AOI21X1  g04638(.A0(new_n7028_), .A1(new_n6887_), .B0(pi0210), .Y(new_n7075_));
  MX2X1    g04639(.A(new_n7026_), .B(new_n6835_), .S0(pi0095), .Y(new_n7076_));
  NOR3X1   g04640(.A(new_n7076_), .B(new_n7075_), .C(new_n5048_), .Y(new_n7077_));
  OAI21X1  g04641(.A0(new_n7077_), .A1(new_n7062_), .B0(new_n3193_), .Y(new_n7078_));
  AND2X1   g04642(.A(new_n7078_), .B(pi0172), .Y(new_n7079_));
  AOI22X1  g04643(.A0(new_n7079_), .A1(new_n7074_), .B0(new_n7069_), .B1(new_n7065_), .Y(new_n7080_));
  OR2X1    g04644(.A(new_n7080_), .B(new_n7060_), .Y(new_n7081_));
  OAI21X1  g04645(.A0(new_n7071_), .A1(new_n6999_), .B0(new_n6998_), .Y(new_n7082_));
  INVX1    g04646(.A(new_n7082_), .Y(new_n7083_));
  INVX1    g04647(.A(pi0172), .Y(new_n7084_));
  OAI21X1  g04648(.A0(new_n7075_), .A1(new_n5048_), .B0(new_n7044_), .Y(new_n7085_));
  NAND2X1  g04649(.A(new_n7085_), .B(new_n7027_), .Y(new_n7086_));
  AOI21X1  g04650(.A0(new_n7086_), .A1(new_n3193_), .B0(new_n7084_), .Y(new_n7087_));
  OAI21X1  g04651(.A0(new_n7083_), .A1(new_n3193_), .B0(new_n7087_), .Y(new_n7088_));
  AND2X1   g04652(.A(new_n6949_), .B(new_n6892_), .Y(new_n7089_));
  AND3X1   g04653(.A(new_n7089_), .B(new_n7063_), .C(new_n5023_), .Y(new_n7090_));
  OR2X1    g04654(.A(new_n7090_), .B(pi0152), .Y(new_n7091_));
  INVX1    g04655(.A(new_n7066_), .Y(new_n7092_));
  AOI21X1  g04656(.A0(new_n7092_), .A1(pi0152), .B0(pi0172), .Y(new_n7093_));
  INVX1    g04657(.A(pi0158), .Y(new_n7094_));
  AND2X1   g04658(.A(pi0299), .B(new_n7094_), .Y(new_n7095_));
  INVX1    g04659(.A(new_n7095_), .Y(new_n7096_));
  OR2X1    g04660(.A(new_n7096_), .B(new_n7062_), .Y(new_n7097_));
  AOI21X1  g04661(.A0(new_n7093_), .A1(new_n7091_), .B0(new_n7097_), .Y(new_n7098_));
  AOI21X1  g04662(.A0(new_n7098_), .A1(new_n7088_), .B0(pi0149), .Y(new_n7099_));
  AND2X1   g04663(.A(new_n7099_), .B(new_n7081_), .Y(new_n7100_));
  INVX1    g04664(.A(pi0149), .Y(new_n7101_));
  OAI21X1  g04665(.A0(new_n7062_), .A1(new_n6979_), .B0(pi0152), .Y(new_n7102_));
  OAI21X1  g04666(.A0(new_n7062_), .A1(new_n6962_), .B0(new_n3193_), .Y(new_n7103_));
  NAND3X1  g04667(.A(new_n7103_), .B(new_n7102_), .C(new_n7084_), .Y(new_n7104_));
  AOI21X1  g04668(.A0(new_n7070_), .A1(new_n7041_), .B0(new_n3193_), .Y(new_n7105_));
  NOR2X1   g04669(.A(new_n7066_), .B(new_n5023_), .Y(new_n7106_));
  NOR3X1   g04670(.A(new_n7106_), .B(new_n6999_), .C(pi0152), .Y(new_n7107_));
  OR3X1    g04671(.A(new_n7107_), .B(new_n7105_), .C(new_n7084_), .Y(new_n7108_));
  AOI21X1  g04672(.A0(new_n7108_), .A1(new_n7104_), .B0(new_n7060_), .Y(new_n7109_));
  OAI21X1  g04673(.A0(new_n7062_), .A1(new_n7016_), .B0(pi0152), .Y(new_n7110_));
  AOI21X1  g04674(.A0(new_n7033_), .A1(new_n5023_), .B0(new_n7062_), .Y(new_n7111_));
  OR2X1    g04675(.A(new_n7111_), .B(pi0152), .Y(new_n7112_));
  NAND3X1  g04676(.A(new_n7112_), .B(new_n7110_), .C(pi0172), .Y(new_n7113_));
  OAI21X1  g04677(.A0(new_n6960_), .A1(pi0095), .B0(new_n6892_), .Y(new_n7114_));
  AND2X1   g04678(.A(new_n7114_), .B(new_n5023_), .Y(new_n7115_));
  OR3X1    g04679(.A(new_n7115_), .B(new_n7106_), .C(pi0152), .Y(new_n7116_));
  INVX1    g04680(.A(new_n7106_), .Y(new_n7117_));
  NAND3X1  g04681(.A(new_n7117_), .B(new_n6975_), .C(pi0152), .Y(new_n7118_));
  NAND3X1  g04682(.A(new_n7118_), .B(new_n7116_), .C(new_n7084_), .Y(new_n7119_));
  AOI21X1  g04683(.A0(new_n7119_), .A1(new_n7113_), .B0(new_n7096_), .Y(new_n7120_));
  NOR3X1   g04684(.A(new_n7120_), .B(new_n7109_), .C(new_n7101_), .Y(new_n7121_));
  OAI22X1  g04685(.A0(new_n7121_), .A1(new_n7100_), .B0(new_n7058_), .B1(pi0299), .Y(new_n7122_));
  OAI21X1  g04686(.A0(new_n6936_), .A1(new_n5009_), .B0(new_n6930_), .Y(new_n7123_));
  NAND2X1  g04687(.A(new_n7123_), .B(new_n5215_), .Y(new_n7124_));
  NAND2X1  g04688(.A(new_n7124_), .B(new_n2939_), .Y(new_n7125_));
  AOI21X1  g04689(.A0(new_n7122_), .A1(pi0232), .B0(new_n7125_), .Y(new_n7126_));
  OAI21X1  g04690(.A0(new_n7126_), .A1(new_n6884_), .B0(new_n2979_), .Y(new_n7127_));
  AOI21X1  g04691(.A0(new_n7127_), .A1(new_n6831_), .B0(pi0100), .Y(new_n7128_));
  AND2X1   g04692(.A(new_n6807_), .B(pi0100), .Y(new_n7129_));
  OR2X1    g04693(.A(new_n7129_), .B(pi0087), .Y(new_n7130_));
  NAND3X1  g04694(.A(new_n6815_), .B(new_n5023_), .C(pi0232), .Y(new_n7131_));
  NOR2X1   g04695(.A(new_n7131_), .B(new_n2979_), .Y(new_n7132_));
  AOI21X1  g04696(.A0(new_n7132_), .A1(new_n3007_), .B0(new_n7129_), .Y(new_n7133_));
  AOI21X1  g04697(.A0(new_n6834_), .A1(new_n3251_), .B0(new_n3131_), .Y(new_n7134_));
  AOI21X1  g04698(.A0(new_n7134_), .A1(new_n7133_), .B0(new_n5295_), .Y(new_n7135_));
  OAI21X1  g04699(.A0(new_n7130_), .A1(new_n7128_), .B0(new_n7135_), .Y(new_n7136_));
  AND2X1   g04700(.A(new_n6807_), .B(pi0075), .Y(new_n7137_));
  AND2X1   g04701(.A(pi0092), .B(new_n3073_), .Y(new_n7138_));
  AND2X1   g04702(.A(new_n6834_), .B(new_n3251_), .Y(new_n7139_));
  INVX1    g04703(.A(new_n7139_), .Y(new_n7140_));
  OR2X1    g04704(.A(pi0087), .B(pi0039), .Y(new_n7141_));
  INVX1    g04705(.A(new_n6843_), .Y(new_n7142_));
  AOI21X1  g04706(.A0(pi0299), .A1(new_n3133_), .B0(new_n5215_), .Y(new_n7143_));
  OR2X1    g04707(.A(pi0299), .B(pi0176), .Y(new_n7144_));
  AND3X1   g04708(.A(new_n7144_), .B(new_n7143_), .C(new_n5023_), .Y(new_n7145_));
  NOR3X1   g04709(.A(new_n7145_), .B(new_n7142_), .C(new_n7141_), .Y(new_n7146_));
  OAI21X1  g04710(.A0(new_n7146_), .A1(new_n7140_), .B0(new_n7133_), .Y(new_n7147_));
  AOI21X1  g04711(.A0(new_n7147_), .A1(new_n7138_), .B0(new_n7137_), .Y(new_n7148_));
  AOI21X1  g04712(.A0(new_n7148_), .A1(new_n7136_), .B0(pi0054), .Y(new_n7149_));
  OAI21X1  g04713(.A0(new_n7149_), .A1(new_n6817_), .B0(new_n4982_), .Y(new_n7150_));
  NAND2X1  g04714(.A(new_n6799_), .B(pi0055), .Y(new_n7151_));
  NOR2X1   g04715(.A(new_n6796_), .B(new_n3091_), .Y(new_n7152_));
  INVX1    g04716(.A(new_n7152_), .Y(new_n7153_));
  AOI21X1  g04717(.A0(new_n6792_), .A1(pi0232), .B0(new_n3073_), .Y(new_n7154_));
  OR2X1    g04718(.A(new_n7154_), .B(pi0092), .Y(new_n7155_));
  INVX1    g04719(.A(new_n3101_), .Y(new_n7156_));
  AOI21X1  g04720(.A0(new_n6819_), .A1(pi0164), .B0(new_n2979_), .Y(new_n7157_));
  NOR2X1   g04721(.A(new_n7157_), .B(new_n7156_), .Y(new_n7158_));
  AOI21X1  g04722(.A0(new_n6819_), .A1(pi0149), .B0(pi0039), .Y(new_n7159_));
  AOI21X1  g04723(.A0(new_n7159_), .A1(new_n6843_), .B0(new_n6835_), .Y(new_n7160_));
  OAI21X1  g04724(.A0(new_n7160_), .A1(pi0038), .B0(new_n7158_), .Y(new_n7161_));
  AOI21X1  g04725(.A0(new_n6792_), .A1(pi0232), .B0(new_n3007_), .Y(new_n7162_));
  NOR2X1   g04726(.A(new_n6834_), .B(pi0038), .Y(new_n7163_));
  NOR4X1   g04727(.A(new_n7163_), .B(new_n7157_), .C(pi0100), .D(new_n3131_), .Y(new_n7164_));
  NOR2X1   g04728(.A(new_n7164_), .B(new_n7162_), .Y(new_n7165_));
  AOI21X1  g04729(.A0(new_n7165_), .A1(new_n7161_), .B0(pi0075), .Y(new_n7166_));
  OR4X1    g04730(.A(new_n7163_), .B(new_n7157_), .C(pi0100), .D(pi0075), .Y(new_n7167_));
  NOR2X1   g04731(.A(new_n6793_), .B(new_n3079_), .Y(new_n7168_));
  AOI21X1  g04732(.A0(new_n7168_), .A1(new_n7167_), .B0(pi0054), .Y(new_n7169_));
  OAI21X1  g04733(.A0(new_n7166_), .A1(new_n7155_), .B0(new_n7169_), .Y(new_n7170_));
  AOI21X1  g04734(.A0(new_n7170_), .A1(new_n7153_), .B0(pi0074), .Y(new_n7171_));
  OAI21X1  g04735(.A0(new_n7171_), .A1(new_n7151_), .B0(new_n3123_), .Y(new_n7172_));
  AOI21X1  g04736(.A0(new_n7150_), .A1(new_n6814_), .B0(new_n7172_), .Y(new_n7173_));
  AND3X1   g04737(.A(new_n6819_), .B(pi0164), .C(pi0038), .Y(new_n7174_));
  AOI21X1  g04738(.A0(new_n7174_), .A1(new_n6794_), .B0(new_n6793_), .Y(new_n7175_));
  OAI21X1  g04739(.A0(new_n6796_), .A1(new_n3091_), .B0(new_n7175_), .Y(new_n7176_));
  NAND2X1  g04740(.A(new_n7176_), .B(new_n4982_), .Y(new_n7177_));
  AOI21X1  g04741(.A0(new_n7177_), .A1(new_n6799_), .B0(new_n3123_), .Y(new_n7178_));
  NOR4X1   g04742(.A(pi0107), .B(pi0063), .C(pi0040), .D(pi0038), .Y(new_n7179_));
  AND3X1   g04743(.A(new_n7179_), .B(new_n6794_), .C(new_n3102_), .Y(new_n7180_));
  AND2X1   g04744(.A(new_n7180_), .B(new_n4975_), .Y(new_n7181_));
  OR3X1    g04745(.A(new_n7181_), .B(new_n7178_), .C(new_n3374_), .Y(new_n7182_));
  OAI21X1  g04746(.A0(new_n7182_), .A1(new_n7173_), .B0(new_n6800_), .Y(new_n7183_));
  OAI21X1  g04747(.A0(new_n6788_), .A1(pi0033), .B0(new_n7183_), .Y(new_n7184_));
  AOI21X1  g04748(.A0(new_n6787_), .A1(new_n6783_), .B0(pi0033), .Y(new_n7185_));
  OR2X1    g04749(.A(new_n7178_), .B(new_n3374_), .Y(new_n7186_));
  INVX1    g04750(.A(new_n6856_), .Y(new_n7187_));
  OAI21X1  g04751(.A0(new_n5236_), .A1(new_n6865_), .B0(pi0154), .Y(new_n7188_));
  NOR4X1   g04752(.A(new_n5239_), .B(new_n5228_), .C(new_n5224_), .D(new_n6865_), .Y(new_n7189_));
  OR2X1    g04753(.A(new_n7189_), .B(pi0154), .Y(new_n7190_));
  AND2X1   g04754(.A(new_n7190_), .B(new_n3193_), .Y(new_n7191_));
  AND2X1   g04755(.A(new_n5947_), .B(pi1091), .Y(new_n7192_));
  AND3X1   g04756(.A(new_n7192_), .B(new_n5059_), .C(new_n5023_), .Y(new_n7193_));
  AND2X1   g04757(.A(pi0154), .B(pi0152), .Y(new_n7194_));
  AOI22X1  g04758(.A0(new_n7194_), .A1(new_n7193_), .B0(new_n7191_), .B1(new_n7188_), .Y(new_n7195_));
  OAI21X1  g04759(.A0(new_n7195_), .A1(new_n7187_), .B0(pi0299), .Y(new_n7196_));
  INVX1    g04760(.A(new_n6833_), .Y(new_n7197_));
  INVX1    g04761(.A(new_n6878_), .Y(new_n7198_));
  OR2X1    g04762(.A(new_n5041_), .B(new_n5048_), .Y(new_n7199_));
  NOR4X1   g04763(.A(new_n5239_), .B(new_n5228_), .C(new_n5224_), .D(new_n7199_), .Y(new_n7200_));
  NAND3X1  g04764(.A(new_n7200_), .B(new_n6848_), .C(new_n6851_), .Y(new_n7201_));
  AND2X1   g04765(.A(new_n7201_), .B(new_n2933_), .Y(new_n7202_));
  INVX1    g04766(.A(new_n6848_), .Y(new_n7203_));
  NOR3X1   g04767(.A(new_n7203_), .B(new_n5236_), .C(new_n7199_), .Y(new_n7204_));
  NAND4X1  g04768(.A(new_n6848_), .B(new_n7192_), .C(new_n5042_), .D(new_n5023_), .Y(new_n7205_));
  OAI21X1  g04769(.A0(new_n7205_), .A1(new_n6851_), .B0(new_n2933_), .Y(new_n7206_));
  AOI21X1  g04770(.A0(new_n7204_), .A1(new_n6851_), .B0(new_n7206_), .Y(new_n7207_));
  OAI22X1  g04771(.A0(new_n7207_), .A1(new_n7198_), .B0(new_n7202_), .B1(new_n7197_), .Y(new_n7208_));
  AND3X1   g04772(.A(new_n7208_), .B(new_n7196_), .C(pi0039), .Y(new_n7209_));
  AOI21X1  g04773(.A0(new_n2477_), .A1(new_n2705_), .B0(new_n2682_), .Y(new_n7210_));
  NOR3X1   g04774(.A(new_n7210_), .B(new_n4992_), .C(new_n2525_), .Y(new_n7211_));
  INVX1    g04775(.A(new_n7211_), .Y(new_n7212_));
  NOR4X1   g04776(.A(new_n2525_), .B(new_n2498_), .C(new_n2493_), .D(pi0090), .Y(new_n7213_));
  AND2X1   g04777(.A(new_n7213_), .B(new_n6895_), .Y(new_n7214_));
  AOI21X1  g04778(.A0(new_n7214_), .A1(new_n6912_), .B0(pi0070), .Y(new_n7215_));
  NOR4X1   g04779(.A(new_n5881_), .B(new_n2848_), .C(pi0096), .D(pi0051), .Y(new_n7216_));
  INVX1    g04780(.A(new_n7216_), .Y(new_n7217_));
  AOI21X1  g04781(.A0(new_n7215_), .A1(new_n7212_), .B0(new_n7217_), .Y(new_n7218_));
  INVX1    g04782(.A(new_n7218_), .Y(new_n7219_));
  NOR2X1   g04783(.A(new_n5174_), .B(pi0095), .Y(new_n7220_));
  NOR2X1   g04784(.A(new_n7217_), .B(new_n7215_), .Y(new_n7221_));
  NOR2X1   g04785(.A(new_n7221_), .B(new_n7220_), .Y(new_n7222_));
  OAI21X1  g04786(.A0(new_n7222_), .A1(pi0198), .B0(new_n7219_), .Y(new_n7223_));
  AND3X1   g04787(.A(new_n6910_), .B(new_n6754_), .C(new_n6895_), .Y(new_n7224_));
  INVX1    g04788(.A(new_n7224_), .Y(new_n7225_));
  AND3X1   g04789(.A(new_n7225_), .B(new_n4991_), .C(new_n2682_), .Y(new_n7226_));
  NOR4X1   g04790(.A(new_n7226_), .B(new_n7210_), .C(new_n6932_), .D(new_n2478_), .Y(new_n7227_));
  NOR2X1   g04791(.A(pi0095), .B(pi0032), .Y(new_n7228_));
  AND3X1   g04792(.A(new_n5023_), .B(new_n7228_), .C(new_n2529_), .Y(new_n7229_));
  AND2X1   g04793(.A(new_n7229_), .B(new_n7227_), .Y(new_n7230_));
  INVX1    g04794(.A(new_n7230_), .Y(new_n7231_));
  OAI21X1  g04795(.A0(new_n7231_), .A1(pi0183), .B0(new_n6851_), .Y(new_n7232_));
  AOI21X1  g04796(.A0(new_n7223_), .A1(new_n6968_), .B0(new_n7232_), .Y(new_n7233_));
  AOI21X1  g04797(.A0(new_n7213_), .A1(new_n6903_), .B0(pi0070), .Y(new_n7234_));
  AOI21X1  g04798(.A0(new_n7234_), .A1(new_n7212_), .B0(new_n7217_), .Y(new_n7235_));
  OR2X1    g04799(.A(new_n7235_), .B(new_n5198_), .Y(new_n7236_));
  AND2X1   g04800(.A(new_n7236_), .B(new_n5023_), .Y(new_n7237_));
  NOR4X1   g04801(.A(new_n7210_), .B(new_n6932_), .C(new_n4992_), .D(new_n2478_), .Y(new_n7238_));
  AND2X1   g04802(.A(new_n7238_), .B(new_n7229_), .Y(new_n7239_));
  INVX1    g04803(.A(new_n7239_), .Y(new_n7240_));
  OAI21X1  g04804(.A0(new_n7240_), .A1(pi0183), .B0(pi0174), .Y(new_n7241_));
  AOI21X1  g04805(.A0(new_n7237_), .A1(pi0183), .B0(new_n7241_), .Y(new_n7242_));
  OAI21X1  g04806(.A0(new_n7242_), .A1(new_n7233_), .B0(pi0193), .Y(new_n7243_));
  NOR2X1   g04807(.A(new_n7221_), .B(new_n5198_), .Y(new_n7244_));
  INVX1    g04808(.A(new_n7234_), .Y(new_n7245_));
  AOI21X1  g04809(.A0(new_n7245_), .A1(new_n7216_), .B0(new_n5198_), .Y(new_n7246_));
  NAND2X1  g04810(.A(new_n7246_), .B(pi0174), .Y(new_n7247_));
  NAND2X1  g04811(.A(new_n7247_), .B(new_n6968_), .Y(new_n7248_));
  AOI21X1  g04812(.A0(new_n7244_), .A1(new_n6851_), .B0(new_n7248_), .Y(new_n7249_));
  INVX1    g04813(.A(new_n7228_), .Y(new_n7250_));
  NAND4X1  g04814(.A(new_n6933_), .B(new_n6910_), .C(new_n6754_), .D(new_n6895_), .Y(new_n7251_));
  NOR3X1   g04815(.A(new_n7251_), .B(new_n6982_), .C(new_n7250_), .Y(new_n7252_));
  AND3X1   g04816(.A(new_n7252_), .B(new_n6802_), .C(new_n6851_), .Y(new_n7253_));
  OR3X1    g04817(.A(new_n7253_), .B(new_n7249_), .C(pi0193), .Y(new_n7254_));
  AND2X1   g04818(.A(new_n5023_), .B(new_n2880_), .Y(new_n7255_));
  INVX1    g04819(.A(new_n7255_), .Y(new_n7256_));
  OAI21X1  g04820(.A0(new_n7256_), .A1(new_n5203_), .B0(new_n2933_), .Y(new_n7257_));
  AOI21X1  g04821(.A0(new_n7254_), .A1(new_n7243_), .B0(new_n7257_), .Y(new_n7258_));
  AND2X1   g04822(.A(pi0232), .B(new_n2939_), .Y(new_n7259_));
  INVX1    g04823(.A(new_n7259_), .Y(new_n7260_));
  NOR3X1   g04824(.A(new_n7221_), .B(new_n5175_), .C(pi0152), .Y(new_n7261_));
  OAI21X1  g04825(.A0(new_n7219_), .A1(new_n7084_), .B0(new_n7261_), .Y(new_n7262_));
  AOI21X1  g04826(.A0(new_n7245_), .A1(new_n7216_), .B0(new_n5175_), .Y(new_n7263_));
  AOI21X1  g04827(.A0(new_n7235_), .A1(pi0172), .B0(new_n3193_), .Y(new_n7264_));
  NAND2X1  g04828(.A(new_n5023_), .B(pi0149), .Y(new_n7265_));
  AOI21X1  g04829(.A0(new_n7264_), .A1(new_n7263_), .B0(new_n7265_), .Y(new_n7266_));
  OAI21X1  g04830(.A0(new_n7231_), .A1(pi0152), .B0(new_n7240_), .Y(new_n7267_));
  AND3X1   g04831(.A(new_n7252_), .B(new_n7084_), .C(new_n3193_), .Y(new_n7268_));
  AOI21X1  g04832(.A0(new_n7267_), .A1(pi0172), .B0(new_n7268_), .Y(new_n7269_));
  AOI21X1  g04833(.A0(new_n7255_), .A1(pi0158), .B0(new_n2933_), .Y(new_n7270_));
  OAI21X1  g04834(.A0(new_n7269_), .A1(pi0149), .B0(new_n7270_), .Y(new_n7271_));
  AOI21X1  g04835(.A0(new_n7266_), .A1(new_n7262_), .B0(new_n7271_), .Y(new_n7272_));
  NOR3X1   g04836(.A(new_n7272_), .B(new_n7260_), .C(new_n7258_), .Y(new_n7273_));
  OAI21X1  g04837(.A0(new_n7273_), .A1(new_n7209_), .B0(new_n2979_), .Y(new_n7274_));
  AND2X1   g04838(.A(new_n6831_), .B(new_n3131_), .Y(new_n7275_));
  OAI21X1  g04839(.A0(new_n7132_), .A1(new_n3131_), .B0(new_n3007_), .Y(new_n7276_));
  AOI21X1  g04840(.A0(new_n7275_), .A1(new_n7274_), .B0(new_n7276_), .Y(new_n7277_));
  OAI21X1  g04841(.A0(new_n7277_), .A1(new_n7129_), .B0(new_n3084_), .Y(new_n7278_));
  INVX1    g04842(.A(new_n7138_), .Y(new_n7279_));
  NOR2X1   g04843(.A(pi0087), .B(pi0038), .Y(new_n7280_));
  NAND4X1  g04844(.A(new_n7280_), .B(new_n7145_), .C(new_n4986_), .D(new_n3007_), .Y(new_n7281_));
  AOI21X1  g04845(.A0(new_n7281_), .A1(new_n7133_), .B0(new_n7279_), .Y(new_n7282_));
  NOR2X1   g04846(.A(new_n7282_), .B(new_n7137_), .Y(new_n7283_));
  AOI21X1  g04847(.A0(new_n7283_), .A1(new_n7278_), .B0(pi0054), .Y(new_n7284_));
  OAI21X1  g04848(.A0(new_n7284_), .A1(new_n6817_), .B0(new_n4982_), .Y(new_n7285_));
  AND3X1   g04849(.A(new_n6819_), .B(new_n4986_), .C(pi0149), .Y(new_n7286_));
  OAI21X1  g04850(.A0(new_n7286_), .A1(pi0038), .B0(new_n7158_), .Y(new_n7287_));
  AND2X1   g04851(.A(new_n3007_), .B(pi0087), .Y(new_n7288_));
  AOI21X1  g04852(.A0(new_n7174_), .A1(new_n7288_), .B0(new_n7162_), .Y(new_n7289_));
  AOI21X1  g04853(.A0(new_n7289_), .A1(new_n7287_), .B0(pi0075), .Y(new_n7290_));
  AOI21X1  g04854(.A0(new_n7175_), .A1(pi0092), .B0(pi0054), .Y(new_n7291_));
  OAI21X1  g04855(.A0(new_n7290_), .A1(new_n7155_), .B0(new_n7291_), .Y(new_n7292_));
  AOI21X1  g04856(.A0(new_n7292_), .A1(new_n7153_), .B0(pi0074), .Y(new_n7293_));
  OAI21X1  g04857(.A0(new_n7293_), .A1(new_n7151_), .B0(new_n3123_), .Y(new_n7294_));
  AOI21X1  g04858(.A0(new_n7285_), .A1(new_n6814_), .B0(new_n7294_), .Y(new_n7295_));
  OAI21X1  g04859(.A0(new_n7295_), .A1(new_n7186_), .B0(new_n6800_), .Y(new_n7296_));
  AOI21X1  g04860(.A0(new_n7296_), .A1(new_n7185_), .B0(pi0954), .Y(new_n7297_));
  INVX1    g04861(.A(pi0033), .Y(new_n7298_));
  NAND2X1  g04862(.A(new_n7183_), .B(new_n7298_), .Y(new_n7299_));
  INVX1    g04863(.A(pi0954), .Y(po1110));
  AOI21X1  g04864(.A0(new_n7296_), .A1(pi0033), .B0(po1110), .Y(new_n7301_));
  AOI22X1  g04865(.A0(new_n7301_), .A1(new_n7299_), .B0(new_n7297_), .B1(new_n7184_), .Y(po0191));
  XOR2X1   g04866(.A(new_n6789_), .B(pi0197), .Y(new_n7303_));
  AND2X1   g04867(.A(new_n5023_), .B(pi0162), .Y(new_n7304_));
  AND3X1   g04868(.A(new_n7304_), .B(new_n6789_), .C(pi0197), .Y(new_n7305_));
  INVX1    g04869(.A(pi0162), .Y(new_n7306_));
  INVX1    g04870(.A(pi0197), .Y(new_n7307_));
  AOI21X1  g04871(.A0(new_n7307_), .A1(new_n7306_), .B0(new_n6791_), .Y(new_n7308_));
  NOR3X1   g04872(.A(new_n7308_), .B(new_n7305_), .C(new_n5048_), .Y(new_n7309_));
  MX2X1    g04873(.A(new_n7309_), .B(new_n7304_), .S0(new_n7303_), .Y(new_n7310_));
  AND3X1   g04874(.A(new_n7310_), .B(new_n6809_), .C(pi0232), .Y(new_n7311_));
  AND3X1   g04875(.A(new_n5023_), .B(pi0232), .C(pi0167), .Y(new_n7312_));
  AND2X1   g04876(.A(new_n7312_), .B(new_n6794_), .Y(new_n7313_));
  NOR3X1   g04877(.A(new_n7313_), .B(new_n7311_), .C(pi0074), .Y(new_n7314_));
  AND2X1   g04878(.A(new_n6795_), .B(pi0148), .Y(new_n7315_));
  NOR3X1   g04879(.A(new_n7315_), .B(new_n7311_), .C(new_n4982_), .Y(new_n7316_));
  NOR2X1   g04880(.A(new_n7316_), .B(new_n7314_), .Y(new_n7317_));
  AND3X1   g04881(.A(new_n7312_), .B(new_n6794_), .C(pi0038), .Y(new_n7318_));
  NOR4X1   g04882(.A(new_n7318_), .B(new_n7311_), .C(pi0074), .D(pi0054), .Y(new_n7319_));
  OR3X1    g04883(.A(new_n7319_), .B(new_n7316_), .C(new_n7314_), .Y(new_n7320_));
  AOI21X1  g04884(.A0(new_n7320_), .A1(new_n4975_), .B0(new_n3374_), .Y(new_n7321_));
  INVX1    g04885(.A(new_n7180_), .Y(new_n7322_));
  AOI21X1  g04886(.A0(new_n7322_), .A1(new_n4975_), .B0(new_n3374_), .Y(new_n7323_));
  OR2X1    g04887(.A(new_n7323_), .B(new_n7321_), .Y(new_n7324_));
  NOR2X1   g04888(.A(new_n7310_), .B(new_n2933_), .Y(new_n7325_));
  AND2X1   g04889(.A(pi0145), .B(pi0140), .Y(new_n7326_));
  NOR2X1   g04890(.A(pi0145), .B(pi0140), .Y(new_n7327_));
  NOR4X1   g04891(.A(new_n7327_), .B(new_n7326_), .C(new_n6803_), .D(new_n5048_), .Y(new_n7328_));
  OAI21X1  g04892(.A0(new_n7327_), .A1(new_n7326_), .B0(new_n6804_), .Y(new_n7329_));
  NAND2X1  g04893(.A(new_n7329_), .B(new_n2933_), .Y(new_n7330_));
  OAI21X1  g04894(.A0(new_n7330_), .A1(new_n7328_), .B0(pi0232), .Y(new_n7331_));
  NOR2X1   g04895(.A(new_n7331_), .B(new_n7325_), .Y(new_n7332_));
  AOI21X1  g04896(.A0(new_n3007_), .A1(new_n3073_), .B0(new_n7332_), .Y(new_n7333_));
  MX2X1    g04897(.A(pi0141), .B(pi0148), .S0(pi0299), .Y(new_n7334_));
  NAND3X1  g04898(.A(new_n7334_), .B(new_n5023_), .C(pi0232), .Y(new_n7335_));
  AOI21X1  g04899(.A0(new_n7335_), .A1(new_n6794_), .B0(new_n7333_), .Y(new_n7336_));
  OAI21X1  g04900(.A0(new_n7336_), .A1(new_n4982_), .B0(new_n3107_), .Y(new_n7337_));
  MX2X1    g04901(.A(pi0188), .B(pi0167), .S0(pi0299), .Y(new_n7338_));
  AND3X1   g04902(.A(new_n7338_), .B(new_n5023_), .C(pi0232), .Y(new_n7339_));
  NOR3X1   g04903(.A(new_n7339_), .B(pi0100), .C(pi0075), .Y(new_n7340_));
  OAI21X1  g04904(.A0(new_n7340_), .A1(new_n7333_), .B0(pi0054), .Y(new_n7341_));
  NOR2X1   g04905(.A(new_n7332_), .B(new_n3007_), .Y(new_n7342_));
  INVX1    g04906(.A(new_n7342_), .Y(new_n7343_));
  INVX1    g04907(.A(pi0144), .Y(new_n7344_));
  AND2X1   g04908(.A(new_n7010_), .B(new_n6989_), .Y(new_n7345_));
  AOI21X1  g04909(.A0(new_n6967_), .A1(pi0142), .B0(pi0140), .Y(new_n7346_));
  OAI21X1  g04910(.A0(new_n7345_), .A1(pi0142), .B0(new_n7346_), .Y(new_n7347_));
  OAI21X1  g04911(.A0(new_n7016_), .A1(new_n6938_), .B0(new_n2953_), .Y(new_n7348_));
  NAND3X1  g04912(.A(new_n7019_), .B(new_n6975_), .C(pi0142), .Y(new_n7349_));
  NAND3X1  g04913(.A(new_n7349_), .B(new_n7348_), .C(pi0140), .Y(new_n7350_));
  AOI21X1  g04914(.A0(new_n7350_), .A1(new_n7347_), .B0(pi0181), .Y(new_n7351_));
  AND2X1   g04915(.A(new_n7039_), .B(new_n2953_), .Y(new_n7352_));
  INVX1    g04916(.A(pi0140), .Y(new_n7353_));
  OAI21X1  g04917(.A0(new_n6985_), .A1(new_n2953_), .B0(new_n7353_), .Y(new_n7354_));
  NOR2X1   g04918(.A(new_n6980_), .B(new_n2953_), .Y(new_n7355_));
  AOI21X1  g04919(.A0(new_n7041_), .A1(new_n6989_), .B0(pi0142), .Y(new_n7356_));
  OR3X1    g04920(.A(new_n7356_), .B(new_n7355_), .C(new_n7353_), .Y(new_n7357_));
  OAI21X1  g04921(.A0(new_n7354_), .A1(new_n7352_), .B0(new_n7357_), .Y(new_n7358_));
  AND2X1   g04922(.A(new_n7358_), .B(pi0181), .Y(new_n7359_));
  NOR3X1   g04923(.A(new_n7359_), .B(new_n7351_), .C(new_n7344_), .Y(new_n7360_));
  AOI21X1  g04924(.A0(new_n7054_), .A1(new_n2953_), .B0(pi0140), .Y(new_n7361_));
  OAI21X1  g04925(.A0(new_n6951_), .A1(new_n2953_), .B0(new_n7361_), .Y(new_n7362_));
  AND3X1   g04926(.A(new_n7019_), .B(new_n7044_), .C(new_n2953_), .Y(new_n7363_));
  OAI21X1  g04927(.A0(new_n6963_), .A1(new_n2953_), .B0(pi0140), .Y(new_n7364_));
  OAI21X1  g04928(.A0(new_n7364_), .A1(new_n7363_), .B0(new_n7362_), .Y(new_n7365_));
  OR2X1    g04929(.A(new_n7031_), .B(pi0142), .Y(new_n7366_));
  AOI21X1  g04930(.A0(new_n7089_), .A1(new_n6948_), .B0(new_n5048_), .Y(new_n7367_));
  NOR2X1   g04931(.A(new_n7367_), .B(new_n2953_), .Y(new_n7368_));
  AOI21X1  g04932(.A0(new_n7368_), .A1(new_n7019_), .B0(pi0140), .Y(new_n7369_));
  NAND2X1  g04933(.A(new_n7034_), .B(new_n2953_), .Y(new_n7370_));
  AOI21X1  g04934(.A0(new_n7114_), .A1(new_n5023_), .B0(new_n2953_), .Y(new_n7371_));
  AOI21X1  g04935(.A0(new_n7371_), .A1(new_n7019_), .B0(new_n7353_), .Y(new_n7372_));
  AOI22X1  g04936(.A0(new_n7372_), .A1(new_n7370_), .B0(new_n7369_), .B1(new_n7366_), .Y(new_n7373_));
  OAI21X1  g04937(.A0(new_n7373_), .A1(pi0181), .B0(new_n7344_), .Y(new_n7374_));
  AOI21X1  g04938(.A0(new_n7365_), .A1(pi0181), .B0(new_n7374_), .Y(new_n7375_));
  NOR3X1   g04939(.A(new_n7375_), .B(new_n7360_), .C(pi0299), .Y(new_n7376_));
  INVX1    g04940(.A(pi0159), .Y(new_n7377_));
  AND2X1   g04941(.A(pi0299), .B(new_n7377_), .Y(new_n7378_));
  INVX1    g04942(.A(new_n7378_), .Y(new_n7379_));
  NOR3X1   g04943(.A(new_n7115_), .B(new_n7106_), .C(new_n2776_), .Y(new_n7380_));
  OAI21X1  g04944(.A0(new_n7111_), .A1(pi0146), .B0(new_n4611_), .Y(new_n7381_));
  AND3X1   g04945(.A(new_n7117_), .B(new_n6975_), .C(pi0146), .Y(new_n7382_));
  OAI21X1  g04946(.A0(new_n7062_), .A1(new_n7016_), .B0(new_n2776_), .Y(new_n7383_));
  NAND2X1  g04947(.A(new_n7383_), .B(pi0161), .Y(new_n7384_));
  OAI22X1  g04948(.A0(new_n7384_), .A1(new_n7382_), .B0(new_n7381_), .B1(new_n7380_), .Y(new_n7385_));
  AOI21X1  g04949(.A0(new_n7086_), .A1(new_n4611_), .B0(pi0146), .Y(new_n7386_));
  OAI21X1  g04950(.A0(new_n7083_), .A1(new_n4611_), .B0(new_n7386_), .Y(new_n7387_));
  OR2X1    g04951(.A(new_n7090_), .B(pi0161), .Y(new_n7388_));
  AOI21X1  g04952(.A0(new_n7092_), .A1(pi0161), .B0(new_n2776_), .Y(new_n7389_));
  OR2X1    g04953(.A(new_n7062_), .B(pi0162), .Y(new_n7390_));
  AOI21X1  g04954(.A0(new_n7389_), .A1(new_n7388_), .B0(new_n7390_), .Y(new_n7391_));
  AOI22X1  g04955(.A0(new_n7391_), .A1(new_n7387_), .B0(new_n7385_), .B1(pi0162), .Y(new_n7392_));
  NAND2X1  g04956(.A(new_n7073_), .B(new_n2776_), .Y(new_n7393_));
  AOI21X1  g04957(.A0(new_n7068_), .A1(pi0146), .B0(new_n4611_), .Y(new_n7394_));
  AND2X1   g04958(.A(new_n7394_), .B(new_n7393_), .Y(new_n7395_));
  OR2X1    g04959(.A(new_n7064_), .B(new_n2776_), .Y(new_n7396_));
  OAI21X1  g04960(.A0(new_n7077_), .A1(new_n7062_), .B0(new_n2776_), .Y(new_n7397_));
  AND3X1   g04961(.A(new_n7397_), .B(new_n7396_), .C(new_n4611_), .Y(new_n7398_));
  NOR3X1   g04962(.A(new_n7398_), .B(new_n7395_), .C(pi0162), .Y(new_n7399_));
  OR3X1    g04963(.A(new_n7106_), .B(new_n6999_), .C(pi0146), .Y(new_n7400_));
  OAI21X1  g04964(.A0(new_n7062_), .A1(new_n6962_), .B0(pi0146), .Y(new_n7401_));
  AND3X1   g04965(.A(new_n7401_), .B(new_n7400_), .C(new_n4611_), .Y(new_n7402_));
  OAI21X1  g04966(.A0(new_n7062_), .A1(new_n6979_), .B0(pi0146), .Y(new_n7403_));
  NOR3X1   g04967(.A(new_n7015_), .B(new_n6886_), .C(new_n5048_), .Y(new_n7404_));
  OAI21X1  g04968(.A0(new_n7062_), .A1(new_n7404_), .B0(new_n2776_), .Y(new_n7405_));
  AND3X1   g04969(.A(new_n7405_), .B(new_n7403_), .C(pi0161), .Y(new_n7406_));
  OR2X1    g04970(.A(new_n7406_), .B(new_n7306_), .Y(new_n7407_));
  AND2X1   g04971(.A(pi0299), .B(pi0159), .Y(new_n7408_));
  OAI21X1  g04972(.A0(new_n7407_), .A1(new_n7402_), .B0(new_n7408_), .Y(new_n7409_));
  OAI22X1  g04973(.A0(new_n7409_), .A1(new_n7399_), .B0(new_n7392_), .B1(new_n7379_), .Y(new_n7410_));
  OAI21X1  g04974(.A0(new_n7410_), .A1(new_n7376_), .B0(pi0232), .Y(new_n7411_));
  AOI21X1  g04975(.A0(new_n7411_), .A1(new_n7124_), .B0(new_n3060_), .Y(new_n7412_));
  OR2X1    g04976(.A(new_n6880_), .B(new_n7344_), .Y(new_n7413_));
  OR2X1    g04977(.A(pi0299), .B(pi0177), .Y(new_n7414_));
  NOR2X1   g04978(.A(new_n6850_), .B(pi0144), .Y(new_n7415_));
  AOI21X1  g04979(.A0(new_n7415_), .A1(new_n6875_), .B0(new_n7414_), .Y(new_n7416_));
  AOI21X1  g04980(.A0(new_n6853_), .A1(new_n6847_), .B0(new_n6849_), .Y(new_n7417_));
  AND2X1   g04981(.A(new_n2933_), .B(pi0177), .Y(new_n7418_));
  INVX1    g04982(.A(new_n7418_), .Y(new_n7419_));
  NOR2X1   g04983(.A(new_n7419_), .B(new_n7415_), .Y(new_n7420_));
  AOI22X1  g04984(.A0(new_n7420_), .A1(new_n7417_), .B0(new_n7416_), .B1(new_n7413_), .Y(new_n7421_));
  OR2X1    g04985(.A(new_n7421_), .B(new_n5215_), .Y(new_n7422_));
  OAI21X1  g04986(.A0(new_n6881_), .A1(pi0232), .B0(new_n7422_), .Y(new_n7423_));
  OR4X1    g04987(.A(new_n6861_), .B(new_n6835_), .C(new_n5048_), .D(pi0161), .Y(new_n7424_));
  AOI21X1  g04988(.A0(new_n7424_), .A1(new_n6860_), .B0(new_n7187_), .Y(new_n7425_));
  NOR2X1   g04989(.A(pi0155), .B(pi0038), .Y(new_n7426_));
  NAND3X1  g04990(.A(new_n7426_), .B(new_n6857_), .C(pi0299), .Y(new_n7427_));
  NAND2X1  g04991(.A(new_n6856_), .B(new_n6847_), .Y(new_n7428_));
  AOI21X1  g04992(.A0(new_n6868_), .A1(pi0161), .B0(new_n7428_), .Y(new_n7429_));
  AND2X1   g04993(.A(pi0155), .B(new_n2979_), .Y(new_n7430_));
  NAND3X1  g04994(.A(new_n7430_), .B(new_n6857_), .C(pi0299), .Y(new_n7431_));
  OAI22X1  g04995(.A0(new_n7431_), .A1(new_n7429_), .B0(new_n7427_), .B1(new_n7425_), .Y(new_n7432_));
  AOI22X1  g04996(.A0(new_n7432_), .A1(pi0232), .B0(new_n7423_), .B1(new_n2979_), .Y(new_n7433_));
  AOI21X1  g04997(.A0(new_n6829_), .A1(pi0188), .B0(pi0167), .Y(new_n7434_));
  INVX1    g04998(.A(new_n7434_), .Y(new_n7435_));
  INVX1    g04999(.A(pi0188), .Y(new_n7436_));
  INVX1    g05000(.A(pi0167), .Y(new_n7437_));
  NOR3X1   g05001(.A(new_n6823_), .B(new_n7436_), .C(new_n7437_), .Y(new_n7438_));
  AOI21X1  g05002(.A0(new_n6822_), .A1(new_n7436_), .B0(new_n7438_), .Y(new_n7439_));
  AOI21X1  g05003(.A0(new_n7439_), .A1(new_n7435_), .B0(new_n2979_), .Y(new_n7440_));
  NOR2X1   g05004(.A(new_n7440_), .B(pi0087), .Y(new_n7441_));
  OAI21X1  g05005(.A0(new_n7433_), .A1(new_n2939_), .B0(new_n7441_), .Y(new_n7442_));
  MX2X1    g05006(.A(new_n7339_), .B(new_n6834_), .S0(new_n2979_), .Y(new_n7443_));
  AOI21X1  g05007(.A0(new_n7443_), .A1(pi0087), .B0(pi0100), .Y(new_n7444_));
  OAI21X1  g05008(.A0(new_n7442_), .A1(new_n7412_), .B0(new_n7444_), .Y(new_n7445_));
  AOI21X1  g05009(.A0(new_n7445_), .A1(new_n7343_), .B0(new_n5295_), .Y(new_n7446_));
  NOR2X1   g05010(.A(new_n7332_), .B(new_n3073_), .Y(new_n7447_));
  INVX1    g05011(.A(new_n7447_), .Y(new_n7448_));
  INVX1    g05012(.A(pi0155), .Y(new_n7449_));
  INVX1    g05013(.A(pi0177), .Y(new_n7450_));
  MX2X1    g05014(.A(new_n7450_), .B(new_n7449_), .S0(pi0299), .Y(new_n7451_));
  AOI21X1  g05015(.A0(new_n7451_), .A1(new_n2979_), .B0(new_n6820_), .Y(new_n7452_));
  OR3X1    g05016(.A(new_n7452_), .B(new_n7142_), .C(new_n7141_), .Y(new_n7453_));
  AOI21X1  g05017(.A0(new_n7453_), .A1(new_n7443_), .B0(pi0100), .Y(new_n7454_));
  OAI21X1  g05018(.A0(new_n7454_), .A1(new_n7342_), .B0(new_n7138_), .Y(new_n7455_));
  NAND2X1  g05019(.A(new_n7455_), .B(new_n7448_), .Y(new_n7456_));
  OAI21X1  g05020(.A0(new_n7456_), .A1(new_n7446_), .B0(new_n3091_), .Y(new_n7457_));
  AOI21X1  g05021(.A0(new_n7457_), .A1(new_n7341_), .B0(pi0074), .Y(new_n7458_));
  NOR2X1   g05022(.A(new_n7316_), .B(new_n3107_), .Y(new_n7459_));
  NOR3X1   g05023(.A(new_n7313_), .B(new_n7311_), .C(new_n3091_), .Y(new_n7460_));
  NAND2X1  g05024(.A(new_n7179_), .B(new_n6794_), .Y(new_n7461_));
  NOR3X1   g05025(.A(new_n7318_), .B(new_n7311_), .C(pi0054), .Y(new_n7462_));
  AOI22X1  g05026(.A0(new_n7462_), .A1(new_n7461_), .B0(new_n3079_), .B1(new_n3091_), .Y(new_n7463_));
  AOI21X1  g05027(.A0(new_n7310_), .A1(pi0232), .B0(new_n3007_), .Y(new_n7464_));
  INVX1    g05028(.A(new_n7179_), .Y(new_n7465_));
  NOR3X1   g05029(.A(new_n7304_), .B(new_n7142_), .C(new_n7141_), .Y(new_n7466_));
  OAI21X1  g05030(.A0(new_n7466_), .A1(new_n7465_), .B0(new_n3007_), .Y(new_n7467_));
  NAND4X1  g05031(.A(new_n6843_), .B(new_n5215_), .C(new_n3131_), .D(new_n2939_), .Y(new_n7468_));
  AOI22X1  g05032(.A0(new_n7468_), .A1(new_n7467_), .B0(new_n7312_), .B1(pi0038), .Y(new_n7469_));
  OAI21X1  g05033(.A0(new_n7469_), .A1(new_n7464_), .B0(new_n3073_), .Y(new_n7470_));
  AOI21X1  g05034(.A0(new_n7310_), .A1(pi0232), .B0(new_n3073_), .Y(new_n7471_));
  NOR2X1   g05035(.A(new_n7471_), .B(pi0092), .Y(new_n7472_));
  AOI21X1  g05036(.A0(new_n7472_), .A1(new_n7470_), .B0(new_n7463_), .Y(new_n7473_));
  OAI21X1  g05037(.A0(new_n7473_), .A1(new_n7460_), .B0(new_n4982_), .Y(new_n7474_));
  AOI21X1  g05038(.A0(new_n7474_), .A1(new_n7459_), .B0(new_n4975_), .Y(new_n7475_));
  OAI21X1  g05039(.A0(new_n7458_), .A1(new_n7337_), .B0(new_n7475_), .Y(new_n7476_));
  AOI22X1  g05040(.A0(new_n7476_), .A1(new_n7324_), .B0(new_n7317_), .B1(new_n3374_), .Y(new_n7477_));
  NAND2X1  g05041(.A(new_n7477_), .B(new_n6783_), .Y(new_n7478_));
  AOI21X1  g05042(.A0(new_n7229_), .A1(new_n7227_), .B0(pi0146), .Y(new_n7479_));
  OAI21X1  g05043(.A0(new_n7252_), .A1(new_n2776_), .B0(new_n4611_), .Y(new_n7480_));
  NAND4X1  g05044(.A(new_n7238_), .B(new_n7229_), .C(pi0161), .D(new_n2776_), .Y(new_n7481_));
  OAI21X1  g05045(.A0(new_n7480_), .A1(new_n7479_), .B0(new_n7481_), .Y(new_n7482_));
  INVX1    g05046(.A(new_n7408_), .Y(new_n7483_));
  AOI21X1  g05047(.A0(new_n7255_), .A1(new_n7306_), .B0(new_n7483_), .Y(new_n7484_));
  OAI22X1  g05048(.A0(new_n7484_), .A1(new_n7378_), .B0(new_n5048_), .B1(new_n7306_), .Y(new_n7485_));
  NOR2X1   g05049(.A(new_n7221_), .B(new_n5175_), .Y(new_n7486_));
  INVX1    g05050(.A(new_n7486_), .Y(new_n7487_));
  AOI21X1  g05051(.A0(new_n7218_), .A1(new_n2776_), .B0(new_n7487_), .Y(new_n7488_));
  INVX1    g05052(.A(new_n7235_), .Y(new_n7489_));
  OAI21X1  g05053(.A0(new_n7489_), .A1(pi0146), .B0(new_n7263_), .Y(new_n7490_));
  OAI21X1  g05054(.A0(new_n5115_), .A1(new_n7377_), .B0(pi0299), .Y(new_n7491_));
  AOI21X1  g05055(.A0(new_n7490_), .A1(pi0161), .B0(new_n7491_), .Y(new_n7492_));
  OAI21X1  g05056(.A0(new_n7488_), .A1(pi0161), .B0(new_n7492_), .Y(new_n7493_));
  AOI22X1  g05057(.A0(new_n7493_), .A1(new_n7485_), .B0(new_n7482_), .B1(new_n7306_), .Y(new_n7494_));
  AOI21X1  g05058(.A0(new_n7252_), .A1(pi0142), .B0(pi0140), .Y(new_n7495_));
  OAI21X1  g05059(.A0(new_n7231_), .A1(pi0142), .B0(new_n7495_), .Y(new_n7496_));
  AND2X1   g05060(.A(new_n7218_), .B(new_n2953_), .Y(new_n7497_));
  OR3X1    g05061(.A(new_n7221_), .B(new_n5198_), .C(new_n7353_), .Y(new_n7498_));
  OAI21X1  g05062(.A0(new_n7498_), .A1(new_n7497_), .B0(new_n7496_), .Y(new_n7499_));
  AOI21X1  g05063(.A0(new_n7239_), .A1(new_n2953_), .B0(pi0140), .Y(new_n7500_));
  AOI21X1  g05064(.A0(new_n7235_), .A1(new_n2953_), .B0(new_n7353_), .Y(new_n7501_));
  AOI21X1  g05065(.A0(new_n7501_), .A1(new_n7246_), .B0(new_n7500_), .Y(new_n7502_));
  OAI22X1  g05066(.A0(new_n7502_), .A1(new_n7344_), .B0(new_n5023_), .B1(new_n7353_), .Y(new_n7503_));
  AOI21X1  g05067(.A0(new_n7499_), .A1(new_n7344_), .B0(new_n7503_), .Y(new_n7504_));
  OAI21X1  g05068(.A0(new_n7256_), .A1(new_n5204_), .B0(new_n2933_), .Y(new_n7505_));
  OAI21X1  g05069(.A0(new_n7505_), .A1(new_n7504_), .B0(pi0232), .Y(new_n7506_));
  OAI21X1  g05070(.A0(new_n7506_), .A1(new_n7494_), .B0(new_n3047_), .Y(new_n7507_));
  NOR2X1   g05071(.A(new_n7193_), .B(new_n4611_), .Y(new_n7508_));
  NOR2X1   g05072(.A(new_n5236_), .B(new_n6865_), .Y(new_n7509_));
  OAI21X1  g05073(.A0(new_n7509_), .A1(pi0161), .B0(new_n6856_), .Y(new_n7510_));
  OR2X1    g05074(.A(new_n7510_), .B(new_n7508_), .Y(new_n7511_));
  NAND3X1  g05075(.A(new_n7189_), .B(new_n6856_), .C(new_n4611_), .Y(new_n7512_));
  AOI22X1  g05076(.A0(new_n7512_), .A1(new_n7426_), .B0(new_n7511_), .B1(new_n7430_), .Y(new_n7513_));
  OAI21X1  g05077(.A0(new_n7205_), .A1(new_n7344_), .B0(new_n7418_), .Y(new_n7514_));
  AOI21X1  g05078(.A0(new_n7204_), .A1(new_n7344_), .B0(new_n7514_), .Y(new_n7515_));
  AND3X1   g05079(.A(new_n7200_), .B(new_n6848_), .C(new_n7344_), .Y(new_n7516_));
  OAI21X1  g05080(.A0(new_n7516_), .A1(new_n7414_), .B0(pi0232), .Y(new_n7517_));
  OAI21X1  g05081(.A0(new_n7517_), .A1(new_n7515_), .B0(new_n2979_), .Y(new_n7518_));
  OAI21X1  g05082(.A0(new_n7513_), .A1(new_n2933_), .B0(new_n7518_), .Y(new_n7519_));
  AOI21X1  g05083(.A0(new_n7519_), .A1(pi0039), .B0(new_n7440_), .Y(new_n7520_));
  AOI21X1  g05084(.A0(new_n7520_), .A1(new_n7507_), .B0(pi0100), .Y(new_n7521_));
  OAI21X1  g05085(.A0(new_n7521_), .A1(new_n7342_), .B0(new_n3131_), .Y(new_n7522_));
  INVX1    g05086(.A(new_n7339_), .Y(new_n7523_));
  OAI21X1  g05087(.A0(new_n7523_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n7524_));
  OAI21X1  g05088(.A0(new_n7332_), .A1(new_n3007_), .B0(new_n7524_), .Y(new_n7525_));
  AND2X1   g05089(.A(new_n7525_), .B(pi0087), .Y(new_n7526_));
  INVX1    g05090(.A(new_n7526_), .Y(new_n7527_));
  AOI21X1  g05091(.A0(new_n7527_), .A1(new_n7522_), .B0(new_n5295_), .Y(new_n7528_));
  NAND2X1  g05092(.A(new_n7338_), .B(pi0038), .Y(new_n7529_));
  OR3X1    g05093(.A(new_n7451_), .B(new_n3060_), .C(new_n2996_), .Y(new_n7530_));
  AOI21X1  g05094(.A0(new_n7530_), .A1(new_n7529_), .B0(new_n6820_), .Y(new_n7531_));
  OAI21X1  g05095(.A0(new_n7531_), .A1(pi0100), .B0(new_n7343_), .Y(new_n7532_));
  AOI21X1  g05096(.A0(new_n7532_), .A1(new_n3131_), .B0(new_n7526_), .Y(new_n7533_));
  OAI21X1  g05097(.A0(new_n7533_), .A1(new_n7279_), .B0(new_n7448_), .Y(new_n7534_));
  OAI21X1  g05098(.A0(new_n7534_), .A1(new_n7528_), .B0(new_n3091_), .Y(new_n7535_));
  AOI21X1  g05099(.A0(new_n7535_), .A1(new_n7341_), .B0(pi0074), .Y(new_n7536_));
  OR2X1    g05100(.A(new_n7311_), .B(pi0054), .Y(new_n7537_));
  NAND4X1  g05101(.A(new_n5023_), .B(pi0232), .C(pi0167), .D(pi0038), .Y(new_n7538_));
  NAND4X1  g05102(.A(new_n7280_), .B(new_n7259_), .C(pi0162), .D(new_n3079_), .Y(new_n7539_));
  OAI21X1  g05103(.A0(new_n7539_), .A1(new_n5431_), .B0(new_n7538_), .Y(new_n7540_));
  AOI21X1  g05104(.A0(new_n7540_), .A1(new_n6794_), .B0(new_n7537_), .Y(new_n7541_));
  OAI21X1  g05105(.A0(new_n7541_), .A1(new_n7460_), .B0(new_n4982_), .Y(new_n7542_));
  AOI21X1  g05106(.A0(new_n7542_), .A1(new_n7459_), .B0(new_n4975_), .Y(new_n7543_));
  OAI21X1  g05107(.A0(new_n7536_), .A1(new_n7337_), .B0(new_n7543_), .Y(new_n7544_));
  AOI22X1  g05108(.A0(new_n7544_), .A1(new_n7321_), .B0(new_n7317_), .B1(new_n3374_), .Y(new_n7545_));
  AOI22X1  g05109(.A0(new_n7545_), .A1(pi0034), .B0(po1110), .B1(new_n7298_), .Y(new_n7546_));
  OAI21X1  g05110(.A0(new_n6787_), .A1(pi0034), .B0(new_n7477_), .Y(new_n7547_));
  OR2X1    g05111(.A(pi0954), .B(pi0033), .Y(new_n7548_));
  NOR2X1   g05112(.A(new_n6787_), .B(pi0034), .Y(new_n7549_));
  AOI21X1  g05113(.A0(new_n7549_), .A1(new_n7545_), .B0(new_n7548_), .Y(new_n7550_));
  AOI22X1  g05114(.A0(new_n7550_), .A1(new_n7547_), .B0(new_n7546_), .B1(new_n7478_), .Y(po0192));
  OR2X1    g05115(.A(pi0074), .B(pi0055), .Y(new_n7552_));
  OR3X1    g05116(.A(new_n6773_), .B(new_n6772_), .C(pi0051), .Y(new_n7553_));
  OR2X1    g05117(.A(new_n5919_), .B(new_n5918_), .Y(new_n7554_));
  AND3X1   g05118(.A(new_n2759_), .B(pi0957), .C(new_n2701_), .Y(new_n7555_));
  NOR3X1   g05119(.A(new_n7555_), .B(new_n5928_), .C(new_n5077_), .Y(new_n7556_));
  NOR3X1   g05120(.A(new_n7556_), .B(new_n5082_), .C(new_n3035_), .Y(new_n7557_));
  AOI22X1  g05121(.A0(new_n5919_), .A1(pi0146), .B0(new_n5918_), .B1(pi0142), .Y(new_n7558_));
  AOI21X1  g05122(.A0(new_n7558_), .A1(new_n7554_), .B0(new_n7557_), .Y(new_n7559_));
  OAI22X1  g05123(.A0(new_n7559_), .A1(new_n5920_), .B0(new_n3035_), .B1(pi0137), .Y(new_n7560_));
  OR4X1    g05124(.A(new_n7557_), .B(new_n5920_), .C(new_n5082_), .D(new_n5072_), .Y(new_n7561_));
  AND2X1   g05125(.A(new_n7561_), .B(new_n7560_), .Y(new_n7562_));
  OAI22X1  g05126(.A0(new_n7562_), .A1(new_n6727_), .B0(new_n6725_), .B1(new_n2452_), .Y(new_n7563_));
  INVX1    g05127(.A(new_n5009_), .Y(new_n7564_));
  OAI21X1  g05128(.A0(new_n4991_), .A1(pi0090), .B0(new_n2516_), .Y(new_n7565_));
  AOI21X1  g05129(.A0(new_n7565_), .A1(new_n5003_), .B0(pi0035), .Y(new_n7566_));
  OAI21X1  g05130(.A0(new_n2706_), .A1(new_n2508_), .B0(new_n6759_), .Y(new_n7567_));
  OR2X1    g05131(.A(new_n7567_), .B(new_n7566_), .Y(new_n7568_));
  INVX1    g05132(.A(new_n2548_), .Y(new_n7569_));
  OR3X1    g05133(.A(new_n6732_), .B(pi0093), .C(new_n2455_), .Y(new_n7570_));
  OR4X1    g05134(.A(new_n7570_), .B(new_n2476_), .C(new_n7569_), .D(pi0841), .Y(new_n7571_));
  OAI21X1  g05135(.A0(new_n7568_), .A1(pi0032), .B0(new_n7571_), .Y(new_n7572_));
  AND3X1   g05136(.A(new_n7572_), .B(new_n7564_), .C(new_n2523_), .Y(new_n7573_));
  AND3X1   g05137(.A(new_n5907_), .B(new_n2703_), .C(pi1093), .Y(new_n7574_));
  AOI21X1  g05138(.A0(new_n7564_), .A1(new_n2452_), .B0(new_n6072_), .Y(new_n7575_));
  NOR2X1   g05139(.A(po0740), .B(pi0122), .Y(new_n7576_));
  AOI21X1  g05140(.A0(new_n7564_), .A1(new_n2452_), .B0(new_n6073_), .Y(new_n7577_));
  AOI22X1  g05141(.A0(new_n7577_), .A1(new_n7576_), .B0(new_n7575_), .B1(new_n7574_), .Y(new_n7578_));
  OAI21X1  g05142(.A0(new_n7566_), .A1(new_n7564_), .B0(new_n7578_), .Y(new_n7579_));
  OR4X1    g05143(.A(new_n6757_), .B(new_n6738_), .C(new_n2484_), .D(new_n2472_), .Y(new_n7580_));
  OR2X1    g05144(.A(new_n7567_), .B(new_n7250_), .Y(new_n7581_));
  AOI21X1  g05145(.A0(new_n7580_), .A1(new_n7566_), .B0(new_n7581_), .Y(new_n7582_));
  AND2X1   g05146(.A(new_n7582_), .B(new_n7579_), .Y(new_n7583_));
  NAND2X1  g05147(.A(new_n2527_), .B(pi0040), .Y(new_n7584_));
  NAND2X1  g05148(.A(new_n7228_), .B(pi1082), .Y(new_n7585_));
  AOI21X1  g05149(.A0(new_n7568_), .A1(new_n7584_), .B0(new_n7585_), .Y(new_n7586_));
  OR4X1    g05150(.A(new_n7586_), .B(new_n7583_), .C(new_n7573_), .D(pi0038), .Y(new_n7587_));
  OR2X1    g05151(.A(pi0100), .B(pi0039), .Y(new_n7588_));
  AOI21X1  g05152(.A0(new_n7553_), .A1(pi0038), .B0(new_n7588_), .Y(new_n7589_));
  AOI22X1  g05153(.A0(new_n7589_), .A1(new_n7587_), .B0(new_n7563_), .B1(new_n6723_), .Y(new_n7590_));
  NOR3X1   g05154(.A(po0840), .B(new_n6775_), .C(new_n2452_), .Y(new_n7591_));
  OAI21X1  g05155(.A0(new_n7591_), .A1(new_n6776_), .B0(new_n6778_), .Y(new_n7592_));
  OAI22X1  g05156(.A0(new_n7592_), .A1(new_n7553_), .B0(new_n7590_), .B1(new_n3080_), .Y(new_n7593_));
  AOI21X1  g05157(.A0(new_n7593_), .A1(new_n3079_), .B0(pi0054), .Y(new_n7594_));
  AOI21X1  g05158(.A0(new_n5809_), .A1(new_n5777_), .B0(new_n3091_), .Y(new_n7595_));
  OR4X1    g05159(.A(new_n7595_), .B(new_n7594_), .C(new_n7552_), .D(new_n4975_), .Y(new_n7596_));
  NOR4X1   g05160(.A(new_n7553_), .B(new_n4975_), .C(new_n3105_), .D(pi0055), .Y(new_n7597_));
  OAI21X1  g05161(.A0(new_n7597_), .A1(new_n3127_), .B0(new_n2436_), .Y(new_n7598_));
  AOI21X1  g05162(.A0(new_n7596_), .A1(new_n3127_), .B0(new_n7598_), .Y(po0193));
  NOR3X1   g05163(.A(new_n2561_), .B(new_n6914_), .C(pi0058), .Y(new_n7600_));
  OR4X1    g05164(.A(new_n6836_), .B(new_n2469_), .C(new_n2558_), .D(pi0065), .Y(new_n7601_));
  OR4X1    g05165(.A(pi0103), .B(pi0071), .C(pi0067), .D(new_n2640_), .Y(new_n7602_));
  NOR3X1   g05166(.A(new_n7602_), .B(new_n7601_), .C(pi0069), .Y(new_n7603_));
  NAND4X1  g05167(.A(new_n7603_), .B(new_n7600_), .C(new_n2643_), .D(new_n2594_), .Y(new_n7604_));
  OAI21X1  g05168(.A0(new_n5931_), .A1(pi0058), .B0(new_n7604_), .Y(new_n7605_));
  AND3X1   g05169(.A(new_n5168_), .B(new_n5010_), .C(new_n2483_), .Y(new_n7606_));
  AND3X1   g05170(.A(new_n5102_), .B(new_n3102_), .C(new_n2436_), .Y(new_n7607_));
  AND3X1   g05171(.A(new_n7607_), .B(new_n3208_), .C(new_n3079_), .Y(new_n7608_));
  AND2X1   g05172(.A(new_n7608_), .B(new_n7606_), .Y(new_n7609_));
  AND3X1   g05173(.A(new_n7609_), .B(new_n7605_), .C(po0740), .Y(po0194));
  NAND4X1  g05174(.A(new_n2984_), .B(new_n2531_), .C(new_n2939_), .D(pi0024), .Y(new_n7611_));
  OR4X1    g05175(.A(new_n2469_), .B(new_n2463_), .C(pi0104), .D(pi0071), .Y(new_n7612_));
  OR4X1    g05176(.A(pi0073), .B(pi0066), .C(pi0049), .D(pi0045), .Y(new_n7613_));
  INVX1    g05177(.A(pi0089), .Y(new_n7614_));
  OR2X1    g05178(.A(pi0065), .B(pi0048), .Y(new_n7615_));
  OR4X1    g05179(.A(new_n7615_), .B(new_n7614_), .C(pi0084), .D(pi0082), .Y(new_n7616_));
  NOR4X1   g05180(.A(new_n7616_), .B(new_n7613_), .C(new_n7612_), .D(new_n6906_), .Y(new_n7617_));
  AOI21X1  g05181(.A0(new_n7617_), .A1(pi0332), .B0(pi0064), .Y(new_n7618_));
  INVX1    g05182(.A(new_n5168_), .Y(new_n7619_));
  INVX1    g05183(.A(new_n6991_), .Y(new_n7620_));
  OR3X1    g05184(.A(new_n7620_), .B(new_n7619_), .C(new_n2504_), .Y(new_n7621_));
  OR4X1    g05185(.A(new_n2457_), .B(pi0841), .C(pi0102), .D(pi0039), .Y(new_n7622_));
  OR4X1    g05186(.A(new_n7622_), .B(new_n7621_), .C(new_n7618_), .D(new_n2526_), .Y(new_n7623_));
  NOR3X1   g05187(.A(new_n7623_), .B(new_n2586_), .C(pi0081), .Y(new_n7624_));
  AND2X1   g05188(.A(new_n6489_), .B(new_n3103_), .Y(new_n7625_));
  OAI21X1  g05189(.A0(new_n7624_), .A1(pi0038), .B0(new_n7625_), .Y(new_n7626_));
  AOI21X1  g05190(.A0(new_n7611_), .A1(pi0038), .B0(new_n7626_), .Y(po0196));
  AND3X1   g05191(.A(new_n6489_), .B(new_n3103_), .C(new_n2979_), .Y(new_n7628_));
  INVX1    g05192(.A(new_n7628_), .Y(new_n7629_));
  OR2X1    g05193(.A(new_n5225_), .B(pi0984), .Y(new_n7630_));
  AOI21X1  g05194(.A0(new_n7630_), .A1(pi0835), .B0(new_n5028_), .Y(new_n7631_));
  NOR3X1   g05195(.A(new_n7631_), .B(new_n5034_), .C(new_n5031_), .Y(new_n7632_));
  NOR2X1   g05196(.A(new_n5028_), .B(new_n5025_), .Y(new_n7633_));
  INVX1    g05197(.A(new_n7633_), .Y(new_n7634_));
  OR4X1    g05198(.A(new_n7634_), .B(new_n2985_), .C(new_n2536_), .D(pi0287), .Y(new_n7635_));
  AOI21X1  g05199(.A0(new_n7632_), .A1(pi1093), .B0(new_n7635_), .Y(new_n7636_));
  NAND2X1  g05200(.A(new_n7636_), .B(new_n2940_), .Y(new_n7637_));
  AND2X1   g05201(.A(new_n7632_), .B(new_n6255_), .Y(new_n7638_));
  NOR3X1   g05202(.A(new_n7638_), .B(new_n7635_), .C(new_n5042_), .Y(new_n7639_));
  NOR4X1   g05203(.A(new_n7631_), .B(new_n5043_), .C(new_n5034_), .D(new_n5031_), .Y(new_n7640_));
  NOR3X1   g05204(.A(new_n7640_), .B(new_n7635_), .C(new_n5041_), .Y(new_n7641_));
  NOR3X1   g05205(.A(new_n7641_), .B(new_n7639_), .C(pi0299), .Y(new_n7642_));
  AND2X1   g05206(.A(new_n7642_), .B(new_n7637_), .Y(new_n7643_));
  AND2X1   g05207(.A(new_n7636_), .B(new_n2934_), .Y(new_n7644_));
  NOR3X1   g05208(.A(new_n7638_), .B(new_n7635_), .C(new_n5059_), .Y(new_n7645_));
  NOR3X1   g05209(.A(new_n7640_), .B(new_n7635_), .C(new_n5058_), .Y(new_n7646_));
  OR4X1    g05210(.A(new_n7646_), .B(new_n7645_), .C(new_n7644_), .D(new_n2933_), .Y(new_n7647_));
  INVX1    g05211(.A(pi0786), .Y(new_n7648_));
  OR2X1    g05212(.A(pi1082), .B(new_n7648_), .Y(new_n7649_));
  NAND2X1  g05213(.A(new_n7649_), .B(new_n7647_), .Y(new_n7650_));
  AOI22X1  g05214(.A0(new_n5946_), .A1(new_n4889_), .B0(new_n5950_), .B1(new_n4769_), .Y(new_n7651_));
  OR4X1    g05215(.A(new_n7651_), .B(new_n7649_), .C(new_n5224_), .D(new_n5912_), .Y(new_n7652_));
  OAI21X1  g05216(.A0(new_n7650_), .A1(new_n7643_), .B0(new_n7652_), .Y(new_n7653_));
  NOR2X1   g05217(.A(pi0095), .B(pi0039), .Y(new_n7654_));
  AOI21X1  g05218(.A0(new_n2562_), .A1(pi0108), .B0(new_n2495_), .Y(new_n7655_));
  INVX1    g05219(.A(pi0097), .Y(new_n7656_));
  OR4X1    g05220(.A(new_n6748_), .B(new_n6745_), .C(new_n2460_), .D(pi0111), .Y(new_n7657_));
  OR4X1    g05221(.A(pi0084), .B(pi0081), .C(pi0066), .D(pi0064), .Y(new_n7658_));
  OR3X1    g05222(.A(new_n7658_), .B(pi0069), .C(pi0065), .Y(new_n7659_));
  OR4X1    g05223(.A(pi0082), .B(pi0068), .C(pi0049), .D(new_n2609_), .Y(new_n7660_));
  OR3X1    g05224(.A(new_n7660_), .B(pi0073), .C(pi0045), .Y(new_n7661_));
  NOR4X1   g05225(.A(new_n7661_), .B(new_n7659_), .C(new_n7657_), .D(new_n7612_), .Y(new_n7662_));
  AND3X1   g05226(.A(new_n2489_), .B(new_n6733_), .C(new_n2705_), .Y(new_n7663_));
  AND3X1   g05227(.A(new_n7663_), .B(new_n7662_), .C(new_n7656_), .Y(new_n7664_));
  OR2X1    g05228(.A(new_n2495_), .B(new_n2837_), .Y(new_n7665_));
  OAI21X1  g05229(.A0(new_n7665_), .A1(new_n2562_), .B0(new_n2550_), .Y(new_n7666_));
  AOI21X1  g05230(.A0(new_n7664_), .A1(new_n7655_), .B0(new_n7666_), .Y(new_n7667_));
  OAI21X1  g05231(.A0(po0740), .A1(pi0986), .B0(pi0252), .Y(new_n7668_));
  AND2X1   g05232(.A(new_n7668_), .B(pi0314), .Y(new_n7669_));
  NAND2X1  g05233(.A(new_n7669_), .B(new_n5000_), .Y(new_n7670_));
  OR4X1    g05234(.A(new_n2470_), .B(new_n2458_), .C(pi0081), .D(new_n2550_), .Y(new_n7671_));
  NAND3X1  g05235(.A(new_n7662_), .B(new_n2705_), .C(new_n2550_), .Y(new_n7672_));
  AND2X1   g05236(.A(new_n7672_), .B(new_n7671_), .Y(new_n7673_));
  OR3X1    g05237(.A(new_n7669_), .B(new_n2503_), .C(new_n4999_), .Y(new_n7674_));
  OAI22X1  g05238(.A0(new_n7674_), .A1(new_n7673_), .B0(new_n7670_), .B1(new_n7667_), .Y(new_n7675_));
  AOI21X1  g05239(.A0(new_n7675_), .A1(new_n2483_), .B0(pi0035), .Y(new_n7676_));
  AOI21X1  g05240(.A0(new_n5173_), .A1(pi0035), .B0(new_n2526_), .Y(new_n7677_));
  NAND2X1  g05241(.A(new_n7677_), .B(new_n2695_), .Y(new_n7678_));
  OAI22X1  g05242(.A0(new_n7678_), .A1(new_n7676_), .B0(new_n5174_), .B1(new_n7564_), .Y(new_n7679_));
  AOI22X1  g05243(.A0(new_n7679_), .A1(new_n7654_), .B0(new_n7653_), .B1(pi0039), .Y(new_n7680_));
  NOR2X1   g05244(.A(new_n7680_), .B(new_n7629_), .Y(po0197));
  INVX1    g05245(.A(pi1082), .Y(new_n7682_));
  OAI21X1  g05246(.A0(new_n2527_), .A1(new_n2529_), .B0(new_n7228_), .Y(new_n7683_));
  OR4X1    g05247(.A(new_n2502_), .B(new_n2457_), .C(new_n2580_), .D(pi0093), .Y(new_n7684_));
  OR4X1    g05248(.A(new_n7684_), .B(new_n6954_), .C(new_n2504_), .D(new_n2471_), .Y(new_n7685_));
  AND2X1   g05249(.A(new_n7685_), .B(new_n2529_), .Y(new_n7686_));
  OAI21X1  g05250(.A0(new_n7686_), .A1(new_n7683_), .B0(new_n7682_), .Y(new_n7687_));
  OAI21X1  g05251(.A0(new_n7685_), .A1(new_n7619_), .B0(pi1082), .Y(new_n7688_));
  AND3X1   g05252(.A(new_n7688_), .B(new_n7687_), .C(new_n7608_), .Y(po0198));
  NOR2X1   g05253(.A(pi0072), .B(pi0041), .Y(new_n7690_));
  NOR2X1   g05254(.A(new_n7690_), .B(new_n6278_), .Y(new_n7691_));
  INVX1    g05255(.A(new_n6278_), .Y(new_n7692_));
  AOI21X1  g05256(.A0(new_n7690_), .A1(new_n2704_), .B0(new_n7692_), .Y(new_n7693_));
  INVX1    g05257(.A(new_n7693_), .Y(new_n7694_));
  INVX1    g05258(.A(new_n6239_), .Y(new_n7695_));
  AND2X1   g05259(.A(new_n5907_), .B(pi1093), .Y(new_n7696_));
  INVX1    g05260(.A(new_n7696_), .Y(new_n7697_));
  OR4X1    g05261(.A(new_n2985_), .B(new_n2536_), .C(pi0101), .D(pi0044), .Y(new_n7698_));
  NOR2X1   g05262(.A(new_n7698_), .B(new_n7697_), .Y(new_n7699_));
  INVX1    g05263(.A(new_n7699_), .Y(new_n7700_));
  OAI21X1  g05264(.A0(new_n7700_), .A1(new_n7695_), .B0(pi0041), .Y(new_n7701_));
  OAI21X1  g05265(.A0(new_n2530_), .A1(pi0041), .B0(new_n2703_), .Y(new_n7702_));
  INVX1    g05266(.A(pi0099), .Y(new_n7703_));
  NAND2X1  g05267(.A(new_n5081_), .B(new_n7703_), .Y(new_n7704_));
  AOI21X1  g05268(.A0(pi0101), .A1(new_n2530_), .B0(pi0041), .Y(new_n7705_));
  INVX1    g05269(.A(new_n7705_), .Y(new_n7706_));
  NAND3X1  g05270(.A(new_n2479_), .B(new_n2477_), .C(new_n5777_), .Y(new_n7707_));
  NAND2X1  g05271(.A(new_n5168_), .B(pi0252), .Y(new_n7708_));
  OR4X1    g05272(.A(new_n7708_), .B(new_n7707_), .C(new_n7697_), .D(pi0044), .Y(new_n7709_));
  NOR2X1   g05273(.A(new_n7709_), .B(new_n7706_), .Y(new_n7710_));
  AOI21X1  g05274(.A0(new_n7710_), .A1(new_n7704_), .B0(new_n7702_), .Y(new_n7711_));
  AOI21X1  g05275(.A0(new_n7711_), .A1(new_n7701_), .B0(new_n7694_), .Y(new_n7712_));
  OAI21X1  g05276(.A0(new_n7712_), .A1(new_n7691_), .B0(new_n2939_), .Y(new_n7713_));
  NOR3X1   g05277(.A(pi0468), .B(pi0332), .C(pi0189), .Y(new_n7714_));
  AND2X1   g05278(.A(new_n7714_), .B(pi0144), .Y(new_n7715_));
  AOI21X1  g05279(.A0(new_n7715_), .A1(new_n6851_), .B0(pi0299), .Y(new_n7716_));
  NOR3X1   g05280(.A(pi0468), .B(pi0332), .C(pi0166), .Y(new_n7717_));
  AND3X1   g05281(.A(new_n7717_), .B(pi0161), .C(new_n3193_), .Y(new_n7718_));
  OAI21X1  g05282(.A0(new_n7718_), .A1(new_n5918_), .B0(pi0232), .Y(new_n7719_));
  NOR2X1   g05283(.A(new_n7719_), .B(new_n7716_), .Y(new_n7720_));
  INVX1    g05284(.A(new_n7720_), .Y(new_n7721_));
  AOI21X1  g05285(.A0(new_n7721_), .A1(new_n2530_), .B0(new_n2939_), .Y(new_n7722_));
  NOR2X1   g05286(.A(new_n7722_), .B(new_n5778_), .Y(new_n7723_));
  NOR2X1   g05287(.A(new_n7690_), .B(pi0039), .Y(new_n7724_));
  NOR2X1   g05288(.A(new_n7724_), .B(new_n7722_), .Y(new_n7725_));
  INVX1    g05289(.A(new_n7725_), .Y(new_n7726_));
  OAI21X1  g05290(.A0(new_n7726_), .A1(new_n3087_), .B0(pi0075), .Y(new_n7727_));
  AOI21X1  g05291(.A0(new_n7723_), .A1(new_n7713_), .B0(new_n7727_), .Y(new_n7728_));
  OR4X1    g05292(.A(new_n5907_), .B(new_n5900_), .C(new_n5881_), .D(pi0096), .Y(new_n7729_));
  AND3X1   g05293(.A(new_n7729_), .B(new_n5909_), .C(new_n5032_), .Y(new_n7730_));
  NOR3X1   g05294(.A(new_n5900_), .B(new_n5881_), .C(pi0096), .Y(new_n7731_));
  AND2X1   g05295(.A(new_n2544_), .B(pi0091), .Y(new_n7732_));
  NOR2X1   g05296(.A(new_n5896_), .B(new_n2732_), .Y(new_n7733_));
  AOI22X1  g05297(.A0(new_n7733_), .A1(new_n2727_), .B0(new_n7732_), .B1(new_n5777_), .Y(new_n7734_));
  OAI21X1  g05298(.A0(new_n7734_), .A1(new_n2502_), .B0(new_n5887_), .Y(new_n7735_));
  AOI21X1  g05299(.A0(new_n7735_), .A1(new_n5885_), .B0(pi0051), .Y(new_n7736_));
  OAI21X1  g05300(.A0(new_n7736_), .A1(new_n2847_), .B0(new_n2513_), .Y(new_n7737_));
  NOR4X1   g05301(.A(new_n5908_), .B(new_n5905_), .C(new_n7619_), .D(pi0072), .Y(new_n7738_));
  AOI22X1  g05302(.A0(new_n7738_), .A1(new_n7737_), .B0(new_n5908_), .B1(new_n7731_), .Y(new_n7739_));
  AND2X1   g05303(.A(new_n7739_), .B(pi1093), .Y(new_n7740_));
  OR4X1    g05304(.A(new_n7740_), .B(new_n7730_), .C(pi0101), .D(pi0044), .Y(new_n7741_));
  NAND2X1  g05305(.A(new_n7741_), .B(pi0041), .Y(new_n7742_));
  INVX1    g05306(.A(pi0101), .Y(new_n7743_));
  OR3X1    g05307(.A(new_n5907_), .B(new_n7731_), .C(pi0072), .Y(new_n7744_));
  OR2X1    g05308(.A(new_n5905_), .B(new_n7619_), .Y(new_n7745_));
  AND2X1   g05309(.A(new_n5907_), .B(new_n2530_), .Y(new_n7746_));
  OAI21X1  g05310(.A0(new_n7745_), .A1(new_n5903_), .B0(new_n7746_), .Y(new_n7747_));
  AND3X1   g05311(.A(new_n7747_), .B(new_n7744_), .C(new_n5032_), .Y(new_n7748_));
  AOI21X1  g05312(.A0(new_n7739_), .A1(new_n2530_), .B0(new_n5032_), .Y(new_n7749_));
  NOR2X1   g05313(.A(new_n7749_), .B(new_n7748_), .Y(new_n7750_));
  MX2X1    g05314(.A(new_n7750_), .B(new_n2530_), .S0(pi0044), .Y(new_n7751_));
  AOI21X1  g05315(.A0(new_n7751_), .A1(new_n7743_), .B0(new_n7706_), .Y(new_n7752_));
  NOR2X1   g05316(.A(new_n7752_), .B(new_n2704_), .Y(new_n7753_));
  NOR3X1   g05317(.A(new_n7748_), .B(new_n7731_), .C(pi0072), .Y(new_n7754_));
  MX2X1    g05318(.A(new_n7754_), .B(new_n2530_), .S0(pi0044), .Y(new_n7755_));
  AOI21X1  g05319(.A0(new_n7755_), .A1(new_n7743_), .B0(new_n7706_), .Y(new_n7756_));
  INVX1    g05320(.A(pi0041), .Y(new_n7757_));
  NOR2X1   g05321(.A(new_n7731_), .B(new_n5032_), .Y(new_n7758_));
  NOR4X1   g05322(.A(new_n7758_), .B(new_n7730_), .C(pi0101), .D(pi0044), .Y(new_n7759_));
  OAI21X1  g05323(.A0(new_n7759_), .A1(new_n7757_), .B0(new_n2704_), .Y(new_n7760_));
  OAI21X1  g05324(.A0(new_n7760_), .A1(new_n7756_), .B0(pi0228), .Y(new_n7761_));
  AOI21X1  g05325(.A0(new_n7753_), .A1(new_n7742_), .B0(new_n7761_), .Y(new_n7762_));
  INVX1    g05326(.A(new_n2479_), .Y(new_n7763_));
  INVX1    g05327(.A(pi0480), .Y(new_n7764_));
  AND2X1   g05328(.A(pi0949), .B(new_n7764_), .Y(new_n7765_));
  NAND4X1  g05329(.A(new_n2569_), .B(new_n2497_), .C(pi0094), .D(new_n2566_), .Y(new_n7766_));
  OR3X1    g05330(.A(new_n7766_), .B(new_n7765_), .C(new_n7763_), .Y(new_n7767_));
  INVX1    g05331(.A(new_n2570_), .Y(new_n7768_));
  OR4X1    g05332(.A(pi0109), .B(pi0108), .C(pi0097), .D(pi0046), .Y(new_n7769_));
  OAI21X1  g05333(.A0(new_n7769_), .A1(new_n7768_), .B0(new_n2547_), .Y(new_n7770_));
  NAND2X1  g05334(.A(new_n7765_), .B(new_n2479_), .Y(new_n7771_));
  NOR4X1   g05335(.A(new_n7771_), .B(new_n2549_), .C(new_n4999_), .D(pi0047), .Y(new_n7772_));
  INVX1    g05336(.A(pi0959), .Y(new_n7773_));
  NAND2X1  g05337(.A(new_n7773_), .B(pi0901), .Y(new_n7774_));
  AOI21X1  g05338(.A0(new_n7772_), .A1(new_n7770_), .B0(new_n7774_), .Y(new_n7775_));
  NOR4X1   g05339(.A(new_n2475_), .B(new_n7569_), .C(new_n2547_), .D(pi0109), .Y(new_n7776_));
  INVX1    g05340(.A(new_n7776_), .Y(new_n7777_));
  OAI21X1  g05341(.A0(new_n7777_), .A1(new_n7771_), .B0(new_n7774_), .Y(new_n7778_));
  INVX1    g05342(.A(pi0250), .Y(new_n7779_));
  AND2X1   g05343(.A(pi0252), .B(new_n7779_), .Y(new_n7780_));
  NAND3X1  g05344(.A(new_n7780_), .B(new_n7778_), .C(new_n5168_), .Y(new_n7781_));
  AOI21X1  g05345(.A0(new_n7775_), .A1(new_n7767_), .B0(new_n7781_), .Y(new_n7782_));
  INVX1    g05346(.A(new_n7780_), .Y(new_n7783_));
  AND2X1   g05347(.A(new_n7783_), .B(new_n7765_), .Y(new_n7784_));
  AND3X1   g05348(.A(new_n7784_), .B(new_n7776_), .C(new_n7606_), .Y(new_n7785_));
  AOI21X1  g05349(.A0(new_n7782_), .A1(new_n2530_), .B0(new_n7785_), .Y(new_n7786_));
  NOR3X1   g05350(.A(new_n7786_), .B(pi0101), .C(pi0044), .Y(new_n7787_));
  NOR2X1   g05351(.A(new_n7787_), .B(new_n7757_), .Y(new_n7788_));
  NOR4X1   g05352(.A(new_n7780_), .B(new_n7777_), .C(new_n7771_), .D(new_n7619_), .Y(new_n7789_));
  NOR3X1   g05353(.A(new_n7789_), .B(new_n7782_), .C(pi0072), .Y(new_n7790_));
  MX2X1    g05354(.A(new_n7790_), .B(new_n2530_), .S0(pi0044), .Y(new_n7791_));
  AOI21X1  g05355(.A0(new_n7791_), .A1(new_n7743_), .B0(new_n7706_), .Y(new_n7792_));
  OAI21X1  g05356(.A0(new_n7792_), .A1(new_n7788_), .B0(new_n2793_), .Y(new_n7793_));
  NAND2X1  g05357(.A(new_n7793_), .B(new_n2939_), .Y(new_n7794_));
  INVX1    g05358(.A(pi0287), .Y(new_n7795_));
  NOR3X1   g05359(.A(new_n2985_), .B(new_n2536_), .C(new_n7795_), .Y(new_n7796_));
  MX2X1    g05360(.A(new_n7796_), .B(new_n2530_), .S0(new_n7721_), .Y(new_n7797_));
  AOI21X1  g05361(.A0(new_n7797_), .A1(pi0039), .B0(new_n3252_), .Y(new_n7798_));
  OAI21X1  g05362(.A0(new_n7794_), .A1(new_n7762_), .B0(new_n7798_), .Y(new_n7799_));
  INVX1    g05363(.A(new_n7722_), .Y(new_n7800_));
  NAND4X1  g05364(.A(new_n5168_), .B(new_n2479_), .C(new_n2477_), .D(new_n5078_), .Y(new_n7801_));
  NOR2X1   g05365(.A(new_n7801_), .B(new_n7706_), .Y(new_n7802_));
  AOI21X1  g05366(.A0(pi0072), .A1(new_n7757_), .B0(new_n7802_), .Y(new_n7803_));
  AOI21X1  g05367(.A0(new_n7697_), .A1(new_n2530_), .B0(new_n7803_), .Y(new_n7804_));
  NAND2X1  g05368(.A(new_n7704_), .B(new_n2703_), .Y(new_n7805_));
  AOI22X1  g05369(.A0(new_n7805_), .A1(new_n7702_), .B0(new_n7804_), .B1(new_n7704_), .Y(new_n7806_));
  OAI21X1  g05370(.A0(new_n7699_), .A1(new_n7757_), .B0(new_n7806_), .Y(new_n7807_));
  AOI21X1  g05371(.A0(new_n7807_), .A1(new_n7693_), .B0(new_n7691_), .Y(new_n7808_));
  OAI21X1  g05372(.A0(new_n7808_), .A1(pi0039), .B0(new_n7800_), .Y(new_n7809_));
  OAI21X1  g05373(.A0(new_n7725_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n7810_));
  AOI21X1  g05374(.A0(new_n7809_), .A1(new_n5074_), .B0(new_n7810_), .Y(new_n7811_));
  NAND2X1  g05375(.A(new_n7698_), .B(pi0041), .Y(new_n7812_));
  NAND3X1  g05376(.A(new_n7812_), .B(new_n7803_), .C(pi0228), .Y(new_n7813_));
  AOI21X1  g05377(.A0(new_n7690_), .A1(new_n2793_), .B0(new_n3132_), .Y(new_n7814_));
  NOR3X1   g05378(.A(new_n7690_), .B(new_n3251_), .C(pi0039), .Y(new_n7815_));
  OR3X1    g05379(.A(new_n7815_), .B(new_n7722_), .C(new_n3131_), .Y(new_n7816_));
  AOI21X1  g05380(.A0(new_n7814_), .A1(new_n7813_), .B0(new_n7816_), .Y(new_n7817_));
  OR2X1    g05381(.A(new_n7817_), .B(pi0075), .Y(new_n7818_));
  AOI21X1  g05382(.A0(new_n7811_), .A1(new_n7799_), .B0(new_n7818_), .Y(new_n7819_));
  OAI21X1  g05383(.A0(new_n7819_), .A1(new_n7728_), .B0(new_n5880_), .Y(new_n7820_));
  AOI21X1  g05384(.A0(new_n7726_), .A1(new_n6295_), .B0(po1038), .Y(new_n7821_));
  AND2X1   g05385(.A(pi0232), .B(pi0039), .Y(new_n7822_));
  OR3X1    g05386(.A(new_n7724_), .B(new_n6489_), .C(pi0072), .Y(new_n7823_));
  AOI21X1  g05387(.A0(new_n7822_), .A1(new_n7718_), .B0(new_n7823_), .Y(new_n7824_));
  AOI21X1  g05388(.A0(new_n7821_), .A1(new_n7820_), .B0(new_n7824_), .Y(po0199));
  AND2X1   g05389(.A(pi0208), .B(pi0207), .Y(new_n7826_));
  INVX1    g05390(.A(new_n7826_), .Y(new_n7827_));
  INVX1    g05391(.A(pi0115), .Y(new_n7828_));
  AND2X1   g05392(.A(new_n2703_), .B(new_n7828_), .Y(new_n7829_));
  INVX1    g05393(.A(pi0114), .Y(new_n7830_));
  NAND2X1  g05394(.A(pi0116), .B(pi0072), .Y(new_n7831_));
  NOR2X1   g05395(.A(pi0099), .B(pi0041), .Y(new_n7832_));
  INVX1    g05396(.A(new_n7832_), .Y(new_n7833_));
  AOI22X1  g05397(.A0(new_n7752_), .A1(new_n7703_), .B0(new_n7833_), .B1(pi0072), .Y(new_n7834_));
  MX2X1    g05398(.A(new_n7834_), .B(new_n2530_), .S0(pi0113), .Y(new_n7835_));
  OAI21X1  g05399(.A0(new_n7835_), .A1(pi0116), .B0(new_n7831_), .Y(new_n7836_));
  AND3X1   g05400(.A(new_n7836_), .B(new_n7830_), .C(pi0042), .Y(new_n7837_));
  AND2X1   g05401(.A(new_n2530_), .B(pi0042), .Y(new_n7838_));
  OR2X1    g05402(.A(pi0116), .B(pi0113), .Y(new_n7839_));
  NOR3X1   g05403(.A(new_n7741_), .B(new_n7839_), .C(new_n7833_), .Y(new_n7840_));
  OAI22X1  g05404(.A0(new_n7840_), .A1(pi0042), .B0(new_n7838_), .B1(new_n7830_), .Y(new_n7841_));
  OAI21X1  g05405(.A0(new_n7841_), .A1(new_n7837_), .B0(new_n7829_), .Y(new_n7842_));
  AOI21X1  g05406(.A0(new_n2530_), .A1(pi0042), .B0(new_n7830_), .Y(new_n7843_));
  NOR2X1   g05407(.A(new_n2703_), .B(pi0115), .Y(new_n7844_));
  AOI22X1  g05408(.A0(new_n7756_), .A1(new_n7703_), .B0(new_n7833_), .B1(pi0072), .Y(new_n7845_));
  MX2X1    g05409(.A(new_n7845_), .B(new_n2530_), .S0(pi0113), .Y(new_n7846_));
  MX2X1    g05410(.A(new_n7846_), .B(new_n2530_), .S0(pi0116), .Y(new_n7847_));
  INVX1    g05411(.A(pi0042), .Y(new_n7848_));
  OR3X1    g05412(.A(new_n7758_), .B(new_n7730_), .C(pi0044), .Y(new_n7849_));
  NOR4X1   g05413(.A(new_n7849_), .B(new_n7839_), .C(new_n7833_), .D(pi0101), .Y(new_n7850_));
  AND2X1   g05414(.A(new_n7850_), .B(new_n7848_), .Y(new_n7851_));
  OR2X1    g05415(.A(new_n7851_), .B(pi0114), .Y(new_n7852_));
  AOI21X1  g05416(.A0(new_n7847_), .A1(pi0042), .B0(new_n7852_), .Y(new_n7853_));
  OAI21X1  g05417(.A0(new_n7853_), .A1(new_n7843_), .B0(new_n7844_), .Y(new_n7854_));
  OAI21X1  g05418(.A0(pi0072), .A1(new_n7848_), .B0(pi0115), .Y(new_n7855_));
  AND3X1   g05419(.A(new_n7855_), .B(new_n7854_), .C(pi0228), .Y(new_n7856_));
  AOI22X1  g05420(.A0(new_n7792_), .A1(new_n7703_), .B0(new_n7833_), .B1(pi0072), .Y(new_n7857_));
  MX2X1    g05421(.A(new_n7857_), .B(new_n2530_), .S0(pi0113), .Y(new_n7858_));
  MX2X1    g05422(.A(new_n7858_), .B(new_n2530_), .S0(pi0116), .Y(new_n7859_));
  OR3X1    g05423(.A(new_n7859_), .B(pi0114), .C(new_n7848_), .Y(new_n7860_));
  INVX1    g05424(.A(pi0113), .Y(new_n7861_));
  INVX1    g05425(.A(pi0116), .Y(new_n7862_));
  NOR4X1   g05426(.A(new_n7786_), .B(new_n7833_), .C(pi0101), .D(pi0044), .Y(new_n7863_));
  AND3X1   g05427(.A(new_n7863_), .B(new_n7862_), .C(new_n7861_), .Y(new_n7864_));
  INVX1    g05428(.A(new_n7864_), .Y(new_n7865_));
  AOI21X1  g05429(.A0(new_n7865_), .A1(new_n7848_), .B0(new_n7843_), .Y(new_n7866_));
  AOI21X1  g05430(.A0(new_n7866_), .A1(new_n7860_), .B0(pi0115), .Y(new_n7867_));
  NAND2X1  g05431(.A(new_n7855_), .B(new_n2793_), .Y(new_n7868_));
  OAI21X1  g05432(.A0(new_n7868_), .A1(new_n7867_), .B0(new_n2939_), .Y(new_n7869_));
  AOI21X1  g05433(.A0(new_n7856_), .A1(new_n7842_), .B0(new_n7869_), .Y(new_n7870_));
  INVX1    g05434(.A(pi0199), .Y(new_n7871_));
  INVX1    g05435(.A(pi0189), .Y(new_n7872_));
  INVX1    g05436(.A(new_n7714_), .Y(new_n7873_));
  NOR4X1   g05437(.A(new_n5048_), .B(new_n2985_), .C(new_n2536_), .D(new_n7795_), .Y(new_n7874_));
  AOI22X1  g05438(.A0(new_n7874_), .A1(new_n7872_), .B0(new_n7873_), .B1(new_n2530_), .Y(new_n7875_));
  AND2X1   g05439(.A(new_n2933_), .B(pi0232), .Y(new_n7876_));
  OAI21X1  g05440(.A0(new_n7875_), .A1(new_n7871_), .B0(new_n7876_), .Y(new_n7877_));
  AOI21X1  g05441(.A0(new_n6819_), .A1(new_n4459_), .B0(pi0072), .Y(new_n7878_));
  OR3X1    g05442(.A(new_n7878_), .B(new_n2933_), .C(new_n5215_), .Y(new_n7879_));
  AOI21X1  g05443(.A0(new_n7796_), .A1(new_n7717_), .B0(new_n7879_), .Y(new_n7880_));
  AOI21X1  g05444(.A0(pi0199), .A1(new_n2530_), .B0(pi0232), .Y(new_n7881_));
  OAI21X1  g05445(.A0(pi0232), .A1(new_n2530_), .B0(pi0299), .Y(new_n7882_));
  AND2X1   g05446(.A(new_n7882_), .B(new_n7881_), .Y(new_n7883_));
  NOR2X1   g05447(.A(new_n7883_), .B(new_n7880_), .Y(new_n7884_));
  AOI21X1  g05448(.A0(new_n7884_), .A1(new_n7877_), .B0(new_n2939_), .Y(new_n7885_));
  OAI21X1  g05449(.A0(new_n7885_), .A1(new_n7870_), .B0(new_n3251_), .Y(new_n7886_));
  INVX1    g05450(.A(new_n7838_), .Y(new_n7887_));
  INVX1    g05451(.A(new_n7829_), .Y(new_n7888_));
  AOI21X1  g05452(.A0(new_n7838_), .A1(new_n7888_), .B0(new_n7692_), .Y(new_n7889_));
  NOR4X1   g05453(.A(new_n7843_), .B(new_n5922_), .C(new_n2702_), .D(pi0115), .Y(new_n7890_));
  NOR3X1   g05454(.A(pi0052), .B(pi0043), .C(pi0042), .Y(new_n7891_));
  NOR4X1   g05455(.A(new_n7698_), .B(new_n7697_), .C(new_n7839_), .D(new_n7833_), .Y(new_n7892_));
  INVX1    g05456(.A(new_n7892_), .Y(new_n7893_));
  NOR4X1   g05457(.A(new_n7893_), .B(new_n7891_), .C(pi0114), .D(pi0042), .Y(new_n7894_));
  INVX1    g05458(.A(new_n5079_), .Y(new_n7895_));
  NOR3X1   g05459(.A(new_n7801_), .B(new_n7839_), .C(new_n7895_), .Y(new_n7896_));
  INVX1    g05460(.A(new_n7896_), .Y(new_n7897_));
  OAI21X1  g05461(.A0(new_n7897_), .A1(new_n7697_), .B0(new_n2530_), .Y(new_n7898_));
  OAI21X1  g05462(.A0(new_n7898_), .A1(new_n7848_), .B0(new_n7830_), .Y(new_n7899_));
  OAI21X1  g05463(.A0(new_n7899_), .A1(new_n7894_), .B0(new_n7890_), .Y(new_n7900_));
  AOI22X1  g05464(.A0(new_n7900_), .A1(new_n7889_), .B0(new_n7887_), .B1(new_n7692_), .Y(new_n7901_));
  NOR2X1   g05465(.A(new_n7881_), .B(pi0299), .Y(new_n7902_));
  NOR3X1   g05466(.A(new_n7714_), .B(new_n7871_), .C(pi0072), .Y(new_n7903_));
  OAI21X1  g05467(.A0(new_n7903_), .A1(new_n5215_), .B0(new_n7902_), .Y(new_n7904_));
  AOI21X1  g05468(.A0(new_n7878_), .A1(pi0299), .B0(new_n2939_), .Y(new_n7905_));
  AND2X1   g05469(.A(new_n7905_), .B(new_n7904_), .Y(new_n7906_));
  INVX1    g05470(.A(new_n7906_), .Y(new_n7907_));
  OAI21X1  g05471(.A0(new_n7901_), .A1(pi0039), .B0(new_n7907_), .Y(new_n7908_));
  AOI22X1  g05472(.A0(new_n7905_), .A1(new_n7904_), .B0(new_n7887_), .B1(new_n2939_), .Y(new_n7909_));
  OAI21X1  g05473(.A0(new_n7909_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n7910_));
  AOI21X1  g05474(.A0(new_n7908_), .A1(new_n5074_), .B0(new_n7910_), .Y(new_n7911_));
  OR4X1    g05475(.A(new_n7698_), .B(new_n7839_), .C(new_n7833_), .D(new_n2793_), .Y(new_n7912_));
  OR4X1    g05476(.A(new_n7912_), .B(pi0115), .C(pi0114), .D(pi0042), .Y(new_n7913_));
  OR3X1    g05477(.A(new_n7801_), .B(new_n7895_), .C(new_n2793_), .Y(new_n7914_));
  OAI21X1  g05478(.A0(new_n7914_), .A1(new_n5080_), .B0(new_n7838_), .Y(new_n7915_));
  AND3X1   g05479(.A(new_n7915_), .B(new_n7913_), .C(new_n3064_), .Y(new_n7916_));
  OAI21X1  g05480(.A0(pi0072), .A1(new_n7848_), .B0(new_n2939_), .Y(new_n7917_));
  OAI21X1  g05481(.A0(new_n7917_), .A1(new_n3251_), .B0(pi0087), .Y(new_n7918_));
  OR2X1    g05482(.A(new_n7918_), .B(new_n7916_), .Y(new_n7919_));
  OAI21X1  g05483(.A0(new_n7919_), .A1(new_n7906_), .B0(new_n3073_), .Y(new_n7920_));
  AOI21X1  g05484(.A0(new_n7911_), .A1(new_n7886_), .B0(new_n7920_), .Y(new_n7921_));
  INVX1    g05485(.A(new_n7889_), .Y(new_n7922_));
  NOR4X1   g05486(.A(new_n7893_), .B(new_n7695_), .C(new_n7891_), .D(pi0114), .Y(new_n7923_));
  NAND2X1  g05487(.A(new_n7923_), .B(new_n7848_), .Y(new_n7924_));
  OR4X1    g05488(.A(new_n7709_), .B(new_n7895_), .C(pi0116), .D(pi0113), .Y(new_n7925_));
  AOI21X1  g05489(.A0(new_n7925_), .A1(new_n7838_), .B0(pi0114), .Y(new_n7926_));
  NAND2X1  g05490(.A(new_n7926_), .B(new_n7924_), .Y(new_n7927_));
  AOI21X1  g05491(.A0(new_n7927_), .A1(new_n7890_), .B0(new_n7922_), .Y(new_n7928_));
  OAI21X1  g05492(.A0(new_n7838_), .A1(new_n6278_), .B0(new_n3087_), .Y(new_n7929_));
  AOI21X1  g05493(.A0(new_n7838_), .A1(new_n5778_), .B0(pi0039), .Y(new_n7930_));
  OAI21X1  g05494(.A0(new_n7929_), .A1(new_n7928_), .B0(new_n7930_), .Y(new_n7931_));
  AOI21X1  g05495(.A0(new_n7931_), .A1(new_n7907_), .B0(new_n3073_), .Y(new_n7932_));
  OR2X1    g05496(.A(new_n7932_), .B(new_n6295_), .Y(new_n7933_));
  OAI21X1  g05497(.A0(new_n7933_), .A1(new_n7921_), .B0(new_n7827_), .Y(new_n7934_));
  AOI21X1  g05498(.A0(pi0200), .A1(new_n2530_), .B0(pi0232), .Y(new_n7935_));
  NOR2X1   g05499(.A(new_n7935_), .B(pi0299), .Y(new_n7936_));
  INVX1    g05500(.A(pi0200), .Y(new_n7937_));
  NOR3X1   g05501(.A(new_n7714_), .B(new_n7937_), .C(pi0072), .Y(new_n7938_));
  OAI21X1  g05502(.A0(new_n7938_), .A1(new_n5215_), .B0(new_n7936_), .Y(new_n7939_));
  AND3X1   g05503(.A(new_n7939_), .B(new_n7904_), .C(pi0039), .Y(new_n7940_));
  AOI21X1  g05504(.A0(new_n7887_), .A1(new_n2939_), .B0(new_n7940_), .Y(new_n7941_));
  AOI21X1  g05505(.A0(new_n7941_), .A1(new_n6295_), .B0(new_n7827_), .Y(new_n7942_));
  OAI21X1  g05506(.A0(new_n7875_), .A1(new_n7871_), .B0(pi0232), .Y(new_n7943_));
  NOR2X1   g05507(.A(new_n7875_), .B(new_n7937_), .Y(new_n7944_));
  OR3X1    g05508(.A(new_n7944_), .B(new_n7943_), .C(pi0299), .Y(new_n7945_));
  OR2X1    g05509(.A(new_n7937_), .B(pi0072), .Y(new_n7946_));
  AOI21X1  g05510(.A0(new_n7946_), .A1(new_n7883_), .B0(new_n7880_), .Y(new_n7947_));
  AOI21X1  g05511(.A0(new_n7947_), .A1(new_n7945_), .B0(new_n2939_), .Y(new_n7948_));
  OAI21X1  g05512(.A0(new_n7948_), .A1(new_n7870_), .B0(new_n3251_), .Y(new_n7949_));
  AND2X1   g05513(.A(new_n7939_), .B(pi0039), .Y(new_n7950_));
  AND2X1   g05514(.A(new_n7950_), .B(new_n7906_), .Y(new_n7951_));
  INVX1    g05515(.A(new_n7951_), .Y(new_n7952_));
  OAI21X1  g05516(.A0(new_n7901_), .A1(pi0039), .B0(new_n7952_), .Y(new_n7953_));
  OAI21X1  g05517(.A0(new_n7941_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n7954_));
  AOI22X1  g05518(.A0(new_n7954_), .A1(new_n7910_), .B0(new_n7953_), .B1(new_n5074_), .Y(new_n7955_));
  OR2X1    g05519(.A(new_n7951_), .B(new_n7918_), .Y(new_n7956_));
  OAI21X1  g05520(.A0(new_n7956_), .A1(new_n7916_), .B0(new_n3073_), .Y(new_n7957_));
  AOI21X1  g05521(.A0(new_n7955_), .A1(new_n7949_), .B0(new_n7957_), .Y(new_n7958_));
  AOI21X1  g05522(.A0(new_n7952_), .A1(new_n7931_), .B0(new_n3073_), .Y(new_n7959_));
  OR2X1    g05523(.A(new_n7959_), .B(new_n6295_), .Y(new_n7960_));
  OAI21X1  g05524(.A0(new_n7960_), .A1(new_n7958_), .B0(new_n7942_), .Y(new_n7961_));
  AND3X1   g05525(.A(pi0214), .B(pi0212), .C(pi0211), .Y(new_n7962_));
  NOR2X1   g05526(.A(new_n7962_), .B(pi0219), .Y(new_n7963_));
  AND2X1   g05527(.A(new_n7909_), .B(new_n6295_), .Y(new_n7964_));
  OR2X1    g05528(.A(new_n7964_), .B(new_n7963_), .Y(new_n7965_));
  AOI21X1  g05529(.A0(new_n7961_), .A1(new_n7934_), .B0(new_n7965_), .Y(new_n7966_));
  INVX1    g05530(.A(new_n7963_), .Y(new_n7967_));
  AOI21X1  g05531(.A0(new_n7943_), .A1(new_n7902_), .B0(new_n2939_), .Y(new_n7968_));
  OAI21X1  g05532(.A0(new_n7968_), .A1(new_n7870_), .B0(new_n3251_), .Y(new_n7969_));
  AND2X1   g05533(.A(new_n7904_), .B(pi0039), .Y(new_n7970_));
  INVX1    g05534(.A(new_n7970_), .Y(new_n7971_));
  OAI21X1  g05535(.A0(new_n7901_), .A1(pi0039), .B0(new_n7971_), .Y(new_n7972_));
  AOI21X1  g05536(.A0(new_n7887_), .A1(new_n2939_), .B0(new_n7970_), .Y(new_n7973_));
  OAI21X1  g05537(.A0(new_n7973_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n7974_));
  AOI21X1  g05538(.A0(new_n7972_), .A1(new_n5074_), .B0(new_n7974_), .Y(new_n7975_));
  OAI21X1  g05539(.A0(new_n7970_), .A1(new_n7919_), .B0(new_n3073_), .Y(new_n7976_));
  AOI21X1  g05540(.A0(new_n7975_), .A1(new_n7969_), .B0(new_n7976_), .Y(new_n7977_));
  AOI21X1  g05541(.A0(new_n7971_), .A1(new_n7931_), .B0(new_n3073_), .Y(new_n7978_));
  OR3X1    g05542(.A(new_n7978_), .B(new_n7977_), .C(new_n6295_), .Y(new_n7979_));
  AOI21X1  g05543(.A0(new_n7973_), .A1(new_n6295_), .B0(new_n7826_), .Y(new_n7980_));
  OAI22X1  g05544(.A0(new_n7944_), .A1(new_n7943_), .B0(new_n7936_), .B1(new_n7902_), .Y(new_n7981_));
  AND2X1   g05545(.A(new_n7981_), .B(pi0039), .Y(new_n7982_));
  OAI21X1  g05546(.A0(new_n7982_), .A1(new_n7870_), .B0(new_n3251_), .Y(new_n7983_));
  INVX1    g05547(.A(new_n7940_), .Y(new_n7984_));
  OAI21X1  g05548(.A0(new_n7901_), .A1(pi0039), .B0(new_n7984_), .Y(new_n7985_));
  AOI21X1  g05549(.A0(new_n7985_), .A1(new_n5074_), .B0(new_n7954_), .Y(new_n7986_));
  OAI21X1  g05550(.A0(new_n7940_), .A1(new_n7919_), .B0(new_n3073_), .Y(new_n7987_));
  AOI21X1  g05551(.A0(new_n7986_), .A1(new_n7983_), .B0(new_n7987_), .Y(new_n7988_));
  AOI21X1  g05552(.A0(new_n7984_), .A1(new_n7931_), .B0(new_n3073_), .Y(new_n7989_));
  OR3X1    g05553(.A(new_n7989_), .B(new_n7988_), .C(new_n6295_), .Y(new_n7990_));
  AOI22X1  g05554(.A0(new_n7990_), .A1(new_n7942_), .B0(new_n7980_), .B1(new_n7979_), .Y(new_n7991_));
  OAI21X1  g05555(.A0(new_n7991_), .A1(new_n7967_), .B0(new_n6489_), .Y(new_n7992_));
  AOI21X1  g05556(.A0(new_n7967_), .A1(new_n7878_), .B0(new_n2939_), .Y(new_n7993_));
  OAI21X1  g05557(.A0(new_n5103_), .A1(pi0057), .B0(new_n7917_), .Y(new_n7994_));
  OAI22X1  g05558(.A0(new_n7994_), .A1(new_n7993_), .B0(new_n7992_), .B1(new_n7966_), .Y(po0200));
  AND2X1   g05559(.A(pi0214), .B(pi0212), .Y(new_n7996_));
  NOR2X1   g05560(.A(pi0219), .B(pi0211), .Y(new_n7997_));
  MX2X1    g05561(.A(pi0211), .B(new_n7997_), .S0(new_n7996_), .Y(new_n7998_));
  INVX1    g05562(.A(new_n7859_), .Y(new_n7999_));
  INVX1    g05563(.A(new_n7847_), .Y(new_n8000_));
  MX2X1    g05564(.A(new_n8000_), .B(new_n7836_), .S0(new_n2703_), .Y(new_n8001_));
  MX2X1    g05565(.A(new_n8001_), .B(new_n7999_), .S0(new_n2793_), .Y(new_n8002_));
  NOR3X1   g05566(.A(pi0115), .B(pi0114), .C(pi0042), .Y(new_n8003_));
  NAND3X1  g05567(.A(new_n8003_), .B(new_n8002_), .C(pi0043), .Y(new_n8004_));
  INVX1    g05568(.A(pi0043), .Y(new_n8005_));
  NAND2X1  g05569(.A(new_n7759_), .B(new_n7832_), .Y(new_n8006_));
  NAND2X1  g05570(.A(new_n8006_), .B(new_n2704_), .Y(new_n8007_));
  OAI21X1  g05571(.A0(new_n7741_), .A1(new_n7833_), .B0(new_n2703_), .Y(new_n8008_));
  NAND2X1  g05572(.A(new_n8008_), .B(new_n8007_), .Y(new_n8009_));
  NOR2X1   g05573(.A(new_n8009_), .B(new_n7839_), .Y(new_n8010_));
  MX2X1    g05574(.A(new_n8010_), .B(new_n7864_), .S0(new_n2793_), .Y(new_n8011_));
  INVX1    g05575(.A(new_n8011_), .Y(new_n8012_));
  AOI21X1  g05576(.A0(new_n2530_), .A1(pi0043), .B0(new_n8003_), .Y(new_n8013_));
  AOI21X1  g05577(.A0(new_n8012_), .A1(new_n8005_), .B0(new_n8013_), .Y(new_n8014_));
  AOI21X1  g05578(.A0(new_n8014_), .A1(new_n8004_), .B0(pi0039), .Y(new_n8015_));
  OAI21X1  g05579(.A0(new_n7875_), .A1(new_n7937_), .B0(pi0232), .Y(new_n8016_));
  AOI21X1  g05580(.A0(new_n8016_), .A1(new_n7936_), .B0(new_n2939_), .Y(new_n8017_));
  OAI21X1  g05581(.A0(new_n8017_), .A1(new_n8015_), .B0(new_n3251_), .Y(new_n8018_));
  AND2X1   g05582(.A(new_n2530_), .B(pi0043), .Y(new_n8019_));
  INVX1    g05583(.A(new_n8019_), .Y(new_n8020_));
  OAI21X1  g05584(.A0(new_n5920_), .A1(new_n2793_), .B0(new_n8020_), .Y(new_n8021_));
  AND2X1   g05585(.A(new_n8003_), .B(new_n2703_), .Y(new_n8022_));
  INVX1    g05586(.A(new_n8022_), .Y(new_n8023_));
  AOI21X1  g05587(.A0(new_n8023_), .A1(new_n8019_), .B0(new_n7692_), .Y(new_n8024_));
  AND2X1   g05588(.A(pi0052), .B(new_n8005_), .Y(new_n8025_));
  NOR2X1   g05589(.A(new_n7898_), .B(new_n8005_), .Y(new_n8026_));
  AOI21X1  g05590(.A0(new_n8025_), .A1(new_n7892_), .B0(new_n8026_), .Y(new_n8027_));
  OAI21X1  g05591(.A0(new_n8027_), .A1(new_n8023_), .B0(new_n8024_), .Y(new_n8028_));
  AOI21X1  g05592(.A0(new_n8028_), .A1(new_n8021_), .B0(pi0039), .Y(new_n8029_));
  OAI21X1  g05593(.A0(new_n8029_), .A1(new_n7950_), .B0(new_n5074_), .Y(new_n8030_));
  AOI21X1  g05594(.A0(new_n2530_), .A1(pi0043), .B0(pi0039), .Y(new_n8031_));
  AOI21X1  g05595(.A0(new_n7939_), .A1(pi0039), .B0(new_n8031_), .Y(new_n8032_));
  OR2X1    g05596(.A(new_n8032_), .B(new_n2979_), .Y(new_n8033_));
  AND3X1   g05597(.A(new_n8033_), .B(new_n8030_), .C(new_n3131_), .Y(new_n8034_));
  NOR3X1   g05598(.A(new_n7698_), .B(new_n7839_), .C(new_n7833_), .Y(new_n8035_));
  OR2X1    g05599(.A(new_n8035_), .B(pi0043), .Y(new_n8036_));
  OAI21X1  g05600(.A0(new_n7896_), .A1(pi0072), .B0(pi0043), .Y(new_n8037_));
  AND2X1   g05601(.A(new_n8003_), .B(pi0228), .Y(new_n8038_));
  AND3X1   g05602(.A(new_n8038_), .B(new_n8037_), .C(new_n8036_), .Y(new_n8039_));
  OAI21X1  g05603(.A0(new_n8038_), .A1(new_n8020_), .B0(new_n3064_), .Y(new_n8040_));
  AOI21X1  g05604(.A0(new_n8031_), .A1(new_n3252_), .B0(new_n3131_), .Y(new_n8041_));
  OAI21X1  g05605(.A0(new_n8040_), .A1(new_n8039_), .B0(new_n8041_), .Y(new_n8042_));
  OAI21X1  g05606(.A0(new_n8042_), .A1(new_n7950_), .B0(new_n3073_), .Y(new_n8043_));
  AOI21X1  g05607(.A0(new_n8034_), .A1(new_n8018_), .B0(new_n8043_), .Y(new_n8044_));
  AND3X1   g05608(.A(new_n7925_), .B(new_n2530_), .C(pi0043), .Y(new_n8045_));
  AND3X1   g05609(.A(new_n8025_), .B(new_n7892_), .C(new_n6239_), .Y(new_n8046_));
  OAI21X1  g05610(.A0(new_n8046_), .A1(new_n8045_), .B0(new_n8022_), .Y(new_n8047_));
  AOI22X1  g05611(.A0(new_n8047_), .A1(new_n8024_), .B0(new_n8020_), .B1(new_n7692_), .Y(new_n8048_));
  OAI21X1  g05612(.A0(new_n8048_), .A1(pi0039), .B0(new_n3087_), .Y(new_n8049_));
  OR2X1    g05613(.A(new_n8031_), .B(new_n3087_), .Y(new_n8050_));
  AOI21X1  g05614(.A0(new_n8050_), .A1(new_n8049_), .B0(new_n7950_), .Y(new_n8051_));
  OAI21X1  g05615(.A0(new_n8051_), .A1(new_n3073_), .B0(new_n5880_), .Y(new_n8052_));
  AOI21X1  g05616(.A0(new_n8032_), .A1(new_n6295_), .B0(new_n7826_), .Y(new_n8053_));
  OAI21X1  g05617(.A0(new_n8052_), .A1(new_n8044_), .B0(new_n8053_), .Y(new_n8054_));
  NOR2X1   g05618(.A(pi0200), .B(pi0199), .Y(new_n8055_));
  OAI21X1  g05619(.A0(new_n8055_), .A1(pi0299), .B0(new_n2530_), .Y(new_n8056_));
  AOI21X1  g05620(.A0(new_n8056_), .A1(new_n5215_), .B0(pi0299), .Y(new_n8057_));
  INVX1    g05621(.A(new_n8055_), .Y(new_n8058_));
  OAI21X1  g05622(.A0(new_n8058_), .A1(new_n7875_), .B0(pi0232), .Y(new_n8059_));
  AOI21X1  g05623(.A0(new_n8059_), .A1(new_n8057_), .B0(new_n2939_), .Y(new_n8060_));
  OAI21X1  g05624(.A0(new_n8060_), .A1(new_n8015_), .B0(new_n3251_), .Y(new_n8061_));
  AND2X1   g05625(.A(new_n8056_), .B(new_n5215_), .Y(new_n8062_));
  NOR4X1   g05626(.A(new_n7714_), .B(pi0200), .C(pi0199), .D(pi0072), .Y(new_n8063_));
  NOR2X1   g05627(.A(new_n8063_), .B(new_n5215_), .Y(new_n8064_));
  NOR3X1   g05628(.A(new_n8064_), .B(new_n8062_), .C(pi0299), .Y(new_n8065_));
  NOR2X1   g05629(.A(new_n8065_), .B(new_n2939_), .Y(new_n8066_));
  OR2X1    g05630(.A(new_n8066_), .B(new_n8029_), .Y(new_n8067_));
  MX2X1    g05631(.A(new_n8065_), .B(new_n8019_), .S0(new_n2939_), .Y(new_n8068_));
  OAI21X1  g05632(.A0(new_n8068_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n8069_));
  AOI21X1  g05633(.A0(new_n8067_), .A1(new_n5074_), .B0(new_n8069_), .Y(new_n8070_));
  NOR2X1   g05634(.A(new_n8068_), .B(new_n3111_), .Y(new_n8071_));
  OAI21X1  g05635(.A0(new_n8071_), .A1(new_n8042_), .B0(new_n3073_), .Y(new_n8072_));
  AOI21X1  g05636(.A0(new_n8070_), .A1(new_n8061_), .B0(new_n8072_), .Y(new_n8073_));
  AOI21X1  g05637(.A0(new_n8050_), .A1(new_n8049_), .B0(new_n8066_), .Y(new_n8074_));
  OAI21X1  g05638(.A0(new_n8074_), .A1(new_n3073_), .B0(new_n5880_), .Y(new_n8075_));
  AOI21X1  g05639(.A0(new_n8068_), .A1(new_n6295_), .B0(new_n7827_), .Y(new_n8076_));
  OAI21X1  g05640(.A0(new_n8075_), .A1(new_n8073_), .B0(new_n8076_), .Y(new_n8077_));
  AOI21X1  g05641(.A0(new_n8077_), .A1(new_n8054_), .B0(new_n7998_), .Y(new_n8078_));
  INVX1    g05642(.A(new_n7998_), .Y(new_n8079_));
  OAI21X1  g05643(.A0(new_n7875_), .A1(new_n7937_), .B0(new_n7876_), .Y(new_n8080_));
  AOI21X1  g05644(.A0(new_n7935_), .A1(new_n7882_), .B0(new_n7880_), .Y(new_n8081_));
  AOI21X1  g05645(.A0(new_n8081_), .A1(new_n8080_), .B0(new_n2939_), .Y(new_n8082_));
  OAI21X1  g05646(.A0(new_n8082_), .A1(new_n8015_), .B0(new_n3251_), .Y(new_n8083_));
  AND2X1   g05647(.A(new_n7939_), .B(new_n7905_), .Y(new_n8084_));
  OAI21X1  g05648(.A0(new_n8084_), .A1(new_n8029_), .B0(new_n5074_), .Y(new_n8085_));
  AOI21X1  g05649(.A0(new_n7939_), .A1(new_n7905_), .B0(new_n8031_), .Y(new_n8086_));
  OR2X1    g05650(.A(new_n8086_), .B(new_n2979_), .Y(new_n8087_));
  AND3X1   g05651(.A(new_n8087_), .B(new_n8085_), .C(new_n3131_), .Y(new_n8088_));
  OAI21X1  g05652(.A0(new_n8084_), .A1(new_n8042_), .B0(new_n3073_), .Y(new_n8089_));
  AOI21X1  g05653(.A0(new_n8088_), .A1(new_n8083_), .B0(new_n8089_), .Y(new_n8090_));
  AOI21X1  g05654(.A0(new_n8050_), .A1(new_n8049_), .B0(new_n8084_), .Y(new_n8091_));
  OAI21X1  g05655(.A0(new_n8091_), .A1(new_n3073_), .B0(new_n5880_), .Y(new_n8092_));
  AOI21X1  g05656(.A0(new_n8086_), .A1(new_n6295_), .B0(new_n7826_), .Y(new_n8093_));
  OAI21X1  g05657(.A0(new_n8092_), .A1(new_n8090_), .B0(new_n8093_), .Y(new_n8094_));
  OAI21X1  g05658(.A0(new_n8058_), .A1(new_n7875_), .B0(new_n7876_), .Y(new_n8095_));
  NOR2X1   g05659(.A(new_n8062_), .B(new_n7880_), .Y(new_n8096_));
  AOI21X1  g05660(.A0(new_n8096_), .A1(new_n8095_), .B0(new_n2939_), .Y(new_n8097_));
  OAI21X1  g05661(.A0(new_n8097_), .A1(new_n8015_), .B0(new_n3251_), .Y(new_n8098_));
  AND2X1   g05662(.A(new_n7878_), .B(pi0299), .Y(new_n8099_));
  NOR3X1   g05663(.A(new_n8065_), .B(new_n8099_), .C(new_n2939_), .Y(new_n8100_));
  OAI21X1  g05664(.A0(new_n8100_), .A1(new_n8029_), .B0(new_n5074_), .Y(new_n8101_));
  OAI21X1  g05665(.A0(new_n8100_), .A1(new_n8031_), .B0(pi0038), .Y(new_n8102_));
  AND3X1   g05666(.A(new_n8102_), .B(new_n8101_), .C(new_n3131_), .Y(new_n8103_));
  OAI21X1  g05667(.A0(new_n8100_), .A1(new_n8042_), .B0(new_n3073_), .Y(new_n8104_));
  AOI21X1  g05668(.A0(new_n8103_), .A1(new_n8098_), .B0(new_n8104_), .Y(new_n8105_));
  AOI21X1  g05669(.A0(new_n8050_), .A1(new_n8049_), .B0(new_n8100_), .Y(new_n8106_));
  OAI21X1  g05670(.A0(new_n8106_), .A1(new_n3073_), .B0(new_n5880_), .Y(new_n8107_));
  OR3X1    g05671(.A(new_n8100_), .B(new_n8031_), .C(new_n5880_), .Y(new_n8108_));
  AND2X1   g05672(.A(new_n8108_), .B(new_n7826_), .Y(new_n8109_));
  OAI21X1  g05673(.A0(new_n8107_), .A1(new_n8105_), .B0(new_n8109_), .Y(new_n8110_));
  AOI21X1  g05674(.A0(new_n8110_), .A1(new_n8094_), .B0(new_n8079_), .Y(new_n8111_));
  OR3X1    g05675(.A(new_n8111_), .B(new_n8078_), .C(po1038), .Y(new_n8112_));
  AOI21X1  g05676(.A0(new_n7998_), .A1(new_n7878_), .B0(new_n2939_), .Y(new_n8113_));
  OR2X1    g05677(.A(new_n8031_), .B(new_n6489_), .Y(new_n8114_));
  OAI21X1  g05678(.A0(new_n8114_), .A1(new_n8113_), .B0(new_n8112_), .Y(po0201));
  AND2X1   g05679(.A(new_n2530_), .B(pi0044), .Y(new_n8116_));
  INVX1    g05680(.A(new_n8116_), .Y(new_n8117_));
  AOI21X1  g05681(.A0(new_n8117_), .A1(new_n7692_), .B0(pi0039), .Y(new_n8118_));
  AOI21X1  g05682(.A0(new_n8116_), .A1(new_n2704_), .B0(new_n7692_), .Y(new_n8119_));
  AND2X1   g05683(.A(pi0072), .B(pi0044), .Y(new_n8120_));
  NOR4X1   g05684(.A(new_n8120_), .B(new_n5082_), .C(new_n5922_), .D(new_n2702_), .Y(new_n8121_));
  INVX1    g05685(.A(new_n8121_), .Y(new_n8122_));
  OR3X1    g05686(.A(new_n7708_), .B(new_n7707_), .C(new_n7697_), .Y(new_n8123_));
  NOR4X1   g05687(.A(new_n7697_), .B(new_n2985_), .C(new_n2536_), .D(pi0044), .Y(new_n8124_));
  AND2X1   g05688(.A(new_n8124_), .B(new_n6239_), .Y(new_n8125_));
  AOI21X1  g05689(.A0(new_n8123_), .A1(pi0044), .B0(new_n8125_), .Y(new_n8126_));
  OAI21X1  g05690(.A0(new_n8126_), .A1(new_n8122_), .B0(new_n8119_), .Y(new_n8127_));
  AND3X1   g05691(.A(new_n5920_), .B(new_n2530_), .C(pi0039), .Y(new_n8128_));
  AOI21X1  g05692(.A0(new_n8127_), .A1(new_n8118_), .B0(new_n8128_), .Y(new_n8129_));
  AOI21X1  g05693(.A0(new_n5920_), .A1(new_n2530_), .B0(new_n2939_), .Y(new_n8130_));
  AOI21X1  g05694(.A0(new_n8117_), .A1(new_n2939_), .B0(new_n8130_), .Y(new_n8131_));
  AOI21X1  g05695(.A0(new_n8131_), .A1(new_n5778_), .B0(new_n3073_), .Y(new_n8132_));
  OAI21X1  g05696(.A0(new_n8129_), .A1(new_n5778_), .B0(new_n8132_), .Y(new_n8133_));
  OR3X1    g05697(.A(new_n7740_), .B(new_n7730_), .C(pi0044), .Y(new_n8134_));
  OR3X1    g05698(.A(new_n7749_), .B(new_n7748_), .C(new_n5078_), .Y(new_n8135_));
  AND3X1   g05699(.A(new_n8135_), .B(new_n8134_), .C(new_n2703_), .Y(new_n8136_));
  OR4X1    g05700(.A(new_n7748_), .B(new_n7731_), .C(pi0072), .D(new_n5078_), .Y(new_n8137_));
  AND3X1   g05701(.A(new_n8137_), .B(new_n7849_), .C(new_n2704_), .Y(new_n8138_));
  OAI21X1  g05702(.A0(new_n8138_), .A1(new_n8136_), .B0(pi0228), .Y(new_n8139_));
  OR2X1    g05703(.A(new_n7786_), .B(pi0044), .Y(new_n8140_));
  AOI21X1  g05704(.A0(new_n7790_), .A1(pi0044), .B0(pi0228), .Y(new_n8141_));
  AOI21X1  g05705(.A0(new_n8141_), .A1(new_n8140_), .B0(pi0039), .Y(new_n8142_));
  AND3X1   g05706(.A(new_n5168_), .B(new_n2479_), .C(new_n2477_), .Y(new_n8143_));
  AOI21X1  g05707(.A0(new_n8143_), .A1(pi0287), .B0(pi0072), .Y(new_n8144_));
  AND3X1   g05708(.A(new_n8144_), .B(new_n5920_), .C(pi0039), .Y(new_n8145_));
  OR2X1    g05709(.A(new_n8145_), .B(new_n3252_), .Y(new_n8146_));
  AOI21X1  g05710(.A0(new_n8142_), .A1(new_n8139_), .B0(new_n8146_), .Y(new_n8147_));
  NAND4X1  g05711(.A(new_n7696_), .B(new_n5168_), .C(new_n2479_), .D(new_n2477_), .Y(new_n8148_));
  AOI21X1  g05712(.A0(new_n8148_), .A1(pi0044), .B0(new_n8124_), .Y(new_n8149_));
  OAI21X1  g05713(.A0(new_n8149_), .A1(new_n8122_), .B0(new_n8119_), .Y(new_n8150_));
  OR2X1    g05714(.A(new_n8128_), .B(new_n5075_), .Y(new_n8151_));
  AOI21X1  g05715(.A0(new_n8150_), .A1(new_n8118_), .B0(new_n8151_), .Y(new_n8152_));
  OAI21X1  g05716(.A0(new_n8131_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n8153_));
  OR2X1    g05717(.A(new_n8153_), .B(new_n8152_), .Y(new_n8154_));
  AND2X1   g05718(.A(new_n3251_), .B(pi0228), .Y(new_n8155_));
  INVX1    g05719(.A(new_n8155_), .Y(new_n8156_));
  NOR4X1   g05720(.A(new_n8156_), .B(new_n2985_), .C(new_n2536_), .D(pi0044), .Y(new_n8157_));
  AOI21X1  g05721(.A0(new_n8155_), .A1(new_n8143_), .B0(new_n8117_), .Y(new_n8158_));
  OR3X1    g05722(.A(new_n8158_), .B(new_n8157_), .C(pi0039), .Y(new_n8159_));
  NOR2X1   g05723(.A(new_n8130_), .B(new_n3131_), .Y(new_n8160_));
  AOI21X1  g05724(.A0(new_n8160_), .A1(new_n8159_), .B0(pi0075), .Y(new_n8161_));
  OAI21X1  g05725(.A0(new_n8154_), .A1(new_n8147_), .B0(new_n8161_), .Y(new_n8162_));
  AOI21X1  g05726(.A0(new_n8162_), .A1(new_n8133_), .B0(new_n6295_), .Y(new_n8163_));
  OAI21X1  g05727(.A0(new_n8131_), .A1(new_n5880_), .B0(new_n6489_), .Y(new_n8164_));
  AND3X1   g05728(.A(new_n5023_), .B(new_n2450_), .C(pi0232), .Y(new_n8165_));
  AOI21X1  g05729(.A0(new_n8165_), .A1(new_n2530_), .B0(new_n2939_), .Y(new_n8166_));
  OAI22X1  g05730(.A0(new_n8116_), .A1(pi0039), .B0(new_n5103_), .B1(pi0057), .Y(new_n8167_));
  OAI22X1  g05731(.A0(new_n8167_), .A1(new_n8166_), .B0(new_n8164_), .B1(new_n8163_), .Y(po0202));
  AND2X1   g05732(.A(pi0039), .B(new_n2979_), .Y(new_n8169_));
  NAND3X1  g05733(.A(new_n8169_), .B(new_n6489_), .C(new_n3103_), .Y(new_n8170_));
  NOR4X1   g05734(.A(new_n8170_), .B(new_n2986_), .C(new_n5026_), .D(pi0287), .Y(po0203));
  INVX1    g05735(.A(new_n6754_), .Y(new_n8172_));
  OR3X1    g05736(.A(pi0111), .B(pi0104), .C(pi0102), .Y(new_n8173_));
  OR4X1    g05737(.A(pi0076), .B(pi0073), .C(pi0068), .D(pi0049), .Y(new_n8174_));
  OR4X1    g05738(.A(new_n8174_), .B(new_n8173_), .C(new_n2469_), .D(pi0071), .Y(new_n8175_));
  NAND4X1  g05739(.A(new_n7614_), .B(new_n2594_), .C(new_n2629_), .D(pi0061), .Y(new_n8176_));
  OR4X1    g05740(.A(new_n8176_), .B(new_n6751_), .C(new_n6749_), .D(new_n5892_), .Y(new_n8177_));
  OR4X1    g05741(.A(new_n8177_), .B(new_n8175_), .C(new_n7659_), .D(new_n8172_), .Y(new_n8178_));
  OR4X1    g05742(.A(new_n2564_), .B(new_n2476_), .C(new_n2473_), .D(new_n2676_), .Y(new_n8179_));
  OAI22X1  g05743(.A0(new_n8179_), .A1(new_n5777_), .B0(new_n8178_), .B1(pi0841), .Y(new_n8180_));
  AND2X1   g05744(.A(new_n8180_), .B(new_n7609_), .Y(po0204));
  NOR2X1   g05745(.A(new_n5931_), .B(pi0058), .Y(new_n8182_));
  OAI21X1  g05746(.A0(new_n2664_), .A1(new_n2663_), .B0(new_n5891_), .Y(new_n8183_));
  NAND3X1  g05747(.A(new_n2601_), .B(pi0104), .C(new_n2603_), .Y(new_n8184_));
  OR4X1    g05748(.A(new_n8184_), .B(new_n7613_), .C(new_n2608_), .D(pi0082), .Y(new_n8185_));
  OR4X1    g05749(.A(pi0107), .B(pi0103), .C(pi0067), .D(pi0063), .Y(new_n8186_));
  OR4X1    g05750(.A(new_n8186_), .B(new_n6836_), .C(new_n6750_), .D(pi0098), .Y(new_n8187_));
  AOI21X1  g05751(.A0(new_n8185_), .A1(new_n2640_), .B0(new_n8187_), .Y(new_n8188_));
  OAI21X1  g05752(.A0(new_n2643_), .A1(new_n2640_), .B0(new_n8188_), .Y(new_n8189_));
  AND2X1   g05753(.A(new_n8189_), .B(new_n2663_), .Y(new_n8190_));
  NOR4X1   g05754(.A(new_n8190_), .B(new_n8183_), .C(new_n2514_), .D(new_n4999_), .Y(new_n8191_));
  OAI21X1  g05755(.A0(new_n8191_), .A1(new_n8182_), .B0(new_n7606_), .Y(new_n8192_));
  AND2X1   g05756(.A(new_n8192_), .B(new_n5970_), .Y(new_n8193_));
  INVX1    g05757(.A(new_n5922_), .Y(new_n8194_));
  OR2X1    g05758(.A(new_n8192_), .B(new_n5225_), .Y(new_n8195_));
  NOR4X1   g05759(.A(new_n7620_), .B(new_n7619_), .C(new_n2526_), .D(new_n2504_), .Y(new_n8196_));
  OR3X1    g05760(.A(new_n8187_), .B(new_n8185_), .C(pi0036), .Y(new_n8197_));
  AOI21X1  g05761(.A0(new_n8197_), .A1(new_n2663_), .B0(new_n8183_), .Y(new_n8198_));
  INVX1    g05762(.A(pi0824), .Y(new_n8199_));
  AND2X1   g05763(.A(new_n5225_), .B(new_n8199_), .Y(new_n8200_));
  NAND3X1  g05764(.A(new_n8200_), .B(new_n8198_), .C(new_n8196_), .Y(new_n8201_));
  AND2X1   g05765(.A(new_n8201_), .B(pi0829), .Y(new_n8202_));
  AND3X1   g05766(.A(new_n8202_), .B(new_n8195_), .C(new_n8194_), .Y(new_n8203_));
  OR2X1    g05767(.A(new_n8203_), .B(new_n8193_), .Y(new_n8204_));
  OR2X1    g05768(.A(new_n8192_), .B(new_n5927_), .Y(new_n8205_));
  AOI22X1  g05769(.A0(new_n8205_), .A1(new_n5237_), .B0(new_n8202_), .B1(new_n8195_), .Y(new_n8206_));
  INVX1    g05770(.A(new_n7608_), .Y(new_n8207_));
  AND2X1   g05771(.A(new_n7606_), .B(new_n5927_), .Y(new_n8208_));
  AOI22X1  g05772(.A0(new_n8208_), .A1(new_n7605_), .B0(new_n5968_), .B1(new_n5238_), .Y(new_n8209_));
  AOI21X1  g05773(.A0(new_n8209_), .A1(new_n8205_), .B0(new_n8207_), .Y(new_n8210_));
  OAI21X1  g05774(.A0(new_n8206_), .A1(pi1093), .B0(new_n8210_), .Y(new_n8211_));
  AOI21X1  g05775(.A0(new_n8204_), .A1(pi1091), .B0(new_n8211_), .Y(po0205));
  NOR3X1   g05776(.A(new_n2707_), .B(new_n2705_), .C(pi0072), .Y(new_n8213_));
  NAND4X1  g05777(.A(new_n8213_), .B(new_n7662_), .C(new_n7608_), .D(new_n2534_), .Y(new_n8214_));
  NOR2X1   g05778(.A(new_n8214_), .B(new_n7621_), .Y(po0206));
  OR2X1    g05779(.A(new_n2469_), .B(new_n2457_), .Y(new_n8216_));
  OR3X1    g05780(.A(new_n7658_), .B(new_n2637_), .C(pi0103), .Y(new_n8217_));
  OR4X1    g05781(.A(new_n8217_), .B(new_n6750_), .C(pi0073), .D(pi0068), .Y(new_n8218_));
  OR3X1    g05782(.A(new_n8173_), .B(new_n2617_), .C(pi0045), .Y(new_n8219_));
  OR3X1    g05783(.A(new_n8219_), .B(new_n8218_), .C(new_n8216_), .Y(new_n8220_));
  NOR3X1   g05784(.A(new_n8220_), .B(new_n2608_), .C(pi0082), .Y(new_n8221_));
  NAND4X1  g05785(.A(new_n8221_), .B(new_n6754_), .C(new_n2534_), .D(new_n2508_), .Y(new_n8222_));
  NAND3X1  g05786(.A(new_n8213_), .B(new_n5168_), .C(new_n2483_), .Y(new_n8223_));
  OAI21X1  g05787(.A0(new_n8223_), .A1(new_n8222_), .B0(new_n4982_), .Y(new_n8224_));
  NAND3X1  g05788(.A(new_n8224_), .B(new_n6489_), .C(new_n5839_), .Y(new_n8225_));
  AOI21X1  g05789(.A0(new_n7553_), .A1(pi0074), .B0(new_n8225_), .Y(po0207));
  AND2X1   g05790(.A(new_n6737_), .B(pi0024), .Y(new_n8227_));
  AOI21X1  g05791(.A0(new_n2570_), .A1(new_n2497_), .B0(new_n8227_), .Y(new_n8228_));
  NAND3X1  g05792(.A(new_n6736_), .B(new_n2572_), .C(pi0024), .Y(new_n8229_));
  MX2X1    g05793(.A(po0840), .B(new_n6728_), .S0(new_n3035_), .Y(new_n8230_));
  NAND3X1  g05794(.A(new_n8230_), .B(new_n8229_), .C(new_n7606_), .Y(new_n8231_));
  AND3X1   g05795(.A(new_n2984_), .B(new_n2517_), .C(new_n2513_), .Y(new_n8232_));
  INVX1    g05796(.A(new_n8232_), .Y(new_n8233_));
  OR4X1    g05797(.A(new_n8233_), .B(new_n8230_), .C(pi0090), .D(new_n5777_), .Y(new_n8234_));
  OR4X1    g05798(.A(new_n8234_), .B(new_n6738_), .C(new_n6736_), .D(pi0093), .Y(new_n8235_));
  OAI21X1  g05799(.A0(new_n8231_), .A1(new_n8228_), .B0(new_n8235_), .Y(new_n8236_));
  AND3X1   g05800(.A(new_n5263_), .B(new_n5072_), .C(pi0100), .Y(new_n8237_));
  AOI21X1  g05801(.A0(new_n8236_), .A1(new_n3007_), .B0(new_n8237_), .Y(new_n8238_));
  OR4X1    g05802(.A(pi0087), .B(pi0075), .C(pi0039), .D(pi0038), .Y(new_n8239_));
  OR3X1    g05803(.A(new_n6779_), .B(new_n5082_), .C(new_n5071_), .Y(new_n8240_));
  OAI22X1  g05804(.A0(new_n8240_), .A1(new_n6774_), .B0(new_n8239_), .B1(new_n8238_), .Y(new_n8241_));
  AND2X1   g05805(.A(new_n8241_), .B(new_n6722_), .Y(po0208));
  INVX1    g05806(.A(new_n7606_), .Y(new_n8243_));
  NOR4X1   g05807(.A(new_n8207_), .B(new_n8243_), .C(new_n2514_), .D(new_n4999_), .Y(new_n8244_));
  OR4X1    g05808(.A(new_n6836_), .B(new_n2469_), .C(new_n2459_), .D(new_n2457_), .Y(new_n8245_));
  OR4X1    g05809(.A(new_n8245_), .B(new_n2637_), .C(new_n2460_), .D(pi0069), .Y(new_n8246_));
  NOR4X1   g05810(.A(new_n8246_), .B(new_n2633_), .C(new_n2602_), .D(new_n2629_), .Y(new_n8247_));
  AND2X1   g05811(.A(new_n8247_), .B(new_n8244_), .Y(po0209));
  OR3X1    g05812(.A(new_n7996_), .B(pi0219), .C(pi0211), .Y(new_n8249_));
  AND3X1   g05813(.A(new_n2530_), .B(pi0052), .C(new_n2939_), .Y(new_n8250_));
  AND2X1   g05814(.A(new_n2530_), .B(pi0052), .Y(new_n8251_));
  NOR4X1   g05815(.A(pi0115), .B(pi0114), .C(pi0043), .D(pi0042), .Y(new_n8252_));
  NAND2X1  g05816(.A(new_n8252_), .B(pi0228), .Y(new_n8253_));
  INVX1    g05817(.A(pi0052), .Y(new_n8254_));
  NOR2X1   g05818(.A(new_n7896_), .B(pi0072), .Y(new_n8255_));
  MX2X1    g05819(.A(new_n8255_), .B(new_n8035_), .S0(new_n8254_), .Y(new_n8256_));
  MX2X1    g05820(.A(new_n8256_), .B(new_n8251_), .S0(new_n8253_), .Y(new_n8257_));
  MX2X1    g05821(.A(new_n8257_), .B(new_n8250_), .S0(pi0038), .Y(new_n8258_));
  NOR2X1   g05822(.A(new_n8250_), .B(new_n3007_), .Y(new_n8259_));
  OR3X1    g05823(.A(pi0100), .B(new_n2939_), .C(pi0038), .Y(new_n8260_));
  NAND2X1  g05824(.A(new_n8260_), .B(pi0087), .Y(new_n8261_));
  NOR2X1   g05825(.A(new_n8261_), .B(new_n8259_), .Y(new_n8262_));
  OAI21X1  g05826(.A0(new_n8258_), .A1(pi0100), .B0(new_n8262_), .Y(new_n8263_));
  OR3X1    g05827(.A(pi0114), .B(pi0043), .C(pi0042), .Y(new_n8264_));
  AOI21X1  g05828(.A0(new_n7840_), .A1(new_n8254_), .B0(new_n7888_), .Y(new_n8265_));
  OAI21X1  g05829(.A0(new_n7836_), .A1(new_n8254_), .B0(new_n8265_), .Y(new_n8266_));
  INVX1    g05830(.A(new_n7844_), .Y(new_n8267_));
  AOI21X1  g05831(.A0(new_n7850_), .A1(new_n8254_), .B0(new_n8267_), .Y(new_n8268_));
  OAI21X1  g05832(.A0(new_n8000_), .A1(new_n8254_), .B0(new_n8268_), .Y(new_n8269_));
  AOI21X1  g05833(.A0(new_n8269_), .A1(new_n8266_), .B0(new_n8264_), .Y(new_n8270_));
  AOI21X1  g05834(.A0(new_n2530_), .A1(pi0052), .B0(new_n8252_), .Y(new_n8271_));
  NOR3X1   g05835(.A(new_n8271_), .B(new_n8270_), .C(new_n2793_), .Y(new_n8272_));
  OAI21X1  g05836(.A0(new_n7865_), .A1(pi0052), .B0(new_n8252_), .Y(new_n8273_));
  AOI21X1  g05837(.A0(new_n7859_), .A1(pi0052), .B0(new_n8273_), .Y(new_n8274_));
  OR2X1    g05838(.A(new_n8271_), .B(pi0228), .Y(new_n8275_));
  OAI21X1  g05839(.A0(new_n8275_), .A1(new_n8274_), .B0(new_n2939_), .Y(new_n8276_));
  OR3X1    g05840(.A(new_n8276_), .B(new_n8272_), .C(pi0100), .Y(new_n8277_));
  NOR4X1   g05841(.A(new_n5920_), .B(new_n2704_), .C(new_n2793_), .D(pi0115), .Y(new_n8278_));
  INVX1    g05842(.A(new_n8278_), .Y(new_n8279_));
  OR3X1    g05843(.A(new_n8279_), .B(new_n8264_), .C(new_n7697_), .Y(new_n8280_));
  OAI21X1  g05844(.A0(new_n8280_), .A1(new_n7897_), .B0(new_n8251_), .Y(new_n8281_));
  AOI21X1  g05845(.A0(new_n8281_), .A1(pi0100), .B0(pi0039), .Y(new_n8282_));
  AOI21X1  g05846(.A0(new_n8282_), .A1(new_n8277_), .B0(pi0038), .Y(new_n8283_));
  OAI21X1  g05847(.A0(new_n8250_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n8284_));
  OAI21X1  g05848(.A0(new_n8284_), .A1(new_n8283_), .B0(new_n8263_), .Y(new_n8285_));
  OR4X1    g05849(.A(new_n8279_), .B(new_n8264_), .C(new_n7925_), .D(new_n5778_), .Y(new_n8286_));
  NAND2X1  g05850(.A(new_n8286_), .B(new_n8250_), .Y(new_n8287_));
  OAI21X1  g05851(.A0(new_n8287_), .A1(new_n3073_), .B0(new_n5880_), .Y(new_n8288_));
  AOI21X1  g05852(.A0(new_n8285_), .A1(new_n3073_), .B0(new_n8288_), .Y(new_n8289_));
  OAI21X1  g05853(.A0(new_n8250_), .A1(new_n5880_), .B0(new_n7826_), .Y(new_n8290_));
  NOR2X1   g05854(.A(new_n8276_), .B(new_n8272_), .Y(new_n8291_));
  OAI21X1  g05855(.A0(new_n8291_), .A1(new_n8060_), .B0(new_n3251_), .Y(new_n8292_));
  AND2X1   g05856(.A(new_n8281_), .B(new_n2939_), .Y(new_n8293_));
  OAI21X1  g05857(.A0(new_n8293_), .A1(new_n8066_), .B0(new_n5074_), .Y(new_n8294_));
  MX2X1    g05858(.A(new_n8251_), .B(new_n8065_), .S0(pi0039), .Y(new_n8295_));
  OR2X1    g05859(.A(new_n8295_), .B(new_n2979_), .Y(new_n8296_));
  AND3X1   g05860(.A(new_n8296_), .B(new_n8294_), .C(new_n3131_), .Y(new_n8297_));
  OR2X1    g05861(.A(new_n8257_), .B(pi0039), .Y(new_n8298_));
  NOR2X1   g05862(.A(new_n8066_), .B(new_n3252_), .Y(new_n8299_));
  AOI22X1  g05863(.A0(new_n8299_), .A1(new_n8298_), .B0(new_n8295_), .B1(new_n3252_), .Y(new_n8300_));
  OAI21X1  g05864(.A0(new_n8300_), .A1(new_n3131_), .B0(new_n3073_), .Y(new_n8301_));
  AOI21X1  g05865(.A0(new_n8297_), .A1(new_n8292_), .B0(new_n8301_), .Y(new_n8302_));
  INVX1    g05866(.A(new_n8251_), .Y(new_n8303_));
  NOR3X1   g05867(.A(new_n8279_), .B(new_n8264_), .C(new_n7925_), .Y(new_n8304_));
  OAI21X1  g05868(.A0(new_n8304_), .A1(new_n8303_), .B0(new_n2939_), .Y(new_n8305_));
  NOR2X1   g05869(.A(new_n8066_), .B(new_n5778_), .Y(new_n8306_));
  AND2X1   g05870(.A(new_n8295_), .B(new_n5778_), .Y(new_n8307_));
  OR2X1    g05871(.A(new_n8307_), .B(new_n3073_), .Y(new_n8308_));
  AOI21X1  g05872(.A0(new_n8306_), .A1(new_n8305_), .B0(new_n8308_), .Y(new_n8309_));
  OR3X1    g05873(.A(new_n8309_), .B(new_n7826_), .C(new_n6295_), .Y(new_n8310_));
  OAI22X1  g05874(.A0(new_n8310_), .A1(new_n8302_), .B0(new_n8290_), .B1(new_n8289_), .Y(new_n8311_));
  NAND2X1  g05875(.A(new_n8311_), .B(new_n8249_), .Y(new_n8312_));
  OAI21X1  g05876(.A0(new_n7882_), .A1(new_n7880_), .B0(pi0039), .Y(new_n8313_));
  OAI21X1  g05877(.A0(new_n8276_), .A1(new_n8272_), .B0(new_n8313_), .Y(new_n8314_));
  AOI21X1  g05878(.A0(new_n8303_), .A1(new_n2939_), .B0(new_n7905_), .Y(new_n8315_));
  AOI21X1  g05879(.A0(new_n8281_), .A1(new_n2939_), .B0(new_n7905_), .Y(new_n8316_));
  OAI22X1  g05880(.A0(new_n8316_), .A1(new_n5075_), .B0(new_n8315_), .B1(new_n2979_), .Y(new_n8317_));
  AOI21X1  g05881(.A0(new_n8314_), .A1(new_n3251_), .B0(new_n8317_), .Y(new_n8318_));
  OR2X1    g05882(.A(new_n8318_), .B(pi0087), .Y(new_n8319_));
  AOI21X1  g05883(.A0(new_n8315_), .A1(new_n3252_), .B0(new_n3131_), .Y(new_n8320_));
  NOR2X1   g05884(.A(new_n7905_), .B(new_n3252_), .Y(new_n8321_));
  OAI21X1  g05885(.A0(new_n8257_), .A1(pi0039), .B0(new_n8321_), .Y(new_n8322_));
  AOI21X1  g05886(.A0(new_n8322_), .A1(new_n8320_), .B0(new_n7827_), .Y(new_n8323_));
  NOR2X1   g05887(.A(new_n8291_), .B(new_n8097_), .Y(new_n8324_));
  NOR2X1   g05888(.A(new_n8324_), .B(new_n3252_), .Y(new_n8325_));
  AOI21X1  g05889(.A0(new_n8281_), .A1(new_n2939_), .B0(new_n8100_), .Y(new_n8326_));
  OAI22X1  g05890(.A0(new_n8326_), .A1(new_n5075_), .B0(new_n8315_), .B1(new_n8296_), .Y(new_n8327_));
  OAI21X1  g05891(.A0(new_n8327_), .A1(new_n8325_), .B0(new_n3131_), .Y(new_n8328_));
  INVX1    g05892(.A(new_n8100_), .Y(new_n8329_));
  NAND3X1  g05893(.A(new_n8298_), .B(new_n8329_), .C(new_n3251_), .Y(new_n8330_));
  NAND2X1  g05894(.A(new_n8295_), .B(new_n3252_), .Y(new_n8331_));
  AND2X1   g05895(.A(new_n8320_), .B(new_n8331_), .Y(new_n8332_));
  AOI21X1  g05896(.A0(new_n8332_), .A1(new_n8330_), .B0(new_n7826_), .Y(new_n8333_));
  AOI22X1  g05897(.A0(new_n8333_), .A1(new_n8328_), .B0(new_n8323_), .B1(new_n8319_), .Y(new_n8334_));
  AOI21X1  g05898(.A0(new_n7905_), .A1(new_n7826_), .B0(new_n3073_), .Y(new_n8335_));
  OAI21X1  g05899(.A0(new_n8329_), .A1(new_n7826_), .B0(new_n8335_), .Y(new_n8336_));
  AOI21X1  g05900(.A0(new_n8287_), .A1(new_n2939_), .B0(new_n8336_), .Y(new_n8337_));
  NOR2X1   g05901(.A(new_n8337_), .B(new_n6295_), .Y(new_n8338_));
  OAI21X1  g05902(.A0(new_n8334_), .A1(pi0075), .B0(new_n8338_), .Y(new_n8339_));
  NOR2X1   g05903(.A(new_n8315_), .B(new_n5880_), .Y(new_n8340_));
  NOR2X1   g05904(.A(new_n8340_), .B(new_n8249_), .Y(new_n8341_));
  AND3X1   g05905(.A(new_n8295_), .B(new_n7827_), .C(new_n6295_), .Y(new_n8342_));
  OR2X1    g05906(.A(new_n8342_), .B(po1038), .Y(new_n8343_));
  AOI21X1  g05907(.A0(new_n8341_), .A1(new_n8339_), .B0(new_n8343_), .Y(new_n8344_));
  NOR4X1   g05908(.A(new_n7996_), .B(pi0219), .C(pi0211), .D(new_n2939_), .Y(new_n8345_));
  OR2X1    g05909(.A(new_n8250_), .B(new_n6489_), .Y(new_n8346_));
  AOI21X1  g05910(.A0(new_n8345_), .A1(new_n7878_), .B0(new_n8346_), .Y(new_n8347_));
  AOI21X1  g05911(.A0(new_n8344_), .A1(new_n8312_), .B0(new_n8347_), .Y(po0210));
  AND2X1   g05912(.A(new_n7606_), .B(pi0024), .Y(new_n8349_));
  NOR4X1   g05913(.A(new_n2498_), .B(new_n2491_), .C(new_n2490_), .D(new_n2485_), .Y(new_n8350_));
  AOI21X1  g05914(.A0(new_n8350_), .A1(new_n8349_), .B0(pi0039), .Y(new_n8351_));
  AND3X1   g05915(.A(new_n5025_), .B(new_n5026_), .C(new_n7795_), .Y(new_n8352_));
  OAI21X1  g05916(.A0(new_n8352_), .A1(new_n2939_), .B0(new_n7628_), .Y(new_n8353_));
  NOR3X1   g05917(.A(new_n8353_), .B(new_n8351_), .C(new_n3169_), .Y(po0211));
  INVX1    g05918(.A(new_n3088_), .Y(new_n8355_));
  OAI21X1  g05919(.A0(new_n7611_), .A1(new_n8355_), .B0(pi0054), .Y(new_n8356_));
  NAND4X1  g05920(.A(new_n6737_), .B(new_n2496_), .C(new_n2489_), .D(new_n2485_), .Y(new_n8357_));
  INVX1    g05921(.A(pi0106), .Y(new_n8358_));
  OR2X1    g05922(.A(pi0085), .B(pi0060), .Y(new_n8359_));
  OR4X1    g05923(.A(pi0111), .B(pi0102), .C(pi0089), .D(pi0082), .Y(new_n8360_));
  OR4X1    g05924(.A(new_n8360_), .B(new_n8359_), .C(new_n8174_), .D(new_n8358_), .Y(new_n8361_));
  OR4X1    g05925(.A(new_n8361_), .B(new_n8217_), .C(new_n8216_), .D(new_n6752_), .Y(new_n8362_));
  NAND4X1  g05926(.A(new_n3084_), .B(new_n3070_), .C(new_n2534_), .D(new_n2508_), .Y(new_n8363_));
  OR4X1    g05927(.A(new_n8363_), .B(new_n6773_), .C(new_n2484_), .D(pi0841), .Y(new_n8364_));
  NOR3X1   g05928(.A(new_n8364_), .B(new_n8362_), .C(new_n8357_), .Y(new_n8365_));
  OR2X1    g05929(.A(new_n8365_), .B(pi0054), .Y(new_n8366_));
  AND3X1   g05930(.A(new_n8366_), .B(new_n8356_), .C(new_n6721_), .Y(po0212));
  OR4X1    g05931(.A(new_n7611_), .B(new_n8355_), .C(pi0074), .D(pi0054), .Y(new_n8368_));
  NAND3X1  g05932(.A(new_n6895_), .B(new_n5122_), .C(pi0045), .Y(new_n8369_));
  OR4X1    g05933(.A(new_n8369_), .B(new_n8218_), .C(new_n2464_), .D(pi0104), .Y(new_n8370_));
  NAND4X1  g05934(.A(new_n6754_), .B(new_n5168_), .C(new_n5010_), .D(new_n2483_), .Y(new_n8371_));
  NOR4X1   g05935(.A(new_n8371_), .B(new_n8370_), .C(new_n3105_), .D(new_n2458_), .Y(new_n8372_));
  OAI21X1  g05936(.A0(new_n8372_), .A1(pi0055), .B0(new_n6720_), .Y(new_n8373_));
  AOI21X1  g05937(.A0(new_n8368_), .A1(pi0055), .B0(new_n8373_), .Y(po0213));
  NOR3X1   g05938(.A(new_n7553_), .B(new_n4975_), .C(new_n3105_), .Y(new_n8375_));
  AND2X1   g05939(.A(new_n3222_), .B(pi0056), .Y(new_n8376_));
  AOI21X1  g05940(.A0(new_n8375_), .A1(pi0055), .B0(new_n8376_), .Y(new_n8377_));
  AND3X1   g05941(.A(new_n3113_), .B(new_n3111_), .C(new_n7228_), .Y(new_n8378_));
  AOI21X1  g05942(.A0(new_n8378_), .A1(new_n5011_), .B0(new_n3118_), .Y(new_n8379_));
  NOR3X1   g05943(.A(new_n8379_), .B(new_n8377_), .C(new_n3374_), .Y(po0214));
  INVX1    g05944(.A(new_n5306_), .Y(new_n8381_));
  OAI21X1  g05945(.A0(new_n8368_), .A1(new_n8381_), .B0(pi0057), .Y(new_n8382_));
  NOR3X1   g05946(.A(new_n5173_), .B(new_n2747_), .C(new_n5172_), .Y(new_n8383_));
  NAND2X1  g05947(.A(new_n8378_), .B(new_n8383_), .Y(new_n8384_));
  INVX1    g05948(.A(pi0924), .Y(new_n8385_));
  AND2X1   g05949(.A(pi0062), .B(new_n3118_), .Y(new_n8386_));
  AOI21X1  g05950(.A0(new_n8386_), .A1(new_n8385_), .B0(new_n8376_), .Y(new_n8387_));
  OAI21X1  g05951(.A0(new_n8387_), .A1(new_n8384_), .B0(new_n2436_), .Y(new_n8388_));
  AND3X1   g05952(.A(new_n8388_), .B(new_n8382_), .C(new_n3127_), .Y(po0215));
  INVX1    g05953(.A(new_n2477_), .Y(new_n8390_));
  NAND3X1  g05954(.A(new_n8232_), .B(new_n7608_), .C(new_n2516_), .Y(new_n8391_));
  NOR4X1   g05955(.A(new_n8391_), .B(new_n8390_), .C(pi0841), .D(new_n2682_), .Y(po0216));
  OAI21X1  g05956(.A0(new_n8368_), .A1(new_n8381_), .B0(pi0059), .Y(new_n8393_));
  NAND4X1  g05957(.A(new_n8386_), .B(new_n8378_), .C(new_n8383_), .D(pi0924), .Y(new_n8394_));
  AOI21X1  g05958(.A0(new_n8394_), .A1(new_n3127_), .B0(pi0057), .Y(new_n8395_));
  AND2X1   g05959(.A(new_n8395_), .B(new_n8393_), .Y(po0217));
  OR4X1    g05960(.A(new_n5027_), .B(new_n5025_), .C(pi0979), .D(new_n2939_), .Y(new_n8397_));
  OR4X1    g05961(.A(new_n8397_), .B(new_n2985_), .C(new_n2536_), .D(pi0287), .Y(new_n8398_));
  OR4X1    g05962(.A(new_n8357_), .B(new_n8243_), .C(pi0039), .D(new_n5777_), .Y(new_n8399_));
  OR2X1    g05963(.A(new_n8399_), .B(new_n2487_), .Y(new_n8400_));
  AOI21X1  g05964(.A0(new_n8400_), .A1(new_n8398_), .B0(new_n7629_), .Y(po0218));
  OR2X1    g05965(.A(new_n8357_), .B(pi0024), .Y(new_n8402_));
  OAI22X1  g05966(.A0(new_n8402_), .A1(new_n2487_), .B0(new_n8178_), .B1(new_n2705_), .Y(new_n8403_));
  AND2X1   g05967(.A(new_n8403_), .B(new_n7609_), .Y(po0219));
  OR2X1    g05968(.A(new_n7597_), .B(new_n2436_), .Y(new_n8405_));
  NAND3X1  g05969(.A(new_n8386_), .B(new_n8378_), .C(new_n5011_), .Y(new_n8406_));
  AOI21X1  g05970(.A0(new_n8406_), .A1(new_n2436_), .B0(pi0059), .Y(new_n8407_));
  AND2X1   g05971(.A(new_n8407_), .B(new_n8405_), .Y(po0220));
  INVX1    g05972(.A(pi0999), .Y(new_n8409_));
  OR4X1    g05973(.A(new_n6837_), .B(new_n8172_), .C(new_n2657_), .D(new_n2468_), .Y(new_n8410_));
  OAI22X1  g05974(.A0(new_n8410_), .A1(new_n8409_), .B0(new_n8179_), .B1(pi0024), .Y(new_n8411_));
  AND2X1   g05975(.A(new_n8411_), .B(new_n7609_), .Y(po0221));
  OR4X1    g05976(.A(new_n2468_), .B(new_n2459_), .C(new_n2587_), .D(pi0063), .Y(new_n8413_));
  AND2X1   g05977(.A(new_n8413_), .B(new_n2584_), .Y(new_n8414_));
  OR4X1    g05978(.A(new_n8414_), .B(new_n2586_), .C(new_n2458_), .D(pi0081), .Y(new_n8415_));
  NOR4X1   g05979(.A(new_n6837_), .B(new_n2468_), .C(new_n2587_), .D(pi0063), .Y(new_n8416_));
  OAI21X1  g05980(.A0(new_n8416_), .A1(pi0841), .B0(new_n8244_), .Y(new_n8417_));
  AOI21X1  g05981(.A0(new_n8415_), .A1(pi0841), .B0(new_n8417_), .Y(po0222));
  NOR3X1   g05982(.A(new_n7646_), .B(new_n7645_), .C(new_n2933_), .Y(new_n8419_));
  OR3X1    g05983(.A(pi1082), .B(new_n7648_), .C(new_n2939_), .Y(new_n8420_));
  NOR4X1   g05984(.A(new_n8420_), .B(new_n8419_), .C(new_n7642_), .D(new_n7629_), .Y(po0223));
  INVX1    g05985(.A(pi0219), .Y(new_n8422_));
  NOR2X1   g05986(.A(pi0299), .B(pi0199), .Y(new_n8423_));
  OR3X1    g05987(.A(new_n8371_), .B(new_n2457_), .C(new_n5117_), .Y(new_n8424_));
  OR4X1    g05988(.A(new_n8424_), .B(new_n2470_), .C(pi0102), .D(new_n2579_), .Y(new_n8425_));
  NOR3X1   g05989(.A(new_n8425_), .B(new_n8423_), .C(new_n3105_), .Y(new_n8426_));
  OR2X1    g05990(.A(new_n8426_), .B(new_n8422_), .Y(new_n8427_));
  NAND3X1  g05991(.A(new_n3102_), .B(new_n3084_), .C(new_n3251_), .Y(new_n8428_));
  OR4X1    g05992(.A(new_n8428_), .B(new_n7141_), .C(pi0299), .D(new_n7871_), .Y(new_n8429_));
  OAI21X1  g05993(.A0(new_n8429_), .A1(new_n8425_), .B0(new_n8422_), .Y(new_n8430_));
  AND3X1   g05994(.A(new_n8430_), .B(new_n8427_), .C(new_n6489_), .Y(po0224));
  OR4X1    g05995(.A(new_n8245_), .B(new_n8207_), .C(pi0103), .D(new_n2594_), .Y(new_n8432_));
  NOR4X1   g05996(.A(new_n8432_), .B(new_n8424_), .C(new_n5130_), .D(new_n2461_), .Y(po0225));
  NOR4X1   g05997(.A(new_n5239_), .B(new_n5228_), .C(new_n5224_), .D(new_n5062_), .Y(new_n8434_));
  NOR4X1   g05998(.A(new_n2933_), .B(pi0221), .C(new_n2438_), .D(pi0215), .Y(new_n8435_));
  NOR4X1   g05999(.A(new_n5239_), .B(new_n5228_), .C(new_n5224_), .D(new_n5049_), .Y(new_n8436_));
  AND3X1   g06000(.A(new_n4769_), .B(pi0224), .C(new_n2941_), .Y(new_n8437_));
  AOI22X1  g06001(.A0(new_n8437_), .A1(new_n8436_), .B0(new_n8435_), .B1(new_n8434_), .Y(new_n8438_));
  NOR2X1   g06002(.A(new_n8438_), .B(new_n8170_), .Y(po0226));
  INVX1    g06003(.A(new_n8244_), .Y(new_n8440_));
  NOR3X1   g06004(.A(new_n2637_), .B(pi0103), .C(new_n2591_), .Y(new_n8441_));
  NAND3X1  g06005(.A(new_n8441_), .B(new_n2643_), .C(new_n2594_), .Y(new_n8442_));
  AND2X1   g06006(.A(new_n8442_), .B(new_n2590_), .Y(new_n8443_));
  OR2X1    g06007(.A(pi0314), .B(pi0081), .Y(new_n8444_));
  OR4X1    g06008(.A(new_n8444_), .B(new_n8443_), .C(new_n5136_), .D(new_n2458_), .Y(new_n8445_));
  NAND3X1  g06009(.A(new_n5891_), .B(pi0314), .C(pi0071), .Y(new_n8446_));
  OR3X1    g06010(.A(new_n8446_), .B(new_n7601_), .C(new_n2468_), .Y(new_n8447_));
  AOI21X1  g06011(.A0(new_n8447_), .A1(new_n8445_), .B0(new_n8440_), .Y(po0227));
  NAND2X1  g06012(.A(new_n2984_), .B(new_n2939_), .Y(new_n8449_));
  OR4X1    g06013(.A(new_n2689_), .B(pi0096), .C(new_n2535_), .D(pi0051), .Y(new_n8450_));
  OR3X1    g06014(.A(new_n8450_), .B(new_n8449_), .C(new_n5777_), .Y(new_n8451_));
  AND2X1   g06015(.A(pi0589), .B(pi0198), .Y(new_n8452_));
  NOR2X1   g06016(.A(new_n5049_), .B(new_n3261_), .Y(new_n8453_));
  AND2X1   g06017(.A(pi0589), .B(pi0210), .Y(new_n8454_));
  OR3X1    g06018(.A(new_n2933_), .B(pi0221), .C(pi0215), .Y(new_n8455_));
  NOR3X1   g06019(.A(new_n8455_), .B(new_n5062_), .C(pi0216), .Y(new_n8456_));
  AOI22X1  g06020(.A0(new_n8456_), .A1(new_n8454_), .B0(new_n8453_), .B1(new_n8452_), .Y(new_n8457_));
  NOR4X1   g06021(.A(new_n8457_), .B(new_n5234_), .C(new_n5223_), .D(pi0593), .Y(new_n8458_));
  OAI21X1  g06022(.A0(new_n8458_), .A1(pi0287), .B0(pi0039), .Y(new_n8459_));
  OR2X1    g06023(.A(new_n8459_), .B(new_n2986_), .Y(new_n8460_));
  AOI21X1  g06024(.A0(new_n8460_), .A1(new_n8451_), .B0(new_n7629_), .Y(po0228));
  AND3X1   g06025(.A(new_n6754_), .B(new_n5141_), .C(new_n6734_), .Y(new_n8462_));
  INVX1    g06026(.A(new_n8462_), .Y(new_n8463_));
  OR4X1    g06027(.A(new_n2465_), .B(new_n2462_), .C(pi0084), .D(pi0068), .Y(new_n8464_));
  OR4X1    g06028(.A(new_n8464_), .B(new_n2622_), .C(new_n2606_), .D(new_n5124_), .Y(new_n8465_));
  NOR4X1   g06029(.A(new_n8465_), .B(new_n8186_), .C(new_n6750_), .D(pi0064), .Y(new_n8466_));
  AND3X1   g06030(.A(new_n2933_), .B(pi0200), .C(new_n7871_), .Y(new_n8467_));
  AND3X1   g06031(.A(pi0299), .B(new_n8422_), .C(pi0211), .Y(new_n8468_));
  NOR2X1   g06032(.A(new_n8468_), .B(new_n8467_), .Y(new_n8469_));
  INVX1    g06033(.A(new_n8469_), .Y(new_n8470_));
  AND3X1   g06034(.A(new_n8470_), .B(new_n7606_), .C(pi0314), .Y(new_n8471_));
  OAI21X1  g06035(.A0(new_n8466_), .A1(pi0081), .B0(new_n8471_), .Y(new_n8472_));
  OR4X1    g06036(.A(new_n8470_), .B(new_n8424_), .C(new_n6836_), .D(new_n6750_), .Y(new_n8473_));
  OR3X1    g06037(.A(new_n8473_), .B(new_n8465_), .C(new_n8186_), .Y(new_n8474_));
  OAI21X1  g06038(.A0(new_n8472_), .A1(new_n8463_), .B0(new_n8474_), .Y(new_n8475_));
  AND2X1   g06039(.A(new_n8475_), .B(new_n7608_), .Y(po0229));
  AND3X1   g06040(.A(new_n2531_), .B(pi0072), .C(pi0024), .Y(new_n8477_));
  INVX1    g06041(.A(new_n2664_), .Y(new_n8478_));
  INVX1    g06042(.A(new_n6933_), .Y(new_n8479_));
  OR4X1    g06043(.A(new_n2561_), .B(new_n6914_), .C(new_n2663_), .D(pi0058), .Y(new_n8480_));
  NOR4X1   g06044(.A(new_n8480_), .B(new_n8479_), .C(new_n5233_), .D(new_n8478_), .Y(new_n8481_));
  OAI21X1  g06045(.A0(new_n8481_), .A1(new_n8477_), .B0(new_n5168_), .Y(new_n8482_));
  NAND2X1  g06046(.A(new_n8482_), .B(new_n2939_), .Y(new_n8483_));
  AND3X1   g06047(.A(new_n8434_), .B(new_n5331_), .C(new_n2438_), .Y(new_n8484_));
  INVX1    g06048(.A(new_n8484_), .Y(new_n8485_));
  AOI21X1  g06049(.A0(new_n8436_), .A1(new_n5951_), .B0(new_n2939_), .Y(new_n8486_));
  AOI21X1  g06050(.A0(new_n8486_), .A1(new_n8485_), .B0(new_n7629_), .Y(new_n8487_));
  AND2X1   g06051(.A(new_n8487_), .B(new_n8483_), .Y(po0230));
  AND2X1   g06052(.A(new_n8436_), .B(new_n6848_), .Y(new_n8489_));
  AOI21X1  g06053(.A0(new_n8434_), .A1(new_n6856_), .B0(new_n2933_), .Y(new_n8490_));
  INVX1    g06054(.A(new_n8490_), .Y(new_n8491_));
  OAI21X1  g06055(.A0(new_n8489_), .A1(pi0299), .B0(new_n8491_), .Y(new_n8492_));
  INVX1    g06056(.A(pi1050), .Y(new_n8493_));
  NAND4X1  g06057(.A(new_n7606_), .B(new_n6910_), .C(new_n6754_), .D(new_n6895_), .Y(new_n8494_));
  NOR3X1   g06058(.A(new_n8494_), .B(new_n8493_), .C(pi0314), .Y(new_n8495_));
  OAI21X1  g06059(.A0(new_n8495_), .A1(pi0039), .B0(new_n7628_), .Y(new_n8496_));
  AOI21X1  g06060(.A0(new_n8492_), .A1(pi0039), .B0(new_n8496_), .Y(po0231));
  OR4X1    g06061(.A(new_n7611_), .B(new_n8355_), .C(new_n4982_), .D(pi0054), .Y(new_n8498_));
  OR4X1    g06062(.A(new_n5932_), .B(new_n2561_), .C(new_n2559_), .D(new_n2518_), .Y(new_n8499_));
  AND2X1   g06063(.A(new_n8499_), .B(new_n2513_), .Y(new_n8500_));
  NAND3X1  g06064(.A(new_n5927_), .B(new_n5032_), .C(new_n2513_), .Y(new_n8501_));
  AND3X1   g06065(.A(new_n5880_), .B(new_n3111_), .C(new_n3077_), .Y(new_n8502_));
  OAI21X1  g06066(.A0(new_n5009_), .A1(pi0096), .B0(pi0479), .Y(new_n8503_));
  NAND4X1  g06067(.A(new_n8503_), .B(new_n8502_), .C(new_n8501_), .D(new_n6741_), .Y(new_n8504_));
  OR4X1    g06068(.A(new_n8504_), .B(new_n8500_), .C(new_n5905_), .D(new_n5881_), .Y(new_n8505_));
  AOI21X1  g06069(.A0(new_n8505_), .A1(new_n8498_), .B0(po1038), .Y(po0232));
  OAI22X1  g06070(.A0(new_n8500_), .A1(new_n2760_), .B0(pi1093), .B1(new_n2513_), .Y(new_n8507_));
  NAND3X1  g06071(.A(new_n8507_), .B(new_n5937_), .C(new_n3070_), .Y(new_n8508_));
  OAI21X1  g06072(.A0(new_n7611_), .A1(new_n5778_), .B0(pi0075), .Y(new_n8509_));
  NAND2X1  g06073(.A(new_n8509_), .B(new_n6722_), .Y(new_n8510_));
  AOI21X1  g06074(.A0(new_n8508_), .A1(new_n3073_), .B0(new_n8510_), .Y(po0233));
  AND2X1   g06075(.A(new_n2761_), .B(pi0252), .Y(new_n8512_));
  OR4X1    g06076(.A(new_n8512_), .B(new_n7766_), .C(new_n5881_), .D(new_n7763_), .Y(new_n8513_));
  NOR2X1   g06077(.A(new_n8513_), .B(pi0137), .Y(new_n8514_));
  AND2X1   g06078(.A(new_n2703_), .B(new_n2452_), .Y(new_n8515_));
  OAI21X1  g06079(.A0(new_n6757_), .A1(new_n2472_), .B0(new_n2572_), .Y(new_n8516_));
  NAND2X1  g06080(.A(new_n8516_), .B(new_n7606_), .Y(new_n8517_));
  AOI21X1  g06081(.A0(new_n7766_), .A1(new_n6738_), .B0(new_n8517_), .Y(new_n8518_));
  NOR2X1   g06082(.A(new_n8518_), .B(new_n2761_), .Y(new_n8519_));
  AND3X1   g06083(.A(new_n8196_), .B(new_n6753_), .C(pi0252), .Y(new_n8520_));
  OR2X1    g06084(.A(new_n8520_), .B(new_n2762_), .Y(new_n8521_));
  AOI21X1  g06085(.A0(new_n8518_), .A1(new_n3035_), .B0(new_n8521_), .Y(new_n8522_));
  NOR2X1   g06086(.A(new_n8522_), .B(new_n8519_), .Y(new_n8523_));
  NOR3X1   g06087(.A(new_n8518_), .B(new_n5928_), .C(new_n2761_), .Y(new_n8524_));
  NOR3X1   g06088(.A(new_n7766_), .B(new_n5881_), .C(new_n7763_), .Y(new_n8525_));
  NOR2X1   g06089(.A(new_n8525_), .B(new_n5882_), .Y(new_n8526_));
  NOR3X1   g06090(.A(new_n8526_), .B(new_n8524_), .C(new_n8522_), .Y(new_n8527_));
  MX2X1    g06091(.A(new_n8527_), .B(new_n8523_), .S0(pi0122), .Y(new_n8528_));
  OR2X1    g06092(.A(new_n8528_), .B(pi1093), .Y(new_n8529_));
  NOR2X1   g06093(.A(new_n8523_), .B(new_n5906_), .Y(new_n8530_));
  AOI21X1  g06094(.A0(new_n8513_), .A1(new_n5906_), .B0(new_n8530_), .Y(new_n8531_));
  OAI21X1  g06095(.A0(new_n8531_), .A1(new_n5032_), .B0(new_n8529_), .Y(new_n8532_));
  AOI21X1  g06096(.A0(new_n8532_), .A1(new_n2703_), .B0(new_n8515_), .Y(new_n8533_));
  OR4X1    g06097(.A(new_n7766_), .B(new_n5881_), .C(new_n7763_), .D(pi0122), .Y(new_n8534_));
  NOR2X1   g06098(.A(new_n8518_), .B(new_n5032_), .Y(new_n8535_));
  OAI21X1  g06099(.A0(new_n8535_), .A1(new_n6243_), .B0(new_n8534_), .Y(new_n8536_));
  AOI21X1  g06100(.A0(new_n8536_), .A1(new_n8529_), .B0(new_n2703_), .Y(new_n8537_));
  NOR2X1   g06101(.A(new_n2703_), .B(pi0137), .Y(new_n8538_));
  NOR2X1   g06102(.A(new_n8538_), .B(new_n8537_), .Y(new_n8539_));
  NAND2X1  g06103(.A(pi1092), .B(pi0252), .Y(new_n8540_));
  NOR2X1   g06104(.A(new_n8540_), .B(pi1093), .Y(new_n8541_));
  INVX1    g06105(.A(new_n8541_), .Y(new_n8542_));
  OAI21X1  g06106(.A0(new_n8542_), .A1(new_n2724_), .B0(new_n2452_), .Y(new_n8543_));
  NOR4X1   g06107(.A(new_n8543_), .B(new_n7766_), .C(new_n5881_), .D(new_n7763_), .Y(new_n8544_));
  OAI22X1  g06108(.A0(new_n8544_), .A1(new_n8539_), .B0(new_n8533_), .B1(new_n8514_), .Y(new_n8545_));
  OR4X1    g06109(.A(new_n7621_), .B(new_n7576_), .C(new_n6757_), .D(new_n2526_), .Y(new_n8546_));
  NOR2X1   g06110(.A(new_n5082_), .B(pi0137), .Y(new_n8547_));
  AOI21X1  g06111(.A0(new_n8546_), .A1(po1057), .B0(new_n8547_), .Y(new_n8548_));
  INVX1    g06112(.A(new_n8548_), .Y(new_n8549_));
  AOI21X1  g06113(.A0(new_n8545_), .A1(new_n5082_), .B0(new_n8549_), .Y(new_n8550_));
  AND2X1   g06114(.A(new_n8532_), .B(new_n2703_), .Y(new_n8551_));
  OR2X1    g06115(.A(new_n8537_), .B(new_n8551_), .Y(new_n8552_));
  MX2X1    g06116(.A(new_n8546_), .B(new_n8552_), .S0(new_n5082_), .Y(new_n8553_));
  INVX1    g06117(.A(new_n8553_), .Y(new_n8554_));
  MX2X1    g06118(.A(new_n8554_), .B(new_n8550_), .S0(new_n2777_), .Y(new_n8555_));
  AND2X1   g06119(.A(new_n7717_), .B(new_n4510_), .Y(new_n8556_));
  MX2X1    g06120(.A(new_n8552_), .B(new_n8545_), .S0(new_n2777_), .Y(new_n8557_));
  AOI21X1  g06121(.A0(new_n8557_), .A1(new_n8556_), .B0(new_n2933_), .Y(new_n8558_));
  OAI21X1  g06122(.A0(new_n8556_), .A1(new_n8555_), .B0(new_n8558_), .Y(new_n8559_));
  MX2X1    g06123(.A(new_n8554_), .B(new_n8550_), .S0(new_n2954_), .Y(new_n8560_));
  AND2X1   g06124(.A(new_n5023_), .B(new_n2961_), .Y(new_n8561_));
  MX2X1    g06125(.A(new_n8552_), .B(new_n8545_), .S0(new_n2954_), .Y(new_n8562_));
  AOI21X1  g06126(.A0(new_n8562_), .A1(new_n8561_), .B0(pi0299), .Y(new_n8563_));
  OAI21X1  g06127(.A0(new_n8561_), .A1(new_n8560_), .B0(new_n8563_), .Y(new_n8564_));
  AOI21X1  g06128(.A0(new_n8564_), .A1(new_n8559_), .B0(new_n5215_), .Y(new_n8565_));
  NOR2X1   g06129(.A(new_n8555_), .B(new_n2933_), .Y(new_n8566_));
  OAI21X1  g06130(.A0(new_n8560_), .A1(pi0299), .B0(new_n5215_), .Y(new_n8567_));
  NOR2X1   g06131(.A(new_n8567_), .B(new_n8566_), .Y(new_n8568_));
  OAI21X1  g06132(.A0(new_n8568_), .A1(new_n8565_), .B0(new_n6072_), .Y(new_n8569_));
  INVX1    g06133(.A(new_n7574_), .Y(new_n8570_));
  INVX1    g06134(.A(new_n8512_), .Y(new_n8571_));
  INVX1    g06135(.A(new_n8519_), .Y(new_n8572_));
  OR2X1    g06136(.A(new_n8525_), .B(new_n2762_), .Y(new_n8573_));
  AND3X1   g06137(.A(new_n8573_), .B(new_n8572_), .C(new_n8571_), .Y(new_n8574_));
  NOR3X1   g06138(.A(new_n8574_), .B(new_n5032_), .C(pi0122), .Y(new_n8575_));
  NOR2X1   g06139(.A(new_n8575_), .B(new_n8530_), .Y(new_n8576_));
  NOR2X1   g06140(.A(new_n8523_), .B(pi1093), .Y(new_n8577_));
  AOI21X1  g06141(.A0(new_n8535_), .A1(new_n2704_), .B0(new_n8577_), .Y(new_n8578_));
  OAI21X1  g06142(.A0(new_n8576_), .A1(new_n2704_), .B0(new_n8578_), .Y(new_n8579_));
  INVX1    g06143(.A(new_n8579_), .Y(new_n8580_));
  AND3X1   g06144(.A(new_n8196_), .B(new_n6753_), .C(po1057), .Y(new_n8581_));
  AOI22X1  g06145(.A0(new_n8581_), .A1(new_n8570_), .B0(new_n8580_), .B1(new_n5082_), .Y(new_n8582_));
  AND2X1   g06146(.A(new_n8196_), .B(new_n6753_), .Y(new_n8583_));
  NOR3X1   g06147(.A(new_n8523_), .B(pi1093), .C(new_n2452_), .Y(new_n8584_));
  NOR3X1   g06148(.A(new_n8574_), .B(pi1093), .C(pi0137), .Y(new_n8585_));
  NOR3X1   g06149(.A(new_n8585_), .B(new_n8584_), .C(new_n8535_), .Y(new_n8586_));
  MX2X1    g06150(.A(new_n8583_), .B(new_n8586_), .S0(new_n5082_), .Y(new_n8587_));
  AOI21X1  g06151(.A0(new_n8547_), .A1(new_n6740_), .B0(new_n2703_), .Y(new_n8588_));
  NOR2X1   g06152(.A(new_n8574_), .B(pi0137), .Y(new_n8589_));
  NOR2X1   g06153(.A(new_n8576_), .B(new_n2452_), .Y(new_n8590_));
  NOR3X1   g06154(.A(new_n8590_), .B(new_n8589_), .C(new_n8584_), .Y(new_n8591_));
  OR2X1    g06155(.A(new_n8591_), .B(po1057), .Y(new_n8592_));
  OAI21X1  g06156(.A0(new_n6243_), .A1(new_n2452_), .B0(new_n2761_), .Y(new_n8593_));
  NAND3X1  g06157(.A(new_n8593_), .B(new_n8196_), .C(new_n6753_), .Y(new_n8594_));
  AOI21X1  g06158(.A0(new_n8594_), .A1(po1057), .B0(new_n2704_), .Y(new_n8595_));
  AOI22X1  g06159(.A0(new_n8595_), .A1(new_n8592_), .B0(new_n8588_), .B1(new_n8587_), .Y(new_n8596_));
  MX2X1    g06160(.A(new_n8596_), .B(new_n8582_), .S0(pi0210), .Y(new_n8597_));
  MX2X1    g06161(.A(new_n8591_), .B(new_n8586_), .S0(new_n2704_), .Y(new_n8598_));
  INVX1    g06162(.A(new_n8556_), .Y(new_n8599_));
  AOI21X1  g06163(.A0(new_n8579_), .A1(pi0210), .B0(new_n8599_), .Y(new_n8600_));
  OAI21X1  g06164(.A0(new_n8598_), .A1(pi0210), .B0(new_n8600_), .Y(new_n8601_));
  AND2X1   g06165(.A(new_n8601_), .B(pi0299), .Y(new_n8602_));
  OAI21X1  g06166(.A0(new_n8597_), .A1(new_n8556_), .B0(new_n8602_), .Y(new_n8603_));
  MX2X1    g06167(.A(new_n8596_), .B(new_n8582_), .S0(pi0198), .Y(new_n8604_));
  MX2X1    g06168(.A(new_n8598_), .B(new_n8580_), .S0(pi0198), .Y(new_n8605_));
  AOI21X1  g06169(.A0(new_n8605_), .A1(new_n8561_), .B0(pi0299), .Y(new_n8606_));
  OAI21X1  g06170(.A0(new_n8604_), .A1(new_n8561_), .B0(new_n8606_), .Y(new_n8607_));
  AOI21X1  g06171(.A0(new_n8607_), .A1(new_n8603_), .B0(new_n5215_), .Y(new_n8608_));
  NOR2X1   g06172(.A(new_n8604_), .B(pi0299), .Y(new_n8609_));
  OAI21X1  g06173(.A0(new_n8597_), .A1(new_n2933_), .B0(new_n5215_), .Y(new_n8610_));
  OAI21X1  g06174(.A0(new_n8610_), .A1(new_n8609_), .B0(new_n6073_), .Y(new_n8611_));
  OR2X1    g06175(.A(new_n8611_), .B(new_n8608_), .Y(new_n8612_));
  AOI21X1  g06176(.A0(new_n8612_), .A1(new_n8569_), .B0(new_n8207_), .Y(po0234));
  OR3X1    g06177(.A(new_n2568_), .B(new_n2559_), .C(new_n2576_), .Y(new_n8614_));
  AND2X1   g06178(.A(new_n8614_), .B(new_n2566_), .Y(new_n8615_));
  NOR3X1   g06179(.A(new_n8615_), .B(new_n5145_), .C(new_n2476_), .Y(new_n8616_));
  INVX1    g06180(.A(new_n8616_), .Y(new_n8617_));
  AND3X1   g06181(.A(new_n6737_), .B(new_n2569_), .C(pi0086), .Y(new_n8618_));
  OAI21X1  g06182(.A0(new_n8618_), .A1(new_n5117_), .B0(new_n7609_), .Y(new_n8619_));
  AOI21X1  g06183(.A0(new_n8617_), .A1(new_n5117_), .B0(new_n8619_), .Y(po0235));
  INVX1    g06184(.A(pi0468), .Y(new_n8621_));
  AND3X1   g06185(.A(new_n8621_), .B(pi0232), .C(pi0119), .Y(po0236));
  INVX1    g06186(.A(pi0163), .Y(new_n8623_));
  OR2X1    g06187(.A(new_n7305_), .B(pi0163), .Y(new_n8624_));
  OAI22X1  g06188(.A0(new_n8624_), .A1(new_n7308_), .B0(new_n7309_), .B1(new_n8623_), .Y(new_n8625_));
  NOR2X1   g06189(.A(new_n8625_), .B(new_n5215_), .Y(new_n8626_));
  AOI21X1  g06190(.A0(new_n3007_), .A1(new_n3073_), .B0(new_n8626_), .Y(new_n8627_));
  AND3X1   g06191(.A(new_n5023_), .B(pi0232), .C(pi0147), .Y(new_n8628_));
  AND2X1   g06192(.A(new_n8628_), .B(new_n6794_), .Y(new_n8629_));
  AOI21X1  g06193(.A0(new_n8626_), .A1(new_n6809_), .B0(new_n4982_), .Y(new_n8630_));
  OR4X1    g06194(.A(new_n8630_), .B(new_n8629_), .C(new_n8627_), .D(new_n3223_), .Y(new_n8631_));
  NOR2X1   g06195(.A(new_n7326_), .B(new_n6803_), .Y(new_n8632_));
  NOR4X1   g06196(.A(new_n7327_), .B(new_n8632_), .C(new_n5048_), .D(pi0184), .Y(new_n8633_));
  INVX1    g06197(.A(pi0184), .Y(new_n8634_));
  NOR3X1   g06198(.A(new_n7327_), .B(new_n8632_), .C(new_n5048_), .Y(new_n8635_));
  NOR3X1   g06199(.A(new_n8635_), .B(new_n5048_), .C(new_n8634_), .Y(new_n8636_));
  NOR3X1   g06200(.A(new_n8636_), .B(new_n8633_), .C(pi0299), .Y(new_n8637_));
  OR2X1    g06201(.A(new_n8637_), .B(new_n5215_), .Y(new_n8638_));
  AOI21X1  g06202(.A0(new_n8625_), .A1(pi0299), .B0(new_n8638_), .Y(new_n8639_));
  AOI21X1  g06203(.A0(new_n8639_), .A1(new_n6809_), .B0(new_n4982_), .Y(new_n8640_));
  NOR2X1   g06204(.A(new_n8640_), .B(pi0055), .Y(new_n8641_));
  MX2X1    g06205(.A(pi0187), .B(pi0147), .S0(pi0299), .Y(new_n8642_));
  AND3X1   g06206(.A(new_n8642_), .B(new_n5023_), .C(pi0232), .Y(new_n8643_));
  OAI21X1  g06207(.A0(new_n8643_), .A1(new_n6809_), .B0(pi0054), .Y(new_n8644_));
  AOI21X1  g06208(.A0(new_n8639_), .A1(new_n6809_), .B0(new_n8644_), .Y(new_n8645_));
  INVX1    g06209(.A(pi0187), .Y(new_n8646_));
  OAI21X1  g06210(.A0(new_n6823_), .A1(new_n8646_), .B0(pi0147), .Y(new_n8647_));
  AOI21X1  g06211(.A0(new_n6822_), .A1(new_n8646_), .B0(new_n8647_), .Y(new_n8648_));
  INVX1    g06212(.A(pi0147), .Y(new_n8649_));
  AND3X1   g06213(.A(new_n6829_), .B(pi0187), .C(new_n8649_), .Y(new_n8650_));
  OAI21X1  g06214(.A0(new_n8650_), .A1(new_n8648_), .B0(pi0038), .Y(new_n8651_));
  OAI21X1  g06215(.A0(new_n6960_), .A1(pi0040), .B0(new_n2523_), .Y(new_n8652_));
  NOR3X1   g06216(.A(new_n6973_), .B(new_n4459_), .C(pi0040), .Y(new_n8653_));
  NOR2X1   g06217(.A(new_n8653_), .B(new_n8652_), .Y(new_n8654_));
  OR2X1    g06218(.A(new_n7001_), .B(new_n5048_), .Y(new_n8655_));
  OAI21X1  g06219(.A0(new_n8655_), .A1(new_n8654_), .B0(new_n2924_), .Y(new_n8656_));
  AND2X1   g06220(.A(new_n7014_), .B(new_n2529_), .Y(new_n8657_));
  OAI21X1  g06221(.A0(new_n8657_), .A1(pi0095), .B0(pi0166), .Y(new_n8658_));
  AOI21X1  g06222(.A0(new_n7717_), .A1(new_n7046_), .B0(new_n2924_), .Y(new_n8659_));
  OAI21X1  g06223(.A0(new_n8658_), .A1(new_n8655_), .B0(new_n8659_), .Y(new_n8660_));
  AND2X1   g06224(.A(new_n8660_), .B(pi0160), .Y(new_n8661_));
  NOR3X1   g06225(.A(new_n8653_), .B(new_n8652_), .C(pi0153), .Y(new_n8662_));
  OR2X1    g06226(.A(new_n7001_), .B(new_n2454_), .Y(new_n8663_));
  OAI21X1  g06227(.A0(new_n6889_), .A1(new_n2469_), .B0(new_n6888_), .Y(new_n8664_));
  AND2X1   g06228(.A(new_n8664_), .B(new_n8663_), .Y(new_n8665_));
  OAI21X1  g06229(.A0(new_n8657_), .A1(pi0095), .B0(new_n8494_), .Y(new_n8666_));
  AND3X1   g06230(.A(new_n8666_), .B(new_n8658_), .C(pi0153), .Y(new_n8667_));
  OR4X1    g06231(.A(new_n8667_), .B(new_n8665_), .C(new_n5048_), .D(pi0160), .Y(new_n8668_));
  OAI21X1  g06232(.A0(new_n8668_), .A1(new_n8662_), .B0(pi0163), .Y(new_n8669_));
  AOI21X1  g06233(.A0(new_n8661_), .A1(new_n8656_), .B0(new_n8669_), .Y(new_n8670_));
  INVX1    g06234(.A(new_n8665_), .Y(new_n8671_));
  NOR2X1   g06235(.A(new_n7067_), .B(pi0040), .Y(new_n8672_));
  OAI21X1  g06236(.A0(new_n8672_), .A1(pi0095), .B0(new_n8671_), .Y(new_n8673_));
  OAI21X1  g06237(.A0(new_n6945_), .A1(pi0040), .B0(new_n2455_), .Y(new_n8674_));
  AOI21X1  g06238(.A0(new_n8674_), .A1(new_n7047_), .B0(pi0095), .Y(new_n8675_));
  OAI21X1  g06239(.A0(new_n8675_), .A1(new_n8665_), .B0(pi0210), .Y(new_n8676_));
  INVX1    g06240(.A(new_n7717_), .Y(new_n8677_));
  AOI21X1  g06241(.A0(new_n8674_), .A1(new_n7004_), .B0(pi0095), .Y(new_n8678_));
  OR2X1    g06242(.A(new_n8678_), .B(new_n8665_), .Y(new_n8679_));
  AOI21X1  g06243(.A0(new_n8679_), .A1(new_n2777_), .B0(new_n8677_), .Y(new_n8680_));
  AOI21X1  g06244(.A0(new_n8680_), .A1(new_n8676_), .B0(pi0153), .Y(new_n8681_));
  OAI21X1  g06245(.A0(new_n8673_), .A1(new_n4459_), .B0(new_n8681_), .Y(new_n8682_));
  OAI21X1  g06246(.A0(new_n6996_), .A1(new_n6990_), .B0(new_n2523_), .Y(new_n8683_));
  AOI21X1  g06247(.A0(new_n8683_), .A1(new_n8671_), .B0(new_n2777_), .Y(new_n8684_));
  AOI21X1  g06248(.A0(new_n8671_), .A1(new_n7006_), .B0(pi0210), .Y(new_n8685_));
  AND2X1   g06249(.A(new_n5023_), .B(pi0166), .Y(new_n8686_));
  INVX1    g06250(.A(new_n8686_), .Y(new_n8687_));
  OR3X1    g06251(.A(new_n8687_), .B(new_n8685_), .C(new_n8684_), .Y(new_n8688_));
  OAI21X1  g06252(.A0(new_n8665_), .A1(new_n7051_), .B0(new_n2777_), .Y(new_n8689_));
  OAI21X1  g06253(.A0(new_n7049_), .A1(pi0095), .B0(new_n8671_), .Y(new_n8690_));
  AOI21X1  g06254(.A0(new_n8690_), .A1(pi0210), .B0(new_n8677_), .Y(new_n8691_));
  AOI21X1  g06255(.A0(new_n8691_), .A1(new_n8689_), .B0(new_n2924_), .Y(new_n8692_));
  AOI21X1  g06256(.A0(new_n8692_), .A1(new_n8688_), .B0(pi0160), .Y(new_n8693_));
  OR2X1    g06257(.A(new_n8678_), .B(new_n7001_), .Y(new_n8694_));
  AND2X1   g06258(.A(new_n8694_), .B(new_n2777_), .Y(new_n8695_));
  OAI21X1  g06259(.A0(new_n8675_), .A1(new_n7001_), .B0(pi0210), .Y(new_n8696_));
  NAND2X1  g06260(.A(new_n8696_), .B(new_n7717_), .Y(new_n8697_));
  OAI21X1  g06261(.A0(new_n8697_), .A1(new_n8695_), .B0(new_n2924_), .Y(new_n8698_));
  AOI21X1  g06262(.A0(new_n8686_), .A1(new_n8672_), .B0(new_n8698_), .Y(new_n8699_));
  NOR2X1   g06263(.A(new_n7050_), .B(new_n2777_), .Y(new_n8700_));
  OAI21X1  g06264(.A0(new_n7052_), .A1(pi0210), .B0(new_n7717_), .Y(new_n8701_));
  NOR2X1   g06265(.A(new_n8701_), .B(new_n8700_), .Y(new_n8702_));
  AOI21X1  g06266(.A0(new_n7006_), .A1(new_n7002_), .B0(pi0210), .Y(new_n8703_));
  AND2X1   g06267(.A(new_n8683_), .B(new_n7002_), .Y(new_n8704_));
  OAI21X1  g06268(.A0(new_n8704_), .A1(new_n2777_), .B0(new_n8686_), .Y(new_n8705_));
  OAI21X1  g06269(.A0(new_n8705_), .A1(new_n8703_), .B0(pi0153), .Y(new_n8706_));
  OAI21X1  g06270(.A0(new_n8706_), .A1(new_n8702_), .B0(pi0160), .Y(new_n8707_));
  OAI21X1  g06271(.A0(new_n8707_), .A1(new_n8699_), .B0(new_n8623_), .Y(new_n8708_));
  AOI21X1  g06272(.A0(new_n8693_), .A1(new_n8682_), .B0(new_n8708_), .Y(new_n8709_));
  OR2X1    g06273(.A(new_n8673_), .B(new_n5023_), .Y(new_n8710_));
  AND2X1   g06274(.A(new_n8710_), .B(pi0299), .Y(new_n8711_));
  OAI21X1  g06275(.A0(new_n8709_), .A1(new_n8670_), .B0(new_n8711_), .Y(new_n8712_));
  OAI21X1  g06276(.A0(new_n6983_), .A1(new_n6937_), .B0(new_n2529_), .Y(new_n8713_));
  AOI21X1  g06277(.A0(new_n8713_), .A1(new_n2523_), .B0(new_n8665_), .Y(new_n8714_));
  NAND2X1  g06278(.A(new_n8714_), .B(new_n5048_), .Y(new_n8715_));
  NOR2X1   g06279(.A(pi0299), .B(pi0175), .Y(new_n8716_));
  INVX1    g06280(.A(new_n8716_), .Y(new_n8717_));
  NOR3X1   g06281(.A(new_n6973_), .B(new_n7872_), .C(pi0040), .Y(new_n8718_));
  AND3X1   g06282(.A(new_n8664_), .B(new_n8663_), .C(new_n5205_), .Y(new_n8719_));
  OAI21X1  g06283(.A0(new_n7002_), .A1(new_n5205_), .B0(new_n5023_), .Y(new_n8720_));
  NOR2X1   g06284(.A(new_n8720_), .B(new_n8719_), .Y(new_n8721_));
  OAI21X1  g06285(.A0(new_n8718_), .A1(new_n8652_), .B0(new_n8721_), .Y(new_n8722_));
  OR3X1    g06286(.A(new_n8713_), .B(new_n5048_), .C(new_n7872_), .Y(new_n8723_));
  OAI21X1  g06287(.A0(new_n8678_), .A1(new_n7001_), .B0(new_n2954_), .Y(new_n8724_));
  OAI21X1  g06288(.A0(new_n8675_), .A1(new_n7001_), .B0(pi0198), .Y(new_n8725_));
  NAND3X1  g06289(.A(new_n8725_), .B(new_n8724_), .C(new_n7714_), .Y(new_n8726_));
  AND3X1   g06290(.A(new_n8726_), .B(new_n8634_), .C(pi0182), .Y(new_n8727_));
  AOI22X1  g06291(.A0(new_n8727_), .A1(new_n8723_), .B0(new_n8722_), .B1(pi0184), .Y(new_n8728_));
  AND2X1   g06292(.A(new_n7714_), .B(new_n7053_), .Y(new_n8729_));
  AOI21X1  g06293(.A0(new_n7006_), .A1(new_n7002_), .B0(pi0198), .Y(new_n8730_));
  AND2X1   g06294(.A(new_n5023_), .B(pi0189), .Y(new_n8731_));
  OAI21X1  g06295(.A0(new_n8704_), .A1(new_n2954_), .B0(new_n8731_), .Y(new_n8732_));
  OAI21X1  g06296(.A0(new_n8732_), .A1(new_n8730_), .B0(pi0182), .Y(new_n8733_));
  AOI21X1  g06297(.A0(new_n8671_), .A1(new_n7006_), .B0(pi0198), .Y(new_n8734_));
  AND2X1   g06298(.A(new_n8683_), .B(new_n8671_), .Y(new_n8735_));
  OAI21X1  g06299(.A0(new_n8735_), .A1(new_n2954_), .B0(new_n8731_), .Y(new_n8736_));
  OAI21X1  g06300(.A0(new_n8736_), .A1(new_n8734_), .B0(new_n5205_), .Y(new_n8737_));
  OAI21X1  g06301(.A0(new_n8733_), .A1(new_n8729_), .B0(new_n8737_), .Y(new_n8738_));
  AND2X1   g06302(.A(new_n5205_), .B(pi0095), .Y(new_n8739_));
  AOI21X1  g06303(.A0(new_n8664_), .A1(new_n8663_), .B0(new_n7873_), .Y(new_n8740_));
  OAI21X1  g06304(.A0(new_n8739_), .A1(new_n7053_), .B0(new_n8740_), .Y(new_n8741_));
  AOI21X1  g06305(.A0(new_n8741_), .A1(new_n8738_), .B0(pi0184), .Y(new_n8742_));
  AND2X1   g06306(.A(new_n2933_), .B(pi0175), .Y(new_n8743_));
  AND2X1   g06307(.A(new_n5023_), .B(pi0184), .Y(new_n8744_));
  OAI21X1  g06308(.A0(new_n7872_), .A1(pi0095), .B0(new_n6895_), .Y(new_n8745_));
  AND3X1   g06309(.A(new_n8745_), .B(new_n7014_), .C(new_n2529_), .Y(new_n8746_));
  OAI21X1  g06310(.A0(new_n8746_), .A1(new_n8739_), .B0(new_n8744_), .Y(new_n8747_));
  OAI21X1  g06311(.A0(new_n8747_), .A1(new_n8719_), .B0(new_n8743_), .Y(new_n8748_));
  OAI22X1  g06312(.A0(new_n8748_), .A1(new_n8742_), .B0(new_n8728_), .B1(new_n8717_), .Y(new_n8749_));
  NAND2X1  g06313(.A(new_n8714_), .B(new_n7873_), .Y(new_n8750_));
  OAI21X1  g06314(.A0(new_n8675_), .A1(new_n8665_), .B0(pi0198), .Y(new_n8751_));
  AOI21X1  g06315(.A0(new_n8679_), .A1(new_n2954_), .B0(new_n7873_), .Y(new_n8752_));
  OR4X1    g06316(.A(pi0299), .B(pi0184), .C(pi0182), .D(pi0175), .Y(new_n8753_));
  AOI21X1  g06317(.A0(new_n8752_), .A1(new_n8751_), .B0(new_n8753_), .Y(new_n8754_));
  AOI22X1  g06318(.A0(new_n8754_), .A1(new_n8750_), .B0(new_n8749_), .B1(new_n8715_), .Y(new_n8755_));
  AOI21X1  g06319(.A0(new_n8755_), .A1(new_n8712_), .B0(new_n5215_), .Y(new_n8756_));
  AND2X1   g06320(.A(new_n8714_), .B(new_n2933_), .Y(new_n8757_));
  OAI21X1  g06321(.A0(new_n8673_), .A1(new_n2933_), .B0(new_n5215_), .Y(new_n8758_));
  OAI21X1  g06322(.A0(new_n8758_), .A1(new_n8757_), .B0(new_n2939_), .Y(new_n8759_));
  NOR2X1   g06323(.A(new_n7046_), .B(new_n6848_), .Y(new_n8760_));
  NOR2X1   g06324(.A(new_n6847_), .B(pi0040), .Y(new_n8761_));
  NOR2X1   g06325(.A(new_n8761_), .B(pi0189), .Y(new_n8762_));
  AOI21X1  g06326(.A0(new_n6867_), .A1(new_n6895_), .B0(new_n6982_), .Y(new_n8763_));
  OAI21X1  g06327(.A0(new_n6846_), .A1(new_n2469_), .B0(new_n2529_), .Y(new_n8764_));
  INVX1    g06328(.A(new_n8764_), .Y(new_n8765_));
  AOI22X1  g06329(.A0(new_n8765_), .A1(new_n6255_), .B0(new_n7046_), .B1(new_n5043_), .Y(new_n8766_));
  INVX1    g06330(.A(new_n8766_), .Y(new_n8767_));
  NOR4X1   g06331(.A(new_n8767_), .B(new_n8763_), .C(new_n5041_), .D(new_n7872_), .Y(new_n8768_));
  OAI21X1  g06332(.A0(new_n8768_), .A1(new_n8762_), .B0(pi0179), .Y(new_n8769_));
  AND2X1   g06333(.A(new_n6843_), .B(new_n5050_), .Y(new_n8770_));
  OAI21X1  g06334(.A0(new_n8770_), .A1(new_n2469_), .B0(new_n6981_), .Y(new_n8771_));
  AOI21X1  g06335(.A0(new_n8771_), .A1(new_n8766_), .B0(pi0189), .Y(new_n8772_));
  INVX1    g06336(.A(new_n7046_), .Y(new_n8773_));
  MX2X1    g06337(.A(new_n8764_), .B(new_n8773_), .S0(new_n5043_), .Y(new_n8774_));
  AOI21X1  g06338(.A0(new_n5040_), .A1(new_n5039_), .B0(pi0179), .Y(new_n8775_));
  OAI21X1  g06339(.A0(new_n8774_), .A1(new_n7872_), .B0(new_n8775_), .Y(new_n8776_));
  OAI22X1  g06340(.A0(new_n8776_), .A1(new_n8772_), .B0(new_n8761_), .B1(new_n5042_), .Y(new_n8777_));
  INVX1    g06341(.A(new_n8777_), .Y(new_n8778_));
  AOI21X1  g06342(.A0(new_n8778_), .A1(new_n8769_), .B0(new_n7203_), .Y(new_n8779_));
  OAI21X1  g06343(.A0(new_n8779_), .A1(new_n8760_), .B0(new_n2933_), .Y(new_n8780_));
  INVX1    g06344(.A(new_n8780_), .Y(new_n8781_));
  OAI21X1  g06345(.A0(new_n8773_), .A1(new_n6856_), .B0(pi0299), .Y(new_n8782_));
  INVX1    g06346(.A(new_n8761_), .Y(new_n8783_));
  MX2X1    g06347(.A(new_n8774_), .B(new_n8783_), .S0(new_n5058_), .Y(new_n8784_));
  OAI21X1  g06348(.A0(new_n5058_), .A1(pi0166), .B0(new_n8784_), .Y(new_n8785_));
  NAND4X1  g06349(.A(new_n8771_), .B(new_n8766_), .C(new_n5059_), .D(new_n4459_), .Y(new_n8786_));
  AND2X1   g06350(.A(new_n8786_), .B(new_n6856_), .Y(new_n8787_));
  AOI21X1  g06351(.A0(new_n8787_), .A1(new_n8785_), .B0(new_n8782_), .Y(new_n8788_));
  INVX1    g06352(.A(pi0156), .Y(new_n8789_));
  AND2X1   g06353(.A(pi0232), .B(new_n8789_), .Y(new_n8790_));
  OAI21X1  g06354(.A0(new_n8788_), .A1(new_n8781_), .B0(new_n8790_), .Y(new_n8791_));
  OR4X1    g06355(.A(new_n8767_), .B(new_n8763_), .C(new_n5058_), .D(new_n4459_), .Y(new_n8792_));
  OAI22X1  g06356(.A0(new_n6847_), .A1(pi0040), .B0(new_n5058_), .B1(new_n4459_), .Y(new_n8793_));
  AND3X1   g06357(.A(new_n8793_), .B(new_n8792_), .C(new_n6856_), .Y(new_n8794_));
  OAI21X1  g06358(.A0(new_n8794_), .A1(new_n8782_), .B0(new_n8780_), .Y(new_n8795_));
  AND2X1   g06359(.A(pi0232), .B(pi0156), .Y(new_n8796_));
  MX2X1    g06360(.A(new_n8774_), .B(new_n8783_), .S0(new_n5041_), .Y(new_n8797_));
  OAI21X1  g06361(.A0(new_n7046_), .A1(new_n6848_), .B0(new_n2933_), .Y(new_n8798_));
  AOI21X1  g06362(.A0(new_n8797_), .A1(new_n6848_), .B0(new_n8798_), .Y(new_n8799_));
  INVX1    g06363(.A(new_n6858_), .Y(new_n8800_));
  OAI21X1  g06364(.A0(new_n8784_), .A1(new_n8800_), .B0(new_n5215_), .Y(new_n8801_));
  OAI21X1  g06365(.A0(new_n8801_), .A1(new_n8799_), .B0(pi0039), .Y(new_n8802_));
  AOI21X1  g06366(.A0(new_n8796_), .A1(new_n8795_), .B0(new_n8802_), .Y(new_n8803_));
  AOI21X1  g06367(.A0(new_n8803_), .A1(new_n8791_), .B0(pi0038), .Y(new_n8804_));
  OAI21X1  g06368(.A0(new_n8759_), .A1(new_n8756_), .B0(new_n8804_), .Y(new_n8805_));
  AOI21X1  g06369(.A0(new_n8805_), .A1(new_n8651_), .B0(new_n7156_), .Y(new_n8806_));
  OAI21X1  g06370(.A0(new_n8643_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n8807_));
  NOR2X1   g06371(.A(pi0040), .B(pi0038), .Y(new_n8808_));
  AND3X1   g06372(.A(new_n8808_), .B(new_n2469_), .C(pi0087), .Y(new_n8809_));
  OR2X1    g06373(.A(new_n8809_), .B(new_n8807_), .Y(new_n8810_));
  OAI22X1  g06374(.A0(new_n8810_), .A1(new_n3131_), .B0(new_n8639_), .B1(new_n3007_), .Y(new_n8811_));
  OAI21X1  g06375(.A0(new_n8811_), .A1(new_n8806_), .B0(new_n3084_), .Y(new_n8812_));
  NOR2X1   g06376(.A(new_n8639_), .B(new_n3073_), .Y(new_n8813_));
  OR2X1    g06377(.A(new_n8639_), .B(new_n3007_), .Y(new_n8814_));
  OAI21X1  g06378(.A0(new_n7046_), .A1(new_n2939_), .B0(new_n7280_), .Y(new_n8815_));
  AOI21X1  g06379(.A0(new_n7142_), .A1(new_n6895_), .B0(pi0040), .Y(new_n8816_));
  MX2X1    g06380(.A(pi0179), .B(pi0156), .S0(pi0299), .Y(new_n8817_));
  NAND3X1  g06381(.A(new_n8817_), .B(new_n5023_), .C(pi0232), .Y(new_n8818_));
  OAI21X1  g06382(.A0(new_n8818_), .A1(new_n2469_), .B0(new_n8816_), .Y(new_n8819_));
  AOI21X1  g06383(.A0(new_n8819_), .A1(new_n2939_), .B0(new_n8815_), .Y(new_n8820_));
  OAI21X1  g06384(.A0(new_n8820_), .A1(new_n8810_), .B0(new_n8814_), .Y(new_n8821_));
  AOI21X1  g06385(.A0(new_n8821_), .A1(new_n7138_), .B0(new_n8813_), .Y(new_n8822_));
  AOI21X1  g06386(.A0(new_n8822_), .A1(new_n8812_), .B0(pi0054), .Y(new_n8823_));
  OAI21X1  g06387(.A0(new_n8823_), .A1(new_n8645_), .B0(new_n4982_), .Y(new_n8824_));
  OR2X1    g06388(.A(new_n8630_), .B(new_n3107_), .Y(new_n8825_));
  OAI21X1  g06389(.A0(new_n8629_), .A1(new_n8627_), .B0(pi0054), .Y(new_n8826_));
  OAI21X1  g06390(.A0(new_n8625_), .A1(new_n5215_), .B0(pi0100), .Y(new_n8827_));
  NAND2X1  g06391(.A(pi0232), .B(pi0163), .Y(new_n8828_));
  OAI21X1  g06392(.A0(new_n7142_), .A1(new_n5023_), .B0(new_n6834_), .Y(new_n8829_));
  OAI21X1  g06393(.A0(new_n8829_), .A1(new_n8828_), .B0(new_n8816_), .Y(new_n8830_));
  AOI21X1  g06394(.A0(new_n8830_), .A1(new_n2939_), .B0(new_n8815_), .Y(new_n8831_));
  OAI21X1  g06395(.A0(new_n8628_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n8832_));
  OR3X1    g06396(.A(new_n8832_), .B(new_n8831_), .C(new_n8809_), .Y(new_n8833_));
  AOI21X1  g06397(.A0(new_n8833_), .A1(new_n8827_), .B0(new_n5295_), .Y(new_n8834_));
  OAI21X1  g06398(.A0(new_n8832_), .A1(new_n8808_), .B0(new_n8827_), .Y(new_n8835_));
  OAI21X1  g06399(.A0(new_n8835_), .A1(new_n7139_), .B0(new_n7138_), .Y(new_n8836_));
  OAI21X1  g06400(.A0(new_n8626_), .A1(new_n3073_), .B0(new_n8836_), .Y(new_n8837_));
  OAI21X1  g06401(.A0(new_n8837_), .A1(new_n8834_), .B0(new_n3091_), .Y(new_n8838_));
  AOI21X1  g06402(.A0(new_n8838_), .A1(new_n8826_), .B0(pi0074), .Y(new_n8839_));
  OAI21X1  g06403(.A0(new_n8839_), .A1(new_n8825_), .B0(new_n3123_), .Y(new_n8840_));
  AOI21X1  g06404(.A0(new_n8824_), .A1(new_n8641_), .B0(new_n8840_), .Y(new_n8841_));
  NOR2X1   g06405(.A(new_n8626_), .B(new_n3073_), .Y(new_n8842_));
  AOI21X1  g06406(.A0(new_n8835_), .A1(new_n3073_), .B0(new_n8842_), .Y(new_n8843_));
  OAI21X1  g06407(.A0(new_n8843_), .A1(pi0054), .B0(new_n8826_), .Y(new_n8844_));
  AOI21X1  g06408(.A0(new_n8844_), .A1(new_n4982_), .B0(new_n8630_), .Y(new_n8845_));
  OAI21X1  g06409(.A0(new_n8845_), .A1(new_n3123_), .B0(new_n3223_), .Y(new_n8846_));
  OR2X1    g06410(.A(new_n8846_), .B(new_n7181_), .Y(new_n8847_));
  OAI21X1  g06411(.A0(new_n8847_), .A1(new_n8841_), .B0(new_n8631_), .Y(new_n8848_));
  NOR2X1   g06412(.A(new_n8848_), .B(pi0079), .Y(new_n8849_));
  INVX1    g06413(.A(pi0160), .Y(new_n8850_));
  INVX1    g06414(.A(new_n2527_), .Y(new_n8851_));
  NOR4X1   g06415(.A(new_n8851_), .B(pi0479), .C(new_n2523_), .D(pi0032), .Y(new_n8852_));
  OR4X1    g06416(.A(new_n8852_), .B(new_n7221_), .C(new_n5175_), .D(pi0040), .Y(new_n8853_));
  AND2X1   g06417(.A(new_n8853_), .B(new_n7717_), .Y(new_n8854_));
  NOR2X1   g06418(.A(new_n7234_), .B(new_n7217_), .Y(new_n8855_));
  NOR4X1   g06419(.A(new_n8852_), .B(new_n8855_), .C(new_n5175_), .D(pi0040), .Y(new_n8856_));
  OAI21X1  g06420(.A0(new_n8856_), .A1(new_n8687_), .B0(new_n2924_), .Y(new_n8857_));
  OAI21X1  g06421(.A0(new_n7221_), .A1(new_n7220_), .B0(new_n2777_), .Y(new_n8858_));
  NOR3X1   g06422(.A(new_n8852_), .B(new_n7218_), .C(pi0040), .Y(new_n8859_));
  AOI21X1  g06423(.A0(new_n8859_), .A1(new_n8858_), .B0(new_n8677_), .Y(new_n8860_));
  AOI21X1  g06424(.A0(new_n8856_), .A1(new_n7489_), .B0(new_n8687_), .Y(new_n8861_));
  OR2X1    g06425(.A(new_n8861_), .B(new_n2924_), .Y(new_n8862_));
  OAI22X1  g06426(.A0(new_n8862_), .A1(new_n8860_), .B0(new_n8857_), .B1(new_n8854_), .Y(new_n8863_));
  OAI21X1  g06427(.A0(pi0468), .A1(pi0332), .B0(pi0040), .Y(new_n8864_));
  AND2X1   g06428(.A(new_n8864_), .B(pi0163), .Y(new_n8865_));
  AOI21X1  g06429(.A0(new_n8865_), .A1(new_n8863_), .B0(new_n8850_), .Y(new_n8866_));
  AOI21X1  g06430(.A0(new_n7218_), .A1(pi0153), .B0(new_n7487_), .Y(new_n8867_));
  OAI21X1  g06431(.A0(new_n7489_), .A1(new_n2924_), .B0(new_n7263_), .Y(new_n8868_));
  OR2X1    g06432(.A(new_n8623_), .B(pi0040), .Y(new_n8869_));
  AOI21X1  g06433(.A0(new_n8868_), .A1(new_n8686_), .B0(new_n8869_), .Y(new_n8870_));
  OAI21X1  g06434(.A0(new_n8867_), .A1(new_n8677_), .B0(new_n8870_), .Y(new_n8871_));
  AND3X1   g06435(.A(new_n5023_), .B(new_n7228_), .C(pi0153), .Y(new_n8872_));
  NOR3X1   g06436(.A(new_n8677_), .B(new_n7251_), .C(new_n7250_), .Y(new_n8873_));
  OR3X1    g06437(.A(new_n8873_), .B(pi0163), .C(pi0040), .Y(new_n8874_));
  AOI21X1  g06438(.A0(new_n8872_), .A1(new_n7238_), .B0(new_n8874_), .Y(new_n8875_));
  NOR2X1   g06439(.A(new_n8875_), .B(pi0160), .Y(new_n8876_));
  AND2X1   g06440(.A(new_n8876_), .B(new_n8871_), .Y(new_n8877_));
  NAND2X1  g06441(.A(new_n8852_), .B(new_n5023_), .Y(new_n8878_));
  AOI21X1  g06442(.A0(new_n8878_), .A1(new_n8875_), .B0(new_n2933_), .Y(new_n8879_));
  OAI21X1  g06443(.A0(new_n8877_), .A1(new_n8866_), .B0(new_n8879_), .Y(new_n8880_));
  OR3X1    g06444(.A(new_n7221_), .B(new_n5198_), .C(new_n8634_), .Y(new_n8881_));
  OAI21X1  g06445(.A0(new_n7251_), .A1(new_n7250_), .B0(new_n8634_), .Y(new_n8882_));
  AND2X1   g06446(.A(new_n8882_), .B(new_n7872_), .Y(new_n8883_));
  NAND2X1  g06447(.A(new_n8852_), .B(pi0182), .Y(new_n8884_));
  NAND2X1  g06448(.A(pi0189), .B(pi0184), .Y(new_n8885_));
  OAI21X1  g06449(.A0(new_n8885_), .A1(new_n7246_), .B0(new_n8884_), .Y(new_n8886_));
  AOI21X1  g06450(.A0(new_n8883_), .A1(new_n8881_), .B0(new_n8886_), .Y(new_n8887_));
  OAI21X1  g06451(.A0(new_n8887_), .A1(new_n5048_), .B0(new_n2529_), .Y(new_n8888_));
  NOR2X1   g06452(.A(new_n7238_), .B(new_n7872_), .Y(new_n8889_));
  OAI21X1  g06453(.A0(new_n7227_), .A1(pi0189), .B0(new_n7228_), .Y(new_n8890_));
  OAI21X1  g06454(.A0(new_n8890_), .A1(new_n8889_), .B0(new_n8884_), .Y(new_n8891_));
  AOI21X1  g06455(.A0(new_n8891_), .A1(new_n5023_), .B0(pi0184), .Y(new_n8892_));
  AND3X1   g06456(.A(new_n7236_), .B(new_n5023_), .C(pi0189), .Y(new_n8893_));
  OR3X1    g06457(.A(new_n8893_), .B(new_n8634_), .C(pi0182), .Y(new_n8894_));
  AOI21X1  g06458(.A0(new_n7714_), .A1(new_n7223_), .B0(new_n8894_), .Y(new_n8895_));
  OAI21X1  g06459(.A0(new_n8895_), .A1(new_n8892_), .B0(new_n2529_), .Y(new_n8896_));
  INVX1    g06460(.A(new_n8743_), .Y(new_n8897_));
  OAI21X1  g06461(.A0(new_n7222_), .A1(pi0198), .B0(new_n8859_), .Y(new_n8898_));
  NAND2X1  g06462(.A(new_n8898_), .B(new_n7714_), .Y(new_n8899_));
  OR4X1    g06463(.A(new_n8852_), .B(new_n7235_), .C(new_n5198_), .D(pi0040), .Y(new_n8900_));
  NAND3X1  g06464(.A(new_n8864_), .B(pi0184), .C(pi0182), .Y(new_n8901_));
  AOI21X1  g06465(.A0(new_n8900_), .A1(new_n8731_), .B0(new_n8901_), .Y(new_n8902_));
  AOI21X1  g06466(.A0(new_n8902_), .A1(new_n8899_), .B0(new_n8897_), .Y(new_n8903_));
  AOI22X1  g06467(.A0(new_n8903_), .A1(new_n8896_), .B0(new_n8888_), .B1(new_n8716_), .Y(new_n8904_));
  AOI21X1  g06468(.A0(new_n8904_), .A1(new_n8880_), .B0(pi0039), .Y(new_n8905_));
  NAND3X1  g06469(.A(new_n5023_), .B(new_n7228_), .C(new_n2527_), .Y(new_n8906_));
  AOI22X1  g06470(.A0(new_n6844_), .A1(new_n4459_), .B0(new_n5050_), .B1(pi0156), .Y(new_n8907_));
  OR4X1    g06471(.A(new_n8907_), .B(new_n8906_), .C(new_n7187_), .D(new_n5058_), .Y(new_n8908_));
  AND3X1   g06472(.A(new_n8908_), .B(pi0299), .C(new_n2529_), .Y(new_n8909_));
  AOI22X1  g06473(.A0(new_n6844_), .A1(new_n7872_), .B0(new_n5050_), .B1(pi0179), .Y(new_n8910_));
  NOR4X1   g06474(.A(new_n8910_), .B(new_n8906_), .C(new_n7203_), .D(new_n5041_), .Y(new_n8911_));
  OR2X1    g06475(.A(pi0299), .B(pi0040), .Y(new_n8912_));
  OAI21X1  g06476(.A0(new_n8912_), .A1(new_n8911_), .B0(pi0039), .Y(new_n8913_));
  OAI21X1  g06477(.A0(new_n8913_), .A1(new_n8909_), .B0(pi0232), .Y(new_n8914_));
  AOI21X1  g06478(.A0(new_n5215_), .A1(new_n2529_), .B0(pi0038), .Y(new_n8915_));
  OAI21X1  g06479(.A0(new_n8914_), .A1(new_n8905_), .B0(new_n8915_), .Y(new_n8916_));
  AOI21X1  g06480(.A0(new_n8916_), .A1(new_n8651_), .B0(new_n7156_), .Y(new_n8917_));
  OAI21X1  g06481(.A0(pi0040), .A1(pi0038), .B0(pi0087), .Y(new_n8918_));
  OAI22X1  g06482(.A0(new_n8918_), .A1(new_n8807_), .B0(new_n8639_), .B1(new_n3007_), .Y(new_n8919_));
  OAI21X1  g06483(.A0(new_n8919_), .A1(new_n8917_), .B0(new_n3084_), .Y(new_n8920_));
  INVX1    g06484(.A(new_n8808_), .Y(new_n8921_));
  NOR3X1   g06485(.A(new_n8818_), .B(new_n7141_), .C(new_n7250_), .Y(new_n8922_));
  AOI21X1  g06486(.A0(new_n8922_), .A1(new_n2527_), .B0(new_n8921_), .Y(new_n8923_));
  OAI21X1  g06487(.A0(new_n8923_), .A1(new_n8807_), .B0(new_n8814_), .Y(new_n8924_));
  AOI21X1  g06488(.A0(new_n8924_), .A1(new_n7138_), .B0(new_n8813_), .Y(new_n8925_));
  AOI21X1  g06489(.A0(new_n8925_), .A1(new_n8920_), .B0(pi0054), .Y(new_n8926_));
  OAI21X1  g06490(.A0(new_n8926_), .A1(new_n8645_), .B0(new_n4982_), .Y(new_n8927_));
  OR4X1    g06491(.A(new_n8906_), .B(new_n8828_), .C(new_n7141_), .D(pi0092), .Y(new_n8928_));
  OR2X1    g06492(.A(new_n8832_), .B(pi0075), .Y(new_n8929_));
  AOI21X1  g06493(.A0(new_n8928_), .A1(new_n8808_), .B0(new_n8929_), .Y(new_n8930_));
  OAI21X1  g06494(.A0(new_n8930_), .A1(new_n8627_), .B0(new_n3091_), .Y(new_n8931_));
  AOI21X1  g06495(.A0(new_n8931_), .A1(new_n8826_), .B0(pi0074), .Y(new_n8932_));
  OAI21X1  g06496(.A0(new_n8932_), .A1(new_n8825_), .B0(new_n3123_), .Y(new_n8933_));
  AOI21X1  g06497(.A0(new_n8927_), .A1(new_n8641_), .B0(new_n8933_), .Y(new_n8934_));
  OAI21X1  g06498(.A0(new_n8934_), .A1(new_n8846_), .B0(new_n8631_), .Y(new_n8935_));
  OAI22X1  g06499(.A0(new_n8935_), .A1(new_n6784_), .B0(new_n7548_), .B1(pi0034), .Y(new_n8936_));
  AOI21X1  g06500(.A0(new_n6786_), .A1(new_n6785_), .B0(pi0079), .Y(new_n8937_));
  NOR2X1   g06501(.A(new_n8937_), .B(new_n8848_), .Y(new_n8938_));
  NOR3X1   g06502(.A(pi0954), .B(pi0034), .C(pi0033), .Y(new_n8939_));
  INVX1    g06503(.A(new_n8937_), .Y(new_n8940_));
  OAI21X1  g06504(.A0(new_n8940_), .A1(new_n8935_), .B0(new_n8939_), .Y(new_n8941_));
  OAI22X1  g06505(.A0(new_n8941_), .A1(new_n8938_), .B0(new_n8936_), .B1(new_n8849_), .Y(po0237));
  INVX1    g06506(.A(new_n6713_), .Y(new_n8943_));
  AND2X1   g06507(.A(pi1092), .B(pi0098), .Y(new_n8944_));
  AOI22X1  g06508(.A0(new_n8944_), .A1(pi1093), .B0(new_n2720_), .B1(new_n5979_), .Y(new_n8945_));
  AOI21X1  g06509(.A0(new_n8945_), .A1(new_n6562_), .B0(new_n6603_), .Y(new_n8946_));
  INVX1    g06510(.A(new_n8946_), .Y(new_n8947_));
  NOR2X1   g06511(.A(new_n8945_), .B(new_n6009_), .Y(new_n8948_));
  AOI21X1  g06512(.A0(new_n2720_), .A1(new_n5979_), .B0(new_n6295_), .Y(new_n8949_));
  NAND3X1  g06513(.A(pi1093), .B(pi1092), .C(pi0098), .Y(new_n8950_));
  NOR2X1   g06514(.A(new_n8950_), .B(new_n2702_), .Y(new_n8951_));
  OR3X1    g06515(.A(new_n7769_), .B(new_n2472_), .C(pi0088), .Y(new_n8952_));
  OR3X1    g06516(.A(new_n8952_), .B(new_n2475_), .C(pi0110), .Y(new_n8953_));
  OR4X1    g06517(.A(new_n8953_), .B(new_n5892_), .C(new_n2567_), .D(pi0094), .Y(new_n8954_));
  NOR4X1   g06518(.A(new_n8954_), .B(new_n5898_), .C(pi0070), .D(new_n2534_), .Y(new_n8955_));
  AND2X1   g06519(.A(pi0093), .B(pi0090), .Y(new_n8956_));
  OR4X1    g06520(.A(new_n8956_), .B(new_n5172_), .C(new_n2483_), .D(pi0841), .Y(new_n8957_));
  NOR2X1   g06521(.A(new_n8957_), .B(new_n8954_), .Y(new_n8958_));
  AND2X1   g06522(.A(pi0950), .B(pi0824), .Y(new_n8959_));
  AND3X1   g06523(.A(new_n8959_), .B(new_n2984_), .C(new_n2513_), .Y(new_n8960_));
  OAI21X1  g06524(.A0(new_n8958_), .A1(new_n8955_), .B0(new_n8960_), .Y(new_n8961_));
  AOI21X1  g06525(.A0(new_n8961_), .A1(new_n5893_), .B0(new_n5024_), .Y(new_n8962_));
  OAI21X1  g06526(.A0(new_n8944_), .A1(new_n2702_), .B0(pi1093), .Y(new_n8963_));
  NOR2X1   g06527(.A(new_n8963_), .B(new_n3074_), .Y(new_n8964_));
  OAI21X1  g06528(.A0(new_n8962_), .A1(new_n8951_), .B0(new_n8964_), .Y(new_n8965_));
  INVX1    g06529(.A(new_n8951_), .Y(new_n8966_));
  NAND4X1  g06530(.A(new_n8959_), .B(new_n2984_), .C(new_n2513_), .D(new_n2534_), .Y(new_n8967_));
  NOR4X1   g06531(.A(new_n8967_), .B(new_n8954_), .C(new_n5898_), .D(pi0070), .Y(new_n8968_));
  OAI21X1  g06532(.A0(new_n8968_), .A1(pi0098), .B0(pi1092), .Y(new_n8969_));
  AND2X1   g06533(.A(new_n8969_), .B(new_n8966_), .Y(new_n8970_));
  NOR2X1   g06534(.A(new_n8963_), .B(new_n5986_), .Y(new_n8971_));
  INVX1    g06535(.A(new_n8971_), .Y(new_n8972_));
  OR2X1    g06536(.A(new_n8972_), .B(new_n8970_), .Y(new_n8973_));
  OR2X1    g06537(.A(new_n8950_), .B(new_n3064_), .Y(new_n8974_));
  AND3X1   g06538(.A(new_n8974_), .B(new_n8973_), .C(new_n8965_), .Y(new_n8975_));
  MX2X1    g06539(.A(new_n8975_), .B(new_n8950_), .S0(pi0075), .Y(new_n8976_));
  OR2X1    g06540(.A(new_n8976_), .B(new_n5979_), .Y(new_n8977_));
  AOI22X1  g06541(.A0(new_n8977_), .A1(new_n8949_), .B0(new_n8945_), .B1(new_n6295_), .Y(new_n8978_));
  AOI21X1  g06542(.A0(new_n8978_), .A1(new_n6009_), .B0(new_n8948_), .Y(new_n8979_));
  INVX1    g06543(.A(new_n8979_), .Y(new_n8980_));
  NOR2X1   g06544(.A(new_n8945_), .B(pi1196), .Y(new_n8981_));
  NOR2X1   g06545(.A(new_n8981_), .B(new_n6518_), .Y(new_n8982_));
  INVX1    g06546(.A(pi0429), .Y(new_n8983_));
  INVX1    g06547(.A(pi0443), .Y(new_n8984_));
  MX2X1    g06548(.A(new_n8979_), .B(new_n8945_), .S0(new_n8984_), .Y(new_n8985_));
  INVX1    g06549(.A(new_n8985_), .Y(new_n8986_));
  MX2X1    g06550(.A(new_n8979_), .B(new_n8945_), .S0(pi0443), .Y(new_n8987_));
  INVX1    g06551(.A(new_n8987_), .Y(new_n8988_));
  MX2X1    g06552(.A(new_n8988_), .B(new_n8986_), .S0(new_n6567_), .Y(new_n8989_));
  AOI21X1  g06553(.A0(new_n8985_), .A1(pi0444), .B0(pi0436), .Y(new_n8990_));
  OAI21X1  g06554(.A0(new_n8988_), .A1(pi0444), .B0(new_n8990_), .Y(new_n8991_));
  AOI21X1  g06555(.A0(new_n8987_), .A1(pi0444), .B0(new_n6527_), .Y(new_n8992_));
  OAI21X1  g06556(.A0(new_n8986_), .A1(pi0444), .B0(new_n8992_), .Y(new_n8993_));
  AND2X1   g06557(.A(new_n8993_), .B(new_n8991_), .Y(new_n8994_));
  INVX1    g06558(.A(new_n8994_), .Y(new_n8995_));
  MX2X1    g06559(.A(new_n8995_), .B(new_n8989_), .S0(pi0435), .Y(new_n8996_));
  NAND2X1  g06560(.A(new_n8996_), .B(new_n8983_), .Y(new_n8997_));
  INVX1    g06561(.A(pi0435), .Y(new_n8998_));
  MX2X1    g06562(.A(new_n8995_), .B(new_n8989_), .S0(new_n8998_), .Y(new_n8999_));
  AOI21X1  g06563(.A0(new_n8999_), .A1(pi0429), .B0(new_n6532_), .Y(new_n9000_));
  AND2X1   g06564(.A(new_n9000_), .B(new_n8997_), .Y(new_n9001_));
  AND2X1   g06565(.A(new_n8999_), .B(new_n8983_), .Y(new_n9002_));
  AND2X1   g06566(.A(new_n8996_), .B(pi0429), .Y(new_n9003_));
  NOR3X1   g06567(.A(new_n9003_), .B(new_n9002_), .C(new_n6533_), .Y(new_n9004_));
  OR3X1    g06568(.A(new_n9004_), .B(new_n9001_), .C(new_n6045_), .Y(new_n9005_));
  AOI22X1  g06569(.A0(new_n9005_), .A1(new_n8982_), .B0(new_n8979_), .B1(new_n6518_), .Y(new_n9006_));
  MX2X1    g06570(.A(new_n9006_), .B(new_n8980_), .S0(pi0428), .Y(new_n9007_));
  MX2X1    g06571(.A(new_n9006_), .B(new_n8980_), .S0(new_n6497_), .Y(new_n9008_));
  MX2X1    g06572(.A(new_n9008_), .B(new_n9007_), .S0(new_n6496_), .Y(new_n9009_));
  MX2X1    g06573(.A(new_n9008_), .B(new_n9007_), .S0(pi0427), .Y(new_n9010_));
  MX2X1    g06574(.A(new_n9010_), .B(new_n9009_), .S0(pi0430), .Y(new_n9011_));
  MX2X1    g06575(.A(new_n9010_), .B(new_n9009_), .S0(new_n6550_), .Y(new_n9012_));
  MX2X1    g06576(.A(new_n9012_), .B(new_n9011_), .S0(pi0426), .Y(new_n9013_));
  MX2X1    g06577(.A(new_n9012_), .B(new_n9011_), .S0(new_n6553_), .Y(new_n9014_));
  MX2X1    g06578(.A(new_n9014_), .B(new_n9013_), .S0(pi0445), .Y(new_n9015_));
  NAND2X1  g06579(.A(new_n9015_), .B(pi0448), .Y(new_n9016_));
  MX2X1    g06580(.A(new_n9014_), .B(new_n9013_), .S0(new_n6557_), .Y(new_n9017_));
  AOI21X1  g06581(.A0(new_n9017_), .A1(new_n6491_), .B0(new_n6591_), .Y(new_n9018_));
  NAND2X1  g06582(.A(new_n9018_), .B(new_n9016_), .Y(new_n9019_));
  NAND2X1  g06583(.A(new_n9017_), .B(pi0448), .Y(new_n9020_));
  AOI21X1  g06584(.A0(new_n9015_), .A1(new_n6491_), .B0(new_n6494_), .Y(new_n9021_));
  AOI21X1  g06585(.A0(new_n9021_), .A1(new_n9020_), .B0(new_n6053_), .Y(new_n9022_));
  AND2X1   g06586(.A(new_n9006_), .B(new_n6053_), .Y(new_n9023_));
  OR2X1    g06587(.A(new_n9023_), .B(new_n6562_), .Y(new_n9024_));
  AOI21X1  g06588(.A0(new_n9022_), .A1(new_n9019_), .B0(new_n9024_), .Y(new_n9025_));
  INVX1    g06589(.A(new_n8945_), .Y(new_n9026_));
  AOI21X1  g06590(.A0(new_n9026_), .A1(pi0591), .B0(new_n6334_), .Y(new_n9027_));
  NOR2X1   g06591(.A(new_n6620_), .B(new_n6023_), .Y(new_n9028_));
  MX2X1    g06592(.A(new_n8979_), .B(new_n8945_), .S0(new_n9028_), .Y(new_n9029_));
  NOR2X1   g06593(.A(new_n8981_), .B(pi1198), .Y(new_n9030_));
  INVX1    g06594(.A(new_n9030_), .Y(new_n9031_));
  MX2X1    g06595(.A(new_n9026_), .B(new_n8980_), .S0(new_n6014_), .Y(new_n9032_));
  MX2X1    g06596(.A(new_n8979_), .B(new_n8945_), .S0(pi0455), .Y(new_n9033_));
  MX2X1    g06597(.A(new_n8979_), .B(new_n8945_), .S0(new_n6032_), .Y(new_n9034_));
  MX2X1    g06598(.A(new_n9034_), .B(new_n9033_), .S0(new_n6030_), .Y(new_n9035_));
  INVX1    g06599(.A(new_n9035_), .Y(new_n9036_));
  MX2X1    g06600(.A(new_n9036_), .B(new_n9032_), .S0(pi0355), .Y(new_n9037_));
  NAND2X1  g06601(.A(new_n9037_), .B(new_n6029_), .Y(new_n9038_));
  MX2X1    g06602(.A(new_n9036_), .B(new_n9032_), .S0(new_n6013_), .Y(new_n9039_));
  AOI21X1  g06603(.A0(new_n9039_), .A1(pi0458), .B0(new_n6020_), .Y(new_n9040_));
  NAND2X1  g06604(.A(new_n9040_), .B(new_n9038_), .Y(new_n9041_));
  NAND2X1  g06605(.A(new_n9039_), .B(new_n6029_), .Y(new_n9042_));
  AOI21X1  g06606(.A0(new_n9037_), .A1(pi0458), .B0(new_n6028_), .Y(new_n9043_));
  AOI21X1  g06607(.A0(new_n9043_), .A1(new_n9042_), .B0(new_n6045_), .Y(new_n9044_));
  AOI21X1  g06608(.A0(new_n9044_), .A1(new_n9041_), .B0(new_n9031_), .Y(new_n9045_));
  AOI21X1  g06609(.A0(new_n9029_), .A1(pi1198), .B0(new_n9045_), .Y(new_n9046_));
  MX2X1    g06610(.A(new_n9046_), .B(new_n8980_), .S0(new_n5879_), .Y(new_n9047_));
  NOR2X1   g06611(.A(new_n8979_), .B(new_n6053_), .Y(new_n9048_));
  AOI22X1  g06612(.A0(new_n9048_), .A1(pi0351), .B0(new_n9047_), .B1(new_n6057_), .Y(new_n9049_));
  AOI22X1  g06613(.A0(new_n9048_), .A1(new_n6050_), .B0(new_n9047_), .B1(new_n6052_), .Y(new_n9050_));
  MX2X1    g06614(.A(new_n9050_), .B(new_n9049_), .S0(new_n5866_), .Y(new_n9051_));
  MX2X1    g06615(.A(new_n9050_), .B(new_n9049_), .S0(pi0461), .Y(new_n9052_));
  MX2X1    g06616(.A(new_n9052_), .B(new_n9051_), .S0(new_n5865_), .Y(new_n9053_));
  MX2X1    g06617(.A(new_n9052_), .B(new_n9051_), .S0(pi0357), .Y(new_n9054_));
  MX2X1    g06618(.A(new_n9054_), .B(new_n9053_), .S0(new_n5864_), .Y(new_n9055_));
  NOR2X1   g06619(.A(new_n9055_), .B(pi0354), .Y(new_n9056_));
  INVX1    g06620(.A(pi0354), .Y(new_n9057_));
  MX2X1    g06621(.A(new_n9054_), .B(new_n9053_), .S0(pi0356), .Y(new_n9058_));
  OAI21X1  g06622(.A0(new_n9058_), .A1(new_n9057_), .B0(new_n5862_), .Y(new_n9059_));
  NOR2X1   g06623(.A(new_n9059_), .B(new_n9056_), .Y(new_n9060_));
  NOR2X1   g06624(.A(new_n9058_), .B(pi0354), .Y(new_n9061_));
  INVX1    g06625(.A(new_n5862_), .Y(new_n9062_));
  OAI21X1  g06626(.A0(new_n9055_), .A1(new_n9057_), .B0(new_n9062_), .Y(new_n9063_));
  OAI21X1  g06627(.A0(new_n9063_), .A1(new_n9061_), .B0(new_n6069_), .Y(new_n9064_));
  OAI21X1  g06628(.A0(new_n9064_), .A1(new_n9060_), .B0(new_n9027_), .Y(new_n9065_));
  AOI21X1  g06629(.A0(new_n6172_), .A1(pi1198), .B0(pi1197), .Y(new_n9066_));
  AOI21X1  g06630(.A0(new_n8945_), .A1(new_n6295_), .B0(new_n6364_), .Y(new_n9067_));
  INVX1    g06631(.A(new_n8962_), .Y(new_n9068_));
  AOI21X1  g06632(.A0(new_n8944_), .A1(new_n6174_), .B0(new_n6181_), .Y(new_n9069_));
  OAI21X1  g06633(.A0(new_n9068_), .A1(new_n6174_), .B0(new_n9069_), .Y(new_n9070_));
  INVX1    g06634(.A(new_n8944_), .Y(new_n9071_));
  OAI21X1  g06635(.A0(new_n9071_), .A1(new_n6174_), .B0(new_n6181_), .Y(new_n9072_));
  AND2X1   g06636(.A(new_n8962_), .B(new_n6174_), .Y(new_n9073_));
  OAI21X1  g06637(.A0(new_n9073_), .A1(new_n9072_), .B0(new_n9070_), .Y(new_n9074_));
  NAND2X1  g06638(.A(new_n9074_), .B(new_n8966_), .Y(new_n9075_));
  OAI21X1  g06639(.A0(new_n8969_), .A1(new_n6174_), .B0(new_n9069_), .Y(new_n9076_));
  INVX1    g06640(.A(new_n9072_), .Y(new_n9077_));
  OAI21X1  g06641(.A0(new_n8969_), .A1(pi0411), .B0(new_n9077_), .Y(new_n9078_));
  AOI21X1  g06642(.A0(new_n9078_), .A1(new_n9076_), .B0(new_n8951_), .Y(new_n9079_));
  OAI21X1  g06643(.A0(new_n9079_), .A1(new_n8972_), .B0(new_n8974_), .Y(new_n9080_));
  AOI21X1  g06644(.A0(new_n9075_), .A1(new_n8964_), .B0(new_n9080_), .Y(new_n9081_));
  MX2X1    g06645(.A(new_n9081_), .B(new_n8950_), .S0(pi0075), .Y(new_n9082_));
  OAI21X1  g06646(.A0(new_n9082_), .A1(new_n5979_), .B0(new_n8949_), .Y(new_n9083_));
  OR3X1    g06647(.A(new_n8981_), .B(new_n8948_), .C(pi1199), .Y(new_n9084_));
  AOI21X1  g06648(.A0(new_n9083_), .A1(new_n9067_), .B0(new_n9084_), .Y(new_n9085_));
  INVX1    g06649(.A(new_n9067_), .Y(new_n9086_));
  OR3X1    g06650(.A(new_n8972_), .B(new_n8970_), .C(new_n6202_), .Y(new_n9087_));
  MX2X1    g06651(.A(new_n9068_), .B(new_n9071_), .S0(new_n6202_), .Y(new_n9088_));
  NOR2X1   g06652(.A(new_n9088_), .B(new_n8965_), .Y(new_n9089_));
  INVX1    g06653(.A(new_n9089_), .Y(new_n9090_));
  AND3X1   g06654(.A(new_n9090_), .B(new_n9087_), .C(new_n9081_), .Y(new_n9091_));
  MX2X1    g06655(.A(new_n8969_), .B(new_n9071_), .S0(new_n6202_), .Y(new_n9092_));
  OAI21X1  g06656(.A0(new_n9092_), .A1(new_n8973_), .B0(new_n8974_), .Y(new_n9093_));
  AOI21X1  g06657(.A0(new_n8945_), .A1(new_n6295_), .B0(new_n6427_), .Y(new_n9094_));
  OAI21X1  g06658(.A0(new_n9093_), .A1(new_n9089_), .B0(new_n9094_), .Y(new_n9095_));
  OAI21X1  g06659(.A0(new_n9091_), .A1(new_n9086_), .B0(new_n9095_), .Y(new_n9096_));
  AND2X1   g06660(.A(pi0567), .B(new_n3073_), .Y(new_n9097_));
  AOI21X1  g06661(.A0(new_n8949_), .A1(new_n6187_), .B0(new_n8945_), .Y(new_n9098_));
  OR2X1    g06662(.A(new_n9098_), .B(new_n6053_), .Y(new_n9099_));
  AOI21X1  g06663(.A0(new_n9097_), .A1(new_n9096_), .B0(new_n9099_), .Y(new_n9100_));
  OR3X1    g06664(.A(new_n9100_), .B(new_n9085_), .C(new_n6173_), .Y(new_n9101_));
  OAI22X1  g06665(.A0(new_n9101_), .A1(pi1197), .B0(new_n9066_), .B1(new_n8979_), .Y(new_n9102_));
  AND2X1   g06666(.A(new_n9102_), .B(new_n6162_), .Y(new_n9103_));
  OAI21X1  g06667(.A0(new_n8979_), .A1(new_n6451_), .B0(new_n9101_), .Y(new_n9104_));
  AOI21X1  g06668(.A0(new_n9104_), .A1(pi0333), .B0(new_n9103_), .Y(new_n9105_));
  OR2X1    g06669(.A(new_n9105_), .B(pi0391), .Y(new_n9106_));
  AND2X1   g06670(.A(new_n9102_), .B(pi0333), .Y(new_n9107_));
  AOI21X1  g06671(.A0(new_n9104_), .A1(new_n6162_), .B0(new_n9107_), .Y(new_n9108_));
  OAI21X1  g06672(.A0(new_n9108_), .A1(new_n6219_), .B0(new_n9106_), .Y(new_n9109_));
  AND2X1   g06673(.A(new_n9109_), .B(new_n6161_), .Y(new_n9110_));
  OR2X1    g06674(.A(new_n9108_), .B(pi0391), .Y(new_n9111_));
  OAI21X1  g06675(.A0(new_n9105_), .A1(new_n6219_), .B0(new_n9111_), .Y(new_n9112_));
  AOI21X1  g06676(.A0(new_n9112_), .A1(pi0392), .B0(new_n9110_), .Y(new_n9113_));
  NOR2X1   g06677(.A(new_n9113_), .B(pi0393), .Y(new_n9114_));
  AND2X1   g06678(.A(new_n9112_), .B(new_n6161_), .Y(new_n9115_));
  AOI21X1  g06679(.A0(new_n9109_), .A1(pi0392), .B0(new_n9115_), .Y(new_n9116_));
  OAI21X1  g06680(.A0(new_n9116_), .A1(new_n6160_), .B0(new_n6677_), .Y(new_n9117_));
  NOR2X1   g06681(.A(new_n9117_), .B(new_n9114_), .Y(new_n9118_));
  NOR2X1   g06682(.A(new_n9116_), .B(pi0393), .Y(new_n9119_));
  OAI21X1  g06683(.A0(new_n9113_), .A1(new_n6160_), .B0(new_n6361_), .Y(new_n9120_));
  OAI21X1  g06684(.A0(new_n9120_), .A1(new_n9119_), .B0(pi0591), .Y(new_n9121_));
  MX2X1    g06685(.A(new_n8978_), .B(new_n9026_), .S0(new_n6009_), .Y(new_n9122_));
  AOI21X1  g06686(.A0(new_n8945_), .A1(new_n6643_), .B0(new_n6053_), .Y(new_n9123_));
  OAI21X1  g06687(.A0(new_n9122_), .A1(new_n6643_), .B0(new_n9123_), .Y(new_n9124_));
  AOI22X1  g06688(.A0(new_n9026_), .A1(new_n5876_), .B0(new_n6087_), .B1(pi1196), .Y(new_n9125_));
  XOR2X1   g06689(.A(new_n6096_), .B(new_n6089_), .Y(new_n9126_));
  XOR2X1   g06690(.A(new_n9126_), .B(pi0367), .Y(new_n9127_));
  AOI21X1  g06691(.A0(new_n9127_), .A1(new_n8945_), .B0(new_n5876_), .Y(new_n9128_));
  OAI21X1  g06692(.A0(new_n9127_), .A1(new_n9122_), .B0(new_n9128_), .Y(new_n9129_));
  AND2X1   g06693(.A(new_n9129_), .B(new_n9125_), .Y(new_n9130_));
  INVX1    g06694(.A(new_n6088_), .Y(new_n9131_));
  OAI21X1  g06695(.A0(new_n9122_), .A1(new_n9131_), .B0(new_n6053_), .Y(new_n9132_));
  OAI21X1  g06696(.A0(new_n9132_), .A1(new_n9130_), .B0(new_n9124_), .Y(new_n9133_));
  MX2X1    g06697(.A(new_n9133_), .B(new_n9122_), .S0(pi1198), .Y(new_n9134_));
  MX2X1    g06698(.A(new_n9134_), .B(new_n9133_), .S0(new_n6079_), .Y(new_n9135_));
  NAND2X1  g06699(.A(new_n9135_), .B(new_n6078_), .Y(new_n9136_));
  XOR2X1   g06700(.A(new_n6338_), .B(pi0371), .Y(new_n9137_));
  XOR2X1   g06701(.A(new_n9137_), .B(new_n6077_), .Y(new_n9138_));
  MX2X1    g06702(.A(new_n9134_), .B(new_n9133_), .S0(pi0374), .Y(new_n9139_));
  AOI21X1  g06703(.A0(new_n9139_), .A1(pi0369), .B0(new_n9138_), .Y(new_n9140_));
  NAND2X1  g06704(.A(new_n9140_), .B(new_n9136_), .Y(new_n9141_));
  NAND2X1  g06705(.A(new_n9135_), .B(pi0369), .Y(new_n9142_));
  INVX1    g06706(.A(new_n9138_), .Y(new_n9143_));
  AOI21X1  g06707(.A0(new_n9139_), .A1(new_n6078_), .B0(new_n9143_), .Y(new_n9144_));
  AOI21X1  g06708(.A0(new_n9144_), .A1(new_n9142_), .B0(pi0591), .Y(new_n9145_));
  AOI21X1  g06709(.A0(new_n9145_), .A1(new_n9141_), .B0(pi0590), .Y(new_n9146_));
  OAI21X1  g06710(.A0(new_n9121_), .A1(new_n9118_), .B0(new_n9146_), .Y(new_n9147_));
  AND2X1   g06711(.A(new_n9147_), .B(new_n6603_), .Y(new_n9148_));
  AOI21X1  g06712(.A0(new_n9148_), .A1(new_n9065_), .B0(new_n6073_), .Y(new_n9149_));
  OAI21X1  g06713(.A0(new_n9025_), .A1(new_n8947_), .B0(new_n9149_), .Y(new_n9150_));
  INVX1    g06714(.A(new_n8948_), .Y(new_n9151_));
  AOI22X1  g06715(.A0(new_n8944_), .A1(pi1093), .B0(new_n6246_), .B1(new_n2702_), .Y(new_n9152_));
  AOI21X1  g06716(.A0(new_n9152_), .A1(new_n5906_), .B0(new_n5968_), .Y(new_n9153_));
  OAI21X1  g06717(.A0(new_n8950_), .A1(new_n2702_), .B0(new_n3064_), .Y(new_n9154_));
  NOR2X1   g06718(.A(new_n9154_), .B(pi0087), .Y(new_n9155_));
  NOR2X1   g06719(.A(new_n9154_), .B(new_n3131_), .Y(new_n9156_));
  AOI22X1  g06720(.A0(new_n9156_), .A1(new_n8969_), .B0(new_n9155_), .B1(new_n9068_), .Y(new_n9157_));
  OAI22X1  g06721(.A0(new_n9157_), .A1(new_n5906_), .B0(new_n9154_), .B1(new_n9153_), .Y(new_n9158_));
  AND2X1   g06722(.A(new_n5880_), .B(pi0567), .Y(new_n9159_));
  OAI21X1  g06723(.A0(new_n3378_), .A1(pi0075), .B0(new_n9152_), .Y(new_n9160_));
  NAND2X1  g06724(.A(new_n9160_), .B(new_n9159_), .Y(new_n9161_));
  AOI21X1  g06725(.A0(new_n9158_), .A1(new_n3073_), .B0(new_n9161_), .Y(new_n9162_));
  OAI22X1  g06726(.A0(new_n9152_), .A1(new_n5880_), .B0(new_n2725_), .B1(pi0567), .Y(new_n9163_));
  OAI21X1  g06727(.A0(new_n9163_), .A1(new_n9162_), .B0(new_n6009_), .Y(new_n9164_));
  AND2X1   g06728(.A(new_n9164_), .B(new_n9151_), .Y(new_n9165_));
  INVX1    g06729(.A(new_n9165_), .Y(new_n9166_));
  MX2X1    g06730(.A(new_n9165_), .B(new_n8945_), .S0(new_n8984_), .Y(new_n9167_));
  INVX1    g06731(.A(new_n9167_), .Y(new_n9168_));
  MX2X1    g06732(.A(new_n9165_), .B(new_n8945_), .S0(pi0443), .Y(new_n9169_));
  INVX1    g06733(.A(new_n9169_), .Y(new_n9170_));
  MX2X1    g06734(.A(new_n9170_), .B(new_n9168_), .S0(new_n6567_), .Y(new_n9171_));
  NAND2X1  g06735(.A(new_n9169_), .B(new_n6520_), .Y(new_n9172_));
  AOI21X1  g06736(.A0(new_n9167_), .A1(pi0444), .B0(pi0436), .Y(new_n9173_));
  NAND2X1  g06737(.A(new_n9167_), .B(new_n6520_), .Y(new_n9174_));
  AOI21X1  g06738(.A0(new_n9169_), .A1(pi0444), .B0(new_n6527_), .Y(new_n9175_));
  AOI22X1  g06739(.A0(new_n9175_), .A1(new_n9174_), .B0(new_n9173_), .B1(new_n9172_), .Y(new_n9176_));
  INVX1    g06740(.A(new_n9176_), .Y(new_n9177_));
  MX2X1    g06741(.A(new_n9177_), .B(new_n9171_), .S0(pi0435), .Y(new_n9178_));
  NAND2X1  g06742(.A(new_n9178_), .B(new_n8983_), .Y(new_n9179_));
  MX2X1    g06743(.A(new_n9177_), .B(new_n9171_), .S0(new_n8998_), .Y(new_n9180_));
  AOI21X1  g06744(.A0(new_n9180_), .A1(pi0429), .B0(new_n6532_), .Y(new_n9181_));
  AND2X1   g06745(.A(new_n9181_), .B(new_n9179_), .Y(new_n9182_));
  AND2X1   g06746(.A(new_n9180_), .B(new_n8983_), .Y(new_n9183_));
  AND2X1   g06747(.A(new_n9178_), .B(pi0429), .Y(new_n9184_));
  NOR3X1   g06748(.A(new_n9184_), .B(new_n9183_), .C(new_n6533_), .Y(new_n9185_));
  NOR3X1   g06749(.A(new_n9185_), .B(new_n9182_), .C(new_n6045_), .Y(new_n9186_));
  NOR3X1   g06750(.A(new_n9186_), .B(new_n8981_), .C(new_n6518_), .Y(new_n9187_));
  AOI21X1  g06751(.A0(new_n9165_), .A1(new_n6518_), .B0(new_n9187_), .Y(new_n9188_));
  MX2X1    g06752(.A(new_n9188_), .B(new_n9166_), .S0(new_n6497_), .Y(new_n9189_));
  MX2X1    g06753(.A(new_n9188_), .B(new_n9166_), .S0(pi0428), .Y(new_n9190_));
  MX2X1    g06754(.A(new_n9190_), .B(new_n9189_), .S0(new_n6496_), .Y(new_n9191_));
  MX2X1    g06755(.A(new_n9190_), .B(new_n9189_), .S0(pi0427), .Y(new_n9192_));
  MX2X1    g06756(.A(new_n9192_), .B(new_n9191_), .S0(pi0430), .Y(new_n9193_));
  MX2X1    g06757(.A(new_n9192_), .B(new_n9191_), .S0(new_n6550_), .Y(new_n9194_));
  MX2X1    g06758(.A(new_n9194_), .B(new_n9193_), .S0(pi0426), .Y(new_n9195_));
  MX2X1    g06759(.A(new_n9194_), .B(new_n9193_), .S0(new_n6553_), .Y(new_n9196_));
  MX2X1    g06760(.A(new_n9196_), .B(new_n9195_), .S0(pi0445), .Y(new_n9197_));
  OR2X1    g06761(.A(new_n9196_), .B(new_n6557_), .Y(new_n9198_));
  OAI21X1  g06762(.A0(new_n9195_), .A1(pi0445), .B0(new_n9198_), .Y(new_n9199_));
  OAI21X1  g06763(.A0(new_n9199_), .A1(pi0448), .B0(new_n6591_), .Y(new_n9200_));
  AOI21X1  g06764(.A0(new_n9197_), .A1(pi0448), .B0(new_n9200_), .Y(new_n9201_));
  AND2X1   g06765(.A(new_n9197_), .B(new_n6491_), .Y(new_n9202_));
  OAI21X1  g06766(.A0(new_n9199_), .A1(new_n6491_), .B0(new_n6494_), .Y(new_n9203_));
  OAI21X1  g06767(.A0(new_n9203_), .A1(new_n9202_), .B0(pi1199), .Y(new_n9204_));
  AOI21X1  g06768(.A0(new_n9188_), .A1(new_n6053_), .B0(new_n6562_), .Y(new_n9205_));
  OAI21X1  g06769(.A0(new_n9204_), .A1(new_n9201_), .B0(new_n9205_), .Y(new_n9206_));
  MX2X1    g06770(.A(new_n9166_), .B(new_n9026_), .S0(new_n9028_), .Y(new_n9207_));
  MX2X1    g06771(.A(new_n9026_), .B(new_n9166_), .S0(new_n6014_), .Y(new_n9208_));
  MX2X1    g06772(.A(new_n9165_), .B(new_n8945_), .S0(pi0455), .Y(new_n9209_));
  MX2X1    g06773(.A(new_n9165_), .B(new_n8945_), .S0(new_n6032_), .Y(new_n9210_));
  MX2X1    g06774(.A(new_n9210_), .B(new_n9209_), .S0(new_n6030_), .Y(new_n9211_));
  INVX1    g06775(.A(new_n9211_), .Y(new_n9212_));
  MX2X1    g06776(.A(new_n9212_), .B(new_n9208_), .S0(new_n6013_), .Y(new_n9213_));
  NAND2X1  g06777(.A(new_n9213_), .B(new_n6029_), .Y(new_n9214_));
  MX2X1    g06778(.A(new_n9212_), .B(new_n9208_), .S0(pi0355), .Y(new_n9215_));
  AOI21X1  g06779(.A0(new_n9215_), .A1(pi0458), .B0(new_n6028_), .Y(new_n9216_));
  NAND2X1  g06780(.A(new_n9216_), .B(new_n9214_), .Y(new_n9217_));
  NAND2X1  g06781(.A(new_n9215_), .B(new_n6029_), .Y(new_n9218_));
  AOI21X1  g06782(.A0(new_n9213_), .A1(pi0458), .B0(new_n6020_), .Y(new_n9219_));
  AOI21X1  g06783(.A0(new_n9219_), .A1(new_n9218_), .B0(new_n6045_), .Y(new_n9220_));
  AND2X1   g06784(.A(new_n9220_), .B(new_n9217_), .Y(new_n9221_));
  OAI22X1  g06785(.A0(new_n9221_), .A1(new_n9031_), .B0(new_n9207_), .B1(new_n6025_), .Y(new_n9222_));
  MX2X1    g06786(.A(new_n9222_), .B(new_n9165_), .S0(new_n5879_), .Y(new_n9223_));
  INVX1    g06787(.A(new_n9223_), .Y(new_n9224_));
  AOI21X1  g06788(.A0(new_n9164_), .A1(new_n9151_), .B0(new_n6053_), .Y(new_n9225_));
  AOI22X1  g06789(.A0(new_n9225_), .A1(pi0351), .B0(new_n9224_), .B1(new_n6057_), .Y(new_n9226_));
  AOI22X1  g06790(.A0(new_n9225_), .A1(new_n6050_), .B0(new_n9224_), .B1(new_n6052_), .Y(new_n9227_));
  MX2X1    g06791(.A(new_n9227_), .B(new_n9226_), .S0(new_n5866_), .Y(new_n9228_));
  MX2X1    g06792(.A(new_n9227_), .B(new_n9226_), .S0(pi0461), .Y(new_n9229_));
  MX2X1    g06793(.A(new_n9229_), .B(new_n9228_), .S0(new_n5865_), .Y(new_n9230_));
  MX2X1    g06794(.A(new_n9229_), .B(new_n9228_), .S0(pi0357), .Y(new_n9231_));
  MX2X1    g06795(.A(new_n9231_), .B(new_n9230_), .S0(new_n5864_), .Y(new_n9232_));
  NOR2X1   g06796(.A(new_n9232_), .B(pi0354), .Y(new_n9233_));
  MX2X1    g06797(.A(new_n9231_), .B(new_n9230_), .S0(pi0356), .Y(new_n9234_));
  OAI21X1  g06798(.A0(new_n9234_), .A1(new_n9057_), .B0(new_n5862_), .Y(new_n9235_));
  OR2X1    g06799(.A(new_n9235_), .B(new_n9233_), .Y(new_n9236_));
  OR2X1    g06800(.A(new_n9234_), .B(pi0354), .Y(new_n9237_));
  OR2X1    g06801(.A(new_n9232_), .B(new_n9057_), .Y(new_n9238_));
  NAND3X1  g06802(.A(new_n9238_), .B(new_n9237_), .C(new_n9062_), .Y(new_n9239_));
  NAND3X1  g06803(.A(new_n9239_), .B(new_n9236_), .C(new_n6069_), .Y(new_n9240_));
  NOR2X1   g06804(.A(new_n9163_), .B(new_n9162_), .Y(new_n9241_));
  MX2X1    g06805(.A(new_n9241_), .B(new_n8945_), .S0(new_n6009_), .Y(new_n9242_));
  INVX1    g06806(.A(new_n9242_), .Y(new_n9243_));
  MX2X1    g06807(.A(new_n9243_), .B(new_n9026_), .S0(pi0367), .Y(new_n9244_));
  MX2X1    g06808(.A(new_n9243_), .B(new_n9026_), .S0(new_n6090_), .Y(new_n9245_));
  MX2X1    g06809(.A(new_n9245_), .B(new_n9244_), .S0(new_n6089_), .Y(new_n9246_));
  AND2X1   g06810(.A(new_n9246_), .B(new_n6092_), .Y(new_n9247_));
  MX2X1    g06811(.A(new_n9244_), .B(new_n9245_), .S0(new_n6089_), .Y(new_n9248_));
  AND2X1   g06812(.A(new_n9248_), .B(new_n6091_), .Y(new_n9249_));
  NOR3X1   g06813(.A(new_n9249_), .B(new_n9247_), .C(new_n6095_), .Y(new_n9250_));
  NAND2X1  g06814(.A(new_n9246_), .B(new_n6091_), .Y(new_n9251_));
  NAND2X1  g06815(.A(new_n9248_), .B(new_n6092_), .Y(new_n9252_));
  AND3X1   g06816(.A(new_n9252_), .B(new_n9251_), .C(new_n6095_), .Y(new_n9253_));
  OR2X1    g06817(.A(new_n9253_), .B(new_n5876_), .Y(new_n9254_));
  OAI21X1  g06818(.A0(new_n9254_), .A1(new_n9250_), .B0(new_n9125_), .Y(new_n9255_));
  AOI21X1  g06819(.A0(new_n9242_), .A1(new_n6088_), .B0(pi1199), .Y(new_n9256_));
  MX2X1    g06820(.A(new_n9243_), .B(new_n9026_), .S0(new_n6643_), .Y(new_n9257_));
  AOI22X1  g06821(.A0(new_n9257_), .A1(pi1199), .B0(new_n9256_), .B1(new_n9255_), .Y(new_n9258_));
  AND3X1   g06822(.A(new_n9256_), .B(new_n9255_), .C(new_n6025_), .Y(new_n9259_));
  AOI22X1  g06823(.A0(new_n9257_), .A1(new_n6129_), .B0(new_n9243_), .B1(pi1198), .Y(new_n9260_));
  INVX1    g06824(.A(new_n9260_), .Y(new_n9261_));
  NOR2X1   g06825(.A(new_n9261_), .B(new_n9259_), .Y(new_n9262_));
  MX2X1    g06826(.A(new_n9262_), .B(new_n9258_), .S0(new_n6079_), .Y(new_n9263_));
  OAI21X1  g06827(.A0(new_n9261_), .A1(new_n9259_), .B0(new_n6079_), .Y(new_n9264_));
  OAI21X1  g06828(.A0(new_n9258_), .A1(new_n6079_), .B0(new_n9264_), .Y(new_n9265_));
  AOI21X1  g06829(.A0(new_n9265_), .A1(new_n6078_), .B0(new_n9143_), .Y(new_n9266_));
  OAI21X1  g06830(.A0(new_n9263_), .A1(new_n6078_), .B0(new_n9266_), .Y(new_n9267_));
  AOI21X1  g06831(.A0(new_n9265_), .A1(pi0369), .B0(new_n9138_), .Y(new_n9268_));
  OAI21X1  g06832(.A0(new_n9263_), .A1(pi0369), .B0(new_n9268_), .Y(new_n9269_));
  AND3X1   g06833(.A(new_n9269_), .B(new_n9267_), .C(new_n6069_), .Y(new_n9270_));
  INVX1    g06834(.A(new_n9066_), .Y(new_n9271_));
  INVX1    g06835(.A(new_n8981_), .Y(new_n9272_));
  INVX1    g06836(.A(pi0412), .Y(new_n9273_));
  XOR2X1   g06837(.A(pi0404), .B(pi0397), .Y(new_n9274_));
  XOR2X1   g06838(.A(new_n9274_), .B(pi0411), .Y(new_n9275_));
  XOR2X1   g06839(.A(new_n9275_), .B(new_n6175_), .Y(new_n9276_));
  OAI21X1  g06840(.A0(new_n9276_), .A1(new_n5928_), .B0(new_n9071_), .Y(new_n9277_));
  AOI21X1  g06841(.A0(new_n9276_), .A1(new_n5927_), .B0(new_n8944_), .Y(new_n9278_));
  OAI21X1  g06842(.A0(new_n9278_), .A1(new_n9273_), .B0(new_n6179_), .Y(new_n9279_));
  AOI21X1  g06843(.A0(new_n9277_), .A1(new_n9273_), .B0(new_n9279_), .Y(new_n9280_));
  INVX1    g06844(.A(new_n6179_), .Y(new_n9281_));
  OAI21X1  g06845(.A0(new_n9278_), .A1(pi0412), .B0(new_n9281_), .Y(new_n9282_));
  AOI21X1  g06846(.A0(new_n9277_), .A1(pi0412), .B0(new_n9282_), .Y(new_n9283_));
  NOR3X1   g06847(.A(new_n9283_), .B(new_n9280_), .C(pi0122), .Y(new_n9284_));
  INVX1    g06848(.A(new_n9284_), .Y(new_n9285_));
  AOI21X1  g06849(.A0(new_n9285_), .A1(new_n9071_), .B0(new_n5968_), .Y(new_n9286_));
  NOR2X1   g06850(.A(new_n9286_), .B(new_n8951_), .Y(new_n9287_));
  MX2X1    g06851(.A(new_n9287_), .B(new_n2725_), .S0(new_n5979_), .Y(new_n9288_));
  NOR2X1   g06852(.A(new_n9288_), .B(new_n8949_), .Y(new_n9289_));
  INVX1    g06853(.A(new_n9155_), .Y(new_n9290_));
  OAI21X1  g06854(.A0(new_n9074_), .A1(new_n5906_), .B0(new_n9285_), .Y(new_n9291_));
  AND2X1   g06855(.A(new_n9291_), .B(new_n5967_), .Y(new_n9292_));
  AND3X1   g06856(.A(new_n9078_), .B(new_n9076_), .C(pi0122), .Y(new_n9293_));
  OAI21X1  g06857(.A0(new_n9293_), .A1(new_n9284_), .B0(new_n5967_), .Y(new_n9294_));
  AOI22X1  g06858(.A0(new_n9294_), .A1(new_n9156_), .B0(new_n9287_), .B1(new_n3132_), .Y(new_n9295_));
  OAI21X1  g06859(.A0(new_n9292_), .A1(new_n9290_), .B0(new_n9295_), .Y(new_n9296_));
  INVX1    g06860(.A(new_n9287_), .Y(new_n9297_));
  OAI21X1  g06861(.A0(new_n9297_), .A1(new_n3073_), .B0(new_n9159_), .Y(new_n9298_));
  AOI21X1  g06862(.A0(new_n9296_), .A1(new_n3073_), .B0(new_n9298_), .Y(new_n9299_));
  OAI21X1  g06863(.A0(new_n9299_), .A1(new_n9289_), .B0(new_n6363_), .Y(new_n9300_));
  AOI21X1  g06864(.A0(new_n9300_), .A1(new_n9272_), .B0(pi1199), .Y(new_n9301_));
  AOI21X1  g06865(.A0(new_n5927_), .A1(new_n5906_), .B0(new_n8944_), .Y(new_n9302_));
  OR2X1    g06866(.A(new_n6202_), .B(new_n5928_), .Y(new_n9303_));
  AND3X1   g06867(.A(new_n9303_), .B(new_n9071_), .C(new_n5906_), .Y(new_n9304_));
  OR3X1    g06868(.A(new_n9304_), .B(new_n9302_), .C(new_n8963_), .Y(new_n9305_));
  MX2X1    g06869(.A(new_n9305_), .B(new_n2725_), .S0(new_n5979_), .Y(new_n9306_));
  INVX1    g06870(.A(new_n9306_), .Y(new_n9307_));
  AOI21X1  g06871(.A0(new_n9297_), .A1(pi0567), .B0(new_n9307_), .Y(new_n9308_));
  NOR2X1   g06872(.A(new_n9308_), .B(new_n8949_), .Y(new_n9309_));
  OAI21X1  g06873(.A0(new_n9304_), .A1(new_n8963_), .B0(new_n3064_), .Y(new_n9310_));
  AND2X1   g06874(.A(new_n9078_), .B(new_n9076_), .Y(new_n9311_));
  INVX1    g06875(.A(new_n9311_), .Y(new_n9312_));
  AND2X1   g06876(.A(new_n9155_), .B(new_n9088_), .Y(new_n9313_));
  INVX1    g06877(.A(new_n6181_), .Y(new_n9314_));
  OAI21X1  g06878(.A0(new_n9073_), .A1(new_n9314_), .B0(new_n9070_), .Y(new_n9315_));
  OR2X1    g06879(.A(new_n8969_), .B(new_n6202_), .Y(new_n9316_));
  AND2X1   g06880(.A(new_n9156_), .B(new_n9316_), .Y(new_n9317_));
  AOI22X1  g06881(.A0(new_n9317_), .A1(new_n9312_), .B0(new_n9315_), .B1(new_n9313_), .Y(new_n9318_));
  OAI21X1  g06882(.A0(new_n9303_), .A1(pi0122), .B0(new_n9285_), .Y(new_n9319_));
  OAI22X1  g06883(.A0(new_n9319_), .A1(new_n9318_), .B0(new_n9310_), .B1(new_n9286_), .Y(new_n9320_));
  OAI21X1  g06884(.A0(new_n3378_), .A1(pi0075), .B0(new_n9305_), .Y(new_n9321_));
  OAI21X1  g06885(.A0(new_n9321_), .A1(new_n9286_), .B0(new_n9159_), .Y(new_n9322_));
  AOI21X1  g06886(.A0(new_n9320_), .A1(new_n3073_), .B0(new_n9322_), .Y(new_n9323_));
  OAI21X1  g06887(.A0(new_n9323_), .A1(new_n9309_), .B0(new_n6363_), .Y(new_n9324_));
  NOR2X1   g06888(.A(new_n9306_), .B(new_n8949_), .Y(new_n9325_));
  AOI22X1  g06889(.A0(new_n9156_), .A1(new_n9092_), .B0(new_n9155_), .B1(new_n9088_), .Y(new_n9326_));
  OAI21X1  g06890(.A0(new_n9326_), .A1(new_n5906_), .B0(new_n9310_), .Y(new_n9327_));
  NAND2X1  g06891(.A(new_n9321_), .B(new_n9159_), .Y(new_n9328_));
  AOI21X1  g06892(.A0(new_n9327_), .A1(new_n3073_), .B0(new_n9328_), .Y(new_n9329_));
  OAI21X1  g06893(.A0(new_n9329_), .A1(new_n9325_), .B0(new_n6426_), .Y(new_n9330_));
  AOI21X1  g06894(.A0(new_n9330_), .A1(new_n9324_), .B0(new_n6053_), .Y(new_n9331_));
  NOR4X1   g06895(.A(new_n9331_), .B(new_n9301_), .C(new_n9271_), .D(new_n8948_), .Y(new_n9332_));
  AOI21X1  g06896(.A0(new_n9165_), .A1(new_n9271_), .B0(new_n9332_), .Y(new_n9333_));
  NOR3X1   g06897(.A(new_n9331_), .B(new_n9301_), .C(new_n8948_), .Y(new_n9334_));
  MX2X1    g06898(.A(new_n9334_), .B(new_n9165_), .S0(new_n6173_), .Y(new_n9335_));
  INVX1    g06899(.A(new_n9335_), .Y(new_n9336_));
  MX2X1    g06900(.A(new_n9336_), .B(new_n9333_), .S0(pi0333), .Y(new_n9337_));
  MX2X1    g06901(.A(new_n9336_), .B(new_n9333_), .S0(new_n6162_), .Y(new_n9338_));
  MX2X1    g06902(.A(new_n9338_), .B(new_n9337_), .S0(pi0391), .Y(new_n9339_));
  MX2X1    g06903(.A(new_n9338_), .B(new_n9337_), .S0(new_n6219_), .Y(new_n9340_));
  MX2X1    g06904(.A(new_n9340_), .B(new_n9339_), .S0(pi0392), .Y(new_n9341_));
  MX2X1    g06905(.A(new_n9340_), .B(new_n9339_), .S0(new_n6161_), .Y(new_n9342_));
  MX2X1    g06906(.A(new_n9342_), .B(new_n9341_), .S0(pi0393), .Y(new_n9343_));
  NOR2X1   g06907(.A(new_n9343_), .B(new_n6361_), .Y(new_n9344_));
  MX2X1    g06908(.A(new_n9342_), .B(new_n9341_), .S0(new_n6160_), .Y(new_n9345_));
  OAI21X1  g06909(.A0(new_n9345_), .A1(new_n6677_), .B0(pi0591), .Y(new_n9346_));
  OAI21X1  g06910(.A0(new_n9346_), .A1(new_n9344_), .B0(new_n6334_), .Y(new_n9347_));
  OAI21X1  g06911(.A0(new_n9347_), .A1(new_n9270_), .B0(new_n6603_), .Y(new_n9348_));
  AOI21X1  g06912(.A0(new_n9240_), .A1(new_n9027_), .B0(new_n9348_), .Y(new_n9349_));
  OR2X1    g06913(.A(new_n9349_), .B(new_n6072_), .Y(new_n9350_));
  AOI21X1  g06914(.A0(new_n9206_), .A1(new_n8946_), .B0(new_n9350_), .Y(new_n9351_));
  NOR3X1   g06915(.A(new_n9351_), .B(po1038), .C(pi0080), .Y(new_n9352_));
  INVX1    g06916(.A(pi0217), .Y(new_n9353_));
  AND2X1   g06917(.A(new_n8945_), .B(new_n6621_), .Y(new_n9354_));
  NOR2X1   g06918(.A(new_n8981_), .B(new_n8948_), .Y(new_n9355_));
  OAI21X1  g06919(.A0(new_n9288_), .A1(new_n6364_), .B0(new_n9355_), .Y(new_n9356_));
  AOI21X1  g06920(.A0(new_n9307_), .A1(new_n6426_), .B0(new_n8948_), .Y(new_n9357_));
  OAI21X1  g06921(.A0(new_n9308_), .A1(new_n6364_), .B0(new_n9357_), .Y(new_n9358_));
  MX2X1    g06922(.A(new_n9358_), .B(new_n9356_), .S0(new_n6053_), .Y(new_n9359_));
  INVX1    g06923(.A(new_n9359_), .Y(new_n9360_));
  MX2X1    g06924(.A(new_n9360_), .B(new_n9354_), .S0(new_n9271_), .Y(new_n9361_));
  MX2X1    g06925(.A(new_n9360_), .B(new_n9354_), .S0(new_n6173_), .Y(new_n9362_));
  MX2X1    g06926(.A(new_n9362_), .B(new_n9361_), .S0(pi0333), .Y(new_n9363_));
  NOR2X1   g06927(.A(new_n9363_), .B(new_n6219_), .Y(new_n9364_));
  XOR2X1   g06928(.A(new_n6362_), .B(pi0392), .Y(new_n9365_));
  MX2X1    g06929(.A(new_n9362_), .B(new_n9361_), .S0(new_n6162_), .Y(new_n9366_));
  NOR2X1   g06930(.A(new_n9366_), .B(pi0391), .Y(new_n9367_));
  NOR3X1   g06931(.A(new_n9367_), .B(new_n9365_), .C(new_n9364_), .Y(new_n9368_));
  NOR2X1   g06932(.A(new_n9366_), .B(new_n6219_), .Y(new_n9369_));
  OAI21X1  g06933(.A0(new_n9363_), .A1(pi0391), .B0(new_n9365_), .Y(new_n9370_));
  OAI21X1  g06934(.A0(new_n9370_), .A1(new_n9369_), .B0(pi0591), .Y(new_n9371_));
  AOI22X1  g06935(.A0(new_n6653_), .A1(new_n6646_), .B0(new_n6604_), .B1(new_n6009_), .Y(new_n9372_));
  OAI21X1  g06936(.A0(new_n6645_), .A1(new_n6605_), .B0(new_n6025_), .Y(new_n9373_));
  NAND2X1  g06937(.A(new_n9373_), .B(new_n6666_), .Y(new_n9374_));
  OAI21X1  g06938(.A0(new_n9374_), .A1(new_n9372_), .B0(new_n8945_), .Y(new_n9375_));
  AOI21X1  g06939(.A0(new_n9375_), .A1(new_n6069_), .B0(pi0590), .Y(new_n9376_));
  OAI21X1  g06940(.A0(new_n9371_), .A1(new_n9368_), .B0(new_n9376_), .Y(new_n9377_));
  NOR3X1   g06941(.A(new_n9026_), .B(new_n6627_), .C(new_n6624_), .Y(new_n9378_));
  AOI21X1  g06942(.A0(new_n9378_), .A1(new_n6057_), .B0(new_n9354_), .Y(new_n9379_));
  AOI21X1  g06943(.A0(new_n9378_), .A1(new_n6052_), .B0(new_n9354_), .Y(new_n9380_));
  MX2X1    g06944(.A(new_n9380_), .B(new_n9379_), .S0(pi0461), .Y(new_n9381_));
  MX2X1    g06945(.A(new_n9380_), .B(new_n9379_), .S0(new_n5866_), .Y(new_n9382_));
  MX2X1    g06946(.A(new_n9382_), .B(new_n9381_), .S0(pi0357), .Y(new_n9383_));
  MX2X1    g06947(.A(new_n9382_), .B(new_n9381_), .S0(new_n5865_), .Y(new_n9384_));
  MX2X1    g06948(.A(new_n9384_), .B(new_n9383_), .S0(pi0356), .Y(new_n9385_));
  INVX1    g06949(.A(new_n9385_), .Y(new_n9386_));
  MX2X1    g06950(.A(new_n9384_), .B(new_n9383_), .S0(new_n5864_), .Y(new_n9387_));
  AOI21X1  g06951(.A0(new_n9387_), .A1(new_n9057_), .B0(new_n9062_), .Y(new_n9388_));
  OAI21X1  g06952(.A0(new_n9386_), .A1(new_n9057_), .B0(new_n9388_), .Y(new_n9389_));
  NAND2X1  g06953(.A(new_n9387_), .B(pi0354), .Y(new_n9390_));
  AOI21X1  g06954(.A0(new_n9385_), .A1(new_n9057_), .B0(new_n5862_), .Y(new_n9391_));
  AOI21X1  g06955(.A0(new_n9391_), .A1(new_n9390_), .B0(pi0591), .Y(new_n9392_));
  NAND2X1  g06956(.A(new_n9392_), .B(new_n9389_), .Y(new_n9393_));
  AOI21X1  g06957(.A0(new_n9393_), .A1(new_n9027_), .B0(pi0588), .Y(new_n9394_));
  AND2X1   g06958(.A(new_n6518_), .B(pi0592), .Y(new_n9395_));
  OAI21X1  g06959(.A0(new_n6690_), .A1(new_n6518_), .B0(new_n6604_), .Y(new_n9396_));
  OAI21X1  g06960(.A0(new_n9396_), .A1(new_n9395_), .B0(new_n8945_), .Y(new_n9397_));
  INVX1    g06961(.A(new_n9397_), .Y(new_n9398_));
  MX2X1    g06962(.A(new_n9398_), .B(new_n9354_), .S0(new_n6497_), .Y(new_n9399_));
  MX2X1    g06963(.A(new_n9398_), .B(new_n9354_), .S0(pi0428), .Y(new_n9400_));
  MX2X1    g06964(.A(new_n9400_), .B(new_n9399_), .S0(new_n6496_), .Y(new_n9401_));
  MX2X1    g06965(.A(new_n9400_), .B(new_n9399_), .S0(pi0427), .Y(new_n9402_));
  MX2X1    g06966(.A(new_n9402_), .B(new_n9401_), .S0(new_n6550_), .Y(new_n9403_));
  MX2X1    g06967(.A(new_n9402_), .B(new_n9401_), .S0(pi0430), .Y(new_n9404_));
  MX2X1    g06968(.A(new_n9404_), .B(new_n9403_), .S0(new_n6553_), .Y(new_n9405_));
  MX2X1    g06969(.A(new_n9404_), .B(new_n9403_), .S0(pi0426), .Y(new_n9406_));
  MX2X1    g06970(.A(new_n9406_), .B(new_n9405_), .S0(new_n6557_), .Y(new_n9407_));
  OR2X1    g06971(.A(new_n9406_), .B(pi0445), .Y(new_n9408_));
  OAI21X1  g06972(.A0(new_n9405_), .A1(new_n6557_), .B0(new_n9408_), .Y(new_n9409_));
  AOI21X1  g06973(.A0(new_n9409_), .A1(new_n6491_), .B0(new_n6591_), .Y(new_n9410_));
  OAI21X1  g06974(.A0(new_n9407_), .A1(new_n6491_), .B0(new_n9410_), .Y(new_n9411_));
  OR2X1    g06975(.A(new_n9407_), .B(pi0448), .Y(new_n9412_));
  AOI21X1  g06976(.A0(new_n9409_), .A1(pi0448), .B0(new_n6494_), .Y(new_n9413_));
  AOI21X1  g06977(.A0(new_n9413_), .A1(new_n9412_), .B0(new_n6053_), .Y(new_n9414_));
  OAI21X1  g06978(.A0(new_n9398_), .A1(pi1199), .B0(new_n6561_), .Y(new_n9415_));
  AOI21X1  g06979(.A0(new_n9414_), .A1(new_n9411_), .B0(new_n9415_), .Y(new_n9416_));
  OAI21X1  g06980(.A0(new_n9416_), .A1(new_n8947_), .B0(new_n6073_), .Y(new_n9417_));
  AOI21X1  g06981(.A0(new_n9394_), .A1(new_n9377_), .B0(new_n9417_), .Y(new_n9418_));
  AOI21X1  g06982(.A0(new_n5102_), .A1(new_n2436_), .B0(pi0080), .Y(new_n9419_));
  OAI21X1  g06983(.A0(new_n9026_), .A1(new_n6073_), .B0(new_n9419_), .Y(new_n9420_));
  OAI21X1  g06984(.A0(new_n9420_), .A1(new_n9418_), .B0(new_n9353_), .Y(new_n9421_));
  AOI21X1  g06985(.A0(new_n9352_), .A1(new_n9150_), .B0(new_n9421_), .Y(new_n9422_));
  INVX1    g06986(.A(pi0080), .Y(new_n9423_));
  AOI21X1  g06987(.A0(new_n9026_), .A1(new_n9423_), .B0(new_n9353_), .Y(new_n9424_));
  NOR3X1   g06988(.A(new_n9424_), .B(new_n9422_), .C(new_n8943_), .Y(po0238));
  NOR4X1   g06989(.A(new_n8371_), .B(po1038), .C(new_n3105_), .D(new_n2458_), .Y(new_n9426_));
  INVX1    g06990(.A(new_n9426_), .Y(new_n9427_));
  OR3X1    g06991(.A(new_n2470_), .B(pi0314), .C(new_n2579_), .Y(new_n9428_));
  INVX1    g06992(.A(pi0068), .Y(new_n9429_));
  OR4X1    g06993(.A(new_n8186_), .B(new_n2465_), .C(pi0081), .D(new_n9429_), .Y(new_n9430_));
  OR4X1    g06994(.A(new_n9430_), .B(new_n6750_), .C(new_n2633_), .D(pi0064), .Y(new_n9431_));
  AOI21X1  g06995(.A0(new_n9431_), .A1(new_n9428_), .B0(new_n9427_), .Y(po0239));
  AND2X1   g06996(.A(pi0314), .B(pi0069), .Y(new_n9433_));
  NOR4X1   g06997(.A(new_n2467_), .B(new_n2461_), .C(pi0073), .D(new_n6907_), .Y(new_n9434_));
  AOI21X1  g06998(.A0(new_n9433_), .A1(new_n2592_), .B0(new_n9434_), .Y(new_n9435_));
  NOR4X1   g06999(.A(new_n9435_), .B(new_n8245_), .C(new_n8440_), .D(new_n2460_), .Y(po0240));
  NOR3X1   g07000(.A(new_n8245_), .B(new_n2476_), .C(new_n2474_), .Y(new_n9437_));
  NOR4X1   g07001(.A(new_n6905_), .B(new_n2604_), .C(new_n2465_), .D(new_n2603_), .Y(new_n9438_));
  OAI21X1  g07002(.A0(new_n9438_), .A1(pi0083), .B0(new_n9437_), .Y(new_n9439_));
  OAI21X1  g07003(.A0(new_n9439_), .A1(new_n2597_), .B0(new_n5117_), .Y(new_n9440_));
  INVX1    g07004(.A(new_n7609_), .Y(new_n9441_));
  NAND4X1  g07005(.A(new_n9438_), .B(new_n9437_), .C(new_n2595_), .D(new_n2594_), .Y(new_n9442_));
  AOI21X1  g07006(.A0(new_n9442_), .A1(pi0314), .B0(new_n9441_), .Y(new_n9443_));
  AND2X1   g07007(.A(new_n9443_), .B(new_n9440_), .Y(po0241));
  NOR2X1   g07008(.A(new_n8055_), .B(pi0299), .Y(new_n9445_));
  AND2X1   g07009(.A(pi0299), .B(pi0211), .Y(new_n9446_));
  AND2X1   g07010(.A(pi0299), .B(pi0219), .Y(new_n9447_));
  NOR3X1   g07011(.A(new_n9447_), .B(new_n9446_), .C(new_n9445_), .Y(new_n9448_));
  INVX1    g07012(.A(new_n9448_), .Y(new_n9449_));
  NOR4X1   g07013(.A(new_n9449_), .B(new_n8425_), .C(po1038), .D(new_n3105_), .Y(po0242));
  NAND2X1  g07014(.A(new_n5131_), .B(pi0067), .Y(new_n9451_));
  OR3X1    g07015(.A(new_n8245_), .B(new_n2460_), .C(pi0069), .Y(new_n9452_));
  OR2X1    g07016(.A(new_n8246_), .B(pi0314), .Y(new_n9453_));
  OAI22X1  g07017(.A0(new_n9453_), .A1(new_n8465_), .B0(new_n9452_), .B1(new_n9451_), .Y(new_n9454_));
  AND2X1   g07018(.A(new_n9454_), .B(new_n8244_), .Y(po0243));
  AND3X1   g07019(.A(new_n5947_), .B(new_n5950_), .C(pi1091), .Y(new_n9456_));
  AOI22X1  g07020(.A0(new_n8437_), .A1(new_n9456_), .B0(new_n8435_), .B1(new_n5948_), .Y(new_n9457_));
  NOR2X1   g07021(.A(new_n9457_), .B(new_n8170_), .Y(po0244));
  OR4X1    g07022(.A(new_n8207_), .B(new_n8243_), .C(new_n2476_), .D(new_n5117_), .Y(new_n9459_));
  NOR4X1   g07023(.A(new_n9459_), .B(new_n8245_), .C(new_n2647_), .D(new_n2474_), .Y(po0245));
  AND3X1   g07024(.A(new_n8198_), .B(new_n8196_), .C(new_n5927_), .Y(new_n9461_));
  INVX1    g07025(.A(new_n7555_), .Y(new_n9462_));
  NOR4X1   g07026(.A(pi0110), .B(pi0091), .C(pi0058), .D(pi0047), .Y(new_n9463_));
  NOR4X1   g07027(.A(new_n8952_), .B(new_n8197_), .C(new_n5892_), .D(pi0094), .Y(new_n9464_));
  AND3X1   g07028(.A(new_n9464_), .B(new_n9463_), .C(new_n8208_), .Y(new_n9465_));
  OR2X1    g07029(.A(new_n9465_), .B(new_n5032_), .Y(new_n9466_));
  AND3X1   g07030(.A(new_n9466_), .B(new_n9462_), .C(new_n3104_), .Y(new_n9467_));
  OAI21X1  g07031(.A0(new_n9461_), .A1(pi1093), .B0(new_n9467_), .Y(new_n9468_));
  NAND4X1  g07032(.A(new_n3103_), .B(new_n3047_), .C(new_n2984_), .D(new_n5032_), .Y(new_n9469_));
  OR3X1    g07033(.A(new_n9469_), .B(new_n5928_), .C(new_n7763_), .Y(new_n9470_));
  NOR4X1   g07034(.A(new_n9470_), .B(new_n8480_), .C(new_n2567_), .D(pi0098), .Y(new_n9471_));
  OAI21X1  g07035(.A0(new_n9471_), .A1(new_n6072_), .B0(new_n6489_), .Y(new_n9472_));
  AOI21X1  g07036(.A0(new_n9468_), .A1(new_n6072_), .B0(new_n9472_), .Y(po0246));
  NOR4X1   g07037(.A(new_n8172_), .B(new_n2458_), .C(pi0081), .D(pi0064), .Y(new_n9474_));
  NAND2X1  g07038(.A(new_n9474_), .B(new_n7617_), .Y(new_n9475_));
  NOR3X1   g07039(.A(new_n9475_), .B(new_n5898_), .C(new_n2705_), .Y(new_n9476_));
  INVX1    g07040(.A(new_n7607_), .Y(new_n9477_));
  NOR4X1   g07041(.A(new_n9477_), .B(new_n3279_), .C(new_n2985_), .D(pi0092), .Y(new_n9478_));
  OAI21X1  g07042(.A0(new_n9476_), .A1(pi0070), .B0(new_n9478_), .Y(new_n9479_));
  AOI21X1  g07043(.A0(new_n6772_), .A1(pi0070), .B0(new_n9479_), .Y(po0247));
  AOI21X1  g07044(.A0(new_n7224_), .A1(new_n8493_), .B0(pi0090), .Y(new_n9481_));
  NOR4X1   g07045(.A(new_n9481_), .B(new_n8391_), .C(new_n5886_), .D(new_n2683_), .Y(po0248));
  INVX1    g07046(.A(new_n7625_), .Y(new_n9483_));
  INVX1    g07047(.A(new_n7732_), .Y(new_n9484_));
  OAI21X1  g07048(.A0(new_n9484_), .A1(pi0058), .B0(new_n7604_), .Y(new_n9485_));
  AND2X1   g07049(.A(new_n7606_), .B(new_n2757_), .Y(new_n9486_));
  OR4X1    g07050(.A(new_n8233_), .B(new_n2757_), .C(new_n2728_), .D(new_n5777_), .Y(new_n9487_));
  OAI21X1  g07051(.A0(new_n9487_), .A1(new_n9484_), .B0(new_n2939_), .Y(new_n9488_));
  AOI21X1  g07052(.A0(new_n9486_), .A1(new_n9485_), .B0(new_n9488_), .Y(new_n9489_));
  NOR3X1   g07053(.A(new_n9489_), .B(new_n9483_), .C(new_n5954_), .Y(po0249));
  NAND4X1  g07054(.A(new_n3111_), .B(new_n3077_), .C(pi1050), .D(new_n5117_), .Y(new_n9491_));
  OR4X1    g07055(.A(new_n9491_), .B(new_n2985_), .C(new_n2536_), .D(new_n3079_), .Y(new_n9492_));
  NOR4X1   g07056(.A(new_n2933_), .B(new_n2437_), .C(new_n2438_), .D(pi0215), .Y(new_n9493_));
  AND3X1   g07057(.A(new_n4769_), .B(pi0224), .C(pi0222), .Y(new_n9494_));
  AOI22X1  g07058(.A0(new_n9494_), .A1(new_n9456_), .B0(new_n9493_), .B1(new_n5948_), .Y(new_n9495_));
  OR3X1    g07059(.A(new_n9495_), .B(new_n8260_), .C(new_n3112_), .Y(new_n9496_));
  AOI21X1  g07060(.A0(new_n9496_), .A1(new_n9492_), .B0(new_n9477_), .Y(po0250));
  OR3X1    g07061(.A(new_n2985_), .B(new_n2536_), .C(pi1050), .Y(new_n9498_));
  AND2X1   g07062(.A(new_n7607_), .B(new_n3208_), .Y(new_n9499_));
  AND3X1   g07063(.A(new_n8232_), .B(new_n5164_), .C(pi0093), .Y(new_n9500_));
  OAI21X1  g07064(.A0(new_n9500_), .A1(pi0092), .B0(new_n9499_), .Y(new_n9501_));
  AOI21X1  g07065(.A0(new_n9498_), .A1(pi0092), .B0(new_n9501_), .Y(po0251));
  NOR4X1   g07066(.A(new_n8222_), .B(new_n6773_), .C(new_n2484_), .D(pi0841), .Y(new_n9503_));
  AOI21X1  g07067(.A0(new_n9503_), .A1(new_n2703_), .B0(new_n5032_), .Y(new_n9504_));
  AOI21X1  g07068(.A0(new_n8221_), .A1(new_n7663_), .B0(new_n2570_), .Y(new_n9505_));
  NAND3X1  g07069(.A(new_n7606_), .B(new_n2497_), .C(pi0252), .Y(new_n9506_));
  OAI22X1  g07070(.A0(new_n9506_), .A1(new_n9505_), .B0(new_n9504_), .B1(new_n2762_), .Y(new_n9507_));
  AND2X1   g07071(.A(new_n9507_), .B(new_n6741_), .Y(new_n9508_));
  OAI22X1  g07072(.A0(new_n9508_), .A1(new_n9503_), .B0(new_n9507_), .B1(new_n3035_), .Y(new_n9509_));
  OAI21X1  g07073(.A0(new_n9503_), .A1(new_n6728_), .B0(new_n7608_), .Y(new_n9510_));
  AOI21X1  g07074(.A0(new_n9509_), .A1(new_n6728_), .B0(new_n9510_), .Y(po0252));
  OAI21X1  g07075(.A0(new_n5235_), .A1(new_n5229_), .B0(new_n5950_), .Y(new_n9512_));
  OR3X1    g07076(.A(new_n9512_), .B(new_n8452_), .C(new_n3261_), .Y(new_n9513_));
  INVX1    g07077(.A(new_n8456_), .Y(new_n9514_));
  NOR3X1   g07078(.A(new_n9514_), .B(new_n8454_), .C(new_n5236_), .Y(new_n9515_));
  NOR2X1   g07079(.A(new_n9515_), .B(new_n2939_), .Y(new_n9516_));
  AND3X1   g07080(.A(new_n2456_), .B(pi0095), .C(new_n2455_), .Y(new_n9517_));
  AND3X1   g07081(.A(new_n9517_), .B(new_n2531_), .C(pi0024), .Y(new_n9518_));
  NAND4X1  g07082(.A(new_n7606_), .B(new_n2483_), .C(new_n2705_), .D(new_n2444_), .Y(new_n9519_));
  OAI21X1  g07083(.A0(new_n9519_), .A1(new_n9475_), .B0(new_n2939_), .Y(new_n9520_));
  OAI21X1  g07084(.A0(new_n9520_), .A1(new_n9518_), .B0(new_n7628_), .Y(new_n9521_));
  AOI21X1  g07085(.A0(new_n9516_), .A1(new_n9513_), .B0(new_n9521_), .Y(po0253));
  NAND4X1  g07086(.A(new_n9517_), .B(new_n2479_), .C(new_n2477_), .D(new_n5777_), .Y(new_n9523_));
  AND2X1   g07087(.A(new_n6741_), .B(pi0479), .Y(new_n9524_));
  INVX1    g07088(.A(new_n2706_), .Y(new_n9525_));
  NAND4X1  g07089(.A(new_n2695_), .B(pi0096), .C(new_n2535_), .D(new_n2508_), .Y(new_n9526_));
  NOR4X1   g07090(.A(new_n9526_), .B(new_n9524_), .C(new_n9525_), .D(new_n2691_), .Y(new_n9527_));
  AOI21X1  g07091(.A0(new_n9524_), .A1(new_n2877_), .B0(new_n9527_), .Y(new_n9528_));
  OAI21X1  g07092(.A0(new_n9528_), .A1(pi0095), .B0(new_n9523_), .Y(new_n9529_));
  AND2X1   g07093(.A(new_n9529_), .B(new_n7608_), .Y(po0254));
  NAND2X1  g07094(.A(pi0593), .B(pi0039), .Y(new_n9531_));
  OR3X1    g07095(.A(new_n9531_), .B(new_n8457_), .C(new_n5236_), .Y(new_n9532_));
  AOI21X1  g07096(.A0(new_n9524_), .A1(new_n5009_), .B0(po0740), .Y(new_n9533_));
  OR4X1    g07097(.A(new_n9533_), .B(new_n8499_), .C(new_n8449_), .D(pi0096), .Y(new_n9534_));
  AOI21X1  g07098(.A0(new_n9534_), .A1(new_n9532_), .B0(new_n7629_), .Y(po0255));
  MX2X1    g07099(.A(new_n8494_), .B(new_n2986_), .S0(pi0092), .Y(new_n9536_));
  NAND4X1  g07100(.A(new_n7607_), .B(new_n3208_), .C(pi1050), .D(pi0314), .Y(new_n9537_));
  NOR2X1   g07101(.A(new_n9537_), .B(new_n9536_), .Y(po0256));
  AND2X1   g07102(.A(pi0099), .B(new_n2530_), .Y(new_n9539_));
  INVX1    g07103(.A(new_n9539_), .Y(new_n9540_));
  OAI21X1  g07104(.A0(new_n5920_), .A1(new_n2793_), .B0(new_n9540_), .Y(new_n9541_));
  AOI21X1  g07105(.A0(new_n9539_), .A1(new_n2704_), .B0(new_n7692_), .Y(new_n9542_));
  NOR2X1   g07106(.A(new_n9540_), .B(new_n7710_), .Y(new_n9543_));
  AOI21X1  g07107(.A0(new_n8125_), .A1(new_n5079_), .B0(new_n9543_), .Y(new_n9544_));
  OAI21X1  g07108(.A0(new_n9544_), .A1(new_n7805_), .B0(new_n9542_), .Y(new_n9545_));
  AOI21X1  g07109(.A0(new_n9545_), .A1(new_n9541_), .B0(pi0039), .Y(new_n9546_));
  NOR4X1   g07110(.A(new_n8677_), .B(new_n4611_), .C(new_n3193_), .D(pi0072), .Y(new_n9547_));
  AND3X1   g07111(.A(new_n2933_), .B(pi0174), .C(new_n2530_), .Y(new_n9548_));
  AOI22X1  g07112(.A0(new_n9548_), .A1(new_n7715_), .B0(new_n9547_), .B1(pi0299), .Y(new_n9549_));
  OAI21X1  g07113(.A0(new_n9549_), .A1(new_n5215_), .B0(pi0039), .Y(new_n9550_));
  NAND2X1  g07114(.A(new_n9550_), .B(new_n3087_), .Y(new_n9551_));
  INVX1    g07115(.A(new_n9550_), .Y(new_n9552_));
  AOI21X1  g07116(.A0(new_n9540_), .A1(new_n2939_), .B0(new_n9552_), .Y(new_n9553_));
  AOI21X1  g07117(.A0(new_n9553_), .A1(new_n5778_), .B0(new_n3073_), .Y(new_n9554_));
  OAI21X1  g07118(.A0(new_n9551_), .A1(new_n9546_), .B0(new_n9554_), .Y(new_n9555_));
  AOI21X1  g07119(.A0(pi0072), .A1(pi0041), .B0(new_n7703_), .Y(new_n9556_));
  INVX1    g07120(.A(new_n9556_), .Y(new_n9557_));
  NOR2X1   g07121(.A(new_n9557_), .B(new_n7752_), .Y(new_n9558_));
  NOR2X1   g07122(.A(new_n9558_), .B(new_n8008_), .Y(new_n9559_));
  INVX1    g07123(.A(new_n7756_), .Y(new_n9560_));
  AOI21X1  g07124(.A0(new_n9556_), .A1(new_n9560_), .B0(new_n8007_), .Y(new_n9561_));
  OAI21X1  g07125(.A0(new_n9561_), .A1(new_n9559_), .B0(pi0228), .Y(new_n9562_));
  NOR2X1   g07126(.A(new_n7863_), .B(pi0228), .Y(new_n9563_));
  OAI21X1  g07127(.A0(new_n9557_), .A1(new_n7792_), .B0(new_n9563_), .Y(new_n9564_));
  AND2X1   g07128(.A(new_n9564_), .B(new_n2939_), .Y(new_n9565_));
  INVX1    g07129(.A(new_n7822_), .Y(new_n9566_));
  OR2X1    g07130(.A(new_n9549_), .B(new_n9566_), .Y(new_n9567_));
  AOI21X1  g07131(.A0(new_n8143_), .A1(pi0287), .B0(new_n9567_), .Y(new_n9568_));
  OR2X1    g07132(.A(new_n9568_), .B(new_n3252_), .Y(new_n9569_));
  AOI21X1  g07133(.A0(new_n9565_), .A1(new_n9562_), .B0(new_n9569_), .Y(new_n9570_));
  NOR2X1   g07134(.A(new_n9540_), .B(new_n7804_), .Y(new_n9571_));
  AOI21X1  g07135(.A0(new_n7699_), .A1(new_n7832_), .B0(new_n9571_), .Y(new_n9572_));
  OAI21X1  g07136(.A0(new_n9572_), .A1(new_n7805_), .B0(new_n9542_), .Y(new_n9573_));
  AOI21X1  g07137(.A0(new_n9573_), .A1(new_n9541_), .B0(pi0039), .Y(new_n9574_));
  OAI21X1  g07138(.A0(new_n9574_), .A1(new_n9552_), .B0(new_n5074_), .Y(new_n9575_));
  INVX1    g07139(.A(new_n9553_), .Y(new_n9576_));
  AOI21X1  g07140(.A0(new_n9576_), .A1(pi0038), .B0(pi0087), .Y(new_n9577_));
  NAND2X1  g07141(.A(new_n9577_), .B(new_n9575_), .Y(new_n9578_));
  NOR3X1   g07142(.A(new_n7698_), .B(new_n7833_), .C(new_n2793_), .Y(new_n9579_));
  AOI21X1  g07143(.A0(new_n7802_), .A1(pi0228), .B0(new_n9540_), .Y(new_n9580_));
  OR3X1    g07144(.A(new_n9580_), .B(new_n9579_), .C(new_n3378_), .Y(new_n9581_));
  AOI21X1  g07145(.A0(new_n9576_), .A1(new_n3378_), .B0(new_n3131_), .Y(new_n9582_));
  AOI21X1  g07146(.A0(new_n9582_), .A1(new_n9581_), .B0(pi0075), .Y(new_n9583_));
  OAI21X1  g07147(.A0(new_n9578_), .A1(new_n9570_), .B0(new_n9583_), .Y(new_n9584_));
  AOI21X1  g07148(.A0(new_n9584_), .A1(new_n9555_), .B0(new_n6295_), .Y(new_n9585_));
  OAI21X1  g07149(.A0(new_n9553_), .A1(new_n5880_), .B0(new_n6489_), .Y(new_n9586_));
  AOI21X1  g07150(.A0(new_n9547_), .A1(pi0232), .B0(new_n2939_), .Y(new_n9587_));
  OAI22X1  g07151(.A0(new_n9539_), .A1(pi0039), .B0(new_n5103_), .B1(pi0057), .Y(new_n9588_));
  OAI22X1  g07152(.A0(new_n9588_), .A1(new_n9587_), .B0(new_n9586_), .B1(new_n9585_), .Y(po0257));
  INVX1    g07153(.A(new_n6722_), .Y(new_n9590_));
  AOI21X1  g07154(.A0(new_n7557_), .A1(new_n6820_), .B0(new_n5083_), .Y(new_n9591_));
  NOR2X1   g07155(.A(new_n5082_), .B(pi0683), .Y(new_n9592_));
  OR2X1    g07156(.A(new_n5086_), .B(new_n9592_), .Y(new_n9593_));
  INVX1    g07157(.A(new_n7558_), .Y(new_n9594_));
  OR2X1    g07158(.A(new_n7557_), .B(new_n5083_), .Y(new_n9595_));
  AOI22X1  g07159(.A0(new_n9595_), .A1(new_n9594_), .B0(new_n9593_), .B1(new_n5072_), .Y(new_n9596_));
  OAI21X1  g07160(.A0(new_n9591_), .A1(new_n7554_), .B0(new_n9596_), .Y(new_n9597_));
  NOR4X1   g07161(.A(new_n7141_), .B(new_n3007_), .C(pi0075), .D(pi0038), .Y(new_n9598_));
  NOR4X1   g07162(.A(new_n6779_), .B(new_n6776_), .C(new_n6741_), .D(pi0024), .Y(new_n9599_));
  AOI21X1  g07163(.A0(new_n9598_), .A1(new_n9597_), .B0(new_n9599_), .Y(new_n9600_));
  NOR3X1   g07164(.A(new_n9600_), .B(new_n9590_), .C(new_n2986_), .Y(po0258));
  AND2X1   g07165(.A(pi0101), .B(new_n2530_), .Y(new_n9602_));
  INVX1    g07166(.A(new_n9602_), .Y(new_n9603_));
  OAI21X1  g07167(.A0(new_n5920_), .A1(new_n2793_), .B0(new_n9603_), .Y(new_n9604_));
  AOI21X1  g07168(.A0(new_n9602_), .A1(new_n2704_), .B0(new_n7692_), .Y(new_n9605_));
  NAND2X1  g07169(.A(new_n5081_), .B(new_n5079_), .Y(new_n9606_));
  NAND2X1  g07170(.A(new_n9606_), .B(new_n2703_), .Y(new_n9607_));
  AOI22X1  g07171(.A0(new_n7709_), .A1(new_n9602_), .B0(new_n7699_), .B1(new_n6239_), .Y(new_n9608_));
  OAI21X1  g07172(.A0(new_n9608_), .A1(new_n9607_), .B0(new_n9605_), .Y(new_n9609_));
  AOI21X1  g07173(.A0(new_n9609_), .A1(new_n9604_), .B0(pi0039), .Y(new_n9610_));
  NOR4X1   g07174(.A(new_n3192_), .B(pi0468), .C(pi0332), .D(new_n3193_), .Y(new_n9611_));
  AOI21X1  g07175(.A0(new_n9611_), .A1(new_n2530_), .B0(new_n2933_), .Y(new_n9612_));
  AND3X1   g07176(.A(new_n7714_), .B(pi0174), .C(new_n7344_), .Y(new_n9613_));
  AOI21X1  g07177(.A0(new_n9613_), .A1(new_n2530_), .B0(pi0299), .Y(new_n9614_));
  OR2X1    g07178(.A(new_n9614_), .B(new_n5215_), .Y(new_n9615_));
  OAI21X1  g07179(.A0(new_n9615_), .A1(new_n9612_), .B0(pi0039), .Y(new_n9616_));
  NAND2X1  g07180(.A(new_n9616_), .B(new_n3087_), .Y(new_n9617_));
  INVX1    g07181(.A(new_n9616_), .Y(new_n9618_));
  AOI21X1  g07182(.A0(new_n9603_), .A1(new_n2939_), .B0(new_n9618_), .Y(new_n9619_));
  AOI21X1  g07183(.A0(new_n9619_), .A1(new_n5778_), .B0(new_n3073_), .Y(new_n9620_));
  OAI21X1  g07184(.A0(new_n9617_), .A1(new_n9610_), .B0(new_n9620_), .Y(new_n9621_));
  NAND2X1  g07185(.A(new_n7741_), .B(new_n2703_), .Y(new_n9622_));
  AOI21X1  g07186(.A0(new_n7751_), .A1(pi0101), .B0(new_n9622_), .Y(new_n9623_));
  OR2X1    g07187(.A(new_n7759_), .B(new_n2703_), .Y(new_n9624_));
  AOI21X1  g07188(.A0(new_n7755_), .A1(pi0101), .B0(new_n9624_), .Y(new_n9625_));
  OAI21X1  g07189(.A0(new_n9625_), .A1(new_n9623_), .B0(pi0228), .Y(new_n9626_));
  NAND2X1  g07190(.A(new_n7791_), .B(pi0101), .Y(new_n9627_));
  NOR2X1   g07191(.A(new_n7787_), .B(pi0228), .Y(new_n9628_));
  AOI21X1  g07192(.A0(new_n9628_), .A1(new_n9627_), .B0(pi0039), .Y(new_n9629_));
  AOI21X1  g07193(.A0(new_n9611_), .A1(new_n8144_), .B0(new_n2933_), .Y(new_n9630_));
  AOI21X1  g07194(.A0(new_n9613_), .A1(new_n8144_), .B0(pi0299), .Y(new_n9631_));
  NOR3X1   g07195(.A(new_n9631_), .B(new_n9630_), .C(new_n9566_), .Y(new_n9632_));
  OR2X1    g07196(.A(new_n9632_), .B(new_n3252_), .Y(new_n9633_));
  AOI21X1  g07197(.A0(new_n9629_), .A1(new_n9626_), .B0(new_n9633_), .Y(new_n9634_));
  INVX1    g07198(.A(new_n9605_), .Y(new_n9635_));
  OAI21X1  g07199(.A0(new_n8148_), .A1(pi0044), .B0(new_n9602_), .Y(new_n9636_));
  AOI21X1  g07200(.A0(new_n9636_), .A1(new_n7700_), .B0(new_n9607_), .Y(new_n9637_));
  OAI21X1  g07201(.A0(new_n9637_), .A1(new_n9635_), .B0(new_n9604_), .Y(new_n9638_));
  AOI21X1  g07202(.A0(new_n9638_), .A1(new_n2939_), .B0(new_n9618_), .Y(new_n9639_));
  OR2X1    g07203(.A(new_n9619_), .B(new_n2979_), .Y(new_n9640_));
  AND2X1   g07204(.A(new_n9640_), .B(new_n3131_), .Y(new_n9641_));
  OAI21X1  g07205(.A0(new_n9639_), .A1(new_n5075_), .B0(new_n9641_), .Y(new_n9642_));
  NAND2X1  g07206(.A(new_n8157_), .B(new_n7743_), .Y(new_n9643_));
  OAI21X1  g07207(.A0(new_n8156_), .A1(new_n7801_), .B0(new_n9602_), .Y(new_n9644_));
  NAND3X1  g07208(.A(new_n9644_), .B(new_n9643_), .C(new_n2939_), .Y(new_n9645_));
  AND2X1   g07209(.A(new_n9616_), .B(pi0087), .Y(new_n9646_));
  AOI21X1  g07210(.A0(new_n9646_), .A1(new_n9645_), .B0(pi0075), .Y(new_n9647_));
  OAI21X1  g07211(.A0(new_n9642_), .A1(new_n9634_), .B0(new_n9647_), .Y(new_n9648_));
  AOI21X1  g07212(.A0(new_n9648_), .A1(new_n9621_), .B0(new_n6295_), .Y(new_n9649_));
  OAI21X1  g07213(.A0(new_n9619_), .A1(new_n5880_), .B0(new_n6489_), .Y(new_n9650_));
  NAND3X1  g07214(.A(new_n9611_), .B(pi0232), .C(new_n2530_), .Y(new_n9651_));
  AND2X1   g07215(.A(new_n9651_), .B(pi0039), .Y(new_n9652_));
  OAI22X1  g07216(.A0(new_n9602_), .A1(pi0039), .B0(new_n5103_), .B1(pi0057), .Y(new_n9653_));
  OAI22X1  g07217(.A0(new_n9653_), .A1(new_n9652_), .B0(new_n9650_), .B1(new_n9649_), .Y(po0259));
  NOR4X1   g07218(.A(new_n6746_), .B(new_n2468_), .C(pi0071), .D(new_n2650_), .Y(new_n9655_));
  AND2X1   g07219(.A(new_n9655_), .B(new_n9426_), .Y(po0260));
  NOR3X1   g07220(.A(new_n8245_), .B(new_n2647_), .C(new_n2474_), .Y(new_n9657_));
  OAI21X1  g07221(.A0(new_n9657_), .A1(pi0109), .B0(new_n5119_), .Y(new_n9658_));
  AND3X1   g07222(.A(new_n7609_), .B(new_n2515_), .C(new_n2494_), .Y(new_n9659_));
  AND3X1   g07223(.A(new_n2555_), .B(new_n2548_), .C(pi0109), .Y(new_n9660_));
  OAI21X1  g07224(.A0(new_n9660_), .A1(new_n5117_), .B0(new_n9659_), .Y(new_n9661_));
  AOI21X1  g07225(.A0(new_n9658_), .A1(new_n5117_), .B0(new_n9661_), .Y(po0261));
  NOR2X1   g07226(.A(new_n7555_), .B(new_n5928_), .Y(new_n9663_));
  OAI21X1  g07227(.A0(new_n6728_), .A1(new_n6073_), .B0(new_n9663_), .Y(new_n9664_));
  NAND3X1  g07228(.A(new_n9664_), .B(new_n7776_), .C(new_n7606_), .Y(new_n9665_));
  AND3X1   g07229(.A(new_n7606_), .B(new_n5927_), .C(new_n2550_), .Y(new_n9666_));
  OAI21X1  g07230(.A0(new_n9464_), .A1(pi0110), .B0(new_n9666_), .Y(new_n9667_));
  OR3X1    g07231(.A(new_n9667_), .B(new_n2549_), .C(new_n4999_), .Y(new_n9668_));
  NOR2X1   g07232(.A(new_n7555_), .B(new_n5920_), .Y(new_n9669_));
  OAI21X1  g07233(.A0(new_n9465_), .A1(new_n5082_), .B0(new_n9669_), .Y(new_n9670_));
  AOI21X1  g07234(.A0(new_n9668_), .A1(new_n5082_), .B0(new_n9670_), .Y(new_n9671_));
  INVX1    g07235(.A(new_n5920_), .Y(new_n9672_));
  NOR3X1   g07236(.A(new_n9668_), .B(new_n7555_), .C(new_n9672_), .Y(new_n9673_));
  OAI21X1  g07237(.A0(new_n9673_), .A1(new_n9671_), .B0(new_n6073_), .Y(new_n9674_));
  AOI21X1  g07238(.A0(new_n9674_), .A1(new_n9665_), .B0(new_n8207_), .Y(po0262));
  NOR3X1   g07239(.A(new_n8362_), .B(new_n8357_), .C(new_n5777_), .Y(new_n9676_));
  AOI21X1  g07240(.A0(new_n8362_), .A1(new_n2485_), .B0(new_n2493_), .Y(new_n9677_));
  AND3X1   g07241(.A(new_n9677_), .B(new_n2497_), .C(new_n5777_), .Y(new_n9678_));
  OAI21X1  g07242(.A0(new_n9678_), .A1(new_n9676_), .B0(pi0841), .Y(new_n9679_));
  NAND3X1  g07243(.A(new_n8350_), .B(new_n2705_), .C(new_n5777_), .Y(new_n9680_));
  AOI21X1  g07244(.A0(new_n9680_), .A1(new_n9679_), .B0(new_n9441_), .Y(po0264));
  NOR3X1   g07245(.A(new_n8410_), .B(new_n9441_), .C(pi0999), .Y(po0265));
  AND2X1   g07246(.A(new_n2562_), .B(pi0108), .Y(new_n9683_));
  AOI21X1  g07247(.A0(new_n5895_), .A1(new_n7656_), .B0(pi0108), .Y(new_n9684_));
  OR4X1    g07248(.A(new_n9684_), .B(new_n9683_), .C(new_n2495_), .D(new_n2475_), .Y(new_n9685_));
  OAI21X1  g07249(.A0(new_n5896_), .A1(new_n2498_), .B0(pi0314), .Y(new_n9686_));
  NAND4X1  g07250(.A(new_n9686_), .B(new_n7668_), .C(new_n5897_), .D(new_n2535_), .Y(new_n9687_));
  AOI21X1  g07251(.A0(new_n9685_), .A1(new_n5117_), .B0(new_n9687_), .Y(new_n9688_));
  OR3X1    g07252(.A(new_n7668_), .B(new_n5898_), .C(pi0070), .Y(new_n9689_));
  OAI21X1  g07253(.A0(new_n9689_), .A1(new_n9685_), .B0(new_n2534_), .Y(new_n9690_));
  NOR4X1   g07254(.A(new_n3132_), .B(new_n5881_), .C(new_n2847_), .D(pi0096), .Y(new_n9691_));
  OAI21X1  g07255(.A0(new_n9690_), .A1(new_n9688_), .B0(new_n9691_), .Y(new_n9692_));
  NAND3X1  g07256(.A(new_n6722_), .B(new_n5090_), .C(new_n3073_), .Y(new_n9693_));
  AOI21X1  g07257(.A0(new_n9692_), .A1(new_n3131_), .B0(new_n9693_), .Y(po0266));
  NOR4X1   g07258(.A(new_n8172_), .B(new_n2559_), .C(new_n2576_), .D(pi0050), .Y(new_n9695_));
  AND3X1   g07259(.A(new_n9695_), .B(new_n7609_), .C(pi0314), .Y(po0267));
  NAND4X1  g07260(.A(new_n9463_), .B(pi0111), .C(new_n2546_), .D(new_n2629_), .Y(new_n9697_));
  NOR3X1   g07261(.A(new_n9697_), .B(new_n8246_), .C(new_n2474_), .Y(new_n9698_));
  AND2X1   g07262(.A(new_n9698_), .B(new_n2631_), .Y(new_n9699_));
  NOR4X1   g07263(.A(new_n7555_), .B(new_n5928_), .C(new_n5920_), .D(new_n5082_), .Y(new_n9700_));
  AOI22X1  g07264(.A0(new_n9700_), .A1(new_n7776_), .B0(new_n9699_), .B1(pi0314), .Y(new_n9701_));
  NOR2X1   g07265(.A(new_n9701_), .B(new_n9441_), .Y(po0268));
  AND3X1   g07266(.A(new_n9698_), .B(new_n2631_), .C(new_n5117_), .Y(new_n9703_));
  INVX1    g07267(.A(new_n9703_), .Y(new_n9704_));
  OAI22X1  g07268(.A0(new_n9704_), .A1(new_n8479_), .B0(new_n7707_), .B1(new_n2530_), .Y(new_n9705_));
  AND3X1   g07269(.A(new_n9705_), .B(new_n7608_), .C(new_n5168_), .Y(po0269));
  NAND2X1  g07270(.A(new_n8621_), .B(pi0124), .Y(po0270));
  AND3X1   g07271(.A(pi0113), .B(new_n2530_), .C(new_n2939_), .Y(new_n9708_));
  INVX1    g07272(.A(new_n7753_), .Y(new_n9709_));
  AOI21X1  g07273(.A0(new_n9560_), .A1(new_n2704_), .B0(pi0099), .Y(new_n9710_));
  OAI21X1  g07274(.A0(new_n7832_), .A1(new_n2530_), .B0(pi0113), .Y(new_n9711_));
  AOI21X1  g07275(.A0(new_n9710_), .A1(new_n9709_), .B0(new_n9711_), .Y(new_n9712_));
  OAI21X1  g07276(.A0(new_n8009_), .A1(pi0113), .B0(pi0228), .Y(new_n9713_));
  NAND2X1  g07277(.A(new_n7857_), .B(pi0113), .Y(new_n9714_));
  AOI21X1  g07278(.A0(new_n7863_), .A1(new_n7861_), .B0(pi0228), .Y(new_n9715_));
  AOI21X1  g07279(.A0(new_n9715_), .A1(new_n9714_), .B0(pi0039), .Y(new_n9716_));
  OAI21X1  g07280(.A0(new_n9713_), .A1(new_n9712_), .B0(new_n9716_), .Y(new_n9717_));
  AND2X1   g07281(.A(pi0113), .B(new_n2530_), .Y(new_n9718_));
  NOR3X1   g07282(.A(new_n5920_), .B(new_n2704_), .C(new_n2793_), .Y(new_n9719_));
  INVX1    g07283(.A(new_n9719_), .Y(new_n9720_));
  NOR2X1   g07284(.A(new_n7801_), .B(new_n7895_), .Y(new_n9721_));
  AOI21X1  g07285(.A0(new_n9721_), .A1(new_n7696_), .B0(new_n5081_), .Y(new_n9722_));
  OAI21X1  g07286(.A0(new_n9722_), .A1(new_n9720_), .B0(new_n9718_), .Y(new_n9723_));
  NOR4X1   g07287(.A(new_n5920_), .B(new_n5081_), .C(new_n2704_), .D(new_n2793_), .Y(new_n9724_));
  INVX1    g07288(.A(new_n9724_), .Y(new_n9725_));
  NOR4X1   g07289(.A(new_n9725_), .B(new_n7700_), .C(new_n7833_), .D(pi0113), .Y(new_n9726_));
  INVX1    g07290(.A(new_n9726_), .Y(new_n9727_));
  AOI21X1  g07291(.A0(new_n9727_), .A1(new_n9723_), .B0(pi0039), .Y(new_n9728_));
  OAI22X1  g07292(.A0(new_n9728_), .A1(new_n5075_), .B0(new_n9708_), .B1(new_n2979_), .Y(new_n9729_));
  AOI21X1  g07293(.A0(new_n9717_), .A1(new_n3251_), .B0(new_n9729_), .Y(new_n9730_));
  AOI22X1  g07294(.A0(new_n9718_), .A1(new_n7914_), .B0(new_n9579_), .B1(new_n7861_), .Y(new_n9731_));
  AOI21X1  g07295(.A0(new_n9708_), .A1(new_n3252_), .B0(new_n3131_), .Y(new_n9732_));
  OAI21X1  g07296(.A0(new_n9731_), .A1(new_n3378_), .B0(new_n9732_), .Y(new_n9733_));
  OAI21X1  g07297(.A0(new_n9730_), .A1(pi0087), .B0(new_n9733_), .Y(new_n9734_));
  NOR2X1   g07298(.A(new_n7709_), .B(new_n7895_), .Y(new_n9735_));
  OAI21X1  g07299(.A0(new_n9735_), .A1(new_n5081_), .B0(new_n9719_), .Y(new_n9736_));
  AOI22X1  g07300(.A0(new_n9736_), .A1(new_n9718_), .B0(new_n9726_), .B1(new_n6239_), .Y(new_n9737_));
  OR2X1    g07301(.A(new_n9737_), .B(new_n3074_), .Y(new_n9738_));
  AOI21X1  g07302(.A0(new_n9708_), .A1(new_n5778_), .B0(new_n3073_), .Y(new_n9739_));
  AOI22X1  g07303(.A0(new_n9739_), .A1(new_n9738_), .B0(new_n9734_), .B1(new_n3073_), .Y(new_n9740_));
  MX2X1    g07304(.A(new_n9740_), .B(new_n9708_), .S0(new_n9590_), .Y(po0271));
  AND3X1   g07305(.A(pi0114), .B(new_n2530_), .C(new_n2939_), .Y(new_n9742_));
  NAND2X1  g07306(.A(new_n7925_), .B(new_n2530_), .Y(new_n9743_));
  OAI21X1  g07307(.A0(new_n9743_), .A1(new_n7830_), .B0(new_n8278_), .Y(new_n9744_));
  AND2X1   g07308(.A(pi0114), .B(new_n2530_), .Y(new_n9745_));
  INVX1    g07309(.A(new_n9745_), .Y(new_n9746_));
  AOI21X1  g07310(.A0(new_n9746_), .A1(new_n8279_), .B0(new_n3074_), .Y(new_n9747_));
  OAI21X1  g07311(.A0(new_n9744_), .A1(new_n7923_), .B0(new_n9747_), .Y(new_n9748_));
  AOI21X1  g07312(.A0(new_n9742_), .A1(new_n5778_), .B0(new_n3073_), .Y(new_n9749_));
  MX2X1    g07313(.A(new_n8012_), .B(new_n8002_), .S0(pi0114), .Y(new_n9750_));
  OAI21X1  g07314(.A0(new_n9745_), .A1(new_n7828_), .B0(new_n2939_), .Y(new_n9751_));
  AOI21X1  g07315(.A0(new_n9750_), .A1(new_n7828_), .B0(new_n9751_), .Y(new_n9752_));
  NOR3X1   g07316(.A(new_n7893_), .B(new_n7891_), .C(pi0114), .Y(new_n9753_));
  OAI21X1  g07317(.A0(new_n7898_), .A1(new_n7830_), .B0(new_n8278_), .Y(new_n9754_));
  AOI21X1  g07318(.A0(new_n9746_), .A1(new_n8279_), .B0(pi0039), .Y(new_n9755_));
  OAI21X1  g07319(.A0(new_n9754_), .A1(new_n9753_), .B0(new_n9755_), .Y(new_n9756_));
  OAI21X1  g07320(.A0(new_n9742_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n9757_));
  AOI21X1  g07321(.A0(new_n9756_), .A1(new_n5074_), .B0(new_n9757_), .Y(new_n9758_));
  OAI21X1  g07322(.A0(new_n9752_), .A1(new_n3252_), .B0(new_n9758_), .Y(new_n9759_));
  NOR3X1   g07323(.A(new_n7912_), .B(pi0115), .C(pi0114), .Y(new_n9760_));
  NOR4X1   g07324(.A(new_n7801_), .B(new_n7839_), .C(new_n7895_), .D(new_n2793_), .Y(new_n9761_));
  AOI21X1  g07325(.A0(new_n9761_), .A1(new_n7828_), .B0(new_n9746_), .Y(new_n9762_));
  OR3X1    g07326(.A(new_n9762_), .B(new_n9760_), .C(new_n3252_), .Y(new_n9763_));
  NOR2X1   g07327(.A(new_n9742_), .B(new_n3251_), .Y(new_n9764_));
  NOR2X1   g07328(.A(new_n9764_), .B(new_n8261_), .Y(new_n9765_));
  AOI21X1  g07329(.A0(new_n9765_), .A1(new_n9763_), .B0(pi0075), .Y(new_n9766_));
  AOI22X1  g07330(.A0(new_n9766_), .A1(new_n9759_), .B0(new_n9749_), .B1(new_n9748_), .Y(new_n9767_));
  MX2X1    g07331(.A(new_n9767_), .B(new_n9742_), .S0(new_n9590_), .Y(po0272));
  AND3X1   g07332(.A(pi0115), .B(new_n2530_), .C(new_n2939_), .Y(new_n9769_));
  NOR4X1   g07333(.A(pi0114), .B(pi0052), .C(pi0043), .D(pi0042), .Y(new_n9770_));
  NOR4X1   g07334(.A(new_n9770_), .B(new_n7893_), .C(new_n7695_), .D(pi0115), .Y(new_n9771_));
  OAI21X1  g07335(.A0(new_n9743_), .A1(new_n7828_), .B0(new_n9719_), .Y(new_n9772_));
  OR2X1    g07336(.A(new_n7828_), .B(pi0072), .Y(new_n9773_));
  AOI21X1  g07337(.A0(new_n9773_), .A1(new_n9720_), .B0(new_n3074_), .Y(new_n9774_));
  OAI21X1  g07338(.A0(new_n9772_), .A1(new_n9771_), .B0(new_n9774_), .Y(new_n9775_));
  AOI21X1  g07339(.A0(new_n9769_), .A1(new_n5778_), .B0(new_n3073_), .Y(new_n9776_));
  OAI21X1  g07340(.A0(new_n8011_), .A1(pi0115), .B0(new_n2939_), .Y(new_n9777_));
  AOI21X1  g07341(.A0(new_n8002_), .A1(pi0115), .B0(new_n9777_), .Y(new_n9778_));
  NOR3X1   g07342(.A(new_n9770_), .B(new_n7893_), .C(pi0115), .Y(new_n9779_));
  OAI21X1  g07343(.A0(new_n7898_), .A1(new_n7828_), .B0(new_n9719_), .Y(new_n9780_));
  AOI21X1  g07344(.A0(new_n9773_), .A1(new_n9720_), .B0(pi0039), .Y(new_n9781_));
  OAI21X1  g07345(.A0(new_n9780_), .A1(new_n9779_), .B0(new_n9781_), .Y(new_n9782_));
  OAI21X1  g07346(.A0(new_n9769_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n9783_));
  AOI21X1  g07347(.A0(new_n9782_), .A1(new_n5074_), .B0(new_n9783_), .Y(new_n9784_));
  OAI21X1  g07348(.A0(new_n9778_), .A1(new_n3252_), .B0(new_n9784_), .Y(new_n9785_));
  NOR2X1   g07349(.A(new_n7912_), .B(pi0115), .Y(new_n9786_));
  OAI21X1  g07350(.A0(new_n9773_), .A1(new_n9761_), .B0(new_n3251_), .Y(new_n9787_));
  NOR2X1   g07351(.A(new_n9769_), .B(new_n3251_), .Y(new_n9788_));
  NOR2X1   g07352(.A(new_n9788_), .B(new_n8261_), .Y(new_n9789_));
  OAI21X1  g07353(.A0(new_n9787_), .A1(new_n9786_), .B0(new_n9789_), .Y(new_n9790_));
  AND2X1   g07354(.A(new_n9790_), .B(new_n3073_), .Y(new_n9791_));
  AOI22X1  g07355(.A0(new_n9791_), .A1(new_n9785_), .B0(new_n9776_), .B1(new_n9775_), .Y(new_n9792_));
  MX2X1    g07356(.A(new_n9792_), .B(new_n9769_), .S0(new_n9590_), .Y(po0273));
  AND3X1   g07357(.A(pi0116), .B(new_n2530_), .C(new_n2939_), .Y(new_n9794_));
  AOI21X1  g07358(.A0(new_n7846_), .A1(pi0116), .B0(new_n2703_), .Y(new_n9795_));
  OR2X1    g07359(.A(new_n7835_), .B(new_n2704_), .Y(new_n9796_));
  AOI21X1  g07360(.A0(new_n9796_), .A1(pi0116), .B0(new_n7840_), .Y(new_n9797_));
  AOI21X1  g07361(.A0(new_n7850_), .A1(new_n2704_), .B0(new_n2793_), .Y(new_n9798_));
  OAI21X1  g07362(.A0(new_n9797_), .A1(new_n9795_), .B0(new_n9798_), .Y(new_n9799_));
  AND2X1   g07363(.A(new_n7858_), .B(pi0116), .Y(new_n9800_));
  OR3X1    g07364(.A(new_n9800_), .B(new_n7864_), .C(pi0228), .Y(new_n9801_));
  AND3X1   g07365(.A(new_n9801_), .B(new_n9799_), .C(new_n2939_), .Y(new_n9802_));
  AND2X1   g07366(.A(pi0116), .B(new_n2530_), .Y(new_n9803_));
  INVX1    g07367(.A(new_n9803_), .Y(new_n9804_));
  NOR2X1   g07368(.A(new_n9804_), .B(new_n9719_), .Y(new_n9805_));
  NOR4X1   g07369(.A(new_n7801_), .B(new_n7697_), .C(new_n7895_), .D(pi0113), .Y(new_n9806_));
  OR2X1    g07370(.A(new_n9806_), .B(new_n9804_), .Y(new_n9807_));
  AOI21X1  g07371(.A0(new_n9807_), .A1(new_n7893_), .B0(new_n9725_), .Y(new_n9808_));
  OAI21X1  g07372(.A0(new_n9808_), .A1(new_n9805_), .B0(new_n2939_), .Y(new_n9809_));
  OAI21X1  g07373(.A0(new_n9794_), .A1(new_n2979_), .B0(new_n3131_), .Y(new_n9810_));
  AOI21X1  g07374(.A0(new_n9809_), .A1(new_n5074_), .B0(new_n9810_), .Y(new_n9811_));
  OAI21X1  g07375(.A0(new_n9802_), .A1(new_n3252_), .B0(new_n9811_), .Y(new_n9812_));
  NOR2X1   g07376(.A(new_n9794_), .B(new_n2979_), .Y(new_n9813_));
  OAI21X1  g07377(.A0(new_n7914_), .A1(pi0113), .B0(new_n9803_), .Y(new_n9814_));
  AND3X1   g07378(.A(new_n9814_), .B(new_n7912_), .C(new_n2979_), .Y(new_n9815_));
  OAI21X1  g07379(.A0(new_n9815_), .A1(new_n9813_), .B0(new_n3007_), .Y(new_n9816_));
  NOR2X1   g07380(.A(new_n9794_), .B(new_n3007_), .Y(new_n9817_));
  NOR2X1   g07381(.A(new_n9817_), .B(new_n8261_), .Y(new_n9818_));
  AOI21X1  g07382(.A0(new_n9818_), .A1(new_n9816_), .B0(pi0075), .Y(new_n9819_));
  NOR3X1   g07383(.A(new_n7709_), .B(new_n7895_), .C(pi0113), .Y(new_n9820_));
  OAI22X1  g07384(.A0(new_n9804_), .A1(new_n9820_), .B0(new_n7893_), .B1(new_n7695_), .Y(new_n9821_));
  AOI21X1  g07385(.A0(new_n9821_), .A1(new_n9724_), .B0(new_n9805_), .Y(new_n9822_));
  OR2X1    g07386(.A(new_n9822_), .B(new_n3074_), .Y(new_n9823_));
  AOI21X1  g07387(.A0(new_n9794_), .A1(new_n5778_), .B0(new_n3073_), .Y(new_n9824_));
  AOI22X1  g07388(.A0(new_n9824_), .A1(new_n9823_), .B0(new_n9819_), .B1(new_n9812_), .Y(new_n9825_));
  MX2X1    g07389(.A(new_n9825_), .B(new_n9794_), .S0(new_n9590_), .Y(po0274));
  AOI22X1  g07390(.A0(new_n5824_), .A1(new_n3388_), .B0(new_n3181_), .B1(new_n3007_), .Y(new_n9827_));
  OAI21X1  g07391(.A0(new_n9827_), .A1(pi0038), .B0(new_n3131_), .Y(new_n9828_));
  AOI21X1  g07392(.A0(new_n9828_), .A1(new_n5091_), .B0(pi0092), .Y(new_n9829_));
  NAND3X1  g07393(.A(new_n5784_), .B(new_n4982_), .C(new_n3091_), .Y(new_n9830_));
  OR2X1    g07394(.A(new_n9830_), .B(new_n9829_), .Y(new_n9831_));
  AOI21X1  g07395(.A0(new_n9831_), .A1(new_n3107_), .B0(new_n5814_), .Y(new_n9832_));
  OAI21X1  g07396(.A0(new_n9832_), .A1(pi0056), .B0(new_n4981_), .Y(new_n9833_));
  OR3X1    g07397(.A(new_n5097_), .B(pi0059), .C(pi0057), .Y(new_n9834_));
  AOI21X1  g07398(.A0(new_n9833_), .A1(new_n3222_), .B0(new_n9834_), .Y(po0275));
  INVX1    g07399(.A(new_n7323_), .Y(new_n9836_));
  INVX1    g07400(.A(pi0150), .Y(new_n9837_));
  OAI21X1  g07401(.A0(new_n5048_), .A1(new_n8623_), .B0(new_n8625_), .Y(new_n9838_));
  NOR4X1   g07402(.A(new_n8624_), .B(new_n7308_), .C(new_n5048_), .D(new_n9837_), .Y(new_n9839_));
  AOI21X1  g07403(.A0(new_n9838_), .A1(new_n9837_), .B0(new_n9839_), .Y(new_n9840_));
  NOR3X1   g07404(.A(new_n9840_), .B(new_n6794_), .C(new_n5215_), .Y(new_n9841_));
  NOR2X1   g07405(.A(new_n9841_), .B(new_n4982_), .Y(new_n9842_));
  INVX1    g07406(.A(new_n9842_), .Y(new_n9843_));
  AOI22X1  g07407(.A0(new_n6819_), .A1(pi0165), .B0(new_n3091_), .B1(new_n2979_), .Y(new_n9844_));
  AND2X1   g07408(.A(new_n9844_), .B(new_n6794_), .Y(new_n9845_));
  OR3X1    g07409(.A(new_n9845_), .B(new_n9841_), .C(pi0074), .Y(new_n9846_));
  AOI21X1  g07410(.A0(new_n9846_), .A1(new_n9843_), .B0(new_n3123_), .Y(new_n9847_));
  OAI21X1  g07411(.A0(new_n9847_), .A1(new_n3374_), .B0(new_n9836_), .Y(new_n9848_));
  AND2X1   g07412(.A(new_n9840_), .B(pi0299), .Y(new_n9849_));
  OAI21X1  g07413(.A0(new_n8635_), .A1(pi0184), .B0(pi0185), .Y(new_n9850_));
  OR3X1    g07414(.A(new_n8635_), .B(pi0185), .C(pi0184), .Y(new_n9851_));
  NAND3X1  g07415(.A(new_n9851_), .B(new_n9850_), .C(new_n5023_), .Y(new_n9852_));
  AND2X1   g07416(.A(new_n9852_), .B(new_n2933_), .Y(new_n9853_));
  NOR4X1   g07417(.A(new_n9853_), .B(new_n9849_), .C(new_n6794_), .D(new_n5215_), .Y(new_n9854_));
  INVX1    g07418(.A(new_n9854_), .Y(new_n9855_));
  AOI21X1  g07419(.A0(new_n9855_), .A1(pi0074), .B0(pi0055), .Y(new_n9856_));
  INVX1    g07420(.A(new_n9856_), .Y(new_n9857_));
  MX2X1    g07421(.A(pi0143), .B(pi0165), .S0(pi0299), .Y(new_n9858_));
  AND3X1   g07422(.A(new_n9858_), .B(new_n5023_), .C(pi0232), .Y(new_n9859_));
  OR2X1    g07423(.A(new_n9859_), .B(new_n6809_), .Y(new_n9860_));
  AND2X1   g07424(.A(new_n9860_), .B(pi0054), .Y(new_n9861_));
  AND2X1   g07425(.A(new_n9861_), .B(new_n9855_), .Y(new_n9862_));
  INVX1    g07426(.A(new_n9862_), .Y(new_n9863_));
  OAI21X1  g07427(.A0(new_n6820_), .A1(new_n5782_), .B0(pi0143), .Y(new_n9864_));
  AND2X1   g07428(.A(new_n9864_), .B(pi0165), .Y(new_n9865_));
  OAI21X1  g07429(.A0(new_n6821_), .A1(pi0143), .B0(new_n9865_), .Y(new_n9866_));
  INVX1    g07430(.A(pi0165), .Y(new_n9867_));
  AND2X1   g07431(.A(new_n9867_), .B(pi0143), .Y(new_n9868_));
  AOI21X1  g07432(.A0(new_n9868_), .A1(new_n6829_), .B0(new_n2979_), .Y(new_n9869_));
  AOI21X1  g07433(.A0(new_n9869_), .A1(new_n9866_), .B0(new_n7156_), .Y(new_n9870_));
  AND2X1   g07434(.A(new_n7033_), .B(new_n5048_), .Y(new_n9871_));
  OR2X1    g07435(.A(pi0168), .B(new_n3347_), .Y(new_n9872_));
  OR2X1    g07436(.A(new_n9872_), .B(new_n7090_), .Y(new_n9873_));
  NAND3X1  g07437(.A(new_n7085_), .B(new_n7027_), .C(new_n4308_), .Y(new_n9874_));
  AND2X1   g07438(.A(new_n9874_), .B(new_n3347_), .Y(new_n9875_));
  OAI21X1  g07439(.A0(new_n7082_), .A1(new_n4308_), .B0(new_n9875_), .Y(new_n9876_));
  AOI21X1  g07440(.A0(new_n9876_), .A1(new_n9873_), .B0(new_n9871_), .Y(new_n9877_));
  MX2X1    g07441(.A(new_n7066_), .B(new_n7033_), .S0(new_n5048_), .Y(new_n9878_));
  NAND2X1  g07442(.A(pi0168), .B(pi0151), .Y(new_n9879_));
  OAI21X1  g07443(.A0(new_n9879_), .A1(new_n9878_), .B0(pi0150), .Y(new_n9880_));
  NOR2X1   g07444(.A(new_n7033_), .B(new_n5023_), .Y(new_n9881_));
  INVX1    g07445(.A(new_n9881_), .Y(new_n9882_));
  AND3X1   g07446(.A(new_n9882_), .B(new_n6975_), .C(pi0168), .Y(new_n9883_));
  INVX1    g07447(.A(new_n7033_), .Y(new_n9884_));
  MX2X1    g07448(.A(new_n7114_), .B(new_n9884_), .S0(new_n5048_), .Y(new_n9885_));
  OAI21X1  g07449(.A0(new_n9885_), .A1(pi0168), .B0(pi0151), .Y(new_n9886_));
  AND2X1   g07450(.A(new_n5023_), .B(pi0168), .Y(new_n9887_));
  INVX1    g07451(.A(new_n9887_), .Y(new_n9888_));
  NAND2X1  g07452(.A(new_n9888_), .B(new_n7033_), .Y(new_n9889_));
  AOI21X1  g07453(.A0(new_n7016_), .A1(pi0168), .B0(pi0151), .Y(new_n9890_));
  AOI21X1  g07454(.A0(new_n9890_), .A1(new_n9889_), .B0(pi0150), .Y(new_n9891_));
  OAI21X1  g07455(.A0(new_n9886_), .A1(new_n9883_), .B0(new_n9891_), .Y(new_n9892_));
  AND2X1   g07456(.A(new_n9892_), .B(pi0299), .Y(new_n9893_));
  OAI21X1  g07457(.A0(new_n9880_), .A1(new_n9877_), .B0(new_n9893_), .Y(new_n9894_));
  INVX1    g07458(.A(new_n9871_), .Y(new_n9895_));
  AOI21X1  g07459(.A0(new_n9895_), .A1(new_n7010_), .B0(pi0173), .Y(new_n9896_));
  NOR2X1   g07460(.A(new_n6967_), .B(new_n5048_), .Y(new_n9897_));
  OAI21X1  g07461(.A0(new_n7033_), .A1(new_n5023_), .B0(pi0173), .Y(new_n9898_));
  OAI21X1  g07462(.A0(new_n9898_), .A1(new_n9897_), .B0(pi0185), .Y(new_n9899_));
  INVX1    g07463(.A(pi0190), .Y(new_n9900_));
  NAND3X1  g07464(.A(new_n9882_), .B(new_n6975_), .C(pi0173), .Y(new_n9901_));
  INVX1    g07465(.A(pi0185), .Y(new_n9902_));
  INVX1    g07466(.A(pi0173), .Y(new_n9903_));
  OAI21X1  g07467(.A0(new_n9871_), .A1(new_n7016_), .B0(new_n9903_), .Y(new_n9904_));
  AND2X1   g07468(.A(new_n9904_), .B(new_n9902_), .Y(new_n9905_));
  AOI21X1  g07469(.A0(new_n9905_), .A1(new_n9901_), .B0(new_n9900_), .Y(new_n9906_));
  OAI21X1  g07470(.A0(new_n9899_), .A1(new_n9896_), .B0(new_n9906_), .Y(new_n9907_));
  AOI21X1  g07471(.A0(new_n7089_), .A1(new_n6948_), .B0(new_n9903_), .Y(new_n9908_));
  OAI21X1  g07472(.A0(new_n7030_), .A1(pi0173), .B0(new_n5023_), .Y(new_n9909_));
  AOI21X1  g07473(.A0(new_n7033_), .A1(new_n5048_), .B0(new_n9902_), .Y(new_n9910_));
  OAI21X1  g07474(.A0(new_n9909_), .A1(new_n9908_), .B0(new_n9910_), .Y(new_n9911_));
  AOI21X1  g07475(.A0(new_n7033_), .A1(new_n9903_), .B0(pi0185), .Y(new_n9912_));
  OAI21X1  g07476(.A0(new_n9885_), .A1(new_n9903_), .B0(new_n9912_), .Y(new_n9913_));
  AND2X1   g07477(.A(new_n9913_), .B(new_n9900_), .Y(new_n9914_));
  AOI21X1  g07478(.A0(new_n9914_), .A1(new_n9911_), .B0(pi0299), .Y(new_n9915_));
  AOI21X1  g07479(.A0(new_n9915_), .A1(new_n9907_), .B0(new_n5215_), .Y(new_n9916_));
  OAI21X1  g07480(.A0(new_n9884_), .A1(pi0232), .B0(new_n2939_), .Y(new_n9917_));
  AOI21X1  g07481(.A0(new_n9916_), .A1(new_n9894_), .B0(new_n9917_), .Y(new_n9918_));
  AOI22X1  g07482(.A0(new_n8770_), .A1(pi0157), .B0(new_n6866_), .B1(pi0168), .Y(new_n9919_));
  NOR4X1   g07483(.A(new_n9919_), .B(new_n7187_), .C(new_n5058_), .D(new_n5048_), .Y(new_n9920_));
  MX2X1    g07484(.A(new_n9920_), .B(pi0178), .S0(new_n2933_), .Y(new_n9921_));
  AOI21X1  g07485(.A0(new_n6875_), .A1(pi0178), .B0(pi0190), .Y(new_n9922_));
  OAI22X1  g07486(.A0(new_n9922_), .A1(pi0299), .B0(new_n9921_), .B1(new_n6835_), .Y(new_n9923_));
  AOI21X1  g07487(.A0(new_n6835_), .A1(new_n5041_), .B0(new_n7203_), .Y(new_n9924_));
  AND3X1   g07488(.A(new_n9924_), .B(new_n6853_), .C(new_n6801_), .Y(new_n9925_));
  AND3X1   g07489(.A(new_n9924_), .B(new_n6879_), .C(pi0178), .Y(new_n9926_));
  OAI21X1  g07490(.A0(new_n6848_), .A1(new_n6835_), .B0(new_n2933_), .Y(new_n9927_));
  OR4X1    g07491(.A(new_n9927_), .B(new_n9926_), .C(new_n9925_), .D(new_n9900_), .Y(new_n9928_));
  AND3X1   g07492(.A(new_n9928_), .B(new_n9923_), .C(pi0232), .Y(new_n9929_));
  OAI21X1  g07493(.A0(new_n6835_), .A1(pi0232), .B0(pi0039), .Y(new_n9930_));
  OAI21X1  g07494(.A0(new_n9930_), .A1(new_n9929_), .B0(new_n2979_), .Y(new_n9931_));
  OAI21X1  g07495(.A0(new_n9931_), .A1(new_n9918_), .B0(new_n9870_), .Y(new_n9932_));
  NOR3X1   g07496(.A(new_n9853_), .B(new_n9849_), .C(new_n5215_), .Y(new_n9933_));
  NOR2X1   g07497(.A(new_n9933_), .B(new_n3007_), .Y(new_n9934_));
  OR2X1    g07498(.A(new_n9859_), .B(new_n2979_), .Y(new_n9935_));
  AND2X1   g07499(.A(new_n9935_), .B(new_n7288_), .Y(new_n9936_));
  AOI21X1  g07500(.A0(new_n9936_), .A1(new_n7465_), .B0(new_n9934_), .Y(new_n9937_));
  AOI21X1  g07501(.A0(new_n9937_), .A1(new_n9932_), .B0(new_n5295_), .Y(new_n9938_));
  AND2X1   g07502(.A(new_n9935_), .B(new_n3007_), .Y(new_n9939_));
  INVX1    g07503(.A(new_n9939_), .Y(new_n9940_));
  MX2X1    g07504(.A(pi0178), .B(pi0157), .S0(pi0299), .Y(new_n9941_));
  AND3X1   g07505(.A(new_n9941_), .B(new_n5023_), .C(pi0232), .Y(new_n9942_));
  NAND4X1  g07506(.A(new_n9942_), .B(new_n6843_), .C(new_n3131_), .D(new_n2939_), .Y(new_n9943_));
  AOI21X1  g07507(.A0(new_n9943_), .A1(new_n7179_), .B0(new_n9940_), .Y(new_n9944_));
  OAI21X1  g07508(.A0(new_n9944_), .A1(new_n9934_), .B0(new_n7138_), .Y(new_n9945_));
  OAI21X1  g07509(.A0(new_n9933_), .A1(new_n3073_), .B0(new_n9945_), .Y(new_n9946_));
  OAI21X1  g07510(.A0(new_n9946_), .A1(new_n9938_), .B0(new_n3091_), .Y(new_n9947_));
  AOI21X1  g07511(.A0(new_n9947_), .A1(new_n9863_), .B0(pi0074), .Y(new_n9948_));
  NOR2X1   g07512(.A(new_n9842_), .B(new_n3107_), .Y(new_n9949_));
  NOR2X1   g07513(.A(new_n9841_), .B(pi0074), .Y(new_n9950_));
  NAND3X1  g07514(.A(new_n5023_), .B(pi0232), .C(pi0150), .Y(new_n9951_));
  OR4X1    g07515(.A(new_n9951_), .B(new_n7142_), .C(new_n7141_), .D(pi0092), .Y(new_n9952_));
  AND3X1   g07516(.A(new_n6834_), .B(new_n3091_), .C(new_n2979_), .Y(new_n9953_));
  AOI21X1  g07517(.A0(new_n9953_), .A1(new_n9952_), .B0(new_n9844_), .Y(new_n9954_));
  OAI21X1  g07518(.A0(new_n9954_), .A1(new_n6809_), .B0(new_n9950_), .Y(new_n9955_));
  AOI21X1  g07519(.A0(new_n9955_), .A1(new_n9949_), .B0(new_n4975_), .Y(new_n9956_));
  OAI21X1  g07520(.A0(new_n9948_), .A1(new_n9857_), .B0(new_n9956_), .Y(new_n9957_));
  OAI21X1  g07521(.A0(new_n9840_), .A1(new_n5215_), .B0(new_n6809_), .Y(new_n9958_));
  NAND4X1  g07522(.A(new_n6794_), .B(new_n5023_), .C(pi0232), .D(pi0165), .Y(new_n9959_));
  AND3X1   g07523(.A(new_n9959_), .B(new_n9958_), .C(new_n3374_), .Y(new_n9960_));
  AND2X1   g07524(.A(new_n9960_), .B(new_n9843_), .Y(new_n9961_));
  AOI21X1  g07525(.A0(new_n9957_), .A1(new_n9848_), .B0(new_n9961_), .Y(new_n9962_));
  NOR4X1   g07526(.A(pi0954), .B(pi0079), .C(pi0034), .D(pi0033), .Y(new_n9963_));
  INVX1    g07527(.A(new_n9963_), .Y(new_n9964_));
  OR2X1    g07528(.A(new_n9847_), .B(new_n3374_), .Y(new_n9965_));
  INVX1    g07529(.A(new_n9961_), .Y(new_n9966_));
  INVX1    g07530(.A(new_n9870_), .Y(new_n9967_));
  INVX1    g07531(.A(pi0157), .Y(new_n9968_));
  AOI21X1  g07532(.A0(new_n7193_), .A1(new_n9968_), .B0(new_n4308_), .Y(new_n9969_));
  OR2X1    g07533(.A(pi0168), .B(pi0157), .Y(new_n9970_));
  OAI22X1  g07534(.A0(new_n9970_), .A1(new_n7509_), .B0(new_n7189_), .B1(new_n9968_), .Y(new_n9971_));
  OAI22X1  g07535(.A0(new_n9971_), .A1(new_n9969_), .B0(new_n5236_), .B1(new_n6256_), .Y(new_n9972_));
  INVX1    g07536(.A(new_n9494_), .Y(new_n9973_));
  NAND4X1  g07537(.A(new_n7192_), .B(new_n5042_), .C(new_n5023_), .D(new_n6801_), .Y(new_n9974_));
  OAI21X1  g07538(.A0(new_n5236_), .A1(new_n6256_), .B0(new_n9974_), .Y(new_n9975_));
  NOR2X1   g07539(.A(new_n7200_), .B(new_n6801_), .Y(new_n9976_));
  OAI21X1  g07540(.A0(new_n5236_), .A1(new_n6256_), .B0(new_n9976_), .Y(new_n9977_));
  AOI21X1  g07541(.A0(new_n9512_), .A1(new_n6801_), .B0(pi0190), .Y(new_n9978_));
  AOI22X1  g07542(.A0(new_n9978_), .A1(new_n9977_), .B0(new_n9975_), .B1(pi0190), .Y(new_n9979_));
  OAI21X1  g07543(.A0(new_n9979_), .A1(new_n9973_), .B0(pi0232), .Y(new_n9980_));
  AOI21X1  g07544(.A0(new_n9972_), .A1(new_n9493_), .B0(new_n9980_), .Y(new_n9981_));
  NOR3X1   g07545(.A(new_n7203_), .B(new_n5787_), .C(new_n5236_), .Y(new_n9982_));
  OR4X1    g07546(.A(new_n5062_), .B(new_n4890_), .C(new_n2437_), .D(new_n2438_), .Y(new_n9983_));
  OAI21X1  g07547(.A0(new_n9983_), .A1(new_n5236_), .B0(new_n5215_), .Y(new_n9984_));
  OAI21X1  g07548(.A0(new_n9984_), .A1(new_n9982_), .B0(pi0039), .Y(new_n9985_));
  NOR2X1   g07549(.A(new_n7238_), .B(new_n4308_), .Y(new_n9986_));
  OAI21X1  g07550(.A0(new_n7227_), .A1(pi0168), .B0(new_n3347_), .Y(new_n9987_));
  OAI22X1  g07551(.A0(new_n9987_), .A1(new_n9986_), .B0(new_n9872_), .B1(new_n7251_), .Y(new_n9988_));
  AOI21X1  g07552(.A0(new_n9988_), .A1(new_n7229_), .B0(new_n9837_), .Y(new_n9989_));
  OAI21X1  g07553(.A0(new_n7219_), .A1(pi0151), .B0(new_n7486_), .Y(new_n9990_));
  NAND2X1  g07554(.A(new_n7235_), .B(new_n3347_), .Y(new_n9991_));
  AOI21X1  g07555(.A0(new_n9991_), .A1(new_n7263_), .B0(new_n9888_), .Y(new_n9992_));
  OR2X1    g07556(.A(new_n9992_), .B(pi0150), .Y(new_n9993_));
  AOI21X1  g07557(.A0(new_n9990_), .A1(new_n4308_), .B0(new_n9993_), .Y(new_n9994_));
  AOI21X1  g07558(.A0(new_n8858_), .A1(new_n7219_), .B0(new_n5023_), .Y(new_n9995_));
  NOR2X1   g07559(.A(new_n9995_), .B(new_n2933_), .Y(new_n9996_));
  OAI21X1  g07560(.A0(new_n9994_), .A1(new_n9989_), .B0(new_n9996_), .Y(new_n9997_));
  NOR2X1   g07561(.A(new_n7251_), .B(new_n7619_), .Y(new_n9998_));
  INVX1    g07562(.A(new_n9998_), .Y(new_n9999_));
  NAND3X1  g07563(.A(new_n7227_), .B(new_n5168_), .C(new_n9903_), .Y(new_n10000_));
  OAI21X1  g07564(.A0(new_n9999_), .A1(new_n9903_), .B0(new_n10000_), .Y(new_n10001_));
  NOR3X1   g07565(.A(pi0468), .B(pi0332), .C(pi0190), .Y(new_n10002_));
  NAND4X1  g07566(.A(new_n7238_), .B(new_n7229_), .C(pi0190), .D(new_n9903_), .Y(new_n10003_));
  NAND2X1  g07567(.A(new_n10003_), .B(pi0185), .Y(new_n10004_));
  AOI21X1  g07568(.A0(new_n10002_), .A1(new_n10001_), .B0(new_n10004_), .Y(new_n10005_));
  OAI21X1  g07569(.A0(new_n7219_), .A1(pi0173), .B0(new_n7244_), .Y(new_n10006_));
  OR3X1    g07570(.A(new_n8855_), .B(new_n5198_), .C(new_n9903_), .Y(new_n10007_));
  NAND4X1  g07571(.A(new_n10007_), .B(new_n7236_), .C(new_n5023_), .D(pi0190), .Y(new_n10008_));
  NAND2X1  g07572(.A(new_n10008_), .B(new_n9902_), .Y(new_n10009_));
  AOI21X1  g07573(.A0(new_n10006_), .A1(new_n9900_), .B0(new_n10009_), .Y(new_n10010_));
  AOI21X1  g07574(.A0(new_n7223_), .A1(new_n5048_), .B0(pi0299), .Y(new_n10011_));
  OAI21X1  g07575(.A0(new_n10010_), .A1(new_n10005_), .B0(new_n10011_), .Y(new_n10012_));
  AOI21X1  g07576(.A0(new_n10012_), .A1(new_n9997_), .B0(new_n5215_), .Y(new_n10013_));
  NOR2X1   g07577(.A(new_n7222_), .B(new_n5009_), .Y(new_n10014_));
  OR2X1    g07578(.A(new_n7218_), .B(pi0232), .Y(new_n10015_));
  OAI21X1  g07579(.A0(new_n10015_), .A1(new_n10014_), .B0(new_n2939_), .Y(new_n10016_));
  OAI22X1  g07580(.A0(new_n10016_), .A1(new_n10013_), .B0(new_n9985_), .B1(new_n9981_), .Y(new_n10017_));
  AOI21X1  g07581(.A0(new_n10017_), .A1(new_n2979_), .B0(new_n9967_), .Y(new_n10018_));
  OR2X1    g07582(.A(new_n9936_), .B(new_n9934_), .Y(new_n10019_));
  OAI21X1  g07583(.A0(new_n10019_), .A1(new_n10018_), .B0(new_n3084_), .Y(new_n10020_));
  NOR2X1   g07584(.A(new_n9933_), .B(new_n3073_), .Y(new_n10021_));
  NOR4X1   g07585(.A(new_n9942_), .B(new_n3060_), .C(new_n2986_), .D(pi0087), .Y(new_n10022_));
  OAI22X1  g07586(.A0(new_n10022_), .A1(new_n9940_), .B0(new_n9933_), .B1(new_n3007_), .Y(new_n10023_));
  AOI21X1  g07587(.A0(new_n10023_), .A1(new_n7138_), .B0(new_n10021_), .Y(new_n10024_));
  AOI21X1  g07588(.A0(new_n10024_), .A1(new_n10020_), .B0(pi0054), .Y(new_n10025_));
  OAI21X1  g07589(.A0(new_n10025_), .A1(new_n9862_), .B0(new_n4982_), .Y(new_n10026_));
  NAND4X1  g07590(.A(new_n5023_), .B(pi0232), .C(pi0165), .D(pi0054), .Y(new_n10027_));
  AND3X1   g07591(.A(new_n6794_), .B(new_n6777_), .C(new_n3079_), .Y(new_n10028_));
  AND3X1   g07592(.A(new_n10028_), .B(new_n10027_), .C(new_n9951_), .Y(new_n10029_));
  AOI21X1  g07593(.A0(new_n10029_), .A1(new_n2987_), .B0(new_n9846_), .Y(new_n10030_));
  NOR3X1   g07594(.A(new_n10030_), .B(new_n9842_), .C(new_n3107_), .Y(new_n10031_));
  OR2X1    g07595(.A(new_n10031_), .B(new_n4975_), .Y(new_n10032_));
  AOI21X1  g07596(.A0(new_n10026_), .A1(new_n9856_), .B0(new_n10032_), .Y(new_n10033_));
  OAI21X1  g07597(.A0(new_n10033_), .A1(new_n9965_), .B0(new_n9966_), .Y(new_n10034_));
  OAI21X1  g07598(.A0(new_n10034_), .A1(pi0118), .B0(new_n9964_), .Y(new_n10035_));
  AOI21X1  g07599(.A0(new_n9962_), .A1(pi0118), .B0(new_n10035_), .Y(new_n10036_));
  NOR2X1   g07600(.A(new_n6786_), .B(pi0118), .Y(new_n10037_));
  OAI21X1  g07601(.A0(new_n10037_), .A1(new_n10034_), .B0(new_n9963_), .Y(new_n10038_));
  AOI21X1  g07602(.A0(new_n10037_), .A1(new_n9962_), .B0(new_n10038_), .Y(new_n10039_));
  OR2X1    g07603(.A(new_n10039_), .B(new_n10036_), .Y(po0276));
  NAND2X1  g07604(.A(pi0228), .B(pi0128), .Y(new_n10041_));
  INVX1    g07605(.A(pi0128), .Y(new_n10042_));
  NAND3X1  g07606(.A(new_n9456_), .B(new_n4769_), .C(new_n2952_), .Y(new_n10043_));
  NOR2X1   g07607(.A(pi0221), .B(pi0216), .Y(new_n10044_));
  INVX1    g07608(.A(new_n10044_), .Y(new_n10045_));
  NAND3X1  g07609(.A(new_n5948_), .B(new_n4889_), .C(new_n10045_), .Y(new_n10046_));
  AOI21X1  g07610(.A0(new_n10046_), .A1(new_n10043_), .B0(new_n2939_), .Y(new_n10047_));
  NAND4X1  g07611(.A(new_n7603_), .B(new_n2643_), .C(new_n2560_), .D(new_n2594_), .Y(new_n10048_));
  AOI21X1  g07612(.A0(new_n10048_), .A1(new_n8615_), .B0(new_n2573_), .Y(new_n10049_));
  NOR4X1   g07613(.A(new_n2831_), .B(new_n2565_), .C(pi0108), .D(pi0046), .Y(new_n10050_));
  OAI21X1  g07614(.A0(new_n10049_), .A1(pi0097), .B0(new_n10050_), .Y(new_n10051_));
  NOR4X1   g07615(.A(new_n8615_), .B(new_n2573_), .C(new_n2473_), .D(pi0046), .Y(new_n10052_));
  MX2X1    g07616(.A(new_n5206_), .B(new_n5114_), .S0(pi0299), .Y(new_n10053_));
  NAND2X1  g07617(.A(new_n10053_), .B(new_n6819_), .Y(new_n10054_));
  AOI22X1  g07618(.A0(new_n10054_), .A1(pi0109), .B0(new_n10052_), .B1(new_n2831_), .Y(new_n10055_));
  MX2X1    g07619(.A(new_n5181_), .B(new_n5153_), .S0(new_n10054_), .Y(new_n10056_));
  AOI21X1  g07620(.A0(new_n10055_), .A1(new_n10051_), .B0(new_n10056_), .Y(new_n10057_));
  AOI21X1  g07621(.A0(new_n5149_), .A1(pi0091), .B0(new_n2728_), .Y(new_n10058_));
  OAI21X1  g07622(.A0(new_n10057_), .A1(pi0091), .B0(new_n10058_), .Y(new_n10059_));
  NAND4X1  g07623(.A(new_n2984_), .B(new_n2517_), .C(new_n2513_), .D(new_n2939_), .Y(new_n10060_));
  AOI21X1  g07624(.A0(new_n10059_), .A1(new_n2541_), .B0(new_n10060_), .Y(new_n10061_));
  OAI21X1  g07625(.A0(new_n10061_), .A1(new_n10047_), .B0(new_n2979_), .Y(new_n10062_));
  MX2X1    g07626(.A(new_n10062_), .B(new_n10042_), .S0(pi0228), .Y(new_n10063_));
  OAI21X1  g07627(.A0(new_n3604_), .A1(new_n3060_), .B0(new_n10041_), .Y(new_n10064_));
  AOI21X1  g07628(.A0(new_n10064_), .A1(pi0100), .B0(pi0087), .Y(new_n10065_));
  OAI21X1  g07629(.A0(new_n10063_), .A1(pi0100), .B0(new_n10065_), .Y(new_n10066_));
  AOI21X1  g07630(.A0(new_n10041_), .A1(pi0087), .B0(pi0075), .Y(new_n10067_));
  AOI22X1  g07631(.A0(new_n6777_), .A1(new_n5827_), .B0(pi0228), .B1(pi0128), .Y(new_n10068_));
  OAI21X1  g07632(.A0(new_n10068_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n10069_));
  AOI21X1  g07633(.A0(new_n10067_), .A1(new_n10066_), .B0(new_n10069_), .Y(new_n10070_));
  NAND2X1  g07634(.A(new_n10041_), .B(pi0092), .Y(new_n10071_));
  OAI21X1  g07635(.A0(new_n10071_), .A1(new_n5834_), .B0(new_n7607_), .Y(new_n10072_));
  OAI22X1  g07636(.A0(new_n10072_), .A1(new_n10070_), .B0(new_n10041_), .B1(new_n7607_), .Y(po0277));
  INVX1    g07637(.A(pi0031), .Y(new_n10074_));
  AND3X1   g07638(.A(pi0818), .B(new_n9423_), .C(new_n10074_), .Y(new_n10075_));
  INVX1    g07639(.A(new_n10075_), .Y(new_n10076_));
  AND2X1   g07640(.A(new_n6246_), .B(new_n2702_), .Y(new_n10077_));
  AOI21X1  g07641(.A0(new_n10077_), .A1(new_n6295_), .B0(new_n6072_), .Y(new_n10078_));
  OR3X1    g07642(.A(new_n5880_), .B(pi1093), .C(pi0120), .Y(new_n10079_));
  AND2X1   g07643(.A(new_n10079_), .B(new_n10078_), .Y(new_n10080_));
  NOR3X1   g07644(.A(new_n5923_), .B(new_n2985_), .C(new_n2536_), .Y(new_n10081_));
  INVX1    g07645(.A(pi0120), .Y(new_n10082_));
  AOI21X1  g07646(.A0(new_n6246_), .A1(new_n2702_), .B0(new_n10082_), .Y(new_n10083_));
  INVX1    g07647(.A(new_n10083_), .Y(new_n10084_));
  OAI21X1  g07648(.A0(new_n10084_), .A1(new_n5960_), .B0(new_n10081_), .Y(new_n10085_));
  AND2X1   g07649(.A(pi1093), .B(new_n10082_), .Y(new_n10086_));
  INVX1    g07650(.A(new_n10086_), .Y(new_n10087_));
  NAND2X1  g07651(.A(new_n10087_), .B(new_n5960_), .Y(new_n10088_));
  NOR3X1   g07652(.A(new_n5920_), .B(new_n3060_), .C(new_n2793_), .Y(new_n10089_));
  INVX1    g07653(.A(new_n10089_), .Y(new_n10090_));
  AOI21X1  g07654(.A0(new_n10088_), .A1(new_n10085_), .B0(new_n10090_), .Y(new_n10091_));
  AND2X1   g07655(.A(new_n5927_), .B(new_n5906_), .Y(new_n10092_));
  AOI21X1  g07656(.A0(new_n10092_), .A1(new_n2702_), .B0(new_n10087_), .Y(new_n10093_));
  NOR2X1   g07657(.A(new_n10093_), .B(new_n10083_), .Y(new_n10094_));
  NOR3X1   g07658(.A(new_n10094_), .B(new_n10091_), .C(new_n3007_), .Y(new_n10095_));
  NAND4X1  g07659(.A(new_n5909_), .B(new_n5902_), .C(new_n5032_), .D(pi0120), .Y(new_n10096_));
  NAND2X1  g07660(.A(new_n10096_), .B(new_n2939_), .Y(new_n10097_));
  INVX1    g07661(.A(new_n2759_), .Y(new_n10098_));
  NAND2X1  g07662(.A(new_n7737_), .B(new_n5937_), .Y(new_n10099_));
  NOR4X1   g07663(.A(new_n5928_), .B(new_n5900_), .C(new_n5881_), .D(pi0096), .Y(new_n10100_));
  AOI21X1  g07664(.A0(new_n10100_), .A1(new_n5237_), .B0(pi0122), .Y(new_n10101_));
  OAI21X1  g07665(.A0(new_n5901_), .A1(new_n5906_), .B0(new_n8194_), .Y(new_n10102_));
  AOI21X1  g07666(.A0(new_n10101_), .A1(new_n10099_), .B0(new_n10102_), .Y(new_n10103_));
  OR3X1    g07667(.A(new_n10100_), .B(new_n10092_), .C(new_n5968_), .Y(new_n10104_));
  OAI21X1  g07668(.A0(new_n10103_), .A1(new_n10098_), .B0(new_n10104_), .Y(new_n10105_));
  INVX1    g07669(.A(new_n10094_), .Y(new_n10106_));
  INVX1    g07670(.A(new_n10093_), .Y(new_n10107_));
  NOR3X1   g07671(.A(new_n5224_), .B(new_n2724_), .C(new_n5922_), .Y(new_n10108_));
  AND3X1   g07672(.A(new_n10108_), .B(pi1092), .C(pi1091), .Y(new_n10109_));
  OAI22X1  g07673(.A0(new_n10109_), .A1(new_n10107_), .B0(new_n10084_), .B1(new_n7192_), .Y(new_n10110_));
  MX2X1    g07674(.A(new_n10110_), .B(new_n10106_), .S0(new_n6256_), .Y(new_n10111_));
  NAND2X1  g07675(.A(new_n10111_), .B(new_n5058_), .Y(new_n10112_));
  MX2X1    g07676(.A(new_n10110_), .B(new_n10106_), .S0(new_n5043_), .Y(new_n10113_));
  AOI21X1  g07677(.A0(new_n10113_), .A1(new_n5059_), .B0(new_n6271_), .Y(new_n10114_));
  OAI21X1  g07678(.A0(new_n10106_), .A1(new_n6270_), .B0(pi0299), .Y(new_n10115_));
  AOI21X1  g07679(.A0(new_n10114_), .A1(new_n10112_), .B0(new_n10115_), .Y(new_n10116_));
  NAND2X1  g07680(.A(new_n10111_), .B(new_n5041_), .Y(new_n10117_));
  AOI21X1  g07681(.A0(new_n10113_), .A1(new_n5042_), .B0(new_n6265_), .Y(new_n10118_));
  OR3X1    g07682(.A(new_n10093_), .B(new_n10083_), .C(new_n6264_), .Y(new_n10119_));
  NAND2X1  g07683(.A(new_n10119_), .B(new_n2933_), .Y(new_n10120_));
  AOI21X1  g07684(.A0(new_n10118_), .A1(new_n10117_), .B0(new_n10120_), .Y(new_n10121_));
  OR3X1    g07685(.A(new_n10121_), .B(new_n10116_), .C(new_n2939_), .Y(new_n10122_));
  OAI21X1  g07686(.A0(new_n10105_), .A1(new_n10097_), .B0(new_n10122_), .Y(new_n10123_));
  INVX1    g07687(.A(new_n10077_), .Y(new_n10124_));
  NOR2X1   g07688(.A(pi1093), .B(pi0120), .Y(new_n10125_));
  AOI21X1  g07689(.A0(new_n10125_), .A1(pi0038), .B0(pi0100), .Y(new_n10126_));
  OAI21X1  g07690(.A0(new_n10124_), .A1(new_n2979_), .B0(new_n10126_), .Y(new_n10127_));
  AOI21X1  g07691(.A0(new_n10123_), .A1(new_n2979_), .B0(new_n10127_), .Y(new_n10128_));
  OAI21X1  g07692(.A0(new_n10128_), .A1(new_n10095_), .B0(new_n3131_), .Y(new_n10129_));
  OR3X1    g07693(.A(new_n10125_), .B(new_n5973_), .C(new_n3131_), .Y(new_n10130_));
  NOR3X1   g07694(.A(new_n10092_), .B(new_n6287_), .C(new_n5968_), .Y(new_n10131_));
  OR3X1    g07695(.A(new_n10131_), .B(new_n5972_), .C(new_n3132_), .Y(new_n10132_));
  NAND3X1  g07696(.A(new_n6246_), .B(new_n3132_), .C(new_n2702_), .Y(new_n10133_));
  NAND3X1  g07697(.A(new_n10133_), .B(new_n10132_), .C(pi0087), .Y(new_n10134_));
  OR2X1    g07698(.A(new_n10134_), .B(new_n10130_), .Y(new_n10135_));
  AOI21X1  g07699(.A0(new_n10135_), .A1(new_n10129_), .B0(pi0075), .Y(new_n10136_));
  NOR2X1   g07700(.A(new_n10107_), .B(new_n5924_), .Y(new_n10137_));
  NOR2X1   g07701(.A(new_n6246_), .B(pi1091), .Y(new_n10138_));
  NOR2X1   g07702(.A(new_n10138_), .B(new_n6240_), .Y(new_n10139_));
  OAI21X1  g07703(.A0(new_n10139_), .A1(new_n10082_), .B0(new_n9672_), .Y(new_n10140_));
  OAI22X1  g07704(.A0(new_n10140_), .A1(new_n10137_), .B0(new_n10106_), .B1(new_n9672_), .Y(new_n10141_));
  OAI21X1  g07705(.A0(new_n10106_), .A1(new_n3070_), .B0(pi0075), .Y(new_n10142_));
  AOI21X1  g07706(.A0(new_n10141_), .A1(new_n3070_), .B0(new_n10142_), .Y(new_n10143_));
  OR2X1    g07707(.A(new_n10143_), .B(new_n6295_), .Y(new_n10144_));
  OAI21X1  g07708(.A0(new_n10144_), .A1(new_n10136_), .B0(new_n10080_), .Y(new_n10145_));
  INVX1    g07709(.A(new_n10126_), .Y(new_n10146_));
  OAI22X1  g07710(.A0(new_n10103_), .A1(new_n10098_), .B0(new_n10100_), .B1(new_n5968_), .Y(new_n10147_));
  OR3X1    g07711(.A(new_n5059_), .B(new_n6255_), .C(new_n5032_), .Y(new_n10148_));
  AOI21X1  g07712(.A0(new_n5059_), .A1(new_n5043_), .B0(new_n6271_), .Y(new_n10149_));
  AND2X1   g07713(.A(new_n10149_), .B(new_n10148_), .Y(new_n10150_));
  OAI21X1  g07714(.A0(pi1093), .A1(pi0120), .B0(pi0299), .Y(new_n10151_));
  AOI21X1  g07715(.A0(new_n10150_), .A1(new_n7192_), .B0(new_n10151_), .Y(new_n10152_));
  OR3X1    g07716(.A(new_n6255_), .B(new_n5042_), .C(new_n5032_), .Y(new_n10153_));
  AOI21X1  g07717(.A0(new_n5043_), .A1(new_n5042_), .B0(new_n6265_), .Y(new_n10154_));
  AND3X1   g07718(.A(new_n10154_), .B(new_n10153_), .C(new_n7192_), .Y(new_n10155_));
  OR2X1    g07719(.A(new_n10125_), .B(pi0299), .Y(new_n10156_));
  OAI21X1  g07720(.A0(new_n10156_), .A1(new_n10155_), .B0(pi0039), .Y(new_n10157_));
  OAI22X1  g07721(.A0(new_n10157_), .A1(new_n10152_), .B0(new_n10147_), .B1(new_n10097_), .Y(new_n10158_));
  AOI21X1  g07722(.A0(new_n10158_), .A1(new_n2979_), .B0(new_n10146_), .Y(new_n10159_));
  MX2X1    g07723(.A(new_n10081_), .B(new_n5960_), .S0(pi0120), .Y(new_n10160_));
  OAI21X1  g07724(.A0(pi1093), .A1(pi0120), .B0(pi0100), .Y(new_n10161_));
  AOI21X1  g07725(.A0(new_n10160_), .A1(new_n10089_), .B0(new_n10161_), .Y(new_n10162_));
  OAI21X1  g07726(.A0(new_n10162_), .A1(new_n10159_), .B0(new_n3131_), .Y(new_n10163_));
  AOI21X1  g07727(.A0(new_n10163_), .A1(new_n10130_), .B0(pi0075), .Y(new_n10164_));
  INVX1    g07728(.A(new_n5981_), .Y(new_n10165_));
  OAI21X1  g07729(.A0(new_n10125_), .A1(new_n10165_), .B0(new_n5880_), .Y(new_n10166_));
  AND2X1   g07730(.A(new_n10079_), .B(new_n6072_), .Y(new_n10167_));
  OAI21X1  g07731(.A0(new_n10166_), .A1(new_n10164_), .B0(new_n10167_), .Y(new_n10168_));
  AOI21X1  g07732(.A0(new_n10168_), .A1(new_n10145_), .B0(new_n10076_), .Y(new_n10169_));
  OR3X1    g07733(.A(new_n10093_), .B(new_n10083_), .C(new_n6072_), .Y(new_n10170_));
  NAND2X1  g07734(.A(new_n10170_), .B(pi0120), .Y(new_n10171_));
  INVX1    g07735(.A(new_n10125_), .Y(new_n10172_));
  AND3X1   g07736(.A(new_n10170_), .B(new_n10172_), .C(new_n10075_), .Y(new_n10173_));
  NOR2X1   g07737(.A(new_n10173_), .B(new_n6489_), .Y(new_n10174_));
  AOI21X1  g07738(.A0(new_n10174_), .A1(new_n10171_), .B0(new_n6713_), .Y(new_n10175_));
  AND3X1   g07739(.A(pi1092), .B(pi0982), .C(pi0951), .Y(new_n10176_));
  AOI21X1  g07740(.A0(new_n10176_), .A1(pi1093), .B0(pi0120), .Y(new_n10177_));
  INVX1    g07741(.A(new_n10177_), .Y(new_n10178_));
  AND2X1   g07742(.A(new_n10178_), .B(new_n10170_), .Y(new_n10179_));
  NOR3X1   g07743(.A(new_n10179_), .B(new_n10173_), .C(new_n6489_), .Y(new_n10180_));
  NOR2X1   g07744(.A(new_n10180_), .B(new_n8943_), .Y(new_n10181_));
  OAI22X1  g07745(.A0(new_n10181_), .A1(new_n10175_), .B0(new_n10169_), .B1(po1038), .Y(new_n10182_));
  INVX1    g07746(.A(new_n10080_), .Y(new_n10183_));
  NAND3X1  g07747(.A(new_n5924_), .B(pi1093), .C(pi0120), .Y(new_n10184_));
  AND3X1   g07748(.A(new_n10176_), .B(pi1093), .C(new_n2702_), .Y(new_n10185_));
  NOR2X1   g07749(.A(new_n10185_), .B(pi0120), .Y(new_n10186_));
  AND2X1   g07750(.A(new_n10176_), .B(new_n2759_), .Y(new_n10187_));
  OR4X1    g07751(.A(pi0122), .B(pi0096), .C(pi0093), .D(pi0072), .Y(new_n10188_));
  OR4X1    g07752(.A(new_n10188_), .B(new_n6731_), .C(new_n2724_), .D(new_n5172_), .Y(new_n10189_));
  OR4X1    g07753(.A(new_n10189_), .B(new_n7708_), .C(new_n5082_), .D(new_n5922_), .Y(new_n10190_));
  OAI21X1  g07754(.A0(new_n10190_), .A1(new_n8390_), .B0(new_n10187_), .Y(new_n10191_));
  NAND2X1  g07755(.A(new_n10191_), .B(new_n10186_), .Y(new_n10192_));
  AOI21X1  g07756(.A0(new_n10192_), .A1(new_n10184_), .B0(new_n5920_), .Y(new_n10193_));
  OAI21X1  g07757(.A0(new_n10178_), .A1(new_n9672_), .B0(new_n3070_), .Y(new_n10194_));
  AOI21X1  g07758(.A0(new_n10178_), .A1(new_n3074_), .B0(new_n3073_), .Y(new_n10195_));
  OAI21X1  g07759(.A0(new_n10194_), .A1(new_n10193_), .B0(new_n10195_), .Y(new_n10196_));
  OR3X1    g07760(.A(new_n2985_), .B(new_n2536_), .C(new_n5084_), .Y(new_n10197_));
  OR4X1    g07761(.A(new_n5082_), .B(new_n5922_), .C(new_n5237_), .D(pi0122), .Y(new_n10198_));
  OAI21X1  g07762(.A0(new_n10198_), .A1(new_n10197_), .B0(new_n10187_), .Y(new_n10199_));
  AOI22X1  g07763(.A0(new_n10199_), .A1(new_n10186_), .B0(new_n5960_), .B1(pi0120), .Y(new_n10200_));
  OR3X1    g07764(.A(new_n5920_), .B(new_n2793_), .C(pi0039), .Y(new_n10201_));
  OAI21X1  g07765(.A0(new_n10201_), .A1(new_n10200_), .B0(pi0100), .Y(new_n10202_));
  AOI22X1  g07766(.A0(new_n10202_), .A1(new_n2979_), .B0(new_n10177_), .B1(new_n10090_), .Y(new_n10203_));
  AOI21X1  g07767(.A0(new_n10177_), .A1(new_n6265_), .B0(pi0299), .Y(new_n10204_));
  OR2X1    g07768(.A(new_n10177_), .B(new_n6377_), .Y(new_n10205_));
  NOR2X1   g07769(.A(new_n10177_), .B(new_n6375_), .Y(new_n10206_));
  AOI21X1  g07770(.A0(new_n10206_), .A1(new_n5041_), .B0(new_n6265_), .Y(new_n10207_));
  OAI21X1  g07771(.A0(new_n10205_), .A1(new_n5041_), .B0(new_n10207_), .Y(new_n10208_));
  AOI21X1  g07772(.A0(new_n10177_), .A1(new_n6271_), .B0(new_n2933_), .Y(new_n10209_));
  AOI21X1  g07773(.A0(new_n10206_), .A1(new_n5058_), .B0(new_n6271_), .Y(new_n10210_));
  OAI21X1  g07774(.A0(new_n10205_), .A1(new_n5058_), .B0(new_n10210_), .Y(new_n10211_));
  AOI22X1  g07775(.A0(new_n10211_), .A1(new_n10209_), .B0(new_n10208_), .B1(new_n10204_), .Y(new_n10212_));
  INVX1    g07776(.A(new_n5926_), .Y(new_n10213_));
  AND2X1   g07777(.A(new_n10176_), .B(pi1093), .Y(new_n10214_));
  INVX1    g07778(.A(new_n10214_), .Y(new_n10215_));
  NOR4X1   g07779(.A(new_n2561_), .B(new_n2567_), .C(new_n5893_), .D(pi0088), .Y(new_n10216_));
  OAI21X1  g07780(.A0(new_n10216_), .A1(pi0097), .B0(new_n2731_), .Y(new_n10217_));
  OR4X1    g07781(.A(new_n10217_), .B(new_n2565_), .C(pi0110), .D(pi0108), .Y(new_n10218_));
  AOI21X1  g07782(.A0(new_n10218_), .A1(new_n5931_), .B0(new_n2502_), .Y(new_n10219_));
  OAI21X1  g07783(.A0(new_n10219_), .A1(new_n5888_), .B0(new_n5885_), .Y(new_n10220_));
  AOI21X1  g07784(.A0(new_n10220_), .A1(new_n2534_), .B0(new_n2847_), .Y(new_n10221_));
  NOR4X1   g07785(.A(new_n5905_), .B(new_n7619_), .C(new_n5084_), .D(pi0072), .Y(new_n10222_));
  OAI21X1  g07786(.A0(new_n10221_), .A1(pi0096), .B0(new_n10222_), .Y(new_n10223_));
  AND3X1   g07787(.A(new_n10176_), .B(pi0829), .C(new_n5906_), .Y(new_n10224_));
  NAND4X1  g07788(.A(new_n10216_), .B(new_n5885_), .C(new_n2497_), .D(new_n2682_), .Y(new_n10225_));
  OR4X1    g07789(.A(new_n5881_), .B(new_n2847_), .C(new_n5084_), .D(pi0096), .Y(new_n10226_));
  AOI21X1  g07790(.A0(new_n10225_), .A1(new_n5889_), .B0(new_n10226_), .Y(new_n10227_));
  NAND3X1  g07791(.A(pi1092), .B(pi0982), .C(pi0951), .Y(new_n10228_));
  AOI21X1  g07792(.A0(new_n10227_), .A1(pi0824), .B0(new_n10228_), .Y(new_n10229_));
  NAND2X1  g07793(.A(new_n10229_), .B(new_n5237_), .Y(new_n10230_));
  NAND3X1  g07794(.A(pi0982), .B(pi0951), .C(pi0122), .Y(new_n10231_));
  OR3X1    g07795(.A(new_n10231_), .B(new_n5024_), .C(new_n5237_), .Y(new_n10232_));
  OAI21X1  g07796(.A0(new_n10232_), .A1(new_n10227_), .B0(new_n10230_), .Y(new_n10233_));
  AOI21X1  g07797(.A0(new_n10224_), .A1(new_n10223_), .B0(new_n10233_), .Y(new_n10234_));
  OAI22X1  g07798(.A0(new_n10234_), .A1(new_n10213_), .B0(new_n10215_), .B1(new_n8194_), .Y(new_n10235_));
  INVX1    g07799(.A(new_n10185_), .Y(new_n10236_));
  AND2X1   g07800(.A(new_n10227_), .B(pi0824), .Y(new_n10237_));
  OAI21X1  g07801(.A0(new_n10237_), .A1(new_n10236_), .B0(new_n10082_), .Y(new_n10238_));
  AOI21X1  g07802(.A0(new_n10235_), .A1(pi1091), .B0(new_n10238_), .Y(new_n10239_));
  AND3X1   g07803(.A(new_n5909_), .B(new_n5902_), .C(new_n5032_), .Y(new_n10240_));
  OR2X1    g07804(.A(new_n10147_), .B(new_n10240_), .Y(new_n10241_));
  OAI21X1  g07805(.A0(new_n10241_), .A1(new_n10082_), .B0(new_n2939_), .Y(new_n10242_));
  OAI22X1  g07806(.A0(new_n10242_), .A1(new_n10239_), .B0(new_n10212_), .B1(new_n2939_), .Y(new_n10243_));
  AOI21X1  g07807(.A0(new_n10243_), .A1(new_n3251_), .B0(new_n10203_), .Y(new_n10244_));
  AOI21X1  g07808(.A0(new_n10177_), .A1(new_n3132_), .B0(new_n3131_), .Y(new_n10245_));
  OAI22X1  g07809(.A0(new_n2758_), .A1(pi0833), .B0(pi0829), .B1(pi0824), .Y(new_n10246_));
  OAI21X1  g07810(.A0(new_n10246_), .A1(new_n10197_), .B0(new_n10187_), .Y(new_n10247_));
  OAI21X1  g07811(.A0(new_n10197_), .A1(new_n8199_), .B0(new_n10185_), .Y(new_n10248_));
  AOI21X1  g07812(.A0(new_n10248_), .A1(new_n10247_), .B0(pi0120), .Y(new_n10249_));
  MX2X1    g07813(.A(new_n5966_), .B(new_n5971_), .S0(new_n5968_), .Y(new_n10250_));
  OAI21X1  g07814(.A0(new_n10250_), .A1(new_n10082_), .B0(new_n3064_), .Y(new_n10251_));
  OAI21X1  g07815(.A0(new_n10251_), .A1(new_n10249_), .B0(new_n10245_), .Y(new_n10252_));
  AND2X1   g07816(.A(new_n10252_), .B(new_n3073_), .Y(new_n10253_));
  OAI21X1  g07817(.A0(new_n10244_), .A1(pi0087), .B0(new_n10253_), .Y(new_n10254_));
  AOI21X1  g07818(.A0(new_n10254_), .A1(new_n10196_), .B0(new_n6295_), .Y(new_n10255_));
  NOR2X1   g07819(.A(new_n10084_), .B(new_n5960_), .Y(new_n10256_));
  NOR4X1   g07820(.A(new_n10228_), .B(new_n10092_), .C(new_n5032_), .D(pi1091), .Y(new_n10257_));
  INVX1    g07821(.A(new_n10257_), .Y(new_n10258_));
  AOI21X1  g07822(.A0(new_n10258_), .A1(new_n10199_), .B0(pi0120), .Y(new_n10259_));
  OAI21X1  g07823(.A0(new_n10259_), .A1(new_n10256_), .B0(new_n6278_), .Y(new_n10260_));
  NOR2X1   g07824(.A(new_n10177_), .B(new_n10094_), .Y(new_n10261_));
  AOI21X1  g07825(.A0(new_n10261_), .A1(new_n7692_), .B0(new_n3060_), .Y(new_n10262_));
  OAI21X1  g07826(.A0(new_n10261_), .A1(new_n3047_), .B0(pi0100), .Y(new_n10263_));
  AOI21X1  g07827(.A0(new_n10262_), .A1(new_n10260_), .B0(new_n10263_), .Y(new_n10264_));
  OR3X1    g07828(.A(new_n10105_), .B(new_n10240_), .C(new_n10082_), .Y(new_n10265_));
  NAND2X1  g07829(.A(new_n10235_), .B(pi1091), .Y(new_n10266_));
  OR4X1    g07830(.A(new_n10237_), .B(new_n10228_), .C(new_n10092_), .D(new_n5968_), .Y(new_n10267_));
  NAND3X1  g07831(.A(new_n10267_), .B(new_n10266_), .C(new_n10082_), .Y(new_n10268_));
  AOI21X1  g07832(.A0(new_n10268_), .A1(new_n10265_), .B0(pi0039), .Y(new_n10269_));
  OR3X1    g07833(.A(new_n10228_), .B(new_n10108_), .C(new_n10098_), .Y(new_n10270_));
  AND2X1   g07834(.A(new_n10270_), .B(new_n10258_), .Y(new_n10271_));
  OAI22X1  g07835(.A0(new_n10271_), .A1(pi0120), .B0(new_n10084_), .B1(new_n7192_), .Y(new_n10272_));
  MX2X1    g07836(.A(new_n10272_), .B(new_n10261_), .S0(new_n6256_), .Y(new_n10273_));
  AND2X1   g07837(.A(new_n10273_), .B(new_n5041_), .Y(new_n10274_));
  NOR3X1   g07838(.A(new_n10177_), .B(new_n10094_), .C(new_n5044_), .Y(new_n10275_));
  AOI21X1  g07839(.A0(new_n10272_), .A1(new_n5044_), .B0(new_n10275_), .Y(new_n10276_));
  OAI21X1  g07840(.A0(new_n10276_), .A1(new_n5041_), .B0(new_n6264_), .Y(new_n10277_));
  AND2X1   g07841(.A(new_n10204_), .B(new_n10119_), .Y(new_n10278_));
  OAI21X1  g07842(.A0(new_n10277_), .A1(new_n10274_), .B0(new_n10278_), .Y(new_n10279_));
  AND2X1   g07843(.A(new_n10273_), .B(new_n5058_), .Y(new_n10280_));
  OAI21X1  g07844(.A0(new_n10276_), .A1(new_n5058_), .B0(new_n6270_), .Y(new_n10281_));
  NAND2X1  g07845(.A(new_n6271_), .B(new_n10077_), .Y(new_n10282_));
  AND2X1   g07846(.A(new_n10282_), .B(new_n10209_), .Y(new_n10283_));
  OAI21X1  g07847(.A0(new_n10281_), .A1(new_n10280_), .B0(new_n10283_), .Y(new_n10284_));
  AND3X1   g07848(.A(new_n10284_), .B(new_n10279_), .C(pi0039), .Y(new_n10285_));
  OAI21X1  g07849(.A0(new_n10285_), .A1(new_n10269_), .B0(new_n2979_), .Y(new_n10286_));
  OAI21X1  g07850(.A0(new_n10177_), .A1(new_n10094_), .B0(pi0038), .Y(new_n10287_));
  AND2X1   g07851(.A(new_n10287_), .B(new_n3007_), .Y(new_n10288_));
  AOI21X1  g07852(.A0(new_n10288_), .A1(new_n10286_), .B0(new_n10264_), .Y(new_n10289_));
  NAND2X1  g07853(.A(new_n10258_), .B(new_n10247_), .Y(new_n10290_));
  AOI22X1  g07854(.A0(new_n10290_), .A1(new_n10249_), .B0(new_n10251_), .B1(new_n10132_), .Y(new_n10291_));
  NAND2X1  g07855(.A(new_n10245_), .B(new_n10133_), .Y(new_n10292_));
  OAI22X1  g07856(.A0(new_n10292_), .A1(new_n10291_), .B0(new_n10289_), .B1(pi0087), .Y(new_n10293_));
  AOI21X1  g07857(.A0(new_n10258_), .A1(new_n10191_), .B0(pi0120), .Y(new_n10294_));
  OAI22X1  g07858(.A0(new_n10294_), .A1(new_n10140_), .B0(new_n10261_), .B1(new_n9672_), .Y(new_n10295_));
  OAI21X1  g07859(.A0(new_n10261_), .A1(new_n3070_), .B0(pi0075), .Y(new_n10296_));
  AOI21X1  g07860(.A0(new_n10295_), .A1(new_n3070_), .B0(new_n10296_), .Y(new_n10297_));
  OR2X1    g07861(.A(new_n10297_), .B(new_n6295_), .Y(new_n10298_));
  AOI21X1  g07862(.A0(new_n10293_), .A1(new_n3073_), .B0(new_n10298_), .Y(new_n10299_));
  OAI22X1  g07863(.A0(new_n10299_), .A1(new_n10183_), .B0(new_n10255_), .B1(new_n6073_), .Y(new_n10300_));
  NOR3X1   g07864(.A(new_n10214_), .B(new_n5880_), .C(pi0120), .Y(new_n10301_));
  NOR3X1   g07865(.A(new_n10301_), .B(new_n10180_), .C(new_n8943_), .Y(new_n10302_));
  INVX1    g07866(.A(new_n10078_), .Y(new_n10303_));
  OAI21X1  g07867(.A0(new_n10105_), .A1(new_n10240_), .B0(new_n2939_), .Y(new_n10304_));
  MX2X1    g07868(.A(new_n6246_), .B(new_n5947_), .S0(pi1091), .Y(new_n10305_));
  OR2X1    g07869(.A(new_n10077_), .B(new_n6255_), .Y(new_n10306_));
  OAI21X1  g07870(.A0(new_n10305_), .A1(new_n6256_), .B0(new_n10306_), .Y(new_n10307_));
  MX2X1    g07871(.A(new_n10305_), .B(new_n10077_), .S0(new_n5043_), .Y(new_n10308_));
  OAI21X1  g07872(.A0(new_n10308_), .A1(new_n5041_), .B0(new_n6264_), .Y(new_n10309_));
  AOI21X1  g07873(.A0(new_n10307_), .A1(new_n5041_), .B0(new_n10309_), .Y(new_n10310_));
  OAI21X1  g07874(.A0(new_n6264_), .A1(new_n10124_), .B0(new_n2933_), .Y(new_n10311_));
  OAI21X1  g07875(.A0(new_n10308_), .A1(new_n5058_), .B0(new_n6270_), .Y(new_n10312_));
  AOI21X1  g07876(.A0(new_n10307_), .A1(new_n5058_), .B0(new_n10312_), .Y(new_n10313_));
  NAND2X1  g07877(.A(new_n10282_), .B(pi0299), .Y(new_n10314_));
  OAI22X1  g07878(.A0(new_n10314_), .A1(new_n10313_), .B0(new_n10311_), .B1(new_n10310_), .Y(new_n10315_));
  AOI21X1  g07879(.A0(new_n10315_), .A1(pi0039), .B0(pi0038), .Y(new_n10316_));
  NAND2X1  g07880(.A(new_n10316_), .B(new_n10304_), .Y(new_n10317_));
  AOI21X1  g07881(.A0(new_n10077_), .A1(pi0038), .B0(pi0100), .Y(new_n10318_));
  AOI22X1  g07882(.A0(new_n10318_), .A1(new_n10317_), .B0(new_n10124_), .B1(new_n5963_), .Y(new_n10319_));
  OAI21X1  g07883(.A0(new_n10319_), .A1(pi0087), .B0(new_n10134_), .Y(new_n10320_));
  OAI21X1  g07884(.A0(new_n10124_), .A1(new_n5921_), .B0(pi0075), .Y(new_n10321_));
  AOI21X1  g07885(.A0(new_n10139_), .A1(new_n5921_), .B0(new_n10321_), .Y(new_n10322_));
  AOI21X1  g07886(.A0(new_n10320_), .A1(new_n3073_), .B0(new_n10322_), .Y(new_n10323_));
  AOI21X1  g07887(.A0(new_n10241_), .A1(new_n2939_), .B0(new_n5954_), .Y(new_n10324_));
  OAI21X1  g07888(.A0(new_n10324_), .A1(pi0100), .B0(new_n5964_), .Y(new_n10325_));
  AOI21X1  g07889(.A0(new_n10325_), .A1(new_n3131_), .B0(new_n5974_), .Y(new_n10326_));
  OAI21X1  g07890(.A0(new_n10326_), .A1(pi0075), .B0(new_n10165_), .Y(new_n10327_));
  AOI21X1  g07891(.A0(new_n6295_), .A1(new_n10082_), .B0(new_n6073_), .Y(new_n10328_));
  AOI22X1  g07892(.A0(new_n10328_), .A1(new_n10327_), .B0(new_n10170_), .B1(new_n6295_), .Y(new_n10329_));
  OAI21X1  g07893(.A0(new_n10323_), .A1(new_n10303_), .B0(new_n10329_), .Y(new_n10330_));
  AND2X1   g07894(.A(new_n10175_), .B(pi0120), .Y(new_n10331_));
  AOI22X1  g07895(.A0(new_n10331_), .A1(new_n10330_), .B0(new_n10302_), .B1(new_n10300_), .Y(new_n10332_));
  OAI21X1  g07896(.A0(new_n10332_), .A1(new_n10075_), .B0(new_n10182_), .Y(po0278));
  OR4X1    g07897(.A(pi0136), .B(pi0135), .C(pi0134), .D(pi0130), .Y(new_n10334_));
  NOR4X1   g07898(.A(new_n10334_), .B(pi0132), .C(pi0126), .D(pi0121), .Y(new_n10335_));
  INVX1    g07899(.A(new_n10335_), .Y(new_n10336_));
  NOR2X1   g07900(.A(pi0133), .B(pi0125), .Y(new_n10337_));
  XOR2X1   g07901(.A(new_n10337_), .B(pi0121), .Y(new_n10338_));
  AND2X1   g07902(.A(new_n10338_), .B(new_n10336_), .Y(new_n10339_));
  NOR4X1   g07903(.A(pi0084), .B(pi0071), .C(pi0068), .D(pi0067), .Y(new_n10340_));
  AND2X1   g07904(.A(new_n10340_), .B(new_n2534_), .Y(new_n10341_));
  INVX1    g07905(.A(new_n10341_), .Y(new_n10342_));
  OR3X1    g07906(.A(new_n10342_), .B(new_n10339_), .C(pi0087), .Y(new_n10343_));
  NAND3X1  g07907(.A(new_n5023_), .B(new_n2776_), .C(pi0051), .Y(new_n10344_));
  AND2X1   g07908(.A(new_n10344_), .B(pi0161), .Y(new_n10345_));
  AND2X1   g07909(.A(pi0146), .B(pi0051), .Y(new_n10346_));
  NOR4X1   g07910(.A(new_n10346_), .B(new_n10345_), .C(new_n10341_), .D(new_n5048_), .Y(new_n10347_));
  AOI21X1  g07911(.A0(new_n5023_), .A1(pi0163), .B0(new_n3131_), .Y(new_n10348_));
  NOR2X1   g07912(.A(new_n10348_), .B(new_n5215_), .Y(new_n10349_));
  OAI21X1  g07913(.A0(new_n10347_), .A1(pi0087), .B0(new_n10349_), .Y(new_n10350_));
  NAND3X1  g07914(.A(new_n10350_), .B(new_n10343_), .C(po1038), .Y(new_n10351_));
  AND3X1   g07915(.A(new_n5023_), .B(new_n2953_), .C(pi0051), .Y(new_n10352_));
  INVX1    g07916(.A(new_n10352_), .Y(new_n10353_));
  NOR2X1   g07917(.A(new_n10341_), .B(new_n5048_), .Y(new_n10354_));
  OAI21X1  g07918(.A0(new_n2953_), .A1(new_n2534_), .B0(new_n10354_), .Y(new_n10355_));
  AOI21X1  g07919(.A0(new_n10353_), .A1(pi0144), .B0(new_n10355_), .Y(new_n10356_));
  NOR2X1   g07920(.A(new_n10356_), .B(pi0299), .Y(new_n10357_));
  NOR2X1   g07921(.A(new_n10347_), .B(new_n2933_), .Y(new_n10358_));
  NOR3X1   g07922(.A(new_n10358_), .B(new_n10357_), .C(new_n5215_), .Y(new_n10359_));
  INVX1    g07923(.A(new_n10359_), .Y(new_n10360_));
  AOI21X1  g07924(.A0(new_n10360_), .A1(pi0038), .B0(pi0100), .Y(new_n10361_));
  AOI21X1  g07925(.A0(new_n10342_), .A1(pi0038), .B0(pi0100), .Y(new_n10362_));
  INVX1    g07926(.A(new_n2560_), .Y(new_n10363_));
  OR3X1    g07927(.A(new_n7601_), .B(new_n2460_), .C(pi0069), .Y(new_n10364_));
  OR4X1    g07928(.A(new_n10364_), .B(new_n2604_), .C(new_n10363_), .D(new_n2465_), .Y(new_n10365_));
  AND3X1   g07929(.A(new_n5897_), .B(new_n2513_), .C(new_n2535_), .Y(new_n10366_));
  NAND4X1  g07930(.A(new_n10366_), .B(new_n2496_), .C(new_n2489_), .D(new_n2494_), .Y(new_n10367_));
  NOR4X1   g07931(.A(new_n10367_), .B(new_n10365_), .C(new_n7619_), .D(new_n2530_), .Y(new_n10368_));
  INVX1    g07932(.A(new_n10366_), .Y(new_n10369_));
  AOI21X1  g07933(.A0(new_n10369_), .A1(new_n10340_), .B0(pi0051), .Y(new_n10370_));
  INVX1    g07934(.A(new_n10370_), .Y(new_n10371_));
  OR3X1    g07935(.A(new_n2472_), .B(new_n2576_), .C(pi0050), .Y(new_n10372_));
  OR4X1    g07936(.A(new_n10372_), .B(new_n10364_), .C(new_n2604_), .D(new_n2465_), .Y(new_n10373_));
  OAI21X1  g07937(.A0(new_n10365_), .A1(new_n2566_), .B0(new_n10373_), .Y(new_n10374_));
  NAND3X1  g07938(.A(new_n6737_), .B(pi0086), .C(new_n5777_), .Y(new_n10375_));
  OAI21X1  g07939(.A0(new_n10375_), .A1(new_n10365_), .B0(new_n10340_), .Y(new_n10376_));
  AOI21X1  g07940(.A0(new_n10374_), .A1(new_n8227_), .B0(new_n10376_), .Y(new_n10377_));
  NOR3X1   g07941(.A(new_n10377_), .B(new_n10371_), .C(new_n5881_), .Y(new_n10378_));
  NAND3X1  g07942(.A(new_n10366_), .B(pi0314), .C(new_n5777_), .Y(new_n10379_));
  NOR4X1   g07943(.A(new_n10379_), .B(new_n10373_), .C(new_n6738_), .D(new_n5881_), .Y(new_n10380_));
  NOR2X1   g07944(.A(new_n10380_), .B(new_n10342_), .Y(new_n10381_));
  INVX1    g07945(.A(new_n10381_), .Y(new_n10382_));
  NOR2X1   g07946(.A(new_n10382_), .B(new_n10378_), .Y(new_n10383_));
  NOR2X1   g07947(.A(new_n10383_), .B(new_n5023_), .Y(new_n10384_));
  OR3X1    g07948(.A(new_n10384_), .B(new_n10368_), .C(new_n10354_), .Y(new_n10385_));
  NOR4X1   g07949(.A(new_n10380_), .B(new_n10378_), .C(new_n10368_), .D(new_n10342_), .Y(new_n10386_));
  AND2X1   g07950(.A(new_n5023_), .B(pi0051), .Y(new_n10387_));
  AOI21X1  g07951(.A0(new_n8143_), .A1(pi0072), .B0(new_n10387_), .Y(new_n10388_));
  MX2X1    g07952(.A(new_n10388_), .B(new_n10386_), .S0(new_n5048_), .Y(new_n10389_));
  INVX1    g07953(.A(new_n10389_), .Y(new_n10390_));
  MX2X1    g07954(.A(new_n10390_), .B(new_n10385_), .S0(pi0144), .Y(new_n10391_));
  AOI21X1  g07955(.A0(new_n10391_), .A1(new_n10353_), .B0(new_n5203_), .Y(new_n10392_));
  INVX1    g07956(.A(new_n9695_), .Y(new_n10393_));
  AND2X1   g07957(.A(new_n5023_), .B(new_n2984_), .Y(new_n10394_));
  INVX1    g07958(.A(new_n10394_), .Y(new_n10395_));
  NOR4X1   g07959(.A(new_n10395_), .B(new_n10379_), .C(new_n10393_), .D(pi0051), .Y(new_n10396_));
  INVX1    g07960(.A(new_n10396_), .Y(new_n10397_));
  NAND3X1  g07961(.A(new_n10397_), .B(new_n10389_), .C(pi0142), .Y(new_n10398_));
  AND2X1   g07962(.A(new_n10386_), .B(new_n5048_), .Y(new_n10399_));
  NOR3X1   g07963(.A(new_n10379_), .B(new_n10393_), .C(pi0051), .Y(new_n10400_));
  OAI21X1  g07964(.A0(new_n10400_), .A1(pi0072), .B0(new_n5169_), .Y(new_n10401_));
  AOI21X1  g07965(.A0(new_n10401_), .A1(new_n5023_), .B0(new_n10399_), .Y(new_n10402_));
  OR2X1    g07966(.A(new_n10402_), .B(pi0142), .Y(new_n10403_));
  AND3X1   g07967(.A(new_n10403_), .B(new_n10398_), .C(new_n7344_), .Y(new_n10404_));
  OR2X1    g07968(.A(new_n10352_), .B(new_n7344_), .Y(new_n10405_));
  NOR4X1   g07969(.A(new_n10384_), .B(new_n10380_), .C(new_n10368_), .D(new_n10354_), .Y(new_n10406_));
  OAI21X1  g07970(.A0(new_n10406_), .A1(new_n10405_), .B0(new_n5203_), .Y(new_n10407_));
  OAI21X1  g07971(.A0(new_n10407_), .A1(new_n10404_), .B0(pi0179), .Y(new_n10408_));
  OR2X1    g07972(.A(new_n10408_), .B(new_n10392_), .Y(new_n10409_));
  NOR2X1   g07973(.A(new_n10386_), .B(new_n5023_), .Y(new_n10410_));
  AND2X1   g07974(.A(new_n8143_), .B(pi0072), .Y(new_n10411_));
  INVX1    g07975(.A(new_n10411_), .Y(new_n10412_));
  MX2X1    g07976(.A(new_n8618_), .B(new_n8616_), .S0(pi0024), .Y(new_n10413_));
  MX2X1    g07977(.A(new_n10413_), .B(new_n8616_), .S0(pi0314), .Y(new_n10414_));
  NOR2X1   g07978(.A(new_n6773_), .B(new_n5898_), .Y(new_n10415_));
  AOI21X1  g07979(.A0(new_n10415_), .A1(new_n10414_), .B0(pi0051), .Y(new_n10416_));
  AOI21X1  g07980(.A0(new_n10416_), .A1(new_n10412_), .B0(new_n5048_), .Y(new_n10417_));
  NOR2X1   g07981(.A(new_n10417_), .B(new_n10410_), .Y(new_n10418_));
  INVX1    g07982(.A(new_n10386_), .Y(new_n10419_));
  AOI21X1  g07983(.A0(new_n10414_), .A1(new_n2479_), .B0(pi0072), .Y(new_n10420_));
  NOR2X1   g07984(.A(new_n10420_), .B(new_n5170_), .Y(new_n10421_));
  MX2X1    g07985(.A(new_n10421_), .B(new_n10419_), .S0(new_n5048_), .Y(new_n10422_));
  OAI21X1  g07986(.A0(new_n10422_), .A1(pi0142), .B0(new_n7344_), .Y(new_n10423_));
  AOI21X1  g07987(.A0(new_n10418_), .A1(pi0142), .B0(new_n10423_), .Y(new_n10424_));
  OAI21X1  g07988(.A0(new_n10386_), .A1(new_n10405_), .B0(new_n5203_), .Y(new_n10425_));
  AOI21X1  g07989(.A0(new_n10413_), .A1(new_n2479_), .B0(pi0072), .Y(new_n10426_));
  NOR2X1   g07990(.A(new_n10426_), .B(new_n5170_), .Y(new_n10427_));
  MX2X1    g07991(.A(new_n10427_), .B(new_n10419_), .S0(new_n5048_), .Y(new_n10428_));
  NOR2X1   g07992(.A(new_n10388_), .B(new_n5048_), .Y(new_n10429_));
  AND3X1   g07993(.A(new_n10413_), .B(new_n10394_), .C(new_n2479_), .Y(new_n10430_));
  NOR3X1   g07994(.A(new_n10430_), .B(new_n10429_), .C(new_n10410_), .Y(new_n10431_));
  AOI21X1  g07995(.A0(new_n10431_), .A1(pi0142), .B0(pi0144), .Y(new_n10432_));
  OAI21X1  g07996(.A0(new_n10428_), .A1(pi0142), .B0(new_n10432_), .Y(new_n10433_));
  MX2X1    g07997(.A(new_n10383_), .B(new_n10341_), .S0(new_n5023_), .Y(new_n10434_));
  NOR3X1   g07998(.A(new_n10378_), .B(new_n10368_), .C(new_n10342_), .Y(new_n10435_));
  NOR3X1   g07999(.A(pi0468), .B(pi0332), .C(pi0051), .Y(new_n10436_));
  INVX1    g08000(.A(new_n10436_), .Y(new_n10437_));
  NOR2X1   g08001(.A(new_n10437_), .B(new_n10435_), .Y(new_n10438_));
  NOR2X1   g08002(.A(new_n10438_), .B(new_n10410_), .Y(new_n10439_));
  OR2X1    g08003(.A(new_n10378_), .B(new_n10342_), .Y(new_n10440_));
  AND2X1   g08004(.A(new_n10440_), .B(new_n5023_), .Y(new_n10441_));
  NOR4X1   g08005(.A(new_n10340_), .B(pi0468), .C(pi0332), .D(pi0051), .Y(new_n10442_));
  OAI21X1  g08006(.A0(new_n10377_), .A1(new_n10371_), .B0(new_n2984_), .Y(new_n10443_));
  OAI21X1  g08007(.A0(new_n10442_), .A1(new_n10394_), .B0(new_n10443_), .Y(new_n10444_));
  INVX1    g08008(.A(new_n10444_), .Y(new_n10445_));
  MX2X1    g08009(.A(new_n10445_), .B(new_n10441_), .S0(new_n2953_), .Y(new_n10446_));
  OAI21X1  g08010(.A0(new_n10446_), .A1(new_n10434_), .B0(new_n10439_), .Y(new_n10447_));
  AOI21X1  g08011(.A0(new_n10447_), .A1(pi0144), .B0(new_n5203_), .Y(new_n10448_));
  AOI21X1  g08012(.A0(new_n10448_), .A1(new_n10433_), .B0(pi0179), .Y(new_n10449_));
  OAI21X1  g08013(.A0(new_n10425_), .A1(new_n10424_), .B0(new_n10449_), .Y(new_n10450_));
  AOI21X1  g08014(.A0(new_n10450_), .A1(new_n10409_), .B0(pi0299), .Y(new_n10451_));
  AND2X1   g08015(.A(new_n10344_), .B(new_n4611_), .Y(new_n10452_));
  INVX1    g08016(.A(new_n10452_), .Y(new_n10453_));
  NOR4X1   g08017(.A(new_n10384_), .B(new_n10368_), .C(new_n10354_), .D(new_n2776_), .Y(new_n10454_));
  INVX1    g08018(.A(new_n10340_), .Y(new_n10455_));
  OAI21X1  g08019(.A0(new_n10368_), .A1(new_n10455_), .B0(new_n10436_), .Y(new_n10456_));
  NAND2X1  g08020(.A(new_n10456_), .B(new_n2776_), .Y(new_n10457_));
  OAI21X1  g08021(.A0(new_n10457_), .A1(new_n10410_), .B0(pi0161), .Y(new_n10458_));
  OAI22X1  g08022(.A0(new_n10458_), .A1(new_n10454_), .B0(new_n10453_), .B1(new_n10389_), .Y(new_n10459_));
  AND3X1   g08023(.A(new_n10397_), .B(new_n10389_), .C(pi0146), .Y(new_n10460_));
  OAI21X1  g08024(.A0(new_n10402_), .A1(pi0146), .B0(new_n4611_), .Y(new_n10461_));
  INVX1    g08025(.A(new_n10387_), .Y(new_n10462_));
  OR4X1    g08026(.A(new_n10437_), .B(new_n10380_), .C(new_n10368_), .D(new_n10455_), .Y(new_n10463_));
  AOI22X1  g08027(.A0(new_n10463_), .A1(new_n10462_), .B0(new_n10342_), .B1(pi0146), .Y(new_n10464_));
  OR2X1    g08028(.A(new_n10464_), .B(new_n4611_), .Y(new_n10465_));
  OAI22X1  g08029(.A0(new_n10465_), .A1(new_n10399_), .B0(new_n10461_), .B1(new_n10460_), .Y(new_n10466_));
  AOI22X1  g08030(.A0(new_n10466_), .A1(new_n7095_), .B0(new_n10459_), .B1(new_n7059_), .Y(new_n10467_));
  AOI21X1  g08031(.A0(new_n10418_), .A1(pi0146), .B0(new_n7096_), .Y(new_n10468_));
  OAI21X1  g08032(.A0(new_n10422_), .A1(pi0146), .B0(new_n10468_), .Y(new_n10469_));
  AOI21X1  g08033(.A0(new_n10431_), .A1(pi0146), .B0(new_n7060_), .Y(new_n10470_));
  OAI21X1  g08034(.A0(new_n10428_), .A1(pi0146), .B0(new_n10470_), .Y(new_n10471_));
  AND3X1   g08035(.A(new_n10471_), .B(new_n10469_), .C(new_n4611_), .Y(new_n10472_));
  MX2X1    g08036(.A(new_n10445_), .B(new_n10441_), .S0(new_n2776_), .Y(new_n10473_));
  OAI21X1  g08037(.A0(new_n10473_), .A1(new_n10434_), .B0(new_n10439_), .Y(new_n10474_));
  NAND2X1  g08038(.A(new_n10344_), .B(new_n7095_), .Y(new_n10475_));
  OAI21X1  g08039(.A0(new_n10475_), .A1(new_n10386_), .B0(pi0161), .Y(new_n10476_));
  AOI21X1  g08040(.A0(new_n10474_), .A1(new_n7059_), .B0(new_n10476_), .Y(new_n10477_));
  OR2X1    g08041(.A(new_n10477_), .B(pi0156), .Y(new_n10478_));
  OAI22X1  g08042(.A0(new_n10478_), .A1(new_n10472_), .B0(new_n10467_), .B1(new_n8789_), .Y(new_n10479_));
  OAI21X1  g08043(.A0(new_n10479_), .A1(new_n10451_), .B0(new_n7259_), .Y(new_n10480_));
  NOR3X1   g08044(.A(new_n10367_), .B(new_n10365_), .C(new_n5881_), .Y(new_n10481_));
  NOR2X1   g08045(.A(new_n10481_), .B(new_n10342_), .Y(new_n10482_));
  INVX1    g08046(.A(new_n10482_), .Y(new_n10483_));
  AOI21X1  g08047(.A0(new_n10483_), .A1(new_n5048_), .B0(new_n5037_), .Y(new_n10484_));
  NOR3X1   g08048(.A(new_n5881_), .B(new_n2536_), .C(pi0096), .Y(new_n10485_));
  NOR2X1   g08049(.A(new_n10485_), .B(pi0051), .Y(new_n10486_));
  MX2X1    g08050(.A(new_n10486_), .B(new_n10482_), .S0(new_n5048_), .Y(new_n10487_));
  INVX1    g08051(.A(new_n10487_), .Y(new_n10488_));
  AOI21X1  g08052(.A0(new_n10488_), .A1(pi0142), .B0(new_n5248_), .Y(new_n10489_));
  OAI21X1  g08053(.A0(new_n10484_), .A1(pi0142), .B0(new_n10489_), .Y(new_n10490_));
  AND2X1   g08054(.A(new_n10490_), .B(new_n7203_), .Y(new_n10491_));
  NOR3X1   g08055(.A(pi0468), .B(pi0332), .C(pi0287), .Y(new_n10492_));
  AOI21X1  g08056(.A0(new_n10492_), .A1(new_n2534_), .B0(new_n10487_), .Y(new_n10493_));
  AND3X1   g08057(.A(new_n10493_), .B(new_n10353_), .C(pi0224), .Y(new_n10494_));
  AOI21X1  g08058(.A0(new_n10353_), .A1(new_n10342_), .B0(new_n5247_), .Y(new_n10495_));
  NOR4X1   g08059(.A(new_n10340_), .B(new_n5247_), .C(new_n5048_), .D(pi0051), .Y(new_n10496_));
  NOR3X1   g08060(.A(new_n10496_), .B(new_n10495_), .C(pi0144), .Y(new_n10497_));
  OAI21X1  g08061(.A0(new_n10494_), .A1(new_n10491_), .B0(new_n10497_), .Y(new_n10498_));
  INVX1    g08062(.A(new_n10442_), .Y(new_n10499_));
  INVX1    g08063(.A(new_n10492_), .Y(new_n10500_));
  NOR2X1   g08064(.A(new_n10482_), .B(pi0051), .Y(new_n10501_));
  INVX1    g08065(.A(new_n10501_), .Y(new_n10502_));
  AOI22X1  g08066(.A0(new_n10502_), .A1(new_n7795_), .B0(new_n10500_), .B1(new_n10499_), .Y(new_n10503_));
  INVX1    g08067(.A(new_n10503_), .Y(new_n10504_));
  AOI21X1  g08068(.A0(new_n10504_), .A1(new_n10355_), .B0(new_n7203_), .Y(new_n10505_));
  NAND2X1  g08069(.A(new_n10505_), .B(new_n10340_), .Y(new_n10506_));
  OR2X1    g08070(.A(new_n10495_), .B(new_n7344_), .Y(new_n10507_));
  MX2X1    g08071(.A(new_n10482_), .B(new_n5023_), .S0(pi0051), .Y(new_n10508_));
  AOI21X1  g08072(.A0(pi0142), .A1(pi0051), .B0(new_n5248_), .Y(new_n10509_));
  AOI21X1  g08073(.A0(new_n10509_), .A1(new_n10508_), .B0(new_n10507_), .Y(new_n10510_));
  AOI21X1  g08074(.A0(new_n10510_), .A1(new_n10506_), .B0(new_n5204_), .Y(new_n10511_));
  OR2X1    g08075(.A(new_n10510_), .B(pi0181), .Y(new_n10512_));
  AOI21X1  g08076(.A0(new_n10497_), .A1(new_n10490_), .B0(new_n10512_), .Y(new_n10513_));
  OR2X1    g08077(.A(new_n10513_), .B(pi0299), .Y(new_n10514_));
  AOI21X1  g08078(.A0(new_n10511_), .A1(new_n10498_), .B0(new_n10514_), .Y(new_n10515_));
  AOI21X1  g08079(.A0(new_n10483_), .A1(new_n10344_), .B0(new_n4611_), .Y(new_n10516_));
  INVX1    g08080(.A(new_n10484_), .Y(new_n10517_));
  OAI21X1  g08081(.A0(new_n10487_), .A1(new_n2776_), .B0(new_n4611_), .Y(new_n10518_));
  AOI21X1  g08082(.A0(new_n10517_), .A1(new_n2776_), .B0(new_n10518_), .Y(new_n10519_));
  OAI21X1  g08083(.A0(new_n10519_), .A1(new_n10516_), .B0(new_n5220_), .Y(new_n10520_));
  INVX1    g08084(.A(new_n10345_), .Y(new_n10521_));
  INVX1    g08085(.A(new_n10493_), .Y(new_n10522_));
  AOI21X1  g08086(.A0(new_n10500_), .A1(new_n10481_), .B0(new_n10342_), .Y(new_n10523_));
  OAI22X1  g08087(.A0(new_n10523_), .A1(new_n10521_), .B0(new_n10522_), .B1(new_n10453_), .Y(new_n10524_));
  AOI22X1  g08088(.A0(new_n10524_), .A1(pi0216), .B0(new_n10520_), .B1(new_n7187_), .Y(new_n10525_));
  OAI21X1  g08089(.A0(new_n10347_), .A1(new_n10341_), .B0(new_n5221_), .Y(new_n10526_));
  NAND2X1  g08090(.A(new_n10526_), .B(new_n7408_), .Y(new_n10527_));
  AND2X1   g08091(.A(new_n10526_), .B(new_n7378_), .Y(new_n10528_));
  AOI21X1  g08092(.A0(new_n10528_), .A1(new_n10520_), .B0(new_n5215_), .Y(new_n10529_));
  OAI21X1  g08093(.A0(new_n10527_), .A1(new_n10525_), .B0(new_n10529_), .Y(new_n10530_));
  AND3X1   g08094(.A(new_n2933_), .B(new_n2940_), .C(pi0222), .Y(new_n10531_));
  OAI21X1  g08095(.A0(new_n10531_), .A1(new_n5331_), .B0(new_n10481_), .Y(new_n10532_));
  AND3X1   g08096(.A(new_n10340_), .B(new_n5215_), .C(new_n2534_), .Y(new_n10533_));
  AOI21X1  g08097(.A0(new_n10533_), .A1(new_n10532_), .B0(new_n2939_), .Y(new_n10534_));
  OAI21X1  g08098(.A0(new_n10530_), .A1(new_n10515_), .B0(new_n10534_), .Y(new_n10535_));
  OR3X1    g08099(.A(new_n10386_), .B(pi0232), .C(pi0039), .Y(new_n10536_));
  AND3X1   g08100(.A(new_n10536_), .B(new_n10535_), .C(new_n10480_), .Y(new_n10537_));
  OAI22X1  g08101(.A0(new_n10537_), .A1(pi0038), .B0(new_n10362_), .B1(new_n10361_), .Y(new_n10538_));
  INVX1    g08102(.A(new_n5813_), .Y(new_n10539_));
  AOI21X1  g08103(.A0(new_n10341_), .A1(pi0100), .B0(new_n10539_), .Y(new_n10540_));
  INVX1    g08104(.A(new_n10540_), .Y(new_n10541_));
  AOI21X1  g08105(.A0(new_n10359_), .A1(pi0100), .B0(new_n10541_), .Y(new_n10542_));
  OR4X1    g08106(.A(pi0092), .B(pi0075), .C(pi0074), .D(pi0054), .Y(new_n10543_));
  AND2X1   g08107(.A(new_n10543_), .B(new_n3131_), .Y(new_n10544_));
  OAI21X1  g08108(.A0(new_n10455_), .A1(pi0051), .B0(new_n10544_), .Y(new_n10545_));
  MX2X1    g08109(.A(new_n8634_), .B(new_n8623_), .S0(pi0299), .Y(new_n10546_));
  OR3X1    g08110(.A(new_n10546_), .B(new_n5048_), .C(new_n5215_), .Y(new_n10547_));
  AOI22X1  g08111(.A0(new_n10547_), .A1(pi0087), .B0(new_n10338_), .B1(new_n10336_), .Y(new_n10548_));
  OAI21X1  g08112(.A0(new_n10545_), .A1(new_n10359_), .B0(new_n10548_), .Y(new_n10549_));
  AOI21X1  g08113(.A0(new_n10542_), .A1(new_n10538_), .B0(new_n10549_), .Y(new_n10550_));
  OR3X1    g08114(.A(new_n10416_), .B(new_n10346_), .C(new_n5048_), .Y(new_n10551_));
  OR3X1    g08115(.A(new_n10383_), .B(new_n5048_), .C(pi0146), .Y(new_n10552_));
  NOR3X1   g08116(.A(new_n10379_), .B(new_n10373_), .C(new_n6738_), .Y(new_n10553_));
  INVX1    g08117(.A(new_n10553_), .Y(new_n10554_));
  NAND4X1  g08118(.A(new_n10554_), .B(new_n10377_), .C(new_n10366_), .D(new_n10340_), .Y(new_n10555_));
  AOI21X1  g08119(.A0(new_n10555_), .A1(new_n10370_), .B0(new_n5881_), .Y(new_n10556_));
  AOI21X1  g08120(.A0(new_n10499_), .A1(new_n10395_), .B0(new_n10556_), .Y(new_n10557_));
  AOI21X1  g08121(.A0(new_n10557_), .A1(pi0146), .B0(pi0161), .Y(new_n10558_));
  AOI22X1  g08122(.A0(new_n10558_), .A1(new_n10552_), .B0(new_n10551_), .B1(pi0161), .Y(new_n10559_));
  OAI22X1  g08123(.A0(new_n10473_), .A1(pi0161), .B0(new_n10430_), .B1(new_n10521_), .Y(new_n10560_));
  AOI21X1  g08124(.A0(new_n10560_), .A1(new_n7095_), .B0(new_n5215_), .Y(new_n10561_));
  OAI21X1  g08125(.A0(new_n10559_), .A1(new_n7060_), .B0(new_n10561_), .Y(new_n10562_));
  AND2X1   g08126(.A(new_n10562_), .B(pi0156), .Y(new_n10563_));
  NOR2X1   g08127(.A(new_n10416_), .B(new_n5048_), .Y(new_n10564_));
  INVX1    g08128(.A(new_n10564_), .Y(new_n10565_));
  AOI21X1  g08129(.A0(pi0142), .A1(pi0051), .B0(new_n10565_), .Y(new_n10566_));
  OR3X1    g08130(.A(new_n10383_), .B(new_n5048_), .C(pi0142), .Y(new_n10567_));
  AOI21X1  g08131(.A0(new_n10557_), .A1(pi0142), .B0(pi0144), .Y(new_n10568_));
  AOI21X1  g08132(.A0(new_n10568_), .A1(new_n10567_), .B0(new_n5203_), .Y(new_n10569_));
  OAI21X1  g08133(.A0(new_n10566_), .A1(new_n7344_), .B0(new_n10569_), .Y(new_n10570_));
  OR2X1    g08134(.A(new_n10446_), .B(pi0144), .Y(new_n10571_));
  AND2X1   g08135(.A(new_n10571_), .B(new_n5203_), .Y(new_n10572_));
  OAI21X1  g08136(.A0(new_n10430_), .A1(new_n10405_), .B0(new_n10572_), .Y(new_n10573_));
  AND2X1   g08137(.A(new_n10573_), .B(pi0179), .Y(new_n10574_));
  NOR2X1   g08138(.A(new_n10396_), .B(new_n10405_), .Y(new_n10575_));
  AOI21X1  g08139(.A0(new_n10554_), .A1(new_n10340_), .B0(pi0051), .Y(new_n10576_));
  OAI22X1  g08140(.A0(new_n10576_), .A1(new_n5881_), .B0(new_n10442_), .B1(new_n10394_), .Y(new_n10577_));
  INVX1    g08141(.A(new_n10577_), .Y(new_n10578_));
  OAI21X1  g08142(.A0(new_n10380_), .A1(new_n10342_), .B0(new_n5023_), .Y(new_n10579_));
  OAI21X1  g08143(.A0(new_n10579_), .A1(pi0142), .B0(new_n7344_), .Y(new_n10580_));
  AOI21X1  g08144(.A0(new_n10578_), .A1(pi0142), .B0(new_n10580_), .Y(new_n10581_));
  OR3X1    g08145(.A(new_n10581_), .B(new_n10575_), .C(new_n5203_), .Y(new_n10582_));
  AOI21X1  g08146(.A0(new_n10356_), .A1(new_n5203_), .B0(pi0179), .Y(new_n10583_));
  AOI22X1  g08147(.A0(new_n10583_), .A1(new_n10582_), .B0(new_n10574_), .B1(new_n10570_), .Y(new_n10584_));
  OAI21X1  g08148(.A0(new_n10584_), .A1(pi0299), .B0(new_n2939_), .Y(new_n10585_));
  OAI21X1  g08149(.A0(new_n2985_), .A1(new_n2536_), .B0(pi0142), .Y(new_n10586_));
  OR2X1    g08150(.A(new_n10485_), .B(pi0142), .Y(new_n10587_));
  AND3X1   g08151(.A(new_n10587_), .B(new_n10492_), .C(new_n6848_), .Y(new_n10588_));
  AOI21X1  g08152(.A0(new_n10588_), .A1(new_n10586_), .B0(new_n10405_), .Y(new_n10589_));
  NAND2X1  g08153(.A(new_n10355_), .B(new_n7344_), .Y(new_n10590_));
  OAI21X1  g08154(.A0(new_n10590_), .A1(new_n10505_), .B0(pi0181), .Y(new_n10591_));
  AOI21X1  g08155(.A0(new_n10356_), .A1(new_n5204_), .B0(pi0299), .Y(new_n10592_));
  OAI21X1  g08156(.A0(new_n10591_), .A1(new_n10589_), .B0(new_n10592_), .Y(new_n10593_));
  NOR4X1   g08157(.A(new_n5048_), .B(new_n2985_), .C(new_n2536_), .D(pi0287), .Y(new_n10594_));
  AOI21X1  g08158(.A0(new_n10504_), .A1(new_n10452_), .B0(new_n7187_), .Y(new_n10595_));
  OAI21X1  g08159(.A0(new_n10594_), .A1(new_n10521_), .B0(new_n10595_), .Y(new_n10596_));
  AOI21X1  g08160(.A0(new_n10347_), .A1(new_n7187_), .B0(new_n7483_), .Y(new_n10597_));
  NOR3X1   g08161(.A(new_n10347_), .B(new_n2933_), .C(pi0159), .Y(new_n10598_));
  OR2X1    g08162(.A(new_n10598_), .B(new_n9566_), .Y(new_n10599_));
  AOI21X1  g08163(.A0(new_n10597_), .A1(new_n10596_), .B0(new_n10599_), .Y(new_n10600_));
  AOI21X1  g08164(.A0(new_n10600_), .A1(new_n10593_), .B0(pi0038), .Y(new_n10601_));
  OAI21X1  g08165(.A0(new_n10585_), .A1(new_n10563_), .B0(new_n10601_), .Y(new_n10602_));
  INVX1    g08166(.A(new_n10361_), .Y(new_n10603_));
  OAI21X1  g08167(.A0(new_n10579_), .A1(pi0146), .B0(new_n4611_), .Y(new_n10604_));
  AOI21X1  g08168(.A0(new_n10578_), .A1(pi0146), .B0(new_n10604_), .Y(new_n10605_));
  AOI21X1  g08169(.A0(new_n10397_), .A1(new_n10345_), .B0(new_n10605_), .Y(new_n10606_));
  AOI21X1  g08170(.A0(new_n10358_), .A1(new_n7094_), .B0(new_n5215_), .Y(new_n10607_));
  OAI21X1  g08171(.A0(new_n10606_), .A1(new_n7060_), .B0(new_n10607_), .Y(new_n10608_));
  NOR3X1   g08172(.A(pi0156), .B(pi0039), .C(pi0038), .Y(new_n10609_));
  AOI21X1  g08173(.A0(new_n10609_), .A1(new_n10608_), .B0(new_n10603_), .Y(new_n10610_));
  OAI21X1  g08174(.A0(new_n10360_), .A1(new_n3007_), .B0(new_n5813_), .Y(new_n10611_));
  AOI21X1  g08175(.A0(new_n10610_), .A1(new_n10602_), .B0(new_n10611_), .Y(new_n10612_));
  INVX1    g08176(.A(new_n10544_), .Y(new_n10613_));
  NAND2X1  g08177(.A(new_n10547_), .B(pi0087), .Y(new_n10614_));
  AND2X1   g08178(.A(new_n10614_), .B(new_n10339_), .Y(new_n10615_));
  OAI21X1  g08179(.A0(new_n10613_), .A1(new_n10359_), .B0(new_n10615_), .Y(new_n10616_));
  OAI21X1  g08180(.A0(new_n10616_), .A1(new_n10612_), .B0(new_n6489_), .Y(new_n10617_));
  OAI21X1  g08181(.A0(new_n10617_), .A1(new_n10550_), .B0(new_n10351_), .Y(po0279));
  AOI21X1  g08182(.A0(new_n10323_), .A1(new_n5880_), .B0(new_n10303_), .Y(new_n10619_));
  OAI21X1  g08183(.A0(new_n10327_), .A1(new_n6295_), .B0(new_n6072_), .Y(new_n10620_));
  NAND2X1  g08184(.A(new_n10620_), .B(new_n6489_), .Y(new_n10621_));
  OAI22X1  g08185(.A0(new_n10621_), .A1(new_n10619_), .B0(new_n6711_), .B1(new_n10124_), .Y(po0280));
  NAND2X1  g08186(.A(new_n6844_), .B(new_n2547_), .Y(new_n10623_));
  OR3X1    g08187(.A(new_n10623_), .B(new_n5221_), .C(new_n5062_), .Y(new_n10624_));
  OR4X1    g08188(.A(new_n8165_), .B(new_n7555_), .C(new_n5928_), .D(new_n2547_), .Y(new_n10625_));
  OAI21X1  g08189(.A0(new_n10625_), .A1(new_n5082_), .B0(new_n2939_), .Y(new_n10626_));
  NAND2X1  g08190(.A(new_n10626_), .B(po1038), .Y(new_n10627_));
  AOI21X1  g08191(.A0(new_n10624_), .A1(pi0039), .B0(new_n10627_), .Y(new_n10628_));
  NOR4X1   g08192(.A(new_n10543_), .B(pi0100), .C(pi0087), .D(pi0038), .Y(new_n10629_));
  OR4X1    g08193(.A(new_n10623_), .B(new_n5221_), .C(new_n5062_), .D(new_n2933_), .Y(new_n10630_));
  OR4X1    g08194(.A(new_n10623_), .B(new_n5248_), .C(new_n5049_), .D(pi0299), .Y(new_n10631_));
  AND3X1   g08195(.A(new_n10631_), .B(new_n10630_), .C(pi0039), .Y(new_n10632_));
  NOR3X1   g08196(.A(new_n2475_), .B(new_n7569_), .C(pi0109), .Y(new_n10633_));
  INVX1    g08197(.A(new_n2597_), .Y(new_n10634_));
  INVX1    g08198(.A(new_n2461_), .Y(new_n10635_));
  NOR2X1   g08199(.A(new_n2632_), .B(pi0036), .Y(new_n10636_));
  OAI21X1  g08200(.A0(new_n5128_), .A1(pi0111), .B0(new_n10636_), .Y(new_n10637_));
  OAI21X1  g08201(.A0(new_n2592_), .A1(new_n2591_), .B0(new_n2641_), .Y(new_n10638_));
  AOI21X1  g08202(.A0(new_n10637_), .A1(new_n10635_), .B0(new_n10638_), .Y(new_n10639_));
  OAI21X1  g08203(.A0(new_n10639_), .A1(pi0083), .B0(new_n10634_), .Y(new_n10640_));
  AOI21X1  g08204(.A0(new_n10640_), .A1(new_n2590_), .B0(new_n5136_), .Y(new_n10641_));
  OAI21X1  g08205(.A0(new_n10641_), .A1(pi0081), .B0(new_n8462_), .Y(new_n10642_));
  AOI21X1  g08206(.A0(new_n10642_), .A1(new_n2682_), .B0(new_n2478_), .Y(new_n10643_));
  NOR2X1   g08207(.A(new_n10633_), .B(new_n2682_), .Y(new_n10644_));
  NOR2X1   g08208(.A(new_n10644_), .B(new_n6932_), .Y(new_n10645_));
  NOR4X1   g08209(.A(new_n2478_), .B(pi0093), .C(pi0090), .D(new_n2530_), .Y(new_n10646_));
  AOI22X1  g08210(.A0(new_n10646_), .A1(new_n10633_), .B0(new_n10645_), .B1(new_n10643_), .Y(new_n10647_));
  OAI21X1  g08211(.A0(new_n10647_), .A1(new_n7619_), .B0(new_n2547_), .Y(new_n10648_));
  NOR2X1   g08212(.A(new_n2683_), .B(pi0093), .Y(new_n10649_));
  AOI21X1  g08213(.A0(new_n10643_), .A1(new_n10649_), .B0(pi0072), .Y(new_n10650_));
  OR2X1    g08214(.A(new_n9700_), .B(new_n5170_), .Y(new_n10651_));
  OAI21X1  g08215(.A0(new_n10651_), .A1(new_n10650_), .B0(new_n2939_), .Y(new_n10652_));
  AOI21X1  g08216(.A0(new_n10648_), .A1(new_n9700_), .B0(new_n10652_), .Y(new_n10653_));
  OAI21X1  g08217(.A0(new_n10653_), .A1(new_n10632_), .B0(new_n10629_), .Y(new_n10654_));
  INVX1    g08218(.A(new_n10629_), .Y(new_n10655_));
  AOI21X1  g08219(.A0(new_n9700_), .A1(pi0110), .B0(pi0039), .Y(new_n10656_));
  OAI21X1  g08220(.A0(new_n10656_), .A1(new_n10632_), .B0(new_n10655_), .Y(new_n10657_));
  AND2X1   g08221(.A(new_n10657_), .B(new_n6489_), .Y(new_n10658_));
  AOI21X1  g08222(.A0(new_n10658_), .A1(new_n10654_), .B0(new_n10628_), .Y(po0281));
  INVX1    g08223(.A(pi0125), .Y(new_n10660_));
  XOR2X1   g08224(.A(pi0133), .B(pi0125), .Y(new_n10661_));
  AOI21X1  g08225(.A0(new_n10335_), .A1(new_n10660_), .B0(new_n10661_), .Y(new_n10662_));
  INVX1    g08226(.A(new_n10662_), .Y(new_n10663_));
  AOI22X1  g08227(.A0(new_n10442_), .A1(new_n3193_), .B0(new_n10387_), .B1(pi0172), .Y(new_n10664_));
  INVX1    g08228(.A(new_n10664_), .Y(new_n10665_));
  AOI22X1  g08229(.A0(new_n10665_), .A1(pi0232), .B0(new_n10663_), .B1(new_n10341_), .Y(new_n10666_));
  AND3X1   g08230(.A(new_n5023_), .B(pi0232), .C(pi0087), .Y(new_n10667_));
  AOI21X1  g08231(.A0(new_n10667_), .A1(pi0162), .B0(new_n6489_), .Y(new_n10668_));
  OAI21X1  g08232(.A0(new_n10666_), .A1(pi0087), .B0(new_n10668_), .Y(new_n10669_));
  INVX1    g08233(.A(new_n7426_), .Y(new_n10670_));
  NOR3X1   g08234(.A(pi0468), .B(pi0332), .C(pi0152), .Y(new_n10671_));
  INVX1    g08235(.A(new_n10671_), .Y(new_n10672_));
  OAI21X1  g08236(.A0(new_n10456_), .A1(pi0152), .B0(new_n7307_), .Y(new_n10673_));
  AOI21X1  g08237(.A0(new_n10672_), .A1(new_n10411_), .B0(new_n10673_), .Y(new_n10674_));
  INVX1    g08238(.A(new_n10380_), .Y(new_n10675_));
  NOR3X1   g08239(.A(new_n10437_), .B(new_n10368_), .C(new_n10455_), .Y(new_n10676_));
  AND3X1   g08240(.A(new_n8143_), .B(new_n5048_), .C(pi0072), .Y(new_n10677_));
  INVX1    g08241(.A(new_n10677_), .Y(new_n10678_));
  AOI22X1  g08242(.A0(new_n10678_), .A1(new_n10437_), .B0(new_n10676_), .B1(new_n10675_), .Y(new_n10679_));
  NOR3X1   g08243(.A(new_n10679_), .B(new_n7307_), .C(pi0152), .Y(new_n10680_));
  OAI22X1  g08244(.A0(new_n10680_), .A1(new_n10674_), .B0(new_n10462_), .B1(new_n7084_), .Y(new_n10681_));
  AOI21X1  g08245(.A0(new_n8143_), .A1(pi0072), .B0(new_n5023_), .Y(new_n10682_));
  AOI21X1  g08246(.A0(new_n10401_), .A1(new_n5023_), .B0(new_n10682_), .Y(new_n10683_));
  AND2X1   g08247(.A(new_n10683_), .B(new_n7084_), .Y(new_n10684_));
  NOR3X1   g08248(.A(new_n10396_), .B(new_n10411_), .C(new_n10387_), .Y(new_n10685_));
  NOR2X1   g08249(.A(new_n10685_), .B(new_n7084_), .Y(new_n10686_));
  OR4X1    g08250(.A(new_n10686_), .B(new_n10684_), .C(new_n7307_), .D(new_n3193_), .Y(new_n10687_));
  AOI21X1  g08251(.A0(new_n10687_), .A1(new_n10681_), .B0(new_n10670_), .Y(new_n10688_));
  MX2X1    g08252(.A(new_n10421_), .B(new_n10411_), .S0(new_n5048_), .Y(new_n10689_));
  INVX1    g08253(.A(new_n10689_), .Y(new_n10690_));
  AOI21X1  g08254(.A0(new_n10416_), .A1(new_n10412_), .B0(new_n10682_), .Y(new_n10691_));
  AOI21X1  g08255(.A0(new_n10691_), .A1(pi0172), .B0(new_n3193_), .Y(new_n10692_));
  OAI21X1  g08256(.A0(new_n10690_), .A1(pi0172), .B0(new_n10692_), .Y(new_n10693_));
  AOI22X1  g08257(.A0(new_n10678_), .A1(new_n10437_), .B0(new_n10386_), .B1(new_n5023_), .Y(new_n10694_));
  INVX1    g08258(.A(new_n10694_), .Y(new_n10695_));
  AOI21X1  g08259(.A0(new_n10387_), .A1(pi0172), .B0(pi0152), .Y(new_n10696_));
  AOI21X1  g08260(.A0(new_n10696_), .A1(new_n10695_), .B0(new_n7307_), .Y(new_n10697_));
  MX2X1    g08261(.A(new_n10427_), .B(new_n10411_), .S0(new_n5048_), .Y(new_n10698_));
  NOR2X1   g08262(.A(new_n10677_), .B(new_n10438_), .Y(new_n10699_));
  OAI21X1  g08263(.A0(new_n10699_), .A1(pi0152), .B0(new_n7084_), .Y(new_n10700_));
  AOI21X1  g08264(.A0(new_n10698_), .A1(pi0152), .B0(new_n10700_), .Y(new_n10701_));
  NOR3X1   g08265(.A(new_n10430_), .B(new_n10411_), .C(new_n10387_), .Y(new_n10702_));
  NOR2X1   g08266(.A(new_n10702_), .B(new_n3193_), .Y(new_n10703_));
  INVX1    g08267(.A(new_n10676_), .Y(new_n10704_));
  NOR4X1   g08268(.A(new_n10704_), .B(new_n10378_), .C(new_n10368_), .D(new_n10342_), .Y(new_n10705_));
  NOR2X1   g08269(.A(new_n10705_), .B(new_n10682_), .Y(new_n10706_));
  INVX1    g08270(.A(new_n10706_), .Y(new_n10707_));
  OAI21X1  g08271(.A0(new_n10707_), .A1(pi0152), .B0(pi0172), .Y(new_n10708_));
  OAI21X1  g08272(.A0(new_n10708_), .A1(new_n10703_), .B0(new_n7307_), .Y(new_n10709_));
  OAI21X1  g08273(.A0(new_n10709_), .A1(new_n10701_), .B0(new_n7430_), .Y(new_n10710_));
  AOI21X1  g08274(.A0(new_n10697_), .A1(new_n10693_), .B0(new_n10710_), .Y(new_n10711_));
  OAI21X1  g08275(.A0(new_n10711_), .A1(new_n10688_), .B0(pi0299), .Y(new_n10712_));
  NAND2X1  g08276(.A(new_n10683_), .B(pi0145), .Y(new_n10713_));
  AOI21X1  g08277(.A0(new_n10411_), .A1(new_n5202_), .B0(new_n6851_), .Y(new_n10714_));
  NAND2X1  g08278(.A(new_n10679_), .B(pi0145), .Y(new_n10715_));
  INVX1    g08279(.A(new_n10456_), .Y(new_n10716_));
  NOR2X1   g08280(.A(new_n10677_), .B(new_n10716_), .Y(new_n10717_));
  INVX1    g08281(.A(new_n10717_), .Y(new_n10718_));
  AOI21X1  g08282(.A0(new_n10718_), .A1(new_n5202_), .B0(pi0174), .Y(new_n10719_));
  AOI22X1  g08283(.A0(new_n10719_), .A1(new_n10715_), .B0(new_n10714_), .B1(new_n10713_), .Y(new_n10720_));
  MX2X1    g08284(.A(new_n10462_), .B(new_n5202_), .S0(new_n10396_), .Y(new_n10721_));
  AOI21X1  g08285(.A0(new_n10721_), .A1(new_n10412_), .B0(new_n6851_), .Y(new_n10722_));
  AOI21X1  g08286(.A0(new_n10675_), .A1(new_n10462_), .B0(new_n5202_), .Y(new_n10723_));
  OAI21X1  g08287(.A0(new_n10723_), .A1(new_n10704_), .B0(new_n6851_), .Y(new_n10724_));
  OAI21X1  g08288(.A0(new_n10724_), .A1(new_n10682_), .B0(pi0193), .Y(new_n10725_));
  OAI22X1  g08289(.A0(new_n10725_), .A1(new_n10722_), .B0(new_n10720_), .B1(pi0193), .Y(new_n10726_));
  AND3X1   g08290(.A(new_n10726_), .B(new_n2933_), .C(new_n7450_), .Y(new_n10727_));
  AOI21X1  g08291(.A0(new_n10698_), .A1(new_n5202_), .B0(pi0193), .Y(new_n10728_));
  OAI21X1  g08292(.A0(new_n10690_), .A1(new_n5202_), .B0(new_n10728_), .Y(new_n10729_));
  NAND2X1  g08293(.A(new_n10691_), .B(pi0145), .Y(new_n10730_));
  INVX1    g08294(.A(new_n10702_), .Y(new_n10731_));
  AOI21X1  g08295(.A0(new_n10731_), .A1(new_n5202_), .B0(new_n6885_), .Y(new_n10732_));
  AOI21X1  g08296(.A0(new_n10732_), .A1(new_n10730_), .B0(new_n6851_), .Y(new_n10733_));
  OAI21X1  g08297(.A0(new_n10699_), .A1(pi0193), .B0(new_n5202_), .Y(new_n10734_));
  AOI21X1  g08298(.A0(new_n10706_), .A1(pi0193), .B0(new_n10734_), .Y(new_n10735_));
  AND3X1   g08299(.A(new_n5023_), .B(pi0193), .C(pi0051), .Y(new_n10736_));
  OR2X1    g08300(.A(new_n10736_), .B(new_n5202_), .Y(new_n10737_));
  OAI21X1  g08301(.A0(new_n10737_), .A1(new_n10694_), .B0(new_n6851_), .Y(new_n10738_));
  OAI21X1  g08302(.A0(new_n10738_), .A1(new_n10735_), .B0(new_n7418_), .Y(new_n10739_));
  AOI21X1  g08303(.A0(new_n10733_), .A1(new_n10729_), .B0(new_n10739_), .Y(new_n10740_));
  OAI21X1  g08304(.A0(new_n10740_), .A1(new_n10727_), .B0(new_n2979_), .Y(new_n10741_));
  AOI21X1  g08305(.A0(new_n10741_), .A1(new_n10712_), .B0(new_n7260_), .Y(new_n10742_));
  MX2X1    g08306(.A(new_n6270_), .B(new_n6264_), .S0(new_n2933_), .Y(new_n10743_));
  AOI21X1  g08307(.A0(new_n10743_), .A1(new_n2987_), .B0(pi0232), .Y(new_n10744_));
  NOR2X1   g08308(.A(new_n10744_), .B(new_n2939_), .Y(new_n10745_));
  INVX1    g08309(.A(new_n10745_), .Y(new_n10746_));
  NOR2X1   g08310(.A(new_n10482_), .B(new_n5048_), .Y(new_n10747_));
  INVX1    g08311(.A(new_n10747_), .Y(new_n10748_));
  OAI21X1  g08312(.A0(new_n5023_), .A1(new_n2986_), .B0(new_n10748_), .Y(new_n10749_));
  OAI21X1  g08313(.A0(new_n10485_), .A1(pi0051), .B0(new_n5023_), .Y(new_n10750_));
  OAI21X1  g08314(.A0(new_n5023_), .A1(new_n2986_), .B0(new_n10750_), .Y(new_n10751_));
  MX2X1    g08315(.A(new_n10751_), .B(new_n10749_), .S0(new_n3193_), .Y(new_n10752_));
  OR2X1    g08316(.A(pi0172), .B(new_n2534_), .Y(new_n10753_));
  AOI21X1  g08317(.A0(new_n10753_), .A1(new_n10752_), .B0(pi0216), .Y(new_n10754_));
  AOI22X1  g08318(.A0(new_n10754_), .A1(new_n5220_), .B0(new_n10664_), .B1(new_n6271_), .Y(new_n10755_));
  OR2X1    g08319(.A(new_n10755_), .B(new_n7096_), .Y(new_n10756_));
  NOR4X1   g08320(.A(new_n10500_), .B(new_n5881_), .C(new_n2536_), .D(pi0096), .Y(new_n10757_));
  NOR2X1   g08321(.A(new_n10757_), .B(new_n10387_), .Y(new_n10758_));
  AOI21X1  g08322(.A0(new_n10758_), .A1(pi0224), .B0(new_n5248_), .Y(new_n10759_));
  OAI21X1  g08323(.A0(new_n10751_), .A1(new_n6265_), .B0(new_n10759_), .Y(new_n10760_));
  NAND2X1  g08324(.A(new_n10760_), .B(new_n10462_), .Y(new_n10761_));
  AOI21X1  g08325(.A0(new_n10492_), .A1(new_n10481_), .B0(new_n2942_), .Y(new_n10762_));
  OAI22X1  g08326(.A0(new_n10762_), .A1(new_n5248_), .B0(new_n10341_), .B1(new_n5048_), .Y(new_n10763_));
  OAI21X1  g08327(.A0(new_n10749_), .A1(new_n6265_), .B0(new_n10763_), .Y(new_n10764_));
  OAI21X1  g08328(.A0(new_n10764_), .A1(pi0174), .B0(pi0193), .Y(new_n10765_));
  AOI21X1  g08329(.A0(new_n10761_), .A1(pi0174), .B0(new_n10765_), .Y(new_n10766_));
  MX2X1    g08330(.A(new_n10502_), .B(new_n2986_), .S0(new_n5048_), .Y(new_n10767_));
  AND2X1   g08331(.A(new_n10767_), .B(new_n2942_), .Y(new_n10768_));
  INVX1    g08332(.A(new_n10768_), .Y(new_n10769_));
  AOI21X1  g08333(.A0(new_n10504_), .A1(pi0224), .B0(new_n5248_), .Y(new_n10770_));
  AOI21X1  g08334(.A0(new_n10770_), .A1(new_n10769_), .B0(new_n10496_), .Y(new_n10771_));
  AOI21X1  g08335(.A0(new_n10492_), .A1(new_n6848_), .B0(new_n6264_), .Y(new_n10772_));
  NOR3X1   g08336(.A(new_n10772_), .B(new_n2985_), .C(new_n2536_), .Y(new_n10773_));
  AOI21X1  g08337(.A0(new_n10773_), .A1(pi0174), .B0(pi0193), .Y(new_n10774_));
  OAI21X1  g08338(.A0(new_n10771_), .A1(pi0174), .B0(new_n10774_), .Y(new_n10775_));
  NAND2X1  g08339(.A(new_n10775_), .B(pi0180), .Y(new_n10776_));
  NOR2X1   g08340(.A(new_n10354_), .B(new_n6264_), .Y(new_n10777_));
  OR2X1    g08341(.A(new_n10777_), .B(new_n10767_), .Y(new_n10778_));
  NOR3X1   g08342(.A(new_n6265_), .B(new_n2985_), .C(new_n2536_), .Y(new_n10779_));
  AOI21X1  g08343(.A0(new_n10779_), .A1(pi0174), .B0(new_n10736_), .Y(new_n10780_));
  OAI21X1  g08344(.A0(new_n10778_), .A1(pi0174), .B0(new_n10780_), .Y(new_n10781_));
  AOI21X1  g08345(.A0(new_n10781_), .A1(new_n5203_), .B0(pi0299), .Y(new_n10782_));
  OAI21X1  g08346(.A0(new_n10776_), .A1(new_n10766_), .B0(new_n10782_), .Y(new_n10783_));
  AOI21X1  g08347(.A0(new_n10492_), .A1(new_n10481_), .B0(new_n10354_), .Y(new_n10784_));
  INVX1    g08348(.A(new_n10784_), .Y(new_n10785_));
  OAI21X1  g08349(.A0(new_n10785_), .A1(pi0152), .B0(pi0172), .Y(new_n10786_));
  AOI21X1  g08350(.A0(new_n10758_), .A1(pi0152), .B0(new_n10786_), .Y(new_n10787_));
  NOR2X1   g08351(.A(new_n10594_), .B(new_n3193_), .Y(new_n10788_));
  OAI21X1  g08352(.A0(new_n10503_), .A1(pi0152), .B0(new_n7084_), .Y(new_n10789_));
  OAI21X1  g08353(.A0(new_n10789_), .A1(new_n10788_), .B0(pi0216), .Y(new_n10790_));
  OAI21X1  g08354(.A0(new_n10790_), .A1(new_n10787_), .B0(new_n5220_), .Y(new_n10791_));
  AOI21X1  g08355(.A0(new_n10665_), .A1(new_n5221_), .B0(new_n7060_), .Y(new_n10792_));
  OAI21X1  g08356(.A0(new_n10791_), .A1(new_n10754_), .B0(new_n10792_), .Y(new_n10793_));
  NAND3X1  g08357(.A(new_n10793_), .B(new_n10783_), .C(new_n10756_), .Y(new_n10794_));
  AOI21X1  g08358(.A0(new_n10794_), .A1(pi0232), .B0(new_n10746_), .Y(new_n10795_));
  AOI21X1  g08359(.A0(new_n10412_), .A1(new_n5215_), .B0(pi0039), .Y(new_n10796_));
  NOR3X1   g08360(.A(new_n10796_), .B(new_n10795_), .C(pi0038), .Y(new_n10797_));
  NAND2X1  g08361(.A(new_n10664_), .B(pi0299), .Y(new_n10798_));
  AND2X1   g08362(.A(new_n10442_), .B(new_n6851_), .Y(new_n10799_));
  OR3X1    g08363(.A(new_n10799_), .B(new_n10736_), .C(pi0299), .Y(new_n10800_));
  AND3X1   g08364(.A(new_n10800_), .B(new_n10798_), .C(pi0232), .Y(new_n10801_));
  OAI21X1  g08365(.A0(new_n10801_), .A1(new_n2979_), .B0(new_n3007_), .Y(new_n10802_));
  OR3X1    g08366(.A(new_n10802_), .B(new_n10797_), .C(new_n10742_), .Y(new_n10803_));
  NAND4X1  g08367(.A(new_n10800_), .B(new_n10798_), .C(pi0232), .D(pi0100), .Y(new_n10804_));
  AND2X1   g08368(.A(new_n10804_), .B(new_n5813_), .Y(new_n10805_));
  MX2X1    g08369(.A(new_n7306_), .B(new_n7353_), .S0(new_n2933_), .Y(new_n10806_));
  OAI21X1  g08370(.A0(new_n10806_), .A1(new_n6820_), .B0(pi0087), .Y(new_n10807_));
  AND2X1   g08371(.A(new_n10807_), .B(new_n10662_), .Y(new_n10808_));
  OAI21X1  g08372(.A0(new_n10801_), .A1(new_n10613_), .B0(new_n10808_), .Y(new_n10809_));
  AOI21X1  g08373(.A0(new_n10805_), .A1(new_n10803_), .B0(new_n10809_), .Y(new_n10810_));
  INVX1    g08374(.A(new_n10384_), .Y(new_n10811_));
  NAND3X1  g08375(.A(new_n10414_), .B(new_n10394_), .C(new_n2479_), .Y(new_n10812_));
  NAND3X1  g08376(.A(new_n10812_), .B(new_n10811_), .C(new_n5202_), .Y(new_n10813_));
  NOR3X1   g08377(.A(new_n10430_), .B(new_n10384_), .C(new_n5202_), .Y(new_n10814_));
  NOR2X1   g08378(.A(new_n10814_), .B(pi0174), .Y(new_n10815_));
  NOR2X1   g08379(.A(new_n10557_), .B(new_n10384_), .Y(new_n10816_));
  NOR2X1   g08380(.A(new_n10381_), .B(new_n5023_), .Y(new_n10817_));
  NOR3X1   g08381(.A(new_n10817_), .B(new_n10378_), .C(new_n10354_), .Y(new_n10818_));
  INVX1    g08382(.A(new_n10818_), .Y(new_n10819_));
  AOI21X1  g08383(.A0(new_n10382_), .A1(new_n5202_), .B0(new_n10819_), .Y(new_n10820_));
  AND2X1   g08384(.A(new_n10820_), .B(new_n2984_), .Y(new_n10821_));
  NOR3X1   g08385(.A(new_n10821_), .B(new_n10816_), .C(new_n6851_), .Y(new_n10822_));
  OR2X1    g08386(.A(new_n10822_), .B(new_n6885_), .Y(new_n10823_));
  AOI21X1  g08387(.A0(new_n10815_), .A1(new_n10813_), .B0(new_n10823_), .Y(new_n10824_));
  OR3X1    g08388(.A(new_n10564_), .B(new_n10384_), .C(pi0145), .Y(new_n10825_));
  AOI21X1  g08389(.A0(new_n10814_), .A1(new_n2534_), .B0(pi0174), .Y(new_n10826_));
  OAI21X1  g08390(.A0(new_n10820_), .A1(new_n6851_), .B0(new_n6885_), .Y(new_n10827_));
  AOI21X1  g08391(.A0(new_n10826_), .A1(new_n10825_), .B0(new_n10827_), .Y(new_n10828_));
  OR3X1    g08392(.A(new_n10828_), .B(new_n10824_), .C(new_n7414_), .Y(new_n10829_));
  MX2X1    g08393(.A(new_n10383_), .B(new_n2534_), .S0(new_n5023_), .Y(new_n10830_));
  AND2X1   g08394(.A(new_n10396_), .B(new_n5202_), .Y(new_n10831_));
  OAI22X1  g08395(.A0(new_n10831_), .A1(pi0174), .B0(new_n10455_), .B1(new_n5202_), .Y(new_n10832_));
  AOI21X1  g08396(.A0(new_n10378_), .A1(new_n5048_), .B0(new_n10382_), .Y(new_n10833_));
  AOI22X1  g08397(.A0(new_n10833_), .A1(pi0174), .B0(new_n10832_), .B1(new_n10830_), .Y(new_n10834_));
  AND2X1   g08398(.A(pi0174), .B(new_n5202_), .Y(new_n10835_));
  AOI22X1  g08399(.A0(new_n10835_), .A1(new_n10577_), .B0(new_n10499_), .B1(pi0145), .Y(new_n10836_));
  OAI21X1  g08400(.A0(new_n10831_), .A1(pi0174), .B0(new_n10836_), .Y(new_n10837_));
  NOR2X1   g08401(.A(new_n10384_), .B(new_n6885_), .Y(new_n10838_));
  AOI21X1  g08402(.A0(new_n10838_), .A1(new_n10837_), .B0(new_n7419_), .Y(new_n10839_));
  OAI21X1  g08403(.A0(new_n10834_), .A1(pi0193), .B0(new_n10839_), .Y(new_n10840_));
  AOI21X1  g08404(.A0(new_n10840_), .A1(new_n10829_), .B0(pi0038), .Y(new_n10841_));
  AND2X1   g08405(.A(new_n10812_), .B(new_n10811_), .Y(new_n10842_));
  OAI21X1  g08406(.A0(new_n10557_), .A1(new_n10384_), .B0(pi0152), .Y(new_n10843_));
  AND2X1   g08407(.A(new_n10843_), .B(pi0172), .Y(new_n10844_));
  OAI21X1  g08408(.A0(new_n10842_), .A1(pi0152), .B0(new_n10844_), .Y(new_n10845_));
  INVX1    g08409(.A(new_n10383_), .Y(new_n10846_));
  AOI21X1  g08410(.A0(new_n10672_), .A1(new_n10846_), .B0(pi0172), .Y(new_n10847_));
  OAI21X1  g08411(.A0(new_n10565_), .A1(pi0152), .B0(new_n10847_), .Y(new_n10848_));
  AOI21X1  g08412(.A0(new_n10848_), .A1(new_n10845_), .B0(pi0197), .Y(new_n10849_));
  INVX1    g08413(.A(new_n10430_), .Y(new_n10850_));
  AOI21X1  g08414(.A0(new_n10850_), .A1(new_n10811_), .B0(pi0152), .Y(new_n10851_));
  NOR3X1   g08415(.A(new_n10445_), .B(new_n10384_), .C(new_n7084_), .Y(new_n10852_));
  OAI21X1  g08416(.A0(new_n10819_), .A1(pi0172), .B0(pi0152), .Y(new_n10853_));
  AOI21X1  g08417(.A0(new_n10387_), .A1(new_n7084_), .B0(new_n7307_), .Y(new_n10854_));
  OAI21X1  g08418(.A0(new_n10853_), .A1(new_n10852_), .B0(new_n10854_), .Y(new_n10855_));
  AND2X1   g08419(.A(new_n7426_), .B(pi0299), .Y(new_n10856_));
  OAI21X1  g08420(.A0(new_n10855_), .A1(new_n10851_), .B0(new_n10856_), .Y(new_n10857_));
  NOR3X1   g08421(.A(new_n10396_), .B(new_n10384_), .C(pi0152), .Y(new_n10858_));
  INVX1    g08422(.A(new_n10833_), .Y(new_n10859_));
  OAI21X1  g08423(.A0(new_n10859_), .A1(new_n3193_), .B0(new_n7084_), .Y(new_n10860_));
  AOI21X1  g08424(.A0(new_n10858_), .A1(new_n10462_), .B0(new_n10860_), .Y(new_n10861_));
  OAI21X1  g08425(.A0(new_n10383_), .A1(new_n5023_), .B0(new_n10577_), .Y(new_n10862_));
  OAI21X1  g08426(.A0(new_n10862_), .A1(new_n3193_), .B0(pi0172), .Y(new_n10863_));
  OAI21X1  g08427(.A0(new_n10863_), .A1(new_n10858_), .B0(new_n7307_), .Y(new_n10864_));
  OAI22X1  g08428(.A0(new_n10499_), .A1(new_n3193_), .B0(new_n10383_), .B1(new_n5023_), .Y(new_n10865_));
  NAND2X1  g08429(.A(new_n10865_), .B(pi0172), .Y(new_n10866_));
  AOI21X1  g08430(.A0(new_n10442_), .A1(new_n3193_), .B0(pi0172), .Y(new_n10867_));
  OAI21X1  g08431(.A0(new_n10384_), .A1(new_n10354_), .B0(new_n10867_), .Y(new_n10868_));
  NAND3X1  g08432(.A(new_n10868_), .B(new_n10866_), .C(pi0197), .Y(new_n10869_));
  AND3X1   g08433(.A(new_n10869_), .B(new_n7430_), .C(pi0299), .Y(new_n10870_));
  OAI21X1  g08434(.A0(new_n10864_), .A1(new_n10861_), .B0(new_n10870_), .Y(new_n10871_));
  OAI21X1  g08435(.A0(new_n10857_), .A1(new_n10849_), .B0(new_n10871_), .Y(new_n10872_));
  OAI21X1  g08436(.A0(new_n10872_), .A1(new_n10841_), .B0(new_n7259_), .Y(new_n10873_));
  INVX1    g08437(.A(new_n10362_), .Y(new_n10874_));
  OAI21X1  g08438(.A0(new_n10665_), .A1(new_n10341_), .B0(new_n7187_), .Y(new_n10875_));
  OAI22X1  g08439(.A0(new_n10671_), .A1(new_n10482_), .B0(new_n10750_), .B1(pi0152), .Y(new_n10876_));
  AND2X1   g08440(.A(new_n10876_), .B(new_n7084_), .Y(new_n10877_));
  INVX1    g08441(.A(new_n10508_), .Y(new_n10878_));
  OAI21X1  g08442(.A0(new_n10878_), .A1(new_n3193_), .B0(pi0172), .Y(new_n10879_));
  AOI21X1  g08443(.A0(new_n10484_), .A1(new_n3193_), .B0(new_n10879_), .Y(new_n10880_));
  NOR3X1   g08444(.A(new_n10880_), .B(new_n10877_), .C(new_n7187_), .Y(new_n10881_));
  OAI21X1  g08445(.A0(new_n10462_), .A1(new_n7084_), .B0(pi0152), .Y(new_n10882_));
  OAI21X1  g08446(.A0(new_n10882_), .A1(new_n10523_), .B0(new_n6856_), .Y(new_n10883_));
  AOI21X1  g08447(.A0(new_n10696_), .A1(new_n10493_), .B0(new_n10883_), .Y(new_n10884_));
  OAI22X1  g08448(.A0(new_n10884_), .A1(new_n7060_), .B0(new_n10881_), .B1(new_n7096_), .Y(new_n10885_));
  NOR2X1   g08449(.A(new_n5023_), .B(new_n2534_), .Y(new_n10886_));
  AOI21X1  g08450(.A0(new_n10455_), .A1(new_n5048_), .B0(new_n6848_), .Y(new_n10887_));
  INVX1    g08451(.A(new_n10887_), .Y(new_n10888_));
  OAI22X1  g08452(.A0(new_n10888_), .A1(new_n10886_), .B0(new_n10517_), .B1(new_n7203_), .Y(new_n10889_));
  AOI21X1  g08453(.A0(new_n10481_), .A1(new_n6848_), .B0(new_n10342_), .Y(new_n10890_));
  NOR2X1   g08454(.A(new_n10890_), .B(new_n10387_), .Y(new_n10891_));
  OAI21X1  g08455(.A0(new_n10891_), .A1(new_n6851_), .B0(new_n5203_), .Y(new_n10892_));
  AOI21X1  g08456(.A0(new_n10889_), .A1(new_n6851_), .B0(new_n10892_), .Y(new_n10893_));
  AOI21X1  g08457(.A0(new_n10483_), .A1(new_n5048_), .B0(new_n7203_), .Y(new_n10894_));
  INVX1    g08458(.A(new_n10894_), .Y(new_n10895_));
  OAI22X1  g08459(.A0(new_n10895_), .A1(new_n7874_), .B0(new_n10888_), .B1(new_n10886_), .Y(new_n10896_));
  NOR2X1   g08460(.A(new_n10523_), .B(pi0051), .Y(new_n10897_));
  NOR2X1   g08461(.A(new_n10897_), .B(new_n5048_), .Y(new_n10898_));
  NOR2X1   g08462(.A(new_n10898_), .B(new_n10890_), .Y(new_n10899_));
  OAI21X1  g08463(.A0(new_n10899_), .A1(new_n6851_), .B0(pi0180), .Y(new_n10900_));
  AOI21X1  g08464(.A0(new_n10896_), .A1(new_n6851_), .B0(new_n10900_), .Y(new_n10901_));
  OR3X1    g08465(.A(new_n10901_), .B(new_n10893_), .C(new_n6885_), .Y(new_n10902_));
  OAI22X1  g08466(.A0(new_n10888_), .A1(pi0051), .B0(new_n10488_), .B1(new_n7203_), .Y(new_n10903_));
  OR4X1    g08467(.A(pi0468), .B(pi0332), .C(pi0287), .D(pi0051), .Y(new_n10904_));
  OAI21X1  g08468(.A0(new_n10904_), .A1(new_n5203_), .B0(new_n6851_), .Y(new_n10905_));
  NAND2X1  g08469(.A(new_n10523_), .B(pi0180), .Y(new_n10906_));
  NOR2X1   g08470(.A(new_n10890_), .B(new_n6851_), .Y(new_n10907_));
  AOI21X1  g08471(.A0(new_n10907_), .A1(new_n10906_), .B0(pi0193), .Y(new_n10908_));
  OAI21X1  g08472(.A0(new_n10905_), .A1(new_n10903_), .B0(new_n10908_), .Y(new_n10909_));
  AND2X1   g08473(.A(new_n10909_), .B(new_n2933_), .Y(new_n10910_));
  AOI22X1  g08474(.A0(new_n10910_), .A1(new_n10902_), .B0(new_n10885_), .B1(new_n10875_), .Y(new_n10911_));
  NOR4X1   g08475(.A(new_n10367_), .B(new_n10365_), .C(new_n7187_), .D(new_n5881_), .Y(new_n10912_));
  NOR2X1   g08476(.A(new_n10912_), .B(new_n10342_), .Y(new_n10913_));
  MX2X1    g08477(.A(new_n10913_), .B(new_n10890_), .S0(new_n2933_), .Y(new_n10914_));
  NOR2X1   g08478(.A(new_n10914_), .B(pi0232), .Y(new_n10915_));
  NOR2X1   g08479(.A(new_n10915_), .B(new_n2939_), .Y(new_n10916_));
  OAI21X1  g08480(.A0(new_n10911_), .A1(new_n5215_), .B0(new_n10916_), .Y(new_n10917_));
  OAI21X1  g08481(.A0(new_n10383_), .A1(pi0232), .B0(new_n2939_), .Y(new_n10918_));
  AND2X1   g08482(.A(new_n10918_), .B(new_n2979_), .Y(new_n10919_));
  AOI22X1  g08483(.A0(new_n10919_), .A1(new_n10917_), .B0(new_n10802_), .B1(new_n10874_), .Y(new_n10920_));
  NAND2X1  g08484(.A(new_n10804_), .B(new_n10540_), .Y(new_n10921_));
  AOI21X1  g08485(.A0(new_n10920_), .A1(new_n10873_), .B0(new_n10921_), .Y(new_n10922_));
  AND2X1   g08486(.A(new_n10807_), .B(new_n10663_), .Y(new_n10923_));
  OAI21X1  g08487(.A0(new_n10801_), .A1(new_n10545_), .B0(new_n10923_), .Y(new_n10924_));
  OAI21X1  g08488(.A0(new_n10924_), .A1(new_n10922_), .B0(new_n6489_), .Y(new_n10925_));
  OAI21X1  g08489(.A0(new_n10925_), .A1(new_n10810_), .B0(new_n10669_), .Y(po0282));
  NAND2X1  g08490(.A(new_n10689_), .B(new_n2924_), .Y(new_n10927_));
  AOI21X1  g08491(.A0(new_n10691_), .A1(pi0153), .B0(new_n9968_), .Y(new_n10928_));
  OAI21X1  g08492(.A0(new_n10685_), .A1(new_n2924_), .B0(new_n9968_), .Y(new_n10929_));
  AOI21X1  g08493(.A0(new_n10683_), .A1(new_n2924_), .B0(new_n10929_), .Y(new_n10930_));
  AOI21X1  g08494(.A0(new_n10928_), .A1(new_n10927_), .B0(new_n10930_), .Y(new_n10931_));
  AND3X1   g08495(.A(new_n5023_), .B(pi0153), .C(pi0051), .Y(new_n10932_));
  OR2X1    g08496(.A(new_n10932_), .B(pi0166), .Y(new_n10933_));
  AOI21X1  g08497(.A0(new_n10679_), .A1(new_n9968_), .B0(new_n10933_), .Y(new_n10934_));
  OAI21X1  g08498(.A0(new_n10695_), .A1(new_n9968_), .B0(new_n10934_), .Y(new_n10935_));
  OAI21X1  g08499(.A0(new_n10931_), .A1(new_n4459_), .B0(new_n10935_), .Y(new_n10936_));
  AND2X1   g08500(.A(new_n10936_), .B(new_n7408_), .Y(new_n10937_));
  MX2X1    g08501(.A(new_n10694_), .B(new_n10689_), .S0(pi0189), .Y(new_n10938_));
  NAND2X1  g08502(.A(new_n10938_), .B(pi0178), .Y(new_n10939_));
  NOR2X1   g08503(.A(new_n10679_), .B(pi0189), .Y(new_n10940_));
  OAI21X1  g08504(.A0(new_n10683_), .A1(new_n7872_), .B0(new_n6801_), .Y(new_n10941_));
  OR2X1    g08505(.A(new_n10941_), .B(new_n10940_), .Y(new_n10942_));
  AOI21X1  g08506(.A0(new_n10942_), .A1(new_n10939_), .B0(new_n5204_), .Y(new_n10943_));
  OAI21X1  g08507(.A0(new_n10699_), .A1(pi0189), .B0(pi0178), .Y(new_n10944_));
  AOI21X1  g08508(.A0(new_n10698_), .A1(pi0189), .B0(new_n10944_), .Y(new_n10945_));
  OAI21X1  g08509(.A0(new_n10412_), .A1(new_n7872_), .B0(new_n6801_), .Y(new_n10946_));
  OAI21X1  g08510(.A0(new_n10677_), .A1(new_n10716_), .B0(new_n7872_), .Y(new_n10947_));
  NOR2X1   g08511(.A(new_n10946_), .B(new_n10387_), .Y(new_n10948_));
  AOI21X1  g08512(.A0(new_n10948_), .A1(new_n10947_), .B0(pi0181), .Y(new_n10949_));
  OAI21X1  g08513(.A0(new_n10946_), .A1(new_n10718_), .B0(new_n10949_), .Y(new_n10950_));
  OAI21X1  g08514(.A0(new_n10950_), .A1(new_n10945_), .B0(new_n8716_), .Y(new_n10951_));
  OAI21X1  g08515(.A0(new_n10707_), .A1(pi0166), .B0(pi0153), .Y(new_n10952_));
  AOI21X1  g08516(.A0(new_n10731_), .A1(pi0166), .B0(new_n10952_), .Y(new_n10953_));
  NAND2X1  g08517(.A(new_n10698_), .B(pi0166), .Y(new_n10954_));
  OAI21X1  g08518(.A0(new_n10677_), .A1(new_n10438_), .B0(new_n4459_), .Y(new_n10955_));
  AND2X1   g08519(.A(new_n10955_), .B(new_n2924_), .Y(new_n10956_));
  AOI21X1  g08520(.A0(new_n10956_), .A1(new_n10954_), .B0(new_n10953_), .Y(new_n10957_));
  OR2X1    g08521(.A(new_n10932_), .B(pi0157), .Y(new_n10958_));
  AOI21X1  g08522(.A0(new_n10411_), .A1(pi0166), .B0(new_n10958_), .Y(new_n10959_));
  OAI21X1  g08523(.A0(new_n10717_), .A1(pi0166), .B0(new_n10959_), .Y(new_n10960_));
  OAI21X1  g08524(.A0(new_n10957_), .A1(new_n9968_), .B0(new_n10960_), .Y(new_n10961_));
  AND2X1   g08525(.A(new_n10416_), .B(new_n10412_), .Y(new_n10962_));
  AND2X1   g08526(.A(new_n10830_), .B(new_n7872_), .Y(new_n10963_));
  NOR3X1   g08527(.A(new_n10963_), .B(new_n10682_), .C(new_n10962_), .Y(new_n10964_));
  OAI21X1  g08528(.A0(new_n10695_), .A1(pi0189), .B0(pi0178), .Y(new_n10965_));
  NOR4X1   g08529(.A(new_n10396_), .B(new_n10411_), .C(new_n10387_), .D(new_n7872_), .Y(new_n10966_));
  NOR3X1   g08530(.A(new_n10679_), .B(new_n10387_), .C(pi0189), .Y(new_n10967_));
  OAI21X1  g08531(.A0(new_n10967_), .A1(new_n10966_), .B0(new_n6801_), .Y(new_n10968_));
  AND2X1   g08532(.A(new_n10968_), .B(pi0181), .Y(new_n10969_));
  OAI21X1  g08533(.A0(new_n10965_), .A1(new_n10964_), .B0(new_n10969_), .Y(new_n10970_));
  AOI21X1  g08534(.A0(new_n10706_), .A1(new_n7872_), .B0(new_n6801_), .Y(new_n10971_));
  OAI21X1  g08535(.A0(new_n10702_), .A1(new_n7872_), .B0(new_n10971_), .Y(new_n10972_));
  AOI21X1  g08536(.A0(new_n10972_), .A1(new_n10949_), .B0(new_n8897_), .Y(new_n10973_));
  AOI22X1  g08537(.A0(new_n10973_), .A1(new_n10970_), .B0(new_n10961_), .B1(new_n7378_), .Y(new_n10974_));
  OAI21X1  g08538(.A0(new_n10951_), .A1(new_n10943_), .B0(new_n10974_), .Y(new_n10975_));
  OAI21X1  g08539(.A0(new_n10975_), .A1(new_n10937_), .B0(pi0232), .Y(new_n10976_));
  NOR3X1   g08540(.A(new_n10334_), .B(pi0132), .C(pi0126), .Y(new_n10977_));
  OR3X1    g08541(.A(pi0133), .B(pi0125), .C(pi0121), .Y(new_n10978_));
  XOR2X1   g08542(.A(new_n10978_), .B(pi0126), .Y(new_n10979_));
  NOR2X1   g08543(.A(new_n10979_), .B(new_n10977_), .Y(new_n10980_));
  AOI21X1  g08544(.A0(new_n10779_), .A1(pi0189), .B0(pi0182), .Y(new_n10981_));
  OAI21X1  g08545(.A0(new_n10778_), .A1(pi0189), .B0(new_n10981_), .Y(new_n10982_));
  NOR2X1   g08546(.A(new_n10982_), .B(new_n10387_), .Y(new_n10983_));
  OAI21X1  g08547(.A0(new_n10764_), .A1(pi0189), .B0(pi0182), .Y(new_n10984_));
  AOI21X1  g08548(.A0(new_n10761_), .A1(pi0189), .B0(new_n10984_), .Y(new_n10985_));
  OAI21X1  g08549(.A0(new_n10985_), .A1(new_n10983_), .B0(new_n8743_), .Y(new_n10986_));
  INVX1    g08550(.A(new_n10594_), .Y(new_n10987_));
  AOI21X1  g08551(.A0(new_n10503_), .A1(new_n4459_), .B0(pi0153), .Y(new_n10988_));
  OAI21X1  g08552(.A0(new_n10987_), .A1(new_n4459_), .B0(new_n10988_), .Y(new_n10989_));
  OAI21X1  g08553(.A0(new_n10757_), .A1(new_n10387_), .B0(pi0166), .Y(new_n10990_));
  AOI21X1  g08554(.A0(new_n10785_), .A1(new_n4459_), .B0(new_n2924_), .Y(new_n10991_));
  AOI21X1  g08555(.A0(new_n10991_), .A1(new_n10990_), .B0(new_n8850_), .Y(new_n10992_));
  AOI21X1  g08556(.A0(new_n10992_), .A1(new_n10989_), .B0(new_n2438_), .Y(new_n10993_));
  MX2X1    g08557(.A(new_n10751_), .B(new_n10749_), .S0(new_n4459_), .Y(new_n10994_));
  OR2X1    g08558(.A(pi0153), .B(new_n2534_), .Y(new_n10995_));
  AOI21X1  g08559(.A0(new_n10995_), .A1(new_n10994_), .B0(pi0216), .Y(new_n10996_));
  OR3X1    g08560(.A(new_n10996_), .B(new_n10993_), .C(new_n5221_), .Y(new_n10997_));
  NOR2X1   g08561(.A(new_n10442_), .B(pi0051), .Y(new_n10998_));
  AOI21X1  g08562(.A0(new_n10455_), .A1(new_n8677_), .B0(pi0051), .Y(new_n10999_));
  NOR2X1   g08563(.A(new_n10999_), .B(new_n10932_), .Y(new_n11000_));
  NOR2X1   g08564(.A(new_n11000_), .B(new_n10998_), .Y(new_n11001_));
  OAI21X1  g08565(.A0(new_n2438_), .A1(pi0160), .B0(new_n5220_), .Y(new_n11002_));
  AOI21X1  g08566(.A0(new_n11002_), .A1(new_n11001_), .B0(new_n2933_), .Y(new_n11003_));
  AOI21X1  g08567(.A0(new_n10773_), .A1(pi0189), .B0(new_n5205_), .Y(new_n11004_));
  OAI21X1  g08568(.A0(new_n10771_), .A1(pi0189), .B0(new_n11004_), .Y(new_n11005_));
  AOI21X1  g08569(.A0(new_n11005_), .A1(new_n10982_), .B0(new_n8717_), .Y(new_n11006_));
  AOI21X1  g08570(.A0(new_n11003_), .A1(new_n10997_), .B0(new_n11006_), .Y(new_n11007_));
  AOI21X1  g08571(.A0(new_n11007_), .A1(new_n10986_), .B0(new_n5215_), .Y(new_n11008_));
  OAI21X1  g08572(.A0(new_n11008_), .A1(new_n10746_), .B0(new_n10980_), .Y(new_n11009_));
  AOI21X1  g08573(.A0(new_n10976_), .A1(new_n10796_), .B0(new_n11009_), .Y(new_n11010_));
  AOI22X1  g08574(.A0(new_n10564_), .A1(new_n7872_), .B0(new_n10846_), .B1(new_n7873_), .Y(new_n11011_));
  OR2X1    g08575(.A(new_n11011_), .B(pi0178), .Y(new_n11012_));
  NAND2X1  g08576(.A(new_n10833_), .B(pi0189), .Y(new_n11013_));
  NOR3X1   g08577(.A(new_n10396_), .B(new_n10384_), .C(pi0189), .Y(new_n11014_));
  AOI21X1  g08578(.A0(new_n11014_), .A1(new_n10963_), .B0(new_n6801_), .Y(new_n11015_));
  AOI21X1  g08579(.A0(new_n11015_), .A1(new_n11013_), .B0(pi0181), .Y(new_n11016_));
  OAI21X1  g08580(.A0(new_n10819_), .A1(new_n7872_), .B0(new_n6801_), .Y(new_n11017_));
  AOI21X1  g08581(.A0(new_n10963_), .A1(new_n10850_), .B0(new_n11017_), .Y(new_n11018_));
  AND2X1   g08582(.A(new_n10434_), .B(pi0189), .Y(new_n11019_));
  NOR3X1   g08583(.A(new_n11019_), .B(new_n10963_), .C(new_n6801_), .Y(new_n11020_));
  OR2X1    g08584(.A(new_n11020_), .B(new_n5204_), .Y(new_n11021_));
  OAI21X1  g08585(.A0(new_n11021_), .A1(new_n11018_), .B0(new_n8716_), .Y(new_n11022_));
  AOI21X1  g08586(.A0(new_n11016_), .A1(new_n11012_), .B0(new_n11022_), .Y(new_n11023_));
  AOI21X1  g08587(.A0(new_n10812_), .A1(new_n10811_), .B0(pi0166), .Y(new_n11024_));
  OAI21X1  g08588(.A0(new_n10816_), .A1(new_n4459_), .B0(pi0153), .Y(new_n11025_));
  NOR3X1   g08589(.A(new_n10416_), .B(new_n5048_), .C(pi0166), .Y(new_n11026_));
  OAI21X1  g08590(.A0(new_n10383_), .A1(new_n7717_), .B0(new_n2924_), .Y(new_n11027_));
  OAI22X1  g08591(.A0(new_n11027_), .A1(new_n11026_), .B0(new_n11025_), .B1(new_n11024_), .Y(new_n11028_));
  AOI21X1  g08592(.A0(new_n10397_), .A1(new_n10811_), .B0(pi0166), .Y(new_n11029_));
  AOI22X1  g08593(.A0(new_n10859_), .A1(pi0166), .B0(new_n7717_), .B1(pi0051), .Y(new_n11030_));
  AND2X1   g08594(.A(pi0166), .B(pi0153), .Y(new_n11031_));
  AOI21X1  g08595(.A0(new_n11031_), .A1(new_n10862_), .B0(new_n9968_), .Y(new_n11032_));
  OAI21X1  g08596(.A0(new_n11030_), .A1(pi0153), .B0(new_n11032_), .Y(new_n11033_));
  OAI21X1  g08597(.A0(new_n11033_), .A1(new_n11029_), .B0(new_n7378_), .Y(new_n11034_));
  AOI21X1  g08598(.A0(new_n11028_), .A1(new_n9968_), .B0(new_n11034_), .Y(new_n11035_));
  NAND3X1  g08599(.A(new_n10812_), .B(new_n10811_), .C(new_n7872_), .Y(new_n11036_));
  AOI21X1  g08600(.A0(new_n10816_), .A1(pi0189), .B0(pi0178), .Y(new_n11037_));
  NAND2X1  g08601(.A(new_n11037_), .B(new_n11036_), .Y(new_n11038_));
  NOR2X1   g08602(.A(new_n11014_), .B(new_n6801_), .Y(new_n11039_));
  OR2X1    g08603(.A(new_n10862_), .B(new_n7872_), .Y(new_n11040_));
  AOI21X1  g08604(.A0(new_n11040_), .A1(new_n11039_), .B0(pi0181), .Y(new_n11041_));
  OAI21X1  g08605(.A0(new_n10445_), .A1(new_n7872_), .B0(new_n6801_), .Y(new_n11042_));
  AOI21X1  g08606(.A0(new_n10850_), .A1(new_n7872_), .B0(new_n11042_), .Y(new_n11043_));
  NOR2X1   g08607(.A(new_n10340_), .B(pi0051), .Y(new_n11044_));
  AND3X1   g08608(.A(new_n11044_), .B(new_n8731_), .C(pi0178), .Y(new_n11045_));
  OR3X1    g08609(.A(new_n11045_), .B(new_n10384_), .C(new_n5204_), .Y(new_n11046_));
  OAI21X1  g08610(.A0(new_n11046_), .A1(new_n11043_), .B0(new_n8743_), .Y(new_n11047_));
  AOI21X1  g08611(.A0(new_n11041_), .A1(new_n11038_), .B0(new_n11047_), .Y(new_n11048_));
  OAI21X1  g08612(.A0(new_n10430_), .A1(new_n10384_), .B0(new_n4459_), .Y(new_n11049_));
  OAI21X1  g08613(.A0(new_n10445_), .A1(new_n10384_), .B0(new_n11031_), .Y(new_n11050_));
  OAI22X1  g08614(.A0(new_n10818_), .A1(new_n4459_), .B0(new_n8677_), .B1(new_n2534_), .Y(new_n11051_));
  AOI21X1  g08615(.A0(new_n11051_), .A1(new_n2924_), .B0(pi0157), .Y(new_n11052_));
  AND2X1   g08616(.A(new_n11052_), .B(new_n11050_), .Y(new_n11053_));
  OAI22X1  g08617(.A0(new_n10499_), .A1(new_n4459_), .B0(new_n10383_), .B1(new_n5023_), .Y(new_n11054_));
  AND2X1   g08618(.A(new_n11054_), .B(pi0153), .Y(new_n11055_));
  OAI21X1  g08619(.A0(new_n11000_), .A1(new_n10998_), .B0(new_n2924_), .Y(new_n11056_));
  OAI21X1  g08620(.A0(new_n11056_), .A1(new_n10434_), .B0(pi0157), .Y(new_n11057_));
  OAI21X1  g08621(.A0(new_n11057_), .A1(new_n11055_), .B0(new_n7408_), .Y(new_n11058_));
  AOI21X1  g08622(.A0(new_n11053_), .A1(new_n11049_), .B0(new_n11058_), .Y(new_n11059_));
  OR4X1    g08623(.A(new_n11059_), .B(new_n11048_), .C(new_n11035_), .D(new_n11023_), .Y(new_n11060_));
  AOI21X1  g08624(.A0(new_n11060_), .A1(pi0232), .B0(new_n10918_), .Y(new_n11061_));
  INVX1    g08625(.A(new_n10916_), .Y(new_n11062_));
  INVX1    g08626(.A(new_n10980_), .Y(new_n11063_));
  MX2X1    g08627(.A(new_n10523_), .B(new_n10522_), .S0(new_n4459_), .Y(new_n11064_));
  NOR3X1   g08628(.A(new_n11064_), .B(new_n10932_), .C(new_n8850_), .Y(new_n11065_));
  OAI22X1  g08629(.A0(new_n10750_), .A1(pi0166), .B0(new_n10482_), .B1(new_n7717_), .Y(new_n11066_));
  OAI21X1  g08630(.A0(new_n10878_), .A1(new_n4459_), .B0(pi0153), .Y(new_n11067_));
  AOI21X1  g08631(.A0(new_n10484_), .A1(new_n4459_), .B0(new_n11067_), .Y(new_n11068_));
  AOI21X1  g08632(.A0(new_n11066_), .A1(new_n2924_), .B0(new_n11068_), .Y(new_n11069_));
  OAI21X1  g08633(.A0(new_n11069_), .A1(pi0160), .B0(new_n6856_), .Y(new_n11070_));
  OAI21X1  g08634(.A0(new_n10999_), .A1(new_n10932_), .B0(new_n7187_), .Y(new_n11071_));
  AND2X1   g08635(.A(new_n11071_), .B(pi0299), .Y(new_n11072_));
  OAI21X1  g08636(.A0(new_n11070_), .A1(new_n11065_), .B0(new_n11072_), .Y(new_n11073_));
  INVX1    g08637(.A(new_n10523_), .Y(new_n11074_));
  NOR2X1   g08638(.A(new_n10890_), .B(new_n7872_), .Y(new_n11075_));
  OAI21X1  g08639(.A0(new_n11074_), .A1(new_n5205_), .B0(new_n11075_), .Y(new_n11076_));
  OAI21X1  g08640(.A0(new_n10904_), .A1(new_n5205_), .B0(new_n7872_), .Y(new_n11077_));
  OAI21X1  g08641(.A0(new_n11077_), .A1(new_n10903_), .B0(new_n11076_), .Y(new_n11078_));
  OAI21X1  g08642(.A0(new_n10891_), .A1(new_n7872_), .B0(new_n5205_), .Y(new_n11079_));
  AOI21X1  g08643(.A0(new_n10889_), .A1(new_n7872_), .B0(new_n11079_), .Y(new_n11080_));
  OAI21X1  g08644(.A0(new_n10899_), .A1(new_n7872_), .B0(pi0182), .Y(new_n11081_));
  AOI21X1  g08645(.A0(new_n10896_), .A1(new_n7872_), .B0(new_n11081_), .Y(new_n11082_));
  OR2X1    g08646(.A(new_n11082_), .B(new_n11080_), .Y(new_n11083_));
  AOI22X1  g08647(.A0(new_n11083_), .A1(new_n8743_), .B0(new_n11078_), .B1(new_n8716_), .Y(new_n11084_));
  AOI21X1  g08648(.A0(new_n11084_), .A1(new_n11073_), .B0(new_n5215_), .Y(new_n11085_));
  OAI21X1  g08649(.A0(new_n11085_), .A1(new_n11062_), .B0(new_n11063_), .Y(new_n11086_));
  OAI21X1  g08650(.A0(new_n11086_), .A1(new_n11061_), .B0(new_n3251_), .Y(new_n11087_));
  OAI21X1  g08651(.A0(new_n11000_), .A1(new_n10998_), .B0(pi0299), .Y(new_n11088_));
  AOI21X1  g08652(.A0(new_n10387_), .A1(pi0175), .B0(pi0299), .Y(new_n11089_));
  OAI21X1  g08653(.A0(new_n10499_), .A1(pi0189), .B0(new_n11089_), .Y(new_n11090_));
  AND3X1   g08654(.A(new_n11090_), .B(new_n11088_), .C(pi0232), .Y(new_n11091_));
  NOR3X1   g08655(.A(new_n10980_), .B(new_n10342_), .C(new_n3251_), .Y(new_n11092_));
  OR2X1    g08656(.A(new_n11092_), .B(new_n10539_), .Y(new_n11093_));
  AOI21X1  g08657(.A0(new_n11091_), .A1(new_n3252_), .B0(new_n11093_), .Y(new_n11094_));
  OAI21X1  g08658(.A0(new_n11087_), .A1(new_n11010_), .B0(new_n11094_), .Y(new_n11095_));
  MX2X1    g08659(.A(pi0185), .B(pi0150), .S0(pi0299), .Y(new_n11096_));
  AND3X1   g08660(.A(new_n11096_), .B(new_n5023_), .C(pi0232), .Y(new_n11097_));
  OAI22X1  g08661(.A0(new_n11097_), .A1(new_n3131_), .B0(new_n11091_), .B1(new_n10613_), .Y(new_n11098_));
  AND3X1   g08662(.A(new_n10340_), .B(new_n3131_), .C(new_n2534_), .Y(new_n11099_));
  OAI21X1  g08663(.A0(new_n10979_), .A1(new_n10977_), .B0(new_n11099_), .Y(new_n11100_));
  AOI21X1  g08664(.A0(new_n11100_), .A1(new_n11098_), .B0(po1038), .Y(new_n11101_));
  INVX1    g08665(.A(new_n10998_), .Y(new_n11102_));
  AOI21X1  g08666(.A0(new_n11102_), .A1(pi0232), .B0(new_n11063_), .Y(new_n11103_));
  OAI22X1  g08667(.A0(new_n10999_), .A1(new_n10932_), .B0(new_n10341_), .B1(pi0232), .Y(new_n11104_));
  OAI21X1  g08668(.A0(new_n11104_), .A1(new_n11103_), .B0(new_n3131_), .Y(new_n11105_));
  AOI21X1  g08669(.A0(new_n9951_), .A1(pi0087), .B0(new_n6489_), .Y(new_n11106_));
  AOI22X1  g08670(.A0(new_n11106_), .A1(new_n11105_), .B0(new_n11101_), .B1(new_n11095_), .Y(po0283));
  NOR4X1   g08671(.A(new_n3115_), .B(new_n2985_), .C(new_n2536_), .D(new_n5083_), .Y(new_n11108_));
  AOI21X1  g08672(.A0(new_n4986_), .A1(pi0129), .B0(new_n2979_), .Y(new_n11109_));
  AOI21X1  g08673(.A0(new_n2833_), .A1(pi0093), .B0(new_n2507_), .Y(new_n11110_));
  INVX1    g08674(.A(new_n2545_), .Y(new_n11111_));
  OR3X1    g08675(.A(new_n2655_), .B(pi0102), .C(pi0081), .Y(new_n11112_));
  AOI21X1  g08676(.A0(new_n11112_), .A1(new_n2583_), .B0(new_n2558_), .Y(new_n11113_));
  OAI21X1  g08677(.A0(new_n11113_), .A1(new_n2666_), .B0(new_n2578_), .Y(new_n11114_));
  AOI21X1  g08678(.A0(new_n11114_), .A1(new_n2670_), .B0(new_n2729_), .Y(new_n11115_));
  NOR2X1   g08679(.A(new_n11115_), .B(new_n2575_), .Y(new_n11116_));
  OAI21X1  g08680(.A0(new_n11116_), .A1(pi0086), .B0(new_n2574_), .Y(new_n11117_));
  AOI21X1  g08681(.A0(new_n11117_), .A1(new_n7656_), .B0(new_n2565_), .Y(new_n11118_));
  OAI21X1  g08682(.A0(new_n11118_), .A1(pi0108), .B0(new_n2563_), .Y(new_n11119_));
  AOI21X1  g08683(.A0(new_n11119_), .A1(new_n2678_), .B0(new_n2557_), .Y(new_n11120_));
  OAI21X1  g08684(.A0(new_n11120_), .A1(new_n2556_), .B0(new_n2554_), .Y(new_n11121_));
  OR2X1    g08685(.A(new_n11121_), .B(new_n5912_), .Y(new_n11122_));
  AND2X1   g08686(.A(new_n11117_), .B(new_n2571_), .Y(new_n11123_));
  OAI21X1  g08687(.A0(new_n11123_), .A1(new_n2565_), .B0(new_n2837_), .Y(new_n11124_));
  AOI21X1  g08688(.A0(new_n11124_), .A1(new_n2563_), .B0(new_n5118_), .Y(new_n11125_));
  OAI21X1  g08689(.A0(new_n11125_), .A1(new_n2557_), .B0(new_n2555_), .Y(new_n11126_));
  NAND3X1  g08690(.A(new_n11126_), .B(new_n5912_), .C(new_n2554_), .Y(new_n11127_));
  NOR4X1   g08691(.A(new_n5920_), .B(new_n5082_), .C(new_n3035_), .D(new_n7779_), .Y(new_n11128_));
  AND3X1   g08692(.A(new_n11128_), .B(new_n11127_), .C(new_n11122_), .Y(new_n11129_));
  OR2X1    g08693(.A(new_n11121_), .B(pi0127), .Y(new_n11130_));
  AND3X1   g08694(.A(new_n11126_), .B(new_n2554_), .C(pi0127), .Y(new_n11131_));
  NOR2X1   g08695(.A(new_n11131_), .B(new_n11128_), .Y(new_n11132_));
  AOI21X1  g08696(.A0(new_n11132_), .A1(new_n11130_), .B0(new_n11129_), .Y(new_n11133_));
  OAI21X1  g08697(.A0(new_n11133_), .A1(new_n11111_), .B0(new_n2835_), .Y(new_n11134_));
  NAND2X1  g08698(.A(new_n11134_), .B(new_n2524_), .Y(new_n11135_));
  AOI21X1  g08699(.A0(new_n11135_), .A1(new_n11110_), .B0(pi0070), .Y(new_n11136_));
  OAI21X1  g08700(.A0(new_n11136_), .A1(new_n2848_), .B0(new_n2534_), .Y(new_n11137_));
  AND2X1   g08701(.A(new_n11137_), .B(new_n2537_), .Y(new_n11138_));
  OAI21X1  g08702(.A0(new_n11138_), .A1(new_n2853_), .B0(new_n2532_), .Y(new_n11139_));
  AOI21X1  g08703(.A0(new_n11139_), .A1(new_n2695_), .B0(new_n3178_), .Y(new_n11140_));
  NOR3X1   g08704(.A(new_n2696_), .B(new_n5083_), .C(pi0039), .Y(new_n11141_));
  OAI21X1  g08705(.A0(new_n11140_), .A1(pi0095), .B0(new_n11141_), .Y(new_n11142_));
  AOI21X1  g08706(.A0(new_n6726_), .A1(pi0039), .B0(pi0038), .Y(new_n11143_));
  AOI21X1  g08707(.A0(new_n11143_), .A1(new_n11142_), .B0(new_n11109_), .Y(new_n11144_));
  OAI21X1  g08708(.A0(new_n6777_), .A1(new_n3064_), .B0(new_n6726_), .Y(new_n11145_));
  AOI21X1  g08709(.A0(new_n11145_), .A1(new_n7156_), .B0(pi0075), .Y(new_n11146_));
  OAI21X1  g08710(.A0(new_n11144_), .A1(new_n7156_), .B0(new_n11146_), .Y(new_n11147_));
  NAND3X1  g08711(.A(new_n5779_), .B(pi0129), .C(pi0075), .Y(new_n11148_));
  AND2X1   g08712(.A(new_n11148_), .B(new_n3079_), .Y(new_n11149_));
  AND2X1   g08713(.A(new_n5784_), .B(new_n3091_), .Y(new_n11150_));
  OAI21X1  g08714(.A0(pi0129), .A1(new_n3079_), .B0(new_n11150_), .Y(new_n11151_));
  AOI21X1  g08715(.A0(new_n11149_), .A1(new_n11147_), .B0(new_n11151_), .Y(new_n11152_));
  AND3X1   g08716(.A(new_n3084_), .B(new_n3070_), .C(pi0054), .Y(new_n11153_));
  INVX1    g08717(.A(new_n11153_), .Y(new_n11154_));
  OAI21X1  g08718(.A0(new_n11154_), .A1(new_n6727_), .B0(new_n4982_), .Y(new_n11155_));
  NAND3X1  g08719(.A(new_n5779_), .B(new_n5299_), .C(pi0129), .Y(new_n11156_));
  AOI21X1  g08720(.A0(new_n11156_), .A1(pi0074), .B0(pi0055), .Y(new_n11157_));
  OAI21X1  g08721(.A0(new_n11155_), .A1(new_n11152_), .B0(new_n11157_), .Y(new_n11158_));
  NOR2X1   g08722(.A(new_n10543_), .B(new_n3107_), .Y(new_n11159_));
  NAND3X1  g08723(.A(new_n11159_), .B(new_n5779_), .C(pi0129), .Y(new_n11160_));
  AOI21X1  g08724(.A0(new_n11160_), .A1(new_n11158_), .B0(pi0056), .Y(new_n11161_));
  XOR2X1   g08725(.A(pi0062), .B(pi0056), .Y(new_n11162_));
  OAI22X1  g08726(.A0(new_n11162_), .A1(new_n11161_), .B0(new_n11108_), .B1(new_n3123_), .Y(new_n11163_));
  AOI21X1  g08727(.A0(new_n11108_), .A1(new_n3123_), .B0(new_n3223_), .Y(new_n11164_));
  OR2X1    g08728(.A(new_n11164_), .B(new_n4973_), .Y(new_n11165_));
  AOI21X1  g08729(.A0(new_n11163_), .A1(new_n3223_), .B0(new_n11165_), .Y(po0284));
  INVX1    g08730(.A(new_n5097_), .Y(new_n11167_));
  NOR2X1   g08731(.A(new_n5814_), .B(new_n4984_), .Y(new_n11168_));
  AOI21X1  g08732(.A0(new_n3387_), .A1(new_n2979_), .B0(new_n4989_), .Y(new_n11169_));
  NOR4X1   g08733(.A(new_n5086_), .B(new_n5075_), .C(new_n2986_), .D(pi0039), .Y(new_n11170_));
  OR2X1    g08734(.A(new_n11170_), .B(pi0087), .Y(new_n11171_));
  OAI21X1  g08735(.A0(new_n11171_), .A1(new_n11169_), .B0(new_n5091_), .Y(new_n11172_));
  NOR4X1   g08736(.A(new_n7783_), .B(new_n5920_), .C(new_n5912_), .D(new_n5082_), .Y(new_n11173_));
  AOI21X1  g08737(.A0(new_n7780_), .A1(new_n6728_), .B0(pi0129), .Y(new_n11174_));
  OR4X1    g08738(.A(new_n11174_), .B(new_n11173_), .C(new_n6779_), .D(new_n2986_), .Y(new_n11175_));
  AND3X1   g08739(.A(new_n11175_), .B(new_n3079_), .C(new_n3091_), .Y(new_n11176_));
  OAI21X1  g08740(.A0(new_n5809_), .A1(new_n3091_), .B0(new_n5784_), .Y(new_n11177_));
  AOI21X1  g08741(.A0(new_n11176_), .A1(new_n11172_), .B0(new_n11177_), .Y(new_n11178_));
  OAI21X1  g08742(.A0(new_n11178_), .A1(new_n7552_), .B0(new_n11168_), .Y(new_n11179_));
  AOI21X1  g08743(.A0(new_n11179_), .A1(new_n3118_), .B0(new_n4980_), .Y(new_n11180_));
  OAI21X1  g08744(.A0(new_n11180_), .A1(pi0062), .B0(new_n11167_), .Y(new_n11181_));
  AOI21X1  g08745(.A0(new_n11181_), .A1(new_n3223_), .B0(new_n4977_), .Y(po0286));
  OAI21X1  g08746(.A0(new_n10914_), .A1(pi0051), .B0(new_n5215_), .Y(new_n11183_));
  AND2X1   g08747(.A(new_n11183_), .B(new_n8169_), .Y(new_n11184_));
  AND2X1   g08748(.A(new_n2933_), .B(pi0191), .Y(new_n11185_));
  NOR2X1   g08749(.A(new_n10903_), .B(pi0051), .Y(new_n11186_));
  INVX1    g08750(.A(new_n11186_), .Y(new_n11187_));
  AND2X1   g08751(.A(new_n10492_), .B(pi0140), .Y(new_n11188_));
  OAI21X1  g08752(.A0(new_n11188_), .A1(new_n11187_), .B0(new_n11185_), .Y(new_n11189_));
  NOR3X1   g08753(.A(new_n10492_), .B(new_n10487_), .C(pi0051), .Y(new_n11190_));
  OAI21X1  g08754(.A0(new_n10523_), .A1(pi0051), .B0(new_n4162_), .Y(new_n11191_));
  AND3X1   g08755(.A(new_n11191_), .B(new_n6856_), .C(pi0162), .Y(new_n11192_));
  OAI21X1  g08756(.A0(new_n11190_), .A1(new_n4162_), .B0(new_n11192_), .Y(new_n11193_));
  AND2X1   g08757(.A(new_n5023_), .B(pi0169), .Y(new_n11194_));
  OAI21X1  g08758(.A0(new_n2985_), .A1(new_n2536_), .B0(new_n11194_), .Y(new_n11195_));
  OAI22X1  g08759(.A0(new_n10482_), .A1(pi0051), .B0(new_n5048_), .B1(new_n4162_), .Y(new_n11196_));
  AND3X1   g08760(.A(new_n11196_), .B(new_n6856_), .C(new_n7306_), .Y(new_n11197_));
  NOR3X1   g08761(.A(new_n10340_), .B(new_n6856_), .C(pi0051), .Y(new_n11198_));
  INVX1    g08762(.A(new_n11198_), .Y(new_n11199_));
  OAI21X1  g08763(.A0(new_n11199_), .A1(new_n11194_), .B0(pi0299), .Y(new_n11200_));
  AOI21X1  g08764(.A0(new_n11197_), .A1(new_n11195_), .B0(new_n11200_), .Y(new_n11201_));
  NOR2X1   g08765(.A(pi0299), .B(pi0191), .Y(new_n11202_));
  INVX1    g08766(.A(new_n10898_), .Y(new_n11203_));
  NOR2X1   g08767(.A(new_n10890_), .B(pi0051), .Y(new_n11204_));
  OAI21X1  g08768(.A0(new_n11203_), .A1(new_n7353_), .B0(new_n11204_), .Y(new_n11205_));
  AOI22X1  g08769(.A0(new_n11205_), .A1(new_n11202_), .B0(new_n11201_), .B1(new_n11193_), .Y(new_n11206_));
  AND2X1   g08770(.A(new_n11206_), .B(new_n11189_), .Y(new_n11207_));
  OAI21X1  g08771(.A0(new_n11207_), .A1(new_n5215_), .B0(new_n11184_), .Y(new_n11208_));
  INVX1    g08772(.A(new_n11044_), .Y(new_n11209_));
  NOR3X1   g08773(.A(new_n6811_), .B(new_n5048_), .C(new_n5215_), .Y(new_n11210_));
  OR3X1    g08774(.A(new_n11210_), .B(new_n11209_), .C(new_n8169_), .Y(new_n11211_));
  AND2X1   g08775(.A(new_n11211_), .B(new_n3007_), .Y(new_n11212_));
  OAI22X1  g08776(.A0(new_n11210_), .A1(new_n11209_), .B0(new_n10442_), .B1(pi0051), .Y(new_n11213_));
  OR2X1    g08777(.A(new_n11213_), .B(new_n3007_), .Y(new_n11214_));
  AND2X1   g08778(.A(new_n11214_), .B(new_n5813_), .Y(new_n11215_));
  OAI21X1  g08779(.A0(new_n10342_), .A1(new_n3007_), .B0(new_n11215_), .Y(new_n11216_));
  AOI21X1  g08780(.A0(new_n11212_), .A1(new_n11208_), .B0(new_n11216_), .Y(new_n11217_));
  AOI22X1  g08781(.A0(new_n11213_), .A1(new_n10544_), .B0(new_n7523_), .B1(pi0087), .Y(new_n11218_));
  INVX1    g08782(.A(pi0130), .Y(new_n11219_));
  INVX1    g08783(.A(pi0132), .Y(new_n11220_));
  NOR4X1   g08784(.A(pi0133), .B(pi0126), .C(pi0125), .D(pi0121), .Y(new_n11221_));
  AOI21X1  g08785(.A0(new_n11221_), .A1(new_n11220_), .B0(new_n11219_), .Y(new_n11222_));
  AND3X1   g08786(.A(new_n11221_), .B(new_n11220_), .C(new_n11219_), .Y(new_n11223_));
  OAI21X1  g08787(.A0(new_n11223_), .A1(new_n11222_), .B0(new_n10334_), .Y(new_n11224_));
  OAI21X1  g08788(.A0(new_n11218_), .A1(new_n11099_), .B0(new_n11224_), .Y(new_n11225_));
  NOR2X1   g08789(.A(new_n10785_), .B(new_n10886_), .Y(new_n11226_));
  MX2X1    g08790(.A(new_n10486_), .B(new_n10482_), .S0(new_n5023_), .Y(new_n11227_));
  MX2X1    g08791(.A(new_n11227_), .B(new_n11226_), .S0(pi0224), .Y(new_n11228_));
  MX2X1    g08792(.A(new_n11228_), .B(new_n10998_), .S0(new_n5248_), .Y(new_n11229_));
  AND2X1   g08793(.A(new_n11229_), .B(pi0140), .Y(new_n11230_));
  MX2X1    g08794(.A(new_n11227_), .B(new_n10998_), .S0(new_n6265_), .Y(new_n11231_));
  INVX1    g08795(.A(new_n11231_), .Y(new_n11232_));
  OAI21X1  g08796(.A0(new_n11232_), .A1(pi0140), .B0(new_n11185_), .Y(new_n11233_));
  OAI22X1  g08797(.A0(new_n11194_), .A1(new_n10486_), .B0(new_n10748_), .B1(new_n4162_), .Y(new_n11234_));
  OR3X1    g08798(.A(new_n10757_), .B(pi0169), .C(pi0051), .Y(new_n11235_));
  NAND2X1  g08799(.A(pi0216), .B(pi0162), .Y(new_n11236_));
  AOI21X1  g08800(.A0(new_n11226_), .A1(pi0169), .B0(new_n11236_), .Y(new_n11237_));
  AOI22X1  g08801(.A0(new_n11237_), .A1(new_n11235_), .B0(new_n11234_), .B1(new_n2438_), .Y(new_n11238_));
  AOI21X1  g08802(.A0(new_n10442_), .A1(pi0169), .B0(pi0051), .Y(new_n11239_));
  AOI21X1  g08803(.A0(pi0216), .A1(new_n7306_), .B0(new_n5221_), .Y(new_n11240_));
  OAI22X1  g08804(.A0(new_n11240_), .A1(new_n11239_), .B0(new_n11238_), .B1(new_n5221_), .Y(new_n11241_));
  AOI21X1  g08805(.A0(new_n10759_), .A1(new_n10485_), .B0(pi0051), .Y(new_n11242_));
  AOI21X1  g08806(.A0(new_n10485_), .A1(new_n6264_), .B0(pi0051), .Y(new_n11243_));
  INVX1    g08807(.A(new_n11243_), .Y(new_n11244_));
  OAI21X1  g08808(.A0(new_n11244_), .A1(pi0140), .B0(new_n11202_), .Y(new_n11245_));
  AOI21X1  g08809(.A0(new_n11242_), .A1(pi0140), .B0(new_n11245_), .Y(new_n11246_));
  AOI21X1  g08810(.A0(new_n11241_), .A1(pi0299), .B0(new_n11246_), .Y(new_n11247_));
  OAI21X1  g08811(.A0(new_n11233_), .A1(new_n11230_), .B0(new_n11247_), .Y(new_n11248_));
  AOI21X1  g08812(.A0(new_n10743_), .A1(new_n10485_), .B0(pi0051), .Y(new_n11249_));
  OAI21X1  g08813(.A0(new_n11249_), .A1(pi0232), .B0(pi0039), .Y(new_n11250_));
  AOI21X1  g08814(.A0(new_n11248_), .A1(pi0232), .B0(new_n11250_), .Y(new_n11251_));
  INVX1    g08815(.A(new_n10962_), .Y(new_n11252_));
  AOI21X1  g08816(.A0(new_n11252_), .A1(new_n5215_), .B0(pi0039), .Y(new_n11253_));
  MX2X1    g08817(.A(new_n11252_), .B(new_n10419_), .S0(new_n5023_), .Y(new_n11254_));
  AOI21X1  g08818(.A0(new_n10962_), .A1(new_n6811_), .B0(new_n5215_), .Y(new_n11255_));
  OAI21X1  g08819(.A0(new_n11254_), .A1(new_n6811_), .B0(new_n11255_), .Y(new_n11256_));
  AOI21X1  g08820(.A0(new_n11256_), .A1(new_n11253_), .B0(new_n11251_), .Y(new_n11257_));
  AOI21X1  g08821(.A0(new_n11213_), .A1(pi0038), .B0(pi0100), .Y(new_n11258_));
  OAI21X1  g08822(.A0(new_n11257_), .A1(pi0038), .B0(new_n11258_), .Y(new_n11259_));
  AND2X1   g08823(.A(new_n11259_), .B(new_n11215_), .Y(new_n11260_));
  OR2X1    g08824(.A(new_n11223_), .B(new_n11222_), .Y(new_n11261_));
  NAND3X1  g08825(.A(new_n11261_), .B(new_n11218_), .C(new_n10334_), .Y(new_n11262_));
  OAI22X1  g08826(.A0(new_n11262_), .A1(new_n11260_), .B0(new_n11225_), .B1(new_n11217_), .Y(new_n11263_));
  AND2X1   g08827(.A(new_n10442_), .B(pi0169), .Y(new_n11264_));
  NOR4X1   g08828(.A(new_n11264_), .B(new_n11224_), .C(pi0087), .D(pi0051), .Y(new_n11265_));
  NAND3X1  g08829(.A(new_n5023_), .B(pi0232), .C(pi0169), .Y(new_n11266_));
  AND3X1   g08830(.A(new_n11266_), .B(new_n11044_), .C(new_n3131_), .Y(new_n11267_));
  OAI22X1  g08831(.A0(new_n7312_), .A1(new_n3131_), .B0(new_n5103_), .B1(pi0057), .Y(new_n11268_));
  NOR3X1   g08832(.A(new_n11268_), .B(new_n11267_), .C(new_n11265_), .Y(new_n11269_));
  AOI21X1  g08833(.A0(new_n11263_), .A1(new_n6489_), .B0(new_n11269_), .Y(po0287));
  OAI21X1  g08834(.A0(new_n5804_), .A1(new_n3007_), .B0(new_n3131_), .Y(new_n11271_));
  AOI21X1  g08835(.A0(new_n10062_), .A1(new_n3007_), .B0(new_n11271_), .Y(new_n11272_));
  OAI21X1  g08836(.A0(new_n11272_), .A1(pi0075), .B0(new_n5781_), .Y(new_n11273_));
  NAND3X1  g08837(.A(new_n6721_), .B(new_n5784_), .C(new_n3091_), .Y(new_n11274_));
  AOI21X1  g08838(.A0(new_n11273_), .A1(new_n3079_), .B0(new_n11274_), .Y(po0288));
  AOI22X1  g08839(.A0(new_n10462_), .A1(new_n9888_), .B0(new_n3347_), .B1(pi0051), .Y(new_n11276_));
  AND2X1   g08840(.A(new_n11276_), .B(new_n10354_), .Y(new_n11277_));
  OR2X1    g08841(.A(new_n10334_), .B(pi0132), .Y(new_n11278_));
  XOR2X1   g08842(.A(new_n11221_), .B(pi0132), .Y(new_n11279_));
  AND2X1   g08843(.A(new_n11279_), .B(new_n11278_), .Y(new_n11280_));
  INVX1    g08844(.A(new_n11280_), .Y(new_n11281_));
  AOI22X1  g08845(.A0(new_n11281_), .A1(new_n10341_), .B0(new_n11277_), .B1(pi0232), .Y(new_n11282_));
  AOI21X1  g08846(.A0(new_n10667_), .A1(pi0164), .B0(new_n6489_), .Y(new_n11283_));
  OAI21X1  g08847(.A0(new_n11282_), .A1(pi0087), .B0(new_n11283_), .Y(new_n11284_));
  AND3X1   g08848(.A(new_n10416_), .B(new_n10412_), .C(pi0151), .Y(new_n11285_));
  OAI21X1  g08849(.A0(new_n10421_), .A1(pi0151), .B0(new_n4308_), .Y(new_n11286_));
  AOI21X1  g08850(.A0(new_n3347_), .A1(pi0051), .B0(new_n4308_), .Y(new_n11287_));
  AOI21X1  g08851(.A0(new_n11287_), .A1(new_n10419_), .B0(new_n5048_), .Y(new_n11288_));
  OAI21X1  g08852(.A0(new_n11286_), .A1(new_n11285_), .B0(new_n11288_), .Y(new_n11289_));
  NOR2X1   g08853(.A(new_n10427_), .B(new_n5023_), .Y(new_n11290_));
  NOR2X1   g08854(.A(new_n11290_), .B(new_n8850_), .Y(new_n11291_));
  NOR3X1   g08855(.A(new_n10426_), .B(new_n5170_), .C(new_n5023_), .Y(new_n11292_));
  OR3X1    g08856(.A(new_n11292_), .B(new_n10430_), .C(new_n10429_), .Y(new_n11293_));
  OR2X1    g08857(.A(new_n10705_), .B(new_n4308_), .Y(new_n11294_));
  OAI21X1  g08858(.A0(new_n11294_), .A1(new_n11290_), .B0(pi0151), .Y(new_n11295_));
  AOI21X1  g08859(.A0(new_n11293_), .A1(new_n4308_), .B0(new_n11295_), .Y(new_n11296_));
  NOR3X1   g08860(.A(new_n10426_), .B(new_n9887_), .C(new_n5170_), .Y(new_n11297_));
  NOR3X1   g08861(.A(new_n10437_), .B(new_n10435_), .C(new_n4308_), .Y(new_n11298_));
  OR2X1    g08862(.A(new_n11298_), .B(pi0151), .Y(new_n11299_));
  OAI21X1  g08863(.A0(new_n11299_), .A1(new_n11297_), .B0(new_n8850_), .Y(new_n11300_));
  OAI21X1  g08864(.A0(new_n11300_), .A1(new_n11296_), .B0(pi0299), .Y(new_n11301_));
  AOI21X1  g08865(.A0(new_n11291_), .A1(new_n11289_), .B0(new_n11301_), .Y(new_n11302_));
  OR2X1    g08866(.A(pi0299), .B(pi0190), .Y(new_n11303_));
  NOR2X1   g08867(.A(new_n10421_), .B(new_n5048_), .Y(new_n11304_));
  OAI21X1  g08868(.A0(new_n10427_), .A1(new_n5023_), .B0(pi0182), .Y(new_n11305_));
  AOI21X1  g08869(.A0(new_n10427_), .A1(new_n5205_), .B0(pi0173), .Y(new_n11306_));
  OAI21X1  g08870(.A0(new_n11305_), .A1(new_n11304_), .B0(new_n11306_), .Y(new_n11307_));
  OAI21X1  g08871(.A0(new_n11292_), .A1(new_n10417_), .B0(pi0182), .Y(new_n11308_));
  AOI21X1  g08872(.A0(new_n11293_), .A1(new_n5205_), .B0(new_n9903_), .Y(new_n11309_));
  NAND2X1  g08873(.A(new_n11309_), .B(new_n11308_), .Y(new_n11310_));
  AOI21X1  g08874(.A0(new_n11310_), .A1(new_n11307_), .B0(new_n11303_), .Y(new_n11311_));
  AND2X1   g08875(.A(new_n2933_), .B(pi0190), .Y(new_n11312_));
  INVX1    g08876(.A(new_n11312_), .Y(new_n11313_));
  NAND2X1  g08877(.A(new_n10380_), .B(pi0182), .Y(new_n11314_));
  OAI21X1  g08878(.A0(pi0173), .A1(new_n2534_), .B0(new_n5023_), .Y(new_n11315_));
  AOI21X1  g08879(.A0(new_n11314_), .A1(new_n10435_), .B0(new_n11315_), .Y(new_n11316_));
  NOR3X1   g08880(.A(new_n11316_), .B(new_n11313_), .C(new_n11292_), .Y(new_n11317_));
  OR4X1    g08881(.A(new_n11317_), .B(new_n11311_), .C(new_n11302_), .D(new_n5215_), .Y(new_n11318_));
  OR3X1    g08882(.A(new_n10426_), .B(new_n5170_), .C(pi0232), .Y(new_n11319_));
  AOI21X1  g08883(.A0(new_n11319_), .A1(new_n11318_), .B0(pi0039), .Y(new_n11320_));
  AOI21X1  g08884(.A0(new_n10503_), .A1(pi0168), .B0(pi0151), .Y(new_n11321_));
  OAI21X1  g08885(.A0(new_n10987_), .A1(pi0168), .B0(new_n11321_), .Y(new_n11322_));
  OAI21X1  g08886(.A0(new_n10757_), .A1(new_n10387_), .B0(new_n4308_), .Y(new_n11323_));
  AOI21X1  g08887(.A0(new_n10785_), .A1(pi0168), .B0(new_n3347_), .Y(new_n11324_));
  AOI21X1  g08888(.A0(new_n11324_), .A1(new_n11323_), .B0(new_n7101_), .Y(new_n11325_));
  AOI21X1  g08889(.A0(new_n11325_), .A1(new_n11322_), .B0(new_n2438_), .Y(new_n11326_));
  OR2X1    g08890(.A(pi0151), .B(new_n2534_), .Y(new_n11327_));
  MX2X1    g08891(.A(new_n10751_), .B(new_n10749_), .S0(pi0168), .Y(new_n11328_));
  AOI21X1  g08892(.A0(new_n11328_), .A1(new_n11327_), .B0(pi0216), .Y(new_n11329_));
  NOR3X1   g08893(.A(new_n11329_), .B(new_n11326_), .C(new_n5221_), .Y(new_n11330_));
  INVX1    g08894(.A(new_n11277_), .Y(new_n11331_));
  AOI21X1  g08895(.A0(pi0216), .A1(new_n7101_), .B0(new_n5221_), .Y(new_n11332_));
  OAI21X1  g08896(.A0(new_n11332_), .A1(new_n11331_), .B0(pi0299), .Y(new_n11333_));
  NOR2X1   g08897(.A(new_n10771_), .B(new_n6802_), .Y(new_n11334_));
  OAI21X1  g08898(.A0(new_n10767_), .A1(pi0183), .B0(new_n9903_), .Y(new_n11335_));
  OAI21X1  g08899(.A0(new_n10749_), .A1(new_n6265_), .B0(new_n6802_), .Y(new_n11336_));
  AND3X1   g08900(.A(new_n11336_), .B(new_n10764_), .C(pi0173), .Y(new_n11337_));
  AOI21X1  g08901(.A0(new_n10777_), .A1(new_n6802_), .B0(new_n11337_), .Y(new_n11338_));
  OAI21X1  g08902(.A0(new_n11335_), .A1(new_n11334_), .B0(new_n11338_), .Y(new_n11339_));
  OR3X1    g08903(.A(new_n10779_), .B(new_n10387_), .C(pi0183), .Y(new_n11340_));
  AND2X1   g08904(.A(new_n11340_), .B(pi0173), .Y(new_n11341_));
  OAI21X1  g08905(.A0(new_n10761_), .A1(new_n6802_), .B0(new_n11341_), .Y(new_n11342_));
  AOI21X1  g08906(.A0(new_n6265_), .A1(new_n6802_), .B0(pi0173), .Y(new_n11343_));
  AOI21X1  g08907(.A0(new_n11343_), .A1(new_n10773_), .B0(new_n11303_), .Y(new_n11344_));
  AOI22X1  g08908(.A0(new_n11344_), .A1(new_n11342_), .B0(new_n11339_), .B1(new_n11312_), .Y(new_n11345_));
  OAI21X1  g08909(.A0(new_n11333_), .A1(new_n11330_), .B0(new_n11345_), .Y(new_n11346_));
  AOI21X1  g08910(.A0(new_n11346_), .A1(pi0232), .B0(new_n10746_), .Y(new_n11347_));
  OAI21X1  g08911(.A0(new_n11347_), .A1(new_n11320_), .B0(new_n3251_), .Y(new_n11348_));
  AND3X1   g08912(.A(new_n5023_), .B(pi0173), .C(pi0051), .Y(new_n11349_));
  NOR2X1   g08913(.A(new_n11349_), .B(pi0299), .Y(new_n11350_));
  OAI21X1  g08914(.A0(new_n10499_), .A1(new_n9900_), .B0(new_n11350_), .Y(new_n11351_));
  OR2X1    g08915(.A(new_n11277_), .B(new_n2933_), .Y(new_n11352_));
  AND3X1   g08916(.A(new_n11352_), .B(new_n11351_), .C(pi0232), .Y(new_n11353_));
  AOI21X1  g08917(.A0(new_n11353_), .A1(new_n3252_), .B0(new_n10539_), .Y(new_n11354_));
  AOI21X1  g08918(.A0(new_n7131_), .A1(pi0087), .B0(new_n11281_), .Y(new_n11355_));
  OAI21X1  g08919(.A0(new_n11353_), .A1(new_n10613_), .B0(new_n11355_), .Y(new_n11356_));
  AOI21X1  g08920(.A0(new_n11354_), .A1(new_n11348_), .B0(new_n11356_), .Y(new_n11357_));
  NOR3X1   g08921(.A(new_n11277_), .B(new_n10341_), .C(new_n2933_), .Y(new_n11358_));
  AOI21X1  g08922(.A0(new_n10878_), .A1(new_n4308_), .B0(new_n3347_), .Y(new_n11359_));
  OAI21X1  g08923(.A0(new_n10484_), .A1(new_n4308_), .B0(new_n11359_), .Y(new_n11360_));
  AOI21X1  g08924(.A0(new_n10483_), .A1(new_n9888_), .B0(pi0151), .Y(new_n11361_));
  OAI21X1  g08925(.A0(new_n10750_), .A1(new_n4308_), .B0(new_n11361_), .Y(new_n11362_));
  AND3X1   g08926(.A(new_n11362_), .B(new_n11360_), .C(new_n7101_), .Y(new_n11363_));
  OAI21X1  g08927(.A0(new_n10757_), .A1(new_n10387_), .B0(new_n11327_), .Y(new_n11364_));
  AOI21X1  g08928(.A0(new_n11364_), .A1(new_n10488_), .B0(new_n4308_), .Y(new_n11365_));
  OAI21X1  g08929(.A0(new_n11276_), .A1(new_n10523_), .B0(new_n4308_), .Y(new_n11366_));
  NAND2X1  g08930(.A(new_n11366_), .B(pi0149), .Y(new_n11367_));
  OAI21X1  g08931(.A0(new_n11367_), .A1(new_n11365_), .B0(new_n6856_), .Y(new_n11368_));
  OAI22X1  g08932(.A0(new_n11368_), .A1(new_n11363_), .B0(new_n11358_), .B1(new_n9493_), .Y(new_n11369_));
  AND2X1   g08933(.A(new_n10889_), .B(new_n6802_), .Y(new_n11370_));
  AND2X1   g08934(.A(new_n10896_), .B(pi0183), .Y(new_n11371_));
  OR2X1    g08935(.A(new_n11371_), .B(new_n9903_), .Y(new_n11372_));
  OAI21X1  g08936(.A0(new_n10904_), .A1(new_n6802_), .B0(new_n9903_), .Y(new_n11373_));
  OAI22X1  g08937(.A0(new_n11373_), .A1(new_n10903_), .B0(new_n11372_), .B1(new_n11370_), .Y(new_n11374_));
  OR3X1    g08938(.A(new_n11349_), .B(new_n11303_), .C(new_n10890_), .Y(new_n11375_));
  AOI21X1  g08939(.A0(new_n10523_), .A1(pi0183), .B0(new_n11375_), .Y(new_n11376_));
  AOI21X1  g08940(.A0(new_n11374_), .A1(new_n11312_), .B0(new_n11376_), .Y(new_n11377_));
  AOI21X1  g08941(.A0(new_n11377_), .A1(new_n11369_), .B0(new_n5215_), .Y(new_n11378_));
  OAI21X1  g08942(.A0(new_n11378_), .A1(new_n10915_), .B0(pi0039), .Y(new_n11379_));
  AOI21X1  g08943(.A0(new_n10382_), .A1(new_n3347_), .B0(pi0168), .Y(new_n11380_));
  OAI21X1  g08944(.A0(new_n10577_), .A1(new_n3347_), .B0(new_n11380_), .Y(new_n11381_));
  OAI21X1  g08945(.A0(new_n10462_), .A1(pi0151), .B0(pi0168), .Y(new_n11382_));
  OAI21X1  g08946(.A0(new_n11382_), .A1(new_n10396_), .B0(new_n11381_), .Y(new_n11383_));
  NOR2X1   g08947(.A(new_n10817_), .B(pi0160), .Y(new_n11384_));
  OAI22X1  g08948(.A0(new_n10499_), .A1(pi0168), .B0(new_n10381_), .B1(new_n5023_), .Y(new_n11385_));
  AOI21X1  g08949(.A0(new_n10380_), .A1(new_n5048_), .B0(new_n10342_), .Y(new_n11386_));
  OR2X1    g08950(.A(new_n11277_), .B(pi0151), .Y(new_n11387_));
  OAI21X1  g08951(.A0(new_n11387_), .A1(new_n11386_), .B0(pi0160), .Y(new_n11388_));
  AOI21X1  g08952(.A0(new_n11385_), .A1(pi0151), .B0(new_n11388_), .Y(new_n11389_));
  OR2X1    g08953(.A(new_n11389_), .B(new_n2933_), .Y(new_n11390_));
  AOI21X1  g08954(.A0(new_n11384_), .A1(new_n11383_), .B0(new_n11390_), .Y(new_n11391_));
  OAI22X1  g08955(.A0(new_n10381_), .A1(new_n5023_), .B0(pi0173), .B1(new_n2534_), .Y(new_n11392_));
  AOI21X1  g08956(.A0(new_n10396_), .A1(new_n5205_), .B0(new_n11392_), .Y(new_n11393_));
  NAND2X1  g08957(.A(new_n11386_), .B(pi0182), .Y(new_n11394_));
  NOR3X1   g08958(.A(new_n11349_), .B(new_n11303_), .C(new_n10381_), .Y(new_n11395_));
  AOI21X1  g08959(.A0(new_n11395_), .A1(new_n11394_), .B0(new_n5215_), .Y(new_n11396_));
  OAI21X1  g08960(.A0(new_n11393_), .A1(new_n11313_), .B0(new_n11396_), .Y(new_n11397_));
  AOI21X1  g08961(.A0(new_n10381_), .A1(new_n5215_), .B0(pi0039), .Y(new_n11398_));
  OAI21X1  g08962(.A0(new_n11397_), .A1(new_n11391_), .B0(new_n11398_), .Y(new_n11399_));
  AND2X1   g08963(.A(new_n11399_), .B(new_n3251_), .Y(new_n11400_));
  AND2X1   g08964(.A(new_n10341_), .B(new_n3252_), .Y(new_n11401_));
  AND2X1   g08965(.A(new_n11353_), .B(new_n3252_), .Y(new_n11402_));
  OR3X1    g08966(.A(new_n11402_), .B(new_n11401_), .C(new_n10539_), .Y(new_n11403_));
  AOI21X1  g08967(.A0(new_n11400_), .A1(new_n11379_), .B0(new_n11403_), .Y(new_n11404_));
  AOI22X1  g08968(.A0(new_n11279_), .A1(new_n11278_), .B0(new_n7131_), .B1(pi0087), .Y(new_n11405_));
  OAI21X1  g08969(.A0(new_n11353_), .A1(new_n10545_), .B0(new_n11405_), .Y(new_n11406_));
  OAI21X1  g08970(.A0(new_n11406_), .A1(new_n11404_), .B0(new_n6489_), .Y(new_n11407_));
  OAI21X1  g08971(.A0(new_n11407_), .A1(new_n11357_), .B0(new_n11284_), .Y(po0289));
  AOI21X1  g08972(.A0(new_n10401_), .A1(new_n5048_), .B0(new_n11304_), .Y(new_n11409_));
  AND2X1   g08973(.A(pi0176), .B(new_n2939_), .Y(new_n11410_));
  OAI21X1  g08974(.A0(new_n10401_), .A1(new_n7143_), .B0(new_n11410_), .Y(new_n11411_));
  AOI21X1  g08975(.A0(new_n11409_), .A1(new_n7143_), .B0(new_n11411_), .Y(new_n11412_));
  AND3X1   g08976(.A(pi0299), .B(pi0232), .C(pi0154), .Y(new_n11413_));
  NOR2X1   g08977(.A(pi0176), .B(pi0039), .Y(new_n11414_));
  OAI21X1  g08978(.A0(new_n11413_), .A1(new_n10401_), .B0(new_n11414_), .Y(new_n11415_));
  AOI21X1  g08979(.A0(new_n11413_), .A1(new_n11409_), .B0(new_n11415_), .Y(new_n11416_));
  INVX1    g08980(.A(new_n10744_), .Y(new_n11417_));
  INVX1    g08981(.A(new_n10772_), .Y(new_n11418_));
  OR2X1    g08982(.A(new_n2437_), .B(pi0216), .Y(new_n11419_));
  NAND2X1  g08983(.A(new_n10492_), .B(pi0197), .Y(new_n11420_));
  NAND2X1  g08984(.A(new_n11420_), .B(new_n11419_), .Y(new_n11421_));
  AOI21X1  g08985(.A0(new_n6265_), .A1(new_n5202_), .B0(pi0299), .Y(new_n11422_));
  AOI22X1  g08986(.A0(new_n11422_), .A1(new_n11418_), .B0(new_n11421_), .B1(new_n5331_), .Y(new_n11423_));
  OAI21X1  g08987(.A0(new_n11423_), .A1(new_n2986_), .B0(pi0232), .Y(new_n11424_));
  AOI21X1  g08988(.A0(new_n11424_), .A1(new_n11417_), .B0(new_n2939_), .Y(new_n11425_));
  OR4X1    g08989(.A(new_n11425_), .B(new_n11416_), .C(new_n11412_), .D(new_n8428_), .Y(new_n11426_));
  AOI21X1  g08990(.A0(new_n10335_), .A1(new_n10660_), .B0(pi0133), .Y(new_n11427_));
  AND2X1   g08991(.A(new_n11427_), .B(new_n3131_), .Y(new_n11428_));
  NOR2X1   g08992(.A(new_n10890_), .B(pi0299), .Y(new_n11429_));
  OAI21X1  g08993(.A0(new_n11074_), .A1(new_n5202_), .B0(new_n11429_), .Y(new_n11430_));
  AOI21X1  g08994(.A0(new_n11420_), .A1(new_n10912_), .B0(new_n10342_), .Y(new_n11431_));
  OR2X1    g08995(.A(new_n11431_), .B(new_n2933_), .Y(new_n11432_));
  AOI21X1  g08996(.A0(new_n11432_), .A1(new_n11430_), .B0(new_n5215_), .Y(new_n11433_));
  OR4X1    g08997(.A(new_n10377_), .B(new_n10371_), .C(new_n7145_), .D(new_n5881_), .Y(new_n11434_));
  AND3X1   g08998(.A(new_n10340_), .B(new_n2534_), .C(new_n2939_), .Y(new_n11435_));
  AOI21X1  g08999(.A0(new_n11435_), .A1(new_n11434_), .B0(pi0038), .Y(new_n11436_));
  OAI21X1  g09000(.A0(new_n11433_), .A1(new_n11062_), .B0(new_n11436_), .Y(new_n11437_));
  AOI21X1  g09001(.A0(new_n11437_), .A1(new_n10362_), .B0(new_n10541_), .Y(new_n11438_));
  AOI21X1  g09002(.A0(new_n10544_), .A1(new_n10342_), .B0(new_n11438_), .Y(new_n11439_));
  MX2X1    g09003(.A(pi0183), .B(pi0149), .S0(pi0299), .Y(new_n11440_));
  AND3X1   g09004(.A(new_n11440_), .B(new_n5023_), .C(pi0232), .Y(new_n11441_));
  OAI22X1  g09005(.A0(new_n11441_), .A1(new_n3131_), .B0(new_n11439_), .B1(new_n11427_), .Y(new_n11442_));
  AOI21X1  g09006(.A0(new_n11428_), .A1(new_n11426_), .B0(new_n11442_), .Y(new_n11443_));
  NOR3X1   g09007(.A(new_n11427_), .B(new_n10342_), .C(pi0087), .Y(new_n11444_));
  NAND4X1  g09008(.A(new_n5023_), .B(pi0232), .C(pi0149), .D(pi0087), .Y(new_n11445_));
  OAI21X1  g09009(.A0(new_n5103_), .A1(pi0057), .B0(new_n11445_), .Y(new_n11446_));
  OAI22X1  g09010(.A0(new_n11446_), .A1(new_n11444_), .B0(new_n11443_), .B1(po1038), .Y(po0290));
  INVX1    g09011(.A(pi0134), .Y(new_n11448_));
  INVX1    g09012(.A(pi0135), .Y(new_n11449_));
  INVX1    g09013(.A(pi0136), .Y(new_n11450_));
  AND3X1   g09014(.A(new_n11223_), .B(new_n11450_), .C(new_n11449_), .Y(new_n11451_));
  NOR2X1   g09015(.A(new_n11451_), .B(new_n11448_), .Y(new_n11452_));
  OR3X1    g09016(.A(new_n6489_), .B(pi0087), .C(pi0051), .Y(new_n11453_));
  NOR4X1   g09017(.A(new_n10340_), .B(pi0468), .C(pi0332), .D(new_n3715_), .Y(new_n11454_));
  AOI21X1  g09018(.A0(new_n11454_), .A1(pi0232), .B0(new_n11453_), .Y(new_n11455_));
  OAI21X1  g09019(.A0(new_n11452_), .A1(new_n10455_), .B0(new_n11455_), .Y(new_n11456_));
  NAND2X1  g09020(.A(pi0186), .B(pi0039), .Y(new_n11457_));
  INVX1    g09021(.A(pi0192), .Y(new_n11458_));
  OR2X1    g09022(.A(pi0299), .B(new_n11458_), .Y(new_n11459_));
  NOR3X1   g09023(.A(new_n10903_), .B(new_n10492_), .C(pi0051), .Y(new_n11460_));
  INVX1    g09024(.A(new_n11204_), .Y(new_n11461_));
  NOR2X1   g09025(.A(pi0299), .B(pi0192), .Y(new_n11462_));
  OAI21X1  g09026(.A0(new_n11461_), .A1(new_n10898_), .B0(new_n11462_), .Y(new_n11463_));
  OAI21X1  g09027(.A0(new_n11460_), .A1(new_n11459_), .B0(new_n11463_), .Y(new_n11464_));
  AND2X1   g09028(.A(new_n5023_), .B(pi0171), .Y(new_n11465_));
  INVX1    g09029(.A(new_n11465_), .Y(new_n11466_));
  AOI21X1  g09030(.A0(new_n11466_), .A1(new_n11198_), .B0(new_n2933_), .Y(new_n11467_));
  INVX1    g09031(.A(new_n11467_), .Y(new_n11468_));
  NAND3X1  g09032(.A(new_n5023_), .B(new_n2986_), .C(pi0171), .Y(new_n11469_));
  AOI21X1  g09033(.A0(new_n11466_), .A1(new_n10502_), .B0(new_n7187_), .Y(new_n11470_));
  AOI21X1  g09034(.A0(new_n11470_), .A1(new_n11469_), .B0(new_n11468_), .Y(new_n11471_));
  OAI21X1  g09035(.A0(new_n11471_), .A1(new_n11464_), .B0(pi0232), .Y(new_n11472_));
  AOI21X1  g09036(.A0(new_n11472_), .A1(new_n11183_), .B0(new_n11457_), .Y(new_n11473_));
  OR2X1    g09037(.A(pi0186), .B(new_n2939_), .Y(new_n11474_));
  INVX1    g09038(.A(new_n11462_), .Y(new_n11475_));
  OAI22X1  g09039(.A0(new_n11475_), .A1(new_n11204_), .B0(new_n11459_), .B1(new_n11186_), .Y(new_n11476_));
  OAI21X1  g09040(.A0(new_n11476_), .A1(new_n11471_), .B0(pi0232), .Y(new_n11477_));
  AOI21X1  g09041(.A0(new_n11477_), .A1(new_n11183_), .B0(new_n11474_), .Y(new_n11478_));
  MX2X1    g09042(.A(new_n11458_), .B(new_n3715_), .S0(pi0299), .Y(new_n11479_));
  OAI21X1  g09043(.A0(new_n11479_), .A1(new_n6820_), .B0(new_n11044_), .Y(new_n11480_));
  AND2X1   g09044(.A(new_n11480_), .B(new_n2939_), .Y(new_n11481_));
  NOR4X1   g09045(.A(new_n11481_), .B(new_n11478_), .C(new_n11473_), .D(pi0164), .Y(new_n11482_));
  OAI21X1  g09046(.A0(new_n10523_), .A1(pi0051), .B0(new_n3715_), .Y(new_n11483_));
  AND2X1   g09047(.A(new_n11483_), .B(new_n6856_), .Y(new_n11484_));
  OAI21X1  g09048(.A0(new_n11190_), .A1(new_n3715_), .B0(new_n11484_), .Y(new_n11485_));
  AND2X1   g09049(.A(new_n11485_), .B(new_n11467_), .Y(new_n11486_));
  OAI21X1  g09050(.A0(new_n11486_), .A1(new_n11464_), .B0(pi0232), .Y(new_n11487_));
  AOI21X1  g09051(.A0(new_n11487_), .A1(new_n11183_), .B0(new_n11457_), .Y(new_n11488_));
  OAI21X1  g09052(.A0(new_n11486_), .A1(new_n11476_), .B0(pi0232), .Y(new_n11489_));
  AOI21X1  g09053(.A0(new_n11489_), .A1(new_n11183_), .B0(new_n11474_), .Y(new_n11490_));
  NOR4X1   g09054(.A(new_n11490_), .B(new_n11488_), .C(new_n11481_), .D(new_n6826_), .Y(new_n11491_));
  OR3X1    g09055(.A(new_n11491_), .B(new_n11482_), .C(new_n3252_), .Y(new_n11492_));
  AND3X1   g09056(.A(new_n11480_), .B(new_n11102_), .C(new_n3252_), .Y(new_n11493_));
  NOR3X1   g09057(.A(new_n11493_), .B(new_n11401_), .C(new_n10539_), .Y(new_n11494_));
  OAI22X1  g09058(.A0(new_n11480_), .A1(new_n10613_), .B0(new_n11451_), .B1(new_n11448_), .Y(new_n11495_));
  AOI21X1  g09059(.A0(new_n11494_), .A1(new_n11492_), .B0(new_n11495_), .Y(new_n11496_));
  OR2X1    g09060(.A(new_n11493_), .B(new_n10539_), .Y(new_n11497_));
  INVX1    g09061(.A(new_n11250_), .Y(new_n11498_));
  NOR2X1   g09062(.A(new_n11454_), .B(pi0051), .Y(new_n11499_));
  AOI21X1  g09063(.A0(pi0216), .A1(new_n6826_), .B0(new_n5221_), .Y(new_n11500_));
  OAI22X1  g09064(.A0(new_n11465_), .A1(new_n10486_), .B0(new_n10748_), .B1(new_n3715_), .Y(new_n11501_));
  OR3X1    g09065(.A(new_n10757_), .B(pi0171), .C(pi0051), .Y(new_n11502_));
  NAND2X1  g09066(.A(pi0216), .B(pi0164), .Y(new_n11503_));
  AOI21X1  g09067(.A0(new_n11226_), .A1(pi0171), .B0(new_n11503_), .Y(new_n11504_));
  AOI22X1  g09068(.A0(new_n11504_), .A1(new_n11502_), .B0(new_n11501_), .B1(new_n2438_), .Y(new_n11505_));
  OAI22X1  g09069(.A0(new_n11505_), .A1(new_n5221_), .B0(new_n11500_), .B1(new_n11499_), .Y(new_n11506_));
  AOI22X1  g09070(.A0(new_n11462_), .A1(new_n11244_), .B0(pi0186), .B1(pi0039), .Y(new_n11507_));
  OAI21X1  g09071(.A0(new_n11459_), .A1(new_n11231_), .B0(new_n11507_), .Y(new_n11508_));
  INVX1    g09072(.A(new_n11242_), .Y(new_n11509_));
  AOI21X1  g09073(.A0(new_n11462_), .A1(new_n11509_), .B0(new_n6818_), .Y(new_n11510_));
  OAI21X1  g09074(.A0(new_n11459_), .A1(new_n11229_), .B0(new_n11510_), .Y(new_n11511_));
  AOI22X1  g09075(.A0(new_n11511_), .A1(new_n11508_), .B0(new_n11506_), .B1(pi0299), .Y(new_n11512_));
  OAI21X1  g09076(.A0(new_n11512_), .A1(new_n5215_), .B0(new_n11498_), .Y(new_n11513_));
  INVX1    g09077(.A(new_n11479_), .Y(new_n11514_));
  NAND3X1  g09078(.A(new_n11514_), .B(new_n11254_), .C(pi0232), .Y(new_n11515_));
  AOI22X1  g09079(.A0(new_n11514_), .A1(pi0232), .B0(new_n10416_), .B1(new_n10412_), .Y(new_n11516_));
  NOR2X1   g09080(.A(new_n11516_), .B(pi0039), .Y(new_n11517_));
  AOI21X1  g09081(.A0(new_n11517_), .A1(new_n11515_), .B0(new_n3252_), .Y(new_n11518_));
  AOI21X1  g09082(.A0(new_n11518_), .A1(new_n11513_), .B0(new_n11497_), .Y(new_n11519_));
  AND2X1   g09083(.A(new_n11480_), .B(new_n11102_), .Y(new_n11520_));
  OAI21X1  g09084(.A0(new_n11520_), .A1(new_n10613_), .B0(new_n11452_), .Y(new_n11521_));
  OAI21X1  g09085(.A0(new_n11521_), .A1(new_n11519_), .B0(new_n6489_), .Y(new_n11522_));
  OAI21X1  g09086(.A0(new_n11522_), .A1(new_n11496_), .B0(new_n11456_), .Y(po0291));
  AND2X1   g09087(.A(pi0299), .B(pi0232), .Y(new_n11524_));
  AND3X1   g09088(.A(new_n11524_), .B(new_n5023_), .C(pi0170), .Y(new_n11525_));
  NOR3X1   g09089(.A(new_n11525_), .B(new_n10340_), .C(pi0051), .Y(new_n11526_));
  INVX1    g09090(.A(new_n11526_), .Y(new_n11527_));
  AOI21X1  g09091(.A0(new_n6827_), .A1(pi0194), .B0(new_n11527_), .Y(new_n11528_));
  NOR2X1   g09092(.A(new_n11528_), .B(new_n10998_), .Y(new_n11529_));
  AOI21X1  g09093(.A0(new_n11529_), .A1(pi0100), .B0(new_n10539_), .Y(new_n11530_));
  AND2X1   g09094(.A(new_n5023_), .B(pi0170), .Y(new_n11531_));
  AOI21X1  g09095(.A0(new_n10747_), .A1(pi0170), .B0(new_n6271_), .Y(new_n11532_));
  OAI21X1  g09096(.A0(new_n11531_), .A1(new_n10486_), .B0(new_n11532_), .Y(new_n11533_));
  NAND2X1  g09097(.A(new_n11533_), .B(new_n7187_), .Y(new_n11534_));
  NOR3X1   g09098(.A(new_n10757_), .B(pi0170), .C(pi0051), .Y(new_n11535_));
  NOR3X1   g09099(.A(new_n10785_), .B(new_n10886_), .C(new_n3865_), .Y(new_n11536_));
  OR2X1    g09100(.A(new_n11536_), .B(new_n2438_), .Y(new_n11537_));
  OAI21X1  g09101(.A0(new_n11537_), .A1(new_n11535_), .B0(new_n11534_), .Y(new_n11538_));
  NAND2X1  g09102(.A(pi0299), .B(pi0150), .Y(new_n11539_));
  AOI21X1  g09103(.A0(new_n11531_), .A1(new_n10455_), .B0(pi0051), .Y(new_n11540_));
  AOI21X1  g09104(.A0(new_n11540_), .A1(new_n5221_), .B0(new_n11539_), .Y(new_n11541_));
  AND2X1   g09105(.A(pi0299), .B(new_n9837_), .Y(new_n11542_));
  INVX1    g09106(.A(new_n11542_), .Y(new_n11543_));
  AOI21X1  g09107(.A0(new_n11540_), .A1(new_n6271_), .B0(new_n11543_), .Y(new_n11544_));
  AOI22X1  g09108(.A0(new_n11544_), .A1(new_n11533_), .B0(new_n11541_), .B1(new_n11538_), .Y(new_n11545_));
  AOI21X1  g09109(.A0(new_n11243_), .A1(new_n9902_), .B0(pi0299), .Y(new_n11546_));
  OAI21X1  g09110(.A0(new_n11509_), .A1(new_n9902_), .B0(new_n11546_), .Y(new_n11547_));
  AOI21X1  g09111(.A0(new_n11547_), .A1(new_n11545_), .B0(new_n5215_), .Y(new_n11548_));
  AOI21X1  g09112(.A0(new_n10416_), .A1(new_n10412_), .B0(pi0299), .Y(new_n11549_));
  NOR2X1   g09113(.A(new_n11254_), .B(new_n3865_), .Y(new_n11550_));
  OAI21X1  g09114(.A0(new_n11252_), .A1(pi0170), .B0(new_n11524_), .Y(new_n11551_));
  OAI21X1  g09115(.A0(new_n11551_), .A1(new_n11550_), .B0(new_n11253_), .Y(new_n11552_));
  OAI22X1  g09116(.A0(new_n11552_), .A1(new_n11549_), .B0(new_n11548_), .B1(new_n11250_), .Y(new_n11553_));
  INVX1    g09117(.A(pi0194), .Y(new_n11554_));
  OAI21X1  g09118(.A0(new_n11526_), .A1(new_n10998_), .B0(pi0038), .Y(new_n11555_));
  NAND2X1  g09119(.A(new_n11555_), .B(new_n11554_), .Y(new_n11556_));
  AOI21X1  g09120(.A0(new_n11553_), .A1(new_n2979_), .B0(new_n11556_), .Y(new_n11557_));
  AND2X1   g09121(.A(new_n11229_), .B(pi0185), .Y(new_n11558_));
  OAI21X1  g09122(.A0(new_n11232_), .A1(pi0185), .B0(new_n2933_), .Y(new_n11559_));
  OAI21X1  g09123(.A0(new_n11559_), .A1(new_n11558_), .B0(new_n11545_), .Y(new_n11560_));
  AND2X1   g09124(.A(new_n11560_), .B(pi0232), .Y(new_n11561_));
  AND2X1   g09125(.A(new_n11254_), .B(new_n7876_), .Y(new_n11562_));
  OAI22X1  g09126(.A0(new_n11562_), .A1(new_n11552_), .B0(new_n11561_), .B1(new_n11250_), .Y(new_n11563_));
  AND3X1   g09127(.A(new_n5023_), .B(pi0232), .C(pi0170), .Y(new_n11564_));
  NOR4X1   g09128(.A(new_n11564_), .B(new_n10340_), .C(new_n6827_), .D(pi0051), .Y(new_n11565_));
  OAI21X1  g09129(.A0(new_n11565_), .A1(new_n10998_), .B0(pi0038), .Y(new_n11566_));
  NAND2X1  g09130(.A(new_n11566_), .B(pi0194), .Y(new_n11567_));
  AOI21X1  g09131(.A0(new_n11563_), .A1(new_n2979_), .B0(new_n11567_), .Y(new_n11568_));
  OAI21X1  g09132(.A0(new_n11568_), .A1(new_n11557_), .B0(new_n3007_), .Y(new_n11569_));
  AOI21X1  g09133(.A0(new_n11223_), .A1(new_n11450_), .B0(new_n11449_), .Y(new_n11570_));
  AOI21X1  g09134(.A0(new_n11451_), .A1(pi0134), .B0(new_n11570_), .Y(new_n11571_));
  INVX1    g09135(.A(new_n11571_), .Y(new_n11572_));
  OAI21X1  g09136(.A0(new_n11529_), .A1(new_n10613_), .B0(new_n11572_), .Y(new_n11573_));
  AOI21X1  g09137(.A0(new_n11569_), .A1(new_n11530_), .B0(new_n11573_), .Y(new_n11574_));
  OAI21X1  g09138(.A0(new_n11527_), .A1(new_n8169_), .B0(new_n11554_), .Y(new_n11575_));
  INVX1    g09139(.A(new_n8169_), .Y(new_n11576_));
  AOI21X1  g09140(.A0(new_n11565_), .A1(new_n11576_), .B0(new_n11554_), .Y(new_n11577_));
  INVX1    g09141(.A(new_n11577_), .Y(new_n11578_));
  AND2X1   g09142(.A(new_n11578_), .B(new_n11575_), .Y(new_n11579_));
  AOI21X1  g09143(.A0(new_n10898_), .A1(pi0185), .B0(new_n11461_), .Y(new_n11580_));
  NOR3X1   g09144(.A(new_n10903_), .B(pi0185), .C(pi0051), .Y(new_n11581_));
  OR3X1    g09145(.A(new_n11578_), .B(new_n11581_), .C(new_n11460_), .Y(new_n11582_));
  OAI21X1  g09146(.A0(new_n11575_), .A1(new_n11580_), .B0(new_n11582_), .Y(new_n11583_));
  NOR2X1   g09147(.A(new_n11190_), .B(new_n3865_), .Y(new_n11584_));
  OAI21X1  g09148(.A0(new_n10897_), .A1(pi0170), .B0(new_n6856_), .Y(new_n11585_));
  NOR2X1   g09149(.A(new_n11585_), .B(new_n11584_), .Y(new_n11586_));
  AND3X1   g09150(.A(new_n5023_), .B(new_n2986_), .C(pi0170), .Y(new_n11587_));
  OAI21X1  g09151(.A0(new_n11531_), .A1(new_n10501_), .B0(new_n6856_), .Y(new_n11588_));
  OAI21X1  g09152(.A0(new_n11588_), .A1(new_n11587_), .B0(new_n11542_), .Y(new_n11589_));
  OAI21X1  g09153(.A0(new_n11586_), .A1(new_n11539_), .B0(new_n11589_), .Y(new_n11590_));
  NOR4X1   g09154(.A(new_n11531_), .B(new_n10340_), .C(new_n6856_), .D(pi0051), .Y(new_n11591_));
  AOI21X1  g09155(.A0(new_n11578_), .A1(new_n11575_), .B0(new_n11591_), .Y(new_n11592_));
  AOI22X1  g09156(.A0(new_n11592_), .A1(new_n11590_), .B0(new_n11583_), .B1(new_n2933_), .Y(new_n11593_));
  OAI22X1  g09157(.A0(new_n11593_), .A1(new_n5215_), .B0(new_n11579_), .B1(new_n11184_), .Y(new_n11594_));
  OAI21X1  g09158(.A0(new_n10342_), .A1(new_n3007_), .B0(new_n11530_), .Y(new_n11595_));
  AOI21X1  g09159(.A0(new_n11594_), .A1(new_n3007_), .B0(new_n11595_), .Y(new_n11596_));
  AND2X1   g09160(.A(new_n11528_), .B(new_n10544_), .Y(new_n11597_));
  OR2X1    g09161(.A(new_n11597_), .B(new_n11572_), .Y(new_n11598_));
  OAI21X1  g09162(.A0(new_n11598_), .A1(new_n11596_), .B0(new_n6489_), .Y(new_n11599_));
  AOI21X1  g09163(.A0(new_n11564_), .A1(new_n10455_), .B0(new_n11453_), .Y(new_n11600_));
  OAI21X1  g09164(.A0(new_n11572_), .A1(new_n10455_), .B0(new_n11600_), .Y(new_n11601_));
  OAI21X1  g09165(.A0(new_n11599_), .A1(new_n11574_), .B0(new_n11601_), .Y(po0292));
  NOR3X1   g09166(.A(pi0136), .B(pi0135), .C(pi0134), .Y(new_n11603_));
  XOR2X1   g09167(.A(new_n11223_), .B(new_n11450_), .Y(new_n11604_));
  NOR2X1   g09168(.A(new_n11604_), .B(new_n11603_), .Y(new_n11605_));
  NAND3X1  g09169(.A(new_n5023_), .B(pi0232), .C(pi0148), .Y(new_n11606_));
  AOI22X1  g09170(.A0(new_n11606_), .A1(new_n10455_), .B0(new_n11605_), .B1(new_n11209_), .Y(new_n11607_));
  AND2X1   g09171(.A(new_n2933_), .B(pi0141), .Y(new_n11608_));
  INVX1    g09172(.A(new_n11608_), .Y(new_n11609_));
  AND2X1   g09173(.A(pi0299), .B(pi0148), .Y(new_n11610_));
  INVX1    g09174(.A(new_n11610_), .Y(new_n11611_));
  AOI21X1  g09175(.A0(new_n11611_), .A1(new_n11609_), .B0(new_n11254_), .Y(new_n11612_));
  OAI21X1  g09176(.A0(new_n11252_), .A1(new_n7334_), .B0(pi0232), .Y(new_n11613_));
  OAI21X1  g09177(.A0(new_n11613_), .A1(new_n11612_), .B0(new_n11253_), .Y(new_n11614_));
  OAI21X1  g09178(.A0(new_n11232_), .A1(pi0184), .B0(new_n11608_), .Y(new_n11615_));
  AOI21X1  g09179(.A0(new_n11229_), .A1(pi0184), .B0(new_n11615_), .Y(new_n11616_));
  AND2X1   g09180(.A(new_n11242_), .B(pi0184), .Y(new_n11617_));
  NOR2X1   g09181(.A(pi0299), .B(pi0141), .Y(new_n11618_));
  OAI21X1  g09182(.A0(new_n11244_), .A1(pi0184), .B0(new_n11618_), .Y(new_n11619_));
  NOR2X1   g09183(.A(new_n11227_), .B(new_n6271_), .Y(new_n11620_));
  NOR4X1   g09184(.A(new_n10785_), .B(new_n10886_), .C(new_n5221_), .D(new_n8623_), .Y(new_n11621_));
  OAI21X1  g09185(.A0(new_n10998_), .A1(new_n6270_), .B0(new_n8623_), .Y(new_n11622_));
  OAI21X1  g09186(.A0(new_n11102_), .A1(new_n5220_), .B0(new_n11622_), .Y(new_n11623_));
  OAI21X1  g09187(.A0(new_n11623_), .A1(new_n11621_), .B0(pi0148), .Y(new_n11624_));
  AND3X1   g09188(.A(new_n5023_), .B(new_n7795_), .C(pi0163), .Y(new_n11625_));
  OR2X1    g09189(.A(new_n11625_), .B(new_n2438_), .Y(new_n11626_));
  AND2X1   g09190(.A(new_n11626_), .B(new_n5220_), .Y(new_n11627_));
  OR2X1    g09191(.A(pi0148), .B(pi0051), .Y(new_n11628_));
  AOI21X1  g09192(.A0(new_n11627_), .A1(new_n10485_), .B0(new_n11628_), .Y(new_n11629_));
  NOR2X1   g09193(.A(new_n11629_), .B(new_n2933_), .Y(new_n11630_));
  OAI21X1  g09194(.A0(new_n11624_), .A1(new_n11620_), .B0(new_n11630_), .Y(new_n11631_));
  OAI21X1  g09195(.A0(new_n11619_), .A1(new_n11617_), .B0(new_n11631_), .Y(new_n11632_));
  OAI21X1  g09196(.A0(new_n11632_), .A1(new_n11616_), .B0(pi0232), .Y(new_n11633_));
  AOI21X1  g09197(.A0(new_n11633_), .A1(new_n11498_), .B0(new_n3252_), .Y(new_n11634_));
  NAND2X1  g09198(.A(new_n11634_), .B(new_n11614_), .Y(new_n11635_));
  OAI21X1  g09199(.A0(new_n10340_), .A1(new_n7335_), .B0(new_n2534_), .Y(new_n11636_));
  AOI21X1  g09200(.A0(new_n11636_), .A1(new_n3252_), .B0(new_n10539_), .Y(new_n11637_));
  OR2X1    g09201(.A(new_n11636_), .B(new_n10613_), .Y(new_n11638_));
  NAND2X1  g09202(.A(new_n11638_), .B(new_n11605_), .Y(new_n11639_));
  AOI21X1  g09203(.A0(new_n11637_), .A1(new_n11635_), .B0(new_n11639_), .Y(new_n11640_));
  NAND4X1  g09204(.A(new_n10455_), .B(new_n8260_), .C(new_n7335_), .D(new_n2534_), .Y(new_n11641_));
  AND2X1   g09205(.A(new_n10492_), .B(pi0184), .Y(new_n11642_));
  OAI21X1  g09206(.A0(new_n11642_), .A1(new_n11187_), .B0(new_n11608_), .Y(new_n11643_));
  NOR3X1   g09207(.A(new_n10487_), .B(new_n7187_), .C(pi0051), .Y(new_n11644_));
  OAI21X1  g09208(.A0(new_n11199_), .A1(new_n5023_), .B0(pi0148), .Y(new_n11645_));
  AOI21X1  g09209(.A0(new_n10912_), .A1(new_n2534_), .B0(pi0148), .Y(new_n11646_));
  OAI22X1  g09210(.A0(new_n11646_), .A1(new_n11625_), .B0(new_n11209_), .B1(pi0148), .Y(new_n11647_));
  OAI21X1  g09211(.A0(new_n11645_), .A1(new_n11644_), .B0(new_n11647_), .Y(new_n11648_));
  OAI21X1  g09212(.A0(new_n11203_), .A1(new_n8634_), .B0(new_n11204_), .Y(new_n11649_));
  AOI22X1  g09213(.A0(new_n11649_), .A1(new_n11618_), .B0(new_n11648_), .B1(pi0299), .Y(new_n11650_));
  AOI21X1  g09214(.A0(new_n11650_), .A1(new_n11643_), .B0(new_n5215_), .Y(new_n11651_));
  NAND3X1  g09215(.A(new_n11183_), .B(new_n8169_), .C(new_n3007_), .Y(new_n11652_));
  OAI21X1  g09216(.A0(new_n11652_), .A1(new_n11651_), .B0(new_n11641_), .Y(new_n11653_));
  OAI22X1  g09217(.A0(new_n11638_), .A1(new_n10340_), .B0(new_n11604_), .B1(new_n11603_), .Y(new_n11654_));
  AOI21X1  g09218(.A0(new_n11653_), .A1(new_n5813_), .B0(new_n11654_), .Y(new_n11655_));
  OR2X1    g09219(.A(new_n11655_), .B(po1038), .Y(new_n11656_));
  OAI22X1  g09220(.A0(new_n11656_), .A1(new_n11640_), .B0(new_n11607_), .B1(new_n11453_), .Y(po0293));
  OR4X1    g09221(.A(new_n10655_), .B(new_n2985_), .C(new_n2536_), .D(new_n7795_), .Y(new_n11658_));
  AND3X1   g09222(.A(new_n8556_), .B(pi0299), .C(new_n2777_), .Y(new_n11659_));
  AND3X1   g09223(.A(new_n5102_), .B(new_n2933_), .C(new_n2436_), .Y(new_n11660_));
  AND3X1   g09224(.A(new_n11660_), .B(new_n8561_), .C(new_n2954_), .Y(new_n11661_));
  OR2X1    g09225(.A(new_n11661_), .B(new_n11659_), .Y(new_n11662_));
  AND3X1   g09226(.A(new_n7717_), .B(new_n4510_), .C(new_n2777_), .Y(new_n11663_));
  AOI22X1  g09227(.A0(new_n11663_), .A1(po1038), .B0(new_n11662_), .B1(new_n11658_), .Y(new_n11664_));
  OAI22X1  g09228(.A0(new_n11664_), .A1(new_n9566_), .B0(new_n2452_), .B1(pi0039), .Y(po0294));
  INVX1    g09229(.A(pi0138), .Y(new_n11666_));
  AND3X1   g09230(.A(new_n6843_), .B(new_n3131_), .C(new_n2939_), .Y(new_n11667_));
  NOR2X1   g09231(.A(new_n7461_), .B(new_n11667_), .Y(new_n11668_));
  OAI21X1  g09232(.A0(new_n11668_), .A1(new_n3079_), .B0(new_n3102_), .Y(new_n11669_));
  NOR2X1   g09233(.A(new_n7134_), .B(pi0075), .Y(new_n11670_));
  AOI21X1  g09234(.A0(new_n7089_), .A1(new_n7063_), .B0(new_n2933_), .Y(new_n11671_));
  AOI21X1  g09235(.A0(new_n7089_), .A1(new_n6948_), .B0(pi0299), .Y(new_n11672_));
  NOR3X1   g09236(.A(new_n11672_), .B(new_n11671_), .C(pi0232), .Y(new_n11673_));
  NOR2X1   g09237(.A(new_n11673_), .B(pi0039), .Y(new_n11674_));
  INVX1    g09238(.A(new_n11674_), .Y(new_n11675_));
  INVX1    g09239(.A(pi0141), .Y(new_n11676_));
  AND2X1   g09240(.A(new_n7089_), .B(new_n6948_), .Y(new_n11677_));
  MX2X1    g09241(.A(new_n11677_), .B(new_n6967_), .S0(new_n5023_), .Y(new_n11678_));
  OR3X1    g09242(.A(new_n11678_), .B(pi0299), .C(new_n11676_), .Y(new_n11679_));
  AND2X1   g09243(.A(new_n7089_), .B(new_n7063_), .Y(new_n11680_));
  NOR2X1   g09244(.A(new_n7066_), .B(new_n5048_), .Y(new_n11681_));
  INVX1    g09245(.A(new_n11681_), .Y(new_n11682_));
  AND2X1   g09246(.A(new_n5023_), .B(pi0148), .Y(new_n11683_));
  OAI22X1  g09247(.A0(new_n11683_), .A1(new_n11680_), .B0(new_n11682_), .B1(new_n4046_), .Y(new_n11684_));
  OR2X1    g09248(.A(new_n11677_), .B(pi0299), .Y(new_n11685_));
  OAI21X1  g09249(.A0(new_n11685_), .A1(pi0141), .B0(pi0232), .Y(new_n11686_));
  AOI21X1  g09250(.A0(new_n11684_), .A1(pi0299), .B0(new_n11686_), .Y(new_n11687_));
  AOI21X1  g09251(.A0(new_n11687_), .A1(new_n11679_), .B0(new_n11675_), .Y(new_n11688_));
  OR2X1    g09252(.A(new_n6861_), .B(new_n6835_), .Y(new_n11689_));
  AOI21X1  g09253(.A0(new_n8829_), .A1(new_n11689_), .B0(new_n6874_), .Y(new_n11690_));
  NOR2X1   g09254(.A(new_n11690_), .B(new_n9927_), .Y(new_n11691_));
  AND2X1   g09255(.A(new_n8829_), .B(new_n11689_), .Y(new_n11692_));
  AND2X1   g09256(.A(new_n11689_), .B(new_n5059_), .Y(new_n11693_));
  NOR3X1   g09257(.A(new_n11693_), .B(new_n11692_), .C(new_n7187_), .Y(new_n11694_));
  NOR2X1   g09258(.A(new_n11694_), .B(new_n8800_), .Y(new_n11695_));
  OAI21X1  g09259(.A0(new_n11695_), .A1(new_n11691_), .B0(new_n5215_), .Y(new_n11696_));
  NOR2X1   g09260(.A(new_n6859_), .B(new_n5058_), .Y(new_n11697_));
  OAI21X1  g09261(.A0(new_n11692_), .A1(new_n11697_), .B0(new_n6857_), .Y(new_n11698_));
  NOR2X1   g09262(.A(new_n11695_), .B(new_n11610_), .Y(new_n11699_));
  AOI21X1  g09263(.A0(new_n11698_), .A1(pi0148), .B0(new_n11699_), .Y(new_n11700_));
  AOI21X1  g09264(.A0(new_n11690_), .A1(new_n6879_), .B0(new_n9927_), .Y(new_n11701_));
  MX2X1    g09265(.A(new_n11701_), .B(new_n11691_), .S0(new_n11676_), .Y(new_n11702_));
  OAI21X1  g09266(.A0(new_n11702_), .A1(new_n11700_), .B0(pi0232), .Y(new_n11703_));
  AOI21X1  g09267(.A0(new_n11703_), .A1(new_n11696_), .B0(new_n2939_), .Y(new_n11704_));
  OR2X1    g09268(.A(new_n11704_), .B(new_n3252_), .Y(new_n11705_));
  OAI21X1  g09269(.A0(new_n11705_), .A1(new_n11688_), .B0(new_n3131_), .Y(new_n11706_));
  AOI21X1  g09270(.A0(new_n11706_), .A1(new_n11670_), .B0(pi0092), .Y(new_n11707_));
  OAI21X1  g09271(.A0(new_n11707_), .A1(new_n11669_), .B0(new_n3107_), .Y(new_n11708_));
  AND2X1   g09272(.A(new_n11667_), .B(new_n3079_), .Y(new_n11709_));
  OAI21X1  g09273(.A0(new_n11709_), .A1(new_n7322_), .B0(pi0055), .Y(new_n11710_));
  AOI21X1  g09274(.A0(new_n11710_), .A1(new_n11708_), .B0(new_n4975_), .Y(new_n11711_));
  OR3X1    g09275(.A(new_n11711_), .B(new_n9836_), .C(new_n11666_), .Y(new_n11712_));
  AND2X1   g09276(.A(new_n8492_), .B(new_n5215_), .Y(new_n11713_));
  INVX1    g09277(.A(new_n11713_), .Y(new_n11714_));
  NOR4X1   g09278(.A(new_n5239_), .B(new_n5228_), .C(new_n5224_), .D(new_n6256_), .Y(new_n11715_));
  AND2X1   g09279(.A(new_n11715_), .B(new_n6848_), .Y(new_n11716_));
  OAI22X1  g09280(.A0(new_n11716_), .A1(new_n11609_), .B0(new_n11611_), .B1(new_n6255_), .Y(new_n11717_));
  AOI21X1  g09281(.A0(new_n8492_), .A1(new_n11609_), .B0(new_n11717_), .Y(new_n11718_));
  OR2X1    g09282(.A(new_n11718_), .B(new_n5215_), .Y(new_n11719_));
  AOI21X1  g09283(.A0(new_n11719_), .A1(new_n11714_), .B0(new_n2939_), .Y(new_n11720_));
  AOI21X1  g09284(.A0(new_n9998_), .A1(new_n7335_), .B0(pi0039), .Y(new_n11721_));
  NOR3X1   g09285(.A(new_n11721_), .B(new_n11720_), .C(new_n7629_), .Y(new_n11722_));
  INVX1    g09286(.A(pi0139), .Y(new_n11723_));
  AND3X1   g09287(.A(new_n9963_), .B(new_n11723_), .C(new_n6785_), .Y(new_n11724_));
  AOI21X1  g09288(.A0(new_n11722_), .A1(new_n11666_), .B0(new_n11724_), .Y(new_n11725_));
  OAI21X1  g09289(.A0(pi0196), .A1(pi0195), .B0(new_n11666_), .Y(new_n11726_));
  OR3X1    g09290(.A(new_n11726_), .B(new_n11711_), .C(new_n9836_), .Y(new_n11727_));
  INVX1    g09291(.A(new_n11724_), .Y(new_n11728_));
  AOI21X1  g09292(.A0(new_n11726_), .A1(new_n11722_), .B0(new_n11728_), .Y(new_n11729_));
  AOI22X1  g09293(.A0(new_n11729_), .A1(new_n11727_), .B0(new_n11725_), .B1(new_n11712_), .Y(po0295));
  OR3X1    g09294(.A(new_n11678_), .B(pi0299), .C(new_n6810_), .Y(new_n11731_));
  OAI22X1  g09295(.A0(new_n11194_), .A1(new_n11680_), .B0(new_n11682_), .B1(new_n4162_), .Y(new_n11732_));
  OAI21X1  g09296(.A0(new_n11685_), .A1(pi0191), .B0(pi0232), .Y(new_n11733_));
  AOI21X1  g09297(.A0(new_n11732_), .A1(pi0299), .B0(new_n11733_), .Y(new_n11734_));
  AOI21X1  g09298(.A0(new_n11734_), .A1(new_n11731_), .B0(new_n11675_), .Y(new_n11735_));
  OAI22X1  g09299(.A0(new_n11692_), .A1(new_n11697_), .B0(new_n11689_), .B1(pi0169), .Y(new_n11736_));
  AOI21X1  g09300(.A0(new_n11736_), .A1(new_n6856_), .B0(new_n8800_), .Y(new_n11737_));
  MX2X1    g09301(.A(new_n11701_), .B(new_n11691_), .S0(new_n6810_), .Y(new_n11738_));
  OAI21X1  g09302(.A0(new_n11738_), .A1(new_n11737_), .B0(pi0232), .Y(new_n11739_));
  AOI21X1  g09303(.A0(new_n11739_), .A1(new_n11696_), .B0(new_n2939_), .Y(new_n11740_));
  OR2X1    g09304(.A(new_n11740_), .B(new_n3252_), .Y(new_n11741_));
  OAI21X1  g09305(.A0(new_n11741_), .A1(new_n11735_), .B0(new_n3131_), .Y(new_n11742_));
  AOI21X1  g09306(.A0(new_n11742_), .A1(new_n11670_), .B0(pi0092), .Y(new_n11743_));
  OAI21X1  g09307(.A0(new_n11743_), .A1(new_n11669_), .B0(new_n3107_), .Y(new_n11744_));
  AOI21X1  g09308(.A0(new_n11744_), .A1(new_n11710_), .B0(new_n4975_), .Y(new_n11745_));
  OR3X1    g09309(.A(new_n11745_), .B(new_n9836_), .C(new_n11723_), .Y(new_n11746_));
  NOR3X1   g09310(.A(new_n6255_), .B(new_n2933_), .C(new_n4162_), .Y(new_n11747_));
  NOR3X1   g09311(.A(new_n8489_), .B(pi0299), .C(pi0191), .Y(new_n11748_));
  NOR3X1   g09312(.A(new_n11716_), .B(pi0299), .C(new_n6810_), .Y(new_n11749_));
  OR4X1    g09313(.A(new_n11749_), .B(new_n11748_), .C(new_n11747_), .D(new_n8490_), .Y(new_n11750_));
  MX2X1    g09314(.A(new_n11750_), .B(new_n8492_), .S0(new_n5215_), .Y(new_n11751_));
  NOR3X1   g09315(.A(new_n11210_), .B(new_n7251_), .C(new_n7619_), .Y(new_n11752_));
  OAI21X1  g09316(.A0(new_n11752_), .A1(pi0039), .B0(new_n7628_), .Y(new_n11753_));
  AOI21X1  g09317(.A0(new_n11751_), .A1(pi0039), .B0(new_n11753_), .Y(new_n11754_));
  AOI22X1  g09318(.A0(new_n11754_), .A1(new_n11723_), .B0(new_n9963_), .B1(new_n6785_), .Y(new_n11755_));
  NOR3X1   g09319(.A(pi0196), .B(pi0195), .C(pi0138), .Y(new_n11756_));
  OR2X1    g09320(.A(new_n11756_), .B(pi0139), .Y(new_n11757_));
  OR3X1    g09321(.A(new_n11757_), .B(new_n11745_), .C(new_n9836_), .Y(new_n11758_));
  NAND2X1  g09322(.A(new_n9963_), .B(new_n6785_), .Y(new_n11759_));
  AOI21X1  g09323(.A0(new_n11757_), .A1(new_n11754_), .B0(new_n11759_), .Y(new_n11760_));
  AOI22X1  g09324(.A0(new_n11760_), .A1(new_n11758_), .B0(new_n11755_), .B1(new_n11746_), .Y(po0296));
  INVX1    g09325(.A(pi1160), .Y(new_n11762_));
  INVX1    g09326(.A(pi0787), .Y(new_n11763_));
  INVX1    g09327(.A(pi0792), .Y(new_n11764_));
  INVX1    g09328(.A(pi0788), .Y(new_n11765_));
  INVX1    g09329(.A(pi0789), .Y(new_n11766_));
  INVX1    g09330(.A(pi0781), .Y(new_n11767_));
  INVX1    g09331(.A(pi0785), .Y(new_n11768_));
  INVX1    g09332(.A(pi0778), .Y(new_n11769_));
  INVX1    g09333(.A(new_n3103_), .Y(new_n11770_));
  INVX1    g09334(.A(pi0738), .Y(new_n11771_));
  INVX1    g09335(.A(pi0761), .Y(new_n11772_));
  AND2X1   g09336(.A(new_n8370_), .B(new_n2580_), .Y(new_n11773_));
  OR4X1    g09337(.A(new_n2472_), .B(pi0088), .C(pi0077), .D(pi0050), .Y(new_n11774_));
  NOR4X1   g09338(.A(new_n11774_), .B(new_n11773_), .C(new_n2582_), .D(pi0098), .Y(new_n11775_));
  AND2X1   g09339(.A(new_n6933_), .B(new_n6737_), .Y(new_n11776_));
  AOI21X1  g09340(.A0(new_n11776_), .A1(new_n11775_), .B0(pi0040), .Y(new_n11777_));
  OAI21X1  g09341(.A0(new_n11777_), .A1(new_n7683_), .B0(new_n3035_), .Y(new_n11778_));
  NOR3X1   g09342(.A(new_n2553_), .B(new_n2728_), .C(pi0091), .Y(new_n11779_));
  NOR3X1   g09343(.A(new_n2495_), .B(new_n2473_), .C(pi0094), .Y(new_n11780_));
  AND2X1   g09344(.A(new_n11775_), .B(new_n11780_), .Y(new_n11781_));
  OR2X1    g09345(.A(new_n11781_), .B(pi0047), .Y(new_n11782_));
  NOR3X1   g09346(.A(new_n7665_), .B(new_n2562_), .C(new_n5117_), .Y(new_n11783_));
  OAI21X1  g09347(.A0(new_n11783_), .A1(new_n11782_), .B0(new_n11779_), .Y(new_n11784_));
  NAND2X1  g09348(.A(new_n7677_), .B(new_n2529_), .Y(new_n11785_));
  AOI21X1  g09349(.A0(new_n11784_), .A1(new_n2508_), .B0(new_n11785_), .Y(new_n11786_));
  NAND2X1  g09350(.A(new_n7584_), .B(pi0252), .Y(new_n11787_));
  OAI21X1  g09351(.A0(new_n11787_), .A1(new_n11786_), .B0(new_n11778_), .Y(new_n11788_));
  NOR4X1   g09352(.A(new_n11788_), .B(new_n8959_), .C(new_n7250_), .D(new_n5024_), .Y(new_n11789_));
  INVX1    g09353(.A(new_n7683_), .Y(new_n11790_));
  OR3X1    g09354(.A(new_n11773_), .B(new_n2582_), .C(pi0098), .Y(new_n11791_));
  AOI21X1  g09355(.A0(new_n11791_), .A1(new_n2663_), .B0(new_n8183_), .Y(new_n11792_));
  AND2X1   g09356(.A(new_n11792_), .B(new_n2552_), .Y(new_n11793_));
  OR2X1    g09357(.A(new_n11783_), .B(pi0047), .Y(new_n11794_));
  OAI21X1  g09358(.A0(new_n11794_), .A1(new_n11793_), .B0(new_n11779_), .Y(new_n11795_));
  AND2X1   g09359(.A(new_n11795_), .B(new_n2508_), .Y(new_n11796_));
  NAND2X1  g09360(.A(new_n7677_), .B(pi0252), .Y(new_n11797_));
  NOR4X1   g09361(.A(new_n8172_), .B(new_n6954_), .C(new_n2484_), .D(pi0252), .Y(new_n11798_));
  AOI21X1  g09362(.A0(new_n11798_), .A1(new_n11792_), .B0(pi0040), .Y(new_n11799_));
  OAI21X1  g09363(.A0(new_n11797_), .A1(new_n11796_), .B0(new_n11799_), .Y(new_n11800_));
  AND3X1   g09364(.A(new_n11800_), .B(new_n11790_), .C(new_n5927_), .Y(new_n11801_));
  OAI21X1  g09365(.A0(new_n11801_), .A1(new_n11789_), .B0(pi1093), .Y(new_n11802_));
  NOR2X1   g09366(.A(new_n11788_), .B(new_n7250_), .Y(new_n11803_));
  AND3X1   g09367(.A(new_n2759_), .B(new_n5922_), .C(pi1092), .Y(po1106));
  AOI21X1  g09368(.A0(po1106), .A1(new_n11803_), .B0(new_n2703_), .Y(new_n11805_));
  AOI21X1  g09369(.A0(new_n11802_), .A1(new_n8194_), .B0(new_n11805_), .Y(new_n11806_));
  NOR2X1   g09370(.A(new_n11802_), .B(pi1091), .Y(new_n11807_));
  OR2X1    g09371(.A(new_n11807_), .B(new_n11806_), .Y(new_n11808_));
  AOI21X1  g09372(.A0(new_n11800_), .A1(new_n3175_), .B0(pi0032), .Y(new_n11809_));
  AND2X1   g09373(.A(new_n5225_), .B(new_n2523_), .Y(new_n11810_));
  OAI21X1  g09374(.A0(new_n8383_), .A1(new_n2455_), .B0(new_n11810_), .Y(new_n11811_));
  NOR3X1   g09375(.A(new_n11811_), .B(new_n11809_), .C(new_n8199_), .Y(new_n11812_));
  OAI21X1  g09376(.A0(new_n11812_), .A1(new_n11789_), .B0(new_n5967_), .Y(new_n11813_));
  AOI21X1  g09377(.A0(new_n11788_), .A1(new_n2455_), .B0(new_n11811_), .Y(new_n11814_));
  AND3X1   g09378(.A(new_n11814_), .B(pi0829), .C(new_n8199_), .Y(new_n11815_));
  OR3X1    g09379(.A(new_n11815_), .B(new_n11812_), .C(new_n11789_), .Y(new_n11816_));
  AOI21X1  g09380(.A0(new_n11816_), .A1(pi1093), .B0(new_n5922_), .Y(new_n11817_));
  OAI21X1  g09381(.A0(new_n11817_), .A1(new_n11805_), .B0(new_n11813_), .Y(new_n11818_));
  MX2X1    g09382(.A(new_n11818_), .B(new_n11808_), .S0(new_n2777_), .Y(new_n11819_));
  MX2X1    g09383(.A(new_n11818_), .B(new_n11808_), .S0(new_n2954_), .Y(new_n11820_));
  MX2X1    g09384(.A(new_n11820_), .B(new_n11819_), .S0(pi0299), .Y(new_n11821_));
  INVX1    g09385(.A(new_n11821_), .Y(new_n11822_));
  OR4X1    g09386(.A(new_n7633_), .B(new_n2985_), .C(new_n2536_), .D(pi0287), .Y(new_n11823_));
  MX2X1    g09387(.A(new_n11823_), .B(new_n2986_), .S0(pi0120), .Y(new_n11824_));
  OR2X1    g09388(.A(new_n11824_), .B(new_n2725_), .Y(new_n11825_));
  NOR4X1   g09389(.A(new_n7633_), .B(new_n2985_), .C(new_n2536_), .D(pi0287), .Y(new_n11826_));
  AOI21X1  g09390(.A0(new_n11826_), .A1(new_n2720_), .B0(pi0120), .Y(new_n11827_));
  NOR3X1   g09391(.A(new_n2985_), .B(new_n2725_), .C(new_n2536_), .Y(new_n11828_));
  OR2X1    g09392(.A(new_n10246_), .B(new_n5030_), .Y(new_n11829_));
  AOI21X1  g09393(.A0(new_n11829_), .A1(new_n11828_), .B0(new_n10082_), .Y(new_n11830_));
  NOR3X1   g09394(.A(new_n11830_), .B(new_n11827_), .C(new_n2702_), .Y(new_n11831_));
  OAI21X1  g09395(.A0(new_n11828_), .A1(new_n10082_), .B0(new_n2702_), .Y(new_n11832_));
  NOR3X1   g09396(.A(new_n5030_), .B(new_n8199_), .C(new_n10082_), .Y(new_n11833_));
  NOR3X1   g09397(.A(new_n11833_), .B(new_n11832_), .C(new_n11827_), .Y(new_n11834_));
  NOR2X1   g09398(.A(new_n11834_), .B(new_n11831_), .Y(new_n11835_));
  MX2X1    g09399(.A(new_n11835_), .B(new_n11825_), .S0(new_n5048_), .Y(new_n11836_));
  INVX1    g09400(.A(new_n11836_), .Y(new_n11837_));
  INVX1    g09401(.A(pi0614), .Y(new_n11838_));
  AND2X1   g09402(.A(new_n5016_), .B(pi0603), .Y(new_n11839_));
  INVX1    g09403(.A(new_n11839_), .Y(new_n11840_));
  AND2X1   g09404(.A(new_n11825_), .B(new_n11840_), .Y(new_n11841_));
  OR3X1    g09405(.A(new_n11834_), .B(new_n11831_), .C(new_n5023_), .Y(new_n11842_));
  OAI21X1  g09406(.A0(new_n11824_), .A1(new_n2725_), .B0(new_n5023_), .Y(new_n11843_));
  AOI21X1  g09407(.A0(new_n11843_), .A1(new_n11842_), .B0(new_n11840_), .Y(new_n11844_));
  OAI21X1  g09408(.A0(new_n11844_), .A1(new_n11841_), .B0(new_n11838_), .Y(new_n11845_));
  OAI21X1  g09409(.A0(new_n11845_), .A1(pi0616), .B0(new_n11837_), .Y(new_n11846_));
  AND2X1   g09410(.A(new_n11846_), .B(pi0681), .Y(new_n11847_));
  INVX1    g09411(.A(pi0661), .Y(new_n11848_));
  INVX1    g09412(.A(pi0662), .Y(new_n11849_));
  AND2X1   g09413(.A(pi0680), .B(new_n11849_), .Y(new_n11850_));
  INVX1    g09414(.A(new_n11850_), .Y(new_n11851_));
  OAI21X1  g09415(.A0(new_n11824_), .A1(new_n2725_), .B0(pi0614), .Y(new_n11852_));
  NAND2X1  g09416(.A(new_n11852_), .B(new_n11845_), .Y(new_n11853_));
  MX2X1    g09417(.A(new_n11853_), .B(new_n11825_), .S0(pi0616), .Y(new_n11854_));
  AND2X1   g09418(.A(new_n11854_), .B(new_n11851_), .Y(new_n11855_));
  NOR3X1   g09419(.A(new_n11834_), .B(new_n11831_), .C(new_n11851_), .Y(new_n11856_));
  OR2X1    g09420(.A(new_n11856_), .B(new_n5023_), .Y(new_n11857_));
  OAI22X1  g09421(.A0(new_n11857_), .A1(new_n11855_), .B0(new_n11835_), .B1(new_n5048_), .Y(new_n11858_));
  INVX1    g09422(.A(pi0681), .Y(new_n11859_));
  OAI21X1  g09423(.A0(new_n11846_), .A1(new_n11848_), .B0(new_n11859_), .Y(new_n11860_));
  AOI21X1  g09424(.A0(new_n11858_), .A1(new_n11848_), .B0(new_n11860_), .Y(new_n11861_));
  NOR2X1   g09425(.A(new_n11861_), .B(new_n11847_), .Y(new_n11862_));
  NOR3X1   g09426(.A(pi0681), .B(pi0662), .C(pi0661), .Y(new_n11863_));
  OR2X1    g09427(.A(new_n11863_), .B(pi0616), .Y(new_n11864_));
  NOR2X1   g09428(.A(new_n11864_), .B(new_n11853_), .Y(new_n11865_));
  AOI21X1  g09429(.A0(new_n11852_), .A1(new_n11845_), .B0(pi0616), .Y(new_n11866_));
  INVX1    g09430(.A(new_n11863_), .Y(new_n11867_));
  AOI21X1  g09431(.A0(new_n11843_), .A1(new_n11842_), .B0(new_n5019_), .Y(new_n11868_));
  OR3X1    g09432(.A(new_n11868_), .B(new_n11867_), .C(pi0616), .Y(new_n11869_));
  AOI21X1  g09433(.A0(new_n11866_), .A1(new_n5019_), .B0(new_n11869_), .Y(new_n11870_));
  INVX1    g09434(.A(pi0616), .Y(new_n11871_));
  AND2X1   g09435(.A(new_n11825_), .B(new_n5019_), .Y(new_n11872_));
  OR3X1    g09436(.A(new_n11872_), .B(new_n11867_), .C(new_n11871_), .Y(new_n11873_));
  OR3X1    g09437(.A(new_n11824_), .B(new_n2725_), .C(new_n11871_), .Y(new_n11874_));
  OAI22X1  g09438(.A0(new_n11874_), .A1(new_n11863_), .B0(new_n11873_), .B1(new_n11868_), .Y(new_n11875_));
  NOR4X1   g09439(.A(new_n11875_), .B(new_n11870_), .C(new_n11865_), .D(pi0681), .Y(new_n11876_));
  AOI21X1  g09440(.A0(new_n11854_), .A1(pi0681), .B0(new_n11876_), .Y(new_n11877_));
  MX2X1    g09441(.A(new_n11877_), .B(new_n11862_), .S0(new_n5042_), .Y(new_n11878_));
  NOR2X1   g09442(.A(new_n11878_), .B(new_n2940_), .Y(new_n11879_));
  INVX1    g09443(.A(new_n11825_), .Y(new_n11880_));
  INVX1    g09444(.A(pi0603), .Y(new_n11881_));
  NOR2X1   g09445(.A(new_n11828_), .B(new_n10082_), .Y(new_n11882_));
  AND2X1   g09446(.A(new_n11823_), .B(new_n8199_), .Y(new_n11883_));
  NOR4X1   g09447(.A(new_n7631_), .B(new_n2985_), .C(new_n2536_), .D(pi0287), .Y(new_n11884_));
  AOI21X1  g09448(.A0(new_n11884_), .A1(pi1092), .B0(new_n8200_), .Y(new_n11885_));
  OR3X1    g09449(.A(new_n11885_), .B(new_n11883_), .C(new_n5032_), .Y(new_n11886_));
  AND2X1   g09450(.A(new_n11886_), .B(new_n10082_), .Y(new_n11887_));
  OR2X1    g09451(.A(new_n11887_), .B(new_n11832_), .Y(new_n11888_));
  OR3X1    g09452(.A(new_n11823_), .B(new_n2725_), .C(new_n8194_), .Y(new_n11889_));
  OR2X1    g09453(.A(new_n11826_), .B(pi0824), .Y(new_n11890_));
  INVX1    g09454(.A(new_n8200_), .Y(new_n11891_));
  OR4X1    g09455(.A(new_n7631_), .B(new_n2985_), .C(new_n2536_), .D(pi0287), .Y(new_n11892_));
  OAI21X1  g09456(.A0(new_n11892_), .A1(new_n5024_), .B0(new_n11891_), .Y(new_n11893_));
  AOI21X1  g09457(.A0(new_n11893_), .A1(new_n11890_), .B0(pi0829), .Y(new_n11894_));
  AOI21X1  g09458(.A0(new_n11884_), .A1(pi1092), .B0(new_n5237_), .Y(new_n11895_));
  OR2X1    g09459(.A(new_n11895_), .B(new_n10213_), .Y(new_n11896_));
  OAI21X1  g09460(.A0(new_n11896_), .A1(new_n11894_), .B0(new_n11889_), .Y(new_n11897_));
  AOI21X1  g09461(.A0(new_n11897_), .A1(pi1091), .B0(pi0120), .Y(new_n11898_));
  OAI21X1  g09462(.A0(new_n11898_), .A1(new_n11882_), .B0(new_n11888_), .Y(new_n11899_));
  MX2X1    g09463(.A(new_n11899_), .B(new_n11880_), .S0(new_n5023_), .Y(new_n11900_));
  MX2X1    g09464(.A(new_n11900_), .B(new_n11880_), .S0(new_n11881_), .Y(new_n11901_));
  OAI22X1  g09465(.A0(new_n11901_), .A1(pi0642), .B0(new_n11880_), .B1(new_n11839_), .Y(new_n11902_));
  MX2X1    g09466(.A(new_n11902_), .B(new_n11825_), .S0(pi0614), .Y(new_n11903_));
  MX2X1    g09467(.A(new_n11903_), .B(new_n11825_), .S0(pi0616), .Y(new_n11904_));
  NOR2X1   g09468(.A(new_n5020_), .B(pi0614), .Y(new_n11905_));
  OAI21X1  g09469(.A0(new_n11880_), .A1(new_n11871_), .B0(new_n11905_), .Y(new_n11906_));
  AOI21X1  g09470(.A0(new_n11902_), .A1(new_n11871_), .B0(new_n11906_), .Y(new_n11907_));
  AND3X1   g09471(.A(new_n11900_), .B(new_n5020_), .C(new_n11838_), .Y(new_n11908_));
  INVX1    g09472(.A(new_n11882_), .Y(new_n11909_));
  AOI21X1  g09473(.A0(new_n11886_), .A1(new_n10082_), .B0(new_n11832_), .Y(new_n11910_));
  AND3X1   g09474(.A(new_n11826_), .B(new_n2720_), .C(new_n5922_), .Y(new_n11911_));
  OAI21X1  g09475(.A0(new_n11885_), .A1(new_n11883_), .B0(new_n5237_), .Y(new_n11912_));
  NOR2X1   g09476(.A(new_n11895_), .B(new_n10213_), .Y(new_n11913_));
  AOI21X1  g09477(.A0(new_n11913_), .A1(new_n11912_), .B0(new_n11911_), .Y(new_n11914_));
  OAI21X1  g09478(.A0(new_n11914_), .A1(new_n2702_), .B0(new_n10082_), .Y(new_n11915_));
  AOI21X1  g09479(.A0(new_n11915_), .A1(new_n11909_), .B0(new_n11910_), .Y(new_n11916_));
  MX2X1    g09480(.A(new_n11916_), .B(new_n11825_), .S0(new_n5023_), .Y(new_n11917_));
  NOR3X1   g09481(.A(new_n11872_), .B(new_n11867_), .C(new_n11838_), .Y(new_n11918_));
  INVX1    g09482(.A(new_n11918_), .Y(new_n11919_));
  AOI21X1  g09483(.A0(new_n11917_), .A1(pi0680), .B0(new_n11919_), .Y(new_n11920_));
  NOR4X1   g09484(.A(new_n11863_), .B(new_n11824_), .C(new_n2725_), .D(new_n11838_), .Y(new_n11921_));
  OR2X1    g09485(.A(new_n11921_), .B(new_n11920_), .Y(new_n11922_));
  NOR4X1   g09486(.A(new_n11922_), .B(new_n11908_), .C(new_n11907_), .D(pi0681), .Y(new_n11923_));
  AOI21X1  g09487(.A0(new_n11904_), .A1(pi0681), .B0(new_n11923_), .Y(new_n11924_));
  MX2X1    g09488(.A(new_n11899_), .B(new_n11880_), .S0(new_n5048_), .Y(new_n11925_));
  MX2X1    g09489(.A(new_n11925_), .B(new_n11899_), .S0(new_n5018_), .Y(new_n11926_));
  NOR2X1   g09490(.A(new_n11926_), .B(new_n11859_), .Y(new_n11927_));
  AND3X1   g09491(.A(pi0680), .B(new_n11849_), .C(new_n11848_), .Y(new_n11928_));
  INVX1    g09492(.A(new_n11928_), .Y(new_n11929_));
  OAI21X1  g09493(.A0(new_n11916_), .A1(new_n11929_), .B0(new_n11859_), .Y(new_n11930_));
  AOI21X1  g09494(.A0(new_n11926_), .A1(new_n11929_), .B0(new_n11930_), .Y(new_n11931_));
  NOR2X1   g09495(.A(new_n11931_), .B(new_n11927_), .Y(new_n11932_));
  MX2X1    g09496(.A(new_n11932_), .B(new_n11924_), .S0(new_n5041_), .Y(new_n11933_));
  NOR3X1   g09497(.A(new_n11824_), .B(new_n2952_), .C(new_n2725_), .Y(new_n11934_));
  OR2X1    g09498(.A(new_n11934_), .B(pi0223), .Y(new_n11935_));
  AOI21X1  g09499(.A0(new_n11933_), .A1(new_n2952_), .B0(new_n11935_), .Y(new_n11936_));
  OAI21X1  g09500(.A0(new_n11936_), .A1(new_n11879_), .B0(new_n2933_), .Y(new_n11937_));
  MX2X1    g09501(.A(new_n11917_), .B(new_n11825_), .S0(new_n11881_), .Y(new_n11938_));
  AOI21X1  g09502(.A0(new_n11938_), .A1(new_n5016_), .B0(new_n11841_), .Y(new_n11939_));
  MX2X1    g09503(.A(new_n11939_), .B(new_n11880_), .S0(pi0614), .Y(new_n11940_));
  MX2X1    g09504(.A(new_n11940_), .B(new_n11880_), .S0(pi0616), .Y(new_n11941_));
  OR4X1    g09505(.A(new_n11922_), .B(new_n11908_), .C(new_n11907_), .D(pi0681), .Y(new_n11942_));
  OAI21X1  g09506(.A0(new_n11941_), .A1(new_n11859_), .B0(new_n11942_), .Y(new_n11943_));
  OAI21X1  g09507(.A0(new_n11932_), .A1(new_n5057_), .B0(new_n5055_), .Y(new_n11944_));
  AOI21X1  g09508(.A0(new_n11943_), .A1(new_n5057_), .B0(new_n11944_), .Y(new_n11945_));
  OR4X1    g09509(.A(new_n11931_), .B(new_n11927_), .C(new_n5055_), .D(new_n10044_), .Y(new_n11946_));
  NOR3X1   g09510(.A(new_n11824_), .B(new_n10045_), .C(new_n2725_), .Y(new_n11947_));
  INVX1    g09511(.A(new_n11947_), .Y(new_n11948_));
  NAND3X1  g09512(.A(new_n11948_), .B(new_n11946_), .C(new_n2934_), .Y(new_n11949_));
  AOI21X1  g09513(.A0(new_n11945_), .A1(new_n10045_), .B0(new_n11949_), .Y(new_n11950_));
  NOR3X1   g09514(.A(new_n11861_), .B(new_n11847_), .C(new_n5055_), .Y(new_n11951_));
  INVX1    g09515(.A(new_n5057_), .Y(new_n11952_));
  OR2X1    g09516(.A(new_n11861_), .B(new_n11847_), .Y(new_n11953_));
  OAI21X1  g09517(.A0(new_n11877_), .A1(new_n11952_), .B0(new_n5055_), .Y(new_n11954_));
  AOI21X1  g09518(.A0(new_n11953_), .A1(new_n11952_), .B0(new_n11954_), .Y(new_n11955_));
  NOR3X1   g09519(.A(new_n11955_), .B(new_n11951_), .C(new_n2934_), .Y(new_n11956_));
  OAI21X1  g09520(.A0(new_n11956_), .A1(new_n11950_), .B0(pi0299), .Y(new_n11957_));
  NAND2X1  g09521(.A(new_n11957_), .B(new_n11937_), .Y(new_n11958_));
  MX2X1    g09522(.A(new_n11958_), .B(new_n11822_), .S0(new_n2939_), .Y(new_n11959_));
  OR3X1    g09523(.A(new_n11807_), .B(new_n11806_), .C(pi0210), .Y(new_n11960_));
  OAI21X1  g09524(.A0(new_n11818_), .A1(new_n2777_), .B0(new_n11960_), .Y(new_n11961_));
  NAND2X1  g09525(.A(new_n11806_), .B(pi0621), .Y(new_n11962_));
  INVX1    g09526(.A(pi0621), .Y(new_n11963_));
  OR3X1    g09527(.A(new_n11817_), .B(new_n11805_), .C(new_n11963_), .Y(new_n11964_));
  MX2X1    g09528(.A(new_n11964_), .B(new_n11962_), .S0(new_n2777_), .Y(new_n11965_));
  AOI21X1  g09529(.A0(new_n11965_), .A1(pi0603), .B0(new_n11961_), .Y(new_n11966_));
  NOR2X1   g09530(.A(new_n11966_), .B(new_n2933_), .Y(new_n11967_));
  MX2X1    g09531(.A(new_n11964_), .B(new_n11962_), .S0(new_n2954_), .Y(new_n11968_));
  AOI21X1  g09532(.A0(new_n11806_), .A1(new_n11963_), .B0(new_n11807_), .Y(new_n11969_));
  NOR2X1   g09533(.A(new_n11969_), .B(pi0198), .Y(new_n11970_));
  NAND2X1  g09534(.A(new_n11813_), .B(pi0621), .Y(new_n11971_));
  AND3X1   g09535(.A(new_n11971_), .B(new_n11818_), .C(pi0198), .Y(new_n11972_));
  OAI21X1  g09536(.A0(new_n11972_), .A1(new_n11970_), .B0(new_n11881_), .Y(new_n11973_));
  AND3X1   g09537(.A(new_n11973_), .B(new_n11968_), .C(new_n2933_), .Y(new_n11974_));
  OR2X1    g09538(.A(new_n11974_), .B(new_n11967_), .Y(new_n11975_));
  MX2X1    g09539(.A(new_n11926_), .B(new_n11899_), .S0(new_n5020_), .Y(new_n11976_));
  NOR3X1   g09540(.A(new_n11824_), .B(new_n5023_), .C(new_n2725_), .Y(new_n11977_));
  AOI21X1  g09541(.A0(new_n11899_), .A1(new_n5023_), .B0(new_n11977_), .Y(new_n11978_));
  AND2X1   g09542(.A(pi1091), .B(pi0621), .Y(new_n11979_));
  INVX1    g09543(.A(new_n11979_), .Y(new_n11980_));
  NOR4X1   g09544(.A(new_n11980_), .B(new_n11898_), .C(new_n11882_), .D(new_n5048_), .Y(new_n11981_));
  NOR4X1   g09545(.A(new_n11980_), .B(new_n11824_), .C(new_n5023_), .D(new_n2725_), .Y(new_n11982_));
  OR2X1    g09546(.A(new_n11982_), .B(new_n11881_), .Y(new_n11983_));
  NOR2X1   g09547(.A(new_n11983_), .B(new_n11981_), .Y(new_n11984_));
  AOI21X1  g09548(.A0(new_n11978_), .A1(new_n11881_), .B0(new_n11984_), .Y(new_n11985_));
  OR3X1    g09549(.A(new_n11980_), .B(new_n11898_), .C(new_n11882_), .Y(new_n11986_));
  OAI21X1  g09550(.A0(new_n11910_), .A1(new_n11963_), .B0(new_n11899_), .Y(new_n11987_));
  OAI21X1  g09551(.A0(new_n11987_), .A1(pi0603), .B0(new_n11986_), .Y(new_n11988_));
  OR2X1    g09552(.A(new_n11988_), .B(new_n11985_), .Y(new_n11989_));
  AOI21X1  g09553(.A0(new_n11989_), .A1(new_n11976_), .B0(new_n5058_), .Y(new_n11990_));
  NOR2X1   g09554(.A(new_n11979_), .B(new_n11881_), .Y(new_n11991_));
  NOR3X1   g09555(.A(new_n11991_), .B(new_n11824_), .C(new_n2725_), .Y(new_n11992_));
  INVX1    g09556(.A(new_n11992_), .Y(new_n11993_));
  OR3X1    g09557(.A(new_n11980_), .B(new_n11824_), .C(new_n2725_), .Y(new_n11994_));
  AND2X1   g09558(.A(new_n11994_), .B(new_n5023_), .Y(new_n11995_));
  AOI21X1  g09559(.A0(new_n11986_), .A1(new_n5048_), .B0(new_n11995_), .Y(new_n11996_));
  OR2X1    g09560(.A(new_n11996_), .B(new_n11881_), .Y(new_n11997_));
  AND2X1   g09561(.A(new_n11997_), .B(new_n11900_), .Y(new_n11998_));
  NOR3X1   g09562(.A(pi0642), .B(pi0616), .C(pi0614), .Y(new_n11999_));
  OR4X1    g09563(.A(new_n11991_), .B(new_n11999_), .C(new_n11824_), .D(new_n2725_), .Y(new_n12000_));
  INVX1    g09564(.A(new_n11999_), .Y(new_n12001_));
  AOI21X1  g09565(.A0(new_n11825_), .A1(new_n11881_), .B0(new_n12001_), .Y(new_n12002_));
  OAI21X1  g09566(.A0(new_n11996_), .A1(new_n11881_), .B0(new_n12002_), .Y(new_n12003_));
  NAND2X1  g09567(.A(new_n12003_), .B(new_n12000_), .Y(new_n12004_));
  MX2X1    g09568(.A(new_n12004_), .B(new_n11998_), .S0(new_n5020_), .Y(new_n12005_));
  OAI21X1  g09569(.A0(new_n12005_), .A1(new_n5059_), .B0(new_n10045_), .Y(new_n12006_));
  OAI22X1  g09570(.A0(new_n12006_), .A1(new_n11990_), .B0(new_n11993_), .B1(new_n10045_), .Y(new_n12007_));
  AND2X1   g09571(.A(new_n11843_), .B(new_n11842_), .Y(new_n12008_));
  OR4X1    g09572(.A(new_n11830_), .B(new_n11827_), .C(new_n2702_), .D(new_n11963_), .Y(new_n12009_));
  AOI21X1  g09573(.A0(new_n12009_), .A1(new_n5048_), .B0(new_n11995_), .Y(new_n12010_));
  OR2X1    g09574(.A(new_n12010_), .B(new_n11881_), .Y(new_n12011_));
  AND3X1   g09575(.A(new_n12011_), .B(new_n12008_), .C(new_n5020_), .Y(new_n12012_));
  INVX1    g09576(.A(new_n12012_), .Y(new_n12013_));
  OAI21X1  g09577(.A0(new_n12010_), .A1(new_n11881_), .B0(new_n12002_), .Y(new_n12014_));
  AND2X1   g09578(.A(new_n12014_), .B(new_n12000_), .Y(new_n12015_));
  OAI21X1  g09579(.A0(new_n12015_), .A1(new_n5020_), .B0(new_n12013_), .Y(new_n12016_));
  OR2X1    g09580(.A(new_n12016_), .B(new_n5059_), .Y(new_n12017_));
  NOR2X1   g09581(.A(new_n11991_), .B(new_n2725_), .Y(new_n12018_));
  INVX1    g09582(.A(new_n12018_), .Y(new_n12019_));
  NOR2X1   g09583(.A(new_n12019_), .B(new_n11836_), .Y(new_n12020_));
  OAI21X1  g09584(.A0(new_n11831_), .A1(new_n5348_), .B0(new_n12020_), .Y(new_n12021_));
  OAI21X1  g09585(.A0(new_n11834_), .A1(new_n11831_), .B0(new_n12018_), .Y(new_n12022_));
  AND2X1   g09586(.A(new_n12022_), .B(new_n5020_), .Y(new_n12023_));
  AOI21X1  g09587(.A0(new_n12021_), .A1(new_n5262_), .B0(new_n12023_), .Y(new_n12024_));
  INVX1    g09588(.A(new_n12024_), .Y(new_n12025_));
  AOI21X1  g09589(.A0(new_n12025_), .A1(new_n5059_), .B0(new_n2934_), .Y(new_n12026_));
  AOI22X1  g09590(.A0(new_n12026_), .A1(new_n12017_), .B0(new_n12007_), .B1(new_n2934_), .Y(new_n12027_));
  AOI21X1  g09591(.A0(new_n11989_), .A1(new_n11976_), .B0(new_n5041_), .Y(new_n12028_));
  OAI21X1  g09592(.A0(new_n12005_), .A1(new_n5042_), .B0(new_n2952_), .Y(new_n12029_));
  OAI22X1  g09593(.A0(new_n12029_), .A1(new_n12028_), .B0(new_n11993_), .B1(new_n2952_), .Y(new_n12030_));
  OR2X1    g09594(.A(new_n12016_), .B(new_n5042_), .Y(new_n12031_));
  AOI21X1  g09595(.A0(new_n12025_), .A1(new_n5042_), .B0(new_n2940_), .Y(new_n12032_));
  AOI22X1  g09596(.A0(new_n12032_), .A1(new_n12031_), .B0(new_n12030_), .B1(new_n2940_), .Y(new_n12033_));
  MX2X1    g09597(.A(new_n12033_), .B(new_n12027_), .S0(pi0299), .Y(new_n12034_));
  AND2X1   g09598(.A(new_n12034_), .B(pi0039), .Y(new_n12035_));
  AOI21X1  g09599(.A0(new_n11975_), .A1(new_n2939_), .B0(new_n12035_), .Y(new_n12036_));
  AOI21X1  g09600(.A0(new_n12036_), .A1(new_n11772_), .B0(pi0140), .Y(new_n12037_));
  OAI21X1  g09601(.A0(new_n11959_), .A1(new_n11772_), .B0(new_n12037_), .Y(new_n12038_));
  OR2X1    g09602(.A(new_n11969_), .B(pi0198), .Y(new_n12039_));
  NAND3X1  g09603(.A(new_n11971_), .B(new_n11818_), .C(pi0198), .Y(new_n12040_));
  AOI21X1  g09604(.A0(new_n12040_), .A1(new_n12039_), .B0(new_n11881_), .Y(new_n12041_));
  AND2X1   g09605(.A(new_n11969_), .B(new_n2777_), .Y(new_n12042_));
  AOI21X1  g09606(.A0(new_n11971_), .A1(new_n11818_), .B0(new_n2777_), .Y(new_n12043_));
  NOR3X1   g09607(.A(new_n12043_), .B(new_n12042_), .C(new_n11881_), .Y(new_n12044_));
  MX2X1    g09608(.A(new_n12044_), .B(new_n12041_), .S0(new_n2933_), .Y(new_n12045_));
  NOR2X1   g09609(.A(new_n12045_), .B(pi0039), .Y(new_n12046_));
  NAND2X1  g09610(.A(new_n11991_), .B(new_n11900_), .Y(new_n12047_));
  INVX1    g09611(.A(new_n11991_), .Y(new_n12048_));
  NOR3X1   g09612(.A(new_n12048_), .B(new_n11824_), .C(new_n2725_), .Y(new_n12049_));
  INVX1    g09613(.A(new_n12049_), .Y(new_n12050_));
  MX2X1    g09614(.A(new_n12050_), .B(new_n12047_), .S0(new_n11999_), .Y(new_n12051_));
  MX2X1    g09615(.A(new_n12051_), .B(new_n12047_), .S0(new_n5020_), .Y(new_n12052_));
  AND2X1   g09616(.A(new_n11991_), .B(new_n11976_), .Y(new_n12053_));
  OAI21X1  g09617(.A0(new_n12053_), .A1(new_n5058_), .B0(new_n10045_), .Y(new_n12054_));
  AOI21X1  g09618(.A0(new_n12052_), .A1(new_n5058_), .B0(new_n12054_), .Y(new_n12055_));
  NOR4X1   g09619(.A(new_n11979_), .B(new_n5032_), .C(new_n5024_), .D(new_n11881_), .Y(new_n12056_));
  INVX1    g09620(.A(new_n12056_), .Y(new_n12057_));
  NOR3X1   g09621(.A(new_n12057_), .B(new_n11824_), .C(new_n10045_), .Y(new_n12058_));
  OR2X1    g09622(.A(new_n12058_), .B(pi0215), .Y(new_n12059_));
  AND2X1   g09623(.A(new_n12049_), .B(new_n11842_), .Y(new_n12060_));
  NOR4X1   g09624(.A(new_n12001_), .B(new_n11834_), .C(new_n11831_), .D(new_n5023_), .Y(new_n12061_));
  NOR4X1   g09625(.A(new_n12061_), .B(new_n12050_), .C(new_n11836_), .D(new_n5020_), .Y(new_n12062_));
  OAI22X1  g09626(.A0(new_n12062_), .A1(new_n12060_), .B0(new_n11837_), .B1(new_n5058_), .Y(new_n12063_));
  AOI21X1  g09627(.A0(new_n12063_), .A1(pi0215), .B0(new_n2933_), .Y(new_n12064_));
  OAI21X1  g09628(.A0(new_n12059_), .A1(new_n12055_), .B0(new_n12064_), .Y(new_n12065_));
  NOR4X1   g09629(.A(new_n12048_), .B(new_n11824_), .C(new_n2952_), .D(new_n2725_), .Y(new_n12066_));
  OR2X1    g09630(.A(new_n12066_), .B(pi0223), .Y(new_n12067_));
  OAI21X1  g09631(.A0(new_n12053_), .A1(new_n5041_), .B0(new_n2952_), .Y(new_n12068_));
  AOI21X1  g09632(.A0(new_n12052_), .A1(new_n5041_), .B0(new_n12068_), .Y(new_n12069_));
  OAI22X1  g09633(.A0(new_n12062_), .A1(new_n12060_), .B0(new_n11837_), .B1(new_n5041_), .Y(new_n12070_));
  AOI21X1  g09634(.A0(new_n12070_), .A1(pi0223), .B0(pi0299), .Y(new_n12071_));
  OAI21X1  g09635(.A0(new_n12069_), .A1(new_n12067_), .B0(new_n12071_), .Y(new_n12072_));
  AND2X1   g09636(.A(new_n12072_), .B(new_n12065_), .Y(new_n12073_));
  AOI21X1  g09637(.A0(new_n12073_), .A1(pi0039), .B0(new_n12046_), .Y(new_n12074_));
  NAND3X1  g09638(.A(new_n12074_), .B(new_n11772_), .C(pi0140), .Y(new_n12075_));
  AND2X1   g09639(.A(new_n12075_), .B(new_n12038_), .Y(new_n12076_));
  NOR4X1   g09640(.A(new_n2985_), .B(new_n2725_), .C(new_n2536_), .D(pi0039), .Y(new_n12077_));
  NOR2X1   g09641(.A(new_n12077_), .B(pi0140), .Y(new_n12078_));
  NOR4X1   g09642(.A(new_n12057_), .B(new_n2985_), .C(new_n2536_), .D(pi0039), .Y(new_n12079_));
  AOI21X1  g09643(.A0(new_n12079_), .A1(new_n11772_), .B0(new_n12078_), .Y(new_n12080_));
  MX2X1    g09644(.A(new_n12080_), .B(new_n12076_), .S0(new_n2979_), .Y(new_n12081_));
  OR2X1    g09645(.A(new_n12081_), .B(new_n11771_), .Y(new_n12082_));
  NOR2X1   g09646(.A(new_n11863_), .B(new_n5019_), .Y(new_n12083_));
  AND2X1   g09647(.A(pi1091), .B(pi0665), .Y(new_n12084_));
  NOR2X1   g09648(.A(new_n12084_), .B(new_n11991_), .Y(new_n12085_));
  OR3X1    g09649(.A(new_n12085_), .B(new_n11824_), .C(new_n2725_), .Y(new_n12086_));
  AND2X1   g09650(.A(new_n12086_), .B(pi0616), .Y(new_n12087_));
  AND2X1   g09651(.A(new_n12086_), .B(pi0614), .Y(new_n12088_));
  INVX1    g09652(.A(new_n12088_), .Y(new_n12089_));
  AND2X1   g09653(.A(new_n12086_), .B(pi0642), .Y(new_n12090_));
  INVX1    g09654(.A(pi0665), .Y(new_n12091_));
  NOR4X1   g09655(.A(new_n11830_), .B(new_n11827_), .C(new_n2702_), .D(new_n12091_), .Y(new_n12092_));
  NOR2X1   g09656(.A(new_n12050_), .B(new_n11835_), .Y(new_n12093_));
  NOR2X1   g09657(.A(new_n12093_), .B(new_n12092_), .Y(new_n12094_));
  INVX1    g09658(.A(new_n12084_), .Y(new_n12095_));
  OR4X1    g09659(.A(new_n12095_), .B(new_n11824_), .C(new_n5023_), .D(new_n2725_), .Y(new_n12096_));
  OAI21X1  g09660(.A0(new_n12096_), .A1(pi0603), .B0(new_n12094_), .Y(new_n12097_));
  NOR3X1   g09661(.A(new_n12095_), .B(new_n11824_), .C(new_n2725_), .Y(new_n12098_));
  MX2X1    g09662(.A(new_n12098_), .B(new_n12092_), .S0(new_n5048_), .Y(new_n12099_));
  NOR4X1   g09663(.A(new_n12099_), .B(new_n12097_), .C(new_n12060_), .D(pi0642), .Y(new_n12100_));
  OAI21X1  g09664(.A0(new_n12100_), .A1(new_n12090_), .B0(new_n11838_), .Y(new_n12101_));
  AOI21X1  g09665(.A0(new_n12101_), .A1(new_n12089_), .B0(pi0616), .Y(new_n12102_));
  OAI21X1  g09666(.A0(new_n12102_), .A1(new_n12087_), .B0(new_n12083_), .Y(new_n12103_));
  NOR3X1   g09667(.A(new_n12099_), .B(new_n12060_), .C(new_n5262_), .Y(new_n12104_));
  AOI21X1  g09668(.A0(new_n11854_), .A1(new_n5019_), .B0(new_n12104_), .Y(new_n12105_));
  AOI21X1  g09669(.A0(new_n12105_), .A1(new_n12103_), .B0(new_n5042_), .Y(new_n12106_));
  AND2X1   g09670(.A(new_n11846_), .B(new_n5019_), .Y(new_n12107_));
  INVX1    g09671(.A(new_n12083_), .Y(new_n12108_));
  OR3X1    g09672(.A(new_n12093_), .B(new_n12092_), .C(new_n5262_), .Y(new_n12109_));
  AOI21X1  g09673(.A0(new_n12084_), .A1(new_n11977_), .B0(new_n12092_), .Y(new_n12110_));
  OAI21X1  g09674(.A0(new_n12050_), .A1(new_n11836_), .B0(new_n12110_), .Y(new_n12111_));
  MX2X1    g09675(.A(new_n12111_), .B(new_n12097_), .S0(new_n11999_), .Y(new_n12112_));
  OAI21X1  g09676(.A0(new_n12112_), .A1(new_n12108_), .B0(new_n12109_), .Y(new_n12113_));
  NOR2X1   g09677(.A(new_n12113_), .B(new_n12107_), .Y(new_n12114_));
  OAI21X1  g09678(.A0(new_n12114_), .A1(new_n5041_), .B0(pi0223), .Y(new_n12115_));
  OR2X1    g09679(.A(new_n12115_), .B(new_n12106_), .Y(new_n12116_));
  INVX1    g09680(.A(new_n12087_), .Y(new_n12117_));
  INVX1    g09681(.A(new_n12090_), .Y(new_n12118_));
  OAI21X1  g09682(.A0(new_n12085_), .A1(new_n11938_), .B0(new_n5016_), .Y(new_n12119_));
  AOI21X1  g09683(.A0(new_n12119_), .A1(new_n12118_), .B0(pi0614), .Y(new_n12120_));
  OAI21X1  g09684(.A0(new_n12120_), .A1(new_n12088_), .B0(new_n11871_), .Y(new_n12121_));
  AOI21X1  g09685(.A0(new_n12121_), .A1(new_n12117_), .B0(new_n12108_), .Y(new_n12122_));
  AND3X1   g09686(.A(new_n12084_), .B(new_n11915_), .C(new_n11909_), .Y(new_n12123_));
  MX2X1    g09687(.A(new_n12123_), .B(new_n12098_), .S0(new_n5023_), .Y(new_n12124_));
  OR2X1    g09688(.A(new_n12124_), .B(pi0603), .Y(new_n12125_));
  AND2X1   g09689(.A(new_n12091_), .B(pi0603), .Y(new_n12126_));
  AOI22X1  g09690(.A0(new_n12126_), .A1(new_n11979_), .B0(new_n11917_), .B1(pi0603), .Y(new_n12127_));
  AOI21X1  g09691(.A0(new_n12127_), .A1(new_n12125_), .B0(new_n5262_), .Y(new_n12128_));
  INVX1    g09692(.A(new_n12128_), .Y(new_n12129_));
  OAI21X1  g09693(.A0(new_n11941_), .A1(pi0680), .B0(new_n12129_), .Y(new_n12130_));
  NOR3X1   g09694(.A(new_n12130_), .B(new_n12122_), .C(new_n5042_), .Y(new_n12131_));
  MX2X1    g09695(.A(new_n11978_), .B(new_n11916_), .S0(new_n5018_), .Y(new_n12132_));
  OAI21X1  g09696(.A0(new_n12085_), .A1(new_n12132_), .B0(new_n12083_), .Y(new_n12133_));
  OR2X1    g09697(.A(new_n11987_), .B(new_n11881_), .Y(new_n12134_));
  AND2X1   g09698(.A(new_n11963_), .B(pi0603), .Y(new_n12135_));
  OR4X1    g09699(.A(new_n12135_), .B(new_n12095_), .C(new_n11898_), .D(new_n11882_), .Y(new_n12136_));
  AND2X1   g09700(.A(new_n12136_), .B(new_n5020_), .Y(new_n12137_));
  AOI22X1  g09701(.A0(new_n12137_), .A1(new_n12134_), .B0(new_n12132_), .B1(new_n5019_), .Y(new_n12138_));
  NAND2X1  g09702(.A(new_n12138_), .B(new_n12133_), .Y(new_n12139_));
  OAI21X1  g09703(.A0(new_n12139_), .A1(new_n5041_), .B0(new_n2952_), .Y(new_n12140_));
  NOR3X1   g09704(.A(new_n12084_), .B(new_n11991_), .C(new_n5019_), .Y(new_n12141_));
  NOR3X1   g09705(.A(new_n12141_), .B(new_n11824_), .C(new_n2725_), .Y(new_n12142_));
  INVX1    g09706(.A(new_n12142_), .Y(new_n12143_));
  AOI21X1  g09707(.A0(new_n12143_), .A1(new_n2951_), .B0(pi0223), .Y(new_n12144_));
  OAI21X1  g09708(.A0(new_n12140_), .A1(new_n12131_), .B0(new_n12144_), .Y(new_n12145_));
  AOI21X1  g09709(.A0(new_n12145_), .A1(new_n12116_), .B0(pi0299), .Y(new_n12146_));
  NAND2X1  g09710(.A(new_n12139_), .B(new_n5059_), .Y(new_n12147_));
  OAI21X1  g09711(.A0(new_n12130_), .A1(new_n12122_), .B0(new_n5058_), .Y(new_n12148_));
  AOI21X1  g09712(.A0(new_n12148_), .A1(new_n12147_), .B0(new_n10044_), .Y(new_n12149_));
  AOI21X1  g09713(.A0(new_n12143_), .A1(new_n10044_), .B0(pi0215), .Y(new_n12150_));
  INVX1    g09714(.A(new_n12150_), .Y(new_n12151_));
  AOI21X1  g09715(.A0(new_n12105_), .A1(new_n12103_), .B0(new_n5059_), .Y(new_n12152_));
  OAI21X1  g09716(.A0(new_n12114_), .A1(new_n5058_), .B0(pi0215), .Y(new_n12153_));
  OAI22X1  g09717(.A0(new_n12153_), .A1(new_n12152_), .B0(new_n12151_), .B1(new_n12149_), .Y(new_n12154_));
  AOI21X1  g09718(.A0(new_n12154_), .A1(pi0299), .B0(new_n12146_), .Y(new_n12155_));
  OAI22X1  g09719(.A0(new_n11983_), .A1(new_n11981_), .B0(new_n11925_), .B1(pi0603), .Y(new_n12156_));
  NOR3X1   g09720(.A(new_n12084_), .B(new_n11824_), .C(new_n2725_), .Y(new_n12157_));
  OR2X1    g09721(.A(new_n11910_), .B(new_n12091_), .Y(new_n12158_));
  AOI21X1  g09722(.A0(new_n12158_), .A1(new_n11899_), .B0(new_n12157_), .Y(new_n12159_));
  NOR2X1   g09723(.A(new_n12159_), .B(new_n12156_), .Y(new_n12160_));
  OR2X1    g09724(.A(new_n12159_), .B(new_n12156_), .Y(new_n12161_));
  NOR4X1   g09725(.A(new_n11980_), .B(new_n11898_), .C(new_n11882_), .D(pi0665), .Y(new_n12162_));
  INVX1    g09726(.A(new_n12162_), .Y(new_n12163_));
  OR2X1    g09727(.A(new_n12159_), .B(new_n11978_), .Y(new_n12164_));
  MX2X1    g09728(.A(new_n12164_), .B(new_n12163_), .S0(pi0603), .Y(new_n12165_));
  AOI21X1  g09729(.A0(new_n12165_), .A1(new_n11999_), .B0(new_n12161_), .Y(new_n12166_));
  NOR2X1   g09730(.A(pi0642), .B(pi0614), .Y(new_n12167_));
  INVX1    g09731(.A(new_n12167_), .Y(new_n12168_));
  OAI21X1  g09732(.A0(new_n12165_), .A1(new_n12168_), .B0(new_n11871_), .Y(new_n12169_));
  OAI22X1  g09733(.A0(new_n12169_), .A1(new_n12166_), .B0(new_n12160_), .B1(new_n11871_), .Y(new_n12170_));
  AND3X1   g09734(.A(new_n12158_), .B(new_n11899_), .C(new_n5020_), .Y(new_n12171_));
  OAI21X1  g09735(.A0(new_n12162_), .A1(new_n11881_), .B0(new_n12171_), .Y(new_n12172_));
  AOI22X1  g09736(.A0(new_n12172_), .A1(new_n12108_), .B0(new_n12170_), .B1(new_n11867_), .Y(new_n12173_));
  NOR4X1   g09737(.A(new_n12084_), .B(new_n11991_), .C(new_n11824_), .D(new_n2725_), .Y(new_n12174_));
  INVX1    g09738(.A(new_n12174_), .Y(new_n12175_));
  AOI21X1  g09739(.A0(new_n12175_), .A1(pi0616), .B0(new_n12108_), .Y(new_n12176_));
  INVX1    g09740(.A(new_n12157_), .Y(new_n12177_));
  MX2X1    g09741(.A(new_n12177_), .B(pi0665), .S0(pi0603), .Y(new_n12178_));
  INVX1    g09742(.A(new_n12178_), .Y(new_n12179_));
  OAI21X1  g09743(.A0(new_n11996_), .A1(new_n11881_), .B0(new_n12179_), .Y(new_n12180_));
  AOI21X1  g09744(.A0(new_n12174_), .A1(new_n12168_), .B0(pi0616), .Y(new_n12181_));
  OAI21X1  g09745(.A0(new_n12180_), .A1(new_n12168_), .B0(new_n12181_), .Y(new_n12182_));
  AOI22X1  g09746(.A0(new_n12182_), .A1(new_n12176_), .B0(new_n12128_), .B1(new_n11900_), .Y(new_n12183_));
  AOI21X1  g09747(.A0(new_n12183_), .A1(new_n5058_), .B0(new_n10044_), .Y(new_n12184_));
  OAI21X1  g09748(.A0(new_n12173_), .A1(new_n5058_), .B0(new_n12184_), .Y(new_n12185_));
  AOI21X1  g09749(.A0(new_n12141_), .A1(new_n11947_), .B0(pi0215), .Y(new_n12186_));
  NOR3X1   g09750(.A(new_n12178_), .B(new_n12019_), .C(new_n11836_), .Y(new_n12187_));
  OR2X1    g09751(.A(new_n12187_), .B(new_n11871_), .Y(new_n12188_));
  OR2X1    g09752(.A(pi0616), .B(new_n11838_), .Y(new_n12189_));
  OR2X1    g09753(.A(new_n12189_), .B(new_n12187_), .Y(new_n12190_));
  INVX1    g09754(.A(new_n12187_), .Y(new_n12191_));
  AOI21X1  g09755(.A0(new_n12179_), .A1(new_n12011_), .B0(pi0642), .Y(new_n12192_));
  OAI21X1  g09756(.A0(new_n12192_), .A1(new_n12191_), .B0(new_n5017_), .Y(new_n12193_));
  NAND3X1  g09757(.A(new_n12193_), .B(new_n12190_), .C(new_n12188_), .Y(new_n12194_));
  INVX1    g09758(.A(new_n11835_), .Y(new_n12195_));
  AOI21X1  g09759(.A0(new_n12141_), .A1(new_n12195_), .B0(new_n12083_), .Y(new_n12196_));
  AOI21X1  g09760(.A0(new_n12194_), .A1(new_n11867_), .B0(new_n12196_), .Y(new_n12197_));
  OAI21X1  g09761(.A0(new_n12084_), .A1(new_n12015_), .B0(new_n11871_), .Y(new_n12198_));
  AOI22X1  g09762(.A0(new_n12198_), .A1(new_n12176_), .B0(new_n12179_), .B1(new_n12012_), .Y(new_n12199_));
  OAI21X1  g09763(.A0(new_n12199_), .A1(new_n5059_), .B0(pi0215), .Y(new_n12200_));
  AOI21X1  g09764(.A0(new_n12197_), .A1(new_n5059_), .B0(new_n12200_), .Y(new_n12201_));
  AOI21X1  g09765(.A0(new_n12186_), .A1(new_n12185_), .B0(new_n12201_), .Y(new_n12202_));
  OAI21X1  g09766(.A0(new_n12183_), .A1(new_n5042_), .B0(new_n2952_), .Y(new_n12203_));
  AOI21X1  g09767(.A0(new_n12173_), .A1(new_n5042_), .B0(new_n12203_), .Y(new_n12204_));
  NOR2X1   g09768(.A(new_n12084_), .B(new_n5019_), .Y(new_n12205_));
  OAI21X1  g09769(.A0(new_n12205_), .A1(new_n11991_), .B0(new_n2720_), .Y(new_n12206_));
  NOR3X1   g09770(.A(new_n12206_), .B(new_n11824_), .C(new_n2725_), .Y(new_n12207_));
  NOR2X1   g09771(.A(new_n12207_), .B(new_n2952_), .Y(new_n12208_));
  NOR3X1   g09772(.A(new_n12208_), .B(new_n12204_), .C(new_n12067_), .Y(new_n12209_));
  AOI21X1  g09773(.A0(new_n12199_), .A1(new_n5041_), .B0(new_n2940_), .Y(new_n12210_));
  OAI21X1  g09774(.A0(new_n12197_), .A1(new_n5041_), .B0(new_n12210_), .Y(new_n12211_));
  NAND2X1  g09775(.A(new_n12211_), .B(new_n2933_), .Y(new_n12212_));
  OAI22X1  g09776(.A0(new_n12212_), .A1(new_n12209_), .B0(new_n12202_), .B1(new_n2933_), .Y(new_n12213_));
  OAI21X1  g09777(.A0(new_n12213_), .A1(new_n7353_), .B0(pi0761), .Y(new_n12214_));
  AOI21X1  g09778(.A0(new_n12155_), .A1(new_n7353_), .B0(new_n12214_), .Y(new_n12215_));
  AOI21X1  g09779(.A0(new_n12165_), .A1(new_n12134_), .B0(new_n12001_), .Y(new_n12216_));
  NOR2X1   g09780(.A(new_n11910_), .B(new_n12091_), .Y(new_n12217_));
  OAI21X1  g09781(.A0(new_n12217_), .A1(new_n11916_), .B0(new_n12177_), .Y(new_n12218_));
  OAI21X1  g09782(.A0(new_n12218_), .A1(new_n11991_), .B0(new_n11925_), .Y(new_n12219_));
  OAI21X1  g09783(.A0(new_n12219_), .A1(new_n11999_), .B0(new_n12083_), .Y(new_n12220_));
  NOR2X1   g09784(.A(new_n12220_), .B(new_n12216_), .Y(new_n12221_));
  NOR3X1   g09785(.A(new_n12171_), .B(new_n12083_), .C(new_n12053_), .Y(new_n12222_));
  OR3X1    g09786(.A(new_n12222_), .B(new_n12221_), .C(new_n5041_), .Y(new_n12223_));
  NOR2X1   g09787(.A(new_n12135_), .B(new_n12095_), .Y(new_n12224_));
  NOR3X1   g09788(.A(new_n12224_), .B(new_n11824_), .C(new_n2725_), .Y(new_n12225_));
  AOI21X1  g09789(.A0(new_n12225_), .A1(new_n12001_), .B0(new_n12108_), .Y(new_n12226_));
  AND2X1   g09790(.A(new_n12180_), .B(new_n12047_), .Y(new_n12227_));
  OAI21X1  g09791(.A0(new_n12227_), .A1(new_n12001_), .B0(new_n12226_), .Y(new_n12228_));
  OR2X1    g09792(.A(new_n12159_), .B(new_n11917_), .Y(new_n12229_));
  AND3X1   g09793(.A(new_n12229_), .B(new_n12047_), .C(new_n5020_), .Y(new_n12230_));
  AOI21X1  g09794(.A0(new_n12051_), .A1(new_n5019_), .B0(new_n12230_), .Y(new_n12231_));
  NAND3X1  g09795(.A(new_n12231_), .B(new_n12228_), .C(new_n5041_), .Y(new_n12232_));
  AND2X1   g09796(.A(new_n12232_), .B(new_n2952_), .Y(new_n12233_));
  AND2X1   g09797(.A(new_n12233_), .B(new_n12223_), .Y(new_n12234_));
  NOR3X1   g09798(.A(new_n12234_), .B(new_n12208_), .C(pi0223), .Y(new_n12235_));
  OAI21X1  g09799(.A0(new_n11842_), .A1(new_n5348_), .B0(new_n12157_), .Y(new_n12236_));
  INVX1    g09800(.A(new_n12236_), .Y(new_n12237_));
  OAI21X1  g09801(.A0(new_n12237_), .A1(new_n12060_), .B0(new_n11999_), .Y(new_n12238_));
  AOI21X1  g09802(.A0(new_n12157_), .A1(new_n11842_), .B0(new_n11867_), .Y(new_n12239_));
  NOR2X1   g09803(.A(new_n12239_), .B(new_n5019_), .Y(new_n12240_));
  NOR3X1   g09804(.A(new_n12240_), .B(new_n12062_), .C(new_n12060_), .Y(new_n12241_));
  AOI21X1  g09805(.A0(new_n12238_), .A1(new_n12226_), .B0(new_n12241_), .Y(new_n12242_));
  NOR2X1   g09806(.A(new_n12242_), .B(new_n5042_), .Y(new_n12243_));
  OR2X1    g09807(.A(new_n12093_), .B(new_n12062_), .Y(new_n12244_));
  NOR2X1   g09808(.A(new_n12177_), .B(new_n11836_), .Y(new_n12245_));
  AND3X1   g09809(.A(new_n12245_), .B(new_n12240_), .C(new_n12237_), .Y(new_n12246_));
  NOR3X1   g09810(.A(new_n12246_), .B(new_n12244_), .C(new_n5041_), .Y(new_n12247_));
  OR2X1    g09811(.A(new_n12247_), .B(new_n2940_), .Y(new_n12248_));
  OAI21X1  g09812(.A0(new_n12248_), .A1(new_n12243_), .B0(new_n2933_), .Y(new_n12249_));
  OR2X1    g09813(.A(new_n12249_), .B(new_n12235_), .Y(new_n12250_));
  NOR3X1   g09814(.A(new_n12222_), .B(new_n12221_), .C(new_n5058_), .Y(new_n12251_));
  AND3X1   g09815(.A(new_n12231_), .B(new_n12228_), .C(new_n5058_), .Y(new_n12252_));
  OAI21X1  g09816(.A0(new_n12252_), .A1(new_n12251_), .B0(new_n10045_), .Y(new_n12253_));
  AOI21X1  g09817(.A0(new_n12207_), .A1(new_n10044_), .B0(pi0215), .Y(new_n12254_));
  NOR2X1   g09818(.A(new_n12246_), .B(new_n12244_), .Y(new_n12255_));
  OAI21X1  g09819(.A0(new_n12255_), .A1(new_n5058_), .B0(pi0215), .Y(new_n12256_));
  AOI21X1  g09820(.A0(new_n12242_), .A1(new_n5058_), .B0(new_n12256_), .Y(new_n12257_));
  AOI21X1  g09821(.A0(new_n12254_), .A1(new_n12253_), .B0(new_n12257_), .Y(new_n12258_));
  OR2X1    g09822(.A(new_n12258_), .B(new_n2933_), .Y(new_n12259_));
  AND2X1   g09823(.A(new_n12259_), .B(new_n12250_), .Y(new_n12260_));
  AOI21X1  g09824(.A0(new_n12048_), .A1(new_n11926_), .B0(pi0680), .Y(new_n12261_));
  INVX1    g09825(.A(new_n12123_), .Y(new_n12262_));
  OAI22X1  g09826(.A0(new_n12262_), .A1(new_n5352_), .B0(new_n12096_), .B1(new_n5018_), .Y(new_n12263_));
  AOI21X1  g09827(.A0(new_n12263_), .A1(new_n12224_), .B0(new_n12108_), .Y(new_n12264_));
  OR4X1    g09828(.A(new_n12264_), .B(new_n12261_), .C(new_n12137_), .D(new_n5041_), .Y(new_n12265_));
  AND3X1   g09829(.A(new_n12003_), .B(new_n12000_), .C(new_n5019_), .Y(new_n12266_));
  OR2X1    g09830(.A(new_n12095_), .B(new_n12003_), .Y(new_n12267_));
  NOR4X1   g09831(.A(new_n12135_), .B(new_n12095_), .C(new_n11824_), .D(new_n2725_), .Y(new_n12268_));
  AOI21X1  g09832(.A0(new_n12268_), .A1(new_n12001_), .B0(new_n12108_), .Y(new_n12269_));
  AND2X1   g09833(.A(new_n12269_), .B(new_n12267_), .Y(new_n12270_));
  AOI21X1  g09834(.A0(new_n12224_), .A1(new_n12124_), .B0(new_n5262_), .Y(new_n12271_));
  OR4X1    g09835(.A(new_n12271_), .B(new_n12270_), .C(new_n12266_), .D(new_n5042_), .Y(new_n12272_));
  AOI21X1  g09836(.A0(new_n12272_), .A1(new_n12265_), .B0(new_n2951_), .Y(new_n12273_));
  OR2X1    g09837(.A(new_n11826_), .B(pi0120), .Y(new_n12274_));
  INVX1    g09838(.A(new_n12205_), .Y(new_n12275_));
  AND3X1   g09839(.A(new_n12275_), .B(new_n12048_), .C(new_n11828_), .Y(new_n12276_));
  NAND3X1  g09840(.A(new_n12276_), .B(new_n12274_), .C(new_n2951_), .Y(new_n12277_));
  AND2X1   g09841(.A(new_n12277_), .B(new_n2940_), .Y(new_n12278_));
  INVX1    g09842(.A(new_n12278_), .Y(new_n12279_));
  INVX1    g09843(.A(new_n12099_), .Y(new_n12280_));
  OR3X1    g09844(.A(new_n12205_), .B(new_n12015_), .C(new_n5020_), .Y(new_n12281_));
  OAI21X1  g09845(.A0(pi0621), .A1(new_n11881_), .B0(new_n5020_), .Y(new_n12282_));
  OAI21X1  g09846(.A0(new_n12282_), .A1(new_n12280_), .B0(new_n12281_), .Y(new_n12283_));
  AND2X1   g09847(.A(new_n12283_), .B(new_n5041_), .Y(new_n12284_));
  OAI21X1  g09848(.A0(new_n12110_), .A1(new_n12015_), .B0(new_n12083_), .Y(new_n12285_));
  OAI22X1  g09849(.A0(new_n12092_), .A1(new_n5019_), .B0(pi0621), .B1(new_n11881_), .Y(new_n12286_));
  AOI22X1  g09850(.A0(new_n12286_), .A1(new_n5020_), .B0(new_n12021_), .B1(new_n5019_), .Y(new_n12287_));
  NAND2X1  g09851(.A(new_n12287_), .B(new_n12285_), .Y(new_n12288_));
  OAI21X1  g09852(.A0(new_n12288_), .A1(new_n5041_), .B0(pi0223), .Y(new_n12289_));
  OAI22X1  g09853(.A0(new_n12289_), .A1(new_n12284_), .B0(new_n12279_), .B1(new_n12273_), .Y(new_n12290_));
  AND2X1   g09854(.A(new_n12290_), .B(new_n2933_), .Y(new_n12291_));
  OR4X1    g09855(.A(new_n12264_), .B(new_n12261_), .C(new_n12137_), .D(new_n5058_), .Y(new_n12292_));
  OR4X1    g09856(.A(new_n12271_), .B(new_n12270_), .C(new_n12266_), .D(new_n5059_), .Y(new_n12293_));
  AOI21X1  g09857(.A0(new_n12293_), .A1(new_n12292_), .B0(new_n10044_), .Y(new_n12294_));
  AND3X1   g09858(.A(new_n12276_), .B(new_n12274_), .C(new_n10044_), .Y(new_n12295_));
  NOR2X1   g09859(.A(new_n12295_), .B(pi0215), .Y(new_n12296_));
  INVX1    g09860(.A(new_n12296_), .Y(new_n12297_));
  AND2X1   g09861(.A(new_n12283_), .B(new_n5058_), .Y(new_n12298_));
  OAI21X1  g09862(.A0(new_n12288_), .A1(new_n5058_), .B0(pi0215), .Y(new_n12299_));
  OAI22X1  g09863(.A0(new_n12299_), .A1(new_n12298_), .B0(new_n12297_), .B1(new_n12294_), .Y(new_n12300_));
  AOI21X1  g09864(.A0(new_n12300_), .A1(pi0299), .B0(new_n12291_), .Y(new_n12301_));
  OAI21X1  g09865(.A0(new_n12301_), .A1(pi0140), .B0(new_n11772_), .Y(new_n12302_));
  AOI21X1  g09866(.A0(new_n12260_), .A1(pi0140), .B0(new_n12302_), .Y(new_n12303_));
  OAI21X1  g09867(.A0(new_n12303_), .A1(new_n12215_), .B0(pi0039), .Y(new_n12304_));
  OR3X1    g09868(.A(new_n11807_), .B(new_n11806_), .C(pi0198), .Y(new_n12305_));
  OAI21X1  g09869(.A0(new_n11818_), .A1(new_n2954_), .B0(new_n12305_), .Y(new_n12306_));
  OR3X1    g09870(.A(new_n11817_), .B(new_n11805_), .C(new_n12091_), .Y(new_n12307_));
  AND2X1   g09871(.A(new_n11806_), .B(pi0665), .Y(new_n12308_));
  INVX1    g09872(.A(new_n12308_), .Y(new_n12309_));
  MX2X1    g09873(.A(new_n12309_), .B(new_n12307_), .S0(pi0198), .Y(new_n12310_));
  AOI21X1  g09874(.A0(new_n12310_), .A1(pi0680), .B0(new_n12306_), .Y(new_n12311_));
  MX2X1    g09875(.A(new_n12309_), .B(new_n12307_), .S0(pi0210), .Y(new_n12312_));
  AOI21X1  g09876(.A0(new_n12312_), .A1(pi0680), .B0(new_n11961_), .Y(new_n12313_));
  MX2X1    g09877(.A(new_n12313_), .B(new_n12311_), .S0(new_n2933_), .Y(new_n12314_));
  AOI21X1  g09878(.A0(new_n12045_), .A1(pi0680), .B0(new_n12314_), .Y(new_n12315_));
  AND2X1   g09879(.A(pi0665), .B(pi0603), .Y(new_n12316_));
  AOI21X1  g09880(.A0(new_n11806_), .A1(new_n12091_), .B0(new_n11807_), .Y(new_n12317_));
  NAND2X1  g09881(.A(new_n12317_), .B(new_n2954_), .Y(new_n12318_));
  OR2X1    g09882(.A(new_n11817_), .B(new_n11805_), .Y(new_n12319_));
  AND2X1   g09883(.A(new_n12319_), .B(new_n11813_), .Y(new_n12320_));
  AND2X1   g09884(.A(new_n11813_), .B(pi0665), .Y(new_n12321_));
  OAI21X1  g09885(.A0(new_n12321_), .A1(new_n12320_), .B0(pi0198), .Y(new_n12322_));
  AOI21X1  g09886(.A0(new_n12322_), .A1(new_n12318_), .B0(pi0603), .Y(new_n12323_));
  AND2X1   g09887(.A(new_n11968_), .B(pi0603), .Y(new_n12324_));
  OR4X1    g09888(.A(new_n12324_), .B(new_n12323_), .C(new_n12316_), .D(new_n5019_), .Y(new_n12325_));
  OAI21X1  g09889(.A0(new_n12321_), .A1(new_n12320_), .B0(pi0210), .Y(new_n12326_));
  NAND2X1  g09890(.A(new_n12317_), .B(new_n2777_), .Y(new_n12327_));
  AOI21X1  g09891(.A0(new_n12327_), .A1(new_n12326_), .B0(pi0603), .Y(new_n12328_));
  AOI21X1  g09892(.A0(new_n11965_), .A1(pi0603), .B0(new_n12316_), .Y(new_n12329_));
  INVX1    g09893(.A(new_n12329_), .Y(new_n12330_));
  OR3X1    g09894(.A(new_n12330_), .B(new_n12328_), .C(new_n5019_), .Y(new_n12331_));
  MX2X1    g09895(.A(new_n12331_), .B(new_n12325_), .S0(new_n2933_), .Y(new_n12332_));
  AOI21X1  g09896(.A0(new_n12332_), .A1(pi0140), .B0(new_n11772_), .Y(new_n12333_));
  OAI21X1  g09897(.A0(new_n12315_), .A1(pi0140), .B0(new_n12333_), .Y(new_n12334_));
  NOR3X1   g09898(.A(new_n11817_), .B(new_n11805_), .C(new_n12091_), .Y(new_n12335_));
  MX2X1    g09899(.A(new_n12308_), .B(new_n12335_), .S0(pi0198), .Y(new_n12336_));
  OAI21X1  g09900(.A0(new_n12336_), .A1(new_n5019_), .B0(new_n11820_), .Y(new_n12337_));
  MX2X1    g09901(.A(new_n12308_), .B(new_n12335_), .S0(pi0210), .Y(new_n12338_));
  OAI21X1  g09902(.A0(new_n12338_), .A1(new_n5019_), .B0(new_n11819_), .Y(new_n12339_));
  MX2X1    g09903(.A(new_n12339_), .B(new_n12337_), .S0(new_n2933_), .Y(new_n12340_));
  OR4X1    g09904(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0140), .Y(new_n12341_));
  AND3X1   g09905(.A(new_n12322_), .B(new_n12318_), .C(pi0680), .Y(new_n12342_));
  AND3X1   g09906(.A(new_n12327_), .B(new_n12326_), .C(pi0680), .Y(new_n12343_));
  MX2X1    g09907(.A(new_n12343_), .B(new_n12342_), .S0(new_n2933_), .Y(new_n12344_));
  OR3X1    g09908(.A(new_n12344_), .B(new_n12045_), .C(new_n7353_), .Y(new_n12345_));
  AND3X1   g09909(.A(new_n12345_), .B(new_n12341_), .C(new_n11772_), .Y(new_n12346_));
  NOR2X1   g09910(.A(new_n12346_), .B(pi0039), .Y(new_n12347_));
  AOI21X1  g09911(.A0(new_n12347_), .A1(new_n12334_), .B0(pi0038), .Y(new_n12348_));
  OR4X1    g09912(.A(new_n12206_), .B(new_n2985_), .C(new_n2536_), .D(new_n7353_), .Y(new_n12349_));
  AND2X1   g09913(.A(new_n12349_), .B(new_n11772_), .Y(new_n12350_));
  OAI21X1  g09914(.A0(new_n12276_), .A1(pi0140), .B0(new_n12350_), .Y(new_n12351_));
  INVX1    g09915(.A(new_n12141_), .Y(new_n12352_));
  NOR4X1   g09916(.A(new_n12352_), .B(new_n2985_), .C(new_n2725_), .D(new_n2536_), .Y(new_n12353_));
  NOR2X1   g09917(.A(new_n12353_), .B(new_n11772_), .Y(new_n12354_));
  OAI21X1  g09918(.A0(new_n11828_), .A1(pi0140), .B0(new_n12354_), .Y(new_n12355_));
  AOI21X1  g09919(.A0(new_n12355_), .A1(new_n12351_), .B0(pi0039), .Y(new_n12356_));
  AND2X1   g09920(.A(pi0140), .B(pi0039), .Y(new_n12357_));
  NOR3X1   g09921(.A(new_n12357_), .B(new_n12356_), .C(new_n2979_), .Y(new_n12358_));
  AOI21X1  g09922(.A0(new_n12348_), .A1(new_n12304_), .B0(new_n12358_), .Y(new_n12359_));
  OR2X1    g09923(.A(new_n12359_), .B(pi0738), .Y(new_n12360_));
  AND2X1   g09924(.A(new_n12360_), .B(new_n3103_), .Y(new_n12361_));
  AOI22X1  g09925(.A0(new_n12361_), .A1(new_n12082_), .B0(new_n11770_), .B1(pi0140), .Y(new_n12362_));
  INVX1    g09926(.A(pi0625), .Y(new_n12363_));
  INVX1    g09927(.A(pi1153), .Y(new_n12364_));
  MX2X1    g09928(.A(new_n12081_), .B(pi0140), .S0(new_n11770_), .Y(new_n12365_));
  OAI21X1  g09929(.A0(new_n12365_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n12366_));
  AOI21X1  g09930(.A0(new_n12362_), .A1(new_n12363_), .B0(new_n12366_), .Y(new_n12367_));
  INVX1    g09931(.A(pi0608), .Y(new_n12368_));
  NOR4X1   g09932(.A(new_n12275_), .B(new_n11824_), .C(new_n2952_), .D(new_n2725_), .Y(new_n12369_));
  MX2X1    g09933(.A(new_n12229_), .B(new_n12177_), .S0(new_n5348_), .Y(new_n12370_));
  OAI21X1  g09934(.A0(new_n12159_), .A1(new_n11917_), .B0(new_n11863_), .Y(new_n12371_));
  NAND2X1  g09935(.A(new_n12371_), .B(pi0680), .Y(new_n12372_));
  AOI21X1  g09936(.A0(new_n12370_), .A1(new_n11867_), .B0(new_n12372_), .Y(new_n12373_));
  OR2X1    g09937(.A(new_n12373_), .B(new_n5042_), .Y(new_n12374_));
  AND2X1   g09938(.A(new_n12205_), .B(new_n11926_), .Y(new_n12375_));
  AOI21X1  g09939(.A0(new_n12375_), .A1(new_n11867_), .B0(new_n12171_), .Y(new_n12376_));
  AOI21X1  g09940(.A0(new_n12376_), .A1(new_n5042_), .B0(new_n2951_), .Y(new_n12377_));
  AOI21X1  g09941(.A0(new_n12377_), .A1(new_n12374_), .B0(new_n12369_), .Y(new_n12378_));
  OR2X1    g09942(.A(new_n12378_), .B(pi0223), .Y(new_n12379_));
  AND2X1   g09943(.A(new_n11836_), .B(new_n5042_), .Y(new_n12380_));
  NOR3X1   g09944(.A(new_n12236_), .B(new_n12380_), .C(new_n5019_), .Y(new_n12381_));
  INVX1    g09945(.A(new_n12381_), .Y(new_n12382_));
  OR3X1    g09946(.A(new_n12382_), .B(new_n12239_), .C(new_n2940_), .Y(new_n12383_));
  AND2X1   g09947(.A(new_n12383_), .B(new_n12379_), .Y(new_n12384_));
  AND2X1   g09948(.A(new_n12376_), .B(new_n5059_), .Y(new_n12385_));
  OAI21X1  g09949(.A0(new_n12373_), .A1(new_n5059_), .B0(new_n10045_), .Y(new_n12386_));
  OR4X1    g09950(.A(new_n12275_), .B(new_n11824_), .C(new_n10045_), .D(new_n2725_), .Y(new_n12387_));
  OAI21X1  g09951(.A0(new_n12386_), .A1(new_n12385_), .B0(new_n12387_), .Y(new_n12388_));
  AND2X1   g09952(.A(new_n11836_), .B(new_n5059_), .Y(new_n12389_));
  NOR3X1   g09953(.A(new_n12236_), .B(new_n12389_), .C(new_n5019_), .Y(new_n12390_));
  INVX1    g09954(.A(new_n12390_), .Y(new_n12391_));
  NOR3X1   g09955(.A(new_n12391_), .B(new_n12239_), .C(new_n2934_), .Y(new_n12392_));
  AOI21X1  g09956(.A0(new_n12388_), .A1(new_n2934_), .B0(new_n12392_), .Y(new_n12393_));
  MX2X1    g09957(.A(new_n12393_), .B(new_n12384_), .S0(new_n2933_), .Y(new_n12394_));
  NOR2X1   g09958(.A(new_n12394_), .B(new_n7353_), .Y(new_n12395_));
  AOI21X1  g09959(.A0(new_n12098_), .A1(new_n5348_), .B0(new_n5019_), .Y(new_n12396_));
  INVX1    g09960(.A(new_n12396_), .Y(new_n12397_));
  AOI21X1  g09961(.A0(new_n12124_), .A1(new_n5018_), .B0(new_n12397_), .Y(new_n12398_));
  INVX1    g09962(.A(new_n12398_), .Y(new_n12399_));
  OAI21X1  g09963(.A0(new_n11941_), .A1(pi0680), .B0(new_n12399_), .Y(new_n12400_));
  OR2X1    g09964(.A(new_n12124_), .B(new_n5019_), .Y(new_n12401_));
  AND2X1   g09965(.A(new_n12401_), .B(new_n11863_), .Y(new_n12402_));
  OAI21X1  g09966(.A0(new_n11941_), .A1(pi0680), .B0(new_n12402_), .Y(new_n12403_));
  OAI21X1  g09967(.A0(new_n12400_), .A1(new_n11863_), .B0(new_n12403_), .Y(new_n12404_));
  NOR2X1   g09968(.A(new_n11926_), .B(pi0680), .Y(new_n12405_));
  OAI21X1  g09969(.A0(new_n12262_), .A1(new_n11867_), .B0(pi0680), .Y(new_n12406_));
  AOI21X1  g09970(.A0(new_n12263_), .A1(new_n11867_), .B0(new_n12406_), .Y(new_n12407_));
  NOR2X1   g09971(.A(new_n12407_), .B(new_n12405_), .Y(new_n12408_));
  OAI21X1  g09972(.A0(new_n12408_), .A1(new_n5041_), .B0(new_n2952_), .Y(new_n12409_));
  INVX1    g09973(.A(new_n12409_), .Y(new_n12410_));
  OAI21X1  g09974(.A0(new_n12404_), .A1(new_n5042_), .B0(new_n12410_), .Y(new_n12411_));
  AOI21X1  g09975(.A0(new_n12275_), .A1(new_n11934_), .B0(pi0223), .Y(new_n12412_));
  AOI21X1  g09976(.A0(new_n12397_), .A1(new_n5262_), .B0(new_n12099_), .Y(new_n12413_));
  AOI21X1  g09977(.A0(new_n11854_), .A1(new_n5019_), .B0(new_n12413_), .Y(new_n12414_));
  AND2X1   g09978(.A(new_n12414_), .B(new_n5041_), .Y(new_n12415_));
  INVX1    g09979(.A(new_n12415_), .Y(new_n12416_));
  NOR2X1   g09980(.A(new_n12096_), .B(new_n5018_), .Y(new_n12417_));
  NOR3X1   g09981(.A(new_n12417_), .B(new_n12092_), .C(new_n5019_), .Y(new_n12418_));
  NOR3X1   g09982(.A(new_n12418_), .B(new_n12413_), .C(new_n12107_), .Y(new_n12419_));
  AOI21X1  g09983(.A0(new_n12419_), .A1(new_n5042_), .B0(new_n2940_), .Y(new_n12420_));
  AOI22X1  g09984(.A0(new_n12420_), .A1(new_n12416_), .B0(new_n12412_), .B1(new_n12411_), .Y(new_n12421_));
  OAI21X1  g09985(.A0(new_n12408_), .A1(new_n5058_), .B0(new_n10045_), .Y(new_n12422_));
  INVX1    g09986(.A(new_n12422_), .Y(new_n12423_));
  OAI21X1  g09987(.A0(new_n12404_), .A1(new_n5059_), .B0(new_n12423_), .Y(new_n12424_));
  NOR2X1   g09988(.A(new_n11824_), .B(new_n10045_), .Y(new_n12425_));
  NOR2X1   g09989(.A(new_n12205_), .B(new_n2725_), .Y(new_n12426_));
  AOI21X1  g09990(.A0(new_n12426_), .A1(new_n12425_), .B0(pi0215), .Y(new_n12427_));
  AND2X1   g09991(.A(new_n12414_), .B(new_n5058_), .Y(new_n12428_));
  INVX1    g09992(.A(new_n12428_), .Y(new_n12429_));
  AOI21X1  g09993(.A0(new_n12419_), .A1(new_n5059_), .B0(new_n2934_), .Y(new_n12430_));
  AOI22X1  g09994(.A0(new_n12430_), .A1(new_n12429_), .B0(new_n12427_), .B1(new_n12424_), .Y(new_n12431_));
  MX2X1    g09995(.A(new_n12431_), .B(new_n12421_), .S0(new_n2933_), .Y(new_n12432_));
  OAI21X1  g09996(.A0(new_n12432_), .A1(pi0140), .B0(pi0039), .Y(new_n12433_));
  OR2X1    g09997(.A(new_n12342_), .B(pi0299), .Y(new_n12434_));
  OAI21X1  g09998(.A0(new_n12343_), .A1(new_n2933_), .B0(new_n12434_), .Y(new_n12435_));
  AOI21X1  g09999(.A0(new_n12340_), .A1(new_n7353_), .B0(pi0039), .Y(new_n12436_));
  OAI21X1  g10000(.A0(new_n12435_), .A1(new_n7353_), .B0(new_n12436_), .Y(new_n12437_));
  OAI21X1  g10001(.A0(new_n12433_), .A1(new_n12395_), .B0(new_n12437_), .Y(new_n12438_));
  NOR4X1   g10002(.A(new_n12084_), .B(new_n5032_), .C(new_n5024_), .D(new_n5019_), .Y(new_n12439_));
  AOI21X1  g10003(.A0(new_n12439_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n12440_));
  INVX1    g10004(.A(new_n12440_), .Y(new_n12441_));
  OAI21X1  g10005(.A0(new_n12441_), .A1(new_n12078_), .B0(new_n11771_), .Y(new_n12442_));
  AOI21X1  g10006(.A0(new_n12438_), .A1(new_n2979_), .B0(new_n12442_), .Y(new_n12443_));
  AND2X1   g10007(.A(new_n11957_), .B(new_n11937_), .Y(new_n12444_));
  MX2X1    g10008(.A(new_n12444_), .B(new_n11821_), .S0(new_n2939_), .Y(new_n12445_));
  AND3X1   g10009(.A(new_n2982_), .B(new_n2720_), .C(new_n2939_), .Y(new_n12446_));
  MX2X1    g10010(.A(new_n12446_), .B(new_n12445_), .S0(new_n2979_), .Y(new_n12447_));
  OR2X1    g10011(.A(new_n11771_), .B(pi0140), .Y(new_n12448_));
  OAI21X1  g10012(.A0(new_n12448_), .A1(new_n12447_), .B0(new_n3103_), .Y(new_n12449_));
  OAI22X1  g10013(.A0(new_n12449_), .A1(new_n12443_), .B0(new_n3103_), .B1(new_n7353_), .Y(new_n12450_));
  AOI21X1  g10014(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0140), .Y(new_n12451_));
  AOI21X1  g10015(.A0(new_n12451_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n12452_));
  OAI21X1  g10016(.A0(new_n12450_), .A1(new_n12363_), .B0(new_n12452_), .Y(new_n12453_));
  NAND2X1  g10017(.A(new_n12453_), .B(new_n12368_), .Y(new_n12454_));
  OAI21X1  g10018(.A0(new_n12365_), .A1(pi0625), .B0(pi1153), .Y(new_n12455_));
  AOI21X1  g10019(.A0(new_n12362_), .A1(pi0625), .B0(new_n12455_), .Y(new_n12456_));
  AOI21X1  g10020(.A0(new_n12451_), .A1(pi0625), .B0(pi1153), .Y(new_n12457_));
  OAI21X1  g10021(.A0(new_n12450_), .A1(pi0625), .B0(new_n12457_), .Y(new_n12458_));
  NAND2X1  g10022(.A(new_n12458_), .B(pi0608), .Y(new_n12459_));
  OAI22X1  g10023(.A0(new_n12459_), .A1(new_n12456_), .B0(new_n12454_), .B1(new_n12367_), .Y(new_n12460_));
  MX2X1    g10024(.A(new_n12460_), .B(new_n12362_), .S0(new_n11769_), .Y(new_n12461_));
  INVX1    g10025(.A(pi0609), .Y(new_n12462_));
  INVX1    g10026(.A(pi1155), .Y(new_n12463_));
  NAND2X1  g10027(.A(new_n12458_), .B(new_n12453_), .Y(new_n12464_));
  MX2X1    g10028(.A(new_n12464_), .B(new_n12450_), .S0(new_n11769_), .Y(new_n12465_));
  OAI21X1  g10029(.A0(new_n12465_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n12466_));
  AOI21X1  g10030(.A0(new_n12461_), .A1(new_n12462_), .B0(new_n12466_), .Y(new_n12467_));
  INVX1    g10031(.A(pi0660), .Y(new_n12468_));
  INVX1    g10032(.A(new_n12451_), .Y(new_n12469_));
  XOR2X1   g10033(.A(pi1153), .B(pi0608), .Y(new_n12470_));
  AOI21X1  g10034(.A0(new_n12470_), .A1(pi0778), .B0(new_n12462_), .Y(new_n12471_));
  INVX1    g10035(.A(new_n12471_), .Y(new_n12472_));
  AND2X1   g10036(.A(new_n12470_), .B(pi0778), .Y(new_n12473_));
  INVX1    g10037(.A(new_n12473_), .Y(new_n12474_));
  AND2X1   g10038(.A(new_n12474_), .B(new_n12365_), .Y(new_n12475_));
  AOI22X1  g10039(.A0(new_n12475_), .A1(pi0609), .B0(new_n12472_), .B1(new_n12469_), .Y(new_n12476_));
  OAI21X1  g10040(.A0(new_n12476_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n12477_));
  OAI21X1  g10041(.A0(new_n12465_), .A1(pi0609), .B0(pi1155), .Y(new_n12478_));
  AOI21X1  g10042(.A0(new_n12461_), .A1(pi0609), .B0(new_n12478_), .Y(new_n12479_));
  AOI21X1  g10043(.A0(new_n12470_), .A1(pi0778), .B0(pi0609), .Y(new_n12480_));
  INVX1    g10044(.A(new_n12480_), .Y(new_n12481_));
  AOI22X1  g10045(.A0(new_n12481_), .A1(new_n12469_), .B0(new_n12475_), .B1(new_n12462_), .Y(new_n12482_));
  OAI21X1  g10046(.A0(new_n12482_), .A1(pi1155), .B0(pi0660), .Y(new_n12483_));
  OAI22X1  g10047(.A0(new_n12483_), .A1(new_n12479_), .B0(new_n12477_), .B1(new_n12467_), .Y(new_n12484_));
  MX2X1    g10048(.A(new_n12484_), .B(new_n12461_), .S0(new_n11768_), .Y(new_n12485_));
  INVX1    g10049(.A(pi0618), .Y(new_n12486_));
  INVX1    g10050(.A(pi1154), .Y(new_n12487_));
  AND2X1   g10051(.A(pi1155), .B(pi0660), .Y(new_n12488_));
  NOR2X1   g10052(.A(pi1155), .B(pi0660), .Y(new_n12489_));
  NOR3X1   g10053(.A(new_n12489_), .B(new_n12488_), .C(new_n11768_), .Y(new_n12490_));
  MX2X1    g10054(.A(new_n12465_), .B(new_n12469_), .S0(new_n12490_), .Y(new_n12491_));
  OAI21X1  g10055(.A0(new_n12491_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n12492_));
  AOI21X1  g10056(.A0(new_n12485_), .A1(new_n12486_), .B0(new_n12492_), .Y(new_n12493_));
  INVX1    g10057(.A(pi0627), .Y(new_n12494_));
  MX2X1    g10058(.A(new_n12469_), .B(new_n12365_), .S0(new_n12474_), .Y(new_n12495_));
  NAND2X1  g10059(.A(new_n12495_), .B(new_n11768_), .Y(new_n12496_));
  MX2X1    g10060(.A(new_n12482_), .B(new_n12476_), .S0(pi1155), .Y(new_n12497_));
  OAI21X1  g10061(.A0(new_n12497_), .A1(new_n11768_), .B0(new_n12496_), .Y(new_n12498_));
  AOI21X1  g10062(.A0(new_n12451_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n12499_));
  OAI21X1  g10063(.A0(new_n12498_), .A1(new_n12486_), .B0(new_n12499_), .Y(new_n12500_));
  NAND2X1  g10064(.A(new_n12500_), .B(new_n12494_), .Y(new_n12501_));
  OAI21X1  g10065(.A0(new_n12491_), .A1(pi0618), .B0(pi1154), .Y(new_n12502_));
  AOI21X1  g10066(.A0(new_n12485_), .A1(pi0618), .B0(new_n12502_), .Y(new_n12503_));
  AOI21X1  g10067(.A0(new_n12451_), .A1(pi0618), .B0(pi1154), .Y(new_n12504_));
  OAI21X1  g10068(.A0(new_n12498_), .A1(pi0618), .B0(new_n12504_), .Y(new_n12505_));
  NAND2X1  g10069(.A(new_n12505_), .B(pi0627), .Y(new_n12506_));
  OAI22X1  g10070(.A0(new_n12506_), .A1(new_n12503_), .B0(new_n12501_), .B1(new_n12493_), .Y(new_n12507_));
  MX2X1    g10071(.A(new_n12507_), .B(new_n12485_), .S0(new_n11767_), .Y(new_n12508_));
  INVX1    g10072(.A(pi0619), .Y(new_n12509_));
  INVX1    g10073(.A(pi1159), .Y(new_n12510_));
  AND2X1   g10074(.A(pi1154), .B(pi0627), .Y(new_n12511_));
  NOR2X1   g10075(.A(pi1154), .B(pi0627), .Y(new_n12512_));
  NOR3X1   g10076(.A(new_n12512_), .B(new_n12511_), .C(new_n11767_), .Y(new_n12513_));
  MX2X1    g10077(.A(new_n12491_), .B(new_n12469_), .S0(new_n12513_), .Y(new_n12514_));
  OAI21X1  g10078(.A0(new_n12514_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n12515_));
  AOI21X1  g10079(.A0(new_n12508_), .A1(new_n12509_), .B0(new_n12515_), .Y(new_n12516_));
  INVX1    g10080(.A(pi0648), .Y(new_n12517_));
  NAND2X1  g10081(.A(new_n12505_), .B(new_n12500_), .Y(new_n12518_));
  MX2X1    g10082(.A(new_n12518_), .B(new_n12498_), .S0(new_n11767_), .Y(new_n12519_));
  AOI21X1  g10083(.A0(new_n12451_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n12520_));
  OAI21X1  g10084(.A0(new_n12519_), .A1(new_n12509_), .B0(new_n12520_), .Y(new_n12521_));
  NAND2X1  g10085(.A(new_n12521_), .B(new_n12517_), .Y(new_n12522_));
  OAI21X1  g10086(.A0(new_n12514_), .A1(pi0619), .B0(pi1159), .Y(new_n12523_));
  AOI21X1  g10087(.A0(new_n12508_), .A1(pi0619), .B0(new_n12523_), .Y(new_n12524_));
  AOI21X1  g10088(.A0(new_n12451_), .A1(pi0619), .B0(pi1159), .Y(new_n12525_));
  OAI21X1  g10089(.A0(new_n12519_), .A1(pi0619), .B0(new_n12525_), .Y(new_n12526_));
  NAND2X1  g10090(.A(new_n12526_), .B(pi0648), .Y(new_n12527_));
  OAI22X1  g10091(.A0(new_n12527_), .A1(new_n12524_), .B0(new_n12522_), .B1(new_n12516_), .Y(new_n12528_));
  MX2X1    g10092(.A(new_n12528_), .B(new_n12508_), .S0(new_n11766_), .Y(new_n12529_));
  XOR2X1   g10093(.A(pi1159), .B(new_n12517_), .Y(new_n12530_));
  NOR2X1   g10094(.A(new_n12530_), .B(new_n11766_), .Y(new_n12531_));
  MX2X1    g10095(.A(new_n12514_), .B(new_n12469_), .S0(new_n12531_), .Y(new_n12532_));
  AOI21X1  g10096(.A0(new_n12532_), .A1(pi0626), .B0(pi0641), .Y(new_n12533_));
  OAI21X1  g10097(.A0(new_n12529_), .A1(pi0626), .B0(new_n12533_), .Y(new_n12534_));
  NOR2X1   g10098(.A(pi1158), .B(pi0641), .Y(new_n12535_));
  AND2X1   g10099(.A(new_n12519_), .B(new_n11766_), .Y(new_n12536_));
  AOI21X1  g10100(.A0(new_n12526_), .A1(new_n12521_), .B0(new_n11766_), .Y(new_n12537_));
  OR3X1    g10101(.A(new_n12537_), .B(new_n12536_), .C(pi0626), .Y(new_n12538_));
  AOI21X1  g10102(.A0(new_n12451_), .A1(pi0626), .B0(pi1158), .Y(new_n12539_));
  AND2X1   g10103(.A(new_n12539_), .B(new_n12538_), .Y(new_n12540_));
  OR2X1    g10104(.A(new_n12540_), .B(new_n12535_), .Y(new_n12541_));
  INVX1    g10105(.A(pi0626), .Y(new_n12542_));
  INVX1    g10106(.A(pi0641), .Y(new_n12543_));
  AOI21X1  g10107(.A0(new_n12532_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n12544_));
  OAI21X1  g10108(.A0(new_n12529_), .A1(new_n12542_), .B0(new_n12544_), .Y(new_n12545_));
  AND2X1   g10109(.A(pi1158), .B(pi0641), .Y(new_n12546_));
  OR3X1    g10110(.A(new_n12537_), .B(new_n12536_), .C(new_n12542_), .Y(new_n12547_));
  INVX1    g10111(.A(pi1158), .Y(new_n12548_));
  AOI21X1  g10112(.A0(new_n12451_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n12549_));
  AND2X1   g10113(.A(new_n12549_), .B(new_n12547_), .Y(new_n12550_));
  OR2X1    g10114(.A(new_n12550_), .B(new_n12546_), .Y(new_n12551_));
  AOI22X1  g10115(.A0(new_n12551_), .A1(new_n12545_), .B0(new_n12541_), .B1(new_n12534_), .Y(new_n12552_));
  MX2X1    g10116(.A(new_n12552_), .B(new_n12529_), .S0(new_n11765_), .Y(new_n12553_));
  INVX1    g10117(.A(pi0628), .Y(new_n12554_));
  INVX1    g10118(.A(pi1156), .Y(new_n12555_));
  AOI22X1  g10119(.A0(new_n12549_), .A1(new_n12547_), .B0(new_n12539_), .B1(new_n12538_), .Y(new_n12556_));
  OAI21X1  g10120(.A0(new_n12537_), .A1(new_n12536_), .B0(new_n11765_), .Y(new_n12557_));
  OAI21X1  g10121(.A0(new_n12556_), .A1(new_n11765_), .B0(new_n12557_), .Y(new_n12558_));
  OAI21X1  g10122(.A0(new_n12558_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n12559_));
  AOI21X1  g10123(.A0(new_n12553_), .A1(new_n12554_), .B0(new_n12559_), .Y(new_n12560_));
  INVX1    g10124(.A(pi0629), .Y(new_n12561_));
  XOR2X1   g10125(.A(pi1158), .B(new_n12543_), .Y(new_n12562_));
  NOR2X1   g10126(.A(new_n12562_), .B(new_n11765_), .Y(new_n12563_));
  MX2X1    g10127(.A(new_n12532_), .B(new_n12469_), .S0(new_n12563_), .Y(new_n12564_));
  AOI21X1  g10128(.A0(new_n12451_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n12565_));
  OAI21X1  g10129(.A0(new_n12564_), .A1(new_n12554_), .B0(new_n12565_), .Y(new_n12566_));
  AND2X1   g10130(.A(new_n12566_), .B(new_n12561_), .Y(new_n12567_));
  INVX1    g10131(.A(new_n12567_), .Y(new_n12568_));
  OAI21X1  g10132(.A0(new_n12558_), .A1(pi0628), .B0(pi1156), .Y(new_n12569_));
  AOI21X1  g10133(.A0(new_n12553_), .A1(pi0628), .B0(new_n12569_), .Y(new_n12570_));
  AOI21X1  g10134(.A0(new_n12451_), .A1(pi0628), .B0(pi1156), .Y(new_n12571_));
  OAI21X1  g10135(.A0(new_n12564_), .A1(pi0628), .B0(new_n12571_), .Y(new_n12572_));
  AND2X1   g10136(.A(new_n12572_), .B(pi0629), .Y(new_n12573_));
  INVX1    g10137(.A(new_n12573_), .Y(new_n12574_));
  OAI22X1  g10138(.A0(new_n12574_), .A1(new_n12570_), .B0(new_n12568_), .B1(new_n12560_), .Y(new_n12575_));
  MX2X1    g10139(.A(new_n12575_), .B(new_n12553_), .S0(new_n11764_), .Y(new_n12576_));
  INVX1    g10140(.A(pi0647), .Y(new_n12577_));
  INVX1    g10141(.A(pi1157), .Y(new_n12578_));
  XOR2X1   g10142(.A(pi1156), .B(pi0629), .Y(new_n12579_));
  AND2X1   g10143(.A(new_n12579_), .B(pi0792), .Y(new_n12580_));
  MX2X1    g10144(.A(new_n12558_), .B(new_n12469_), .S0(new_n12580_), .Y(new_n12581_));
  OAI21X1  g10145(.A0(new_n12581_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n12582_));
  AOI21X1  g10146(.A0(new_n12576_), .A1(new_n12577_), .B0(new_n12582_), .Y(new_n12583_));
  AOI21X1  g10147(.A0(new_n12572_), .A1(new_n12566_), .B0(new_n11764_), .Y(new_n12584_));
  AOI21X1  g10148(.A0(new_n12564_), .A1(new_n11764_), .B0(new_n12584_), .Y(new_n12585_));
  OAI21X1  g10149(.A0(new_n12469_), .A1(pi0647), .B0(pi1157), .Y(new_n12586_));
  AOI21X1  g10150(.A0(new_n12585_), .A1(pi0647), .B0(new_n12586_), .Y(new_n12587_));
  NOR2X1   g10151(.A(new_n12587_), .B(pi0630), .Y(new_n12588_));
  INVX1    g10152(.A(new_n12588_), .Y(new_n12589_));
  OAI21X1  g10153(.A0(new_n12581_), .A1(pi0647), .B0(pi1157), .Y(new_n12590_));
  AOI21X1  g10154(.A0(new_n12576_), .A1(pi0647), .B0(new_n12590_), .Y(new_n12591_));
  INVX1    g10155(.A(pi0630), .Y(new_n12592_));
  OAI21X1  g10156(.A0(new_n12469_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n12593_));
  AOI21X1  g10157(.A0(new_n12585_), .A1(new_n12577_), .B0(new_n12593_), .Y(new_n12594_));
  NOR2X1   g10158(.A(new_n12594_), .B(new_n12592_), .Y(new_n12595_));
  INVX1    g10159(.A(new_n12595_), .Y(new_n12596_));
  OAI22X1  g10160(.A0(new_n12596_), .A1(new_n12591_), .B0(new_n12589_), .B1(new_n12583_), .Y(new_n12597_));
  MX2X1    g10161(.A(new_n12597_), .B(new_n12576_), .S0(new_n11763_), .Y(new_n12598_));
  OAI21X1  g10162(.A0(new_n12594_), .A1(new_n12587_), .B0(pi0787), .Y(new_n12599_));
  OAI21X1  g10163(.A0(new_n12585_), .A1(pi0787), .B0(new_n12599_), .Y(new_n12600_));
  OAI21X1  g10164(.A0(new_n12600_), .A1(pi0644), .B0(pi0715), .Y(new_n12601_));
  AOI21X1  g10165(.A0(new_n12598_), .A1(pi0644), .B0(new_n12601_), .Y(new_n12602_));
  XOR2X1   g10166(.A(pi1157), .B(new_n12592_), .Y(new_n12603_));
  NOR2X1   g10167(.A(new_n12603_), .B(new_n11763_), .Y(new_n12604_));
  INVX1    g10168(.A(new_n12604_), .Y(new_n12605_));
  NOR2X1   g10169(.A(new_n12605_), .B(new_n12451_), .Y(new_n12606_));
  AOI21X1  g10170(.A0(new_n12605_), .A1(new_n12581_), .B0(new_n12606_), .Y(new_n12607_));
  INVX1    g10171(.A(pi0715), .Y(new_n12608_));
  OAI21X1  g10172(.A0(new_n12469_), .A1(pi0644), .B0(new_n12608_), .Y(new_n12609_));
  AOI21X1  g10173(.A0(new_n12607_), .A1(pi0644), .B0(new_n12609_), .Y(new_n12610_));
  NOR3X1   g10174(.A(new_n12610_), .B(new_n12602_), .C(new_n11762_), .Y(new_n12611_));
  INVX1    g10175(.A(pi0644), .Y(new_n12612_));
  OAI21X1  g10176(.A0(new_n12600_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n12613_));
  AOI21X1  g10177(.A0(new_n12598_), .A1(new_n12612_), .B0(new_n12613_), .Y(new_n12614_));
  OAI21X1  g10178(.A0(new_n12469_), .A1(new_n12612_), .B0(pi0715), .Y(new_n12615_));
  AOI21X1  g10179(.A0(new_n12607_), .A1(new_n12612_), .B0(new_n12615_), .Y(new_n12616_));
  OR2X1    g10180(.A(new_n12616_), .B(pi1160), .Y(new_n12617_));
  OAI21X1  g10181(.A0(new_n12617_), .A1(new_n12614_), .B0(pi0790), .Y(new_n12618_));
  OR2X1    g10182(.A(new_n12598_), .B(pi0790), .Y(new_n12619_));
  AND2X1   g10183(.A(new_n12619_), .B(new_n6489_), .Y(new_n12620_));
  OAI21X1  g10184(.A0(new_n12618_), .A1(new_n12611_), .B0(new_n12620_), .Y(new_n12621_));
  AOI21X1  g10185(.A0(po1038), .A1(new_n7353_), .B0(pi0832), .Y(new_n12622_));
  AOI21X1  g10186(.A0(pi1093), .A1(pi1092), .B0(pi0140), .Y(new_n12623_));
  AOI21X1  g10187(.A0(new_n12439_), .A1(new_n11771_), .B0(new_n12623_), .Y(new_n12624_));
  AND3X1   g10188(.A(new_n12439_), .B(new_n11771_), .C(new_n12363_), .Y(new_n12625_));
  NOR2X1   g10189(.A(new_n12625_), .B(new_n12624_), .Y(new_n12626_));
  OR2X1    g10190(.A(new_n12623_), .B(pi1153), .Y(new_n12627_));
  OAI22X1  g10191(.A0(new_n12627_), .A1(new_n12625_), .B0(new_n12626_), .B1(new_n12364_), .Y(new_n12628_));
  MX2X1    g10192(.A(new_n12628_), .B(new_n12624_), .S0(new_n11769_), .Y(new_n12629_));
  AND2X1   g10193(.A(new_n12490_), .B(new_n2720_), .Y(new_n12630_));
  AND2X1   g10194(.A(new_n12513_), .B(new_n2720_), .Y(new_n12631_));
  NOR3X1   g10195(.A(new_n12631_), .B(new_n12630_), .C(new_n12629_), .Y(new_n12632_));
  NOR3X1   g10196(.A(new_n12530_), .B(new_n2725_), .C(new_n11766_), .Y(new_n12633_));
  INVX1    g10197(.A(new_n12633_), .Y(new_n12634_));
  XOR2X1   g10198(.A(pi1158), .B(pi0626), .Y(new_n12635_));
  XOR2X1   g10199(.A(pi0641), .B(pi0626), .Y(new_n12636_));
  AND2X1   g10200(.A(new_n12636_), .B(new_n12635_), .Y(new_n12637_));
  AND3X1   g10201(.A(new_n12637_), .B(new_n12634_), .C(new_n12632_), .Y(new_n12638_));
  INVX1    g10202(.A(new_n12562_), .Y(new_n12639_));
  AOI21X1  g10203(.A0(new_n12056_), .A1(new_n11772_), .B0(new_n12623_), .Y(new_n12640_));
  AOI21X1  g10204(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n12640_), .Y(new_n12641_));
  NOR2X1   g10205(.A(new_n12471_), .B(new_n2725_), .Y(new_n12642_));
  OAI21X1  g10206(.A0(new_n12642_), .A1(new_n12640_), .B0(pi1155), .Y(new_n12643_));
  INVX1    g10207(.A(new_n12643_), .Y(new_n12644_));
  AND3X1   g10208(.A(pi1093), .B(pi1092), .C(pi0609), .Y(new_n12645_));
  INVX1    g10209(.A(new_n12645_), .Y(new_n12646_));
  AOI21X1  g10210(.A0(new_n12646_), .A1(new_n12641_), .B0(pi1155), .Y(new_n12647_));
  OAI21X1  g10211(.A0(new_n12647_), .A1(new_n12644_), .B0(pi0785), .Y(new_n12648_));
  OAI21X1  g10212(.A0(new_n12641_), .A1(pi0785), .B0(new_n12648_), .Y(new_n12649_));
  INVX1    g10213(.A(new_n12649_), .Y(new_n12650_));
  AND2X1   g10214(.A(new_n2720_), .B(new_n12486_), .Y(new_n12651_));
  INVX1    g10215(.A(new_n12651_), .Y(new_n12652_));
  AOI21X1  g10216(.A0(new_n12652_), .A1(new_n12650_), .B0(new_n12487_), .Y(new_n12653_));
  AND3X1   g10217(.A(pi1093), .B(pi1092), .C(pi0618), .Y(new_n12654_));
  INVX1    g10218(.A(new_n12654_), .Y(new_n12655_));
  AOI21X1  g10219(.A0(new_n12655_), .A1(new_n12650_), .B0(pi1154), .Y(new_n12656_));
  NOR2X1   g10220(.A(new_n12656_), .B(new_n12653_), .Y(new_n12657_));
  MX2X1    g10221(.A(new_n12657_), .B(new_n12650_), .S0(new_n11767_), .Y(new_n12658_));
  NOR2X1   g10222(.A(new_n12658_), .B(pi0789), .Y(new_n12659_));
  INVX1    g10223(.A(new_n12658_), .Y(new_n12660_));
  AOI21X1  g10224(.A0(new_n12623_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n12661_));
  OAI21X1  g10225(.A0(new_n12660_), .A1(new_n12509_), .B0(new_n12661_), .Y(new_n12662_));
  AOI21X1  g10226(.A0(new_n12623_), .A1(pi0619), .B0(pi1159), .Y(new_n12663_));
  OAI21X1  g10227(.A0(new_n12660_), .A1(pi0619), .B0(new_n12663_), .Y(new_n12664_));
  AOI21X1  g10228(.A0(new_n12664_), .A1(new_n12662_), .B0(new_n11766_), .Y(new_n12665_));
  NOR2X1   g10229(.A(new_n12665_), .B(new_n12659_), .Y(new_n12666_));
  INVX1    g10230(.A(new_n12666_), .Y(new_n12667_));
  AOI21X1  g10231(.A0(new_n12623_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n12668_));
  OAI21X1  g10232(.A0(new_n12667_), .A1(new_n12542_), .B0(new_n12668_), .Y(new_n12669_));
  AOI21X1  g10233(.A0(new_n12623_), .A1(pi0626), .B0(pi1158), .Y(new_n12670_));
  OAI21X1  g10234(.A0(new_n12667_), .A1(pi0626), .B0(new_n12670_), .Y(new_n12671_));
  AND3X1   g10235(.A(new_n12671_), .B(new_n12669_), .C(new_n12639_), .Y(new_n12672_));
  OAI21X1  g10236(.A0(new_n12672_), .A1(new_n12638_), .B0(pi0788), .Y(new_n12673_));
  OAI21X1  g10237(.A0(new_n12624_), .A1(new_n11991_), .B0(new_n12640_), .Y(new_n12674_));
  OR3X1    g10238(.A(new_n12624_), .B(new_n11991_), .C(new_n12363_), .Y(new_n12675_));
  AOI21X1  g10239(.A0(new_n12674_), .A1(new_n12675_), .B0(new_n12627_), .Y(new_n12676_));
  OAI21X1  g10240(.A0(new_n12626_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n12677_));
  AND3X1   g10241(.A(new_n12675_), .B(new_n12640_), .C(pi1153), .Y(new_n12678_));
  OAI21X1  g10242(.A0(new_n12627_), .A1(new_n12625_), .B0(pi0608), .Y(new_n12679_));
  OAI22X1  g10243(.A0(new_n12679_), .A1(new_n12678_), .B0(new_n12677_), .B1(new_n12676_), .Y(new_n12680_));
  MX2X1    g10244(.A(new_n12680_), .B(new_n12674_), .S0(new_n11769_), .Y(new_n12681_));
  OAI21X1  g10245(.A0(new_n12629_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n12682_));
  AOI21X1  g10246(.A0(new_n12681_), .A1(new_n12462_), .B0(new_n12682_), .Y(new_n12683_));
  NAND2X1  g10247(.A(new_n12643_), .B(new_n12468_), .Y(new_n12684_));
  OAI21X1  g10248(.A0(new_n12629_), .A1(pi0609), .B0(pi1155), .Y(new_n12685_));
  AOI21X1  g10249(.A0(new_n12681_), .A1(pi0609), .B0(new_n12685_), .Y(new_n12686_));
  OR2X1    g10250(.A(new_n12647_), .B(new_n12468_), .Y(new_n12687_));
  OAI22X1  g10251(.A0(new_n12687_), .A1(new_n12686_), .B0(new_n12684_), .B1(new_n12683_), .Y(new_n12688_));
  MX2X1    g10252(.A(new_n12688_), .B(new_n12681_), .S0(new_n11768_), .Y(new_n12689_));
  OR2X1    g10253(.A(new_n12630_), .B(new_n12629_), .Y(new_n12690_));
  OAI21X1  g10254(.A0(new_n12690_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n12691_));
  AOI21X1  g10255(.A0(new_n12689_), .A1(new_n12486_), .B0(new_n12691_), .Y(new_n12692_));
  OR2X1    g10256(.A(new_n12653_), .B(pi0627), .Y(new_n12693_));
  OAI21X1  g10257(.A0(new_n12690_), .A1(pi0618), .B0(pi1154), .Y(new_n12694_));
  AOI21X1  g10258(.A0(new_n12689_), .A1(pi0618), .B0(new_n12694_), .Y(new_n12695_));
  OR2X1    g10259(.A(new_n12656_), .B(new_n12494_), .Y(new_n12696_));
  OAI22X1  g10260(.A0(new_n12696_), .A1(new_n12695_), .B0(new_n12693_), .B1(new_n12692_), .Y(new_n12697_));
  MX2X1    g10261(.A(new_n12697_), .B(new_n12689_), .S0(new_n11767_), .Y(new_n12698_));
  NAND2X1  g10262(.A(new_n12698_), .B(new_n12509_), .Y(new_n12699_));
  AOI21X1  g10263(.A0(new_n12632_), .A1(pi0619), .B0(pi1159), .Y(new_n12700_));
  NAND2X1  g10264(.A(new_n12662_), .B(new_n12517_), .Y(new_n12701_));
  AOI21X1  g10265(.A0(new_n12700_), .A1(new_n12699_), .B0(new_n12701_), .Y(new_n12702_));
  NAND2X1  g10266(.A(new_n12698_), .B(pi0619), .Y(new_n12703_));
  AOI21X1  g10267(.A0(new_n12632_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n12704_));
  NAND2X1  g10268(.A(new_n12664_), .B(pi0648), .Y(new_n12705_));
  AOI21X1  g10269(.A0(new_n12704_), .A1(new_n12703_), .B0(new_n12705_), .Y(new_n12706_));
  NOR3X1   g10270(.A(new_n12706_), .B(new_n12702_), .C(new_n11766_), .Y(new_n12707_));
  AND2X1   g10271(.A(new_n12635_), .B(pi0788), .Y(new_n12708_));
  NOR2X1   g10272(.A(new_n12708_), .B(new_n12563_), .Y(new_n12709_));
  OAI21X1  g10273(.A0(new_n12698_), .A1(pi0789), .B0(new_n12709_), .Y(new_n12710_));
  OAI21X1  g10274(.A0(new_n12710_), .A1(new_n12707_), .B0(new_n12673_), .Y(new_n12711_));
  AND2X1   g10275(.A(new_n12671_), .B(new_n12669_), .Y(new_n12712_));
  MX2X1    g10276(.A(new_n12712_), .B(new_n12666_), .S0(new_n11765_), .Y(new_n12713_));
  INVX1    g10277(.A(new_n12713_), .Y(new_n12714_));
  OAI21X1  g10278(.A0(new_n12714_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n12715_));
  AOI21X1  g10279(.A0(new_n12711_), .A1(new_n12554_), .B0(new_n12715_), .Y(new_n12716_));
  NOR3X1   g10280(.A(new_n12562_), .B(new_n2725_), .C(new_n11765_), .Y(new_n12717_));
  INVX1    g10281(.A(new_n12717_), .Y(new_n12718_));
  AND3X1   g10282(.A(new_n12718_), .B(new_n12634_), .C(new_n12632_), .Y(new_n12719_));
  INVX1    g10283(.A(new_n12719_), .Y(new_n12720_));
  AOI21X1  g10284(.A0(new_n2720_), .A1(new_n12554_), .B0(new_n12720_), .Y(new_n12721_));
  OAI21X1  g10285(.A0(new_n12721_), .A1(new_n12555_), .B0(new_n12561_), .Y(new_n12722_));
  OAI21X1  g10286(.A0(new_n12714_), .A1(pi0628), .B0(pi1156), .Y(new_n12723_));
  AOI21X1  g10287(.A0(new_n12711_), .A1(pi0628), .B0(new_n12723_), .Y(new_n12724_));
  AOI21X1  g10288(.A0(new_n2720_), .A1(pi0628), .B0(new_n12720_), .Y(new_n12725_));
  OAI21X1  g10289(.A0(new_n12725_), .A1(pi1156), .B0(pi0629), .Y(new_n12726_));
  OAI22X1  g10290(.A0(new_n12726_), .A1(new_n12724_), .B0(new_n12722_), .B1(new_n12716_), .Y(new_n12727_));
  MX2X1    g10291(.A(new_n12727_), .B(new_n12711_), .S0(new_n11764_), .Y(new_n12728_));
  INVX1    g10292(.A(new_n12623_), .Y(new_n12729_));
  MX2X1    g10293(.A(new_n12714_), .B(new_n12729_), .S0(new_n12580_), .Y(new_n12730_));
  OAI21X1  g10294(.A0(new_n12730_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n12731_));
  AOI21X1  g10295(.A0(new_n12728_), .A1(new_n12577_), .B0(new_n12731_), .Y(new_n12732_));
  AND2X1   g10296(.A(pi1156), .B(new_n12554_), .Y(new_n12733_));
  INVX1    g10297(.A(new_n12733_), .Y(new_n12734_));
  AND2X1   g10298(.A(new_n12555_), .B(pi0628), .Y(new_n12735_));
  INVX1    g10299(.A(new_n12735_), .Y(new_n12736_));
  AOI21X1  g10300(.A0(new_n12736_), .A1(new_n12734_), .B0(new_n11764_), .Y(new_n12737_));
  AND2X1   g10301(.A(new_n12737_), .B(new_n2720_), .Y(new_n12738_));
  INVX1    g10302(.A(new_n12738_), .Y(new_n12739_));
  AND2X1   g10303(.A(new_n12739_), .B(new_n12719_), .Y(new_n12740_));
  OAI21X1  g10304(.A0(new_n12729_), .A1(pi0647), .B0(pi1157), .Y(new_n12741_));
  AOI21X1  g10305(.A0(new_n12740_), .A1(pi0647), .B0(new_n12741_), .Y(new_n12742_));
  OR2X1    g10306(.A(new_n12742_), .B(pi0630), .Y(new_n12743_));
  OAI21X1  g10307(.A0(new_n12730_), .A1(pi0647), .B0(pi1157), .Y(new_n12744_));
  AOI21X1  g10308(.A0(new_n12728_), .A1(pi0647), .B0(new_n12744_), .Y(new_n12745_));
  OAI21X1  g10309(.A0(new_n12729_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n12746_));
  AOI21X1  g10310(.A0(new_n12740_), .A1(new_n12577_), .B0(new_n12746_), .Y(new_n12747_));
  OR2X1    g10311(.A(new_n12747_), .B(new_n12592_), .Y(new_n12748_));
  OAI22X1  g10312(.A0(new_n12748_), .A1(new_n12745_), .B0(new_n12743_), .B1(new_n12732_), .Y(new_n12749_));
  MX2X1    g10313(.A(new_n12749_), .B(new_n12728_), .S0(new_n11763_), .Y(new_n12750_));
  OAI21X1  g10314(.A0(new_n12747_), .A1(new_n12742_), .B0(pi0787), .Y(new_n12751_));
  OAI21X1  g10315(.A0(new_n12740_), .A1(pi0787), .B0(new_n12751_), .Y(new_n12752_));
  OAI21X1  g10316(.A0(new_n12752_), .A1(pi0644), .B0(pi0715), .Y(new_n12753_));
  AOI21X1  g10317(.A0(new_n12750_), .A1(pi0644), .B0(new_n12753_), .Y(new_n12754_));
  NOR3X1   g10318(.A(new_n12623_), .B(new_n12603_), .C(new_n11763_), .Y(new_n12755_));
  AOI21X1  g10319(.A0(new_n12730_), .A1(new_n12605_), .B0(new_n12755_), .Y(new_n12756_));
  OAI21X1  g10320(.A0(new_n12729_), .A1(pi0644), .B0(new_n12608_), .Y(new_n12757_));
  AOI21X1  g10321(.A0(new_n12756_), .A1(pi0644), .B0(new_n12757_), .Y(new_n12758_));
  NOR3X1   g10322(.A(new_n12758_), .B(new_n12754_), .C(new_n11762_), .Y(new_n12759_));
  OAI21X1  g10323(.A0(new_n12752_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n12760_));
  AOI21X1  g10324(.A0(new_n12750_), .A1(new_n12612_), .B0(new_n12760_), .Y(new_n12761_));
  OAI21X1  g10325(.A0(new_n12729_), .A1(new_n12612_), .B0(pi0715), .Y(new_n12762_));
  AOI21X1  g10326(.A0(new_n12756_), .A1(new_n12612_), .B0(new_n12762_), .Y(new_n12763_));
  NOR3X1   g10327(.A(new_n12763_), .B(new_n12761_), .C(pi1160), .Y(new_n12764_));
  OAI21X1  g10328(.A0(new_n12764_), .A1(new_n12759_), .B0(pi0790), .Y(new_n12765_));
  INVX1    g10329(.A(pi0790), .Y(new_n12766_));
  INVX1    g10330(.A(pi0832), .Y(new_n12767_));
  AOI21X1  g10331(.A0(new_n12750_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n12768_));
  AOI22X1  g10332(.A0(new_n12768_), .A1(new_n12765_), .B0(new_n12622_), .B1(new_n12621_), .Y(po0297));
  NOR2X1   g10333(.A(new_n3103_), .B(new_n11676_), .Y(new_n12770_));
  INVX1    g10334(.A(new_n12077_), .Y(new_n12771_));
  AOI22X1  g10335(.A0(new_n12079_), .A1(pi0749), .B0(new_n12771_), .B1(new_n11676_), .Y(new_n12772_));
  OR2X1    g10336(.A(new_n12772_), .B(new_n2979_), .Y(new_n12773_));
  INVX1    g10337(.A(pi0749), .Y(new_n12774_));
  AOI22X1  g10338(.A0(new_n12073_), .A1(pi0141), .B0(new_n12444_), .B1(new_n12774_), .Y(new_n12775_));
  MX2X1    g10339(.A(new_n12034_), .B(new_n11975_), .S0(new_n2939_), .Y(new_n12776_));
  AOI21X1  g10340(.A0(new_n12046_), .A1(pi0141), .B0(new_n12774_), .Y(new_n12777_));
  OAI21X1  g10341(.A0(new_n12776_), .A1(pi0141), .B0(new_n12777_), .Y(new_n12778_));
  AND2X1   g10342(.A(new_n11821_), .B(new_n2939_), .Y(new_n12779_));
  OR3X1    g10343(.A(new_n12779_), .B(pi0749), .C(pi0141), .Y(new_n12780_));
  AOI21X1  g10344(.A0(new_n12780_), .A1(new_n12778_), .B0(pi0038), .Y(new_n12781_));
  OAI21X1  g10345(.A0(new_n12775_), .A1(new_n2939_), .B0(new_n12781_), .Y(new_n12782_));
  AND2X1   g10346(.A(new_n12782_), .B(new_n12773_), .Y(new_n12783_));
  OR2X1    g10347(.A(new_n12783_), .B(pi0706), .Y(new_n12784_));
  OAI21X1  g10348(.A0(new_n12213_), .A1(new_n11676_), .B0(new_n12774_), .Y(new_n12785_));
  AOI21X1  g10349(.A0(new_n12155_), .A1(new_n11676_), .B0(new_n12785_), .Y(new_n12786_));
  OAI22X1  g10350(.A0(new_n12258_), .A1(new_n2933_), .B0(new_n12249_), .B1(new_n12235_), .Y(new_n12787_));
  MX2X1    g10351(.A(new_n12300_), .B(new_n12290_), .S0(new_n2933_), .Y(new_n12788_));
  AOI21X1  g10352(.A0(new_n12788_), .A1(new_n11676_), .B0(new_n12774_), .Y(new_n12789_));
  OAI21X1  g10353(.A0(new_n12787_), .A1(new_n11676_), .B0(new_n12789_), .Y(new_n12790_));
  NAND2X1  g10354(.A(new_n12790_), .B(pi0039), .Y(new_n12791_));
  INVX1    g10355(.A(new_n12315_), .Y(new_n12792_));
  NOR4X1   g10356(.A(new_n12324_), .B(new_n12323_), .C(new_n12316_), .D(new_n5019_), .Y(new_n12793_));
  NOR3X1   g10357(.A(new_n12330_), .B(new_n12328_), .C(new_n5019_), .Y(new_n12794_));
  MX2X1    g10358(.A(new_n12794_), .B(new_n12793_), .S0(new_n2933_), .Y(new_n12795_));
  AOI21X1  g10359(.A0(new_n12795_), .A1(pi0141), .B0(pi0749), .Y(new_n12796_));
  OAI21X1  g10360(.A0(new_n12792_), .A1(pi0141), .B0(new_n12796_), .Y(new_n12797_));
  NOR3X1   g10361(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .Y(new_n12798_));
  OR2X1    g10362(.A(new_n12798_), .B(pi0141), .Y(new_n12799_));
  OR2X1    g10363(.A(new_n12344_), .B(new_n12045_), .Y(new_n12800_));
  AOI21X1  g10364(.A0(new_n12800_), .A1(pi0141), .B0(new_n12774_), .Y(new_n12801_));
  AOI21X1  g10365(.A0(new_n12801_), .A1(new_n12799_), .B0(pi0039), .Y(new_n12802_));
  AOI21X1  g10366(.A0(new_n12802_), .A1(new_n12797_), .B0(pi0038), .Y(new_n12803_));
  OAI21X1  g10367(.A0(new_n12791_), .A1(new_n12786_), .B0(new_n12803_), .Y(new_n12804_));
  INVX1    g10368(.A(pi0706), .Y(new_n12805_));
  AOI21X1  g10369(.A0(new_n12353_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n12806_));
  AOI21X1  g10370(.A0(new_n12806_), .A1(new_n12772_), .B0(new_n12805_), .Y(new_n12807_));
  AOI21X1  g10371(.A0(new_n12807_), .A1(new_n12804_), .B0(new_n11770_), .Y(new_n12808_));
  AOI21X1  g10372(.A0(new_n12808_), .A1(new_n12784_), .B0(new_n12770_), .Y(new_n12809_));
  MX2X1    g10373(.A(new_n12783_), .B(pi0141), .S0(new_n11770_), .Y(new_n12810_));
  OAI21X1  g10374(.A0(new_n12810_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n12811_));
  AOI21X1  g10375(.A0(new_n12809_), .A1(new_n12363_), .B0(new_n12811_), .Y(new_n12812_));
  NAND2X1  g10376(.A(new_n11904_), .B(new_n5019_), .Y(new_n12813_));
  AOI21X1  g10377(.A0(new_n11904_), .A1(new_n5019_), .B0(new_n12398_), .Y(new_n12814_));
  AOI22X1  g10378(.A0(new_n12402_), .A1(new_n12813_), .B0(new_n12814_), .B1(new_n11867_), .Y(new_n12815_));
  AOI21X1  g10379(.A0(new_n12815_), .A1(new_n5041_), .B0(new_n12409_), .Y(new_n12816_));
  INVX1    g10380(.A(new_n12412_), .Y(new_n12817_));
  INVX1    g10381(.A(new_n12420_), .Y(new_n12818_));
  OAI22X1  g10382(.A0(new_n12818_), .A1(new_n12415_), .B0(new_n12817_), .B1(new_n12816_), .Y(new_n12819_));
  AOI21X1  g10383(.A0(new_n12815_), .A1(new_n5058_), .B0(new_n12422_), .Y(new_n12820_));
  INVX1    g10384(.A(new_n12427_), .Y(new_n12821_));
  INVX1    g10385(.A(new_n12430_), .Y(new_n12822_));
  OAI22X1  g10386(.A0(new_n12822_), .A1(new_n12428_), .B0(new_n12821_), .B1(new_n12820_), .Y(new_n12823_));
  MX2X1    g10387(.A(new_n12823_), .B(new_n12819_), .S0(new_n2933_), .Y(new_n12824_));
  MX2X1    g10388(.A(new_n12824_), .B(new_n12340_), .S0(new_n2939_), .Y(new_n12825_));
  MX2X1    g10389(.A(new_n12394_), .B(new_n12435_), .S0(new_n2939_), .Y(new_n12826_));
  OAI21X1  g10390(.A0(new_n12826_), .A1(new_n11676_), .B0(new_n2979_), .Y(new_n12827_));
  AOI21X1  g10391(.A0(new_n12825_), .A1(new_n11676_), .B0(new_n12827_), .Y(new_n12828_));
  AOI21X1  g10392(.A0(new_n12771_), .A1(new_n11676_), .B0(new_n12441_), .Y(new_n12829_));
  OR3X1    g10393(.A(new_n12829_), .B(new_n12828_), .C(new_n12805_), .Y(new_n12830_));
  INVX1    g10394(.A(new_n12446_), .Y(new_n12831_));
  MX2X1    g10395(.A(new_n12831_), .B(new_n11959_), .S0(new_n2979_), .Y(new_n12832_));
  NOR2X1   g10396(.A(pi0706), .B(pi0141), .Y(new_n12833_));
  AOI21X1  g10397(.A0(new_n12833_), .A1(new_n12832_), .B0(new_n11770_), .Y(new_n12834_));
  AOI21X1  g10398(.A0(new_n12834_), .A1(new_n12830_), .B0(new_n12770_), .Y(new_n12835_));
  OAI21X1  g10399(.A0(new_n12832_), .A1(new_n11770_), .B0(new_n11676_), .Y(new_n12836_));
  OAI21X1  g10400(.A0(new_n12836_), .A1(pi0625), .B0(pi1153), .Y(new_n12837_));
  AOI21X1  g10401(.A0(new_n12835_), .A1(pi0625), .B0(new_n12837_), .Y(new_n12838_));
  OR3X1    g10402(.A(new_n12838_), .B(new_n12812_), .C(pi0608), .Y(new_n12839_));
  OAI21X1  g10403(.A0(new_n12810_), .A1(pi0625), .B0(pi1153), .Y(new_n12840_));
  AOI21X1  g10404(.A0(new_n12809_), .A1(pi0625), .B0(new_n12840_), .Y(new_n12841_));
  OAI21X1  g10405(.A0(new_n12836_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n12842_));
  AOI21X1  g10406(.A0(new_n12835_), .A1(new_n12363_), .B0(new_n12842_), .Y(new_n12843_));
  OR3X1    g10407(.A(new_n12843_), .B(new_n12841_), .C(new_n12368_), .Y(new_n12844_));
  AOI21X1  g10408(.A0(new_n12844_), .A1(new_n12839_), .B0(new_n11769_), .Y(new_n12845_));
  AOI21X1  g10409(.A0(new_n12809_), .A1(new_n11769_), .B0(new_n12845_), .Y(new_n12846_));
  NOR2X1   g10410(.A(new_n12843_), .B(new_n12838_), .Y(new_n12847_));
  MX2X1    g10411(.A(new_n12847_), .B(new_n12835_), .S0(new_n11769_), .Y(new_n12848_));
  AOI21X1  g10412(.A0(new_n12848_), .A1(pi0609), .B0(pi1155), .Y(new_n12849_));
  OAI21X1  g10413(.A0(new_n12846_), .A1(pi0609), .B0(new_n12849_), .Y(new_n12850_));
  AND2X1   g10414(.A(new_n12810_), .B(new_n12474_), .Y(new_n12851_));
  AOI22X1  g10415(.A0(new_n12851_), .A1(pi0609), .B0(new_n12836_), .B1(new_n12472_), .Y(new_n12852_));
  OR2X1    g10416(.A(new_n12852_), .B(new_n12463_), .Y(new_n12853_));
  AND2X1   g10417(.A(new_n12853_), .B(new_n12468_), .Y(new_n12854_));
  AOI21X1  g10418(.A0(new_n12848_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n12855_));
  OAI21X1  g10419(.A0(new_n12846_), .A1(new_n12462_), .B0(new_n12855_), .Y(new_n12856_));
  AOI22X1  g10420(.A0(new_n12851_), .A1(new_n12462_), .B0(new_n12836_), .B1(new_n12481_), .Y(new_n12857_));
  OR2X1    g10421(.A(new_n12857_), .B(pi1155), .Y(new_n12858_));
  AND2X1   g10422(.A(new_n12858_), .B(pi0660), .Y(new_n12859_));
  AOI22X1  g10423(.A0(new_n12859_), .A1(new_n12856_), .B0(new_n12854_), .B1(new_n12850_), .Y(new_n12860_));
  OR2X1    g10424(.A(new_n12846_), .B(pi0785), .Y(new_n12861_));
  OAI21X1  g10425(.A0(new_n12860_), .A1(new_n11768_), .B0(new_n12861_), .Y(new_n12862_));
  NAND2X1  g10426(.A(new_n12836_), .B(new_n12490_), .Y(new_n12863_));
  OAI21X1  g10427(.A0(new_n12848_), .A1(new_n12490_), .B0(new_n12863_), .Y(new_n12864_));
  OAI21X1  g10428(.A0(new_n12864_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n12865_));
  AOI21X1  g10429(.A0(new_n12862_), .A1(new_n12486_), .B0(new_n12865_), .Y(new_n12866_));
  MX2X1    g10430(.A(new_n12836_), .B(new_n12810_), .S0(new_n12474_), .Y(new_n12867_));
  NAND2X1  g10431(.A(new_n12858_), .B(new_n12853_), .Y(new_n12868_));
  MX2X1    g10432(.A(new_n12868_), .B(new_n12867_), .S0(new_n11768_), .Y(new_n12869_));
  INVX1    g10433(.A(new_n12836_), .Y(new_n12870_));
  AOI21X1  g10434(.A0(new_n12870_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n12871_));
  OAI21X1  g10435(.A0(new_n12869_), .A1(new_n12486_), .B0(new_n12871_), .Y(new_n12872_));
  NAND2X1  g10436(.A(new_n12872_), .B(new_n12494_), .Y(new_n12873_));
  OAI21X1  g10437(.A0(new_n12864_), .A1(pi0618), .B0(pi1154), .Y(new_n12874_));
  AOI21X1  g10438(.A0(new_n12862_), .A1(pi0618), .B0(new_n12874_), .Y(new_n12875_));
  AOI21X1  g10439(.A0(new_n12870_), .A1(pi0618), .B0(pi1154), .Y(new_n12876_));
  OAI21X1  g10440(.A0(new_n12869_), .A1(pi0618), .B0(new_n12876_), .Y(new_n12877_));
  NAND2X1  g10441(.A(new_n12877_), .B(pi0627), .Y(new_n12878_));
  OAI22X1  g10442(.A0(new_n12878_), .A1(new_n12875_), .B0(new_n12873_), .B1(new_n12866_), .Y(new_n12879_));
  MX2X1    g10443(.A(new_n12879_), .B(new_n12862_), .S0(new_n11767_), .Y(new_n12880_));
  MX2X1    g10444(.A(new_n12864_), .B(new_n12836_), .S0(new_n12513_), .Y(new_n12881_));
  OAI21X1  g10445(.A0(new_n12881_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n12882_));
  AOI21X1  g10446(.A0(new_n12880_), .A1(new_n12509_), .B0(new_n12882_), .Y(new_n12883_));
  NAND2X1  g10447(.A(new_n12877_), .B(new_n12872_), .Y(new_n12884_));
  MX2X1    g10448(.A(new_n12884_), .B(new_n12869_), .S0(new_n11767_), .Y(new_n12885_));
  AOI21X1  g10449(.A0(new_n12870_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n12886_));
  OAI21X1  g10450(.A0(new_n12885_), .A1(new_n12509_), .B0(new_n12886_), .Y(new_n12887_));
  NAND2X1  g10451(.A(new_n12887_), .B(new_n12517_), .Y(new_n12888_));
  OAI21X1  g10452(.A0(new_n12881_), .A1(pi0619), .B0(pi1159), .Y(new_n12889_));
  AOI21X1  g10453(.A0(new_n12880_), .A1(pi0619), .B0(new_n12889_), .Y(new_n12890_));
  AOI21X1  g10454(.A0(new_n12870_), .A1(pi0619), .B0(pi1159), .Y(new_n12891_));
  OAI21X1  g10455(.A0(new_n12885_), .A1(pi0619), .B0(new_n12891_), .Y(new_n12892_));
  NAND2X1  g10456(.A(new_n12892_), .B(pi0648), .Y(new_n12893_));
  OAI22X1  g10457(.A0(new_n12893_), .A1(new_n12890_), .B0(new_n12888_), .B1(new_n12883_), .Y(new_n12894_));
  MX2X1    g10458(.A(new_n12894_), .B(new_n12880_), .S0(new_n11766_), .Y(new_n12895_));
  MX2X1    g10459(.A(new_n12881_), .B(new_n12836_), .S0(new_n12531_), .Y(new_n12896_));
  AOI21X1  g10460(.A0(new_n12896_), .A1(pi0626), .B0(pi0641), .Y(new_n12897_));
  OAI21X1  g10461(.A0(new_n12895_), .A1(pi0626), .B0(new_n12897_), .Y(new_n12898_));
  AND2X1   g10462(.A(new_n12885_), .B(new_n11766_), .Y(new_n12899_));
  AOI21X1  g10463(.A0(new_n12892_), .A1(new_n12887_), .B0(new_n11766_), .Y(new_n12900_));
  NOR2X1   g10464(.A(new_n12900_), .B(new_n12899_), .Y(new_n12901_));
  OAI21X1  g10465(.A0(new_n12836_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n12902_));
  AOI21X1  g10466(.A0(new_n12901_), .A1(new_n12542_), .B0(new_n12902_), .Y(new_n12903_));
  OR2X1    g10467(.A(new_n12903_), .B(new_n12535_), .Y(new_n12904_));
  AOI21X1  g10468(.A0(new_n12896_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n12905_));
  OAI21X1  g10469(.A0(new_n12895_), .A1(new_n12542_), .B0(new_n12905_), .Y(new_n12906_));
  OAI21X1  g10470(.A0(new_n12836_), .A1(pi0626), .B0(pi1158), .Y(new_n12907_));
  AOI21X1  g10471(.A0(new_n12901_), .A1(pi0626), .B0(new_n12907_), .Y(new_n12908_));
  OR2X1    g10472(.A(new_n12908_), .B(new_n12546_), .Y(new_n12909_));
  AOI22X1  g10473(.A0(new_n12909_), .A1(new_n12906_), .B0(new_n12904_), .B1(new_n12898_), .Y(new_n12910_));
  MX2X1    g10474(.A(new_n12910_), .B(new_n12895_), .S0(new_n11765_), .Y(new_n12911_));
  OAI21X1  g10475(.A0(new_n12908_), .A1(new_n12903_), .B0(pi0788), .Y(new_n12912_));
  OAI21X1  g10476(.A0(new_n12901_), .A1(pi0788), .B0(new_n12912_), .Y(new_n12913_));
  OAI21X1  g10477(.A0(new_n12913_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n12914_));
  AOI21X1  g10478(.A0(new_n12911_), .A1(new_n12554_), .B0(new_n12914_), .Y(new_n12915_));
  MX2X1    g10479(.A(new_n12896_), .B(new_n12836_), .S0(new_n12563_), .Y(new_n12916_));
  AOI21X1  g10480(.A0(new_n12870_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n12917_));
  OAI21X1  g10481(.A0(new_n12916_), .A1(new_n12554_), .B0(new_n12917_), .Y(new_n12918_));
  NAND2X1  g10482(.A(new_n12918_), .B(new_n12561_), .Y(new_n12919_));
  OAI21X1  g10483(.A0(new_n12913_), .A1(pi0628), .B0(pi1156), .Y(new_n12920_));
  AOI21X1  g10484(.A0(new_n12911_), .A1(pi0628), .B0(new_n12920_), .Y(new_n12921_));
  AOI21X1  g10485(.A0(new_n12870_), .A1(pi0628), .B0(pi1156), .Y(new_n12922_));
  OAI21X1  g10486(.A0(new_n12916_), .A1(pi0628), .B0(new_n12922_), .Y(new_n12923_));
  NAND2X1  g10487(.A(new_n12923_), .B(pi0629), .Y(new_n12924_));
  OAI22X1  g10488(.A0(new_n12924_), .A1(new_n12921_), .B0(new_n12919_), .B1(new_n12915_), .Y(new_n12925_));
  MX2X1    g10489(.A(new_n12925_), .B(new_n12911_), .S0(new_n11764_), .Y(new_n12926_));
  MX2X1    g10490(.A(new_n12913_), .B(new_n12836_), .S0(new_n12580_), .Y(new_n12927_));
  OAI21X1  g10491(.A0(new_n12927_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n12928_));
  AOI21X1  g10492(.A0(new_n12926_), .A1(new_n12577_), .B0(new_n12928_), .Y(new_n12929_));
  INVX1    g10493(.A(new_n12916_), .Y(new_n12930_));
  AND2X1   g10494(.A(new_n12923_), .B(new_n12918_), .Y(new_n12931_));
  MX2X1    g10495(.A(new_n12931_), .B(new_n12930_), .S0(new_n11764_), .Y(new_n12932_));
  INVX1    g10496(.A(new_n12932_), .Y(new_n12933_));
  AOI21X1  g10497(.A0(new_n12870_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n12934_));
  OAI21X1  g10498(.A0(new_n12933_), .A1(new_n12577_), .B0(new_n12934_), .Y(new_n12935_));
  AND2X1   g10499(.A(new_n12935_), .B(new_n12592_), .Y(new_n12936_));
  INVX1    g10500(.A(new_n12936_), .Y(new_n12937_));
  OAI21X1  g10501(.A0(new_n12927_), .A1(pi0647), .B0(pi1157), .Y(new_n12938_));
  AOI21X1  g10502(.A0(new_n12926_), .A1(pi0647), .B0(new_n12938_), .Y(new_n12939_));
  AOI21X1  g10503(.A0(new_n12870_), .A1(pi0647), .B0(pi1157), .Y(new_n12940_));
  OAI21X1  g10504(.A0(new_n12933_), .A1(pi0647), .B0(new_n12940_), .Y(new_n12941_));
  AND2X1   g10505(.A(new_n12941_), .B(pi0630), .Y(new_n12942_));
  INVX1    g10506(.A(new_n12942_), .Y(new_n12943_));
  OAI22X1  g10507(.A0(new_n12943_), .A1(new_n12939_), .B0(new_n12937_), .B1(new_n12929_), .Y(new_n12944_));
  MX2X1    g10508(.A(new_n12944_), .B(new_n12926_), .S0(new_n11763_), .Y(new_n12945_));
  NAND2X1  g10509(.A(new_n12945_), .B(pi0644), .Y(new_n12946_));
  AND2X1   g10510(.A(new_n12941_), .B(new_n12935_), .Y(new_n12947_));
  MX2X1    g10511(.A(new_n12947_), .B(new_n12932_), .S0(new_n11763_), .Y(new_n12948_));
  AOI21X1  g10512(.A0(new_n12948_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n12949_));
  AND2X1   g10513(.A(new_n12836_), .B(new_n12604_), .Y(new_n12950_));
  AOI21X1  g10514(.A0(new_n12927_), .A1(new_n12605_), .B0(new_n12950_), .Y(new_n12951_));
  OAI21X1  g10515(.A0(new_n12836_), .A1(pi0644), .B0(new_n12608_), .Y(new_n12952_));
  AOI21X1  g10516(.A0(new_n12951_), .A1(pi0644), .B0(new_n12952_), .Y(new_n12953_));
  OR2X1    g10517(.A(new_n12953_), .B(new_n11762_), .Y(new_n12954_));
  AOI21X1  g10518(.A0(new_n12949_), .A1(new_n12946_), .B0(new_n12954_), .Y(new_n12955_));
  AND2X1   g10519(.A(new_n12948_), .B(pi0644), .Y(new_n12956_));
  OR2X1    g10520(.A(new_n12956_), .B(pi0715), .Y(new_n12957_));
  AOI21X1  g10521(.A0(new_n12945_), .A1(new_n12612_), .B0(new_n12957_), .Y(new_n12958_));
  OAI21X1  g10522(.A0(new_n12836_), .A1(new_n12612_), .B0(pi0715), .Y(new_n12959_));
  AOI21X1  g10523(.A0(new_n12951_), .A1(new_n12612_), .B0(new_n12959_), .Y(new_n12960_));
  OR2X1    g10524(.A(new_n12960_), .B(pi1160), .Y(new_n12961_));
  OAI21X1  g10525(.A0(new_n12961_), .A1(new_n12958_), .B0(pi0790), .Y(new_n12962_));
  OR2X1    g10526(.A(new_n12945_), .B(pi0790), .Y(new_n12963_));
  AND2X1   g10527(.A(new_n12963_), .B(new_n6489_), .Y(new_n12964_));
  OAI21X1  g10528(.A0(new_n12962_), .A1(new_n12955_), .B0(new_n12964_), .Y(new_n12965_));
  AOI21X1  g10529(.A0(po1038), .A1(new_n11676_), .B0(pi0832), .Y(new_n12966_));
  AOI21X1  g10530(.A0(pi1093), .A1(pi1092), .B0(pi0141), .Y(new_n12967_));
  AOI21X1  g10531(.A0(new_n12439_), .A1(pi0706), .B0(new_n12967_), .Y(new_n12968_));
  AND3X1   g10532(.A(new_n12439_), .B(pi0706), .C(new_n12363_), .Y(new_n12969_));
  NOR2X1   g10533(.A(new_n12969_), .B(new_n12968_), .Y(new_n12970_));
  OR2X1    g10534(.A(new_n12967_), .B(pi1153), .Y(new_n12971_));
  OAI22X1  g10535(.A0(new_n12971_), .A1(new_n12969_), .B0(new_n12970_), .B1(new_n12364_), .Y(new_n12972_));
  MX2X1    g10536(.A(new_n12972_), .B(new_n12968_), .S0(new_n11769_), .Y(new_n12973_));
  NOR3X1   g10537(.A(new_n12973_), .B(new_n12631_), .C(new_n12630_), .Y(new_n12974_));
  AND3X1   g10538(.A(new_n12974_), .B(new_n12637_), .C(new_n12634_), .Y(new_n12975_));
  AOI21X1  g10539(.A0(new_n12056_), .A1(pi0749), .B0(new_n12967_), .Y(new_n12976_));
  AOI21X1  g10540(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n12976_), .Y(new_n12977_));
  OAI21X1  g10541(.A0(new_n12976_), .A1(new_n12642_), .B0(pi1155), .Y(new_n12978_));
  INVX1    g10542(.A(new_n12978_), .Y(new_n12979_));
  AOI21X1  g10543(.A0(new_n12977_), .A1(new_n12646_), .B0(pi1155), .Y(new_n12980_));
  OAI21X1  g10544(.A0(new_n12980_), .A1(new_n12979_), .B0(pi0785), .Y(new_n12981_));
  OAI21X1  g10545(.A0(new_n12977_), .A1(pi0785), .B0(new_n12981_), .Y(new_n12982_));
  INVX1    g10546(.A(new_n12982_), .Y(new_n12983_));
  AOI21X1  g10547(.A0(new_n12983_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n12984_));
  AOI21X1  g10548(.A0(new_n12983_), .A1(new_n12655_), .B0(pi1154), .Y(new_n12985_));
  NOR2X1   g10549(.A(new_n12985_), .B(new_n12984_), .Y(new_n12986_));
  MX2X1    g10550(.A(new_n12986_), .B(new_n12983_), .S0(new_n11767_), .Y(new_n12987_));
  NOR2X1   g10551(.A(new_n12987_), .B(pi0789), .Y(new_n12988_));
  INVX1    g10552(.A(new_n12987_), .Y(new_n12989_));
  AOI21X1  g10553(.A0(new_n12967_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n12990_));
  OAI21X1  g10554(.A0(new_n12989_), .A1(new_n12509_), .B0(new_n12990_), .Y(new_n12991_));
  AOI21X1  g10555(.A0(new_n12967_), .A1(pi0619), .B0(pi1159), .Y(new_n12992_));
  OAI21X1  g10556(.A0(new_n12989_), .A1(pi0619), .B0(new_n12992_), .Y(new_n12993_));
  AOI21X1  g10557(.A0(new_n12993_), .A1(new_n12991_), .B0(new_n11766_), .Y(new_n12994_));
  NOR2X1   g10558(.A(new_n12994_), .B(new_n12988_), .Y(new_n12995_));
  INVX1    g10559(.A(new_n12995_), .Y(new_n12996_));
  AOI21X1  g10560(.A0(new_n12967_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n12997_));
  OAI21X1  g10561(.A0(new_n12996_), .A1(new_n12542_), .B0(new_n12997_), .Y(new_n12998_));
  AOI21X1  g10562(.A0(new_n12967_), .A1(pi0626), .B0(pi1158), .Y(new_n12999_));
  OAI21X1  g10563(.A0(new_n12996_), .A1(pi0626), .B0(new_n12999_), .Y(new_n13000_));
  AND3X1   g10564(.A(new_n13000_), .B(new_n12998_), .C(new_n12639_), .Y(new_n13001_));
  OAI21X1  g10565(.A0(new_n13001_), .A1(new_n12975_), .B0(pi0788), .Y(new_n13002_));
  OAI21X1  g10566(.A0(new_n12968_), .A1(new_n11991_), .B0(new_n12976_), .Y(new_n13003_));
  OR3X1    g10567(.A(new_n12968_), .B(new_n11991_), .C(new_n12363_), .Y(new_n13004_));
  AOI21X1  g10568(.A0(new_n13003_), .A1(new_n13004_), .B0(new_n12971_), .Y(new_n13005_));
  OAI21X1  g10569(.A0(new_n12970_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n13006_));
  AND3X1   g10570(.A(new_n13004_), .B(new_n12976_), .C(pi1153), .Y(new_n13007_));
  OAI21X1  g10571(.A0(new_n12971_), .A1(new_n12969_), .B0(pi0608), .Y(new_n13008_));
  OAI22X1  g10572(.A0(new_n13008_), .A1(new_n13007_), .B0(new_n13006_), .B1(new_n13005_), .Y(new_n13009_));
  MX2X1    g10573(.A(new_n13009_), .B(new_n13003_), .S0(new_n11769_), .Y(new_n13010_));
  OAI21X1  g10574(.A0(new_n12973_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n13011_));
  AOI21X1  g10575(.A0(new_n13010_), .A1(new_n12462_), .B0(new_n13011_), .Y(new_n13012_));
  NAND2X1  g10576(.A(new_n12978_), .B(new_n12468_), .Y(new_n13013_));
  OAI21X1  g10577(.A0(new_n12973_), .A1(pi0609), .B0(pi1155), .Y(new_n13014_));
  AOI21X1  g10578(.A0(new_n13010_), .A1(pi0609), .B0(new_n13014_), .Y(new_n13015_));
  OR2X1    g10579(.A(new_n12980_), .B(new_n12468_), .Y(new_n13016_));
  OAI22X1  g10580(.A0(new_n13016_), .A1(new_n13015_), .B0(new_n13013_), .B1(new_n13012_), .Y(new_n13017_));
  MX2X1    g10581(.A(new_n13017_), .B(new_n13010_), .S0(new_n11768_), .Y(new_n13018_));
  OR2X1    g10582(.A(new_n12973_), .B(new_n12630_), .Y(new_n13019_));
  OAI21X1  g10583(.A0(new_n13019_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13020_));
  AOI21X1  g10584(.A0(new_n13018_), .A1(new_n12486_), .B0(new_n13020_), .Y(new_n13021_));
  OR2X1    g10585(.A(new_n12984_), .B(pi0627), .Y(new_n13022_));
  OAI21X1  g10586(.A0(new_n13019_), .A1(pi0618), .B0(pi1154), .Y(new_n13023_));
  AOI21X1  g10587(.A0(new_n13018_), .A1(pi0618), .B0(new_n13023_), .Y(new_n13024_));
  OR2X1    g10588(.A(new_n12985_), .B(new_n12494_), .Y(new_n13025_));
  OAI22X1  g10589(.A0(new_n13025_), .A1(new_n13024_), .B0(new_n13022_), .B1(new_n13021_), .Y(new_n13026_));
  MX2X1    g10590(.A(new_n13026_), .B(new_n13018_), .S0(new_n11767_), .Y(new_n13027_));
  NAND2X1  g10591(.A(new_n13027_), .B(new_n12509_), .Y(new_n13028_));
  AOI21X1  g10592(.A0(new_n12974_), .A1(pi0619), .B0(pi1159), .Y(new_n13029_));
  NAND2X1  g10593(.A(new_n12991_), .B(new_n12517_), .Y(new_n13030_));
  AOI21X1  g10594(.A0(new_n13029_), .A1(new_n13028_), .B0(new_n13030_), .Y(new_n13031_));
  NAND2X1  g10595(.A(new_n13027_), .B(pi0619), .Y(new_n13032_));
  AOI21X1  g10596(.A0(new_n12974_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13033_));
  NAND2X1  g10597(.A(new_n12993_), .B(pi0648), .Y(new_n13034_));
  AOI21X1  g10598(.A0(new_n13033_), .A1(new_n13032_), .B0(new_n13034_), .Y(new_n13035_));
  NOR3X1   g10599(.A(new_n13035_), .B(new_n13031_), .C(new_n11766_), .Y(new_n13036_));
  OAI21X1  g10600(.A0(new_n13027_), .A1(pi0789), .B0(new_n12709_), .Y(new_n13037_));
  OAI21X1  g10601(.A0(new_n13037_), .A1(new_n13036_), .B0(new_n13002_), .Y(new_n13038_));
  AND2X1   g10602(.A(new_n13000_), .B(new_n12998_), .Y(new_n13039_));
  MX2X1    g10603(.A(new_n13039_), .B(new_n12995_), .S0(new_n11765_), .Y(new_n13040_));
  INVX1    g10604(.A(new_n13040_), .Y(new_n13041_));
  OAI21X1  g10605(.A0(new_n13041_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13042_));
  AOI21X1  g10606(.A0(new_n13038_), .A1(new_n12554_), .B0(new_n13042_), .Y(new_n13043_));
  AND3X1   g10607(.A(new_n12974_), .B(new_n12718_), .C(new_n12634_), .Y(new_n13044_));
  INVX1    g10608(.A(new_n13044_), .Y(new_n13045_));
  AOI21X1  g10609(.A0(new_n2720_), .A1(new_n12554_), .B0(new_n13045_), .Y(new_n13046_));
  OAI21X1  g10610(.A0(new_n13046_), .A1(new_n12555_), .B0(new_n12561_), .Y(new_n13047_));
  OAI21X1  g10611(.A0(new_n13041_), .A1(pi0628), .B0(pi1156), .Y(new_n13048_));
  AOI21X1  g10612(.A0(new_n13038_), .A1(pi0628), .B0(new_n13048_), .Y(new_n13049_));
  AOI21X1  g10613(.A0(new_n2720_), .A1(pi0628), .B0(new_n13045_), .Y(new_n13050_));
  OAI21X1  g10614(.A0(new_n13050_), .A1(pi1156), .B0(pi0629), .Y(new_n13051_));
  OAI22X1  g10615(.A0(new_n13051_), .A1(new_n13049_), .B0(new_n13047_), .B1(new_n13043_), .Y(new_n13052_));
  MX2X1    g10616(.A(new_n13052_), .B(new_n13038_), .S0(new_n11764_), .Y(new_n13053_));
  INVX1    g10617(.A(new_n12967_), .Y(new_n13054_));
  MX2X1    g10618(.A(new_n13041_), .B(new_n13054_), .S0(new_n12580_), .Y(new_n13055_));
  OAI21X1  g10619(.A0(new_n13055_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13056_));
  AOI21X1  g10620(.A0(new_n13053_), .A1(new_n12577_), .B0(new_n13056_), .Y(new_n13057_));
  AND2X1   g10621(.A(new_n13044_), .B(new_n12739_), .Y(new_n13058_));
  OAI21X1  g10622(.A0(new_n13054_), .A1(pi0647), .B0(pi1157), .Y(new_n13059_));
  AOI21X1  g10623(.A0(new_n13058_), .A1(pi0647), .B0(new_n13059_), .Y(new_n13060_));
  OR2X1    g10624(.A(new_n13060_), .B(pi0630), .Y(new_n13061_));
  OAI21X1  g10625(.A0(new_n13055_), .A1(pi0647), .B0(pi1157), .Y(new_n13062_));
  AOI21X1  g10626(.A0(new_n13053_), .A1(pi0647), .B0(new_n13062_), .Y(new_n13063_));
  OAI21X1  g10627(.A0(new_n13054_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13064_));
  AOI21X1  g10628(.A0(new_n13058_), .A1(new_n12577_), .B0(new_n13064_), .Y(new_n13065_));
  OR2X1    g10629(.A(new_n13065_), .B(new_n12592_), .Y(new_n13066_));
  OAI22X1  g10630(.A0(new_n13066_), .A1(new_n13063_), .B0(new_n13061_), .B1(new_n13057_), .Y(new_n13067_));
  MX2X1    g10631(.A(new_n13067_), .B(new_n13053_), .S0(new_n11763_), .Y(new_n13068_));
  OAI21X1  g10632(.A0(new_n13065_), .A1(new_n13060_), .B0(pi0787), .Y(new_n13069_));
  OAI21X1  g10633(.A0(new_n13058_), .A1(pi0787), .B0(new_n13069_), .Y(new_n13070_));
  OAI21X1  g10634(.A0(new_n13070_), .A1(pi0644), .B0(pi0715), .Y(new_n13071_));
  AOI21X1  g10635(.A0(new_n13068_), .A1(pi0644), .B0(new_n13071_), .Y(new_n13072_));
  NOR3X1   g10636(.A(new_n12967_), .B(new_n12603_), .C(new_n11763_), .Y(new_n13073_));
  AOI21X1  g10637(.A0(new_n13055_), .A1(new_n12605_), .B0(new_n13073_), .Y(new_n13074_));
  OAI21X1  g10638(.A0(new_n13054_), .A1(pi0644), .B0(new_n12608_), .Y(new_n13075_));
  AOI21X1  g10639(.A0(new_n13074_), .A1(pi0644), .B0(new_n13075_), .Y(new_n13076_));
  NOR3X1   g10640(.A(new_n13076_), .B(new_n13072_), .C(new_n11762_), .Y(new_n13077_));
  OAI21X1  g10641(.A0(new_n13070_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n13078_));
  AOI21X1  g10642(.A0(new_n13068_), .A1(new_n12612_), .B0(new_n13078_), .Y(new_n13079_));
  OAI21X1  g10643(.A0(new_n13054_), .A1(new_n12612_), .B0(pi0715), .Y(new_n13080_));
  AOI21X1  g10644(.A0(new_n13074_), .A1(new_n12612_), .B0(new_n13080_), .Y(new_n13081_));
  NOR3X1   g10645(.A(new_n13081_), .B(new_n13079_), .C(pi1160), .Y(new_n13082_));
  OAI21X1  g10646(.A0(new_n13082_), .A1(new_n13077_), .B0(pi0790), .Y(new_n13083_));
  AOI21X1  g10647(.A0(new_n13068_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n13084_));
  AOI22X1  g10648(.A0(new_n13084_), .A1(new_n13083_), .B0(new_n12966_), .B1(new_n12965_), .Y(po0298));
  INVX1    g10649(.A(pi0743), .Y(new_n13086_));
  NAND2X1  g10650(.A(new_n11973_), .B(new_n11968_), .Y(new_n13087_));
  NAND3X1  g10651(.A(new_n12311_), .B(new_n13087_), .C(pi0142), .Y(new_n13088_));
  OR3X1    g10652(.A(new_n12342_), .B(new_n12041_), .C(pi0142), .Y(new_n13089_));
  AOI21X1  g10653(.A0(new_n13089_), .A1(new_n13088_), .B0(new_n13086_), .Y(new_n13090_));
  OR3X1    g10654(.A(new_n12311_), .B(new_n12041_), .C(new_n2953_), .Y(new_n13091_));
  NAND2X1  g10655(.A(new_n13091_), .B(new_n13086_), .Y(new_n13092_));
  AOI21X1  g10656(.A0(new_n12793_), .A1(new_n2953_), .B0(new_n13092_), .Y(new_n13093_));
  NOR3X1   g10657(.A(new_n13093_), .B(new_n13090_), .C(pi0299), .Y(new_n13094_));
  OR3X1    g10658(.A(new_n12343_), .B(new_n12044_), .C(pi0142), .Y(new_n13095_));
  AND2X1   g10659(.A(new_n11966_), .B(pi0142), .Y(new_n13096_));
  OAI21X1  g10660(.A0(new_n12338_), .A1(new_n5019_), .B0(new_n13096_), .Y(new_n13097_));
  AOI21X1  g10661(.A0(new_n13097_), .A1(new_n13095_), .B0(new_n13086_), .Y(new_n13098_));
  OR4X1    g10662(.A(new_n12330_), .B(new_n12328_), .C(new_n5019_), .D(pi0142), .Y(new_n13099_));
  OR3X1    g10663(.A(new_n12313_), .B(new_n12044_), .C(new_n2953_), .Y(new_n13100_));
  AND3X1   g10664(.A(new_n13100_), .B(new_n13099_), .C(new_n13086_), .Y(new_n13101_));
  NOR3X1   g10665(.A(new_n13101_), .B(new_n13098_), .C(new_n2933_), .Y(new_n13102_));
  OR2X1    g10666(.A(new_n13102_), .B(new_n13094_), .Y(new_n13103_));
  OAI21X1  g10667(.A0(new_n12041_), .A1(pi0142), .B0(pi0743), .Y(new_n13104_));
  AOI21X1  g10668(.A0(new_n13087_), .A1(pi0142), .B0(new_n13104_), .Y(new_n13105_));
  OR2X1    g10669(.A(pi0743), .B(new_n2953_), .Y(new_n13106_));
  OAI21X1  g10670(.A0(new_n13106_), .A1(new_n11820_), .B0(new_n2933_), .Y(new_n13107_));
  NOR2X1   g10671(.A(new_n12044_), .B(pi0142), .Y(new_n13108_));
  AOI21X1  g10672(.A0(new_n11961_), .A1(pi0142), .B0(pi0743), .Y(new_n13109_));
  NOR3X1   g10673(.A(new_n13109_), .B(new_n13096_), .C(new_n13108_), .Y(new_n13110_));
  OAI22X1  g10674(.A0(new_n13110_), .A1(new_n2933_), .B0(new_n13107_), .B1(new_n13105_), .Y(new_n13111_));
  OAI21X1  g10675(.A0(new_n13111_), .A1(pi0735), .B0(new_n2939_), .Y(new_n13112_));
  AOI21X1  g10676(.A0(new_n13103_), .A1(pi0735), .B0(new_n13112_), .Y(new_n13113_));
  NAND3X1  g10677(.A(new_n12287_), .B(new_n12285_), .C(pi0142), .Y(new_n13114_));
  AOI21X1  g10678(.A0(new_n12255_), .A1(new_n2953_), .B0(new_n13086_), .Y(new_n13115_));
  OR2X1    g10679(.A(new_n12197_), .B(pi0142), .Y(new_n13116_));
  AOI21X1  g10680(.A0(new_n12114_), .A1(pi0142), .B0(pi0743), .Y(new_n13117_));
  AOI22X1  g10681(.A0(new_n13117_), .A1(new_n13116_), .B0(new_n13115_), .B1(new_n13114_), .Y(new_n13118_));
  OAI21X1  g10682(.A0(new_n11861_), .A1(new_n11847_), .B0(pi0142), .Y(new_n13119_));
  NAND2X1  g10683(.A(new_n13119_), .B(new_n13086_), .Y(new_n13120_));
  NOR3X1   g10684(.A(new_n12093_), .B(new_n12062_), .C(new_n13086_), .Y(new_n13121_));
  OAI21X1  g10685(.A0(new_n12024_), .A1(new_n2953_), .B0(new_n13121_), .Y(new_n13122_));
  NAND2X1  g10686(.A(new_n13122_), .B(new_n13120_), .Y(new_n13123_));
  MX2X1    g10687(.A(new_n13123_), .B(new_n13118_), .S0(pi0735), .Y(new_n13124_));
  AOI21X1  g10688(.A0(new_n12283_), .A1(pi0142), .B0(new_n13086_), .Y(new_n13125_));
  OAI21X1  g10689(.A0(new_n12242_), .A1(pi0142), .B0(new_n13125_), .Y(new_n13126_));
  AND3X1   g10690(.A(new_n12105_), .B(new_n12103_), .C(pi0142), .Y(new_n13127_));
  AND2X1   g10691(.A(new_n12199_), .B(new_n2953_), .Y(new_n13128_));
  OR2X1    g10692(.A(new_n13128_), .B(pi0743), .Y(new_n13129_));
  OAI21X1  g10693(.A0(new_n13129_), .A1(new_n13127_), .B0(new_n13126_), .Y(new_n13130_));
  OAI21X1  g10694(.A0(new_n11877_), .A1(new_n2953_), .B0(new_n13086_), .Y(new_n13131_));
  NOR3X1   g10695(.A(new_n12062_), .B(new_n12060_), .C(new_n13086_), .Y(new_n13132_));
  OAI21X1  g10696(.A0(new_n12016_), .A1(new_n2953_), .B0(new_n13132_), .Y(new_n13133_));
  AND2X1   g10697(.A(new_n13133_), .B(new_n13131_), .Y(new_n13134_));
  MX2X1    g10698(.A(new_n13134_), .B(new_n13130_), .S0(pi0735), .Y(new_n13135_));
  OAI21X1  g10699(.A0(new_n13135_), .A1(new_n5042_), .B0(pi0223), .Y(new_n13136_));
  AOI21X1  g10700(.A0(new_n13124_), .A1(new_n5042_), .B0(new_n13136_), .Y(new_n13137_));
  OR4X1    g10701(.A(new_n12271_), .B(new_n12270_), .C(new_n12266_), .D(new_n2953_), .Y(new_n13138_));
  AOI21X1  g10702(.A0(new_n12231_), .A1(new_n12228_), .B0(pi0142), .Y(new_n13139_));
  NOR2X1   g10703(.A(new_n13139_), .B(new_n13086_), .Y(new_n13140_));
  OR3X1    g10704(.A(new_n12130_), .B(new_n12122_), .C(new_n2953_), .Y(new_n13141_));
  AOI21X1  g10705(.A0(new_n12183_), .A1(new_n2953_), .B0(pi0743), .Y(new_n13142_));
  AOI22X1  g10706(.A0(new_n13142_), .A1(new_n13141_), .B0(new_n13140_), .B1(new_n13138_), .Y(new_n13143_));
  MX2X1    g10707(.A(new_n12052_), .B(new_n12005_), .S0(pi0142), .Y(new_n13144_));
  OR2X1    g10708(.A(new_n11924_), .B(new_n2953_), .Y(new_n13145_));
  MX2X1    g10709(.A(new_n13145_), .B(new_n13144_), .S0(pi0743), .Y(new_n13146_));
  MX2X1    g10710(.A(new_n13146_), .B(new_n13143_), .S0(pi0735), .Y(new_n13147_));
  OR2X1    g10711(.A(new_n13147_), .B(new_n5042_), .Y(new_n13148_));
  OAI21X1  g10712(.A0(new_n12222_), .A1(new_n12221_), .B0(new_n2953_), .Y(new_n13149_));
  OR4X1    g10713(.A(new_n12264_), .B(new_n12261_), .C(new_n12137_), .D(new_n2953_), .Y(new_n13150_));
  AND3X1   g10714(.A(new_n13150_), .B(new_n13149_), .C(pi0743), .Y(new_n13151_));
  NOR2X1   g10715(.A(new_n12162_), .B(new_n11881_), .Y(new_n13152_));
  AOI21X1  g10716(.A0(new_n12164_), .A1(new_n11881_), .B0(new_n13152_), .Y(new_n13153_));
  OAI21X1  g10717(.A0(new_n13153_), .A1(new_n12001_), .B0(new_n12160_), .Y(new_n13154_));
  AOI21X1  g10718(.A0(new_n13153_), .A1(new_n12167_), .B0(pi0616), .Y(new_n13155_));
  AOI22X1  g10719(.A0(new_n13155_), .A1(new_n13154_), .B0(new_n12161_), .B1(pi0616), .Y(new_n13156_));
  OAI21X1  g10720(.A0(new_n11863_), .A1(new_n5019_), .B0(new_n12172_), .Y(new_n13157_));
  OAI21X1  g10721(.A0(new_n13156_), .A1(new_n11863_), .B0(new_n13157_), .Y(new_n13158_));
  OAI21X1  g10722(.A0(new_n12139_), .A1(new_n2953_), .B0(new_n13086_), .Y(new_n13159_));
  AOI21X1  g10723(.A0(new_n13158_), .A1(new_n2953_), .B0(new_n13159_), .Y(new_n13160_));
  OAI21X1  g10724(.A0(new_n13160_), .A1(new_n13151_), .B0(pi0735), .Y(new_n13161_));
  OAI21X1  g10725(.A0(new_n11931_), .A1(new_n11927_), .B0(pi0142), .Y(new_n13162_));
  NAND2X1  g10726(.A(new_n13162_), .B(new_n13086_), .Y(new_n13163_));
  AOI21X1  g10727(.A0(new_n11989_), .A1(new_n11976_), .B0(new_n2953_), .Y(new_n13164_));
  MX2X1    g10728(.A(new_n12132_), .B(new_n11916_), .S0(new_n5020_), .Y(new_n13165_));
  OAI21X1  g10729(.A0(new_n12048_), .A1(new_n13165_), .B0(pi0743), .Y(new_n13166_));
  OR2X1    g10730(.A(new_n13166_), .B(new_n13164_), .Y(new_n13167_));
  NAND2X1  g10731(.A(new_n13167_), .B(new_n13163_), .Y(new_n13168_));
  OAI21X1  g10732(.A0(new_n13168_), .A1(pi0735), .B0(new_n13161_), .Y(new_n13169_));
  AOI21X1  g10733(.A0(new_n13169_), .A1(new_n5042_), .B0(new_n2951_), .Y(new_n13170_));
  INVX1    g10734(.A(pi0735), .Y(new_n13171_));
  AND2X1   g10735(.A(new_n11825_), .B(pi0142), .Y(new_n13172_));
  INVX1    g10736(.A(new_n13172_), .Y(new_n13173_));
  AOI22X1  g10737(.A0(new_n12049_), .A1(pi0743), .B0(new_n11825_), .B1(pi0142), .Y(new_n13174_));
  INVX1    g10738(.A(new_n11828_), .Y(new_n13175_));
  AND2X1   g10739(.A(new_n12056_), .B(pi0743), .Y(new_n13176_));
  AOI22X1  g10740(.A0(new_n13176_), .A1(new_n2987_), .B0(new_n13175_), .B1(pi0142), .Y(new_n13177_));
  OAI21X1  g10741(.A0(new_n12352_), .A1(new_n13175_), .B0(new_n13177_), .Y(new_n13178_));
  AOI21X1  g10742(.A0(new_n13178_), .A1(new_n12274_), .B0(new_n13171_), .Y(new_n13179_));
  AOI22X1  g10743(.A0(new_n13179_), .A1(new_n13173_), .B0(new_n13174_), .B1(new_n13171_), .Y(new_n13180_));
  OAI21X1  g10744(.A0(new_n13180_), .A1(new_n2952_), .B0(new_n2940_), .Y(new_n13181_));
  AOI21X1  g10745(.A0(new_n13170_), .A1(new_n13148_), .B0(new_n13181_), .Y(new_n13182_));
  OAI21X1  g10746(.A0(new_n13182_), .A1(new_n13137_), .B0(new_n2933_), .Y(new_n13183_));
  OAI21X1  g10747(.A0(new_n13135_), .A1(new_n5059_), .B0(pi0215), .Y(new_n13184_));
  AOI21X1  g10748(.A0(new_n13124_), .A1(new_n5059_), .B0(new_n13184_), .Y(new_n13185_));
  OR2X1    g10749(.A(new_n13147_), .B(new_n5059_), .Y(new_n13186_));
  AOI21X1  g10750(.A0(new_n13169_), .A1(new_n5059_), .B0(new_n10044_), .Y(new_n13187_));
  OAI21X1  g10751(.A0(new_n13180_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n13188_));
  AOI21X1  g10752(.A0(new_n13187_), .A1(new_n13186_), .B0(new_n13188_), .Y(new_n13189_));
  OAI21X1  g10753(.A0(new_n13189_), .A1(new_n13185_), .B0(pi0299), .Y(new_n13190_));
  AND3X1   g10754(.A(new_n13190_), .B(new_n13183_), .C(pi0039), .Y(new_n13191_));
  OAI21X1  g10755(.A0(new_n13191_), .A1(new_n13113_), .B0(new_n2979_), .Y(new_n13192_));
  AOI21X1  g10756(.A0(pi0142), .A1(pi0039), .B0(new_n2979_), .Y(new_n13193_));
  INVX1    g10757(.A(new_n13177_), .Y(new_n13194_));
  AND2X1   g10758(.A(new_n12353_), .B(pi0735), .Y(new_n13195_));
  OAI21X1  g10759(.A0(new_n13195_), .A1(new_n13194_), .B0(new_n2939_), .Y(new_n13196_));
  AOI21X1  g10760(.A0(new_n13196_), .A1(new_n13193_), .B0(new_n11770_), .Y(new_n13197_));
  AOI22X1  g10761(.A0(new_n13197_), .A1(new_n13192_), .B0(new_n11770_), .B1(pi0142), .Y(new_n13198_));
  OR2X1    g10762(.A(new_n3103_), .B(new_n2953_), .Y(new_n13199_));
  MX2X1    g10763(.A(new_n13168_), .B(new_n13146_), .S0(new_n5058_), .Y(new_n13200_));
  NOR2X1   g10764(.A(new_n13200_), .B(new_n10044_), .Y(new_n13201_));
  OAI21X1  g10765(.A0(new_n13174_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n13202_));
  AOI21X1  g10766(.A0(new_n13134_), .A1(new_n5058_), .B0(new_n2934_), .Y(new_n13203_));
  OAI21X1  g10767(.A0(new_n13123_), .A1(new_n5058_), .B0(new_n13203_), .Y(new_n13204_));
  OAI21X1  g10768(.A0(new_n13202_), .A1(new_n13201_), .B0(new_n13204_), .Y(new_n13205_));
  NAND3X1  g10769(.A(new_n13167_), .B(new_n13163_), .C(new_n5042_), .Y(new_n13206_));
  AND2X1   g10770(.A(new_n13206_), .B(new_n2952_), .Y(new_n13207_));
  OAI21X1  g10771(.A0(new_n13146_), .A1(new_n5042_), .B0(new_n13207_), .Y(new_n13208_));
  AOI21X1  g10772(.A0(new_n13174_), .A1(new_n2951_), .B0(pi0223), .Y(new_n13209_));
  AOI21X1  g10773(.A0(new_n13122_), .A1(new_n13120_), .B0(new_n5041_), .Y(new_n13210_));
  OAI21X1  g10774(.A0(new_n13134_), .A1(new_n5042_), .B0(pi0223), .Y(new_n13211_));
  OAI21X1  g10775(.A0(new_n13211_), .A1(new_n13210_), .B0(new_n2933_), .Y(new_n13212_));
  AOI21X1  g10776(.A0(new_n13209_), .A1(new_n13208_), .B0(new_n13212_), .Y(new_n13213_));
  OR2X1    g10777(.A(new_n13213_), .B(new_n2939_), .Y(new_n13214_));
  AOI21X1  g10778(.A0(new_n13205_), .A1(pi0299), .B0(new_n13214_), .Y(new_n13215_));
  OAI21X1  g10779(.A0(new_n13111_), .A1(pi0039), .B0(new_n2979_), .Y(new_n13216_));
  OAI21X1  g10780(.A0(new_n13177_), .A1(pi0039), .B0(new_n13193_), .Y(new_n13217_));
  AND2X1   g10781(.A(new_n13217_), .B(new_n3103_), .Y(new_n13218_));
  OAI21X1  g10782(.A0(new_n13216_), .A1(new_n13215_), .B0(new_n13218_), .Y(new_n13219_));
  NAND2X1  g10783(.A(new_n13219_), .B(new_n13199_), .Y(new_n13220_));
  OAI21X1  g10784(.A0(new_n13220_), .A1(pi0625), .B0(pi1153), .Y(new_n13221_));
  AOI21X1  g10785(.A0(new_n13198_), .A1(pi0625), .B0(new_n13221_), .Y(new_n13222_));
  NOR2X1   g10786(.A(new_n11924_), .B(new_n2953_), .Y(new_n13223_));
  MX2X1    g10787(.A(new_n12815_), .B(new_n12373_), .S0(new_n2953_), .Y(new_n13224_));
  MX2X1    g10788(.A(new_n13224_), .B(new_n13223_), .S0(new_n13171_), .Y(new_n13225_));
  MX2X1    g10789(.A(new_n12408_), .B(new_n12376_), .S0(new_n2953_), .Y(new_n13226_));
  MX2X1    g10790(.A(new_n13226_), .B(new_n13162_), .S0(new_n13171_), .Y(new_n13227_));
  OAI21X1  g10791(.A0(new_n13227_), .A1(new_n5058_), .B0(new_n10045_), .Y(new_n13228_));
  AOI21X1  g10792(.A0(new_n13225_), .A1(new_n5058_), .B0(new_n13228_), .Y(new_n13229_));
  AND2X1   g10793(.A(new_n12439_), .B(pi0735), .Y(new_n13230_));
  INVX1    g10794(.A(new_n13230_), .Y(new_n13231_));
  OAI22X1  g10795(.A0(new_n13231_), .A1(new_n11824_), .B0(new_n11880_), .B1(new_n2953_), .Y(new_n13232_));
  OAI21X1  g10796(.A0(new_n13232_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n13233_));
  NOR2X1   g10797(.A(new_n12419_), .B(new_n2953_), .Y(new_n13234_));
  INVX1    g10798(.A(new_n12245_), .Y(new_n13235_));
  OR4X1    g10799(.A(new_n12239_), .B(new_n12236_), .C(new_n5019_), .D(pi0142), .Y(new_n13236_));
  OAI21X1  g10800(.A0(new_n13236_), .A1(new_n13235_), .B0(pi0735), .Y(new_n13237_));
  NOR2X1   g10801(.A(new_n13237_), .B(new_n13234_), .Y(new_n13238_));
  AOI21X1  g10802(.A0(new_n13119_), .A1(new_n13171_), .B0(new_n13238_), .Y(new_n13239_));
  NOR2X1   g10803(.A(new_n11877_), .B(new_n2953_), .Y(new_n13240_));
  AND2X1   g10804(.A(new_n13236_), .B(pi0735), .Y(new_n13241_));
  OAI21X1  g10805(.A0(new_n12414_), .A1(new_n2953_), .B0(new_n13241_), .Y(new_n13242_));
  OAI21X1  g10806(.A0(new_n13240_), .A1(pi0735), .B0(new_n13242_), .Y(new_n13243_));
  AOI21X1  g10807(.A0(new_n13243_), .A1(new_n5058_), .B0(new_n2934_), .Y(new_n13244_));
  OAI21X1  g10808(.A0(new_n13239_), .A1(new_n5058_), .B0(new_n13244_), .Y(new_n13245_));
  AND2X1   g10809(.A(new_n13245_), .B(pi0299), .Y(new_n13246_));
  OAI21X1  g10810(.A0(new_n13233_), .A1(new_n13229_), .B0(new_n13246_), .Y(new_n13247_));
  OAI21X1  g10811(.A0(new_n13227_), .A1(new_n5041_), .B0(new_n2952_), .Y(new_n13248_));
  AOI21X1  g10812(.A0(new_n13225_), .A1(new_n5041_), .B0(new_n13248_), .Y(new_n13249_));
  OAI21X1  g10813(.A0(new_n13232_), .A1(new_n2952_), .B0(new_n2940_), .Y(new_n13250_));
  AOI21X1  g10814(.A0(new_n13243_), .A1(new_n5041_), .B0(new_n2940_), .Y(new_n13251_));
  OAI21X1  g10815(.A0(new_n13239_), .A1(new_n5041_), .B0(new_n13251_), .Y(new_n13252_));
  AND2X1   g10816(.A(new_n13252_), .B(new_n2933_), .Y(new_n13253_));
  OAI21X1  g10817(.A0(new_n13250_), .A1(new_n13249_), .B0(new_n13253_), .Y(new_n13254_));
  NAND3X1  g10818(.A(new_n13254_), .B(new_n13247_), .C(pi0039), .Y(new_n13255_));
  OAI21X1  g10819(.A0(new_n12340_), .A1(new_n2953_), .B0(pi0735), .Y(new_n13256_));
  AOI21X1  g10820(.A0(new_n12435_), .A1(new_n2953_), .B0(new_n13256_), .Y(new_n13257_));
  NOR3X1   g10821(.A(new_n11821_), .B(pi0735), .C(new_n2953_), .Y(new_n13258_));
  OAI21X1  g10822(.A0(new_n13258_), .A1(new_n13257_), .B0(new_n2939_), .Y(new_n13259_));
  NAND3X1  g10823(.A(new_n13259_), .B(new_n13255_), .C(new_n2979_), .Y(new_n13260_));
  AOI22X1  g10824(.A0(new_n13230_), .A1(new_n2987_), .B0(new_n13175_), .B1(pi0142), .Y(new_n13261_));
  OAI21X1  g10825(.A0(new_n13261_), .A1(pi0039), .B0(new_n13193_), .Y(new_n13262_));
  NAND3X1  g10826(.A(new_n13262_), .B(new_n13260_), .C(new_n3103_), .Y(new_n13263_));
  AND3X1   g10827(.A(new_n13263_), .B(new_n13199_), .C(new_n12363_), .Y(new_n13264_));
  NOR2X1   g10828(.A(new_n12446_), .B(new_n2979_), .Y(new_n13265_));
  NOR2X1   g10829(.A(new_n13265_), .B(new_n11770_), .Y(new_n13266_));
  NAND2X1  g10830(.A(new_n11937_), .B(pi0039), .Y(new_n13267_));
  AOI21X1  g10831(.A0(new_n11821_), .A1(new_n2939_), .B0(new_n2953_), .Y(new_n13268_));
  AND2X1   g10832(.A(new_n13119_), .B(new_n5059_), .Y(new_n13269_));
  OAI21X1  g10833(.A0(new_n13240_), .A1(new_n5059_), .B0(pi0215), .Y(new_n13270_));
  NAND2X1  g10834(.A(new_n13162_), .B(new_n5059_), .Y(new_n13271_));
  OAI21X1  g10835(.A0(new_n11924_), .A1(new_n2953_), .B0(new_n5058_), .Y(new_n13272_));
  AOI21X1  g10836(.A0(new_n13272_), .A1(new_n13271_), .B0(new_n10044_), .Y(new_n13273_));
  OAI21X1  g10837(.A0(new_n13172_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n13274_));
  OAI22X1  g10838(.A0(new_n13274_), .A1(new_n13273_), .B0(new_n13270_), .B1(new_n13269_), .Y(new_n13275_));
  AND3X1   g10839(.A(new_n13275_), .B(pi0299), .C(pi0039), .Y(new_n13276_));
  AOI21X1  g10840(.A0(new_n13268_), .A1(new_n13267_), .B0(new_n13276_), .Y(new_n13277_));
  OAI22X1  g10841(.A0(new_n13277_), .A1(new_n10655_), .B0(new_n13266_), .B1(new_n2953_), .Y(new_n13278_));
  OAI21X1  g10842(.A0(new_n13278_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n13279_));
  OAI21X1  g10843(.A0(new_n13279_), .A1(new_n13264_), .B0(pi0608), .Y(new_n13280_));
  OAI21X1  g10844(.A0(new_n13220_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n13281_));
  AOI21X1  g10845(.A0(new_n13198_), .A1(new_n12363_), .B0(new_n13281_), .Y(new_n13282_));
  AND3X1   g10846(.A(new_n13263_), .B(new_n13199_), .C(pi0625), .Y(new_n13283_));
  OAI21X1  g10847(.A0(new_n13278_), .A1(pi0625), .B0(pi1153), .Y(new_n13284_));
  OAI21X1  g10848(.A0(new_n13284_), .A1(new_n13283_), .B0(new_n12368_), .Y(new_n13285_));
  OAI22X1  g10849(.A0(new_n13285_), .A1(new_n13282_), .B0(new_n13280_), .B1(new_n13222_), .Y(new_n13286_));
  MX2X1    g10850(.A(new_n13286_), .B(new_n13198_), .S0(new_n11769_), .Y(new_n13287_));
  NAND2X1  g10851(.A(new_n13263_), .B(new_n13199_), .Y(new_n13288_));
  OAI22X1  g10852(.A0(new_n13284_), .A1(new_n13283_), .B0(new_n13279_), .B1(new_n13264_), .Y(new_n13289_));
  MX2X1    g10853(.A(new_n13289_), .B(new_n13288_), .S0(new_n11769_), .Y(new_n13290_));
  OAI21X1  g10854(.A0(new_n13290_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n13291_));
  AOI21X1  g10855(.A0(new_n13287_), .A1(new_n12462_), .B0(new_n13291_), .Y(new_n13292_));
  AOI21X1  g10856(.A0(new_n13219_), .A1(new_n13199_), .B0(new_n12473_), .Y(new_n13293_));
  AOI22X1  g10857(.A0(new_n13293_), .A1(pi0609), .B0(new_n13278_), .B1(new_n12472_), .Y(new_n13294_));
  OAI21X1  g10858(.A0(new_n13294_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n13295_));
  OAI21X1  g10859(.A0(new_n13290_), .A1(pi0609), .B0(pi1155), .Y(new_n13296_));
  AOI21X1  g10860(.A0(new_n13287_), .A1(pi0609), .B0(new_n13296_), .Y(new_n13297_));
  AOI22X1  g10861(.A0(new_n13293_), .A1(new_n12462_), .B0(new_n13278_), .B1(new_n12481_), .Y(new_n13298_));
  OAI21X1  g10862(.A0(new_n13298_), .A1(pi1155), .B0(pi0660), .Y(new_n13299_));
  OAI22X1  g10863(.A0(new_n13299_), .A1(new_n13297_), .B0(new_n13295_), .B1(new_n13292_), .Y(new_n13300_));
  MX2X1    g10864(.A(new_n13300_), .B(new_n13287_), .S0(new_n11768_), .Y(new_n13301_));
  MX2X1    g10865(.A(new_n13290_), .B(new_n13278_), .S0(new_n12490_), .Y(new_n13302_));
  OAI21X1  g10866(.A0(new_n13302_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13303_));
  AOI21X1  g10867(.A0(new_n13301_), .A1(new_n12486_), .B0(new_n13303_), .Y(new_n13304_));
  AOI21X1  g10868(.A0(new_n13278_), .A1(new_n12473_), .B0(new_n13293_), .Y(new_n13305_));
  MX2X1    g10869(.A(new_n13298_), .B(new_n13294_), .S0(pi1155), .Y(new_n13306_));
  MX2X1    g10870(.A(new_n13306_), .B(new_n13305_), .S0(new_n11768_), .Y(new_n13307_));
  OAI21X1  g10871(.A0(new_n13278_), .A1(pi0618), .B0(pi1154), .Y(new_n13308_));
  AOI21X1  g10872(.A0(new_n13307_), .A1(pi0618), .B0(new_n13308_), .Y(new_n13309_));
  OR2X1    g10873(.A(new_n13309_), .B(pi0627), .Y(new_n13310_));
  OAI21X1  g10874(.A0(new_n13302_), .A1(pi0618), .B0(pi1154), .Y(new_n13311_));
  AOI21X1  g10875(.A0(new_n13301_), .A1(pi0618), .B0(new_n13311_), .Y(new_n13312_));
  OAI21X1  g10876(.A0(new_n13278_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13313_));
  AOI21X1  g10877(.A0(new_n13307_), .A1(new_n12486_), .B0(new_n13313_), .Y(new_n13314_));
  OR2X1    g10878(.A(new_n13314_), .B(new_n12494_), .Y(new_n13315_));
  OAI22X1  g10879(.A0(new_n13315_), .A1(new_n13312_), .B0(new_n13310_), .B1(new_n13304_), .Y(new_n13316_));
  MX2X1    g10880(.A(new_n13316_), .B(new_n13301_), .S0(new_n11767_), .Y(new_n13317_));
  MX2X1    g10881(.A(new_n13302_), .B(new_n13278_), .S0(new_n12513_), .Y(new_n13318_));
  OAI21X1  g10882(.A0(new_n13318_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13319_));
  AOI21X1  g10883(.A0(new_n13317_), .A1(new_n12509_), .B0(new_n13319_), .Y(new_n13320_));
  OR2X1    g10884(.A(new_n13307_), .B(pi0781), .Y(new_n13321_));
  OAI21X1  g10885(.A0(new_n13314_), .A1(new_n13309_), .B0(pi0781), .Y(new_n13322_));
  AND2X1   g10886(.A(new_n13322_), .B(new_n13321_), .Y(new_n13323_));
  OAI21X1  g10887(.A0(new_n13278_), .A1(pi0619), .B0(pi1159), .Y(new_n13324_));
  AOI21X1  g10888(.A0(new_n13323_), .A1(pi0619), .B0(new_n13324_), .Y(new_n13325_));
  OR2X1    g10889(.A(new_n13325_), .B(pi0648), .Y(new_n13326_));
  OAI21X1  g10890(.A0(new_n13318_), .A1(pi0619), .B0(pi1159), .Y(new_n13327_));
  AOI21X1  g10891(.A0(new_n13317_), .A1(pi0619), .B0(new_n13327_), .Y(new_n13328_));
  OAI21X1  g10892(.A0(new_n13278_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13329_));
  AOI21X1  g10893(.A0(new_n13323_), .A1(new_n12509_), .B0(new_n13329_), .Y(new_n13330_));
  OR2X1    g10894(.A(new_n13330_), .B(new_n12517_), .Y(new_n13331_));
  OAI22X1  g10895(.A0(new_n13331_), .A1(new_n13328_), .B0(new_n13326_), .B1(new_n13320_), .Y(new_n13332_));
  MX2X1    g10896(.A(new_n13332_), .B(new_n13317_), .S0(new_n11766_), .Y(new_n13333_));
  MX2X1    g10897(.A(new_n13318_), .B(new_n13278_), .S0(new_n12531_), .Y(new_n13334_));
  AOI21X1  g10898(.A0(new_n13334_), .A1(pi0626), .B0(pi0641), .Y(new_n13335_));
  OAI21X1  g10899(.A0(new_n13333_), .A1(pi0626), .B0(new_n13335_), .Y(new_n13336_));
  INVX1    g10900(.A(new_n12535_), .Y(new_n13337_));
  OAI21X1  g10901(.A0(new_n13330_), .A1(new_n13325_), .B0(pi0789), .Y(new_n13338_));
  OAI21X1  g10902(.A0(new_n13323_), .A1(pi0789), .B0(new_n13338_), .Y(new_n13339_));
  INVX1    g10903(.A(new_n13278_), .Y(new_n13340_));
  AOI21X1  g10904(.A0(new_n13340_), .A1(pi0626), .B0(pi1158), .Y(new_n13341_));
  OAI21X1  g10905(.A0(new_n13339_), .A1(pi0626), .B0(new_n13341_), .Y(new_n13342_));
  NAND2X1  g10906(.A(new_n13342_), .B(new_n13337_), .Y(new_n13343_));
  AOI21X1  g10907(.A0(new_n13334_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n13344_));
  OAI21X1  g10908(.A0(new_n13333_), .A1(new_n12542_), .B0(new_n13344_), .Y(new_n13345_));
  INVX1    g10909(.A(new_n12546_), .Y(new_n13346_));
  AOI21X1  g10910(.A0(new_n13340_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n13347_));
  OAI21X1  g10911(.A0(new_n13339_), .A1(new_n12542_), .B0(new_n13347_), .Y(new_n13348_));
  NAND2X1  g10912(.A(new_n13348_), .B(new_n13346_), .Y(new_n13349_));
  AOI22X1  g10913(.A0(new_n13349_), .A1(new_n13345_), .B0(new_n13343_), .B1(new_n13336_), .Y(new_n13350_));
  MX2X1    g10914(.A(new_n13350_), .B(new_n13333_), .S0(new_n11765_), .Y(new_n13351_));
  NAND2X1  g10915(.A(new_n13348_), .B(new_n13342_), .Y(new_n13352_));
  MX2X1    g10916(.A(new_n13352_), .B(new_n13339_), .S0(new_n11765_), .Y(new_n13353_));
  OAI21X1  g10917(.A0(new_n13353_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13354_));
  AOI21X1  g10918(.A0(new_n13351_), .A1(new_n12554_), .B0(new_n13354_), .Y(new_n13355_));
  INVX1    g10919(.A(new_n12563_), .Y(new_n13356_));
  OR2X1    g10920(.A(new_n13278_), .B(new_n13356_), .Y(new_n13357_));
  OAI21X1  g10921(.A0(new_n13334_), .A1(new_n12563_), .B0(new_n13357_), .Y(new_n13358_));
  OAI21X1  g10922(.A0(new_n13278_), .A1(pi0628), .B0(pi1156), .Y(new_n13359_));
  AOI21X1  g10923(.A0(new_n13358_), .A1(pi0628), .B0(new_n13359_), .Y(new_n13360_));
  OR2X1    g10924(.A(new_n13360_), .B(pi0629), .Y(new_n13361_));
  OAI21X1  g10925(.A0(new_n13353_), .A1(pi0628), .B0(pi1156), .Y(new_n13362_));
  AOI21X1  g10926(.A0(new_n13351_), .A1(pi0628), .B0(new_n13362_), .Y(new_n13363_));
  OAI21X1  g10927(.A0(new_n13278_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13364_));
  AOI21X1  g10928(.A0(new_n13358_), .A1(new_n12554_), .B0(new_n13364_), .Y(new_n13365_));
  OR2X1    g10929(.A(new_n13365_), .B(new_n12561_), .Y(new_n13366_));
  OAI22X1  g10930(.A0(new_n13366_), .A1(new_n13363_), .B0(new_n13361_), .B1(new_n13355_), .Y(new_n13367_));
  MX2X1    g10931(.A(new_n13367_), .B(new_n13351_), .S0(new_n11764_), .Y(new_n13368_));
  MX2X1    g10932(.A(new_n13353_), .B(new_n13278_), .S0(new_n12580_), .Y(new_n13369_));
  OAI21X1  g10933(.A0(new_n13369_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13370_));
  AOI21X1  g10934(.A0(new_n13368_), .A1(new_n12577_), .B0(new_n13370_), .Y(new_n13371_));
  OAI21X1  g10935(.A0(new_n13365_), .A1(new_n13360_), .B0(pi0792), .Y(new_n13372_));
  OAI21X1  g10936(.A0(new_n13358_), .A1(pi0792), .B0(new_n13372_), .Y(new_n13373_));
  NOR2X1   g10937(.A(new_n13373_), .B(new_n12577_), .Y(new_n13374_));
  OAI21X1  g10938(.A0(new_n13278_), .A1(pi0647), .B0(pi1157), .Y(new_n13375_));
  OAI21X1  g10939(.A0(new_n13375_), .A1(new_n13374_), .B0(new_n12592_), .Y(new_n13376_));
  OAI21X1  g10940(.A0(new_n13369_), .A1(pi0647), .B0(pi1157), .Y(new_n13377_));
  AOI21X1  g10941(.A0(new_n13368_), .A1(pi0647), .B0(new_n13377_), .Y(new_n13378_));
  NOR2X1   g10942(.A(new_n13373_), .B(pi0647), .Y(new_n13379_));
  OAI21X1  g10943(.A0(new_n13278_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13380_));
  OAI21X1  g10944(.A0(new_n13380_), .A1(new_n13379_), .B0(pi0630), .Y(new_n13381_));
  OAI22X1  g10945(.A0(new_n13381_), .A1(new_n13378_), .B0(new_n13376_), .B1(new_n13371_), .Y(new_n13382_));
  MX2X1    g10946(.A(new_n13382_), .B(new_n13368_), .S0(new_n11763_), .Y(new_n13383_));
  OAI22X1  g10947(.A0(new_n13380_), .A1(new_n13379_), .B0(new_n13375_), .B1(new_n13374_), .Y(new_n13384_));
  MX2X1    g10948(.A(new_n13384_), .B(new_n13373_), .S0(new_n11763_), .Y(new_n13385_));
  OAI21X1  g10949(.A0(new_n13385_), .A1(pi0644), .B0(pi0715), .Y(new_n13386_));
  AOI21X1  g10950(.A0(new_n13383_), .A1(pi0644), .B0(new_n13386_), .Y(new_n13387_));
  AND2X1   g10951(.A(new_n13278_), .B(new_n12604_), .Y(new_n13388_));
  AOI21X1  g10952(.A0(new_n13369_), .A1(new_n12605_), .B0(new_n13388_), .Y(new_n13389_));
  OAI21X1  g10953(.A0(new_n13278_), .A1(pi0644), .B0(new_n12608_), .Y(new_n13390_));
  AOI21X1  g10954(.A0(new_n13389_), .A1(pi0644), .B0(new_n13390_), .Y(new_n13391_));
  OR3X1    g10955(.A(new_n13391_), .B(new_n13387_), .C(new_n11762_), .Y(new_n13392_));
  OAI21X1  g10956(.A0(new_n13385_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n13393_));
  AOI21X1  g10957(.A0(new_n13383_), .A1(new_n12612_), .B0(new_n13393_), .Y(new_n13394_));
  OAI21X1  g10958(.A0(new_n13278_), .A1(new_n12612_), .B0(pi0715), .Y(new_n13395_));
  AOI21X1  g10959(.A0(new_n13389_), .A1(new_n12612_), .B0(new_n13395_), .Y(new_n13396_));
  OR3X1    g10960(.A(new_n13396_), .B(new_n13394_), .C(pi1160), .Y(new_n13397_));
  AND3X1   g10961(.A(new_n13397_), .B(new_n13392_), .C(pi0790), .Y(new_n13398_));
  OAI21X1  g10962(.A0(new_n13383_), .A1(pi0790), .B0(new_n5102_), .Y(new_n13399_));
  AOI21X1  g10963(.A0(new_n5103_), .A1(new_n2953_), .B0(pi0057), .Y(new_n13400_));
  OAI21X1  g10964(.A0(new_n13399_), .A1(new_n13398_), .B0(new_n13400_), .Y(new_n13401_));
  AOI21X1  g10965(.A0(pi0142), .A1(pi0057), .B0(pi0832), .Y(new_n13402_));
  AND2X1   g10966(.A(new_n13176_), .B(new_n12474_), .Y(new_n13403_));
  AND3X1   g10967(.A(new_n13176_), .B(new_n12474_), .C(pi0609), .Y(new_n13404_));
  NOR2X1   g10968(.A(new_n2720_), .B(new_n2953_), .Y(new_n13405_));
  NOR3X1   g10969(.A(new_n13405_), .B(new_n13404_), .C(new_n12463_), .Y(new_n13406_));
  AND3X1   g10970(.A(new_n13176_), .B(new_n12474_), .C(new_n12462_), .Y(new_n13407_));
  NOR3X1   g10971(.A(new_n13407_), .B(new_n13405_), .C(pi1155), .Y(new_n13408_));
  OAI21X1  g10972(.A0(new_n13408_), .A1(new_n13406_), .B0(pi0785), .Y(new_n13409_));
  NOR2X1   g10973(.A(new_n13405_), .B(pi0785), .Y(new_n13410_));
  INVX1    g10974(.A(new_n13410_), .Y(new_n13411_));
  OAI21X1  g10975(.A0(new_n13411_), .A1(new_n13403_), .B0(new_n13409_), .Y(new_n13412_));
  AND2X1   g10976(.A(new_n13412_), .B(new_n11767_), .Y(new_n13413_));
  AOI21X1  g10977(.A0(new_n13405_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13414_));
  OAI21X1  g10978(.A0(new_n13412_), .A1(new_n12486_), .B0(new_n13414_), .Y(new_n13415_));
  AOI21X1  g10979(.A0(new_n13405_), .A1(pi0618), .B0(pi1154), .Y(new_n13416_));
  OAI21X1  g10980(.A0(new_n13412_), .A1(pi0618), .B0(new_n13416_), .Y(new_n13417_));
  AOI21X1  g10981(.A0(new_n13417_), .A1(new_n13415_), .B0(new_n11767_), .Y(new_n13418_));
  NOR2X1   g10982(.A(new_n13418_), .B(new_n13413_), .Y(new_n13419_));
  INVX1    g10983(.A(new_n13419_), .Y(new_n13420_));
  AOI21X1  g10984(.A0(new_n13405_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13421_));
  OAI21X1  g10985(.A0(new_n13420_), .A1(new_n12509_), .B0(new_n13421_), .Y(new_n13422_));
  AOI21X1  g10986(.A0(new_n13405_), .A1(pi0619), .B0(pi1159), .Y(new_n13423_));
  OAI21X1  g10987(.A0(new_n13420_), .A1(pi0619), .B0(new_n13423_), .Y(new_n13424_));
  AND2X1   g10988(.A(new_n13424_), .B(new_n13422_), .Y(new_n13425_));
  MX2X1    g10989(.A(new_n13425_), .B(new_n13419_), .S0(new_n11766_), .Y(new_n13426_));
  NAND2X1  g10990(.A(new_n13426_), .B(pi0626), .Y(new_n13427_));
  AOI21X1  g10991(.A0(new_n13405_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n13428_));
  NAND2X1  g10992(.A(new_n13426_), .B(new_n12542_), .Y(new_n13429_));
  AOI21X1  g10993(.A0(new_n13405_), .A1(pi0626), .B0(pi1158), .Y(new_n13430_));
  AOI22X1  g10994(.A0(new_n13430_), .A1(new_n13429_), .B0(new_n13428_), .B1(new_n13427_), .Y(new_n13431_));
  XOR2X1   g10995(.A(pi1153), .B(pi0625), .Y(new_n13432_));
  AND2X1   g10996(.A(new_n13432_), .B(pi0778), .Y(new_n13433_));
  INVX1    g10997(.A(new_n13433_), .Y(new_n13434_));
  AOI21X1  g10998(.A0(new_n13434_), .A1(new_n13230_), .B0(new_n13405_), .Y(new_n13435_));
  NOR3X1   g10999(.A(new_n13435_), .B(new_n12513_), .C(new_n12490_), .Y(new_n13436_));
  NOR2X1   g11000(.A(new_n13436_), .B(new_n13405_), .Y(new_n13437_));
  INVX1    g11001(.A(new_n13437_), .Y(new_n13438_));
  INVX1    g11002(.A(new_n12637_), .Y(new_n13439_));
  INVX1    g11003(.A(new_n13405_), .Y(new_n13440_));
  AOI21X1  g11004(.A0(new_n13440_), .A1(new_n12531_), .B0(new_n13439_), .Y(new_n13441_));
  AOI22X1  g11005(.A0(new_n13441_), .A1(new_n13438_), .B0(new_n13431_), .B1(new_n12639_), .Y(new_n13442_));
  NOR4X1   g11006(.A(new_n12084_), .B(new_n11991_), .C(new_n2725_), .D(new_n5019_), .Y(new_n13443_));
  AND2X1   g11007(.A(new_n13443_), .B(pi0735), .Y(new_n13444_));
  NOR3X1   g11008(.A(new_n13444_), .B(new_n13405_), .C(new_n13176_), .Y(new_n13445_));
  AND3X1   g11009(.A(new_n13443_), .B(pi0735), .C(pi0625), .Y(new_n13446_));
  OAI21X1  g11010(.A0(new_n13445_), .A1(new_n13446_), .B0(new_n12364_), .Y(new_n13447_));
  NAND3X1  g11011(.A(new_n12439_), .B(pi0735), .C(pi0625), .Y(new_n13448_));
  NOR2X1   g11012(.A(new_n13405_), .B(new_n12364_), .Y(new_n13449_));
  AOI21X1  g11013(.A0(new_n13449_), .A1(new_n13448_), .B0(pi0608), .Y(new_n13450_));
  OAI21X1  g11014(.A0(new_n13446_), .A1(new_n13176_), .B0(pi1153), .Y(new_n13451_));
  NAND4X1  g11015(.A(new_n12439_), .B(new_n12364_), .C(pi0735), .D(new_n12363_), .Y(new_n13452_));
  NAND3X1  g11016(.A(new_n13452_), .B(new_n13451_), .C(new_n13440_), .Y(new_n13453_));
  AOI22X1  g11017(.A0(new_n13453_), .A1(pi0608), .B0(new_n13450_), .B1(new_n13447_), .Y(new_n13454_));
  MX2X1    g11018(.A(new_n13454_), .B(new_n13445_), .S0(new_n11769_), .Y(new_n13455_));
  INVX1    g11019(.A(new_n13455_), .Y(new_n13456_));
  OAI21X1  g11020(.A0(new_n13435_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n13457_));
  AOI21X1  g11021(.A0(new_n13456_), .A1(new_n12462_), .B0(new_n13457_), .Y(new_n13458_));
  NOR3X1   g11022(.A(new_n13458_), .B(new_n13406_), .C(pi0660), .Y(new_n13459_));
  OAI21X1  g11023(.A0(new_n13435_), .A1(pi0609), .B0(pi1155), .Y(new_n13460_));
  AOI21X1  g11024(.A0(new_n13456_), .A1(pi0609), .B0(new_n13460_), .Y(new_n13461_));
  NOR3X1   g11025(.A(new_n13461_), .B(new_n13408_), .C(new_n12468_), .Y(new_n13462_));
  NOR2X1   g11026(.A(new_n13462_), .B(new_n13459_), .Y(new_n13463_));
  MX2X1    g11027(.A(new_n13463_), .B(new_n13455_), .S0(new_n11768_), .Y(new_n13464_));
  OAI21X1  g11028(.A0(new_n13435_), .A1(new_n12490_), .B0(new_n13440_), .Y(new_n13465_));
  AOI21X1  g11029(.A0(new_n13465_), .A1(pi0618), .B0(pi1154), .Y(new_n13466_));
  OAI21X1  g11030(.A0(new_n13464_), .A1(pi0618), .B0(new_n13466_), .Y(new_n13467_));
  AND2X1   g11031(.A(new_n13415_), .B(new_n12494_), .Y(new_n13468_));
  AOI21X1  g11032(.A0(new_n13465_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13469_));
  OAI21X1  g11033(.A0(new_n13464_), .A1(new_n12486_), .B0(new_n13469_), .Y(new_n13470_));
  AND2X1   g11034(.A(new_n13417_), .B(pi0627), .Y(new_n13471_));
  AOI22X1  g11035(.A0(new_n13471_), .A1(new_n13470_), .B0(new_n13468_), .B1(new_n13467_), .Y(new_n13472_));
  MX2X1    g11036(.A(new_n13472_), .B(new_n13464_), .S0(new_n11767_), .Y(new_n13473_));
  AOI21X1  g11037(.A0(new_n13438_), .A1(pi0619), .B0(pi1159), .Y(new_n13474_));
  OAI21X1  g11038(.A0(new_n13473_), .A1(pi0619), .B0(new_n13474_), .Y(new_n13475_));
  AND3X1   g11039(.A(new_n13475_), .B(new_n13422_), .C(new_n12517_), .Y(new_n13476_));
  AOI21X1  g11040(.A0(new_n13438_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13477_));
  OAI21X1  g11041(.A0(new_n13473_), .A1(new_n12509_), .B0(new_n13477_), .Y(new_n13478_));
  AND3X1   g11042(.A(new_n13478_), .B(new_n13424_), .C(pi0648), .Y(new_n13479_));
  NOR3X1   g11043(.A(new_n13479_), .B(new_n13476_), .C(new_n11766_), .Y(new_n13480_));
  INVX1    g11044(.A(new_n12709_), .Y(new_n13481_));
  AOI21X1  g11045(.A0(new_n13473_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n13482_));
  INVX1    g11046(.A(new_n13482_), .Y(new_n13483_));
  OAI22X1  g11047(.A0(new_n13483_), .A1(new_n13480_), .B0(new_n13442_), .B1(new_n11765_), .Y(new_n13484_));
  MX2X1    g11048(.A(new_n13431_), .B(new_n13426_), .S0(new_n11765_), .Y(new_n13485_));
  INVX1    g11049(.A(new_n13485_), .Y(new_n13486_));
  AOI21X1  g11050(.A0(new_n13486_), .A1(pi0628), .B0(pi1156), .Y(new_n13487_));
  OAI21X1  g11051(.A0(new_n13484_), .A1(pi0628), .B0(new_n13487_), .Y(new_n13488_));
  OR4X1    g11052(.A(new_n12563_), .B(new_n12531_), .C(new_n12513_), .D(new_n12490_), .Y(new_n13489_));
  OR3X1    g11053(.A(new_n13489_), .B(new_n13435_), .C(new_n12554_), .Y(new_n13490_));
  AOI21X1  g11054(.A0(new_n13490_), .A1(new_n13440_), .B0(new_n12555_), .Y(new_n13491_));
  OR2X1    g11055(.A(new_n13491_), .B(pi0629), .Y(new_n13492_));
  INVX1    g11056(.A(new_n13492_), .Y(new_n13493_));
  AOI21X1  g11057(.A0(new_n13486_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13494_));
  OAI21X1  g11058(.A0(new_n13484_), .A1(new_n12554_), .B0(new_n13494_), .Y(new_n13495_));
  NOR3X1   g11059(.A(new_n13489_), .B(new_n13435_), .C(pi0628), .Y(new_n13496_));
  OAI21X1  g11060(.A0(new_n13496_), .A1(new_n13405_), .B0(new_n12555_), .Y(new_n13497_));
  NAND2X1  g11061(.A(new_n13497_), .B(pi0629), .Y(new_n13498_));
  INVX1    g11062(.A(new_n13498_), .Y(new_n13499_));
  AOI22X1  g11063(.A0(new_n13499_), .A1(new_n13495_), .B0(new_n13493_), .B1(new_n13488_), .Y(new_n13500_));
  MX2X1    g11064(.A(new_n13500_), .B(new_n13484_), .S0(new_n11764_), .Y(new_n13501_));
  INVX1    g11065(.A(new_n13501_), .Y(new_n13502_));
  MX2X1    g11066(.A(new_n13486_), .B(new_n13440_), .S0(new_n12580_), .Y(new_n13503_));
  INVX1    g11067(.A(new_n13503_), .Y(new_n13504_));
  AOI21X1  g11068(.A0(new_n13504_), .A1(pi0647), .B0(pi1157), .Y(new_n13505_));
  OAI21X1  g11069(.A0(new_n13502_), .A1(pi0647), .B0(new_n13505_), .Y(new_n13506_));
  OAI21X1  g11070(.A0(pi1156), .A1(pi0628), .B0(pi0792), .Y(new_n13507_));
  AOI21X1  g11071(.A0(pi1156), .A1(pi0628), .B0(new_n13507_), .Y(new_n13508_));
  NOR4X1   g11072(.A(new_n13508_), .B(new_n13489_), .C(new_n13435_), .D(new_n12577_), .Y(new_n13509_));
  OR3X1    g11073(.A(new_n13509_), .B(new_n13405_), .C(new_n12578_), .Y(new_n13510_));
  AND2X1   g11074(.A(new_n13510_), .B(new_n12592_), .Y(new_n13511_));
  AOI21X1  g11075(.A0(new_n13504_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13512_));
  OAI21X1  g11076(.A0(new_n13502_), .A1(new_n12577_), .B0(new_n13512_), .Y(new_n13513_));
  NOR4X1   g11077(.A(new_n13508_), .B(new_n13489_), .C(new_n13435_), .D(pi0647), .Y(new_n13514_));
  OR3X1    g11078(.A(new_n13514_), .B(new_n13405_), .C(pi1157), .Y(new_n13515_));
  AND2X1   g11079(.A(new_n13515_), .B(pi0630), .Y(new_n13516_));
  AOI22X1  g11080(.A0(new_n13516_), .A1(new_n13513_), .B0(new_n13511_), .B1(new_n13506_), .Y(new_n13517_));
  MX2X1    g11081(.A(new_n13517_), .B(new_n13502_), .S0(new_n11763_), .Y(new_n13518_));
  XOR2X1   g11082(.A(pi1157), .B(new_n12577_), .Y(new_n13519_));
  NOR2X1   g11083(.A(new_n13519_), .B(new_n11763_), .Y(new_n13520_));
  NOR4X1   g11084(.A(new_n13520_), .B(new_n13508_), .C(new_n13489_), .D(new_n13435_), .Y(new_n13521_));
  OR2X1    g11085(.A(new_n13521_), .B(new_n13405_), .Y(new_n13522_));
  AOI21X1  g11086(.A0(new_n13522_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n13523_));
  OAI21X1  g11087(.A0(new_n13518_), .A1(new_n12612_), .B0(new_n13523_), .Y(new_n13524_));
  MX2X1    g11088(.A(new_n13503_), .B(new_n13440_), .S0(new_n12604_), .Y(new_n13525_));
  AOI21X1  g11089(.A0(new_n13405_), .A1(new_n12612_), .B0(pi0715), .Y(new_n13526_));
  OAI21X1  g11090(.A0(new_n13525_), .A1(new_n12612_), .B0(new_n13526_), .Y(new_n13527_));
  AND3X1   g11091(.A(new_n13527_), .B(new_n13524_), .C(pi1160), .Y(new_n13528_));
  AOI21X1  g11092(.A0(new_n13522_), .A1(pi0644), .B0(pi0715), .Y(new_n13529_));
  OAI21X1  g11093(.A0(new_n13518_), .A1(pi0644), .B0(new_n13529_), .Y(new_n13530_));
  AOI21X1  g11094(.A0(new_n13405_), .A1(pi0644), .B0(new_n12608_), .Y(new_n13531_));
  OAI21X1  g11095(.A0(new_n13525_), .A1(pi0644), .B0(new_n13531_), .Y(new_n13532_));
  AND3X1   g11096(.A(new_n13532_), .B(new_n13530_), .C(new_n11762_), .Y(new_n13533_));
  OAI21X1  g11097(.A0(new_n13533_), .A1(new_n13528_), .B0(pi0790), .Y(new_n13534_));
  OR2X1    g11098(.A(new_n13518_), .B(pi0790), .Y(new_n13535_));
  AND2X1   g11099(.A(new_n13535_), .B(pi0832), .Y(new_n13536_));
  AOI22X1  g11100(.A0(new_n13536_), .A1(new_n13534_), .B0(new_n13402_), .B1(new_n13401_), .Y(po0299));
  INVX1    g11101(.A(pi0687), .Y(new_n13538_));
  INVX1    g11102(.A(pi0143), .Y(new_n13539_));
  AND2X1   g11103(.A(new_n12352_), .B(new_n12077_), .Y(new_n13540_));
  INVX1    g11104(.A(new_n13540_), .Y(new_n13541_));
  MX2X1    g11105(.A(new_n12315_), .B(new_n12155_), .S0(pi0039), .Y(new_n13542_));
  MX2X1    g11106(.A(new_n13542_), .B(new_n13541_), .S0(pi0038), .Y(new_n13543_));
  MX2X1    g11107(.A(new_n12332_), .B(new_n12213_), .S0(pi0039), .Y(new_n13544_));
  OR2X1    g11108(.A(new_n13544_), .B(pi0038), .Y(new_n13545_));
  INVX1    g11109(.A(pi0774), .Y(new_n13546_));
  AND3X1   g11110(.A(new_n12353_), .B(new_n2939_), .C(pi0038), .Y(new_n13547_));
  NOR2X1   g11111(.A(new_n13547_), .B(new_n13546_), .Y(new_n13548_));
  OAI21X1  g11112(.A0(new_n13545_), .A1(new_n13539_), .B0(new_n13548_), .Y(new_n13549_));
  AOI21X1  g11113(.A0(new_n13543_), .A1(new_n13539_), .B0(new_n13549_), .Y(new_n13550_));
  NOR4X1   g11114(.A(new_n12206_), .B(new_n2985_), .C(new_n2536_), .D(pi0039), .Y(new_n13551_));
  NOR3X1   g11115(.A(new_n12344_), .B(new_n12045_), .C(pi0039), .Y(new_n13552_));
  AOI21X1  g11116(.A0(new_n12787_), .A1(pi0039), .B0(new_n13552_), .Y(new_n13553_));
  MX2X1    g11117(.A(new_n13553_), .B(new_n13551_), .S0(pi0038), .Y(new_n13554_));
  AND2X1   g11118(.A(new_n12788_), .B(pi0039), .Y(new_n13555_));
  OR3X1    g11119(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .Y(new_n13556_));
  AND3X1   g11120(.A(new_n13556_), .B(new_n2939_), .C(new_n2979_), .Y(new_n13557_));
  AOI21X1  g11121(.A0(new_n12276_), .A1(new_n2939_), .B0(new_n2979_), .Y(new_n13558_));
  NOR3X1   g11122(.A(new_n13558_), .B(new_n13557_), .C(new_n13555_), .Y(new_n13559_));
  OAI21X1  g11123(.A0(new_n13559_), .A1(pi0143), .B0(new_n13546_), .Y(new_n13560_));
  AOI21X1  g11124(.A0(new_n13554_), .A1(pi0143), .B0(new_n13560_), .Y(new_n13561_));
  OR3X1    g11125(.A(new_n13561_), .B(new_n13550_), .C(new_n13538_), .Y(new_n13562_));
  OAI21X1  g11126(.A0(new_n12447_), .A1(pi0143), .B0(pi0774), .Y(new_n13563_));
  AND3X1   g11127(.A(new_n12056_), .B(new_n2982_), .C(new_n2939_), .Y(new_n13564_));
  AND2X1   g11128(.A(new_n13564_), .B(pi0038), .Y(new_n13565_));
  AOI21X1  g11129(.A0(new_n12074_), .A1(new_n2979_), .B0(new_n13539_), .Y(new_n13566_));
  AOI21X1  g11130(.A0(new_n12018_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n13567_));
  AOI21X1  g11131(.A0(new_n12776_), .A1(new_n2979_), .B0(new_n13567_), .Y(new_n13568_));
  NOR2X1   g11132(.A(pi0774), .B(pi0143), .Y(new_n13569_));
  AOI21X1  g11133(.A0(new_n13569_), .A1(new_n13568_), .B0(new_n13566_), .Y(new_n13570_));
  OR2X1    g11134(.A(new_n13570_), .B(new_n13565_), .Y(new_n13571_));
  AND2X1   g11135(.A(new_n13571_), .B(new_n13563_), .Y(new_n13572_));
  AOI21X1  g11136(.A0(new_n13572_), .A1(new_n13538_), .B0(new_n11770_), .Y(new_n13573_));
  AOI22X1  g11137(.A0(new_n13573_), .A1(new_n13562_), .B0(new_n11770_), .B1(pi0143), .Y(new_n13574_));
  NAND2X1  g11138(.A(new_n13571_), .B(new_n13563_), .Y(new_n13575_));
  MX2X1    g11139(.A(new_n13575_), .B(pi0143), .S0(new_n11770_), .Y(new_n13576_));
  OAI21X1  g11140(.A0(new_n13576_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n13577_));
  AOI21X1  g11141(.A0(new_n13574_), .A1(new_n12363_), .B0(new_n13577_), .Y(new_n13578_));
  AND3X1   g11142(.A(new_n12832_), .B(new_n13538_), .C(new_n13539_), .Y(new_n13579_));
  OAI21X1  g11143(.A0(new_n12826_), .A1(new_n13539_), .B0(new_n2979_), .Y(new_n13580_));
  AOI21X1  g11144(.A0(new_n12825_), .A1(new_n13539_), .B0(new_n13580_), .Y(new_n13581_));
  OAI21X1  g11145(.A0(new_n12077_), .A1(pi0143), .B0(new_n12440_), .Y(new_n13582_));
  NAND2X1  g11146(.A(new_n13582_), .B(pi0687), .Y(new_n13583_));
  OAI21X1  g11147(.A0(new_n13583_), .A1(new_n13581_), .B0(new_n3103_), .Y(new_n13584_));
  OAI22X1  g11148(.A0(new_n13584_), .A1(new_n13579_), .B0(new_n3103_), .B1(new_n13539_), .Y(new_n13585_));
  AOI21X1  g11149(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0143), .Y(new_n13586_));
  AOI21X1  g11150(.A0(new_n13586_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n13587_));
  OAI21X1  g11151(.A0(new_n13585_), .A1(new_n12363_), .B0(new_n13587_), .Y(new_n13588_));
  NAND2X1  g11152(.A(new_n13588_), .B(new_n12368_), .Y(new_n13589_));
  OAI21X1  g11153(.A0(new_n13576_), .A1(pi0625), .B0(pi1153), .Y(new_n13590_));
  AOI21X1  g11154(.A0(new_n13574_), .A1(pi0625), .B0(new_n13590_), .Y(new_n13591_));
  AOI21X1  g11155(.A0(new_n13586_), .A1(pi0625), .B0(pi1153), .Y(new_n13592_));
  OAI21X1  g11156(.A0(new_n13585_), .A1(pi0625), .B0(new_n13592_), .Y(new_n13593_));
  NAND2X1  g11157(.A(new_n13593_), .B(pi0608), .Y(new_n13594_));
  OAI22X1  g11158(.A0(new_n13594_), .A1(new_n13591_), .B0(new_n13589_), .B1(new_n13578_), .Y(new_n13595_));
  MX2X1    g11159(.A(new_n13595_), .B(new_n13574_), .S0(new_n11769_), .Y(new_n13596_));
  NAND2X1  g11160(.A(new_n13593_), .B(new_n13588_), .Y(new_n13597_));
  MX2X1    g11161(.A(new_n13597_), .B(new_n13585_), .S0(new_n11769_), .Y(new_n13598_));
  OAI21X1  g11162(.A0(new_n13598_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n13599_));
  AOI21X1  g11163(.A0(new_n13596_), .A1(new_n12462_), .B0(new_n13599_), .Y(new_n13600_));
  INVX1    g11164(.A(new_n13586_), .Y(new_n13601_));
  AND2X1   g11165(.A(new_n13576_), .B(new_n12474_), .Y(new_n13602_));
  AOI22X1  g11166(.A0(new_n13602_), .A1(pi0609), .B0(new_n13601_), .B1(new_n12472_), .Y(new_n13603_));
  OAI21X1  g11167(.A0(new_n13603_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n13604_));
  OAI21X1  g11168(.A0(new_n13598_), .A1(pi0609), .B0(pi1155), .Y(new_n13605_));
  AOI21X1  g11169(.A0(new_n13596_), .A1(pi0609), .B0(new_n13605_), .Y(new_n13606_));
  AOI22X1  g11170(.A0(new_n13602_), .A1(new_n12462_), .B0(new_n13601_), .B1(new_n12481_), .Y(new_n13607_));
  OAI21X1  g11171(.A0(new_n13607_), .A1(pi1155), .B0(pi0660), .Y(new_n13608_));
  OAI22X1  g11172(.A0(new_n13608_), .A1(new_n13606_), .B0(new_n13604_), .B1(new_n13600_), .Y(new_n13609_));
  MX2X1    g11173(.A(new_n13609_), .B(new_n13596_), .S0(new_n11768_), .Y(new_n13610_));
  MX2X1    g11174(.A(new_n13598_), .B(new_n13601_), .S0(new_n12490_), .Y(new_n13611_));
  OAI21X1  g11175(.A0(new_n13611_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13612_));
  AOI21X1  g11176(.A0(new_n13610_), .A1(new_n12486_), .B0(new_n13612_), .Y(new_n13613_));
  AOI21X1  g11177(.A0(new_n13601_), .A1(new_n12473_), .B0(new_n13602_), .Y(new_n13614_));
  MX2X1    g11178(.A(new_n13607_), .B(new_n13603_), .S0(pi1155), .Y(new_n13615_));
  MX2X1    g11179(.A(new_n13615_), .B(new_n13614_), .S0(new_n11768_), .Y(new_n13616_));
  OAI21X1  g11180(.A0(new_n13601_), .A1(pi0618), .B0(pi1154), .Y(new_n13617_));
  AOI21X1  g11181(.A0(new_n13616_), .A1(pi0618), .B0(new_n13617_), .Y(new_n13618_));
  OR2X1    g11182(.A(new_n13618_), .B(pi0627), .Y(new_n13619_));
  OAI21X1  g11183(.A0(new_n13611_), .A1(pi0618), .B0(pi1154), .Y(new_n13620_));
  AOI21X1  g11184(.A0(new_n13610_), .A1(pi0618), .B0(new_n13620_), .Y(new_n13621_));
  OAI21X1  g11185(.A0(new_n13601_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13622_));
  AOI21X1  g11186(.A0(new_n13616_), .A1(new_n12486_), .B0(new_n13622_), .Y(new_n13623_));
  OR2X1    g11187(.A(new_n13623_), .B(new_n12494_), .Y(new_n13624_));
  OAI22X1  g11188(.A0(new_n13624_), .A1(new_n13621_), .B0(new_n13619_), .B1(new_n13613_), .Y(new_n13625_));
  MX2X1    g11189(.A(new_n13625_), .B(new_n13610_), .S0(new_n11767_), .Y(new_n13626_));
  MX2X1    g11190(.A(new_n13611_), .B(new_n13601_), .S0(new_n12513_), .Y(new_n13627_));
  OAI21X1  g11191(.A0(new_n13627_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13628_));
  AOI21X1  g11192(.A0(new_n13626_), .A1(new_n12509_), .B0(new_n13628_), .Y(new_n13629_));
  NOR2X1   g11193(.A(new_n13623_), .B(new_n13618_), .Y(new_n13630_));
  MX2X1    g11194(.A(new_n13630_), .B(new_n13616_), .S0(new_n11767_), .Y(new_n13631_));
  OAI21X1  g11195(.A0(new_n13601_), .A1(pi0619), .B0(pi1159), .Y(new_n13632_));
  AOI21X1  g11196(.A0(new_n13631_), .A1(pi0619), .B0(new_n13632_), .Y(new_n13633_));
  OR2X1    g11197(.A(new_n13633_), .B(pi0648), .Y(new_n13634_));
  OAI21X1  g11198(.A0(new_n13627_), .A1(pi0619), .B0(pi1159), .Y(new_n13635_));
  AOI21X1  g11199(.A0(new_n13626_), .A1(pi0619), .B0(new_n13635_), .Y(new_n13636_));
  OAI21X1  g11200(.A0(new_n13601_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13637_));
  AOI21X1  g11201(.A0(new_n13631_), .A1(new_n12509_), .B0(new_n13637_), .Y(new_n13638_));
  OR2X1    g11202(.A(new_n13638_), .B(new_n12517_), .Y(new_n13639_));
  OAI22X1  g11203(.A0(new_n13639_), .A1(new_n13636_), .B0(new_n13634_), .B1(new_n13629_), .Y(new_n13640_));
  MX2X1    g11204(.A(new_n13640_), .B(new_n13626_), .S0(new_n11766_), .Y(new_n13641_));
  MX2X1    g11205(.A(new_n13627_), .B(new_n13601_), .S0(new_n12531_), .Y(new_n13642_));
  AOI21X1  g11206(.A0(new_n13642_), .A1(pi0626), .B0(pi0641), .Y(new_n13643_));
  OAI21X1  g11207(.A0(new_n13641_), .A1(pi0626), .B0(new_n13643_), .Y(new_n13644_));
  OR2X1    g11208(.A(new_n13631_), .B(pi0789), .Y(new_n13645_));
  OAI21X1  g11209(.A0(new_n13638_), .A1(new_n13633_), .B0(pi0789), .Y(new_n13646_));
  NAND3X1  g11210(.A(new_n13646_), .B(new_n13645_), .C(new_n12542_), .Y(new_n13647_));
  AOI21X1  g11211(.A0(new_n13586_), .A1(pi0626), .B0(pi1158), .Y(new_n13648_));
  AND2X1   g11212(.A(new_n13648_), .B(new_n13647_), .Y(new_n13649_));
  OR2X1    g11213(.A(new_n13649_), .B(new_n12535_), .Y(new_n13650_));
  AOI21X1  g11214(.A0(new_n13642_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n13651_));
  OAI21X1  g11215(.A0(new_n13641_), .A1(new_n12542_), .B0(new_n13651_), .Y(new_n13652_));
  NAND3X1  g11216(.A(new_n13646_), .B(new_n13645_), .C(pi0626), .Y(new_n13653_));
  AOI21X1  g11217(.A0(new_n13586_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n13654_));
  AND2X1   g11218(.A(new_n13654_), .B(new_n13653_), .Y(new_n13655_));
  OR2X1    g11219(.A(new_n13655_), .B(new_n12546_), .Y(new_n13656_));
  AOI22X1  g11220(.A0(new_n13656_), .A1(new_n13652_), .B0(new_n13650_), .B1(new_n13644_), .Y(new_n13657_));
  MX2X1    g11221(.A(new_n13657_), .B(new_n13641_), .S0(new_n11765_), .Y(new_n13658_));
  NAND2X1  g11222(.A(new_n13646_), .B(new_n13645_), .Y(new_n13659_));
  OR2X1    g11223(.A(new_n13655_), .B(new_n13649_), .Y(new_n13660_));
  MX2X1    g11224(.A(new_n13660_), .B(new_n13659_), .S0(new_n11765_), .Y(new_n13661_));
  OAI21X1  g11225(.A0(new_n13661_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13662_));
  AOI21X1  g11226(.A0(new_n13658_), .A1(new_n12554_), .B0(new_n13662_), .Y(new_n13663_));
  MX2X1    g11227(.A(new_n13642_), .B(new_n13601_), .S0(new_n12563_), .Y(new_n13664_));
  AOI21X1  g11228(.A0(new_n13586_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13665_));
  OAI21X1  g11229(.A0(new_n13664_), .A1(new_n12554_), .B0(new_n13665_), .Y(new_n13666_));
  AND2X1   g11230(.A(new_n13666_), .B(new_n12561_), .Y(new_n13667_));
  INVX1    g11231(.A(new_n13667_), .Y(new_n13668_));
  OAI21X1  g11232(.A0(new_n13661_), .A1(pi0628), .B0(pi1156), .Y(new_n13669_));
  AOI21X1  g11233(.A0(new_n13658_), .A1(pi0628), .B0(new_n13669_), .Y(new_n13670_));
  AOI21X1  g11234(.A0(new_n13586_), .A1(pi0628), .B0(pi1156), .Y(new_n13671_));
  OAI21X1  g11235(.A0(new_n13664_), .A1(pi0628), .B0(new_n13671_), .Y(new_n13672_));
  AND2X1   g11236(.A(new_n13672_), .B(pi0629), .Y(new_n13673_));
  INVX1    g11237(.A(new_n13673_), .Y(new_n13674_));
  OAI22X1  g11238(.A0(new_n13674_), .A1(new_n13670_), .B0(new_n13668_), .B1(new_n13663_), .Y(new_n13675_));
  MX2X1    g11239(.A(new_n13675_), .B(new_n13658_), .S0(new_n11764_), .Y(new_n13676_));
  MX2X1    g11240(.A(new_n13661_), .B(new_n13601_), .S0(new_n12580_), .Y(new_n13677_));
  OAI21X1  g11241(.A0(new_n13677_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13678_));
  AOI21X1  g11242(.A0(new_n13676_), .A1(new_n12577_), .B0(new_n13678_), .Y(new_n13679_));
  AOI21X1  g11243(.A0(new_n13672_), .A1(new_n13666_), .B0(new_n11764_), .Y(new_n13680_));
  AOI21X1  g11244(.A0(new_n13664_), .A1(new_n11764_), .B0(new_n13680_), .Y(new_n13681_));
  OAI21X1  g11245(.A0(new_n13601_), .A1(pi0647), .B0(pi1157), .Y(new_n13682_));
  AOI21X1  g11246(.A0(new_n13681_), .A1(pi0647), .B0(new_n13682_), .Y(new_n13683_));
  NOR2X1   g11247(.A(new_n13683_), .B(pi0630), .Y(new_n13684_));
  INVX1    g11248(.A(new_n13684_), .Y(new_n13685_));
  OAI21X1  g11249(.A0(new_n13677_), .A1(pi0647), .B0(pi1157), .Y(new_n13686_));
  AOI21X1  g11250(.A0(new_n13676_), .A1(pi0647), .B0(new_n13686_), .Y(new_n13687_));
  OAI21X1  g11251(.A0(new_n13601_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13688_));
  AOI21X1  g11252(.A0(new_n13681_), .A1(new_n12577_), .B0(new_n13688_), .Y(new_n13689_));
  NOR2X1   g11253(.A(new_n13689_), .B(new_n12592_), .Y(new_n13690_));
  INVX1    g11254(.A(new_n13690_), .Y(new_n13691_));
  OAI22X1  g11255(.A0(new_n13691_), .A1(new_n13687_), .B0(new_n13685_), .B1(new_n13679_), .Y(new_n13692_));
  MX2X1    g11256(.A(new_n13692_), .B(new_n13676_), .S0(new_n11763_), .Y(new_n13693_));
  OAI21X1  g11257(.A0(new_n13689_), .A1(new_n13683_), .B0(pi0787), .Y(new_n13694_));
  OAI21X1  g11258(.A0(new_n13681_), .A1(pi0787), .B0(new_n13694_), .Y(new_n13695_));
  OAI21X1  g11259(.A0(new_n13695_), .A1(pi0644), .B0(pi0715), .Y(new_n13696_));
  AOI21X1  g11260(.A0(new_n13693_), .A1(pi0644), .B0(new_n13696_), .Y(new_n13697_));
  NOR2X1   g11261(.A(new_n13586_), .B(new_n12605_), .Y(new_n13698_));
  AOI21X1  g11262(.A0(new_n13677_), .A1(new_n12605_), .B0(new_n13698_), .Y(new_n13699_));
  OAI21X1  g11263(.A0(new_n13601_), .A1(pi0644), .B0(new_n12608_), .Y(new_n13700_));
  AOI21X1  g11264(.A0(new_n13699_), .A1(pi0644), .B0(new_n13700_), .Y(new_n13701_));
  NOR3X1   g11265(.A(new_n13701_), .B(new_n13697_), .C(new_n11762_), .Y(new_n13702_));
  OAI21X1  g11266(.A0(new_n13695_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n13703_));
  AOI21X1  g11267(.A0(new_n13693_), .A1(new_n12612_), .B0(new_n13703_), .Y(new_n13704_));
  OAI21X1  g11268(.A0(new_n13601_), .A1(new_n12612_), .B0(pi0715), .Y(new_n13705_));
  AOI21X1  g11269(.A0(new_n13699_), .A1(new_n12612_), .B0(new_n13705_), .Y(new_n13706_));
  OR2X1    g11270(.A(new_n13706_), .B(pi1160), .Y(new_n13707_));
  OAI21X1  g11271(.A0(new_n13707_), .A1(new_n13704_), .B0(pi0790), .Y(new_n13708_));
  OR2X1    g11272(.A(new_n13693_), .B(pi0790), .Y(new_n13709_));
  AND2X1   g11273(.A(new_n13709_), .B(new_n6489_), .Y(new_n13710_));
  OAI21X1  g11274(.A0(new_n13708_), .A1(new_n13702_), .B0(new_n13710_), .Y(new_n13711_));
  AOI21X1  g11275(.A0(po1038), .A1(new_n13539_), .B0(pi0832), .Y(new_n13712_));
  AOI21X1  g11276(.A0(pi1093), .A1(pi1092), .B0(pi0143), .Y(new_n13713_));
  AOI21X1  g11277(.A0(new_n12439_), .A1(pi0687), .B0(new_n13713_), .Y(new_n13714_));
  AND3X1   g11278(.A(new_n12439_), .B(pi0687), .C(new_n12363_), .Y(new_n13715_));
  NOR2X1   g11279(.A(new_n13715_), .B(new_n13714_), .Y(new_n13716_));
  OR2X1    g11280(.A(new_n13713_), .B(pi1153), .Y(new_n13717_));
  OAI22X1  g11281(.A0(new_n13717_), .A1(new_n13715_), .B0(new_n13716_), .B1(new_n12364_), .Y(new_n13718_));
  MX2X1    g11282(.A(new_n13718_), .B(new_n13714_), .S0(new_n11769_), .Y(new_n13719_));
  NOR3X1   g11283(.A(new_n13719_), .B(new_n12631_), .C(new_n12630_), .Y(new_n13720_));
  AND3X1   g11284(.A(new_n13720_), .B(new_n12637_), .C(new_n12634_), .Y(new_n13721_));
  AOI21X1  g11285(.A0(new_n12056_), .A1(new_n13546_), .B0(new_n13713_), .Y(new_n13722_));
  AOI21X1  g11286(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n13722_), .Y(new_n13723_));
  OAI21X1  g11287(.A0(new_n13722_), .A1(new_n12642_), .B0(pi1155), .Y(new_n13724_));
  INVX1    g11288(.A(new_n13724_), .Y(new_n13725_));
  AOI21X1  g11289(.A0(new_n13723_), .A1(new_n12646_), .B0(pi1155), .Y(new_n13726_));
  OAI21X1  g11290(.A0(new_n13726_), .A1(new_n13725_), .B0(pi0785), .Y(new_n13727_));
  OAI21X1  g11291(.A0(new_n13723_), .A1(pi0785), .B0(new_n13727_), .Y(new_n13728_));
  INVX1    g11292(.A(new_n13728_), .Y(new_n13729_));
  AOI21X1  g11293(.A0(new_n13729_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n13730_));
  AOI21X1  g11294(.A0(new_n13729_), .A1(new_n12655_), .B0(pi1154), .Y(new_n13731_));
  NOR2X1   g11295(.A(new_n13731_), .B(new_n13730_), .Y(new_n13732_));
  MX2X1    g11296(.A(new_n13732_), .B(new_n13729_), .S0(new_n11767_), .Y(new_n13733_));
  NOR2X1   g11297(.A(new_n13733_), .B(pi0789), .Y(new_n13734_));
  INVX1    g11298(.A(new_n13733_), .Y(new_n13735_));
  AOI21X1  g11299(.A0(new_n13713_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13736_));
  OAI21X1  g11300(.A0(new_n13735_), .A1(new_n12509_), .B0(new_n13736_), .Y(new_n13737_));
  AOI21X1  g11301(.A0(new_n13713_), .A1(pi0619), .B0(pi1159), .Y(new_n13738_));
  OAI21X1  g11302(.A0(new_n13735_), .A1(pi0619), .B0(new_n13738_), .Y(new_n13739_));
  AOI21X1  g11303(.A0(new_n13739_), .A1(new_n13737_), .B0(new_n11766_), .Y(new_n13740_));
  NOR2X1   g11304(.A(new_n13740_), .B(new_n13734_), .Y(new_n13741_));
  INVX1    g11305(.A(new_n13741_), .Y(new_n13742_));
  AOI21X1  g11306(.A0(new_n13713_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n13743_));
  OAI21X1  g11307(.A0(new_n13742_), .A1(new_n12542_), .B0(new_n13743_), .Y(new_n13744_));
  AOI21X1  g11308(.A0(new_n13713_), .A1(pi0626), .B0(pi1158), .Y(new_n13745_));
  OAI21X1  g11309(.A0(new_n13742_), .A1(pi0626), .B0(new_n13745_), .Y(new_n13746_));
  AND3X1   g11310(.A(new_n13746_), .B(new_n13744_), .C(new_n12639_), .Y(new_n13747_));
  OAI21X1  g11311(.A0(new_n13747_), .A1(new_n13721_), .B0(pi0788), .Y(new_n13748_));
  OAI21X1  g11312(.A0(new_n13714_), .A1(new_n11991_), .B0(new_n13722_), .Y(new_n13749_));
  OR3X1    g11313(.A(new_n13714_), .B(new_n11991_), .C(new_n12363_), .Y(new_n13750_));
  AOI21X1  g11314(.A0(new_n13749_), .A1(new_n13750_), .B0(new_n13717_), .Y(new_n13751_));
  OAI21X1  g11315(.A0(new_n13716_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n13752_));
  AND3X1   g11316(.A(new_n13750_), .B(new_n13722_), .C(pi1153), .Y(new_n13753_));
  OAI21X1  g11317(.A0(new_n13717_), .A1(new_n13715_), .B0(pi0608), .Y(new_n13754_));
  OAI22X1  g11318(.A0(new_n13754_), .A1(new_n13753_), .B0(new_n13752_), .B1(new_n13751_), .Y(new_n13755_));
  MX2X1    g11319(.A(new_n13755_), .B(new_n13749_), .S0(new_n11769_), .Y(new_n13756_));
  OAI21X1  g11320(.A0(new_n13719_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n13757_));
  AOI21X1  g11321(.A0(new_n13756_), .A1(new_n12462_), .B0(new_n13757_), .Y(new_n13758_));
  NAND2X1  g11322(.A(new_n13724_), .B(new_n12468_), .Y(new_n13759_));
  OAI21X1  g11323(.A0(new_n13719_), .A1(pi0609), .B0(pi1155), .Y(new_n13760_));
  AOI21X1  g11324(.A0(new_n13756_), .A1(pi0609), .B0(new_n13760_), .Y(new_n13761_));
  OR2X1    g11325(.A(new_n13726_), .B(new_n12468_), .Y(new_n13762_));
  OAI22X1  g11326(.A0(new_n13762_), .A1(new_n13761_), .B0(new_n13759_), .B1(new_n13758_), .Y(new_n13763_));
  MX2X1    g11327(.A(new_n13763_), .B(new_n13756_), .S0(new_n11768_), .Y(new_n13764_));
  OR2X1    g11328(.A(new_n13719_), .B(new_n12630_), .Y(new_n13765_));
  OAI21X1  g11329(.A0(new_n13765_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13766_));
  AOI21X1  g11330(.A0(new_n13764_), .A1(new_n12486_), .B0(new_n13766_), .Y(new_n13767_));
  OR2X1    g11331(.A(new_n13730_), .B(pi0627), .Y(new_n13768_));
  OAI21X1  g11332(.A0(new_n13765_), .A1(pi0618), .B0(pi1154), .Y(new_n13769_));
  AOI21X1  g11333(.A0(new_n13764_), .A1(pi0618), .B0(new_n13769_), .Y(new_n13770_));
  OR2X1    g11334(.A(new_n13731_), .B(new_n12494_), .Y(new_n13771_));
  OAI22X1  g11335(.A0(new_n13771_), .A1(new_n13770_), .B0(new_n13768_), .B1(new_n13767_), .Y(new_n13772_));
  MX2X1    g11336(.A(new_n13772_), .B(new_n13764_), .S0(new_n11767_), .Y(new_n13773_));
  NAND2X1  g11337(.A(new_n13773_), .B(new_n12509_), .Y(new_n13774_));
  AOI21X1  g11338(.A0(new_n13720_), .A1(pi0619), .B0(pi1159), .Y(new_n13775_));
  NAND2X1  g11339(.A(new_n13737_), .B(new_n12517_), .Y(new_n13776_));
  AOI21X1  g11340(.A0(new_n13775_), .A1(new_n13774_), .B0(new_n13776_), .Y(new_n13777_));
  NAND2X1  g11341(.A(new_n13773_), .B(pi0619), .Y(new_n13778_));
  AOI21X1  g11342(.A0(new_n13720_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13779_));
  NAND2X1  g11343(.A(new_n13739_), .B(pi0648), .Y(new_n13780_));
  AOI21X1  g11344(.A0(new_n13779_), .A1(new_n13778_), .B0(new_n13780_), .Y(new_n13781_));
  NOR3X1   g11345(.A(new_n13781_), .B(new_n13777_), .C(new_n11766_), .Y(new_n13782_));
  OAI21X1  g11346(.A0(new_n13773_), .A1(pi0789), .B0(new_n12709_), .Y(new_n13783_));
  OAI21X1  g11347(.A0(new_n13783_), .A1(new_n13782_), .B0(new_n13748_), .Y(new_n13784_));
  AND2X1   g11348(.A(new_n13746_), .B(new_n13744_), .Y(new_n13785_));
  MX2X1    g11349(.A(new_n13785_), .B(new_n13741_), .S0(new_n11765_), .Y(new_n13786_));
  INVX1    g11350(.A(new_n13786_), .Y(new_n13787_));
  OAI21X1  g11351(.A0(new_n13787_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13788_));
  AOI21X1  g11352(.A0(new_n13784_), .A1(new_n12554_), .B0(new_n13788_), .Y(new_n13789_));
  AND3X1   g11353(.A(new_n13720_), .B(new_n12718_), .C(new_n12634_), .Y(new_n13790_));
  INVX1    g11354(.A(new_n13790_), .Y(new_n13791_));
  AOI21X1  g11355(.A0(new_n2720_), .A1(new_n12554_), .B0(new_n13791_), .Y(new_n13792_));
  OAI21X1  g11356(.A0(new_n13792_), .A1(new_n12555_), .B0(new_n12561_), .Y(new_n13793_));
  OAI21X1  g11357(.A0(new_n13787_), .A1(pi0628), .B0(pi1156), .Y(new_n13794_));
  AOI21X1  g11358(.A0(new_n13784_), .A1(pi0628), .B0(new_n13794_), .Y(new_n13795_));
  AOI21X1  g11359(.A0(new_n2720_), .A1(pi0628), .B0(new_n13791_), .Y(new_n13796_));
  OAI21X1  g11360(.A0(new_n13796_), .A1(pi1156), .B0(pi0629), .Y(new_n13797_));
  OAI22X1  g11361(.A0(new_n13797_), .A1(new_n13795_), .B0(new_n13793_), .B1(new_n13789_), .Y(new_n13798_));
  MX2X1    g11362(.A(new_n13798_), .B(new_n13784_), .S0(new_n11764_), .Y(new_n13799_));
  INVX1    g11363(.A(new_n13713_), .Y(new_n13800_));
  MX2X1    g11364(.A(new_n13787_), .B(new_n13800_), .S0(new_n12580_), .Y(new_n13801_));
  OAI21X1  g11365(.A0(new_n13801_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13802_));
  AOI21X1  g11366(.A0(new_n13799_), .A1(new_n12577_), .B0(new_n13802_), .Y(new_n13803_));
  AND2X1   g11367(.A(new_n13790_), .B(new_n12739_), .Y(new_n13804_));
  OAI21X1  g11368(.A0(new_n13800_), .A1(pi0647), .B0(pi1157), .Y(new_n13805_));
  AOI21X1  g11369(.A0(new_n13804_), .A1(pi0647), .B0(new_n13805_), .Y(new_n13806_));
  OR2X1    g11370(.A(new_n13806_), .B(pi0630), .Y(new_n13807_));
  OAI21X1  g11371(.A0(new_n13801_), .A1(pi0647), .B0(pi1157), .Y(new_n13808_));
  AOI21X1  g11372(.A0(new_n13799_), .A1(pi0647), .B0(new_n13808_), .Y(new_n13809_));
  OAI21X1  g11373(.A0(new_n13800_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13810_));
  AOI21X1  g11374(.A0(new_n13804_), .A1(new_n12577_), .B0(new_n13810_), .Y(new_n13811_));
  OR2X1    g11375(.A(new_n13811_), .B(new_n12592_), .Y(new_n13812_));
  OAI22X1  g11376(.A0(new_n13812_), .A1(new_n13809_), .B0(new_n13807_), .B1(new_n13803_), .Y(new_n13813_));
  MX2X1    g11377(.A(new_n13813_), .B(new_n13799_), .S0(new_n11763_), .Y(new_n13814_));
  OAI21X1  g11378(.A0(new_n13811_), .A1(new_n13806_), .B0(pi0787), .Y(new_n13815_));
  OAI21X1  g11379(.A0(new_n13804_), .A1(pi0787), .B0(new_n13815_), .Y(new_n13816_));
  OAI21X1  g11380(.A0(new_n13816_), .A1(pi0644), .B0(pi0715), .Y(new_n13817_));
  AOI21X1  g11381(.A0(new_n13814_), .A1(pi0644), .B0(new_n13817_), .Y(new_n13818_));
  NOR3X1   g11382(.A(new_n13713_), .B(new_n12603_), .C(new_n11763_), .Y(new_n13819_));
  AOI21X1  g11383(.A0(new_n13801_), .A1(new_n12605_), .B0(new_n13819_), .Y(new_n13820_));
  OAI21X1  g11384(.A0(new_n13800_), .A1(pi0644), .B0(new_n12608_), .Y(new_n13821_));
  AOI21X1  g11385(.A0(new_n13820_), .A1(pi0644), .B0(new_n13821_), .Y(new_n13822_));
  NOR3X1   g11386(.A(new_n13822_), .B(new_n13818_), .C(new_n11762_), .Y(new_n13823_));
  OAI21X1  g11387(.A0(new_n13816_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n13824_));
  AOI21X1  g11388(.A0(new_n13814_), .A1(new_n12612_), .B0(new_n13824_), .Y(new_n13825_));
  OAI21X1  g11389(.A0(new_n13800_), .A1(new_n12612_), .B0(pi0715), .Y(new_n13826_));
  AOI21X1  g11390(.A0(new_n13820_), .A1(new_n12612_), .B0(new_n13826_), .Y(new_n13827_));
  NOR3X1   g11391(.A(new_n13827_), .B(new_n13825_), .C(pi1160), .Y(new_n13828_));
  OAI21X1  g11392(.A0(new_n13828_), .A1(new_n13823_), .B0(pi0790), .Y(new_n13829_));
  AOI21X1  g11393(.A0(new_n13814_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n13830_));
  AOI22X1  g11394(.A0(new_n13830_), .A1(new_n13829_), .B0(new_n13712_), .B1(new_n13711_), .Y(po0300));
  INVX1    g11395(.A(pi0736), .Y(new_n13832_));
  AOI21X1  g11396(.A0(new_n11957_), .A1(new_n11937_), .B0(pi0758), .Y(new_n13833_));
  AND2X1   g11397(.A(new_n12034_), .B(pi0758), .Y(new_n13834_));
  OAI21X1  g11398(.A0(new_n13834_), .A1(new_n13833_), .B0(pi0039), .Y(new_n13835_));
  INVX1    g11399(.A(pi0758), .Y(new_n13836_));
  AOI21X1  g11400(.A0(new_n11821_), .A1(new_n13836_), .B0(pi0039), .Y(new_n13837_));
  OAI21X1  g11401(.A0(new_n11975_), .A1(new_n13836_), .B0(new_n13837_), .Y(new_n13838_));
  AOI21X1  g11402(.A0(new_n13838_), .A1(new_n13835_), .B0(new_n7344_), .Y(new_n13839_));
  AND3X1   g11403(.A(new_n12074_), .B(pi0758), .C(new_n7344_), .Y(new_n13840_));
  OAI21X1  g11404(.A0(new_n13840_), .A1(new_n13839_), .B0(new_n2979_), .Y(new_n13841_));
  NOR2X1   g11405(.A(new_n12077_), .B(pi0144), .Y(new_n13842_));
  AOI21X1  g11406(.A0(new_n11991_), .A1(pi0758), .B0(new_n12771_), .Y(new_n13843_));
  NOR3X1   g11407(.A(new_n13843_), .B(new_n13842_), .C(new_n2979_), .Y(new_n13844_));
  INVX1    g11408(.A(new_n13844_), .Y(new_n13845_));
  AND3X1   g11409(.A(new_n13845_), .B(new_n13841_), .C(new_n13832_), .Y(new_n13846_));
  AOI21X1  g11410(.A0(new_n12213_), .A1(new_n7344_), .B0(pi0758), .Y(new_n13847_));
  OAI21X1  g11411(.A0(new_n12155_), .A1(new_n7344_), .B0(new_n13847_), .Y(new_n13848_));
  AOI21X1  g11412(.A0(new_n12301_), .A1(pi0144), .B0(new_n13836_), .Y(new_n13849_));
  OAI21X1  g11413(.A0(new_n12260_), .A1(pi0144), .B0(new_n13849_), .Y(new_n13850_));
  AND3X1   g11414(.A(new_n13850_), .B(new_n13848_), .C(pi0039), .Y(new_n13851_));
  OAI21X1  g11415(.A0(new_n12315_), .A1(new_n7344_), .B0(new_n13836_), .Y(new_n13852_));
  AOI21X1  g11416(.A0(new_n12332_), .A1(new_n7344_), .B0(new_n13852_), .Y(new_n13853_));
  NOR4X1   g11417(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(new_n7344_), .Y(new_n13854_));
  OAI21X1  g11418(.A0(new_n12800_), .A1(pi0144), .B0(pi0758), .Y(new_n13855_));
  OAI21X1  g11419(.A0(new_n13855_), .A1(new_n13854_), .B0(new_n2939_), .Y(new_n13856_));
  OAI21X1  g11420(.A0(new_n13856_), .A1(new_n13853_), .B0(new_n2979_), .Y(new_n13857_));
  NOR3X1   g11421(.A(new_n13844_), .B(new_n13547_), .C(new_n13832_), .Y(new_n13858_));
  OAI21X1  g11422(.A0(new_n13857_), .A1(new_n13851_), .B0(new_n13858_), .Y(new_n13859_));
  NAND2X1  g11423(.A(new_n13859_), .B(new_n3103_), .Y(new_n13860_));
  OAI22X1  g11424(.A0(new_n13860_), .A1(new_n13846_), .B0(new_n3103_), .B1(new_n7344_), .Y(new_n13861_));
  OR2X1    g11425(.A(new_n13861_), .B(pi0625), .Y(new_n13862_));
  AND2X1   g11426(.A(new_n13845_), .B(new_n13841_), .Y(new_n13863_));
  MX2X1    g11427(.A(new_n13863_), .B(new_n7344_), .S0(new_n11770_), .Y(new_n13864_));
  AOI21X1  g11428(.A0(new_n13864_), .A1(pi0625), .B0(pi1153), .Y(new_n13865_));
  AOI21X1  g11429(.A0(new_n12447_), .A1(new_n3103_), .B0(new_n7344_), .Y(new_n13866_));
  NOR4X1   g11430(.A(new_n10543_), .B(new_n13832_), .C(pi0100), .D(pi0087), .Y(new_n13867_));
  MX2X1    g11431(.A(new_n12432_), .B(new_n12314_), .S0(new_n2939_), .Y(new_n13868_));
  NAND2X1  g11432(.A(new_n12344_), .B(new_n2939_), .Y(new_n13869_));
  OAI21X1  g11433(.A0(new_n12394_), .A1(new_n2939_), .B0(new_n13869_), .Y(new_n13870_));
  OAI21X1  g11434(.A0(new_n13870_), .A1(pi0144), .B0(new_n2979_), .Y(new_n13871_));
  AOI21X1  g11435(.A0(new_n13868_), .A1(pi0144), .B0(new_n13871_), .Y(new_n13872_));
  AOI21X1  g11436(.A0(new_n12275_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n13873_));
  INVX1    g11437(.A(new_n13873_), .Y(new_n13874_));
  OAI21X1  g11438(.A0(new_n13874_), .A1(new_n13842_), .B0(new_n13867_), .Y(new_n13875_));
  OAI22X1  g11439(.A0(new_n13875_), .A1(new_n13872_), .B0(new_n13867_), .B1(new_n13866_), .Y(new_n13876_));
  OAI21X1  g11440(.A0(new_n13866_), .A1(pi0625), .B0(pi1153), .Y(new_n13877_));
  AOI21X1  g11441(.A0(new_n13876_), .A1(pi0625), .B0(new_n13877_), .Y(new_n13878_));
  OR2X1    g11442(.A(new_n13878_), .B(pi0608), .Y(new_n13879_));
  AOI21X1  g11443(.A0(new_n13865_), .A1(new_n13862_), .B0(new_n13879_), .Y(new_n13880_));
  OR2X1    g11444(.A(new_n13861_), .B(new_n12363_), .Y(new_n13881_));
  AOI21X1  g11445(.A0(new_n13864_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n13882_));
  OAI21X1  g11446(.A0(new_n13866_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n13883_));
  AOI21X1  g11447(.A0(new_n13876_), .A1(new_n12363_), .B0(new_n13883_), .Y(new_n13884_));
  OR2X1    g11448(.A(new_n13884_), .B(new_n12368_), .Y(new_n13885_));
  AOI21X1  g11449(.A0(new_n13882_), .A1(new_n13881_), .B0(new_n13885_), .Y(new_n13886_));
  OAI21X1  g11450(.A0(new_n13886_), .A1(new_n13880_), .B0(pi0778), .Y(new_n13887_));
  OR2X1    g11451(.A(new_n13861_), .B(pi0778), .Y(new_n13888_));
  AOI21X1  g11452(.A0(new_n13888_), .A1(new_n13887_), .B0(pi0609), .Y(new_n13889_));
  OR2X1    g11453(.A(new_n13876_), .B(pi0778), .Y(new_n13890_));
  NOR2X1   g11454(.A(new_n13884_), .B(new_n13878_), .Y(new_n13891_));
  OAI21X1  g11455(.A0(new_n13891_), .A1(new_n11769_), .B0(new_n13890_), .Y(new_n13892_));
  OAI21X1  g11456(.A0(new_n13892_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n13893_));
  NOR2X1   g11457(.A(new_n13866_), .B(new_n12474_), .Y(new_n13894_));
  AOI21X1  g11458(.A0(new_n13864_), .A1(new_n12474_), .B0(new_n13894_), .Y(new_n13895_));
  INVX1    g11459(.A(new_n13866_), .Y(new_n13896_));
  AOI21X1  g11460(.A0(new_n13896_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n13897_));
  OAI21X1  g11461(.A0(new_n13895_), .A1(new_n12462_), .B0(new_n13897_), .Y(new_n13898_));
  AND2X1   g11462(.A(new_n13898_), .B(new_n12468_), .Y(new_n13899_));
  OAI21X1  g11463(.A0(new_n13893_), .A1(new_n13889_), .B0(new_n13899_), .Y(new_n13900_));
  AOI21X1  g11464(.A0(new_n13888_), .A1(new_n13887_), .B0(new_n12462_), .Y(new_n13901_));
  OAI21X1  g11465(.A0(new_n13892_), .A1(pi0609), .B0(pi1155), .Y(new_n13902_));
  AOI21X1  g11466(.A0(new_n13896_), .A1(pi0609), .B0(pi1155), .Y(new_n13903_));
  OAI21X1  g11467(.A0(new_n13895_), .A1(pi0609), .B0(new_n13903_), .Y(new_n13904_));
  AND2X1   g11468(.A(new_n13904_), .B(pi0660), .Y(new_n13905_));
  OAI21X1  g11469(.A0(new_n13902_), .A1(new_n13901_), .B0(new_n13905_), .Y(new_n13906_));
  AOI21X1  g11470(.A0(new_n13906_), .A1(new_n13900_), .B0(new_n11768_), .Y(new_n13907_));
  AOI21X1  g11471(.A0(new_n13888_), .A1(new_n13887_), .B0(pi0785), .Y(new_n13908_));
  OAI21X1  g11472(.A0(new_n13908_), .A1(new_n13907_), .B0(new_n12486_), .Y(new_n13909_));
  INVX1    g11473(.A(new_n12490_), .Y(new_n13910_));
  OR2X1    g11474(.A(new_n13866_), .B(new_n13910_), .Y(new_n13911_));
  OAI21X1  g11475(.A0(new_n13892_), .A1(new_n12490_), .B0(new_n13911_), .Y(new_n13912_));
  AOI21X1  g11476(.A0(new_n13912_), .A1(pi0618), .B0(pi1154), .Y(new_n13913_));
  AOI21X1  g11477(.A0(new_n13904_), .A1(new_n13898_), .B0(new_n11768_), .Y(new_n13914_));
  AOI21X1  g11478(.A0(new_n13895_), .A1(new_n11768_), .B0(new_n13914_), .Y(new_n13915_));
  OAI21X1  g11479(.A0(new_n13866_), .A1(pi0618), .B0(pi1154), .Y(new_n13916_));
  AOI21X1  g11480(.A0(new_n13915_), .A1(pi0618), .B0(new_n13916_), .Y(new_n13917_));
  OR2X1    g11481(.A(new_n13917_), .B(pi0627), .Y(new_n13918_));
  AOI21X1  g11482(.A0(new_n13913_), .A1(new_n13909_), .B0(new_n13918_), .Y(new_n13919_));
  OAI21X1  g11483(.A0(new_n13908_), .A1(new_n13907_), .B0(pi0618), .Y(new_n13920_));
  AOI21X1  g11484(.A0(new_n13912_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13921_));
  OAI21X1  g11485(.A0(new_n13866_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n13922_));
  AOI21X1  g11486(.A0(new_n13915_), .A1(new_n12486_), .B0(new_n13922_), .Y(new_n13923_));
  OR2X1    g11487(.A(new_n13923_), .B(new_n12494_), .Y(new_n13924_));
  AOI21X1  g11488(.A0(new_n13921_), .A1(new_n13920_), .B0(new_n13924_), .Y(new_n13925_));
  OAI21X1  g11489(.A0(new_n13925_), .A1(new_n13919_), .B0(pi0781), .Y(new_n13926_));
  OAI21X1  g11490(.A0(new_n13908_), .A1(new_n13907_), .B0(new_n11767_), .Y(new_n13927_));
  AOI21X1  g11491(.A0(new_n13927_), .A1(new_n13926_), .B0(pi0619), .Y(new_n13928_));
  MX2X1    g11492(.A(new_n13912_), .B(new_n13896_), .S0(new_n12513_), .Y(new_n13929_));
  INVX1    g11493(.A(new_n13929_), .Y(new_n13930_));
  OAI21X1  g11494(.A0(new_n13930_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13931_));
  OAI21X1  g11495(.A0(new_n13923_), .A1(new_n13917_), .B0(pi0781), .Y(new_n13932_));
  OAI21X1  g11496(.A0(new_n13915_), .A1(pi0781), .B0(new_n13932_), .Y(new_n13933_));
  AOI21X1  g11497(.A0(new_n13896_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n13934_));
  OAI21X1  g11498(.A0(new_n13933_), .A1(new_n12509_), .B0(new_n13934_), .Y(new_n13935_));
  AND2X1   g11499(.A(new_n13935_), .B(new_n12517_), .Y(new_n13936_));
  OAI21X1  g11500(.A0(new_n13931_), .A1(new_n13928_), .B0(new_n13936_), .Y(new_n13937_));
  AOI21X1  g11501(.A0(new_n13927_), .A1(new_n13926_), .B0(new_n12509_), .Y(new_n13938_));
  OAI21X1  g11502(.A0(new_n13930_), .A1(pi0619), .B0(pi1159), .Y(new_n13939_));
  AOI21X1  g11503(.A0(new_n13896_), .A1(pi0619), .B0(pi1159), .Y(new_n13940_));
  OAI21X1  g11504(.A0(new_n13933_), .A1(pi0619), .B0(new_n13940_), .Y(new_n13941_));
  AND2X1   g11505(.A(new_n13941_), .B(pi0648), .Y(new_n13942_));
  OAI21X1  g11506(.A0(new_n13939_), .A1(new_n13938_), .B0(new_n13942_), .Y(new_n13943_));
  AOI21X1  g11507(.A0(new_n13943_), .A1(new_n13937_), .B0(new_n11766_), .Y(new_n13944_));
  AOI21X1  g11508(.A0(new_n13927_), .A1(new_n13926_), .B0(pi0789), .Y(new_n13945_));
  OR3X1    g11509(.A(new_n13945_), .B(new_n13944_), .C(pi0788), .Y(new_n13946_));
  OR3X1    g11510(.A(new_n13945_), .B(new_n13944_), .C(pi0626), .Y(new_n13947_));
  MX2X1    g11511(.A(new_n13930_), .B(new_n13866_), .S0(new_n12531_), .Y(new_n13948_));
  AOI21X1  g11512(.A0(new_n13948_), .A1(pi0626), .B0(pi0641), .Y(new_n13949_));
  NAND2X1  g11513(.A(new_n13941_), .B(new_n13935_), .Y(new_n13950_));
  MX2X1    g11514(.A(new_n13950_), .B(new_n13933_), .S0(new_n11766_), .Y(new_n13951_));
  AOI21X1  g11515(.A0(new_n13896_), .A1(pi0626), .B0(pi1158), .Y(new_n13952_));
  OAI21X1  g11516(.A0(new_n13951_), .A1(pi0626), .B0(new_n13952_), .Y(new_n13953_));
  AOI22X1  g11517(.A0(new_n13953_), .A1(new_n13337_), .B0(new_n13949_), .B1(new_n13947_), .Y(new_n13954_));
  OR3X1    g11518(.A(new_n13945_), .B(new_n13944_), .C(new_n12542_), .Y(new_n13955_));
  AOI21X1  g11519(.A0(new_n13948_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n13956_));
  AOI21X1  g11520(.A0(new_n13896_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n13957_));
  OAI21X1  g11521(.A0(new_n13951_), .A1(new_n12542_), .B0(new_n13957_), .Y(new_n13958_));
  AOI22X1  g11522(.A0(new_n13958_), .A1(new_n13346_), .B0(new_n13956_), .B1(new_n13955_), .Y(new_n13959_));
  OAI21X1  g11523(.A0(new_n13959_), .A1(new_n13954_), .B0(pi0788), .Y(new_n13960_));
  AND3X1   g11524(.A(new_n13960_), .B(new_n13946_), .C(new_n12554_), .Y(new_n13961_));
  AOI21X1  g11525(.A0(new_n13958_), .A1(new_n13953_), .B0(new_n11765_), .Y(new_n13962_));
  AND2X1   g11526(.A(new_n13951_), .B(new_n11765_), .Y(new_n13963_));
  NOR2X1   g11527(.A(new_n13963_), .B(new_n13962_), .Y(new_n13964_));
  INVX1    g11528(.A(new_n13964_), .Y(new_n13965_));
  OAI21X1  g11529(.A0(new_n13965_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13966_));
  AND2X1   g11530(.A(new_n13866_), .B(new_n12563_), .Y(new_n13967_));
  AOI21X1  g11531(.A0(new_n13948_), .A1(new_n13356_), .B0(new_n13967_), .Y(new_n13968_));
  OAI21X1  g11532(.A0(new_n13866_), .A1(pi0628), .B0(pi1156), .Y(new_n13969_));
  AOI21X1  g11533(.A0(new_n13968_), .A1(pi0628), .B0(new_n13969_), .Y(new_n13970_));
  NOR2X1   g11534(.A(new_n13970_), .B(pi0629), .Y(new_n13971_));
  OAI21X1  g11535(.A0(new_n13966_), .A1(new_n13961_), .B0(new_n13971_), .Y(new_n13972_));
  AND3X1   g11536(.A(new_n13960_), .B(new_n13946_), .C(pi0628), .Y(new_n13973_));
  OAI21X1  g11537(.A0(new_n13965_), .A1(pi0628), .B0(pi1156), .Y(new_n13974_));
  OAI21X1  g11538(.A0(new_n13866_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n13975_));
  AOI21X1  g11539(.A0(new_n13968_), .A1(new_n12554_), .B0(new_n13975_), .Y(new_n13976_));
  NOR2X1   g11540(.A(new_n13976_), .B(new_n12561_), .Y(new_n13977_));
  OAI21X1  g11541(.A0(new_n13974_), .A1(new_n13973_), .B0(new_n13977_), .Y(new_n13978_));
  AOI21X1  g11542(.A0(new_n13978_), .A1(new_n13972_), .B0(new_n11764_), .Y(new_n13979_));
  AND3X1   g11543(.A(new_n13960_), .B(new_n13946_), .C(new_n11764_), .Y(new_n13980_));
  OAI21X1  g11544(.A0(new_n13980_), .A1(new_n13979_), .B0(new_n12577_), .Y(new_n13981_));
  MX2X1    g11545(.A(new_n13964_), .B(new_n13896_), .S0(new_n12580_), .Y(new_n13982_));
  AOI21X1  g11546(.A0(new_n13982_), .A1(pi0647), .B0(pi1157), .Y(new_n13983_));
  NOR2X1   g11547(.A(new_n13976_), .B(new_n13970_), .Y(new_n13984_));
  MX2X1    g11548(.A(new_n13984_), .B(new_n13968_), .S0(new_n11764_), .Y(new_n13985_));
  OAI21X1  g11549(.A0(new_n13866_), .A1(pi0647), .B0(pi1157), .Y(new_n13986_));
  AOI21X1  g11550(.A0(new_n13985_), .A1(pi0647), .B0(new_n13986_), .Y(new_n13987_));
  OR2X1    g11551(.A(new_n13987_), .B(pi0630), .Y(new_n13988_));
  AOI21X1  g11552(.A0(new_n13983_), .A1(new_n13981_), .B0(new_n13988_), .Y(new_n13989_));
  OAI21X1  g11553(.A0(new_n13980_), .A1(new_n13979_), .B0(pi0647), .Y(new_n13990_));
  AOI21X1  g11554(.A0(new_n13982_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13991_));
  OAI21X1  g11555(.A0(new_n13866_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n13992_));
  AOI21X1  g11556(.A0(new_n13985_), .A1(new_n12577_), .B0(new_n13992_), .Y(new_n13993_));
  OR2X1    g11557(.A(new_n13993_), .B(new_n12592_), .Y(new_n13994_));
  AOI21X1  g11558(.A0(new_n13991_), .A1(new_n13990_), .B0(new_n13994_), .Y(new_n13995_));
  OAI21X1  g11559(.A0(new_n13995_), .A1(new_n13989_), .B0(pi0787), .Y(new_n13996_));
  OAI21X1  g11560(.A0(new_n13980_), .A1(new_n13979_), .B0(new_n11763_), .Y(new_n13997_));
  AOI21X1  g11561(.A0(new_n13997_), .A1(new_n13996_), .B0(new_n12612_), .Y(new_n13998_));
  OAI21X1  g11562(.A0(new_n13993_), .A1(new_n13987_), .B0(pi0787), .Y(new_n13999_));
  OAI21X1  g11563(.A0(new_n13985_), .A1(pi0787), .B0(new_n13999_), .Y(new_n14000_));
  OAI21X1  g11564(.A0(new_n14000_), .A1(pi0644), .B0(pi0715), .Y(new_n14001_));
  NOR2X1   g11565(.A(new_n13866_), .B(new_n12605_), .Y(new_n14002_));
  AOI21X1  g11566(.A0(new_n13982_), .A1(new_n12605_), .B0(new_n14002_), .Y(new_n14003_));
  AOI21X1  g11567(.A0(new_n13896_), .A1(new_n12612_), .B0(pi0715), .Y(new_n14004_));
  OAI21X1  g11568(.A0(new_n14003_), .A1(new_n12612_), .B0(new_n14004_), .Y(new_n14005_));
  AND2X1   g11569(.A(new_n14005_), .B(pi1160), .Y(new_n14006_));
  OAI21X1  g11570(.A0(new_n14001_), .A1(new_n13998_), .B0(new_n14006_), .Y(new_n14007_));
  AOI21X1  g11571(.A0(new_n13997_), .A1(new_n13996_), .B0(pi0644), .Y(new_n14008_));
  OAI21X1  g11572(.A0(new_n14000_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n14009_));
  AOI21X1  g11573(.A0(new_n13896_), .A1(pi0644), .B0(new_n12608_), .Y(new_n14010_));
  OAI21X1  g11574(.A0(new_n14003_), .A1(pi0644), .B0(new_n14010_), .Y(new_n14011_));
  AND2X1   g11575(.A(new_n14011_), .B(new_n11762_), .Y(new_n14012_));
  OAI21X1  g11576(.A0(new_n14009_), .A1(new_n14008_), .B0(new_n14012_), .Y(new_n14013_));
  AND3X1   g11577(.A(new_n14013_), .B(new_n14007_), .C(pi0790), .Y(new_n14014_));
  AND3X1   g11578(.A(new_n13997_), .B(new_n13996_), .C(new_n12766_), .Y(new_n14015_));
  OR2X1    g11579(.A(new_n14015_), .B(new_n5103_), .Y(new_n14016_));
  AOI21X1  g11580(.A0(new_n5103_), .A1(new_n7344_), .B0(pi0057), .Y(new_n14017_));
  OAI21X1  g11581(.A0(new_n14016_), .A1(new_n14014_), .B0(new_n14017_), .Y(new_n14018_));
  AOI21X1  g11582(.A0(pi0144), .A1(pi0057), .B0(pi0832), .Y(new_n14019_));
  NOR2X1   g11583(.A(new_n2720_), .B(new_n7344_), .Y(new_n14020_));
  AOI21X1  g11584(.A0(new_n12439_), .A1(pi0736), .B0(new_n14020_), .Y(new_n14021_));
  NAND2X1  g11585(.A(new_n14021_), .B(new_n11769_), .Y(new_n14022_));
  AND3X1   g11586(.A(new_n12439_), .B(pi0736), .C(pi0625), .Y(new_n14023_));
  OAI21X1  g11587(.A0(new_n14023_), .A1(new_n14021_), .B0(new_n12364_), .Y(new_n14024_));
  INVX1    g11588(.A(new_n14024_), .Y(new_n14025_));
  NOR3X1   g11589(.A(new_n14023_), .B(new_n14020_), .C(new_n12364_), .Y(new_n14026_));
  OAI21X1  g11590(.A0(new_n14026_), .A1(new_n14025_), .B0(pi0778), .Y(new_n14027_));
  AND2X1   g11591(.A(new_n14027_), .B(new_n14022_), .Y(new_n14028_));
  INVX1    g11592(.A(new_n14028_), .Y(new_n14029_));
  NOR2X1   g11593(.A(new_n14029_), .B(new_n13489_), .Y(new_n14030_));
  AOI21X1  g11594(.A0(new_n14030_), .A1(new_n12554_), .B0(new_n12561_), .Y(new_n14031_));
  NOR2X1   g11595(.A(pi1155), .B(pi0609), .Y(new_n14032_));
  AND2X1   g11596(.A(pi1155), .B(pi0609), .Y(new_n14033_));
  NOR3X1   g11597(.A(new_n14033_), .B(new_n14032_), .C(new_n11768_), .Y(new_n14034_));
  XOR2X1   g11598(.A(pi1159), .B(pi0619), .Y(new_n14035_));
  AND2X1   g11599(.A(new_n14035_), .B(pi0789), .Y(new_n14036_));
  NOR2X1   g11600(.A(pi1154), .B(pi0618), .Y(new_n14037_));
  AND2X1   g11601(.A(pi1154), .B(pi0618), .Y(new_n14038_));
  NOR3X1   g11602(.A(new_n14038_), .B(new_n14037_), .C(new_n11767_), .Y(new_n14039_));
  OR3X1    g11603(.A(new_n14039_), .B(new_n14036_), .C(new_n12473_), .Y(new_n14040_));
  OR4X1    g11604(.A(new_n14040_), .B(new_n14034_), .C(new_n12057_), .D(new_n13836_), .Y(new_n14041_));
  NOR2X1   g11605(.A(new_n14041_), .B(new_n12708_), .Y(new_n14042_));
  NOR2X1   g11606(.A(new_n14042_), .B(new_n12554_), .Y(new_n14043_));
  OAI21X1  g11607(.A0(new_n14043_), .A1(new_n14031_), .B0(new_n12555_), .Y(new_n14044_));
  OR3X1    g11608(.A(new_n14029_), .B(new_n13489_), .C(new_n12554_), .Y(new_n14045_));
  OAI21X1  g11609(.A0(new_n14042_), .A1(pi0628), .B0(pi0629), .Y(new_n14046_));
  NAND3X1  g11610(.A(new_n14046_), .B(new_n14045_), .C(pi1156), .Y(new_n14047_));
  AOI21X1  g11611(.A0(new_n14047_), .A1(new_n14044_), .B0(new_n14020_), .Y(new_n14048_));
  AND2X1   g11612(.A(pi1158), .B(new_n12542_), .Y(new_n14049_));
  INVX1    g11613(.A(new_n14049_), .Y(new_n14050_));
  INVX1    g11614(.A(new_n12531_), .Y(new_n14051_));
  INVX1    g11615(.A(new_n14020_), .Y(new_n14052_));
  INVX1    g11616(.A(new_n12513_), .Y(new_n14053_));
  NAND4X1  g11617(.A(new_n14027_), .B(new_n14022_), .C(new_n14053_), .D(new_n13910_), .Y(new_n14054_));
  AND2X1   g11618(.A(new_n14054_), .B(new_n14052_), .Y(new_n14055_));
  INVX1    g11619(.A(new_n14055_), .Y(new_n14056_));
  OAI21X1  g11620(.A0(new_n14020_), .A1(new_n14051_), .B0(new_n14056_), .Y(new_n14057_));
  OAI21X1  g11621(.A0(new_n14041_), .A1(pi0626), .B0(new_n14052_), .Y(new_n14058_));
  AOI21X1  g11622(.A0(new_n14058_), .A1(new_n12548_), .B0(new_n12543_), .Y(new_n14059_));
  OAI21X1  g11623(.A0(new_n14057_), .A1(new_n14050_), .B0(new_n14059_), .Y(new_n14060_));
  AND2X1   g11624(.A(new_n12548_), .B(pi0626), .Y(new_n14061_));
  INVX1    g11625(.A(new_n14061_), .Y(new_n14062_));
  OAI21X1  g11626(.A0(new_n14041_), .A1(new_n12542_), .B0(new_n14052_), .Y(new_n14063_));
  AOI21X1  g11627(.A0(new_n14063_), .A1(pi1158), .B0(pi0641), .Y(new_n14064_));
  OAI21X1  g11628(.A0(new_n14057_), .A1(new_n14062_), .B0(new_n14064_), .Y(new_n14065_));
  AND3X1   g11629(.A(new_n14065_), .B(new_n14060_), .C(pi0788), .Y(new_n14066_));
  INVX1    g11630(.A(new_n14066_), .Y(new_n14067_));
  INVX1    g11631(.A(new_n13443_), .Y(new_n14068_));
  AOI21X1  g11632(.A0(new_n12056_), .A1(pi0758), .B0(new_n14020_), .Y(new_n14069_));
  OAI21X1  g11633(.A0(new_n14068_), .A1(new_n13832_), .B0(new_n14069_), .Y(new_n14070_));
  NAND3X1  g11634(.A(new_n13443_), .B(pi0736), .C(pi0625), .Y(new_n14071_));
  AOI21X1  g11635(.A0(new_n14071_), .A1(new_n14070_), .B0(pi1153), .Y(new_n14072_));
  NOR3X1   g11636(.A(new_n14072_), .B(new_n14026_), .C(pi0608), .Y(new_n14073_));
  AND3X1   g11637(.A(new_n14071_), .B(new_n14069_), .C(pi1153), .Y(new_n14074_));
  NOR3X1   g11638(.A(new_n14074_), .B(new_n14025_), .C(new_n12368_), .Y(new_n14075_));
  OR2X1    g11639(.A(new_n14075_), .B(new_n14073_), .Y(new_n14076_));
  MX2X1    g11640(.A(new_n14076_), .B(new_n14070_), .S0(new_n11769_), .Y(new_n14077_));
  INVX1    g11641(.A(new_n14077_), .Y(new_n14078_));
  AOI21X1  g11642(.A0(new_n14028_), .A1(pi0609), .B0(pi1155), .Y(new_n14079_));
  OAI21X1  g11643(.A0(new_n14078_), .A1(pi0609), .B0(new_n14079_), .Y(new_n14080_));
  NAND3X1  g11644(.A(new_n12471_), .B(new_n12056_), .C(pi0758), .Y(new_n14081_));
  NOR2X1   g11645(.A(new_n14020_), .B(new_n12463_), .Y(new_n14082_));
  AOI21X1  g11646(.A0(new_n14082_), .A1(new_n14081_), .B0(pi0660), .Y(new_n14083_));
  AOI21X1  g11647(.A0(new_n14028_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n14084_));
  OAI21X1  g11648(.A0(new_n14078_), .A1(new_n12462_), .B0(new_n14084_), .Y(new_n14085_));
  NAND3X1  g11649(.A(new_n12480_), .B(new_n12056_), .C(pi0758), .Y(new_n14086_));
  NOR2X1   g11650(.A(new_n14020_), .B(pi1155), .Y(new_n14087_));
  AOI21X1  g11651(.A0(new_n14087_), .A1(new_n14086_), .B0(new_n12468_), .Y(new_n14088_));
  AOI22X1  g11652(.A0(new_n14088_), .A1(new_n14085_), .B0(new_n14083_), .B1(new_n14080_), .Y(new_n14089_));
  MX2X1    g11653(.A(new_n14089_), .B(new_n14078_), .S0(new_n11768_), .Y(new_n14090_));
  AOI21X1  g11654(.A0(new_n14028_), .A1(new_n13910_), .B0(new_n14020_), .Y(new_n14091_));
  INVX1    g11655(.A(new_n14091_), .Y(new_n14092_));
  AOI21X1  g11656(.A0(new_n14092_), .A1(pi0618), .B0(pi1154), .Y(new_n14093_));
  OAI21X1  g11657(.A0(new_n14090_), .A1(pi0618), .B0(new_n14093_), .Y(new_n14094_));
  OR3X1    g11658(.A(new_n14034_), .B(new_n12057_), .C(new_n13836_), .Y(new_n14095_));
  NOR3X1   g11659(.A(new_n14095_), .B(new_n12473_), .C(new_n12486_), .Y(new_n14096_));
  OR3X1    g11660(.A(new_n14096_), .B(new_n14020_), .C(new_n12487_), .Y(new_n14097_));
  AND2X1   g11661(.A(new_n14097_), .B(new_n12494_), .Y(new_n14098_));
  AOI21X1  g11662(.A0(new_n14092_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n14099_));
  OAI21X1  g11663(.A0(new_n14090_), .A1(new_n12486_), .B0(new_n14099_), .Y(new_n14100_));
  NOR3X1   g11664(.A(new_n14095_), .B(new_n12473_), .C(pi0618), .Y(new_n14101_));
  OR3X1    g11665(.A(new_n14101_), .B(new_n14020_), .C(pi1154), .Y(new_n14102_));
  AND2X1   g11666(.A(new_n14102_), .B(pi0627), .Y(new_n14103_));
  AOI22X1  g11667(.A0(new_n14103_), .A1(new_n14100_), .B0(new_n14098_), .B1(new_n14094_), .Y(new_n14104_));
  MX2X1    g11668(.A(new_n14104_), .B(new_n14090_), .S0(new_n11767_), .Y(new_n14105_));
  AOI21X1  g11669(.A0(new_n14056_), .A1(pi0619), .B0(pi1159), .Y(new_n14106_));
  OAI21X1  g11670(.A0(new_n14105_), .A1(pi0619), .B0(new_n14106_), .Y(new_n14107_));
  NOR4X1   g11671(.A(new_n14039_), .B(new_n14095_), .C(new_n12473_), .D(new_n12509_), .Y(new_n14108_));
  OR3X1    g11672(.A(new_n14108_), .B(new_n14020_), .C(new_n12510_), .Y(new_n14109_));
  AND3X1   g11673(.A(new_n14109_), .B(new_n14107_), .C(new_n12517_), .Y(new_n14110_));
  AOI21X1  g11674(.A0(new_n14056_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n14111_));
  OAI21X1  g11675(.A0(new_n14105_), .A1(new_n12509_), .B0(new_n14111_), .Y(new_n14112_));
  NOR4X1   g11676(.A(new_n14039_), .B(new_n14095_), .C(new_n12473_), .D(pi0619), .Y(new_n14113_));
  OR3X1    g11677(.A(new_n14113_), .B(new_n14020_), .C(pi1159), .Y(new_n14114_));
  AND2X1   g11678(.A(new_n14114_), .B(pi0648), .Y(new_n14115_));
  AOI21X1  g11679(.A0(new_n14115_), .A1(new_n14112_), .B0(new_n11766_), .Y(new_n14116_));
  INVX1    g11680(.A(new_n14116_), .Y(new_n14117_));
  AOI21X1  g11681(.A0(new_n14105_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n14118_));
  OAI21X1  g11682(.A0(new_n14117_), .A1(new_n14110_), .B0(new_n14118_), .Y(new_n14119_));
  AOI22X1  g11683(.A0(new_n14119_), .A1(new_n14067_), .B0(new_n14048_), .B1(pi0792), .Y(new_n14120_));
  AOI21X1  g11684(.A0(new_n13519_), .A1(new_n12603_), .B0(new_n11763_), .Y(new_n14121_));
  INVX1    g11685(.A(new_n14121_), .Y(new_n14122_));
  AND3X1   g11686(.A(pi1156), .B(pi0629), .C(pi0628), .Y(new_n14123_));
  NOR3X1   g11687(.A(pi1156), .B(pi0629), .C(pi0628), .Y(new_n14124_));
  NOR3X1   g11688(.A(new_n14124_), .B(new_n14123_), .C(new_n11764_), .Y(new_n14125_));
  INVX1    g11689(.A(new_n14125_), .Y(new_n14126_));
  OAI21X1  g11690(.A0(new_n14126_), .A1(new_n14048_), .B0(new_n14122_), .Y(new_n14127_));
  OR2X1    g11691(.A(new_n14127_), .B(new_n14120_), .Y(new_n14128_));
  NOR3X1   g11692(.A(new_n14041_), .B(new_n12708_), .C(new_n12580_), .Y(new_n14129_));
  AOI21X1  g11693(.A0(new_n14129_), .A1(new_n12592_), .B0(new_n12577_), .Y(new_n14130_));
  NOR3X1   g11694(.A(new_n14029_), .B(new_n13508_), .C(new_n13489_), .Y(new_n14131_));
  INVX1    g11695(.A(new_n14131_), .Y(new_n14132_));
  AOI21X1  g11696(.A0(new_n14132_), .A1(pi0630), .B0(new_n14130_), .Y(new_n14133_));
  AOI21X1  g11697(.A0(new_n14132_), .A1(new_n12592_), .B0(new_n12577_), .Y(new_n14134_));
  AOI21X1  g11698(.A0(new_n14129_), .A1(pi0630), .B0(new_n12578_), .Y(new_n14135_));
  INVX1    g11699(.A(new_n14135_), .Y(new_n14136_));
  OAI22X1  g11700(.A0(new_n14136_), .A1(new_n14134_), .B0(new_n14133_), .B1(pi1157), .Y(new_n14137_));
  NAND3X1  g11701(.A(new_n14137_), .B(new_n14052_), .C(pi0787), .Y(new_n14138_));
  AND2X1   g11702(.A(new_n14138_), .B(new_n14128_), .Y(new_n14139_));
  INVX1    g11703(.A(new_n13520_), .Y(new_n14140_));
  AOI21X1  g11704(.A0(new_n14131_), .A1(new_n14140_), .B0(new_n14020_), .Y(new_n14141_));
  OAI21X1  g11705(.A0(new_n14141_), .A1(pi0644), .B0(pi0715), .Y(new_n14142_));
  AOI21X1  g11706(.A0(new_n14139_), .A1(pi0644), .B0(new_n14142_), .Y(new_n14143_));
  AND3X1   g11707(.A(new_n14129_), .B(new_n12605_), .C(pi0644), .Y(new_n14144_));
  OAI21X1  g11708(.A0(new_n2720_), .A1(new_n7344_), .B0(new_n12608_), .Y(new_n14145_));
  OAI21X1  g11709(.A0(new_n14145_), .A1(new_n14144_), .B0(pi1160), .Y(new_n14146_));
  OAI21X1  g11710(.A0(new_n14141_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n14147_));
  AOI21X1  g11711(.A0(new_n14139_), .A1(new_n12612_), .B0(new_n14147_), .Y(new_n14148_));
  AND3X1   g11712(.A(new_n14129_), .B(new_n12605_), .C(new_n12612_), .Y(new_n14149_));
  OAI21X1  g11713(.A0(new_n2720_), .A1(new_n7344_), .B0(pi0715), .Y(new_n14150_));
  OAI21X1  g11714(.A0(new_n14150_), .A1(new_n14149_), .B0(new_n11762_), .Y(new_n14151_));
  OAI22X1  g11715(.A0(new_n14151_), .A1(new_n14148_), .B0(new_n14146_), .B1(new_n14143_), .Y(new_n14152_));
  AND3X1   g11716(.A(new_n14138_), .B(new_n14128_), .C(new_n12766_), .Y(new_n14153_));
  OR2X1    g11717(.A(new_n14153_), .B(new_n12767_), .Y(new_n14154_));
  AOI21X1  g11718(.A0(new_n14152_), .A1(pi0790), .B0(new_n14154_), .Y(new_n14155_));
  AOI21X1  g11719(.A0(new_n14019_), .A1(new_n14018_), .B0(new_n14155_), .Y(po0301));
  AOI21X1  g11720(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0145), .Y(new_n14157_));
  INVX1    g11721(.A(new_n14157_), .Y(new_n14158_));
  OAI21X1  g11722(.A0(new_n11770_), .A1(pi0698), .B0(new_n14157_), .Y(new_n14159_));
  OAI21X1  g11723(.A0(new_n12826_), .A1(new_n5202_), .B0(new_n2979_), .Y(new_n14160_));
  AOI22X1  g11724(.A0(new_n14160_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n5202_), .Y(new_n14161_));
  AOI21X1  g11725(.A0(new_n12771_), .A1(new_n5202_), .B0(new_n12441_), .Y(new_n14162_));
  OR3X1    g11726(.A(new_n14162_), .B(new_n14161_), .C(pi0698), .Y(new_n14163_));
  NAND3X1  g11727(.A(new_n14163_), .B(new_n14159_), .C(new_n11769_), .Y(new_n14164_));
  AOI21X1  g11728(.A0(new_n14163_), .A1(new_n14159_), .B0(new_n12363_), .Y(new_n14165_));
  OAI21X1  g11729(.A0(new_n14158_), .A1(pi0625), .B0(pi1153), .Y(new_n14166_));
  NOR2X1   g11730(.A(new_n14166_), .B(new_n14165_), .Y(new_n14167_));
  AOI21X1  g11731(.A0(new_n14163_), .A1(new_n14159_), .B0(pi0625), .Y(new_n14168_));
  OAI21X1  g11732(.A0(new_n14158_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n14169_));
  NOR2X1   g11733(.A(new_n14169_), .B(new_n14168_), .Y(new_n14170_));
  OAI21X1  g11734(.A0(new_n14170_), .A1(new_n14167_), .B0(pi0778), .Y(new_n14171_));
  AND2X1   g11735(.A(new_n14171_), .B(new_n14164_), .Y(new_n14172_));
  MX2X1    g11736(.A(new_n14172_), .B(new_n14157_), .S0(new_n12490_), .Y(new_n14173_));
  INVX1    g11737(.A(new_n14173_), .Y(new_n14174_));
  MX2X1    g11738(.A(new_n14174_), .B(new_n14158_), .S0(new_n12513_), .Y(new_n14175_));
  INVX1    g11739(.A(new_n14175_), .Y(new_n14176_));
  MX2X1    g11740(.A(new_n14176_), .B(new_n14157_), .S0(new_n12531_), .Y(new_n14177_));
  INVX1    g11741(.A(new_n14177_), .Y(new_n14178_));
  MX2X1    g11742(.A(new_n14178_), .B(new_n14158_), .S0(new_n12563_), .Y(new_n14179_));
  AOI21X1  g11743(.A0(new_n14157_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n14180_));
  OAI21X1  g11744(.A0(new_n14179_), .A1(new_n12554_), .B0(new_n14180_), .Y(new_n14181_));
  AOI21X1  g11745(.A0(new_n14157_), .A1(pi0628), .B0(pi1156), .Y(new_n14182_));
  OAI21X1  g11746(.A0(new_n14179_), .A1(pi0628), .B0(new_n14182_), .Y(new_n14183_));
  AOI21X1  g11747(.A0(new_n14183_), .A1(new_n14181_), .B0(new_n11764_), .Y(new_n14184_));
  AOI21X1  g11748(.A0(new_n14179_), .A1(new_n11764_), .B0(new_n14184_), .Y(new_n14185_));
  MX2X1    g11749(.A(new_n14185_), .B(new_n14157_), .S0(pi0647), .Y(new_n14186_));
  MX2X1    g11750(.A(new_n14185_), .B(new_n14157_), .S0(new_n12577_), .Y(new_n14187_));
  MX2X1    g11751(.A(new_n14187_), .B(new_n14186_), .S0(new_n12578_), .Y(new_n14188_));
  MX2X1    g11752(.A(new_n14188_), .B(new_n14185_), .S0(new_n11763_), .Y(new_n14189_));
  AOI21X1  g11753(.A0(new_n14189_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n14190_));
  INVX1    g11754(.A(pi0767), .Y(new_n14191_));
  AOI21X1  g11755(.A0(new_n11959_), .A1(new_n5202_), .B0(new_n14191_), .Y(new_n14192_));
  NOR2X1   g11756(.A(pi0767), .B(pi0145), .Y(new_n14193_));
  INVX1    g11757(.A(new_n14193_), .Y(new_n14194_));
  OAI22X1  g11758(.A0(new_n14194_), .A1(new_n12776_), .B0(new_n12074_), .B1(new_n5202_), .Y(new_n14195_));
  OAI21X1  g11759(.A0(new_n14195_), .A1(new_n14192_), .B0(new_n2979_), .Y(new_n14196_));
  INVX1    g11760(.A(new_n12079_), .Y(new_n14197_));
  AOI21X1  g11761(.A0(new_n12771_), .A1(new_n5202_), .B0(new_n2979_), .Y(new_n14198_));
  OAI21X1  g11762(.A0(new_n14197_), .A1(pi0767), .B0(new_n14198_), .Y(new_n14199_));
  NAND2X1  g11763(.A(new_n14199_), .B(new_n14196_), .Y(new_n14200_));
  MX2X1    g11764(.A(new_n14200_), .B(pi0145), .S0(new_n11770_), .Y(new_n14201_));
  AND2X1   g11765(.A(new_n14201_), .B(new_n12474_), .Y(new_n14202_));
  AOI21X1  g11766(.A0(new_n14158_), .A1(new_n12473_), .B0(new_n14202_), .Y(new_n14203_));
  AOI22X1  g11767(.A0(new_n14202_), .A1(pi0609), .B0(new_n14158_), .B1(new_n12472_), .Y(new_n14204_));
  NOR2X1   g11768(.A(new_n14204_), .B(new_n12463_), .Y(new_n14205_));
  AOI22X1  g11769(.A0(new_n14202_), .A1(new_n12462_), .B0(new_n14158_), .B1(new_n12481_), .Y(new_n14206_));
  NOR2X1   g11770(.A(new_n14206_), .B(pi1155), .Y(new_n14207_));
  OAI21X1  g11771(.A0(new_n14207_), .A1(new_n14205_), .B0(pi0785), .Y(new_n14208_));
  OAI21X1  g11772(.A0(new_n14203_), .A1(pi0785), .B0(new_n14208_), .Y(new_n14209_));
  AOI21X1  g11773(.A0(new_n14157_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n14210_));
  OAI21X1  g11774(.A0(new_n14209_), .A1(new_n12486_), .B0(new_n14210_), .Y(new_n14211_));
  AOI21X1  g11775(.A0(new_n14157_), .A1(pi0618), .B0(pi1154), .Y(new_n14212_));
  OAI21X1  g11776(.A0(new_n14209_), .A1(pi0618), .B0(new_n14212_), .Y(new_n14213_));
  NAND2X1  g11777(.A(new_n14213_), .B(new_n14211_), .Y(new_n14214_));
  MX2X1    g11778(.A(new_n14214_), .B(new_n14209_), .S0(new_n11767_), .Y(new_n14215_));
  AND2X1   g11779(.A(new_n14215_), .B(new_n11766_), .Y(new_n14216_));
  AOI21X1  g11780(.A0(new_n14157_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n14217_));
  OAI21X1  g11781(.A0(new_n14215_), .A1(new_n12509_), .B0(new_n14217_), .Y(new_n14218_));
  AOI21X1  g11782(.A0(new_n14157_), .A1(pi0619), .B0(pi1159), .Y(new_n14219_));
  OAI21X1  g11783(.A0(new_n14215_), .A1(pi0619), .B0(new_n14219_), .Y(new_n14220_));
  AOI21X1  g11784(.A0(new_n14220_), .A1(new_n14218_), .B0(new_n11766_), .Y(new_n14221_));
  OR2X1    g11785(.A(new_n14221_), .B(new_n14216_), .Y(new_n14222_));
  AND2X1   g11786(.A(new_n14222_), .B(new_n11765_), .Y(new_n14223_));
  NOR3X1   g11787(.A(new_n14221_), .B(new_n14216_), .C(new_n12542_), .Y(new_n14224_));
  AOI21X1  g11788(.A0(new_n14157_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n14225_));
  INVX1    g11789(.A(new_n14225_), .Y(new_n14226_));
  NOR3X1   g11790(.A(new_n14221_), .B(new_n14216_), .C(pi0626), .Y(new_n14227_));
  AOI21X1  g11791(.A0(new_n14157_), .A1(pi0626), .B0(pi1158), .Y(new_n14228_));
  INVX1    g11792(.A(new_n14228_), .Y(new_n14229_));
  OAI22X1  g11793(.A0(new_n14229_), .A1(new_n14227_), .B0(new_n14226_), .B1(new_n14224_), .Y(new_n14230_));
  AOI21X1  g11794(.A0(new_n14230_), .A1(pi0788), .B0(new_n14223_), .Y(new_n14231_));
  MX2X1    g11795(.A(new_n14231_), .B(new_n14157_), .S0(new_n12580_), .Y(new_n14232_));
  MX2X1    g11796(.A(new_n14232_), .B(new_n14157_), .S0(new_n12604_), .Y(new_n14233_));
  OAI21X1  g11797(.A0(new_n14158_), .A1(pi0644), .B0(new_n12608_), .Y(new_n14234_));
  AOI21X1  g11798(.A0(new_n14233_), .A1(pi0644), .B0(new_n14234_), .Y(new_n14235_));
  OR3X1    g11799(.A(new_n14235_), .B(new_n14190_), .C(new_n11762_), .Y(new_n14236_));
  AND3X1   g11800(.A(pi1157), .B(new_n12577_), .C(pi0630), .Y(new_n14237_));
  AND3X1   g11801(.A(new_n12578_), .B(pi0647), .C(new_n12592_), .Y(new_n14238_));
  NOR2X1   g11802(.A(new_n14238_), .B(new_n14237_), .Y(new_n14239_));
  NOR2X1   g11803(.A(new_n14239_), .B(new_n14232_), .Y(new_n14240_));
  AND2X1   g11804(.A(pi1157), .B(new_n12592_), .Y(new_n14241_));
  INVX1    g11805(.A(new_n14241_), .Y(new_n14242_));
  AND2X1   g11806(.A(new_n12578_), .B(pi0630), .Y(new_n14243_));
  INVX1    g11807(.A(new_n14243_), .Y(new_n14244_));
  OAI22X1  g11808(.A0(new_n14187_), .A1(new_n14242_), .B0(new_n14186_), .B1(new_n14244_), .Y(new_n14245_));
  OAI21X1  g11809(.A0(new_n14245_), .A1(new_n14240_), .B0(pi0787), .Y(new_n14246_));
  AND2X1   g11810(.A(pi0629), .B(new_n12554_), .Y(new_n14247_));
  AND2X1   g11811(.A(new_n12561_), .B(pi0628), .Y(new_n14248_));
  MX2X1    g11812(.A(new_n14248_), .B(new_n14247_), .S0(pi1156), .Y(new_n14249_));
  INVX1    g11813(.A(new_n14249_), .Y(new_n14250_));
  MX2X1    g11814(.A(new_n14183_), .B(new_n14181_), .S0(new_n12561_), .Y(new_n14251_));
  OAI21X1  g11815(.A0(new_n14250_), .A1(new_n14231_), .B0(new_n14251_), .Y(new_n14252_));
  NAND3X1  g11816(.A(new_n14199_), .B(new_n14196_), .C(pi0698), .Y(new_n14253_));
  OAI21X1  g11817(.A0(new_n12213_), .A1(new_n5202_), .B0(pi0767), .Y(new_n14254_));
  AOI21X1  g11818(.A0(new_n12155_), .A1(new_n5202_), .B0(new_n14254_), .Y(new_n14255_));
  AOI21X1  g11819(.A0(new_n12788_), .A1(new_n5202_), .B0(pi0767), .Y(new_n14256_));
  OAI21X1  g11820(.A0(new_n12787_), .A1(new_n5202_), .B0(new_n14256_), .Y(new_n14257_));
  NAND2X1  g11821(.A(new_n14257_), .B(pi0039), .Y(new_n14258_));
  AND2X1   g11822(.A(new_n12332_), .B(pi0145), .Y(new_n14259_));
  OAI21X1  g11823(.A0(new_n12315_), .A1(pi0145), .B0(pi0767), .Y(new_n14260_));
  NOR4X1   g11824(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0145), .Y(new_n14261_));
  OAI21X1  g11825(.A0(new_n12800_), .A1(new_n5202_), .B0(new_n14191_), .Y(new_n14262_));
  OAI22X1  g11826(.A0(new_n14262_), .A1(new_n14261_), .B0(new_n14260_), .B1(new_n14259_), .Y(new_n14263_));
  AOI21X1  g11827(.A0(new_n14263_), .A1(new_n2939_), .B0(pi0038), .Y(new_n14264_));
  OAI21X1  g11828(.A0(new_n14258_), .A1(new_n14255_), .B0(new_n14264_), .Y(new_n14265_));
  OAI21X1  g11829(.A0(new_n12276_), .A1(pi0767), .B0(new_n13540_), .Y(new_n14266_));
  NAND2X1  g11830(.A(new_n14266_), .B(new_n5202_), .Y(new_n14267_));
  AOI21X1  g11831(.A0(new_n12056_), .A1(new_n14191_), .B0(new_n13443_), .Y(new_n14268_));
  NOR2X1   g11832(.A(new_n14268_), .B(new_n5202_), .Y(new_n14269_));
  AOI21X1  g11833(.A0(new_n14269_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n14270_));
  AOI21X1  g11834(.A0(new_n14270_), .A1(new_n14267_), .B0(pi0698), .Y(new_n14271_));
  AOI21X1  g11835(.A0(new_n14271_), .A1(new_n14265_), .B0(new_n11770_), .Y(new_n14272_));
  AOI22X1  g11836(.A0(new_n14272_), .A1(new_n14253_), .B0(new_n11770_), .B1(pi0145), .Y(new_n14273_));
  OAI21X1  g11837(.A0(new_n14201_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n14274_));
  AOI21X1  g11838(.A0(new_n14273_), .A1(new_n12363_), .B0(new_n14274_), .Y(new_n14275_));
  OR3X1    g11839(.A(new_n14275_), .B(new_n14167_), .C(pi0608), .Y(new_n14276_));
  OAI21X1  g11840(.A0(new_n14201_), .A1(pi0625), .B0(pi1153), .Y(new_n14277_));
  AOI21X1  g11841(.A0(new_n14273_), .A1(pi0625), .B0(new_n14277_), .Y(new_n14278_));
  OR3X1    g11842(.A(new_n14278_), .B(new_n14170_), .C(new_n12368_), .Y(new_n14279_));
  AOI21X1  g11843(.A0(new_n14279_), .A1(new_n14276_), .B0(new_n11769_), .Y(new_n14280_));
  AOI21X1  g11844(.A0(new_n14273_), .A1(new_n11769_), .B0(new_n14280_), .Y(new_n14281_));
  AOI21X1  g11845(.A0(new_n14172_), .A1(pi0609), .B0(pi1155), .Y(new_n14282_));
  OAI21X1  g11846(.A0(new_n14281_), .A1(pi0609), .B0(new_n14282_), .Y(new_n14283_));
  NOR2X1   g11847(.A(new_n14205_), .B(pi0660), .Y(new_n14284_));
  AOI21X1  g11848(.A0(new_n14172_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n14285_));
  OAI21X1  g11849(.A0(new_n14281_), .A1(new_n12462_), .B0(new_n14285_), .Y(new_n14286_));
  NOR2X1   g11850(.A(new_n14207_), .B(new_n12468_), .Y(new_n14287_));
  AOI22X1  g11851(.A0(new_n14287_), .A1(new_n14286_), .B0(new_n14284_), .B1(new_n14283_), .Y(new_n14288_));
  OR2X1    g11852(.A(new_n14281_), .B(pi0785), .Y(new_n14289_));
  OAI21X1  g11853(.A0(new_n14288_), .A1(new_n11768_), .B0(new_n14289_), .Y(new_n14290_));
  OAI21X1  g11854(.A0(new_n14174_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n14291_));
  AOI21X1  g11855(.A0(new_n14290_), .A1(new_n12486_), .B0(new_n14291_), .Y(new_n14292_));
  NAND2X1  g11856(.A(new_n14211_), .B(new_n12494_), .Y(new_n14293_));
  OAI21X1  g11857(.A0(new_n14174_), .A1(pi0618), .B0(pi1154), .Y(new_n14294_));
  AOI21X1  g11858(.A0(new_n14290_), .A1(pi0618), .B0(new_n14294_), .Y(new_n14295_));
  NAND2X1  g11859(.A(new_n14213_), .B(pi0627), .Y(new_n14296_));
  OAI22X1  g11860(.A0(new_n14296_), .A1(new_n14295_), .B0(new_n14293_), .B1(new_n14292_), .Y(new_n14297_));
  MX2X1    g11861(.A(new_n14297_), .B(new_n14290_), .S0(new_n11767_), .Y(new_n14298_));
  NAND2X1  g11862(.A(new_n14298_), .B(new_n12509_), .Y(new_n14299_));
  AOI21X1  g11863(.A0(new_n14176_), .A1(pi0619), .B0(pi1159), .Y(new_n14300_));
  NAND2X1  g11864(.A(new_n14218_), .B(new_n12517_), .Y(new_n14301_));
  AOI21X1  g11865(.A0(new_n14300_), .A1(new_n14299_), .B0(new_n14301_), .Y(new_n14302_));
  NAND2X1  g11866(.A(new_n14298_), .B(pi0619), .Y(new_n14303_));
  AOI21X1  g11867(.A0(new_n14176_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n14304_));
  NAND2X1  g11868(.A(new_n14220_), .B(pi0648), .Y(new_n14305_));
  AOI21X1  g11869(.A0(new_n14304_), .A1(new_n14303_), .B0(new_n14305_), .Y(new_n14306_));
  NOR3X1   g11870(.A(new_n14306_), .B(new_n14302_), .C(new_n11766_), .Y(new_n14307_));
  OAI21X1  g11871(.A0(new_n14298_), .A1(pi0789), .B0(new_n12709_), .Y(new_n14308_));
  OR2X1    g11872(.A(new_n14308_), .B(new_n14307_), .Y(new_n14309_));
  OAI22X1  g11873(.A0(new_n14230_), .A1(new_n12562_), .B0(new_n14178_), .B1(new_n13439_), .Y(new_n14310_));
  AOI21X1  g11874(.A0(new_n14310_), .A1(pi0788), .B0(new_n14125_), .Y(new_n14311_));
  AOI22X1  g11875(.A0(new_n14311_), .A1(new_n14309_), .B0(new_n14252_), .B1(pi0792), .Y(new_n14312_));
  OAI21X1  g11876(.A0(new_n14312_), .A1(new_n14121_), .B0(new_n14246_), .Y(new_n14313_));
  NOR2X1   g11877(.A(new_n14313_), .B(pi0644), .Y(new_n14314_));
  AND2X1   g11878(.A(new_n14189_), .B(pi0644), .Y(new_n14315_));
  OR2X1    g11879(.A(new_n14315_), .B(pi0715), .Y(new_n14316_));
  OAI21X1  g11880(.A0(new_n14158_), .A1(new_n12612_), .B0(pi0715), .Y(new_n14317_));
  AOI21X1  g11881(.A0(new_n14233_), .A1(new_n12612_), .B0(new_n14317_), .Y(new_n14318_));
  NOR2X1   g11882(.A(new_n14318_), .B(pi1160), .Y(new_n14319_));
  OAI21X1  g11883(.A0(new_n14316_), .A1(new_n14314_), .B0(new_n14319_), .Y(new_n14320_));
  AOI21X1  g11884(.A0(new_n14320_), .A1(new_n14236_), .B0(new_n12766_), .Y(new_n14321_));
  OR3X1    g11885(.A(new_n14235_), .B(new_n11762_), .C(new_n12612_), .Y(new_n14322_));
  AOI21X1  g11886(.A0(new_n14322_), .A1(pi0790), .B0(new_n14313_), .Y(new_n14323_));
  OAI21X1  g11887(.A0(new_n14323_), .A1(new_n14321_), .B0(new_n6489_), .Y(new_n14324_));
  AOI21X1  g11888(.A0(po1038), .A1(new_n5202_), .B0(pi0832), .Y(new_n14325_));
  INVX1    g11889(.A(new_n14239_), .Y(new_n14326_));
  INVX1    g11890(.A(new_n12580_), .Y(new_n14327_));
  AOI21X1  g11891(.A0(pi1093), .A1(pi1092), .B0(pi0145), .Y(new_n14328_));
  AOI21X1  g11892(.A0(new_n12056_), .A1(new_n14191_), .B0(new_n14328_), .Y(new_n14329_));
  AOI21X1  g11893(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n14329_), .Y(new_n14330_));
  INVX1    g11894(.A(new_n12642_), .Y(new_n14331_));
  INVX1    g11895(.A(new_n14329_), .Y(new_n14332_));
  AOI21X1  g11896(.A0(new_n14332_), .A1(new_n14331_), .B0(new_n12463_), .Y(new_n14333_));
  AOI21X1  g11897(.A0(new_n14330_), .A1(new_n12646_), .B0(pi1155), .Y(new_n14334_));
  OAI21X1  g11898(.A0(new_n14334_), .A1(new_n14333_), .B0(pi0785), .Y(new_n14335_));
  OAI21X1  g11899(.A0(new_n14330_), .A1(pi0785), .B0(new_n14335_), .Y(new_n14336_));
  INVX1    g11900(.A(new_n14336_), .Y(new_n14337_));
  AOI21X1  g11901(.A0(new_n14337_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n14338_));
  AOI21X1  g11902(.A0(new_n14337_), .A1(new_n12655_), .B0(pi1154), .Y(new_n14339_));
  NOR2X1   g11903(.A(new_n14339_), .B(new_n14338_), .Y(new_n14340_));
  MX2X1    g11904(.A(new_n14340_), .B(new_n14337_), .S0(new_n11767_), .Y(new_n14341_));
  NOR2X1   g11905(.A(new_n14341_), .B(pi0789), .Y(new_n14342_));
  INVX1    g11906(.A(new_n14341_), .Y(new_n14343_));
  AOI21X1  g11907(.A0(new_n14328_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n14344_));
  OAI21X1  g11908(.A0(new_n14343_), .A1(new_n12509_), .B0(new_n14344_), .Y(new_n14345_));
  AOI21X1  g11909(.A0(new_n14328_), .A1(pi0619), .B0(pi1159), .Y(new_n14346_));
  OAI21X1  g11910(.A0(new_n14343_), .A1(pi0619), .B0(new_n14346_), .Y(new_n14347_));
  AOI21X1  g11911(.A0(new_n14347_), .A1(new_n14345_), .B0(new_n11766_), .Y(new_n14348_));
  NOR2X1   g11912(.A(new_n14348_), .B(new_n14342_), .Y(new_n14349_));
  INVX1    g11913(.A(new_n14349_), .Y(new_n14350_));
  AOI21X1  g11914(.A0(new_n14328_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n14351_));
  OAI21X1  g11915(.A0(new_n14350_), .A1(new_n12542_), .B0(new_n14351_), .Y(new_n14352_));
  AOI21X1  g11916(.A0(new_n14328_), .A1(pi0626), .B0(pi1158), .Y(new_n14353_));
  OAI21X1  g11917(.A0(new_n14350_), .A1(pi0626), .B0(new_n14353_), .Y(new_n14354_));
  AND2X1   g11918(.A(new_n14354_), .B(new_n14352_), .Y(new_n14355_));
  MX2X1    g11919(.A(new_n14355_), .B(new_n14349_), .S0(new_n11765_), .Y(new_n14356_));
  AND3X1   g11920(.A(new_n14328_), .B(new_n12579_), .C(pi0792), .Y(new_n14357_));
  AOI21X1  g11921(.A0(new_n14356_), .A1(new_n14327_), .B0(new_n14357_), .Y(new_n14358_));
  INVX1    g11922(.A(pi0698), .Y(new_n14359_));
  AOI21X1  g11923(.A0(new_n12439_), .A1(new_n14359_), .B0(new_n14328_), .Y(new_n14360_));
  INVX1    g11924(.A(new_n14360_), .Y(new_n14361_));
  AND3X1   g11925(.A(new_n12439_), .B(new_n14359_), .C(new_n12363_), .Y(new_n14362_));
  NOR2X1   g11926(.A(new_n14362_), .B(new_n14360_), .Y(new_n14363_));
  INVX1    g11927(.A(new_n14363_), .Y(new_n14364_));
  NOR2X1   g11928(.A(new_n14328_), .B(pi1153), .Y(new_n14365_));
  INVX1    g11929(.A(new_n14365_), .Y(new_n14366_));
  NOR2X1   g11930(.A(new_n14366_), .B(new_n14362_), .Y(new_n14367_));
  AOI21X1  g11931(.A0(new_n14364_), .A1(pi1153), .B0(new_n14367_), .Y(new_n14368_));
  MX2X1    g11932(.A(new_n14368_), .B(new_n14361_), .S0(new_n11769_), .Y(new_n14369_));
  INVX1    g11933(.A(new_n14369_), .Y(new_n14370_));
  NOR3X1   g11934(.A(new_n14370_), .B(new_n12631_), .C(new_n12630_), .Y(new_n14371_));
  AND3X1   g11935(.A(new_n14371_), .B(new_n12718_), .C(new_n12634_), .Y(new_n14372_));
  AND2X1   g11936(.A(new_n14372_), .B(new_n12739_), .Y(new_n14373_));
  INVX1    g11937(.A(new_n14373_), .Y(new_n14374_));
  AOI21X1  g11938(.A0(new_n14328_), .A1(pi0647), .B0(pi1157), .Y(new_n14375_));
  OAI21X1  g11939(.A0(new_n14374_), .A1(pi0647), .B0(new_n14375_), .Y(new_n14376_));
  MX2X1    g11940(.A(new_n14373_), .B(new_n14328_), .S0(new_n12577_), .Y(new_n14377_));
  OAI22X1  g11941(.A0(new_n14377_), .A1(new_n14242_), .B0(new_n14376_), .B1(new_n12592_), .Y(new_n14378_));
  AOI21X1  g11942(.A0(new_n14358_), .A1(new_n14326_), .B0(new_n14378_), .Y(new_n14379_));
  AND3X1   g11943(.A(new_n14371_), .B(new_n12637_), .C(new_n12634_), .Y(new_n14380_));
  AND3X1   g11944(.A(new_n14354_), .B(new_n14352_), .C(new_n12639_), .Y(new_n14381_));
  OAI21X1  g11945(.A0(new_n14381_), .A1(new_n14380_), .B0(pi0788), .Y(new_n14382_));
  NOR2X1   g11946(.A(new_n14360_), .B(new_n11991_), .Y(new_n14383_));
  MX2X1    g11947(.A(new_n14332_), .B(new_n12363_), .S0(new_n14383_), .Y(new_n14384_));
  AOI21X1  g11948(.A0(new_n14364_), .A1(pi1153), .B0(pi0608), .Y(new_n14385_));
  OAI21X1  g11949(.A0(new_n14384_), .A1(new_n14366_), .B0(new_n14385_), .Y(new_n14386_));
  NOR3X1   g11950(.A(new_n14360_), .B(new_n11991_), .C(new_n12363_), .Y(new_n14387_));
  NOR3X1   g11951(.A(new_n14387_), .B(new_n14332_), .C(new_n12364_), .Y(new_n14388_));
  NOR3X1   g11952(.A(new_n14388_), .B(new_n14367_), .C(new_n12368_), .Y(new_n14389_));
  INVX1    g11953(.A(new_n14389_), .Y(new_n14390_));
  AOI21X1  g11954(.A0(new_n14390_), .A1(new_n14386_), .B0(new_n11769_), .Y(new_n14391_));
  OR2X1    g11955(.A(new_n14360_), .B(new_n11991_), .Y(new_n14392_));
  AOI21X1  g11956(.A0(new_n14392_), .A1(new_n14329_), .B0(pi0778), .Y(new_n14393_));
  NOR2X1   g11957(.A(new_n14393_), .B(new_n14391_), .Y(new_n14394_));
  OAI21X1  g11958(.A0(new_n14393_), .A1(new_n14391_), .B0(new_n12462_), .Y(new_n14395_));
  AOI21X1  g11959(.A0(new_n14369_), .A1(pi0609), .B0(pi1155), .Y(new_n14396_));
  OR2X1    g11960(.A(new_n14333_), .B(pi0660), .Y(new_n14397_));
  AOI21X1  g11961(.A0(new_n14396_), .A1(new_n14395_), .B0(new_n14397_), .Y(new_n14398_));
  OAI21X1  g11962(.A0(new_n14393_), .A1(new_n14391_), .B0(pi0609), .Y(new_n14399_));
  AOI21X1  g11963(.A0(new_n14369_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n14400_));
  OR2X1    g11964(.A(new_n14334_), .B(new_n12468_), .Y(new_n14401_));
  AOI21X1  g11965(.A0(new_n14400_), .A1(new_n14399_), .B0(new_n14401_), .Y(new_n14402_));
  NOR2X1   g11966(.A(new_n14402_), .B(new_n14398_), .Y(new_n14403_));
  MX2X1    g11967(.A(new_n14403_), .B(new_n14394_), .S0(new_n11768_), .Y(new_n14404_));
  OR3X1    g11968(.A(new_n14370_), .B(new_n12630_), .C(new_n12486_), .Y(new_n14405_));
  AND2X1   g11969(.A(new_n14405_), .B(new_n12487_), .Y(new_n14406_));
  OAI21X1  g11970(.A0(new_n14404_), .A1(pi0618), .B0(new_n14406_), .Y(new_n14407_));
  NOR2X1   g11971(.A(new_n14338_), .B(pi0627), .Y(new_n14408_));
  NOR3X1   g11972(.A(new_n14370_), .B(new_n12630_), .C(pi0618), .Y(new_n14409_));
  NOR2X1   g11973(.A(new_n14409_), .B(new_n12487_), .Y(new_n14410_));
  OAI21X1  g11974(.A0(new_n14404_), .A1(new_n12486_), .B0(new_n14410_), .Y(new_n14411_));
  NOR2X1   g11975(.A(new_n14339_), .B(new_n12494_), .Y(new_n14412_));
  AOI22X1  g11976(.A0(new_n14412_), .A1(new_n14411_), .B0(new_n14408_), .B1(new_n14407_), .Y(new_n14413_));
  MX2X1    g11977(.A(new_n14413_), .B(new_n14404_), .S0(new_n11767_), .Y(new_n14414_));
  AOI21X1  g11978(.A0(new_n14371_), .A1(pi0619), .B0(pi1159), .Y(new_n14415_));
  OAI21X1  g11979(.A0(new_n14414_), .A1(pi0619), .B0(new_n14415_), .Y(new_n14416_));
  AND3X1   g11980(.A(new_n14416_), .B(new_n14345_), .C(new_n12517_), .Y(new_n14417_));
  AOI21X1  g11981(.A0(new_n14371_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n14418_));
  OAI21X1  g11982(.A0(new_n14414_), .A1(new_n12509_), .B0(new_n14418_), .Y(new_n14419_));
  AND2X1   g11983(.A(new_n14347_), .B(pi0648), .Y(new_n14420_));
  AOI21X1  g11984(.A0(new_n14420_), .A1(new_n14419_), .B0(new_n11766_), .Y(new_n14421_));
  INVX1    g11985(.A(new_n14421_), .Y(new_n14422_));
  AOI21X1  g11986(.A0(new_n14414_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n14423_));
  OAI21X1  g11987(.A0(new_n14422_), .A1(new_n14417_), .B0(new_n14423_), .Y(new_n14424_));
  AOI21X1  g11988(.A0(new_n14424_), .A1(new_n14382_), .B0(new_n14125_), .Y(new_n14425_));
  AOI21X1  g11989(.A0(new_n2720_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n14426_));
  AOI22X1  g11990(.A0(new_n14426_), .A1(new_n14372_), .B0(new_n14356_), .B1(new_n12735_), .Y(new_n14427_));
  AOI21X1  g11991(.A0(new_n2720_), .A1(pi0628), .B0(pi1156), .Y(new_n14428_));
  AOI22X1  g11992(.A0(new_n14428_), .A1(new_n14372_), .B0(new_n14356_), .B1(new_n12733_), .Y(new_n14429_));
  MX2X1    g11993(.A(new_n14429_), .B(new_n14427_), .S0(new_n12561_), .Y(new_n14430_));
  OAI21X1  g11994(.A0(new_n14430_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n14431_));
  OAI22X1  g11995(.A0(new_n14431_), .A1(new_n14425_), .B0(new_n14379_), .B1(new_n11763_), .Y(new_n14432_));
  INVX1    g11996(.A(new_n14432_), .Y(new_n14433_));
  OAI21X1  g11997(.A0(new_n14377_), .A1(new_n12578_), .B0(new_n14376_), .Y(new_n14434_));
  MX2X1    g11998(.A(new_n14434_), .B(new_n14374_), .S0(new_n11763_), .Y(new_n14435_));
  OAI21X1  g11999(.A0(new_n14435_), .A1(pi0644), .B0(pi0715), .Y(new_n14436_));
  AOI21X1  g12000(.A0(new_n14433_), .A1(pi0644), .B0(new_n14436_), .Y(new_n14437_));
  INVX1    g12001(.A(new_n14328_), .Y(new_n14438_));
  OR3X1    g12002(.A(new_n14438_), .B(new_n12603_), .C(new_n11763_), .Y(new_n14439_));
  OAI21X1  g12003(.A0(new_n14358_), .A1(new_n12604_), .B0(new_n14439_), .Y(new_n14440_));
  OAI21X1  g12004(.A0(new_n14438_), .A1(pi0644), .B0(new_n12608_), .Y(new_n14441_));
  AOI21X1  g12005(.A0(new_n14440_), .A1(pi0644), .B0(new_n14441_), .Y(new_n14442_));
  OR2X1    g12006(.A(new_n14442_), .B(new_n11762_), .Y(new_n14443_));
  OAI21X1  g12007(.A0(new_n14435_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n14444_));
  AOI21X1  g12008(.A0(new_n14433_), .A1(new_n12612_), .B0(new_n14444_), .Y(new_n14445_));
  OAI21X1  g12009(.A0(new_n14438_), .A1(new_n12612_), .B0(pi0715), .Y(new_n14446_));
  AOI21X1  g12010(.A0(new_n14440_), .A1(new_n12612_), .B0(new_n14446_), .Y(new_n14447_));
  OR2X1    g12011(.A(new_n14447_), .B(pi1160), .Y(new_n14448_));
  OAI22X1  g12012(.A0(new_n14448_), .A1(new_n14445_), .B0(new_n14443_), .B1(new_n14437_), .Y(new_n14449_));
  OAI21X1  g12013(.A0(new_n14432_), .A1(pi0790), .B0(pi0832), .Y(new_n14450_));
  AOI21X1  g12014(.A0(new_n14449_), .A1(pi0790), .B0(new_n14450_), .Y(new_n14451_));
  AOI21X1  g12015(.A0(new_n14325_), .A1(new_n14324_), .B0(new_n14451_), .Y(po0302));
  AND2X1   g12016(.A(new_n5362_), .B(pi0907), .Y(new_n14453_));
  AOI22X1  g12017(.A0(new_n14453_), .A1(pi0735), .B0(pi0947), .B1(pi0743), .Y(new_n14454_));
  AND2X1   g12018(.A(new_n14454_), .B(new_n2720_), .Y(new_n14455_));
  NOR4X1   g12019(.A(new_n5056_), .B(pi0963), .C(pi0960), .D(pi0907), .Y(new_n14456_));
  NOR3X1   g12020(.A(new_n14456_), .B(new_n11932_), .C(new_n2776_), .Y(new_n14457_));
  INVX1    g12021(.A(new_n14456_), .Y(new_n14458_));
  OR3X1    g12022(.A(new_n14458_), .B(new_n11924_), .C(new_n2776_), .Y(new_n14459_));
  OR4X1    g12023(.A(new_n11931_), .B(new_n11927_), .C(new_n5277_), .D(new_n13171_), .Y(new_n14460_));
  AND2X1   g12024(.A(new_n14460_), .B(new_n5362_), .Y(new_n14461_));
  OAI21X1  g12025(.A0(new_n11931_), .A1(new_n11927_), .B0(pi0146), .Y(new_n14462_));
  OR3X1    g12026(.A(new_n11931_), .B(new_n11927_), .C(new_n13086_), .Y(new_n14463_));
  AND3X1   g12027(.A(new_n14463_), .B(new_n14462_), .C(pi0947), .Y(new_n14464_));
  AOI21X1  g12028(.A0(new_n14461_), .A1(new_n14459_), .B0(new_n14464_), .Y(new_n14465_));
  OAI21X1  g12029(.A0(new_n14465_), .A1(new_n14457_), .B0(new_n10045_), .Y(new_n14466_));
  INVX1    g12030(.A(new_n14454_), .Y(new_n14467_));
  MX2X1    g12031(.A(new_n14467_), .B(pi0146), .S0(new_n11825_), .Y(new_n14468_));
  AOI21X1  g12032(.A0(new_n14468_), .A1(new_n10044_), .B0(pi0215), .Y(new_n14469_));
  OR3X1    g12033(.A(new_n11955_), .B(new_n11951_), .C(new_n2776_), .Y(new_n14470_));
  AOI21X1  g12034(.A0(new_n14467_), .A1(new_n11862_), .B0(new_n2934_), .Y(new_n14471_));
  AOI22X1  g12035(.A0(new_n14471_), .A1(new_n14470_), .B0(new_n14469_), .B1(new_n14466_), .Y(new_n14472_));
  NOR3X1   g12036(.A(new_n14454_), .B(new_n11931_), .C(new_n11927_), .Y(new_n14473_));
  NAND2X1  g12037(.A(new_n14462_), .B(new_n5042_), .Y(new_n14474_));
  AND2X1   g12038(.A(new_n14467_), .B(new_n11924_), .Y(new_n14475_));
  OAI21X1  g12039(.A0(new_n11924_), .A1(new_n2776_), .B0(new_n5041_), .Y(new_n14476_));
  OAI22X1  g12040(.A0(new_n14476_), .A1(new_n14475_), .B0(new_n14474_), .B1(new_n14473_), .Y(new_n14477_));
  OAI21X1  g12041(.A0(new_n14468_), .A1(new_n2952_), .B0(new_n2940_), .Y(new_n14478_));
  AOI21X1  g12042(.A0(new_n14477_), .A1(new_n2952_), .B0(new_n14478_), .Y(new_n14479_));
  MX2X1    g12043(.A(pi0146), .B(new_n14467_), .S0(new_n11862_), .Y(new_n14480_));
  OR2X1    g12044(.A(new_n11877_), .B(pi0146), .Y(new_n14481_));
  AOI21X1  g12045(.A0(new_n14454_), .A1(new_n11877_), .B0(new_n5042_), .Y(new_n14482_));
  AOI22X1  g12046(.A0(new_n14482_), .A1(new_n14481_), .B0(new_n14480_), .B1(new_n5042_), .Y(new_n14483_));
  OAI21X1  g12047(.A0(new_n14483_), .A1(new_n2940_), .B0(new_n2933_), .Y(new_n14484_));
  OAI22X1  g12048(.A0(new_n14484_), .A1(new_n14479_), .B0(new_n14472_), .B1(new_n2933_), .Y(new_n14485_));
  OAI21X1  g12049(.A0(new_n14467_), .A1(new_n11961_), .B0(pi0299), .Y(new_n14486_));
  AOI21X1  g12050(.A0(new_n11961_), .A1(new_n2776_), .B0(new_n14486_), .Y(new_n14487_));
  AND2X1   g12051(.A(new_n12306_), .B(new_n2776_), .Y(new_n14488_));
  OAI21X1  g12052(.A0(new_n14467_), .A1(new_n12306_), .B0(new_n2933_), .Y(new_n14489_));
  OAI21X1  g12053(.A0(new_n14489_), .A1(new_n14488_), .B0(new_n2939_), .Y(new_n14490_));
  OAI21X1  g12054(.A0(new_n14490_), .A1(new_n14487_), .B0(new_n2979_), .Y(new_n14491_));
  AOI21X1  g12055(.A0(new_n14485_), .A1(pi0039), .B0(new_n14491_), .Y(new_n14492_));
  OR2X1    g12056(.A(new_n12077_), .B(pi0146), .Y(new_n14493_));
  AOI21X1  g12057(.A0(new_n14455_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n14494_));
  AND2X1   g12058(.A(new_n14494_), .B(new_n14493_), .Y(new_n14495_));
  NOR3X1   g12059(.A(new_n14495_), .B(new_n14492_), .C(new_n9483_), .Y(new_n14496_));
  OAI21X1  g12060(.A0(new_n7625_), .A1(pi0146), .B0(new_n12767_), .Y(new_n14497_));
  OAI21X1  g12061(.A0(new_n2720_), .A1(pi0146), .B0(pi0832), .Y(new_n14498_));
  OAI22X1  g12062(.A0(new_n14498_), .A1(new_n14455_), .B0(new_n14497_), .B1(new_n14496_), .Y(po0303));
  INVX1    g12063(.A(pi0726), .Y(new_n14500_));
  INVX1    g12064(.A(new_n14453_), .Y(new_n14501_));
  OAI22X1  g12065(.A0(new_n14501_), .A1(new_n14500_), .B0(new_n5362_), .B1(pi0770), .Y(new_n14502_));
  OAI21X1  g12066(.A0(new_n2720_), .A1(pi0147), .B0(pi0832), .Y(new_n14503_));
  AOI21X1  g12067(.A0(new_n14502_), .A1(new_n2720_), .B0(new_n14503_), .Y(new_n14504_));
  AOI21X1  g12068(.A0(new_n11821_), .A1(new_n5362_), .B0(pi0039), .Y(new_n14505_));
  NOR4X1   g12069(.A(new_n11936_), .B(new_n11879_), .C(new_n5362_), .D(pi0299), .Y(new_n14506_));
  INVX1    g12070(.A(new_n14506_), .Y(new_n14507_));
  NOR2X1   g12071(.A(new_n11936_), .B(new_n11879_), .Y(new_n14508_));
  OR4X1    g12072(.A(new_n11824_), .B(new_n10045_), .C(new_n2725_), .D(pi0947), .Y(new_n14509_));
  AOI21X1  g12073(.A0(new_n14453_), .A1(new_n11932_), .B0(new_n11945_), .Y(new_n14510_));
  NOR2X1   g12074(.A(new_n14510_), .B(new_n10044_), .Y(new_n14511_));
  NOR2X1   g12075(.A(new_n14511_), .B(pi0215), .Y(new_n14512_));
  NOR3X1   g12076(.A(new_n14501_), .B(new_n11861_), .C(new_n11847_), .Y(new_n14513_));
  NOR3X1   g12077(.A(new_n14513_), .B(new_n11955_), .C(new_n2934_), .Y(new_n14514_));
  AOI21X1  g12078(.A0(new_n14512_), .A1(new_n14509_), .B0(new_n14514_), .Y(new_n14515_));
  MX2X1    g12079(.A(new_n14515_), .B(new_n14508_), .S0(new_n2933_), .Y(new_n14516_));
  AOI21X1  g12080(.A0(new_n14516_), .A1(new_n14507_), .B0(new_n2939_), .Y(new_n14517_));
  NOR3X1   g12081(.A(new_n14517_), .B(new_n14505_), .C(pi0038), .Y(new_n14518_));
  AND3X1   g12082(.A(new_n12446_), .B(new_n5362_), .C(pi0038), .Y(new_n14519_));
  NOR2X1   g12083(.A(new_n14519_), .B(new_n14518_), .Y(new_n14520_));
  MX2X1    g12084(.A(new_n14520_), .B(new_n12832_), .S0(pi0770), .Y(new_n14521_));
  INVX1    g12085(.A(pi0770), .Y(new_n14522_));
  NOR2X1   g12086(.A(new_n14519_), .B(new_n13265_), .Y(new_n14523_));
  AOI21X1  g12087(.A0(new_n11821_), .A1(pi0947), .B0(pi0039), .Y(new_n14524_));
  NOR3X1   g12088(.A(new_n11936_), .B(new_n11879_), .C(new_n5362_), .Y(new_n14525_));
  NOR2X1   g12089(.A(new_n14525_), .B(pi0299), .Y(new_n14526_));
  NOR4X1   g12090(.A(new_n11861_), .B(new_n11847_), .C(new_n5362_), .D(new_n2934_), .Y(new_n14527_));
  OR3X1    g12091(.A(new_n11931_), .B(new_n11927_), .C(new_n5362_), .Y(new_n14528_));
  NOR3X1   g12092(.A(new_n11824_), .B(new_n2725_), .C(new_n5362_), .Y(new_n14529_));
  OAI21X1  g12093(.A0(new_n14529_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n14530_));
  AOI21X1  g12094(.A0(new_n14528_), .A1(new_n10045_), .B0(new_n14530_), .Y(new_n14531_));
  NOR3X1   g12095(.A(new_n14531_), .B(new_n14527_), .C(new_n2933_), .Y(new_n14532_));
  NOR2X1   g12096(.A(new_n14532_), .B(new_n14526_), .Y(new_n14533_));
  INVX1    g12097(.A(new_n14533_), .Y(new_n14534_));
  AOI21X1  g12098(.A0(new_n14534_), .A1(pi0039), .B0(new_n14524_), .Y(new_n14535_));
  OR2X1    g12099(.A(new_n14535_), .B(pi0038), .Y(new_n14536_));
  NAND4X1  g12100(.A(new_n14536_), .B(new_n14523_), .C(new_n14522_), .D(pi0147), .Y(new_n14537_));
  NAND2X1  g12101(.A(new_n14537_), .B(new_n14500_), .Y(new_n14538_));
  AOI21X1  g12102(.A0(new_n14521_), .A1(new_n8649_), .B0(new_n14538_), .Y(new_n14539_));
  NOR2X1   g12103(.A(new_n11955_), .B(new_n2934_), .Y(new_n14540_));
  INVX1    g12104(.A(new_n14540_), .Y(new_n14541_));
  AOI21X1  g12105(.A0(new_n11932_), .A1(pi0947), .B0(new_n11945_), .Y(new_n14542_));
  OAI21X1  g12106(.A0(new_n14542_), .A1(new_n10044_), .B0(new_n2934_), .Y(new_n14543_));
  AOI21X1  g12107(.A0(new_n14501_), .A1(new_n11947_), .B0(new_n14543_), .Y(new_n14544_));
  INVX1    g12108(.A(new_n14544_), .Y(new_n14545_));
  AOI21X1  g12109(.A0(new_n14545_), .A1(new_n14541_), .B0(new_n2933_), .Y(new_n14546_));
  INVX1    g12110(.A(new_n5055_), .Y(new_n14547_));
  AOI22X1  g12111(.A0(new_n11934_), .A1(new_n2987_), .B0(new_n11933_), .B1(new_n2952_), .Y(new_n14548_));
  OAI21X1  g12112(.A0(new_n14548_), .A1(new_n14547_), .B0(new_n2940_), .Y(new_n14549_));
  AOI21X1  g12113(.A0(new_n11878_), .A1(new_n5362_), .B0(new_n2940_), .Y(new_n14550_));
  AOI21X1  g12114(.A0(new_n14501_), .A1(new_n11878_), .B0(new_n2940_), .Y(new_n14551_));
  NOR2X1   g12115(.A(new_n14551_), .B(new_n14550_), .Y(new_n14552_));
  AOI21X1  g12116(.A0(new_n14552_), .A1(new_n14549_), .B0(pi0299), .Y(new_n14553_));
  AND2X1   g12117(.A(pi0947), .B(pi0299), .Y(new_n14554_));
  NOR3X1   g12118(.A(new_n14554_), .B(new_n14553_), .C(new_n14546_), .Y(new_n14555_));
  AOI21X1  g12119(.A0(new_n11821_), .A1(new_n14547_), .B0(pi0039), .Y(new_n14556_));
  AOI22X1  g12120(.A0(new_n14556_), .A1(new_n11821_), .B0(new_n14555_), .B1(pi0039), .Y(new_n14557_));
  INVX1    g12121(.A(new_n14557_), .Y(new_n14558_));
  OR4X1    g12122(.A(new_n11936_), .B(new_n11879_), .C(new_n5055_), .D(pi0299), .Y(new_n14559_));
  NOR3X1   g12123(.A(new_n11824_), .B(new_n5055_), .C(new_n2725_), .Y(new_n14560_));
  AOI21X1  g12124(.A0(new_n14560_), .A1(new_n10044_), .B0(pi0215), .Y(new_n14561_));
  AOI21X1  g12125(.A0(new_n14561_), .A1(new_n11946_), .B0(new_n2933_), .Y(new_n14562_));
  OAI21X1  g12126(.A0(new_n11951_), .A1(new_n2934_), .B0(new_n14562_), .Y(new_n14563_));
  AND2X1   g12127(.A(new_n14563_), .B(new_n14559_), .Y(new_n14564_));
  AOI21X1  g12128(.A0(new_n14564_), .A1(pi0039), .B0(new_n14556_), .Y(new_n14565_));
  AOI21X1  g12129(.A0(new_n14565_), .A1(pi0147), .B0(pi0038), .Y(new_n14566_));
  OAI21X1  g12130(.A0(new_n14558_), .A1(pi0147), .B0(new_n14566_), .Y(new_n14567_));
  AND2X1   g12131(.A(new_n12446_), .B(new_n5055_), .Y(new_n14568_));
  AOI21X1  g12132(.A0(new_n12077_), .A1(new_n14547_), .B0(new_n2979_), .Y(new_n14569_));
  OAI21X1  g12133(.A0(new_n14568_), .A1(pi0147), .B0(new_n14569_), .Y(new_n14570_));
  AND2X1   g12134(.A(new_n14570_), .B(new_n14522_), .Y(new_n14571_));
  AOI21X1  g12135(.A0(new_n14545_), .A1(new_n14541_), .B0(new_n14527_), .Y(new_n14572_));
  OR4X1    g12136(.A(new_n14453_), .B(new_n11936_), .C(new_n11879_), .D(pi0299), .Y(new_n14573_));
  OAI21X1  g12137(.A0(new_n14572_), .A1(new_n2933_), .B0(new_n14573_), .Y(new_n14574_));
  AND2X1   g12138(.A(new_n14501_), .B(new_n11821_), .Y(new_n14575_));
  MX2X1    g12139(.A(new_n14575_), .B(new_n14574_), .S0(pi0039), .Y(new_n14576_));
  INVX1    g12140(.A(new_n14576_), .Y(new_n14577_));
  AOI21X1  g12141(.A0(new_n14453_), .A1(new_n11932_), .B0(new_n10044_), .Y(new_n14578_));
  NOR3X1   g12142(.A(new_n11824_), .B(new_n2725_), .C(new_n5277_), .Y(new_n14579_));
  AOI21X1  g12143(.A0(new_n14579_), .A1(new_n5362_), .B0(new_n10045_), .Y(new_n14580_));
  OAI21X1  g12144(.A0(new_n14580_), .A1(new_n14578_), .B0(new_n2934_), .Y(new_n14581_));
  OAI21X1  g12145(.A0(new_n14513_), .A1(new_n2934_), .B0(new_n14581_), .Y(new_n14582_));
  AND2X1   g12146(.A(new_n14582_), .B(pi0299), .Y(new_n14583_));
  OR3X1    g12147(.A(new_n14501_), .B(new_n11936_), .C(new_n11879_), .Y(new_n14584_));
  AOI21X1  g12148(.A0(new_n14584_), .A1(new_n2933_), .B0(new_n14583_), .Y(new_n14585_));
  AND2X1   g12149(.A(new_n14453_), .B(new_n11821_), .Y(new_n14586_));
  MX2X1    g12150(.A(new_n14586_), .B(new_n14585_), .S0(pi0039), .Y(new_n14587_));
  INVX1    g12151(.A(new_n14587_), .Y(new_n14588_));
  OAI21X1  g12152(.A0(new_n14588_), .A1(new_n8649_), .B0(new_n2979_), .Y(new_n14589_));
  AOI21X1  g12153(.A0(new_n14577_), .A1(new_n8649_), .B0(new_n14589_), .Y(new_n14590_));
  AOI21X1  g12154(.A0(new_n14453_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n14591_));
  OAI21X1  g12155(.A0(new_n12077_), .A1(pi0147), .B0(new_n14591_), .Y(new_n14592_));
  NAND2X1  g12156(.A(new_n14592_), .B(pi0770), .Y(new_n14593_));
  OAI21X1  g12157(.A0(new_n14593_), .A1(new_n14590_), .B0(pi0726), .Y(new_n14594_));
  AOI21X1  g12158(.A0(new_n14571_), .A1(new_n14567_), .B0(new_n14594_), .Y(new_n14595_));
  OR3X1    g12159(.A(new_n14595_), .B(new_n14539_), .C(new_n9483_), .Y(new_n14596_));
  AOI21X1  g12160(.A0(new_n9483_), .A1(new_n8649_), .B0(pi0832), .Y(new_n14597_));
  AOI21X1  g12161(.A0(new_n14597_), .A1(new_n14596_), .B0(new_n14504_), .Y(po0304));
  INVX1    g12162(.A(new_n14508_), .Y(new_n14599_));
  AOI21X1  g12163(.A0(new_n14599_), .A1(new_n2933_), .B0(new_n14583_), .Y(new_n14600_));
  OAI21X1  g12164(.A0(new_n14600_), .A1(new_n4046_), .B0(new_n12774_), .Y(new_n14601_));
  AOI21X1  g12165(.A0(new_n14574_), .A1(new_n11611_), .B0(new_n14601_), .Y(new_n14602_));
  INVX1    g12166(.A(new_n14564_), .Y(new_n14603_));
  OAI21X1  g12167(.A0(new_n14603_), .A1(new_n4046_), .B0(pi0749), .Y(new_n14604_));
  AOI21X1  g12168(.A0(new_n14555_), .A1(new_n4046_), .B0(new_n14604_), .Y(new_n14605_));
  NOR3X1   g12169(.A(new_n14605_), .B(new_n14602_), .C(new_n2939_), .Y(new_n14606_));
  OAI21X1  g12170(.A0(new_n11821_), .A1(pi0148), .B0(new_n2939_), .Y(new_n14607_));
  AND2X1   g12171(.A(pi0947), .B(new_n12774_), .Y(new_n14608_));
  NOR3X1   g12172(.A(new_n14608_), .B(new_n11822_), .C(new_n5055_), .Y(new_n14609_));
  OAI21X1  g12173(.A0(new_n14609_), .A1(new_n14607_), .B0(new_n2979_), .Y(new_n14610_));
  NAND2X1  g12174(.A(new_n12077_), .B(new_n14547_), .Y(new_n14611_));
  OAI22X1  g12175(.A0(new_n14608_), .A1(new_n14611_), .B0(new_n12077_), .B1(pi0148), .Y(new_n14612_));
  AOI21X1  g12176(.A0(new_n14612_), .A1(pi0038), .B0(new_n12805_), .Y(new_n14613_));
  OAI21X1  g12177(.A0(new_n14610_), .A1(new_n14606_), .B0(new_n14613_), .Y(new_n14614_));
  AND2X1   g12178(.A(new_n5102_), .B(new_n3103_), .Y(new_n14615_));
  INVX1    g12179(.A(new_n14615_), .Y(new_n14616_));
  OR2X1    g12180(.A(new_n14531_), .B(new_n14527_), .Y(new_n14617_));
  AOI21X1  g12181(.A0(new_n14617_), .A1(pi0148), .B0(new_n2933_), .Y(new_n14618_));
  OAI21X1  g12182(.A0(new_n14515_), .A1(pi0148), .B0(new_n14618_), .Y(new_n14619_));
  OAI21X1  g12183(.A0(new_n11936_), .A1(new_n11879_), .B0(new_n4046_), .Y(new_n14620_));
  AOI21X1  g12184(.A0(new_n14620_), .A1(new_n14526_), .B0(new_n12774_), .Y(new_n14621_));
  OR2X1    g12185(.A(pi0749), .B(pi0148), .Y(new_n14622_));
  OAI21X1  g12186(.A0(new_n14622_), .A1(new_n12444_), .B0(pi0039), .Y(new_n14623_));
  AOI21X1  g12187(.A0(new_n14621_), .A1(new_n14619_), .B0(new_n14623_), .Y(new_n14624_));
  AND2X1   g12188(.A(pi0947), .B(pi0749), .Y(new_n14625_));
  AOI21X1  g12189(.A0(new_n14625_), .A1(new_n11821_), .B0(new_n14607_), .Y(new_n14626_));
  OR3X1    g12190(.A(new_n14626_), .B(new_n14624_), .C(pi0038), .Y(new_n14627_));
  INVX1    g12191(.A(new_n14625_), .Y(new_n14628_));
  AOI21X1  g12192(.A0(new_n14628_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n14629_));
  OAI21X1  g12193(.A0(new_n12446_), .A1(new_n4046_), .B0(new_n14629_), .Y(new_n14630_));
  AND2X1   g12194(.A(new_n14630_), .B(new_n12805_), .Y(new_n14631_));
  AOI21X1  g12195(.A0(new_n14631_), .A1(new_n14627_), .B0(new_n14616_), .Y(new_n14632_));
  OAI21X1  g12196(.A0(new_n14615_), .A1(pi0148), .B0(new_n2436_), .Y(new_n14633_));
  AOI21X1  g12197(.A0(new_n14632_), .A1(new_n14614_), .B0(new_n14633_), .Y(new_n14634_));
  OAI21X1  g12198(.A0(new_n4046_), .A1(new_n2436_), .B0(new_n12767_), .Y(new_n14635_));
  OAI21X1  g12199(.A0(new_n5362_), .A1(new_n12774_), .B0(new_n2720_), .Y(new_n14636_));
  AOI21X1  g12200(.A0(new_n14453_), .A1(pi0706), .B0(new_n14636_), .Y(new_n14637_));
  OAI21X1  g12201(.A0(new_n2720_), .A1(new_n4046_), .B0(pi0832), .Y(new_n14638_));
  OAI22X1  g12202(.A0(new_n14638_), .A1(new_n14637_), .B0(new_n14635_), .B1(new_n14634_), .Y(po0305));
  INVX1    g12203(.A(pi0755), .Y(new_n14640_));
  AND2X1   g12204(.A(pi0947), .B(new_n14640_), .Y(new_n14641_));
  INVX1    g12205(.A(new_n14641_), .Y(new_n14642_));
  OAI21X1  g12206(.A0(new_n14501_), .A1(pi0725), .B0(new_n14642_), .Y(new_n14643_));
  OAI21X1  g12207(.A0(new_n2720_), .A1(pi0149), .B0(pi0832), .Y(new_n14644_));
  AOI21X1  g12208(.A0(new_n14643_), .A1(new_n2720_), .B0(new_n14644_), .Y(new_n14645_));
  AOI21X1  g12209(.A0(new_n14642_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n14646_));
  OAI21X1  g12210(.A0(new_n12446_), .A1(new_n7101_), .B0(new_n14646_), .Y(new_n14647_));
  AND2X1   g12211(.A(pi0299), .B(new_n7101_), .Y(new_n14648_));
  OAI22X1  g12212(.A0(new_n14532_), .A1(new_n14648_), .B0(new_n14515_), .B1(pi0149), .Y(new_n14649_));
  OAI21X1  g12213(.A0(new_n11936_), .A1(new_n11879_), .B0(new_n7101_), .Y(new_n14650_));
  AOI21X1  g12214(.A0(new_n14650_), .A1(new_n14526_), .B0(pi0755), .Y(new_n14651_));
  OR2X1    g12215(.A(new_n14640_), .B(pi0149), .Y(new_n14652_));
  OAI21X1  g12216(.A0(new_n14652_), .A1(new_n12444_), .B0(pi0039), .Y(new_n14653_));
  AOI21X1  g12217(.A0(new_n14651_), .A1(new_n14649_), .B0(new_n14653_), .Y(new_n14654_));
  AOI21X1  g12218(.A0(new_n14641_), .A1(new_n11821_), .B0(pi0039), .Y(new_n14655_));
  OAI21X1  g12219(.A0(new_n11821_), .A1(pi0149), .B0(new_n14655_), .Y(new_n14656_));
  NAND2X1  g12220(.A(new_n14656_), .B(new_n2979_), .Y(new_n14657_));
  OAI21X1  g12221(.A0(new_n14657_), .A1(new_n14654_), .B0(new_n14647_), .Y(new_n14658_));
  AND2X1   g12222(.A(new_n14658_), .B(pi0725), .Y(new_n14659_));
  OAI21X1  g12223(.A0(new_n14603_), .A1(new_n7101_), .B0(new_n14640_), .Y(new_n14660_));
  AOI21X1  g12224(.A0(new_n14555_), .A1(new_n7101_), .B0(new_n14660_), .Y(new_n14661_));
  NOR3X1   g12225(.A(new_n14572_), .B(new_n2933_), .C(pi0149), .Y(new_n14662_));
  AND2X1   g12226(.A(new_n14573_), .B(pi0755), .Y(new_n14663_));
  OAI21X1  g12227(.A0(new_n14600_), .A1(new_n7101_), .B0(new_n14663_), .Y(new_n14664_));
  OAI21X1  g12228(.A0(new_n14664_), .A1(new_n14662_), .B0(pi0039), .Y(new_n14665_));
  OAI22X1  g12229(.A0(new_n14665_), .A1(new_n14661_), .B0(new_n14656_), .B1(new_n14586_), .Y(new_n14666_));
  INVX1    g12230(.A(pi0725), .Y(new_n14667_));
  NOR2X1   g12231(.A(new_n12077_), .B(pi0149), .Y(new_n14668_));
  OR4X1    g12232(.A(new_n5055_), .B(new_n2985_), .C(new_n2725_), .D(new_n2536_), .Y(new_n14669_));
  OAI21X1  g12233(.A0(new_n5362_), .A1(new_n14640_), .B0(new_n2939_), .Y(new_n14670_));
  OAI21X1  g12234(.A0(new_n14670_), .A1(new_n14669_), .B0(pi0038), .Y(new_n14671_));
  OAI21X1  g12235(.A0(new_n14671_), .A1(new_n14668_), .B0(new_n14667_), .Y(new_n14672_));
  AOI21X1  g12236(.A0(new_n14666_), .A1(new_n2979_), .B0(new_n14672_), .Y(new_n14673_));
  OAI21X1  g12237(.A0(new_n14673_), .A1(new_n14659_), .B0(new_n7625_), .Y(new_n14674_));
  AOI21X1  g12238(.A0(new_n9483_), .A1(new_n7101_), .B0(pi0832), .Y(new_n14675_));
  AOI21X1  g12239(.A0(new_n14675_), .A1(new_n14674_), .B0(new_n14645_), .Y(po0306));
  AND2X1   g12240(.A(new_n14516_), .B(new_n14507_), .Y(new_n14677_));
  INVX1    g12241(.A(pi0751), .Y(new_n14678_));
  OAI21X1  g12242(.A0(new_n14533_), .A1(new_n9837_), .B0(new_n14678_), .Y(new_n14679_));
  AOI21X1  g12243(.A0(new_n14677_), .A1(new_n9837_), .B0(new_n14679_), .Y(new_n14680_));
  NOR3X1   g12244(.A(new_n12444_), .B(new_n14678_), .C(pi0150), .Y(new_n14681_));
  OAI21X1  g12245(.A0(new_n14681_), .A1(new_n14680_), .B0(pi0039), .Y(new_n14682_));
  MX2X1    g12246(.A(new_n9837_), .B(new_n14678_), .S0(new_n11821_), .Y(new_n14683_));
  AOI21X1  g12247(.A0(new_n14683_), .A1(new_n14505_), .B0(pi0038), .Y(new_n14684_));
  OR2X1    g12248(.A(new_n5362_), .B(pi0751), .Y(new_n14685_));
  AOI22X1  g12249(.A0(new_n14685_), .A1(new_n12077_), .B0(new_n12831_), .B1(pi0150), .Y(new_n14686_));
  OAI21X1  g12250(.A0(new_n14686_), .A1(new_n2979_), .B0(pi0701), .Y(new_n14687_));
  AOI21X1  g12251(.A0(new_n14684_), .A1(new_n14682_), .B0(new_n14687_), .Y(new_n14688_));
  OAI21X1  g12252(.A0(new_n14585_), .A1(new_n9837_), .B0(pi0751), .Y(new_n14689_));
  AOI21X1  g12253(.A0(new_n14574_), .A1(new_n9837_), .B0(new_n14689_), .Y(new_n14690_));
  OAI21X1  g12254(.A0(new_n14603_), .A1(new_n9837_), .B0(new_n14678_), .Y(new_n14691_));
  AOI21X1  g12255(.A0(new_n14555_), .A1(new_n9837_), .B0(new_n14691_), .Y(new_n14692_));
  OAI21X1  g12256(.A0(new_n14692_), .A1(new_n14690_), .B0(pi0039), .Y(new_n14693_));
  NAND3X1  g12257(.A(new_n14685_), .B(new_n14501_), .C(new_n11821_), .Y(new_n14694_));
  AOI21X1  g12258(.A0(new_n11822_), .A1(pi0150), .B0(pi0039), .Y(new_n14695_));
  AOI21X1  g12259(.A0(new_n14695_), .A1(new_n14694_), .B0(pi0038), .Y(new_n14696_));
  INVX1    g12260(.A(pi0701), .Y(new_n14697_));
  NOR2X1   g12261(.A(new_n12077_), .B(pi0150), .Y(new_n14698_));
  OAI21X1  g12262(.A0(new_n5362_), .A1(new_n14678_), .B0(new_n2939_), .Y(new_n14699_));
  OAI21X1  g12263(.A0(new_n14699_), .A1(new_n14669_), .B0(pi0038), .Y(new_n14700_));
  OAI21X1  g12264(.A0(new_n14700_), .A1(new_n14698_), .B0(new_n14697_), .Y(new_n14701_));
  AOI21X1  g12265(.A0(new_n14696_), .A1(new_n14693_), .B0(new_n14701_), .Y(new_n14702_));
  OAI21X1  g12266(.A0(new_n14702_), .A1(new_n14688_), .B0(new_n7625_), .Y(new_n14703_));
  AOI21X1  g12267(.A0(new_n9483_), .A1(new_n9837_), .B0(pi0832), .Y(new_n14704_));
  OAI21X1  g12268(.A0(new_n14501_), .A1(pi0701), .B0(new_n14685_), .Y(new_n14705_));
  OAI21X1  g12269(.A0(new_n2720_), .A1(pi0150), .B0(pi0832), .Y(new_n14706_));
  AOI21X1  g12270(.A0(new_n14705_), .A1(new_n2720_), .B0(new_n14706_), .Y(new_n14707_));
  AOI21X1  g12271(.A0(new_n14704_), .A1(new_n14703_), .B0(new_n14707_), .Y(po0307));
  OR2X1    g12272(.A(new_n5362_), .B(pi0745), .Y(new_n14709_));
  OAI21X1  g12273(.A0(new_n14501_), .A1(pi0723), .B0(new_n14709_), .Y(new_n14710_));
  OAI21X1  g12274(.A0(new_n2720_), .A1(pi0151), .B0(pi0832), .Y(new_n14711_));
  AOI21X1  g12275(.A0(new_n14710_), .A1(new_n2720_), .B0(new_n14711_), .Y(new_n14712_));
  AOI21X1  g12276(.A0(new_n14453_), .A1(new_n11821_), .B0(pi0039), .Y(new_n14713_));
  INVX1    g12277(.A(new_n14713_), .Y(new_n14714_));
  INVX1    g12278(.A(pi0745), .Y(new_n14715_));
  NAND3X1  g12279(.A(new_n11821_), .B(pi0947), .C(new_n14715_), .Y(new_n14716_));
  OAI21X1  g12280(.A0(new_n11821_), .A1(pi0151), .B0(new_n14716_), .Y(new_n14717_));
  NOR3X1   g12281(.A(new_n14513_), .B(new_n11955_), .C(pi0151), .Y(new_n14718_));
  OR2X1    g12282(.A(new_n14718_), .B(new_n11951_), .Y(new_n14719_));
  NOR3X1   g12283(.A(new_n11931_), .B(new_n11927_), .C(new_n5055_), .Y(new_n14720_));
  NOR3X1   g12284(.A(new_n14720_), .B(new_n10044_), .C(new_n3347_), .Y(new_n14721_));
  AOI21X1  g12285(.A0(new_n11945_), .A1(new_n10045_), .B0(new_n14721_), .Y(new_n14722_));
  INVX1    g12286(.A(new_n14580_), .Y(new_n14723_));
  AND2X1   g12287(.A(new_n11825_), .B(new_n3347_), .Y(new_n14724_));
  OR3X1    g12288(.A(new_n14724_), .B(new_n14723_), .C(new_n14560_), .Y(new_n14725_));
  AND2X1   g12289(.A(new_n14725_), .B(new_n2934_), .Y(new_n14726_));
  AOI22X1  g12290(.A0(new_n14726_), .A1(new_n14722_), .B0(new_n14719_), .B1(pi0215), .Y(new_n14727_));
  OR2X1    g12291(.A(new_n14727_), .B(new_n2933_), .Y(new_n14728_));
  NOR3X1   g12292(.A(new_n11936_), .B(new_n11879_), .C(new_n5055_), .Y(new_n14729_));
  OAI21X1  g12293(.A0(new_n14729_), .A1(new_n3347_), .B0(new_n14553_), .Y(new_n14730_));
  AOI21X1  g12294(.A0(new_n14730_), .A1(new_n14728_), .B0(pi0745), .Y(new_n14731_));
  INVX1    g12295(.A(new_n14527_), .Y(new_n14732_));
  AND2X1   g12296(.A(new_n14719_), .B(pi0215), .Y(new_n14733_));
  OAI21X1  g12297(.A0(new_n14724_), .A1(new_n14723_), .B0(new_n14722_), .Y(new_n14734_));
  NOR2X1   g12298(.A(new_n14734_), .B(new_n14543_), .Y(new_n14735_));
  OAI21X1  g12299(.A0(new_n14735_), .A1(new_n14733_), .B0(new_n14732_), .Y(new_n14736_));
  NAND2X1  g12300(.A(new_n14584_), .B(new_n2933_), .Y(new_n14737_));
  NOR2X1   g12301(.A(new_n14508_), .B(pi0151), .Y(new_n14738_));
  OAI21X1  g12302(.A0(new_n14738_), .A1(new_n14737_), .B0(pi0745), .Y(new_n14739_));
  AOI21X1  g12303(.A0(new_n14736_), .A1(pi0299), .B0(new_n14739_), .Y(new_n14740_));
  OR3X1    g12304(.A(new_n14740_), .B(new_n14731_), .C(new_n2939_), .Y(new_n14741_));
  OAI21X1  g12305(.A0(new_n14717_), .A1(new_n14714_), .B0(new_n14741_), .Y(new_n14742_));
  INVX1    g12306(.A(pi0723), .Y(new_n14743_));
  NOR2X1   g12307(.A(new_n12077_), .B(pi0151), .Y(new_n14744_));
  OAI21X1  g12308(.A0(new_n5362_), .A1(new_n14715_), .B0(new_n2939_), .Y(new_n14745_));
  OAI21X1  g12309(.A0(new_n14745_), .A1(new_n14669_), .B0(pi0038), .Y(new_n14746_));
  OAI21X1  g12310(.A0(new_n14746_), .A1(new_n14744_), .B0(new_n14743_), .Y(new_n14747_));
  AOI21X1  g12311(.A0(new_n14742_), .A1(new_n2979_), .B0(new_n14747_), .Y(new_n14748_));
  NAND2X1  g12312(.A(new_n11937_), .B(new_n14715_), .Y(new_n14749_));
  AND3X1   g12313(.A(new_n14749_), .B(new_n11958_), .C(new_n3347_), .Y(new_n14750_));
  NOR2X1   g12314(.A(new_n14529_), .B(new_n10045_), .Y(new_n14751_));
  INVX1    g12315(.A(new_n14751_), .Y(new_n14752_));
  OAI21X1  g12316(.A0(new_n14724_), .A1(new_n14752_), .B0(new_n14722_), .Y(new_n14753_));
  OR3X1    g12317(.A(new_n14753_), .B(new_n14511_), .C(pi0215), .Y(new_n14754_));
  NOR2X1   g12318(.A(new_n14513_), .B(new_n2934_), .Y(new_n14755_));
  AOI21X1  g12319(.A0(new_n14719_), .A1(new_n14755_), .B0(new_n2933_), .Y(new_n14756_));
  OAI21X1  g12320(.A0(new_n14525_), .A1(pi0299), .B0(new_n14715_), .Y(new_n14757_));
  AOI21X1  g12321(.A0(new_n14756_), .A1(new_n14754_), .B0(new_n14757_), .Y(new_n14758_));
  OAI21X1  g12322(.A0(new_n14758_), .A1(new_n14750_), .B0(pi0039), .Y(new_n14759_));
  AOI21X1  g12323(.A0(new_n14717_), .A1(new_n2939_), .B0(pi0038), .Y(new_n14760_));
  AOI22X1  g12324(.A0(new_n14709_), .A1(new_n12077_), .B0(new_n12831_), .B1(pi0151), .Y(new_n14761_));
  OAI21X1  g12325(.A0(new_n14761_), .A1(new_n2979_), .B0(pi0723), .Y(new_n14762_));
  AOI21X1  g12326(.A0(new_n14760_), .A1(new_n14759_), .B0(new_n14762_), .Y(new_n14763_));
  OAI21X1  g12327(.A0(new_n14763_), .A1(new_n14748_), .B0(new_n7625_), .Y(new_n14764_));
  AOI21X1  g12328(.A0(new_n9483_), .A1(new_n3347_), .B0(pi0832), .Y(new_n14765_));
  AOI21X1  g12329(.A0(new_n14765_), .A1(new_n14764_), .B0(new_n14712_), .Y(po0308));
  INVX1    g12330(.A(pi0759), .Y(new_n14767_));
  MX2X1    g12331(.A(new_n5055_), .B(new_n3193_), .S0(new_n11825_), .Y(new_n14768_));
  AOI21X1  g12332(.A0(new_n14768_), .A1(new_n10044_), .B0(pi0215), .Y(new_n14769_));
  INVX1    g12333(.A(new_n14542_), .Y(new_n14770_));
  OAI21X1  g12334(.A0(new_n14770_), .A1(new_n3193_), .B0(new_n14578_), .Y(new_n14771_));
  OAI21X1  g12335(.A0(new_n14771_), .A1(new_n14720_), .B0(new_n14769_), .Y(new_n14772_));
  OAI21X1  g12336(.A0(new_n11951_), .A1(pi0152), .B0(new_n14540_), .Y(new_n14773_));
  AND3X1   g12337(.A(new_n14773_), .B(new_n14772_), .C(pi0299), .Y(new_n14774_));
  NOR2X1   g12338(.A(new_n11933_), .B(pi0152), .Y(new_n14775_));
  AOI21X1  g12339(.A0(new_n11933_), .A1(new_n5362_), .B0(new_n2951_), .Y(new_n14776_));
  INVX1    g12340(.A(new_n14776_), .Y(new_n14777_));
  NOR2X1   g12341(.A(new_n14777_), .B(new_n14775_), .Y(new_n14778_));
  INVX1    g12342(.A(new_n11933_), .Y(new_n14779_));
  OAI21X1  g12343(.A0(new_n14779_), .A1(new_n5055_), .B0(new_n2952_), .Y(new_n14780_));
  OR2X1    g12344(.A(new_n14780_), .B(new_n14778_), .Y(new_n14781_));
  AOI21X1  g12345(.A0(new_n14768_), .A1(new_n2951_), .B0(pi0223), .Y(new_n14782_));
  INVX1    g12346(.A(new_n14551_), .Y(new_n14783_));
  NOR2X1   g12347(.A(new_n11878_), .B(pi0152), .Y(new_n14784_));
  OAI21X1  g12348(.A0(new_n11878_), .A1(pi0152), .B0(new_n14550_), .Y(new_n14785_));
  AND2X1   g12349(.A(new_n14785_), .B(new_n2933_), .Y(new_n14786_));
  OAI21X1  g12350(.A0(new_n14784_), .A1(new_n14783_), .B0(new_n14786_), .Y(new_n14787_));
  AOI21X1  g12351(.A0(new_n14782_), .A1(new_n14781_), .B0(new_n14787_), .Y(new_n14788_));
  OR3X1    g12352(.A(new_n14788_), .B(new_n14774_), .C(new_n14767_), .Y(new_n14789_));
  AOI22X1  g12353(.A0(new_n14579_), .A1(new_n5362_), .B0(new_n11825_), .B1(pi0152), .Y(new_n14790_));
  OAI21X1  g12354(.A0(new_n14453_), .A1(new_n14779_), .B0(new_n2952_), .Y(new_n14791_));
  OAI22X1  g12355(.A0(new_n14791_), .A1(new_n14775_), .B0(new_n14790_), .B1(new_n2952_), .Y(new_n14792_));
  OAI21X1  g12356(.A0(new_n14784_), .A1(new_n14783_), .B0(new_n2933_), .Y(new_n14793_));
  AOI21X1  g12357(.A0(new_n14792_), .A1(new_n2940_), .B0(new_n14793_), .Y(new_n14794_));
  OR4X1    g12358(.A(new_n14453_), .B(new_n11824_), .C(new_n10045_), .D(new_n2725_), .Y(new_n14795_));
  AND2X1   g12359(.A(new_n14769_), .B(new_n14795_), .Y(new_n14796_));
  NOR2X1   g12360(.A(new_n11951_), .B(new_n2934_), .Y(new_n14797_));
  NOR2X1   g12361(.A(new_n14797_), .B(new_n14453_), .Y(new_n14798_));
  OAI21X1  g12362(.A0(new_n14798_), .A1(new_n14773_), .B0(pi0299), .Y(new_n14799_));
  AOI21X1  g12363(.A0(new_n14796_), .A1(new_n14771_), .B0(new_n14799_), .Y(new_n14800_));
  OR3X1    g12364(.A(new_n14800_), .B(new_n14794_), .C(pi0759), .Y(new_n14801_));
  AND3X1   g12365(.A(new_n14801_), .B(new_n14789_), .C(pi0039), .Y(new_n14802_));
  NOR2X1   g12366(.A(new_n11821_), .B(pi0039), .Y(new_n14803_));
  AOI21X1  g12367(.A0(pi0947), .A1(pi0759), .B0(pi0039), .Y(new_n14804_));
  OAI22X1  g12368(.A0(new_n14804_), .A1(new_n14803_), .B0(new_n11821_), .B1(new_n3193_), .Y(new_n14805_));
  OAI21X1  g12369(.A0(new_n14805_), .A1(new_n14586_), .B0(new_n2979_), .Y(new_n14806_));
  INVX1    g12370(.A(pi0696), .Y(new_n14807_));
  OR2X1    g12371(.A(new_n12077_), .B(pi0152), .Y(new_n14808_));
  NOR4X1   g12372(.A(new_n14453_), .B(new_n2985_), .C(new_n2725_), .D(new_n2536_), .Y(new_n14809_));
  AOI21X1  g12373(.A0(new_n14809_), .A1(new_n14804_), .B0(new_n2979_), .Y(new_n14810_));
  AOI21X1  g12374(.A0(new_n14810_), .A1(new_n14808_), .B0(new_n14807_), .Y(new_n14811_));
  OAI21X1  g12375(.A0(new_n14806_), .A1(new_n14802_), .B0(new_n14811_), .Y(new_n14812_));
  INVX1    g12376(.A(new_n14511_), .Y(new_n14813_));
  AOI22X1  g12377(.A0(new_n14771_), .A1(new_n14813_), .B0(new_n11932_), .B1(pi0947), .Y(new_n14814_));
  MX2X1    g12378(.A(pi0947), .B(pi0152), .S0(new_n11825_), .Y(new_n14815_));
  OAI21X1  g12379(.A0(new_n14815_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n14816_));
  OR2X1    g12380(.A(new_n14527_), .B(new_n2933_), .Y(new_n14817_));
  AOI21X1  g12381(.A0(new_n14514_), .A1(pi0152), .B0(new_n14817_), .Y(new_n14818_));
  OAI21X1  g12382(.A0(new_n14816_), .A1(new_n14814_), .B0(new_n14818_), .Y(new_n14819_));
  AND2X1   g12383(.A(new_n14815_), .B(new_n2951_), .Y(new_n14820_));
  OAI21X1  g12384(.A0(new_n14820_), .A1(new_n14778_), .B0(new_n2940_), .Y(new_n14821_));
  AOI21X1  g12385(.A0(new_n14821_), .A1(new_n14786_), .B0(new_n14767_), .Y(new_n14822_));
  AOI21X1  g12386(.A0(new_n11957_), .A1(new_n11937_), .B0(pi0759), .Y(new_n14823_));
  AND2X1   g12387(.A(new_n14823_), .B(pi0152), .Y(new_n14824_));
  OR2X1    g12388(.A(new_n14824_), .B(new_n2939_), .Y(new_n14825_));
  AOI21X1  g12389(.A0(new_n14822_), .A1(new_n14819_), .B0(new_n14825_), .Y(new_n14826_));
  NAND2X1  g12390(.A(new_n14805_), .B(new_n2979_), .Y(new_n14827_));
  NAND2X1  g12391(.A(pi0947), .B(pi0759), .Y(new_n14828_));
  AOI21X1  g12392(.A0(new_n14828_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n14829_));
  OAI21X1  g12393(.A0(new_n12446_), .A1(pi0152), .B0(new_n14829_), .Y(new_n14830_));
  AND2X1   g12394(.A(new_n14830_), .B(new_n14807_), .Y(new_n14831_));
  OAI21X1  g12395(.A0(new_n14827_), .A1(new_n14826_), .B0(new_n14831_), .Y(new_n14832_));
  AOI21X1  g12396(.A0(new_n14832_), .A1(new_n14812_), .B0(new_n9483_), .Y(new_n14833_));
  OAI21X1  g12397(.A0(new_n7625_), .A1(pi0152), .B0(new_n12767_), .Y(new_n14834_));
  NAND2X1  g12398(.A(new_n14828_), .B(new_n2720_), .Y(new_n14835_));
  AOI21X1  g12399(.A0(new_n14453_), .A1(pi0696), .B0(new_n14835_), .Y(new_n14836_));
  OAI21X1  g12400(.A0(new_n2720_), .A1(pi0152), .B0(pi0832), .Y(new_n14837_));
  OAI22X1  g12401(.A0(new_n14837_), .A1(new_n14836_), .B0(new_n14834_), .B1(new_n14833_), .Y(po0309));
  AOI21X1  g12402(.A0(pi0947), .A1(pi0766), .B0(new_n2725_), .Y(new_n14839_));
  INVX1    g12403(.A(pi0700), .Y(new_n14840_));
  OR3X1    g12404(.A(pi0947), .B(new_n5277_), .C(new_n14840_), .Y(new_n14841_));
  OAI21X1  g12405(.A0(new_n2720_), .A1(new_n2924_), .B0(pi0832), .Y(new_n14842_));
  AOI21X1  g12406(.A0(new_n14841_), .A1(new_n14839_), .B0(new_n14842_), .Y(new_n14843_));
  INVX1    g12407(.A(pi0766), .Y(new_n14844_));
  AND3X1   g12408(.A(new_n11821_), .B(new_n14844_), .C(new_n2939_), .Y(new_n14845_));
  OAI22X1  g12409(.A0(new_n14845_), .A1(new_n14524_), .B0(new_n11821_), .B1(pi0153), .Y(new_n14846_));
  NOR2X1   g12410(.A(new_n11951_), .B(new_n2924_), .Y(new_n14847_));
  NOR3X1   g12411(.A(new_n14847_), .B(new_n11955_), .C(new_n2934_), .Y(new_n14848_));
  INVX1    g12412(.A(new_n14720_), .Y(new_n14849_));
  NOR2X1   g12413(.A(new_n10044_), .B(new_n2924_), .Y(new_n14850_));
  AOI22X1  g12414(.A0(new_n14850_), .A1(new_n14849_), .B0(new_n11945_), .B1(new_n10045_), .Y(new_n14851_));
  INVX1    g12415(.A(new_n14579_), .Y(new_n14852_));
  AND2X1   g12416(.A(new_n11825_), .B(new_n2924_), .Y(new_n14853_));
  NOR3X1   g12417(.A(new_n14853_), .B(new_n14529_), .C(new_n10045_), .Y(new_n14854_));
  AOI21X1  g12418(.A0(new_n14854_), .A1(new_n14852_), .B0(pi0215), .Y(new_n14855_));
  AOI21X1  g12419(.A0(new_n14855_), .A1(new_n14851_), .B0(new_n14848_), .Y(new_n14856_));
  OR2X1    g12420(.A(new_n14856_), .B(new_n2933_), .Y(new_n14857_));
  OAI21X1  g12421(.A0(new_n14729_), .A1(new_n2924_), .B0(new_n14553_), .Y(new_n14858_));
  AOI21X1  g12422(.A0(new_n14858_), .A1(new_n14857_), .B0(new_n14844_), .Y(new_n14859_));
  INVX1    g12423(.A(new_n14851_), .Y(new_n14860_));
  OAI22X1  g12424(.A0(new_n14853_), .A1(new_n14723_), .B0(new_n14542_), .B1(new_n10044_), .Y(new_n14861_));
  OAI21X1  g12425(.A0(new_n14861_), .A1(new_n14860_), .B0(new_n2934_), .Y(new_n14862_));
  OR3X1    g12426(.A(new_n14848_), .B(new_n11951_), .C(new_n2934_), .Y(new_n14863_));
  AND2X1   g12427(.A(new_n14863_), .B(new_n14732_), .Y(new_n14864_));
  AOI21X1  g12428(.A0(new_n14864_), .A1(new_n14862_), .B0(new_n2933_), .Y(new_n14865_));
  NOR2X1   g12429(.A(new_n14508_), .B(pi0153), .Y(new_n14866_));
  OAI21X1  g12430(.A0(new_n14866_), .A1(new_n14737_), .B0(new_n14844_), .Y(new_n14867_));
  OAI21X1  g12431(.A0(new_n14867_), .A1(new_n14865_), .B0(pi0039), .Y(new_n14868_));
  OAI22X1  g12432(.A0(new_n14868_), .A1(new_n14859_), .B0(new_n14846_), .B1(new_n14586_), .Y(new_n14869_));
  OAI21X1  g12433(.A0(new_n5362_), .A1(pi0766), .B0(new_n2939_), .Y(new_n14870_));
  OAI21X1  g12434(.A0(new_n14870_), .A1(new_n14669_), .B0(pi0038), .Y(new_n14871_));
  AOI21X1  g12435(.A0(new_n12771_), .A1(new_n2924_), .B0(new_n14871_), .Y(new_n14872_));
  AOI21X1  g12436(.A0(new_n14869_), .A1(new_n2979_), .B0(new_n14872_), .Y(new_n14873_));
  NOR3X1   g12437(.A(new_n14866_), .B(new_n14525_), .C(pi0299), .Y(new_n14874_));
  NOR4X1   g12438(.A(new_n14854_), .B(new_n14860_), .C(new_n14511_), .D(pi0215), .Y(new_n14875_));
  INVX1    g12439(.A(new_n14514_), .Y(new_n14876_));
  OAI21X1  g12440(.A0(new_n14847_), .A1(new_n14876_), .B0(pi0299), .Y(new_n14877_));
  OAI21X1  g12441(.A0(new_n14877_), .A1(new_n14875_), .B0(pi0766), .Y(new_n14878_));
  NOR2X1   g12442(.A(new_n14878_), .B(new_n14874_), .Y(new_n14879_));
  OR2X1    g12443(.A(pi0766), .B(pi0153), .Y(new_n14880_));
  OAI21X1  g12444(.A0(new_n14880_), .A1(new_n12444_), .B0(pi0039), .Y(new_n14881_));
  AND2X1   g12445(.A(new_n14846_), .B(new_n2979_), .Y(new_n14882_));
  OAI21X1  g12446(.A0(new_n14881_), .A1(new_n14879_), .B0(new_n14882_), .Y(new_n14883_));
  AOI21X1  g12447(.A0(new_n14839_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n14884_));
  OAI21X1  g12448(.A0(new_n12446_), .A1(new_n2924_), .B0(new_n14884_), .Y(new_n14885_));
  AND2X1   g12449(.A(new_n14885_), .B(new_n14840_), .Y(new_n14886_));
  AOI21X1  g12450(.A0(new_n14886_), .A1(new_n14883_), .B0(new_n14616_), .Y(new_n14887_));
  OAI21X1  g12451(.A0(new_n14873_), .A1(new_n14840_), .B0(new_n14887_), .Y(new_n14888_));
  AOI21X1  g12452(.A0(new_n14616_), .A1(new_n2924_), .B0(pi0057), .Y(new_n14889_));
  OAI21X1  g12453(.A0(new_n2924_), .A1(new_n2436_), .B0(new_n12767_), .Y(new_n14890_));
  AOI21X1  g12454(.A0(new_n14889_), .A1(new_n14888_), .B0(new_n14890_), .Y(new_n14891_));
  OR2X1    g12455(.A(new_n14891_), .B(new_n14843_), .Y(po0310));
  OAI22X1  g12456(.A0(new_n14501_), .A1(pi0704), .B0(new_n5362_), .B1(pi0742), .Y(new_n14893_));
  OAI21X1  g12457(.A0(new_n2720_), .A1(pi0154), .B0(pi0832), .Y(new_n14894_));
  AOI21X1  g12458(.A0(new_n14893_), .A1(new_n2720_), .B0(new_n14894_), .Y(new_n14895_));
  INVX1    g12459(.A(pi0704), .Y(new_n14896_));
  INVX1    g12460(.A(pi0742), .Y(new_n14897_));
  OR2X1    g12461(.A(new_n11821_), .B(pi0154), .Y(new_n14898_));
  AND2X1   g12462(.A(new_n14898_), .B(new_n14713_), .Y(new_n14899_));
  INVX1    g12463(.A(new_n14899_), .Y(new_n14900_));
  AOI21X1  g12464(.A0(new_n14585_), .A1(pi0154), .B0(new_n2939_), .Y(new_n14901_));
  OAI21X1  g12465(.A0(new_n14574_), .A1(pi0154), .B0(new_n14901_), .Y(new_n14902_));
  AOI21X1  g12466(.A0(new_n14902_), .A1(new_n14900_), .B0(pi0038), .Y(new_n14903_));
  OR2X1    g12467(.A(new_n12077_), .B(pi0154), .Y(new_n14904_));
  AND2X1   g12468(.A(new_n14904_), .B(new_n14591_), .Y(new_n14905_));
  OR3X1    g12469(.A(new_n14905_), .B(new_n14903_), .C(new_n14897_), .Y(new_n14906_));
  AND2X1   g12470(.A(new_n11821_), .B(new_n14547_), .Y(new_n14907_));
  INVX1    g12471(.A(new_n14907_), .Y(new_n14908_));
  OR2X1    g12472(.A(new_n14555_), .B(pi0154), .Y(new_n14909_));
  AOI21X1  g12473(.A0(new_n14603_), .A1(pi0154), .B0(new_n2939_), .Y(new_n14910_));
  AOI22X1  g12474(.A0(new_n14910_), .A1(new_n14909_), .B0(new_n14899_), .B1(new_n14908_), .Y(new_n14911_));
  AOI21X1  g12475(.A0(new_n14904_), .A1(new_n14569_), .B0(pi0742), .Y(new_n14912_));
  OAI21X1  g12476(.A0(new_n14911_), .A1(pi0038), .B0(new_n14912_), .Y(new_n14913_));
  AND3X1   g12477(.A(new_n14913_), .B(new_n14906_), .C(new_n14896_), .Y(new_n14914_));
  AND2X1   g12478(.A(new_n14898_), .B(new_n14524_), .Y(new_n14915_));
  AOI21X1  g12479(.A0(new_n14516_), .A1(new_n14507_), .B0(pi0154), .Y(new_n14916_));
  OAI21X1  g12480(.A0(new_n14534_), .A1(new_n3133_), .B0(pi0039), .Y(new_n14917_));
  NOR2X1   g12481(.A(new_n14917_), .B(new_n14916_), .Y(new_n14918_));
  OAI21X1  g12482(.A0(new_n14918_), .A1(new_n14915_), .B0(new_n2979_), .Y(new_n14919_));
  OAI22X1  g12483(.A0(new_n14519_), .A1(new_n13265_), .B0(new_n12446_), .B1(pi0154), .Y(new_n14920_));
  AND2X1   g12484(.A(new_n14920_), .B(new_n14897_), .Y(new_n14921_));
  OR2X1    g12485(.A(new_n14897_), .B(pi0154), .Y(new_n14922_));
  OAI21X1  g12486(.A0(new_n14922_), .A1(new_n12447_), .B0(pi0704), .Y(new_n14923_));
  AOI21X1  g12487(.A0(new_n14921_), .A1(new_n14919_), .B0(new_n14923_), .Y(new_n14924_));
  OR3X1    g12488(.A(new_n14924_), .B(new_n14914_), .C(new_n9483_), .Y(new_n14925_));
  AOI21X1  g12489(.A0(new_n9483_), .A1(new_n3133_), .B0(pi0832), .Y(new_n14926_));
  AOI21X1  g12490(.A0(new_n14926_), .A1(new_n14925_), .B0(new_n14895_), .Y(po0311));
  INVX1    g12491(.A(pi0757), .Y(new_n14928_));
  INVX1    g12492(.A(new_n14565_), .Y(new_n14929_));
  AOI21X1  g12493(.A0(new_n14929_), .A1(new_n2979_), .B0(new_n14569_), .Y(new_n14930_));
  NAND2X1  g12494(.A(new_n14930_), .B(new_n14928_), .Y(new_n14931_));
  AOI21X1  g12495(.A0(new_n14588_), .A1(new_n2979_), .B0(new_n14591_), .Y(new_n14932_));
  AOI21X1  g12496(.A0(new_n14932_), .A1(pi0757), .B0(pi0686), .Y(new_n14933_));
  AND2X1   g12497(.A(new_n14933_), .B(new_n14931_), .Y(new_n14934_));
  INVX1    g12498(.A(pi0686), .Y(new_n14935_));
  AND2X1   g12499(.A(new_n14536_), .B(new_n14523_), .Y(new_n14936_));
  AOI21X1  g12500(.A0(new_n14936_), .A1(new_n14928_), .B0(new_n14935_), .Y(new_n14937_));
  NOR3X1   g12501(.A(new_n14937_), .B(new_n14934_), .C(new_n9483_), .Y(new_n14938_));
  MX2X1    g12502(.A(new_n14568_), .B(new_n14558_), .S0(new_n2979_), .Y(new_n14939_));
  OR2X1    g12503(.A(new_n14939_), .B(pi0757), .Y(new_n14940_));
  AOI22X1  g12504(.A0(new_n14591_), .A1(new_n12077_), .B0(new_n14576_), .B1(new_n2979_), .Y(new_n14941_));
  AOI21X1  g12505(.A0(new_n14941_), .A1(pi0757), .B0(pi0686), .Y(new_n14942_));
  OAI21X1  g12506(.A0(new_n12447_), .A1(new_n14928_), .B0(pi0686), .Y(new_n14943_));
  AOI21X1  g12507(.A0(new_n14520_), .A1(new_n14928_), .B0(new_n14943_), .Y(new_n14944_));
  AOI21X1  g12508(.A0(new_n14942_), .A1(new_n14940_), .B0(new_n14944_), .Y(new_n14945_));
  NAND3X1  g12509(.A(new_n6489_), .B(new_n3103_), .C(new_n7449_), .Y(new_n14946_));
  OAI22X1  g12510(.A0(new_n14946_), .A1(new_n14945_), .B0(new_n14938_), .B1(new_n7449_), .Y(new_n14947_));
  OAI22X1  g12511(.A0(new_n14501_), .A1(pi0686), .B0(new_n5362_), .B1(pi0757), .Y(new_n14948_));
  OAI21X1  g12512(.A0(new_n2720_), .A1(pi0155), .B0(pi0832), .Y(new_n14949_));
  AOI21X1  g12513(.A0(new_n14948_), .A1(new_n2720_), .B0(new_n14949_), .Y(new_n14950_));
  AOI21X1  g12514(.A0(new_n14947_), .A1(new_n12767_), .B0(new_n14950_), .Y(po0312));
  OAI22X1  g12515(.A0(new_n14501_), .A1(pi0724), .B0(new_n5362_), .B1(pi0741), .Y(new_n14952_));
  OAI21X1  g12516(.A0(new_n2720_), .A1(pi0156), .B0(pi0832), .Y(new_n14953_));
  AOI21X1  g12517(.A0(new_n14952_), .A1(new_n2720_), .B0(new_n14953_), .Y(new_n14954_));
  INVX1    g12518(.A(pi0741), .Y(new_n14955_));
  INVX1    g12519(.A(pi0724), .Y(new_n14956_));
  OAI21X1  g12520(.A0(new_n14941_), .A1(new_n14955_), .B0(new_n14956_), .Y(new_n14957_));
  AOI21X1  g12521(.A0(new_n14939_), .A1(new_n14955_), .B0(new_n14957_), .Y(new_n14958_));
  AOI21X1  g12522(.A0(new_n12447_), .A1(pi0741), .B0(new_n14956_), .Y(new_n14959_));
  OAI21X1  g12523(.A0(new_n14520_), .A1(pi0741), .B0(new_n14959_), .Y(new_n14960_));
  NAND2X1  g12524(.A(new_n14960_), .B(new_n7625_), .Y(new_n14961_));
  OAI21X1  g12525(.A0(new_n14961_), .A1(new_n14958_), .B0(new_n8789_), .Y(new_n14962_));
  NOR2X1   g12526(.A(new_n14930_), .B(pi0741), .Y(new_n14963_));
  OAI21X1  g12527(.A0(new_n14932_), .A1(new_n14955_), .B0(new_n14956_), .Y(new_n14964_));
  NAND4X1  g12528(.A(new_n14536_), .B(new_n14523_), .C(new_n14955_), .D(pi0724), .Y(new_n14965_));
  OAI21X1  g12529(.A0(new_n14964_), .A1(new_n14963_), .B0(new_n14965_), .Y(new_n14966_));
  AND3X1   g12530(.A(new_n6489_), .B(new_n3103_), .C(pi0156), .Y(new_n14967_));
  AOI21X1  g12531(.A0(new_n14967_), .A1(new_n14966_), .B0(pi0832), .Y(new_n14968_));
  AOI21X1  g12532(.A0(new_n14968_), .A1(new_n14962_), .B0(new_n14954_), .Y(po0313));
  INVX1    g12533(.A(pi0760), .Y(new_n14970_));
  AND2X1   g12534(.A(pi0947), .B(new_n14970_), .Y(new_n14971_));
  INVX1    g12535(.A(new_n14971_), .Y(new_n14972_));
  OAI21X1  g12536(.A0(new_n14501_), .A1(pi0688), .B0(new_n14972_), .Y(new_n14973_));
  OAI21X1  g12537(.A0(new_n2720_), .A1(pi0157), .B0(pi0832), .Y(new_n14974_));
  AOI21X1  g12538(.A0(new_n14973_), .A1(new_n2720_), .B0(new_n14974_), .Y(new_n14975_));
  AOI21X1  g12539(.A0(new_n14972_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n14976_));
  OAI21X1  g12540(.A0(new_n12446_), .A1(new_n9968_), .B0(new_n14976_), .Y(new_n14977_));
  AND2X1   g12541(.A(pi0299), .B(new_n9968_), .Y(new_n14978_));
  OAI22X1  g12542(.A0(new_n14532_), .A1(new_n14978_), .B0(new_n14515_), .B1(pi0157), .Y(new_n14979_));
  OAI21X1  g12543(.A0(new_n11936_), .A1(new_n11879_), .B0(new_n9968_), .Y(new_n14980_));
  AOI21X1  g12544(.A0(new_n14980_), .A1(new_n14526_), .B0(pi0760), .Y(new_n14981_));
  OR2X1    g12545(.A(new_n14970_), .B(pi0157), .Y(new_n14982_));
  OAI21X1  g12546(.A0(new_n14982_), .A1(new_n12444_), .B0(pi0039), .Y(new_n14983_));
  AOI21X1  g12547(.A0(new_n14981_), .A1(new_n14979_), .B0(new_n14983_), .Y(new_n14984_));
  AOI21X1  g12548(.A0(new_n14971_), .A1(new_n11821_), .B0(pi0039), .Y(new_n14985_));
  OAI21X1  g12549(.A0(new_n11821_), .A1(pi0157), .B0(new_n14985_), .Y(new_n14986_));
  NAND2X1  g12550(.A(new_n14986_), .B(new_n2979_), .Y(new_n14987_));
  OAI21X1  g12551(.A0(new_n14987_), .A1(new_n14984_), .B0(new_n14977_), .Y(new_n14988_));
  AND2X1   g12552(.A(new_n14988_), .B(pi0688), .Y(new_n14989_));
  NOR4X1   g12553(.A(new_n14554_), .B(new_n14553_), .C(new_n14546_), .D(pi0760), .Y(new_n14990_));
  OR2X1    g12554(.A(new_n14990_), .B(pi0157), .Y(new_n14991_));
  AOI21X1  g12555(.A0(new_n14574_), .A1(pi0760), .B0(new_n14991_), .Y(new_n14992_));
  AND3X1   g12556(.A(new_n14563_), .B(new_n14559_), .C(new_n14970_), .Y(new_n14993_));
  OAI21X1  g12557(.A0(new_n14585_), .A1(new_n14970_), .B0(pi0157), .Y(new_n14994_));
  OAI21X1  g12558(.A0(new_n14994_), .A1(new_n14993_), .B0(pi0039), .Y(new_n14995_));
  OAI22X1  g12559(.A0(new_n14995_), .A1(new_n14992_), .B0(new_n14986_), .B1(new_n14586_), .Y(new_n14996_));
  INVX1    g12560(.A(pi0688), .Y(new_n14997_));
  NOR2X1   g12561(.A(new_n12077_), .B(pi0157), .Y(new_n14998_));
  OAI21X1  g12562(.A0(new_n5362_), .A1(new_n14970_), .B0(new_n2939_), .Y(new_n14999_));
  OAI21X1  g12563(.A0(new_n14999_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15000_));
  OAI21X1  g12564(.A0(new_n15000_), .A1(new_n14998_), .B0(new_n14997_), .Y(new_n15001_));
  AOI21X1  g12565(.A0(new_n14996_), .A1(new_n2979_), .B0(new_n15001_), .Y(new_n15002_));
  OAI21X1  g12566(.A0(new_n15002_), .A1(new_n14989_), .B0(new_n7625_), .Y(new_n15003_));
  AOI21X1  g12567(.A0(new_n9483_), .A1(new_n9968_), .B0(pi0832), .Y(new_n15004_));
  AOI21X1  g12568(.A0(new_n15004_), .A1(new_n15003_), .B0(new_n14975_), .Y(po0314));
  INVX1    g12569(.A(pi0753), .Y(new_n15006_));
  OAI21X1  g12570(.A0(new_n14533_), .A1(new_n7094_), .B0(new_n15006_), .Y(new_n15007_));
  AOI21X1  g12571(.A0(new_n14677_), .A1(new_n7094_), .B0(new_n15007_), .Y(new_n15008_));
  NOR3X1   g12572(.A(new_n12444_), .B(new_n15006_), .C(pi0158), .Y(new_n15009_));
  OAI21X1  g12573(.A0(new_n15009_), .A1(new_n15008_), .B0(pi0039), .Y(new_n15010_));
  MX2X1    g12574(.A(new_n7094_), .B(new_n15006_), .S0(new_n11821_), .Y(new_n15011_));
  AOI21X1  g12575(.A0(new_n15011_), .A1(new_n14505_), .B0(pi0038), .Y(new_n15012_));
  OR2X1    g12576(.A(new_n5362_), .B(pi0753), .Y(new_n15013_));
  AOI22X1  g12577(.A0(new_n15013_), .A1(new_n12077_), .B0(new_n12831_), .B1(pi0158), .Y(new_n15014_));
  OAI21X1  g12578(.A0(new_n15014_), .A1(new_n2979_), .B0(pi0702), .Y(new_n15015_));
  AOI21X1  g12579(.A0(new_n15012_), .A1(new_n15010_), .B0(new_n15015_), .Y(new_n15016_));
  OAI21X1  g12580(.A0(new_n14585_), .A1(new_n7094_), .B0(pi0753), .Y(new_n15017_));
  AOI21X1  g12581(.A0(new_n14574_), .A1(new_n7094_), .B0(new_n15017_), .Y(new_n15018_));
  OAI21X1  g12582(.A0(new_n14603_), .A1(new_n7094_), .B0(new_n15006_), .Y(new_n15019_));
  AOI21X1  g12583(.A0(new_n14555_), .A1(new_n7094_), .B0(new_n15019_), .Y(new_n15020_));
  OAI21X1  g12584(.A0(new_n15020_), .A1(new_n15018_), .B0(pi0039), .Y(new_n15021_));
  NAND3X1  g12585(.A(new_n15013_), .B(new_n14501_), .C(new_n11821_), .Y(new_n15022_));
  AOI21X1  g12586(.A0(new_n11822_), .A1(pi0158), .B0(pi0039), .Y(new_n15023_));
  AOI21X1  g12587(.A0(new_n15023_), .A1(new_n15022_), .B0(pi0038), .Y(new_n15024_));
  INVX1    g12588(.A(pi0702), .Y(new_n15025_));
  NOR2X1   g12589(.A(new_n12077_), .B(pi0158), .Y(new_n15026_));
  OAI21X1  g12590(.A0(new_n5362_), .A1(new_n15006_), .B0(new_n2939_), .Y(new_n15027_));
  OAI21X1  g12591(.A0(new_n15027_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15028_));
  OAI21X1  g12592(.A0(new_n15028_), .A1(new_n15026_), .B0(new_n15025_), .Y(new_n15029_));
  AOI21X1  g12593(.A0(new_n15024_), .A1(new_n15021_), .B0(new_n15029_), .Y(new_n15030_));
  OAI21X1  g12594(.A0(new_n15030_), .A1(new_n15016_), .B0(new_n7625_), .Y(new_n15031_));
  AOI21X1  g12595(.A0(new_n9483_), .A1(new_n7094_), .B0(pi0832), .Y(new_n15032_));
  OAI21X1  g12596(.A0(new_n14501_), .A1(pi0702), .B0(new_n15013_), .Y(new_n15033_));
  OAI21X1  g12597(.A0(new_n2720_), .A1(pi0158), .B0(pi0832), .Y(new_n15034_));
  AOI21X1  g12598(.A0(new_n15033_), .A1(new_n2720_), .B0(new_n15034_), .Y(new_n15035_));
  AOI21X1  g12599(.A0(new_n15032_), .A1(new_n15031_), .B0(new_n15035_), .Y(po0315));
  INVX1    g12600(.A(pi0754), .Y(new_n15037_));
  OAI21X1  g12601(.A0(new_n14533_), .A1(new_n7377_), .B0(new_n15037_), .Y(new_n15038_));
  AOI21X1  g12602(.A0(new_n14677_), .A1(new_n7377_), .B0(new_n15038_), .Y(new_n15039_));
  NOR3X1   g12603(.A(new_n12444_), .B(new_n15037_), .C(pi0159), .Y(new_n15040_));
  OAI21X1  g12604(.A0(new_n15040_), .A1(new_n15039_), .B0(pi0039), .Y(new_n15041_));
  MX2X1    g12605(.A(new_n7377_), .B(new_n15037_), .S0(new_n11821_), .Y(new_n15042_));
  AOI21X1  g12606(.A0(new_n15042_), .A1(new_n14505_), .B0(pi0038), .Y(new_n15043_));
  OR2X1    g12607(.A(new_n5362_), .B(pi0754), .Y(new_n15044_));
  AOI22X1  g12608(.A0(new_n15044_), .A1(new_n12077_), .B0(new_n12831_), .B1(pi0159), .Y(new_n15045_));
  OAI21X1  g12609(.A0(new_n15045_), .A1(new_n2979_), .B0(pi0709), .Y(new_n15046_));
  AOI21X1  g12610(.A0(new_n15043_), .A1(new_n15041_), .B0(new_n15046_), .Y(new_n15047_));
  OAI21X1  g12611(.A0(new_n14585_), .A1(new_n7377_), .B0(pi0754), .Y(new_n15048_));
  AOI21X1  g12612(.A0(new_n14574_), .A1(new_n7377_), .B0(new_n15048_), .Y(new_n15049_));
  OAI21X1  g12613(.A0(new_n14603_), .A1(new_n7377_), .B0(new_n15037_), .Y(new_n15050_));
  AOI21X1  g12614(.A0(new_n14555_), .A1(new_n7377_), .B0(new_n15050_), .Y(new_n15051_));
  OAI21X1  g12615(.A0(new_n15051_), .A1(new_n15049_), .B0(pi0039), .Y(new_n15052_));
  NAND3X1  g12616(.A(new_n15044_), .B(new_n14501_), .C(new_n11821_), .Y(new_n15053_));
  AOI21X1  g12617(.A0(new_n11822_), .A1(pi0159), .B0(pi0039), .Y(new_n15054_));
  AOI21X1  g12618(.A0(new_n15054_), .A1(new_n15053_), .B0(pi0038), .Y(new_n15055_));
  INVX1    g12619(.A(pi0709), .Y(new_n15056_));
  NOR2X1   g12620(.A(new_n12077_), .B(pi0159), .Y(new_n15057_));
  OAI21X1  g12621(.A0(new_n5362_), .A1(new_n15037_), .B0(new_n2939_), .Y(new_n15058_));
  OAI21X1  g12622(.A0(new_n15058_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15059_));
  OAI21X1  g12623(.A0(new_n15059_), .A1(new_n15057_), .B0(new_n15056_), .Y(new_n15060_));
  AOI21X1  g12624(.A0(new_n15055_), .A1(new_n15052_), .B0(new_n15060_), .Y(new_n15061_));
  OAI21X1  g12625(.A0(new_n15061_), .A1(new_n15047_), .B0(new_n7625_), .Y(new_n15062_));
  AOI21X1  g12626(.A0(new_n9483_), .A1(new_n7377_), .B0(pi0832), .Y(new_n15063_));
  OAI21X1  g12627(.A0(new_n14501_), .A1(pi0709), .B0(new_n15044_), .Y(new_n15064_));
  OAI21X1  g12628(.A0(new_n2720_), .A1(pi0159), .B0(pi0832), .Y(new_n15065_));
  AOI21X1  g12629(.A0(new_n15064_), .A1(new_n2720_), .B0(new_n15065_), .Y(new_n15066_));
  AOI21X1  g12630(.A0(new_n15063_), .A1(new_n15062_), .B0(new_n15066_), .Y(po0316));
  INVX1    g12631(.A(pi0756), .Y(new_n15068_));
  AND2X1   g12632(.A(pi0947), .B(new_n15068_), .Y(new_n15069_));
  INVX1    g12633(.A(new_n15069_), .Y(new_n15070_));
  OAI21X1  g12634(.A0(new_n14501_), .A1(pi0734), .B0(new_n15070_), .Y(new_n15071_));
  OAI21X1  g12635(.A0(new_n2720_), .A1(pi0160), .B0(pi0832), .Y(new_n15072_));
  AOI21X1  g12636(.A0(new_n15071_), .A1(new_n2720_), .B0(new_n15072_), .Y(new_n15073_));
  AOI21X1  g12637(.A0(new_n15070_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n15074_));
  OAI21X1  g12638(.A0(new_n12446_), .A1(new_n8850_), .B0(new_n15074_), .Y(new_n15075_));
  AOI21X1  g12639(.A0(new_n14617_), .A1(pi0160), .B0(new_n2933_), .Y(new_n15076_));
  OAI21X1  g12640(.A0(new_n14515_), .A1(pi0160), .B0(new_n15076_), .Y(new_n15077_));
  OAI21X1  g12641(.A0(new_n11936_), .A1(new_n11879_), .B0(new_n8850_), .Y(new_n15078_));
  AOI21X1  g12642(.A0(new_n15078_), .A1(new_n14526_), .B0(pi0756), .Y(new_n15079_));
  OR2X1    g12643(.A(new_n15068_), .B(pi0160), .Y(new_n15080_));
  OAI21X1  g12644(.A0(new_n15080_), .A1(new_n12444_), .B0(pi0039), .Y(new_n15081_));
  AOI21X1  g12645(.A0(new_n15079_), .A1(new_n15077_), .B0(new_n15081_), .Y(new_n15082_));
  AOI21X1  g12646(.A0(new_n15069_), .A1(new_n11821_), .B0(pi0039), .Y(new_n15083_));
  OAI21X1  g12647(.A0(new_n11821_), .A1(pi0160), .B0(new_n15083_), .Y(new_n15084_));
  NAND2X1  g12648(.A(new_n15084_), .B(new_n2979_), .Y(new_n15085_));
  OAI21X1  g12649(.A0(new_n15085_), .A1(new_n15082_), .B0(new_n15075_), .Y(new_n15086_));
  AND2X1   g12650(.A(new_n15086_), .B(pi0734), .Y(new_n15087_));
  OAI21X1  g12651(.A0(new_n14603_), .A1(new_n8850_), .B0(new_n15068_), .Y(new_n15088_));
  AOI21X1  g12652(.A0(new_n14555_), .A1(new_n8850_), .B0(new_n15088_), .Y(new_n15089_));
  NOR3X1   g12653(.A(new_n14572_), .B(new_n2933_), .C(pi0160), .Y(new_n15090_));
  AND2X1   g12654(.A(new_n14573_), .B(pi0756), .Y(new_n15091_));
  OAI21X1  g12655(.A0(new_n14600_), .A1(new_n8850_), .B0(new_n15091_), .Y(new_n15092_));
  OAI21X1  g12656(.A0(new_n15092_), .A1(new_n15090_), .B0(pi0039), .Y(new_n15093_));
  OAI22X1  g12657(.A0(new_n15093_), .A1(new_n15089_), .B0(new_n15084_), .B1(new_n14586_), .Y(new_n15094_));
  INVX1    g12658(.A(pi0734), .Y(new_n15095_));
  NOR2X1   g12659(.A(new_n12077_), .B(pi0160), .Y(new_n15096_));
  OAI21X1  g12660(.A0(new_n5362_), .A1(new_n15068_), .B0(new_n2939_), .Y(new_n15097_));
  OAI21X1  g12661(.A0(new_n15097_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15098_));
  OAI21X1  g12662(.A0(new_n15098_), .A1(new_n15096_), .B0(new_n15095_), .Y(new_n15099_));
  AOI21X1  g12663(.A0(new_n15094_), .A1(new_n2979_), .B0(new_n15099_), .Y(new_n15100_));
  OAI21X1  g12664(.A0(new_n15100_), .A1(new_n15087_), .B0(new_n7625_), .Y(new_n15101_));
  AOI21X1  g12665(.A0(new_n9483_), .A1(new_n8850_), .B0(pi0832), .Y(new_n15102_));
  AOI21X1  g12666(.A0(new_n15102_), .A1(new_n15101_), .B0(new_n15073_), .Y(po0317));
  MX2X1    g12667(.A(new_n5055_), .B(new_n4611_), .S0(new_n11825_), .Y(new_n15104_));
  AOI21X1  g12668(.A0(new_n15104_), .A1(new_n10044_), .B0(pi0215), .Y(new_n15105_));
  OAI21X1  g12669(.A0(new_n14770_), .A1(new_n4611_), .B0(new_n14578_), .Y(new_n15106_));
  OAI21X1  g12670(.A0(new_n15106_), .A1(new_n14720_), .B0(new_n15105_), .Y(new_n15107_));
  OAI21X1  g12671(.A0(new_n11951_), .A1(pi0161), .B0(new_n14540_), .Y(new_n15108_));
  AND3X1   g12672(.A(new_n15108_), .B(new_n15107_), .C(pi0299), .Y(new_n15109_));
  NOR2X1   g12673(.A(new_n11933_), .B(pi0161), .Y(new_n15110_));
  NOR2X1   g12674(.A(new_n15110_), .B(new_n14777_), .Y(new_n15111_));
  OR2X1    g12675(.A(new_n15111_), .B(new_n14780_), .Y(new_n15112_));
  AOI21X1  g12676(.A0(new_n15104_), .A1(new_n2951_), .B0(pi0223), .Y(new_n15113_));
  NOR2X1   g12677(.A(new_n11878_), .B(pi0161), .Y(new_n15114_));
  OAI21X1  g12678(.A0(new_n11878_), .A1(pi0161), .B0(new_n14550_), .Y(new_n15115_));
  AND2X1   g12679(.A(new_n15115_), .B(new_n2933_), .Y(new_n15116_));
  OAI21X1  g12680(.A0(new_n15114_), .A1(new_n14783_), .B0(new_n15116_), .Y(new_n15117_));
  AOI21X1  g12681(.A0(new_n15113_), .A1(new_n15112_), .B0(new_n15117_), .Y(new_n15118_));
  OR3X1    g12682(.A(new_n15118_), .B(new_n15109_), .C(new_n13836_), .Y(new_n15119_));
  AOI22X1  g12683(.A0(new_n14579_), .A1(new_n5362_), .B0(new_n11825_), .B1(pi0161), .Y(new_n15120_));
  OAI22X1  g12684(.A0(new_n15120_), .A1(new_n2952_), .B0(new_n15110_), .B1(new_n14791_), .Y(new_n15121_));
  OAI21X1  g12685(.A0(new_n15114_), .A1(new_n14783_), .B0(new_n2933_), .Y(new_n15122_));
  AOI21X1  g12686(.A0(new_n15121_), .A1(new_n2940_), .B0(new_n15122_), .Y(new_n15123_));
  AND2X1   g12687(.A(new_n15105_), .B(new_n14795_), .Y(new_n15124_));
  OAI21X1  g12688(.A0(new_n15108_), .A1(new_n14798_), .B0(pi0299), .Y(new_n15125_));
  AOI21X1  g12689(.A0(new_n15124_), .A1(new_n15106_), .B0(new_n15125_), .Y(new_n15126_));
  OR3X1    g12690(.A(new_n15126_), .B(new_n15123_), .C(pi0758), .Y(new_n15127_));
  AND3X1   g12691(.A(new_n15127_), .B(new_n15119_), .C(pi0039), .Y(new_n15128_));
  AND2X1   g12692(.A(pi0947), .B(pi0758), .Y(new_n15129_));
  INVX1    g12693(.A(new_n15129_), .Y(new_n15130_));
  AOI21X1  g12694(.A0(new_n11822_), .A1(pi0161), .B0(pi0039), .Y(new_n15131_));
  OAI21X1  g12695(.A0(new_n15130_), .A1(new_n11822_), .B0(new_n15131_), .Y(new_n15132_));
  OAI21X1  g12696(.A0(new_n15132_), .A1(new_n14586_), .B0(new_n2979_), .Y(new_n15133_));
  OR2X1    g12697(.A(new_n12077_), .B(pi0161), .Y(new_n15134_));
  AOI21X1  g12698(.A0(pi0947), .A1(pi0758), .B0(pi0039), .Y(new_n15135_));
  AOI21X1  g12699(.A0(new_n15135_), .A1(new_n14809_), .B0(new_n2979_), .Y(new_n15136_));
  AOI21X1  g12700(.A0(new_n15136_), .A1(new_n15134_), .B0(new_n13832_), .Y(new_n15137_));
  OAI21X1  g12701(.A0(new_n15133_), .A1(new_n15128_), .B0(new_n15137_), .Y(new_n15138_));
  AOI22X1  g12702(.A0(new_n15106_), .A1(new_n14813_), .B0(new_n11932_), .B1(pi0947), .Y(new_n15139_));
  MX2X1    g12703(.A(pi0947), .B(pi0161), .S0(new_n11825_), .Y(new_n15140_));
  OAI21X1  g12704(.A0(new_n15140_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n15141_));
  AOI21X1  g12705(.A0(new_n14514_), .A1(pi0161), .B0(new_n14817_), .Y(new_n15142_));
  OAI21X1  g12706(.A0(new_n15141_), .A1(new_n15139_), .B0(new_n15142_), .Y(new_n15143_));
  AND2X1   g12707(.A(new_n15140_), .B(new_n2951_), .Y(new_n15144_));
  OAI21X1  g12708(.A0(new_n15144_), .A1(new_n15111_), .B0(new_n2940_), .Y(new_n15145_));
  AOI21X1  g12709(.A0(new_n15145_), .A1(new_n15116_), .B0(new_n13836_), .Y(new_n15146_));
  AND2X1   g12710(.A(new_n13833_), .B(pi0161), .Y(new_n15147_));
  OR2X1    g12711(.A(new_n15147_), .B(new_n2939_), .Y(new_n15148_));
  AOI21X1  g12712(.A0(new_n15146_), .A1(new_n15143_), .B0(new_n15148_), .Y(new_n15149_));
  NAND2X1  g12713(.A(new_n15132_), .B(new_n2979_), .Y(new_n15150_));
  AOI21X1  g12714(.A0(new_n15130_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n15151_));
  OAI21X1  g12715(.A0(new_n12446_), .A1(pi0161), .B0(new_n15151_), .Y(new_n15152_));
  AND2X1   g12716(.A(new_n15152_), .B(new_n13832_), .Y(new_n15153_));
  OAI21X1  g12717(.A0(new_n15150_), .A1(new_n15149_), .B0(new_n15153_), .Y(new_n15154_));
  AOI21X1  g12718(.A0(new_n15154_), .A1(new_n15138_), .B0(new_n9483_), .Y(new_n15155_));
  OAI21X1  g12719(.A0(new_n7625_), .A1(pi0161), .B0(new_n12767_), .Y(new_n15156_));
  OAI21X1  g12720(.A0(new_n5362_), .A1(new_n13836_), .B0(new_n2720_), .Y(new_n15157_));
  AOI21X1  g12721(.A0(new_n14453_), .A1(pi0736), .B0(new_n15157_), .Y(new_n15158_));
  OAI21X1  g12722(.A0(new_n2720_), .A1(pi0161), .B0(pi0832), .Y(new_n15159_));
  OAI22X1  g12723(.A0(new_n15159_), .A1(new_n15158_), .B0(new_n15156_), .B1(new_n15155_), .Y(po0318));
  AND2X1   g12724(.A(pi0947), .B(new_n11772_), .Y(new_n15161_));
  INVX1    g12725(.A(new_n15161_), .Y(new_n15162_));
  AOI21X1  g12726(.A0(new_n15162_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n15163_));
  OAI21X1  g12727(.A0(new_n12446_), .A1(new_n7306_), .B0(new_n15163_), .Y(new_n15164_));
  OAI21X1  g12728(.A0(new_n11958_), .A1(new_n11772_), .B0(new_n7306_), .Y(new_n15165_));
  AOI21X1  g12729(.A0(new_n14516_), .A1(new_n11772_), .B0(new_n15165_), .Y(new_n15166_));
  AND2X1   g12730(.A(pi0299), .B(pi0162), .Y(new_n15167_));
  AOI21X1  g12731(.A0(new_n14617_), .A1(new_n15167_), .B0(new_n14506_), .Y(new_n15168_));
  OAI21X1  g12732(.A0(new_n15168_), .A1(pi0761), .B0(pi0039), .Y(new_n15169_));
  AOI21X1  g12733(.A0(new_n15161_), .A1(new_n11821_), .B0(pi0039), .Y(new_n15170_));
  OAI21X1  g12734(.A0(new_n11821_), .A1(pi0162), .B0(new_n15170_), .Y(new_n15171_));
  AND2X1   g12735(.A(new_n15171_), .B(new_n2979_), .Y(new_n15172_));
  OAI21X1  g12736(.A0(new_n15169_), .A1(new_n15166_), .B0(new_n15172_), .Y(new_n15173_));
  AOI21X1  g12737(.A0(new_n15173_), .A1(new_n15164_), .B0(new_n11771_), .Y(new_n15174_));
  INVX1    g12738(.A(new_n15167_), .Y(new_n15175_));
  OAI21X1  g12739(.A0(new_n14600_), .A1(new_n7306_), .B0(pi0761), .Y(new_n15176_));
  AOI21X1  g12740(.A0(new_n14574_), .A1(new_n15175_), .B0(new_n15176_), .Y(new_n15177_));
  NOR4X1   g12741(.A(new_n14554_), .B(new_n14553_), .C(new_n14546_), .D(pi0162), .Y(new_n15178_));
  OAI21X1  g12742(.A0(new_n14603_), .A1(new_n7306_), .B0(new_n11772_), .Y(new_n15179_));
  OAI21X1  g12743(.A0(new_n15179_), .A1(new_n15178_), .B0(pi0039), .Y(new_n15180_));
  OAI22X1  g12744(.A0(new_n15180_), .A1(new_n15177_), .B0(new_n15171_), .B1(new_n14586_), .Y(new_n15181_));
  NOR2X1   g12745(.A(new_n12077_), .B(pi0162), .Y(new_n15182_));
  OAI21X1  g12746(.A0(new_n5362_), .A1(new_n11772_), .B0(new_n2939_), .Y(new_n15183_));
  OAI21X1  g12747(.A0(new_n15183_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15184_));
  OAI21X1  g12748(.A0(new_n15184_), .A1(new_n15182_), .B0(new_n11771_), .Y(new_n15185_));
  AOI21X1  g12749(.A0(new_n15181_), .A1(new_n2979_), .B0(new_n15185_), .Y(new_n15186_));
  OAI21X1  g12750(.A0(new_n15186_), .A1(new_n15174_), .B0(new_n7625_), .Y(new_n15187_));
  AOI21X1  g12751(.A0(new_n9483_), .A1(new_n7306_), .B0(pi0832), .Y(new_n15188_));
  OAI21X1  g12752(.A0(new_n14501_), .A1(pi0738), .B0(new_n15162_), .Y(new_n15189_));
  OAI21X1  g12753(.A0(new_n2720_), .A1(pi0162), .B0(pi0832), .Y(new_n15190_));
  AOI21X1  g12754(.A0(new_n15189_), .A1(new_n2720_), .B0(new_n15190_), .Y(new_n15191_));
  AOI21X1  g12755(.A0(new_n15188_), .A1(new_n15187_), .B0(new_n15191_), .Y(po0319));
  INVX1    g12756(.A(pi0777), .Y(new_n15193_));
  AND2X1   g12757(.A(pi0947), .B(new_n15193_), .Y(new_n15194_));
  INVX1    g12758(.A(new_n15194_), .Y(new_n15195_));
  OAI21X1  g12759(.A0(new_n14501_), .A1(pi0737), .B0(new_n15195_), .Y(new_n15196_));
  OAI21X1  g12760(.A0(new_n2720_), .A1(pi0163), .B0(pi0832), .Y(new_n15197_));
  AOI21X1  g12761(.A0(new_n15196_), .A1(new_n2720_), .B0(new_n15197_), .Y(new_n15198_));
  AOI21X1  g12762(.A0(new_n15195_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n15199_));
  OAI21X1  g12763(.A0(new_n12446_), .A1(new_n8623_), .B0(new_n15199_), .Y(new_n15200_));
  AND2X1   g12764(.A(pi0299), .B(new_n8623_), .Y(new_n15201_));
  OAI22X1  g12765(.A0(new_n14532_), .A1(new_n15201_), .B0(new_n14515_), .B1(pi0163), .Y(new_n15202_));
  OAI21X1  g12766(.A0(new_n11936_), .A1(new_n11879_), .B0(new_n8623_), .Y(new_n15203_));
  AOI21X1  g12767(.A0(new_n15203_), .A1(new_n14526_), .B0(pi0777), .Y(new_n15204_));
  OR2X1    g12768(.A(new_n15193_), .B(pi0163), .Y(new_n15205_));
  OAI21X1  g12769(.A0(new_n15205_), .A1(new_n12444_), .B0(pi0039), .Y(new_n15206_));
  AOI21X1  g12770(.A0(new_n15204_), .A1(new_n15202_), .B0(new_n15206_), .Y(new_n15207_));
  AOI21X1  g12771(.A0(new_n15194_), .A1(new_n11821_), .B0(pi0039), .Y(new_n15208_));
  OAI21X1  g12772(.A0(new_n11821_), .A1(pi0163), .B0(new_n15208_), .Y(new_n15209_));
  NAND2X1  g12773(.A(new_n15209_), .B(new_n2979_), .Y(new_n15210_));
  OAI21X1  g12774(.A0(new_n15210_), .A1(new_n15207_), .B0(new_n15200_), .Y(new_n15211_));
  AND2X1   g12775(.A(new_n15211_), .B(pi0737), .Y(new_n15212_));
  OAI21X1  g12776(.A0(new_n14603_), .A1(new_n8623_), .B0(new_n15193_), .Y(new_n15213_));
  AOI21X1  g12777(.A0(new_n14555_), .A1(new_n8623_), .B0(new_n15213_), .Y(new_n15214_));
  NOR3X1   g12778(.A(new_n14572_), .B(new_n2933_), .C(pi0163), .Y(new_n15215_));
  AND2X1   g12779(.A(new_n14573_), .B(pi0777), .Y(new_n15216_));
  OAI21X1  g12780(.A0(new_n14600_), .A1(new_n8623_), .B0(new_n15216_), .Y(new_n15217_));
  OAI21X1  g12781(.A0(new_n15217_), .A1(new_n15215_), .B0(pi0039), .Y(new_n15218_));
  OAI22X1  g12782(.A0(new_n15218_), .A1(new_n15214_), .B0(new_n15209_), .B1(new_n14586_), .Y(new_n15219_));
  INVX1    g12783(.A(pi0737), .Y(new_n15220_));
  NOR2X1   g12784(.A(new_n12077_), .B(pi0163), .Y(new_n15221_));
  OAI21X1  g12785(.A0(new_n5362_), .A1(new_n15193_), .B0(new_n2939_), .Y(new_n15222_));
  OAI21X1  g12786(.A0(new_n15222_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15223_));
  OAI21X1  g12787(.A0(new_n15223_), .A1(new_n15221_), .B0(new_n15220_), .Y(new_n15224_));
  AOI21X1  g12788(.A0(new_n15219_), .A1(new_n2979_), .B0(new_n15224_), .Y(new_n15225_));
  OAI21X1  g12789(.A0(new_n15225_), .A1(new_n15212_), .B0(new_n7625_), .Y(new_n15226_));
  AOI21X1  g12790(.A0(new_n9483_), .A1(new_n8623_), .B0(pi0832), .Y(new_n15227_));
  AOI21X1  g12791(.A0(new_n15227_), .A1(new_n15226_), .B0(new_n15198_), .Y(po0320));
  INVX1    g12792(.A(pi0703), .Y(new_n15229_));
  OAI22X1  g12793(.A0(new_n14501_), .A1(new_n15229_), .B0(new_n5362_), .B1(pi0752), .Y(new_n15230_));
  OAI21X1  g12794(.A0(new_n2720_), .A1(pi0164), .B0(pi0832), .Y(new_n15231_));
  AOI21X1  g12795(.A0(new_n15230_), .A1(new_n2720_), .B0(new_n15231_), .Y(new_n15232_));
  OAI21X1  g12796(.A0(new_n14929_), .A1(new_n6826_), .B0(new_n2979_), .Y(new_n15233_));
  AOI21X1  g12797(.A0(new_n14557_), .A1(new_n6826_), .B0(new_n15233_), .Y(new_n15234_));
  INVX1    g12798(.A(pi0752), .Y(new_n15235_));
  OAI21X1  g12799(.A0(new_n14568_), .A1(pi0164), .B0(new_n14569_), .Y(new_n15236_));
  NAND2X1  g12800(.A(new_n15236_), .B(new_n15235_), .Y(new_n15237_));
  OAI21X1  g12801(.A0(new_n14588_), .A1(new_n6826_), .B0(new_n2979_), .Y(new_n15238_));
  AOI21X1  g12802(.A0(new_n14577_), .A1(new_n6826_), .B0(new_n15238_), .Y(new_n15239_));
  OAI21X1  g12803(.A0(new_n12077_), .A1(pi0164), .B0(new_n14591_), .Y(new_n15240_));
  NAND2X1  g12804(.A(new_n15240_), .B(pi0752), .Y(new_n15241_));
  OAI22X1  g12805(.A0(new_n15241_), .A1(new_n15239_), .B0(new_n15237_), .B1(new_n15234_), .Y(new_n15242_));
  OAI21X1  g12806(.A0(new_n14519_), .A1(new_n6826_), .B0(new_n15235_), .Y(new_n15243_));
  OR2X1    g12807(.A(new_n15243_), .B(new_n14520_), .Y(new_n15244_));
  NAND3X1  g12808(.A(new_n14536_), .B(new_n14523_), .C(new_n15235_), .Y(new_n15245_));
  OAI21X1  g12809(.A0(new_n12832_), .A1(new_n15235_), .B0(new_n15229_), .Y(new_n15246_));
  AOI21X1  g12810(.A0(new_n15245_), .A1(pi0164), .B0(new_n15246_), .Y(new_n15247_));
  AOI22X1  g12811(.A0(new_n15247_), .A1(new_n15244_), .B0(new_n15242_), .B1(pi0703), .Y(new_n15248_));
  OR2X1    g12812(.A(new_n15248_), .B(new_n9483_), .Y(new_n15249_));
  AOI21X1  g12813(.A0(new_n9483_), .A1(new_n6826_), .B0(pi0832), .Y(new_n15250_));
  AOI21X1  g12814(.A0(new_n15250_), .A1(new_n15249_), .B0(new_n15232_), .Y(po0321));
  OAI22X1  g12815(.A0(new_n14501_), .A1(new_n13538_), .B0(new_n5362_), .B1(pi0774), .Y(new_n15252_));
  OAI21X1  g12816(.A0(new_n2720_), .A1(pi0165), .B0(pi0832), .Y(new_n15253_));
  AOI21X1  g12817(.A0(new_n15252_), .A1(new_n2720_), .B0(new_n15253_), .Y(new_n15254_));
  OAI21X1  g12818(.A0(new_n14929_), .A1(new_n9867_), .B0(new_n2979_), .Y(new_n15255_));
  AOI21X1  g12819(.A0(new_n14557_), .A1(new_n9867_), .B0(new_n15255_), .Y(new_n15256_));
  OAI21X1  g12820(.A0(new_n14568_), .A1(pi0165), .B0(new_n14569_), .Y(new_n15257_));
  NAND2X1  g12821(.A(new_n15257_), .B(new_n13546_), .Y(new_n15258_));
  OAI21X1  g12822(.A0(new_n14588_), .A1(new_n9867_), .B0(new_n2979_), .Y(new_n15259_));
  AOI21X1  g12823(.A0(new_n14577_), .A1(new_n9867_), .B0(new_n15259_), .Y(new_n15260_));
  OAI21X1  g12824(.A0(new_n12077_), .A1(pi0165), .B0(new_n14591_), .Y(new_n15261_));
  NAND2X1  g12825(.A(new_n15261_), .B(pi0774), .Y(new_n15262_));
  OAI22X1  g12826(.A0(new_n15262_), .A1(new_n15260_), .B0(new_n15258_), .B1(new_n15256_), .Y(new_n15263_));
  OAI21X1  g12827(.A0(new_n14519_), .A1(new_n9867_), .B0(new_n13546_), .Y(new_n15264_));
  OR2X1    g12828(.A(new_n15264_), .B(new_n14520_), .Y(new_n15265_));
  NAND3X1  g12829(.A(new_n14536_), .B(new_n14523_), .C(new_n13546_), .Y(new_n15266_));
  OAI21X1  g12830(.A0(new_n12832_), .A1(new_n13546_), .B0(new_n13538_), .Y(new_n15267_));
  AOI21X1  g12831(.A0(new_n15266_), .A1(pi0165), .B0(new_n15267_), .Y(new_n15268_));
  AOI22X1  g12832(.A0(new_n15268_), .A1(new_n15265_), .B0(new_n15263_), .B1(pi0687), .Y(new_n15269_));
  OR2X1    g12833(.A(new_n15269_), .B(new_n9483_), .Y(new_n15270_));
  AOI21X1  g12834(.A0(new_n9483_), .A1(new_n9867_), .B0(pi0832), .Y(new_n15271_));
  AOI21X1  g12835(.A0(new_n15271_), .A1(new_n15270_), .B0(new_n15254_), .Y(po0322));
  OAI21X1  g12836(.A0(new_n14770_), .A1(new_n4459_), .B0(new_n14578_), .Y(new_n15273_));
  AOI22X1  g12837(.A0(new_n15273_), .A1(new_n14813_), .B0(new_n11932_), .B1(pi0947), .Y(new_n15274_));
  MX2X1    g12838(.A(pi0947), .B(pi0166), .S0(new_n11825_), .Y(new_n15275_));
  OAI21X1  g12839(.A0(new_n15275_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n15276_));
  AOI21X1  g12840(.A0(new_n14514_), .A1(pi0166), .B0(new_n14817_), .Y(new_n15277_));
  OAI21X1  g12841(.A0(new_n15276_), .A1(new_n15274_), .B0(new_n15277_), .Y(new_n15278_));
  OR2X1    g12842(.A(new_n11878_), .B(pi0166), .Y(new_n15279_));
  AOI21X1  g12843(.A0(new_n15279_), .A1(new_n14550_), .B0(pi0299), .Y(new_n15280_));
  OR2X1    g12844(.A(new_n11933_), .B(pi0166), .Y(new_n15281_));
  AOI22X1  g12845(.A0(new_n15281_), .A1(new_n14776_), .B0(new_n15275_), .B1(new_n2951_), .Y(new_n15282_));
  OAI21X1  g12846(.A0(new_n15282_), .A1(pi0223), .B0(new_n15280_), .Y(new_n15283_));
  AND2X1   g12847(.A(new_n15283_), .B(pi0772), .Y(new_n15284_));
  AOI21X1  g12848(.A0(new_n11957_), .A1(new_n11937_), .B0(pi0772), .Y(new_n15285_));
  AND2X1   g12849(.A(new_n15285_), .B(pi0166), .Y(new_n15286_));
  OR2X1    g12850(.A(new_n15286_), .B(new_n2939_), .Y(new_n15287_));
  AOI21X1  g12851(.A0(new_n15284_), .A1(new_n15278_), .B0(new_n15287_), .Y(new_n15288_));
  AOI21X1  g12852(.A0(pi0947), .A1(pi0772), .B0(pi0039), .Y(new_n15289_));
  OAI22X1  g12853(.A0(new_n15289_), .A1(new_n14803_), .B0(new_n11821_), .B1(new_n4459_), .Y(new_n15290_));
  NAND2X1  g12854(.A(new_n15290_), .B(new_n2979_), .Y(new_n15291_));
  INVX1    g12855(.A(pi0727), .Y(new_n15292_));
  AND2X1   g12856(.A(pi0947), .B(pi0772), .Y(new_n15293_));
  INVX1    g12857(.A(new_n15293_), .Y(new_n15294_));
  AOI21X1  g12858(.A0(new_n15294_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n15295_));
  OAI21X1  g12859(.A0(new_n12446_), .A1(pi0166), .B0(new_n15295_), .Y(new_n15296_));
  AND2X1   g12860(.A(new_n15296_), .B(new_n15292_), .Y(new_n15297_));
  OAI21X1  g12861(.A0(new_n15291_), .A1(new_n15288_), .B0(new_n15297_), .Y(new_n15298_));
  MX2X1    g12862(.A(new_n5055_), .B(new_n4459_), .S0(new_n11825_), .Y(new_n15299_));
  AND2X1   g12863(.A(new_n15299_), .B(new_n10044_), .Y(new_n15300_));
  OR2X1    g12864(.A(new_n15300_), .B(pi0215), .Y(new_n15301_));
  NOR2X1   g12865(.A(new_n15273_), .B(new_n14720_), .Y(new_n15302_));
  NOR2X1   g12866(.A(new_n15302_), .B(new_n15301_), .Y(new_n15303_));
  OAI21X1  g12867(.A0(new_n11951_), .A1(pi0166), .B0(new_n14540_), .Y(new_n15304_));
  NAND2X1  g12868(.A(new_n15304_), .B(pi0299), .Y(new_n15305_));
  INVX1    g12869(.A(pi0772), .Y(new_n15306_));
  AOI21X1  g12870(.A0(new_n15299_), .A1(new_n2951_), .B0(pi0223), .Y(new_n15307_));
  MX2X1    g12871(.A(pi0166), .B(new_n14453_), .S0(new_n11933_), .Y(new_n15308_));
  OAI21X1  g12872(.A0(new_n15308_), .A1(new_n14780_), .B0(new_n15307_), .Y(new_n15309_));
  AND2X1   g12873(.A(new_n11878_), .B(new_n14547_), .Y(new_n15310_));
  OAI21X1  g12874(.A0(new_n15310_), .A1(pi0166), .B0(new_n14551_), .Y(new_n15311_));
  AND2X1   g12875(.A(new_n15311_), .B(new_n15280_), .Y(new_n15312_));
  AOI21X1  g12876(.A0(new_n15312_), .A1(new_n15309_), .B0(new_n15306_), .Y(new_n15313_));
  OAI21X1  g12877(.A0(new_n15305_), .A1(new_n15303_), .B0(new_n15313_), .Y(new_n15314_));
  OR4X1    g12878(.A(new_n11824_), .B(new_n2952_), .C(new_n2725_), .D(new_n5362_), .Y(new_n15315_));
  AND2X1   g12879(.A(new_n15315_), .B(new_n15307_), .Y(new_n15316_));
  OAI21X1  g12880(.A0(new_n15308_), .A1(new_n2951_), .B0(new_n15316_), .Y(new_n15317_));
  AND3X1   g12881(.A(new_n15317_), .B(new_n15311_), .C(new_n2933_), .Y(new_n15318_));
  AOI21X1  g12882(.A0(new_n14501_), .A1(new_n11947_), .B0(new_n15301_), .Y(new_n15319_));
  OAI21X1  g12883(.A0(new_n15304_), .A1(new_n14798_), .B0(pi0299), .Y(new_n15320_));
  AOI21X1  g12884(.A0(new_n15319_), .A1(new_n15273_), .B0(new_n15320_), .Y(new_n15321_));
  OR3X1    g12885(.A(new_n15321_), .B(new_n15318_), .C(pi0772), .Y(new_n15322_));
  AND3X1   g12886(.A(new_n15322_), .B(new_n15314_), .C(pi0039), .Y(new_n15323_));
  OAI21X1  g12887(.A0(new_n15290_), .A1(new_n14586_), .B0(new_n2979_), .Y(new_n15324_));
  NAND2X1  g12888(.A(new_n15289_), .B(new_n14809_), .Y(new_n15325_));
  AOI21X1  g12889(.A0(new_n12771_), .A1(new_n4459_), .B0(new_n2979_), .Y(new_n15326_));
  AOI21X1  g12890(.A0(new_n15326_), .A1(new_n15325_), .B0(new_n15292_), .Y(new_n15327_));
  OAI21X1  g12891(.A0(new_n15324_), .A1(new_n15323_), .B0(new_n15327_), .Y(new_n15328_));
  AOI21X1  g12892(.A0(new_n15328_), .A1(new_n15298_), .B0(new_n9483_), .Y(new_n15329_));
  OAI21X1  g12893(.A0(new_n7625_), .A1(pi0166), .B0(new_n12767_), .Y(new_n15330_));
  OAI21X1  g12894(.A0(new_n5362_), .A1(new_n15306_), .B0(new_n2720_), .Y(new_n15331_));
  AOI21X1  g12895(.A0(new_n14453_), .A1(pi0727), .B0(new_n15331_), .Y(new_n15332_));
  OAI21X1  g12896(.A0(new_n2720_), .A1(pi0166), .B0(pi0832), .Y(new_n15333_));
  OAI22X1  g12897(.A0(new_n15333_), .A1(new_n15332_), .B0(new_n15330_), .B1(new_n15329_), .Y(po0323));
  INVX1    g12898(.A(pi0705), .Y(new_n15335_));
  OAI22X1  g12899(.A0(new_n14501_), .A1(new_n15335_), .B0(new_n5362_), .B1(pi0768), .Y(new_n15336_));
  OAI21X1  g12900(.A0(new_n2720_), .A1(pi0167), .B0(pi0832), .Y(new_n15337_));
  AOI21X1  g12901(.A0(new_n15336_), .A1(new_n2720_), .B0(new_n15337_), .Y(new_n15338_));
  AOI21X1  g12902(.A0(new_n14587_), .A1(pi0167), .B0(pi0038), .Y(new_n15339_));
  OAI21X1  g12903(.A0(new_n14576_), .A1(pi0167), .B0(new_n15339_), .Y(new_n15340_));
  OAI21X1  g12904(.A0(new_n12077_), .A1(pi0167), .B0(new_n14591_), .Y(new_n15341_));
  AND3X1   g12905(.A(new_n15341_), .B(new_n15340_), .C(pi0768), .Y(new_n15342_));
  OAI21X1  g12906(.A0(new_n14929_), .A1(new_n7437_), .B0(new_n2979_), .Y(new_n15343_));
  AOI21X1  g12907(.A0(new_n14557_), .A1(new_n7437_), .B0(new_n15343_), .Y(new_n15344_));
  INVX1    g12908(.A(pi0768), .Y(new_n15345_));
  OAI21X1  g12909(.A0(new_n14568_), .A1(pi0167), .B0(new_n14569_), .Y(new_n15346_));
  NAND2X1  g12910(.A(new_n15346_), .B(new_n15345_), .Y(new_n15347_));
  OAI21X1  g12911(.A0(new_n15347_), .A1(new_n15344_), .B0(pi0705), .Y(new_n15348_));
  OAI21X1  g12912(.A0(new_n14517_), .A1(new_n14505_), .B0(new_n7437_), .Y(new_n15349_));
  AOI21X1  g12913(.A0(new_n14535_), .A1(pi0167), .B0(pi0038), .Y(new_n15350_));
  AND2X1   g12914(.A(new_n15350_), .B(new_n15349_), .Y(new_n15351_));
  AOI21X1  g12915(.A0(new_n12831_), .A1(new_n7437_), .B0(new_n14523_), .Y(new_n15352_));
  OR3X1    g12916(.A(new_n15352_), .B(new_n15351_), .C(pi0768), .Y(new_n15353_));
  OR3X1    g12917(.A(new_n12447_), .B(new_n15345_), .C(pi0167), .Y(new_n15354_));
  AND2X1   g12918(.A(new_n15354_), .B(new_n15335_), .Y(new_n15355_));
  AOI21X1  g12919(.A0(new_n15355_), .A1(new_n15353_), .B0(new_n9483_), .Y(new_n15356_));
  OAI21X1  g12920(.A0(new_n15348_), .A1(new_n15342_), .B0(new_n15356_), .Y(new_n15357_));
  AOI21X1  g12921(.A0(new_n9483_), .A1(new_n7437_), .B0(pi0832), .Y(new_n15358_));
  AOI21X1  g12922(.A0(new_n15358_), .A1(new_n15357_), .B0(new_n15338_), .Y(po0324));
  AOI21X1  g12923(.A0(pi0947), .A1(pi0763), .B0(new_n2725_), .Y(new_n15360_));
  INVX1    g12924(.A(pi0699), .Y(new_n15361_));
  OR3X1    g12925(.A(pi0947), .B(new_n5277_), .C(new_n15361_), .Y(new_n15362_));
  OAI21X1  g12926(.A0(new_n2720_), .A1(new_n4308_), .B0(pi0832), .Y(new_n15363_));
  AOI21X1  g12927(.A0(new_n15362_), .A1(new_n15360_), .B0(new_n15363_), .Y(new_n15364_));
  INVX1    g12928(.A(pi0763), .Y(new_n15365_));
  AND3X1   g12929(.A(new_n11821_), .B(new_n15365_), .C(new_n2939_), .Y(new_n15366_));
  OAI22X1  g12930(.A0(new_n15366_), .A1(new_n14524_), .B0(new_n11821_), .B1(pi0168), .Y(new_n15367_));
  NOR2X1   g12931(.A(new_n11951_), .B(new_n4308_), .Y(new_n15368_));
  NOR3X1   g12932(.A(new_n15368_), .B(new_n11955_), .C(new_n2934_), .Y(new_n15369_));
  NOR2X1   g12933(.A(new_n10044_), .B(new_n4308_), .Y(new_n15370_));
  AOI22X1  g12934(.A0(new_n15370_), .A1(new_n14849_), .B0(new_n11945_), .B1(new_n10045_), .Y(new_n15371_));
  AND2X1   g12935(.A(new_n11825_), .B(new_n4308_), .Y(new_n15372_));
  NOR3X1   g12936(.A(new_n15372_), .B(new_n14529_), .C(new_n10045_), .Y(new_n15373_));
  AOI21X1  g12937(.A0(new_n15373_), .A1(new_n14852_), .B0(pi0215), .Y(new_n15374_));
  AOI21X1  g12938(.A0(new_n15374_), .A1(new_n15371_), .B0(new_n15369_), .Y(new_n15375_));
  OR2X1    g12939(.A(new_n15375_), .B(new_n2933_), .Y(new_n15376_));
  OAI21X1  g12940(.A0(new_n14729_), .A1(new_n4308_), .B0(new_n14553_), .Y(new_n15377_));
  AOI21X1  g12941(.A0(new_n15377_), .A1(new_n15376_), .B0(new_n15365_), .Y(new_n15378_));
  INVX1    g12942(.A(new_n15371_), .Y(new_n15379_));
  OAI22X1  g12943(.A0(new_n15372_), .A1(new_n14723_), .B0(new_n14542_), .B1(new_n10044_), .Y(new_n15380_));
  OAI21X1  g12944(.A0(new_n15380_), .A1(new_n15379_), .B0(new_n2934_), .Y(new_n15381_));
  OR3X1    g12945(.A(new_n15369_), .B(new_n11951_), .C(new_n2934_), .Y(new_n15382_));
  AND2X1   g12946(.A(new_n15382_), .B(new_n14732_), .Y(new_n15383_));
  AOI21X1  g12947(.A0(new_n15383_), .A1(new_n15381_), .B0(new_n2933_), .Y(new_n15384_));
  NOR2X1   g12948(.A(new_n14508_), .B(pi0168), .Y(new_n15385_));
  OAI21X1  g12949(.A0(new_n15385_), .A1(new_n14737_), .B0(new_n15365_), .Y(new_n15386_));
  OAI21X1  g12950(.A0(new_n15386_), .A1(new_n15384_), .B0(pi0039), .Y(new_n15387_));
  OAI22X1  g12951(.A0(new_n15387_), .A1(new_n15378_), .B0(new_n15367_), .B1(new_n14586_), .Y(new_n15388_));
  OAI21X1  g12952(.A0(new_n5362_), .A1(pi0763), .B0(new_n2939_), .Y(new_n15389_));
  OAI21X1  g12953(.A0(new_n15389_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15390_));
  AOI21X1  g12954(.A0(new_n12771_), .A1(new_n4308_), .B0(new_n15390_), .Y(new_n15391_));
  AOI21X1  g12955(.A0(new_n15388_), .A1(new_n2979_), .B0(new_n15391_), .Y(new_n15392_));
  NOR3X1   g12956(.A(new_n15385_), .B(new_n14525_), .C(pi0299), .Y(new_n15393_));
  NOR4X1   g12957(.A(new_n15373_), .B(new_n15379_), .C(new_n14511_), .D(pi0215), .Y(new_n15394_));
  OAI21X1  g12958(.A0(new_n15368_), .A1(new_n14876_), .B0(pi0299), .Y(new_n15395_));
  OAI21X1  g12959(.A0(new_n15395_), .A1(new_n15394_), .B0(pi0763), .Y(new_n15396_));
  NOR2X1   g12960(.A(new_n15396_), .B(new_n15393_), .Y(new_n15397_));
  OR2X1    g12961(.A(pi0763), .B(pi0168), .Y(new_n15398_));
  OAI21X1  g12962(.A0(new_n15398_), .A1(new_n12444_), .B0(pi0039), .Y(new_n15399_));
  AND2X1   g12963(.A(new_n15367_), .B(new_n2979_), .Y(new_n15400_));
  OAI21X1  g12964(.A0(new_n15399_), .A1(new_n15397_), .B0(new_n15400_), .Y(new_n15401_));
  AOI21X1  g12965(.A0(new_n15360_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n15402_));
  OAI21X1  g12966(.A0(new_n12446_), .A1(new_n4308_), .B0(new_n15402_), .Y(new_n15403_));
  AND2X1   g12967(.A(new_n15403_), .B(new_n15361_), .Y(new_n15404_));
  AOI21X1  g12968(.A0(new_n15404_), .A1(new_n15401_), .B0(new_n14616_), .Y(new_n15405_));
  OAI21X1  g12969(.A0(new_n15392_), .A1(new_n15361_), .B0(new_n15405_), .Y(new_n15406_));
  AOI21X1  g12970(.A0(new_n14616_), .A1(new_n4308_), .B0(pi0057), .Y(new_n15407_));
  OAI21X1  g12971(.A0(new_n4308_), .A1(new_n2436_), .B0(new_n12767_), .Y(new_n15408_));
  AOI21X1  g12972(.A0(new_n15407_), .A1(new_n15406_), .B0(new_n15408_), .Y(new_n15409_));
  OR2X1    g12973(.A(new_n15409_), .B(new_n15364_), .Y(po0325));
  AOI21X1  g12974(.A0(pi0947), .A1(pi0746), .B0(new_n2725_), .Y(new_n15411_));
  INVX1    g12975(.A(pi0729), .Y(new_n15412_));
  OR3X1    g12976(.A(pi0947), .B(new_n5277_), .C(new_n15412_), .Y(new_n15413_));
  OAI21X1  g12977(.A0(new_n2720_), .A1(new_n4162_), .B0(pi0832), .Y(new_n15414_));
  AOI21X1  g12978(.A0(new_n15413_), .A1(new_n15411_), .B0(new_n15414_), .Y(new_n15415_));
  INVX1    g12979(.A(pi0746), .Y(new_n15416_));
  AND3X1   g12980(.A(new_n11821_), .B(new_n15416_), .C(new_n2939_), .Y(new_n15417_));
  OAI22X1  g12981(.A0(new_n15417_), .A1(new_n14524_), .B0(new_n11821_), .B1(pi0169), .Y(new_n15418_));
  NOR2X1   g12982(.A(new_n11951_), .B(new_n4162_), .Y(new_n15419_));
  NOR3X1   g12983(.A(new_n15419_), .B(new_n11955_), .C(new_n2934_), .Y(new_n15420_));
  NOR2X1   g12984(.A(new_n10044_), .B(new_n4162_), .Y(new_n15421_));
  AOI22X1  g12985(.A0(new_n15421_), .A1(new_n14849_), .B0(new_n11945_), .B1(new_n10045_), .Y(new_n15422_));
  AND2X1   g12986(.A(new_n11825_), .B(new_n4162_), .Y(new_n15423_));
  NOR3X1   g12987(.A(new_n15423_), .B(new_n14529_), .C(new_n10045_), .Y(new_n15424_));
  AOI21X1  g12988(.A0(new_n15424_), .A1(new_n14852_), .B0(pi0215), .Y(new_n15425_));
  AOI21X1  g12989(.A0(new_n15425_), .A1(new_n15422_), .B0(new_n15420_), .Y(new_n15426_));
  OR2X1    g12990(.A(new_n15426_), .B(new_n2933_), .Y(new_n15427_));
  OAI21X1  g12991(.A0(new_n14729_), .A1(new_n4162_), .B0(new_n14553_), .Y(new_n15428_));
  AOI21X1  g12992(.A0(new_n15428_), .A1(new_n15427_), .B0(new_n15416_), .Y(new_n15429_));
  INVX1    g12993(.A(new_n15422_), .Y(new_n15430_));
  OAI22X1  g12994(.A0(new_n15423_), .A1(new_n14723_), .B0(new_n14542_), .B1(new_n10044_), .Y(new_n15431_));
  OAI21X1  g12995(.A0(new_n15431_), .A1(new_n15430_), .B0(new_n2934_), .Y(new_n15432_));
  OR3X1    g12996(.A(new_n15420_), .B(new_n11951_), .C(new_n2934_), .Y(new_n15433_));
  AND2X1   g12997(.A(new_n15433_), .B(new_n14732_), .Y(new_n15434_));
  AOI21X1  g12998(.A0(new_n15434_), .A1(new_n15432_), .B0(new_n2933_), .Y(new_n15435_));
  NOR2X1   g12999(.A(new_n14508_), .B(pi0169), .Y(new_n15436_));
  OAI21X1  g13000(.A0(new_n15436_), .A1(new_n14737_), .B0(new_n15416_), .Y(new_n15437_));
  OAI21X1  g13001(.A0(new_n15437_), .A1(new_n15435_), .B0(pi0039), .Y(new_n15438_));
  OAI22X1  g13002(.A0(new_n15438_), .A1(new_n15429_), .B0(new_n15418_), .B1(new_n14586_), .Y(new_n15439_));
  OAI21X1  g13003(.A0(new_n5362_), .A1(pi0746), .B0(new_n2939_), .Y(new_n15440_));
  OAI21X1  g13004(.A0(new_n15440_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15441_));
  AOI21X1  g13005(.A0(new_n12771_), .A1(new_n4162_), .B0(new_n15441_), .Y(new_n15442_));
  AOI21X1  g13006(.A0(new_n15439_), .A1(new_n2979_), .B0(new_n15442_), .Y(new_n15443_));
  NOR3X1   g13007(.A(new_n15436_), .B(new_n14525_), .C(pi0299), .Y(new_n15444_));
  NOR4X1   g13008(.A(new_n15424_), .B(new_n15430_), .C(new_n14511_), .D(pi0215), .Y(new_n15445_));
  OAI21X1  g13009(.A0(new_n15419_), .A1(new_n14876_), .B0(pi0299), .Y(new_n15446_));
  OAI21X1  g13010(.A0(new_n15446_), .A1(new_n15445_), .B0(pi0746), .Y(new_n15447_));
  NOR2X1   g13011(.A(new_n15447_), .B(new_n15444_), .Y(new_n15448_));
  OR2X1    g13012(.A(pi0746), .B(pi0169), .Y(new_n15449_));
  OAI21X1  g13013(.A0(new_n15449_), .A1(new_n12444_), .B0(pi0039), .Y(new_n15450_));
  AND2X1   g13014(.A(new_n15418_), .B(new_n2979_), .Y(new_n15451_));
  OAI21X1  g13015(.A0(new_n15450_), .A1(new_n15448_), .B0(new_n15451_), .Y(new_n15452_));
  AOI21X1  g13016(.A0(new_n15411_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n15453_));
  OAI21X1  g13017(.A0(new_n12446_), .A1(new_n4162_), .B0(new_n15453_), .Y(new_n15454_));
  AND2X1   g13018(.A(new_n15454_), .B(new_n15412_), .Y(new_n15455_));
  AOI21X1  g13019(.A0(new_n15455_), .A1(new_n15452_), .B0(new_n14616_), .Y(new_n15456_));
  OAI21X1  g13020(.A0(new_n15443_), .A1(new_n15412_), .B0(new_n15456_), .Y(new_n15457_));
  AOI21X1  g13021(.A0(new_n14616_), .A1(new_n4162_), .B0(pi0057), .Y(new_n15458_));
  OAI21X1  g13022(.A0(new_n4162_), .A1(new_n2436_), .B0(new_n12767_), .Y(new_n15459_));
  AOI21X1  g13023(.A0(new_n15458_), .A1(new_n15457_), .B0(new_n15459_), .Y(new_n15460_));
  OR2X1    g13024(.A(new_n15460_), .B(new_n15415_), .Y(po0326));
  INVX1    g13025(.A(pi0748), .Y(new_n15462_));
  OAI21X1  g13026(.A0(new_n5362_), .A1(new_n15462_), .B0(new_n2720_), .Y(new_n15463_));
  AOI21X1  g13027(.A0(new_n14453_), .A1(pi0730), .B0(new_n15463_), .Y(new_n15464_));
  OAI21X1  g13028(.A0(new_n2720_), .A1(new_n3865_), .B0(pi0832), .Y(new_n15465_));
  INVX1    g13029(.A(pi0730), .Y(new_n15466_));
  NOR2X1   g13030(.A(new_n14542_), .B(new_n10044_), .Y(new_n15467_));
  NOR2X1   g13031(.A(new_n10044_), .B(new_n3865_), .Y(new_n15468_));
  AOI22X1  g13032(.A0(new_n15468_), .A1(new_n14849_), .B0(new_n11945_), .B1(new_n10045_), .Y(new_n15469_));
  INVX1    g13033(.A(new_n15469_), .Y(new_n15470_));
  AOI21X1  g13034(.A0(new_n11825_), .A1(new_n3865_), .B0(new_n14723_), .Y(new_n15471_));
  NOR3X1   g13035(.A(new_n15471_), .B(new_n15470_), .C(new_n15467_), .Y(new_n15472_));
  NOR2X1   g13036(.A(new_n11951_), .B(new_n3865_), .Y(new_n15473_));
  NOR3X1   g13037(.A(new_n15473_), .B(new_n11955_), .C(new_n2934_), .Y(new_n15474_));
  OR3X1    g13038(.A(new_n15474_), .B(new_n11951_), .C(new_n2934_), .Y(new_n15475_));
  AND2X1   g13039(.A(new_n15475_), .B(new_n14732_), .Y(new_n15476_));
  OAI21X1  g13040(.A0(new_n15472_), .A1(pi0215), .B0(new_n15476_), .Y(new_n15477_));
  AOI21X1  g13041(.A0(new_n14599_), .A1(new_n3865_), .B0(pi0299), .Y(new_n15478_));
  AOI22X1  g13042(.A0(new_n15478_), .A1(new_n14584_), .B0(new_n15477_), .B1(pi0299), .Y(new_n15479_));
  NOR2X1   g13043(.A(new_n11821_), .B(pi0170), .Y(new_n15480_));
  OAI22X1  g13044(.A0(new_n15480_), .A1(new_n14714_), .B0(new_n15479_), .B1(new_n2939_), .Y(new_n15481_));
  OAI21X1  g13045(.A0(new_n12077_), .A1(pi0170), .B0(new_n14591_), .Y(new_n15482_));
  NAND2X1  g13046(.A(new_n15482_), .B(new_n15462_), .Y(new_n15483_));
  AOI21X1  g13047(.A0(new_n15481_), .A1(new_n2979_), .B0(new_n15483_), .Y(new_n15484_));
  NOR3X1   g13048(.A(new_n15480_), .B(new_n14907_), .C(pi0039), .Y(new_n15485_));
  OR2X1    g13049(.A(new_n14729_), .B(new_n3865_), .Y(new_n15486_));
  AOI21X1  g13050(.A0(new_n11825_), .A1(new_n3865_), .B0(new_n14752_), .Y(new_n15487_));
  AOI21X1  g13051(.A0(new_n15487_), .A1(new_n14852_), .B0(pi0215), .Y(new_n15488_));
  AOI21X1  g13052(.A0(new_n15488_), .A1(new_n15469_), .B0(new_n15474_), .Y(new_n15489_));
  OAI21X1  g13053(.A0(new_n15489_), .A1(new_n2933_), .B0(pi0039), .Y(new_n15490_));
  AOI21X1  g13054(.A0(new_n15486_), .A1(new_n14553_), .B0(new_n15490_), .Y(new_n15491_));
  OAI21X1  g13055(.A0(new_n15491_), .A1(new_n15485_), .B0(new_n2979_), .Y(new_n15492_));
  OAI21X1  g13056(.A0(new_n12077_), .A1(pi0170), .B0(new_n14569_), .Y(new_n15493_));
  AND3X1   g13057(.A(new_n15493_), .B(new_n15492_), .C(pi0748), .Y(new_n15494_));
  OR3X1    g13058(.A(new_n15494_), .B(new_n15484_), .C(new_n15466_), .Y(new_n15495_));
  INVX1    g13059(.A(new_n15480_), .Y(new_n15496_));
  NOR4X1   g13060(.A(new_n15487_), .B(new_n15470_), .C(new_n14511_), .D(pi0215), .Y(new_n15497_));
  OAI21X1  g13061(.A0(new_n15473_), .A1(new_n14876_), .B0(pi0299), .Y(new_n15498_));
  OAI21X1  g13062(.A0(new_n14599_), .A1(new_n5362_), .B0(new_n15478_), .Y(new_n15499_));
  OAI21X1  g13063(.A0(new_n15498_), .A1(new_n15497_), .B0(new_n15499_), .Y(new_n15500_));
  AOI22X1  g13064(.A0(new_n15500_), .A1(pi0039), .B0(new_n15496_), .B1(new_n14524_), .Y(new_n15501_));
  OAI22X1  g13065(.A0(new_n14519_), .A1(new_n13265_), .B0(new_n12446_), .B1(pi0170), .Y(new_n15502_));
  AND2X1   g13066(.A(new_n15502_), .B(pi0748), .Y(new_n15503_));
  OAI21X1  g13067(.A0(new_n15501_), .A1(pi0038), .B0(new_n15503_), .Y(new_n15504_));
  NOR2X1   g13068(.A(pi0748), .B(pi0170), .Y(new_n15505_));
  AOI21X1  g13069(.A0(new_n15505_), .A1(new_n12832_), .B0(pi0730), .Y(new_n15506_));
  AOI21X1  g13070(.A0(new_n15506_), .A1(new_n15504_), .B0(new_n14616_), .Y(new_n15507_));
  OAI21X1  g13071(.A0(new_n14615_), .A1(pi0170), .B0(new_n2436_), .Y(new_n15508_));
  AOI21X1  g13072(.A0(new_n15507_), .A1(new_n15495_), .B0(new_n15508_), .Y(new_n15509_));
  OAI21X1  g13073(.A0(new_n3865_), .A1(new_n2436_), .B0(new_n12767_), .Y(new_n15510_));
  OAI22X1  g13074(.A0(new_n15510_), .A1(new_n15509_), .B0(new_n15465_), .B1(new_n15464_), .Y(po0327));
  AOI21X1  g13075(.A0(pi0947), .A1(pi0764), .B0(new_n2725_), .Y(new_n15512_));
  INVX1    g13076(.A(pi0691), .Y(new_n15513_));
  OR3X1    g13077(.A(pi0947), .B(new_n5277_), .C(new_n15513_), .Y(new_n15514_));
  OAI21X1  g13078(.A0(new_n2720_), .A1(new_n3715_), .B0(pi0832), .Y(new_n15515_));
  AOI21X1  g13079(.A0(new_n15514_), .A1(new_n15512_), .B0(new_n15515_), .Y(new_n15516_));
  INVX1    g13080(.A(pi0764), .Y(new_n15517_));
  AND3X1   g13081(.A(new_n11821_), .B(new_n15517_), .C(new_n2939_), .Y(new_n15518_));
  OAI22X1  g13082(.A0(new_n15518_), .A1(new_n14524_), .B0(new_n11821_), .B1(pi0171), .Y(new_n15519_));
  NOR2X1   g13083(.A(new_n11951_), .B(new_n3715_), .Y(new_n15520_));
  NOR3X1   g13084(.A(new_n15520_), .B(new_n11955_), .C(new_n2934_), .Y(new_n15521_));
  NOR2X1   g13085(.A(new_n10044_), .B(new_n3715_), .Y(new_n15522_));
  AOI22X1  g13086(.A0(new_n15522_), .A1(new_n14849_), .B0(new_n11945_), .B1(new_n10045_), .Y(new_n15523_));
  AND2X1   g13087(.A(new_n11825_), .B(new_n3715_), .Y(new_n15524_));
  NOR3X1   g13088(.A(new_n15524_), .B(new_n14529_), .C(new_n10045_), .Y(new_n15525_));
  AOI21X1  g13089(.A0(new_n15525_), .A1(new_n14852_), .B0(pi0215), .Y(new_n15526_));
  AOI21X1  g13090(.A0(new_n15526_), .A1(new_n15523_), .B0(new_n15521_), .Y(new_n15527_));
  OR2X1    g13091(.A(new_n15527_), .B(new_n2933_), .Y(new_n15528_));
  OAI21X1  g13092(.A0(new_n14729_), .A1(new_n3715_), .B0(new_n14553_), .Y(new_n15529_));
  AOI21X1  g13093(.A0(new_n15529_), .A1(new_n15528_), .B0(new_n15517_), .Y(new_n15530_));
  INVX1    g13094(.A(new_n15523_), .Y(new_n15531_));
  OAI22X1  g13095(.A0(new_n15524_), .A1(new_n14723_), .B0(new_n14542_), .B1(new_n10044_), .Y(new_n15532_));
  OAI21X1  g13096(.A0(new_n15532_), .A1(new_n15531_), .B0(new_n2934_), .Y(new_n15533_));
  OR3X1    g13097(.A(new_n15521_), .B(new_n11951_), .C(new_n2934_), .Y(new_n15534_));
  AND2X1   g13098(.A(new_n15534_), .B(new_n14732_), .Y(new_n15535_));
  AOI21X1  g13099(.A0(new_n15535_), .A1(new_n15533_), .B0(new_n2933_), .Y(new_n15536_));
  NOR2X1   g13100(.A(new_n14508_), .B(pi0171), .Y(new_n15537_));
  OAI21X1  g13101(.A0(new_n15537_), .A1(new_n14737_), .B0(new_n15517_), .Y(new_n15538_));
  OAI21X1  g13102(.A0(new_n15538_), .A1(new_n15536_), .B0(pi0039), .Y(new_n15539_));
  OAI22X1  g13103(.A0(new_n15539_), .A1(new_n15530_), .B0(new_n15519_), .B1(new_n14586_), .Y(new_n15540_));
  OAI21X1  g13104(.A0(new_n5362_), .A1(pi0764), .B0(new_n2939_), .Y(new_n15541_));
  OAI21X1  g13105(.A0(new_n15541_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15542_));
  AOI21X1  g13106(.A0(new_n12771_), .A1(new_n3715_), .B0(new_n15542_), .Y(new_n15543_));
  AOI21X1  g13107(.A0(new_n15540_), .A1(new_n2979_), .B0(new_n15543_), .Y(new_n15544_));
  NOR3X1   g13108(.A(new_n15537_), .B(new_n14525_), .C(pi0299), .Y(new_n15545_));
  NOR4X1   g13109(.A(new_n15525_), .B(new_n15531_), .C(new_n14511_), .D(pi0215), .Y(new_n15546_));
  OAI21X1  g13110(.A0(new_n15520_), .A1(new_n14876_), .B0(pi0299), .Y(new_n15547_));
  OAI21X1  g13111(.A0(new_n15547_), .A1(new_n15546_), .B0(pi0764), .Y(new_n15548_));
  NOR2X1   g13112(.A(new_n15548_), .B(new_n15545_), .Y(new_n15549_));
  OR2X1    g13113(.A(pi0764), .B(pi0171), .Y(new_n15550_));
  OAI21X1  g13114(.A0(new_n15550_), .A1(new_n12444_), .B0(pi0039), .Y(new_n15551_));
  AND2X1   g13115(.A(new_n15519_), .B(new_n2979_), .Y(new_n15552_));
  OAI21X1  g13116(.A0(new_n15551_), .A1(new_n15549_), .B0(new_n15552_), .Y(new_n15553_));
  AOI21X1  g13117(.A0(new_n15512_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n15554_));
  OAI21X1  g13118(.A0(new_n12446_), .A1(new_n3715_), .B0(new_n15554_), .Y(new_n15555_));
  AND2X1   g13119(.A(new_n15555_), .B(new_n15513_), .Y(new_n15556_));
  AOI21X1  g13120(.A0(new_n15556_), .A1(new_n15553_), .B0(new_n14616_), .Y(new_n15557_));
  OAI21X1  g13121(.A0(new_n15544_), .A1(new_n15513_), .B0(new_n15557_), .Y(new_n15558_));
  AOI21X1  g13122(.A0(new_n14616_), .A1(new_n3715_), .B0(pi0057), .Y(new_n15559_));
  OAI21X1  g13123(.A0(new_n3715_), .A1(new_n2436_), .B0(new_n12767_), .Y(new_n15560_));
  AOI21X1  g13124(.A0(new_n15559_), .A1(new_n15558_), .B0(new_n15560_), .Y(new_n15561_));
  OR2X1    g13125(.A(new_n15561_), .B(new_n15516_), .Y(po0328));
  AND2X1   g13126(.A(pi0947), .B(pi0739), .Y(new_n15563_));
  NOR3X1   g13127(.A(new_n15563_), .B(new_n5032_), .C(new_n5024_), .Y(new_n15564_));
  INVX1    g13128(.A(pi0690), .Y(new_n15565_));
  OR3X1    g13129(.A(pi0947), .B(new_n5277_), .C(new_n15565_), .Y(new_n15566_));
  OAI21X1  g13130(.A0(new_n2720_), .A1(new_n7084_), .B0(pi0832), .Y(new_n15567_));
  AOI21X1  g13131(.A0(new_n15566_), .A1(new_n15564_), .B0(new_n15567_), .Y(new_n15568_));
  AOI21X1  g13132(.A0(new_n15563_), .A1(new_n11821_), .B0(pi0039), .Y(new_n15569_));
  OAI21X1  g13133(.A0(new_n11821_), .A1(pi0172), .B0(new_n15569_), .Y(new_n15570_));
  INVX1    g13134(.A(pi0739), .Y(new_n15571_));
  NOR2X1   g13135(.A(new_n11951_), .B(new_n7084_), .Y(new_n15572_));
  NOR3X1   g13136(.A(new_n15572_), .B(new_n11955_), .C(new_n2934_), .Y(new_n15573_));
  NOR3X1   g13137(.A(new_n14720_), .B(new_n10044_), .C(new_n7084_), .Y(new_n15574_));
  AOI21X1  g13138(.A0(new_n11945_), .A1(new_n10045_), .B0(new_n15574_), .Y(new_n15575_));
  AND2X1   g13139(.A(new_n11825_), .B(new_n7084_), .Y(new_n15576_));
  NOR3X1   g13140(.A(new_n15576_), .B(new_n14529_), .C(new_n10045_), .Y(new_n15577_));
  AOI21X1  g13141(.A0(new_n15577_), .A1(new_n14852_), .B0(pi0215), .Y(new_n15578_));
  AOI21X1  g13142(.A0(new_n15578_), .A1(new_n15575_), .B0(new_n15573_), .Y(new_n15579_));
  OR2X1    g13143(.A(new_n15579_), .B(new_n2933_), .Y(new_n15580_));
  OAI21X1  g13144(.A0(new_n14729_), .A1(new_n7084_), .B0(new_n14553_), .Y(new_n15581_));
  AOI21X1  g13145(.A0(new_n15581_), .A1(new_n15580_), .B0(new_n15571_), .Y(new_n15582_));
  INVX1    g13146(.A(new_n15575_), .Y(new_n15583_));
  OAI22X1  g13147(.A0(new_n15576_), .A1(new_n14723_), .B0(new_n14542_), .B1(new_n10044_), .Y(new_n15584_));
  OAI21X1  g13148(.A0(new_n15584_), .A1(new_n15583_), .B0(new_n2934_), .Y(new_n15585_));
  OR3X1    g13149(.A(new_n15573_), .B(new_n11951_), .C(new_n2934_), .Y(new_n15586_));
  AND2X1   g13150(.A(new_n15586_), .B(new_n14732_), .Y(new_n15587_));
  AOI21X1  g13151(.A0(new_n15587_), .A1(new_n15585_), .B0(new_n2933_), .Y(new_n15588_));
  NOR2X1   g13152(.A(new_n14508_), .B(pi0172), .Y(new_n15589_));
  OAI21X1  g13153(.A0(new_n15589_), .A1(new_n14737_), .B0(new_n15571_), .Y(new_n15590_));
  OAI21X1  g13154(.A0(new_n15590_), .A1(new_n15588_), .B0(pi0039), .Y(new_n15591_));
  OAI22X1  g13155(.A0(new_n15591_), .A1(new_n15582_), .B0(new_n15570_), .B1(new_n14586_), .Y(new_n15592_));
  OAI21X1  g13156(.A0(new_n5362_), .A1(pi0739), .B0(new_n2939_), .Y(new_n15593_));
  OAI21X1  g13157(.A0(new_n15593_), .A1(new_n14669_), .B0(pi0038), .Y(new_n15594_));
  AOI21X1  g13158(.A0(new_n12771_), .A1(new_n7084_), .B0(new_n15594_), .Y(new_n15595_));
  AOI21X1  g13159(.A0(new_n15592_), .A1(new_n2979_), .B0(new_n15595_), .Y(new_n15596_));
  NOR3X1   g13160(.A(new_n15589_), .B(new_n14525_), .C(pi0299), .Y(new_n15597_));
  NOR4X1   g13161(.A(new_n15577_), .B(new_n15583_), .C(new_n14511_), .D(pi0215), .Y(new_n15598_));
  OAI21X1  g13162(.A0(new_n15572_), .A1(new_n14876_), .B0(pi0299), .Y(new_n15599_));
  OAI21X1  g13163(.A0(new_n15599_), .A1(new_n15598_), .B0(pi0739), .Y(new_n15600_));
  NOR2X1   g13164(.A(new_n15600_), .B(new_n15597_), .Y(new_n15601_));
  OR2X1    g13165(.A(pi0739), .B(pi0172), .Y(new_n15602_));
  OAI21X1  g13166(.A0(new_n15602_), .A1(new_n12444_), .B0(pi0039), .Y(new_n15603_));
  AND2X1   g13167(.A(new_n15570_), .B(new_n2979_), .Y(new_n15604_));
  OAI21X1  g13168(.A0(new_n15603_), .A1(new_n15601_), .B0(new_n15604_), .Y(new_n15605_));
  AOI21X1  g13169(.A0(new_n15564_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n15606_));
  OAI21X1  g13170(.A0(new_n12446_), .A1(new_n7084_), .B0(new_n15606_), .Y(new_n15607_));
  AND2X1   g13171(.A(new_n15607_), .B(new_n15565_), .Y(new_n15608_));
  AOI21X1  g13172(.A0(new_n15608_), .A1(new_n15605_), .B0(new_n14616_), .Y(new_n15609_));
  OAI21X1  g13173(.A0(new_n15596_), .A1(new_n15565_), .B0(new_n15609_), .Y(new_n15610_));
  AOI21X1  g13174(.A0(new_n14616_), .A1(new_n7084_), .B0(pi0057), .Y(new_n15611_));
  OAI21X1  g13175(.A0(new_n7084_), .A1(new_n2436_), .B0(new_n12767_), .Y(new_n15612_));
  AOI21X1  g13176(.A0(new_n15611_), .A1(new_n15610_), .B0(new_n15612_), .Y(new_n15613_));
  OR2X1    g13177(.A(new_n15613_), .B(new_n15568_), .Y(po0329));
  AOI21X1  g13178(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0173), .Y(new_n15615_));
  INVX1    g13179(.A(new_n15615_), .Y(new_n15616_));
  OAI21X1  g13180(.A0(new_n11770_), .A1(pi0723), .B0(new_n15615_), .Y(new_n15617_));
  OAI21X1  g13181(.A0(new_n12826_), .A1(new_n9903_), .B0(new_n2979_), .Y(new_n15618_));
  AOI22X1  g13182(.A0(new_n15618_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n9903_), .Y(new_n15619_));
  AOI21X1  g13183(.A0(new_n12771_), .A1(new_n9903_), .B0(new_n12441_), .Y(new_n15620_));
  OR3X1    g13184(.A(new_n15620_), .B(new_n15619_), .C(pi0723), .Y(new_n15621_));
  NAND3X1  g13185(.A(new_n15621_), .B(new_n15617_), .C(new_n11769_), .Y(new_n15622_));
  AOI21X1  g13186(.A0(new_n15621_), .A1(new_n15617_), .B0(new_n12363_), .Y(new_n15623_));
  OAI21X1  g13187(.A0(new_n15616_), .A1(pi0625), .B0(pi1153), .Y(new_n15624_));
  NOR2X1   g13188(.A(new_n15624_), .B(new_n15623_), .Y(new_n15625_));
  AOI21X1  g13189(.A0(new_n15621_), .A1(new_n15617_), .B0(pi0625), .Y(new_n15626_));
  OAI21X1  g13190(.A0(new_n15616_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n15627_));
  NOR2X1   g13191(.A(new_n15627_), .B(new_n15626_), .Y(new_n15628_));
  OAI21X1  g13192(.A0(new_n15628_), .A1(new_n15625_), .B0(pi0778), .Y(new_n15629_));
  AND2X1   g13193(.A(new_n15629_), .B(new_n15622_), .Y(new_n15630_));
  MX2X1    g13194(.A(new_n15630_), .B(new_n15615_), .S0(new_n12490_), .Y(new_n15631_));
  INVX1    g13195(.A(new_n15631_), .Y(new_n15632_));
  MX2X1    g13196(.A(new_n15632_), .B(new_n15616_), .S0(new_n12513_), .Y(new_n15633_));
  INVX1    g13197(.A(new_n15633_), .Y(new_n15634_));
  MX2X1    g13198(.A(new_n15634_), .B(new_n15615_), .S0(new_n12531_), .Y(new_n15635_));
  INVX1    g13199(.A(new_n15635_), .Y(new_n15636_));
  MX2X1    g13200(.A(new_n15636_), .B(new_n15616_), .S0(new_n12563_), .Y(new_n15637_));
  AOI21X1  g13201(.A0(new_n15615_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n15638_));
  OAI21X1  g13202(.A0(new_n15637_), .A1(new_n12554_), .B0(new_n15638_), .Y(new_n15639_));
  AOI21X1  g13203(.A0(new_n15615_), .A1(pi0628), .B0(pi1156), .Y(new_n15640_));
  OAI21X1  g13204(.A0(new_n15637_), .A1(pi0628), .B0(new_n15640_), .Y(new_n15641_));
  AOI21X1  g13205(.A0(new_n15641_), .A1(new_n15639_), .B0(new_n11764_), .Y(new_n15642_));
  AOI21X1  g13206(.A0(new_n15637_), .A1(new_n11764_), .B0(new_n15642_), .Y(new_n15643_));
  MX2X1    g13207(.A(new_n15643_), .B(new_n15615_), .S0(pi0647), .Y(new_n15644_));
  MX2X1    g13208(.A(new_n15643_), .B(new_n15615_), .S0(new_n12577_), .Y(new_n15645_));
  MX2X1    g13209(.A(new_n15645_), .B(new_n15644_), .S0(new_n12578_), .Y(new_n15646_));
  MX2X1    g13210(.A(new_n15646_), .B(new_n15643_), .S0(new_n11763_), .Y(new_n15647_));
  AOI21X1  g13211(.A0(new_n15647_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n15648_));
  AOI21X1  g13212(.A0(new_n11959_), .A1(new_n9903_), .B0(new_n14715_), .Y(new_n15649_));
  NOR2X1   g13213(.A(pi0745), .B(pi0173), .Y(new_n15650_));
  INVX1    g13214(.A(new_n15650_), .Y(new_n15651_));
  OAI22X1  g13215(.A0(new_n15651_), .A1(new_n12776_), .B0(new_n12074_), .B1(new_n9903_), .Y(new_n15652_));
  OAI21X1  g13216(.A0(new_n15652_), .A1(new_n15649_), .B0(new_n2979_), .Y(new_n15653_));
  AOI21X1  g13217(.A0(new_n12771_), .A1(new_n9903_), .B0(new_n2979_), .Y(new_n15654_));
  OAI21X1  g13218(.A0(new_n14197_), .A1(pi0745), .B0(new_n15654_), .Y(new_n15655_));
  NAND2X1  g13219(.A(new_n15655_), .B(new_n15653_), .Y(new_n15656_));
  MX2X1    g13220(.A(new_n15656_), .B(pi0173), .S0(new_n11770_), .Y(new_n15657_));
  AND2X1   g13221(.A(new_n15657_), .B(new_n12474_), .Y(new_n15658_));
  AOI21X1  g13222(.A0(new_n15616_), .A1(new_n12473_), .B0(new_n15658_), .Y(new_n15659_));
  AOI22X1  g13223(.A0(new_n15658_), .A1(pi0609), .B0(new_n15616_), .B1(new_n12472_), .Y(new_n15660_));
  NOR2X1   g13224(.A(new_n15660_), .B(new_n12463_), .Y(new_n15661_));
  AOI22X1  g13225(.A0(new_n15658_), .A1(new_n12462_), .B0(new_n15616_), .B1(new_n12481_), .Y(new_n15662_));
  NOR2X1   g13226(.A(new_n15662_), .B(pi1155), .Y(new_n15663_));
  OAI21X1  g13227(.A0(new_n15663_), .A1(new_n15661_), .B0(pi0785), .Y(new_n15664_));
  OAI21X1  g13228(.A0(new_n15659_), .A1(pi0785), .B0(new_n15664_), .Y(new_n15665_));
  AOI21X1  g13229(.A0(new_n15615_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n15666_));
  OAI21X1  g13230(.A0(new_n15665_), .A1(new_n12486_), .B0(new_n15666_), .Y(new_n15667_));
  AOI21X1  g13231(.A0(new_n15615_), .A1(pi0618), .B0(pi1154), .Y(new_n15668_));
  OAI21X1  g13232(.A0(new_n15665_), .A1(pi0618), .B0(new_n15668_), .Y(new_n15669_));
  NAND2X1  g13233(.A(new_n15669_), .B(new_n15667_), .Y(new_n15670_));
  MX2X1    g13234(.A(new_n15670_), .B(new_n15665_), .S0(new_n11767_), .Y(new_n15671_));
  AND2X1   g13235(.A(new_n15671_), .B(new_n11766_), .Y(new_n15672_));
  AOI21X1  g13236(.A0(new_n15615_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n15673_));
  OAI21X1  g13237(.A0(new_n15671_), .A1(new_n12509_), .B0(new_n15673_), .Y(new_n15674_));
  AOI21X1  g13238(.A0(new_n15615_), .A1(pi0619), .B0(pi1159), .Y(new_n15675_));
  OAI21X1  g13239(.A0(new_n15671_), .A1(pi0619), .B0(new_n15675_), .Y(new_n15676_));
  AOI21X1  g13240(.A0(new_n15676_), .A1(new_n15674_), .B0(new_n11766_), .Y(new_n15677_));
  OR2X1    g13241(.A(new_n15677_), .B(new_n15672_), .Y(new_n15678_));
  AND2X1   g13242(.A(new_n15678_), .B(new_n11765_), .Y(new_n15679_));
  NOR3X1   g13243(.A(new_n15677_), .B(new_n15672_), .C(new_n12542_), .Y(new_n15680_));
  AOI21X1  g13244(.A0(new_n15615_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n15681_));
  INVX1    g13245(.A(new_n15681_), .Y(new_n15682_));
  NOR3X1   g13246(.A(new_n15677_), .B(new_n15672_), .C(pi0626), .Y(new_n15683_));
  AOI21X1  g13247(.A0(new_n15615_), .A1(pi0626), .B0(pi1158), .Y(new_n15684_));
  INVX1    g13248(.A(new_n15684_), .Y(new_n15685_));
  OAI22X1  g13249(.A0(new_n15685_), .A1(new_n15683_), .B0(new_n15682_), .B1(new_n15680_), .Y(new_n15686_));
  AOI21X1  g13250(.A0(new_n15686_), .A1(pi0788), .B0(new_n15679_), .Y(new_n15687_));
  MX2X1    g13251(.A(new_n15687_), .B(new_n15615_), .S0(new_n12580_), .Y(new_n15688_));
  MX2X1    g13252(.A(new_n15688_), .B(new_n15615_), .S0(new_n12604_), .Y(new_n15689_));
  OAI21X1  g13253(.A0(new_n15616_), .A1(pi0644), .B0(new_n12608_), .Y(new_n15690_));
  AOI21X1  g13254(.A0(new_n15689_), .A1(pi0644), .B0(new_n15690_), .Y(new_n15691_));
  OR3X1    g13255(.A(new_n15691_), .B(new_n15648_), .C(new_n11762_), .Y(new_n15692_));
  NOR2X1   g13256(.A(new_n15688_), .B(new_n14239_), .Y(new_n15693_));
  OAI22X1  g13257(.A0(new_n15645_), .A1(new_n14242_), .B0(new_n15644_), .B1(new_n14244_), .Y(new_n15694_));
  OAI21X1  g13258(.A0(new_n15694_), .A1(new_n15693_), .B0(pi0787), .Y(new_n15695_));
  MX2X1    g13259(.A(new_n15641_), .B(new_n15639_), .S0(new_n12561_), .Y(new_n15696_));
  OAI21X1  g13260(.A0(new_n15687_), .A1(new_n14250_), .B0(new_n15696_), .Y(new_n15697_));
  NAND3X1  g13261(.A(new_n15655_), .B(new_n15653_), .C(pi0723), .Y(new_n15698_));
  OAI21X1  g13262(.A0(new_n12213_), .A1(new_n9903_), .B0(pi0745), .Y(new_n15699_));
  AOI21X1  g13263(.A0(new_n12155_), .A1(new_n9903_), .B0(new_n15699_), .Y(new_n15700_));
  AOI21X1  g13264(.A0(new_n12788_), .A1(new_n9903_), .B0(pi0745), .Y(new_n15701_));
  OAI21X1  g13265(.A0(new_n12787_), .A1(new_n9903_), .B0(new_n15701_), .Y(new_n15702_));
  NAND2X1  g13266(.A(new_n15702_), .B(pi0039), .Y(new_n15703_));
  AND2X1   g13267(.A(new_n12332_), .B(pi0173), .Y(new_n15704_));
  OAI21X1  g13268(.A0(new_n12315_), .A1(pi0173), .B0(pi0745), .Y(new_n15705_));
  NOR4X1   g13269(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0173), .Y(new_n15706_));
  OAI21X1  g13270(.A0(new_n12800_), .A1(new_n9903_), .B0(new_n14715_), .Y(new_n15707_));
  OAI22X1  g13271(.A0(new_n15707_), .A1(new_n15706_), .B0(new_n15705_), .B1(new_n15704_), .Y(new_n15708_));
  AOI21X1  g13272(.A0(new_n15708_), .A1(new_n2939_), .B0(pi0038), .Y(new_n15709_));
  OAI21X1  g13273(.A0(new_n15703_), .A1(new_n15700_), .B0(new_n15709_), .Y(new_n15710_));
  OAI21X1  g13274(.A0(new_n12276_), .A1(pi0745), .B0(new_n13540_), .Y(new_n15711_));
  NAND2X1  g13275(.A(new_n15711_), .B(new_n9903_), .Y(new_n15712_));
  AOI21X1  g13276(.A0(new_n12056_), .A1(new_n14715_), .B0(new_n13443_), .Y(new_n15713_));
  NOR2X1   g13277(.A(new_n15713_), .B(new_n9903_), .Y(new_n15714_));
  AOI21X1  g13278(.A0(new_n15714_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n15715_));
  AOI21X1  g13279(.A0(new_n15715_), .A1(new_n15712_), .B0(pi0723), .Y(new_n15716_));
  AOI21X1  g13280(.A0(new_n15716_), .A1(new_n15710_), .B0(new_n11770_), .Y(new_n15717_));
  AOI22X1  g13281(.A0(new_n15717_), .A1(new_n15698_), .B0(new_n11770_), .B1(pi0173), .Y(new_n15718_));
  OAI21X1  g13282(.A0(new_n15657_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n15719_));
  AOI21X1  g13283(.A0(new_n15718_), .A1(new_n12363_), .B0(new_n15719_), .Y(new_n15720_));
  OR3X1    g13284(.A(new_n15720_), .B(new_n15625_), .C(pi0608), .Y(new_n15721_));
  OAI21X1  g13285(.A0(new_n15657_), .A1(pi0625), .B0(pi1153), .Y(new_n15722_));
  AOI21X1  g13286(.A0(new_n15718_), .A1(pi0625), .B0(new_n15722_), .Y(new_n15723_));
  OR3X1    g13287(.A(new_n15723_), .B(new_n15628_), .C(new_n12368_), .Y(new_n15724_));
  AOI21X1  g13288(.A0(new_n15724_), .A1(new_n15721_), .B0(new_n11769_), .Y(new_n15725_));
  AOI21X1  g13289(.A0(new_n15718_), .A1(new_n11769_), .B0(new_n15725_), .Y(new_n15726_));
  AOI21X1  g13290(.A0(new_n15630_), .A1(pi0609), .B0(pi1155), .Y(new_n15727_));
  OAI21X1  g13291(.A0(new_n15726_), .A1(pi0609), .B0(new_n15727_), .Y(new_n15728_));
  NOR2X1   g13292(.A(new_n15661_), .B(pi0660), .Y(new_n15729_));
  AOI21X1  g13293(.A0(new_n15630_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n15730_));
  OAI21X1  g13294(.A0(new_n15726_), .A1(new_n12462_), .B0(new_n15730_), .Y(new_n15731_));
  NOR2X1   g13295(.A(new_n15663_), .B(new_n12468_), .Y(new_n15732_));
  AOI22X1  g13296(.A0(new_n15732_), .A1(new_n15731_), .B0(new_n15729_), .B1(new_n15728_), .Y(new_n15733_));
  OR2X1    g13297(.A(new_n15726_), .B(pi0785), .Y(new_n15734_));
  OAI21X1  g13298(.A0(new_n15733_), .A1(new_n11768_), .B0(new_n15734_), .Y(new_n15735_));
  OAI21X1  g13299(.A0(new_n15632_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n15736_));
  AOI21X1  g13300(.A0(new_n15735_), .A1(new_n12486_), .B0(new_n15736_), .Y(new_n15737_));
  NAND2X1  g13301(.A(new_n15667_), .B(new_n12494_), .Y(new_n15738_));
  OAI21X1  g13302(.A0(new_n15632_), .A1(pi0618), .B0(pi1154), .Y(new_n15739_));
  AOI21X1  g13303(.A0(new_n15735_), .A1(pi0618), .B0(new_n15739_), .Y(new_n15740_));
  NAND2X1  g13304(.A(new_n15669_), .B(pi0627), .Y(new_n15741_));
  OAI22X1  g13305(.A0(new_n15741_), .A1(new_n15740_), .B0(new_n15738_), .B1(new_n15737_), .Y(new_n15742_));
  MX2X1    g13306(.A(new_n15742_), .B(new_n15735_), .S0(new_n11767_), .Y(new_n15743_));
  NAND2X1  g13307(.A(new_n15743_), .B(new_n12509_), .Y(new_n15744_));
  AOI21X1  g13308(.A0(new_n15634_), .A1(pi0619), .B0(pi1159), .Y(new_n15745_));
  NAND2X1  g13309(.A(new_n15674_), .B(new_n12517_), .Y(new_n15746_));
  AOI21X1  g13310(.A0(new_n15745_), .A1(new_n15744_), .B0(new_n15746_), .Y(new_n15747_));
  NAND2X1  g13311(.A(new_n15743_), .B(pi0619), .Y(new_n15748_));
  AOI21X1  g13312(.A0(new_n15634_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n15749_));
  NAND2X1  g13313(.A(new_n15676_), .B(pi0648), .Y(new_n15750_));
  AOI21X1  g13314(.A0(new_n15749_), .A1(new_n15748_), .B0(new_n15750_), .Y(new_n15751_));
  NOR3X1   g13315(.A(new_n15751_), .B(new_n15747_), .C(new_n11766_), .Y(new_n15752_));
  OAI21X1  g13316(.A0(new_n15743_), .A1(pi0789), .B0(new_n12709_), .Y(new_n15753_));
  OR2X1    g13317(.A(new_n15753_), .B(new_n15752_), .Y(new_n15754_));
  OAI22X1  g13318(.A0(new_n15686_), .A1(new_n12562_), .B0(new_n15636_), .B1(new_n13439_), .Y(new_n15755_));
  AOI21X1  g13319(.A0(new_n15755_), .A1(pi0788), .B0(new_n14125_), .Y(new_n15756_));
  AOI22X1  g13320(.A0(new_n15756_), .A1(new_n15754_), .B0(new_n15697_), .B1(pi0792), .Y(new_n15757_));
  OAI21X1  g13321(.A0(new_n15757_), .A1(new_n14121_), .B0(new_n15695_), .Y(new_n15758_));
  NOR2X1   g13322(.A(new_n15758_), .B(pi0644), .Y(new_n15759_));
  AND2X1   g13323(.A(new_n15647_), .B(pi0644), .Y(new_n15760_));
  OR2X1    g13324(.A(new_n15760_), .B(pi0715), .Y(new_n15761_));
  OAI21X1  g13325(.A0(new_n15616_), .A1(new_n12612_), .B0(pi0715), .Y(new_n15762_));
  AOI21X1  g13326(.A0(new_n15689_), .A1(new_n12612_), .B0(new_n15762_), .Y(new_n15763_));
  NOR2X1   g13327(.A(new_n15763_), .B(pi1160), .Y(new_n15764_));
  OAI21X1  g13328(.A0(new_n15761_), .A1(new_n15759_), .B0(new_n15764_), .Y(new_n15765_));
  AOI21X1  g13329(.A0(new_n15765_), .A1(new_n15692_), .B0(new_n12766_), .Y(new_n15766_));
  OR3X1    g13330(.A(new_n15691_), .B(new_n11762_), .C(new_n12612_), .Y(new_n15767_));
  AOI21X1  g13331(.A0(new_n15767_), .A1(pi0790), .B0(new_n15758_), .Y(new_n15768_));
  OAI21X1  g13332(.A0(new_n15768_), .A1(new_n15766_), .B0(new_n6489_), .Y(new_n15769_));
  AOI21X1  g13333(.A0(po1038), .A1(new_n9903_), .B0(pi0832), .Y(new_n15770_));
  NAND3X1  g13334(.A(new_n12470_), .B(new_n2720_), .C(pi0778), .Y(new_n15771_));
  AOI21X1  g13335(.A0(pi1093), .A1(pi1092), .B0(pi0173), .Y(new_n15772_));
  AOI21X1  g13336(.A0(new_n12056_), .A1(new_n14715_), .B0(new_n15772_), .Y(new_n15773_));
  INVX1    g13337(.A(new_n15773_), .Y(new_n15774_));
  NAND2X1  g13338(.A(new_n15774_), .B(new_n15771_), .Y(new_n15775_));
  AND3X1   g13339(.A(new_n12480_), .B(new_n12056_), .C(new_n14715_), .Y(new_n15776_));
  OAI21X1  g13340(.A0(new_n15776_), .A1(new_n15775_), .B0(pi1155), .Y(new_n15777_));
  OR3X1    g13341(.A(new_n15776_), .B(new_n15772_), .C(pi1155), .Y(new_n15778_));
  AOI21X1  g13342(.A0(new_n15778_), .A1(new_n15777_), .B0(new_n11768_), .Y(new_n15779_));
  AOI21X1  g13343(.A0(new_n15775_), .A1(new_n11768_), .B0(new_n15779_), .Y(new_n15780_));
  AOI21X1  g13344(.A0(new_n15780_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n15781_));
  AOI21X1  g13345(.A0(new_n15780_), .A1(new_n12655_), .B0(pi1154), .Y(new_n15782_));
  NOR2X1   g13346(.A(new_n15782_), .B(new_n15781_), .Y(new_n15783_));
  MX2X1    g13347(.A(new_n15783_), .B(new_n15780_), .S0(new_n11767_), .Y(new_n15784_));
  NOR2X1   g13348(.A(new_n15784_), .B(pi0789), .Y(new_n15785_));
  AND2X1   g13349(.A(new_n2720_), .B(new_n12509_), .Y(new_n15786_));
  INVX1    g13350(.A(new_n15786_), .Y(new_n15787_));
  AOI21X1  g13351(.A0(new_n15787_), .A1(new_n15784_), .B0(new_n12510_), .Y(new_n15788_));
  AND3X1   g13352(.A(pi1093), .B(pi1092), .C(pi0619), .Y(new_n15789_));
  INVX1    g13353(.A(new_n15789_), .Y(new_n15790_));
  AOI21X1  g13354(.A0(new_n15790_), .A1(new_n15784_), .B0(pi1159), .Y(new_n15791_));
  OR2X1    g13355(.A(new_n15791_), .B(new_n15788_), .Y(new_n15792_));
  AOI21X1  g13356(.A0(new_n15792_), .A1(pi0789), .B0(new_n15785_), .Y(new_n15793_));
  INVX1    g13357(.A(new_n15793_), .Y(new_n15794_));
  AOI21X1  g13358(.A0(new_n15772_), .A1(new_n12542_), .B0(new_n12548_), .Y(new_n15795_));
  OAI21X1  g13359(.A0(new_n15794_), .A1(new_n12542_), .B0(new_n15795_), .Y(new_n15796_));
  AOI21X1  g13360(.A0(new_n15772_), .A1(pi0626), .B0(pi1158), .Y(new_n15797_));
  OAI21X1  g13361(.A0(new_n15794_), .A1(pi0626), .B0(new_n15797_), .Y(new_n15798_));
  AND2X1   g13362(.A(new_n15798_), .B(new_n15796_), .Y(new_n15799_));
  MX2X1    g13363(.A(new_n15799_), .B(new_n15793_), .S0(new_n11765_), .Y(new_n15800_));
  AND3X1   g13364(.A(new_n15772_), .B(new_n12579_), .C(pi0792), .Y(new_n15801_));
  AOI21X1  g13365(.A0(new_n15800_), .A1(new_n14327_), .B0(new_n15801_), .Y(new_n15802_));
  AOI21X1  g13366(.A0(new_n12439_), .A1(new_n14743_), .B0(new_n15772_), .Y(new_n15803_));
  OR2X1    g13367(.A(new_n15803_), .B(pi0778), .Y(new_n15804_));
  INVX1    g13368(.A(new_n15803_), .Y(new_n15805_));
  AND3X1   g13369(.A(new_n12439_), .B(new_n14743_), .C(new_n12363_), .Y(new_n15806_));
  INVX1    g13370(.A(new_n15806_), .Y(new_n15807_));
  AOI21X1  g13371(.A0(new_n15807_), .A1(new_n15805_), .B0(new_n12364_), .Y(new_n15808_));
  NOR3X1   g13372(.A(new_n15806_), .B(new_n15772_), .C(pi1153), .Y(new_n15809_));
  OR3X1    g13373(.A(new_n15809_), .B(new_n15808_), .C(new_n11769_), .Y(new_n15810_));
  AND2X1   g13374(.A(new_n15810_), .B(new_n15804_), .Y(new_n15811_));
  NOR3X1   g13375(.A(new_n15811_), .B(new_n12631_), .C(new_n12630_), .Y(new_n15812_));
  AND3X1   g13376(.A(new_n15812_), .B(new_n12718_), .C(new_n12634_), .Y(new_n15813_));
  AND2X1   g13377(.A(new_n15813_), .B(new_n12739_), .Y(new_n15814_));
  INVX1    g13378(.A(new_n15814_), .Y(new_n15815_));
  AOI21X1  g13379(.A0(new_n15772_), .A1(pi0647), .B0(pi1157), .Y(new_n15816_));
  OAI21X1  g13380(.A0(new_n15815_), .A1(pi0647), .B0(new_n15816_), .Y(new_n15817_));
  MX2X1    g13381(.A(new_n15814_), .B(new_n15772_), .S0(new_n12577_), .Y(new_n15818_));
  OAI22X1  g13382(.A0(new_n15818_), .A1(new_n14242_), .B0(new_n15817_), .B1(new_n12592_), .Y(new_n15819_));
  AOI21X1  g13383(.A0(new_n15802_), .A1(new_n14326_), .B0(new_n15819_), .Y(new_n15820_));
  AND3X1   g13384(.A(new_n15812_), .B(new_n12637_), .C(new_n12634_), .Y(new_n15821_));
  AND3X1   g13385(.A(new_n15798_), .B(new_n15796_), .C(new_n12639_), .Y(new_n15822_));
  OR2X1    g13386(.A(new_n15822_), .B(new_n15821_), .Y(new_n15823_));
  AOI21X1  g13387(.A0(new_n15805_), .A1(new_n12048_), .B0(new_n15774_), .Y(new_n15824_));
  NOR2X1   g13388(.A(new_n15772_), .B(pi1153), .Y(new_n15825_));
  NOR3X1   g13389(.A(new_n15803_), .B(new_n11991_), .C(new_n12363_), .Y(new_n15826_));
  OAI21X1  g13390(.A0(new_n15824_), .A1(new_n15826_), .B0(new_n15825_), .Y(new_n15827_));
  NOR2X1   g13391(.A(new_n15808_), .B(pi0608), .Y(new_n15828_));
  NOR3X1   g13392(.A(new_n15826_), .B(new_n15774_), .C(new_n12364_), .Y(new_n15829_));
  NOR3X1   g13393(.A(new_n15829_), .B(new_n15809_), .C(new_n12368_), .Y(new_n15830_));
  AOI21X1  g13394(.A0(new_n15828_), .A1(new_n15827_), .B0(new_n15830_), .Y(new_n15831_));
  OR2X1    g13395(.A(new_n15831_), .B(new_n11769_), .Y(new_n15832_));
  OAI21X1  g13396(.A0(new_n15824_), .A1(pi0778), .B0(new_n15832_), .Y(new_n15833_));
  INVX1    g13397(.A(new_n15833_), .Y(new_n15834_));
  INVX1    g13398(.A(new_n15811_), .Y(new_n15835_));
  AOI21X1  g13399(.A0(new_n15835_), .A1(pi0609), .B0(pi1155), .Y(new_n15836_));
  OAI21X1  g13400(.A0(new_n15834_), .A1(pi0609), .B0(new_n15836_), .Y(new_n15837_));
  AND3X1   g13401(.A(new_n15837_), .B(new_n15777_), .C(new_n12468_), .Y(new_n15838_));
  AOI21X1  g13402(.A0(new_n15835_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n15839_));
  OAI21X1  g13403(.A0(new_n15834_), .A1(new_n12462_), .B0(new_n15839_), .Y(new_n15840_));
  AND3X1   g13404(.A(new_n15840_), .B(new_n15778_), .C(pi0660), .Y(new_n15841_));
  NOR2X1   g13405(.A(new_n15841_), .B(new_n15838_), .Y(new_n15842_));
  MX2X1    g13406(.A(new_n15842_), .B(new_n15834_), .S0(new_n11768_), .Y(new_n15843_));
  AOI21X1  g13407(.A0(new_n15810_), .A1(new_n15804_), .B0(new_n12630_), .Y(new_n15844_));
  AOI21X1  g13408(.A0(new_n15844_), .A1(pi0618), .B0(pi1154), .Y(new_n15845_));
  OAI21X1  g13409(.A0(new_n15843_), .A1(pi0618), .B0(new_n15845_), .Y(new_n15846_));
  NOR2X1   g13410(.A(new_n15781_), .B(pi0627), .Y(new_n15847_));
  AOI21X1  g13411(.A0(new_n15844_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n15848_));
  OAI21X1  g13412(.A0(new_n15843_), .A1(new_n12486_), .B0(new_n15848_), .Y(new_n15849_));
  NOR2X1   g13413(.A(new_n15782_), .B(new_n12494_), .Y(new_n15850_));
  AOI22X1  g13414(.A0(new_n15850_), .A1(new_n15849_), .B0(new_n15847_), .B1(new_n15846_), .Y(new_n15851_));
  MX2X1    g13415(.A(new_n15851_), .B(new_n15843_), .S0(new_n11767_), .Y(new_n15852_));
  AOI21X1  g13416(.A0(new_n15812_), .A1(pi0619), .B0(pi1159), .Y(new_n15853_));
  OAI21X1  g13417(.A0(new_n15852_), .A1(pi0619), .B0(new_n15853_), .Y(new_n15854_));
  NOR2X1   g13418(.A(new_n15788_), .B(pi0648), .Y(new_n15855_));
  AND2X1   g13419(.A(new_n15855_), .B(new_n15854_), .Y(new_n15856_));
  AOI21X1  g13420(.A0(new_n15812_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n15857_));
  OAI21X1  g13421(.A0(new_n15852_), .A1(new_n12509_), .B0(new_n15857_), .Y(new_n15858_));
  NOR2X1   g13422(.A(new_n15791_), .B(new_n12517_), .Y(new_n15859_));
  AND2X1   g13423(.A(new_n15859_), .B(new_n15858_), .Y(new_n15860_));
  OR3X1    g13424(.A(new_n15860_), .B(new_n15856_), .C(new_n11766_), .Y(new_n15861_));
  AOI21X1  g13425(.A0(new_n15852_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n15862_));
  AOI22X1  g13426(.A0(new_n15862_), .A1(new_n15861_), .B0(new_n15823_), .B1(pi0788), .Y(new_n15863_));
  NOR2X1   g13427(.A(new_n15863_), .B(new_n14125_), .Y(new_n15864_));
  AOI22X1  g13428(.A0(new_n15813_), .A1(new_n14426_), .B0(new_n15800_), .B1(new_n12735_), .Y(new_n15865_));
  AOI22X1  g13429(.A0(new_n15813_), .A1(new_n14428_), .B0(new_n15800_), .B1(new_n12733_), .Y(new_n15866_));
  MX2X1    g13430(.A(new_n15866_), .B(new_n15865_), .S0(new_n12561_), .Y(new_n15867_));
  OAI21X1  g13431(.A0(new_n15867_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n15868_));
  OAI22X1  g13432(.A0(new_n15868_), .A1(new_n15864_), .B0(new_n15820_), .B1(new_n11763_), .Y(new_n15869_));
  INVX1    g13433(.A(new_n15869_), .Y(new_n15870_));
  OAI21X1  g13434(.A0(new_n15818_), .A1(new_n12578_), .B0(new_n15817_), .Y(new_n15871_));
  MX2X1    g13435(.A(new_n15871_), .B(new_n15815_), .S0(new_n11763_), .Y(new_n15872_));
  OAI21X1  g13436(.A0(new_n15872_), .A1(pi0644), .B0(pi0715), .Y(new_n15873_));
  AOI21X1  g13437(.A0(new_n15870_), .A1(pi0644), .B0(new_n15873_), .Y(new_n15874_));
  INVX1    g13438(.A(new_n15772_), .Y(new_n15875_));
  OR3X1    g13439(.A(new_n15875_), .B(new_n12603_), .C(new_n11763_), .Y(new_n15876_));
  OAI21X1  g13440(.A0(new_n15802_), .A1(new_n12604_), .B0(new_n15876_), .Y(new_n15877_));
  OAI21X1  g13441(.A0(new_n15875_), .A1(pi0644), .B0(new_n12608_), .Y(new_n15878_));
  AOI21X1  g13442(.A0(new_n15877_), .A1(pi0644), .B0(new_n15878_), .Y(new_n15879_));
  OR2X1    g13443(.A(new_n15879_), .B(new_n11762_), .Y(new_n15880_));
  OAI21X1  g13444(.A0(new_n15872_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n15881_));
  AOI21X1  g13445(.A0(new_n15870_), .A1(new_n12612_), .B0(new_n15881_), .Y(new_n15882_));
  OAI21X1  g13446(.A0(new_n15875_), .A1(new_n12612_), .B0(pi0715), .Y(new_n15883_));
  AOI21X1  g13447(.A0(new_n15877_), .A1(new_n12612_), .B0(new_n15883_), .Y(new_n15884_));
  OR2X1    g13448(.A(new_n15884_), .B(pi1160), .Y(new_n15885_));
  OAI22X1  g13449(.A0(new_n15885_), .A1(new_n15882_), .B0(new_n15880_), .B1(new_n15874_), .Y(new_n15886_));
  OAI21X1  g13450(.A0(new_n15869_), .A1(pi0790), .B0(pi0832), .Y(new_n15887_));
  AOI21X1  g13451(.A0(new_n15886_), .A1(pi0790), .B0(new_n15887_), .Y(new_n15888_));
  AOI21X1  g13452(.A0(new_n15770_), .A1(new_n15769_), .B0(new_n15888_), .Y(po0330));
  AND2X1   g13453(.A(new_n12034_), .B(pi0759), .Y(new_n15890_));
  OAI21X1  g13454(.A0(new_n15890_), .A1(new_n14823_), .B0(pi0039), .Y(new_n15891_));
  AOI21X1  g13455(.A0(new_n11821_), .A1(new_n14767_), .B0(pi0039), .Y(new_n15892_));
  OAI21X1  g13456(.A0(new_n11975_), .A1(new_n14767_), .B0(new_n15892_), .Y(new_n15893_));
  AOI21X1  g13457(.A0(new_n15893_), .A1(new_n15891_), .B0(new_n6851_), .Y(new_n15894_));
  AND3X1   g13458(.A(new_n12074_), .B(pi0759), .C(new_n6851_), .Y(new_n15895_));
  OAI21X1  g13459(.A0(new_n15895_), .A1(new_n15894_), .B0(new_n2979_), .Y(new_n15896_));
  NOR2X1   g13460(.A(new_n12077_), .B(pi0174), .Y(new_n15897_));
  AOI21X1  g13461(.A0(new_n11991_), .A1(pi0759), .B0(new_n12771_), .Y(new_n15898_));
  NOR3X1   g13462(.A(new_n15898_), .B(new_n15897_), .C(new_n2979_), .Y(new_n15899_));
  INVX1    g13463(.A(new_n15899_), .Y(new_n15900_));
  AND3X1   g13464(.A(new_n15900_), .B(new_n15896_), .C(new_n14807_), .Y(new_n15901_));
  AOI21X1  g13465(.A0(new_n12213_), .A1(new_n6851_), .B0(pi0759), .Y(new_n15902_));
  OAI21X1  g13466(.A0(new_n12155_), .A1(new_n6851_), .B0(new_n15902_), .Y(new_n15903_));
  AOI21X1  g13467(.A0(new_n12301_), .A1(pi0174), .B0(new_n14767_), .Y(new_n15904_));
  OAI21X1  g13468(.A0(new_n12260_), .A1(pi0174), .B0(new_n15904_), .Y(new_n15905_));
  AND3X1   g13469(.A(new_n15905_), .B(new_n15903_), .C(pi0039), .Y(new_n15906_));
  OAI21X1  g13470(.A0(new_n12315_), .A1(new_n6851_), .B0(new_n14767_), .Y(new_n15907_));
  AOI21X1  g13471(.A0(new_n12332_), .A1(new_n6851_), .B0(new_n15907_), .Y(new_n15908_));
  NOR4X1   g13472(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(new_n6851_), .Y(new_n15909_));
  OAI21X1  g13473(.A0(new_n12800_), .A1(pi0174), .B0(pi0759), .Y(new_n15910_));
  OAI21X1  g13474(.A0(new_n15910_), .A1(new_n15909_), .B0(new_n2939_), .Y(new_n15911_));
  OAI21X1  g13475(.A0(new_n15911_), .A1(new_n15908_), .B0(new_n2979_), .Y(new_n15912_));
  NOR3X1   g13476(.A(new_n15899_), .B(new_n13547_), .C(new_n14807_), .Y(new_n15913_));
  OAI21X1  g13477(.A0(new_n15912_), .A1(new_n15906_), .B0(new_n15913_), .Y(new_n15914_));
  NAND2X1  g13478(.A(new_n15914_), .B(new_n3103_), .Y(new_n15915_));
  OAI22X1  g13479(.A0(new_n15915_), .A1(new_n15901_), .B0(new_n3103_), .B1(new_n6851_), .Y(new_n15916_));
  OR2X1    g13480(.A(new_n15916_), .B(pi0625), .Y(new_n15917_));
  AND2X1   g13481(.A(new_n15900_), .B(new_n15896_), .Y(new_n15918_));
  MX2X1    g13482(.A(new_n15918_), .B(new_n6851_), .S0(new_n11770_), .Y(new_n15919_));
  AOI21X1  g13483(.A0(new_n15919_), .A1(pi0625), .B0(pi1153), .Y(new_n15920_));
  AOI21X1  g13484(.A0(new_n12447_), .A1(new_n3103_), .B0(new_n6851_), .Y(new_n15921_));
  NOR4X1   g13485(.A(new_n10543_), .B(new_n14807_), .C(pi0100), .D(pi0087), .Y(new_n15922_));
  OAI21X1  g13486(.A0(new_n13870_), .A1(pi0174), .B0(new_n2979_), .Y(new_n15923_));
  AOI21X1  g13487(.A0(new_n13868_), .A1(pi0174), .B0(new_n15923_), .Y(new_n15924_));
  OAI21X1  g13488(.A0(new_n15897_), .A1(new_n13874_), .B0(new_n15922_), .Y(new_n15925_));
  OAI22X1  g13489(.A0(new_n15925_), .A1(new_n15924_), .B0(new_n15922_), .B1(new_n15921_), .Y(new_n15926_));
  OAI21X1  g13490(.A0(new_n15921_), .A1(pi0625), .B0(pi1153), .Y(new_n15927_));
  AOI21X1  g13491(.A0(new_n15926_), .A1(pi0625), .B0(new_n15927_), .Y(new_n15928_));
  OR2X1    g13492(.A(new_n15928_), .B(pi0608), .Y(new_n15929_));
  AOI21X1  g13493(.A0(new_n15920_), .A1(new_n15917_), .B0(new_n15929_), .Y(new_n15930_));
  OR2X1    g13494(.A(new_n15916_), .B(new_n12363_), .Y(new_n15931_));
  AOI21X1  g13495(.A0(new_n15919_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n15932_));
  OAI21X1  g13496(.A0(new_n15921_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n15933_));
  AOI21X1  g13497(.A0(new_n15926_), .A1(new_n12363_), .B0(new_n15933_), .Y(new_n15934_));
  OR2X1    g13498(.A(new_n15934_), .B(new_n12368_), .Y(new_n15935_));
  AOI21X1  g13499(.A0(new_n15932_), .A1(new_n15931_), .B0(new_n15935_), .Y(new_n15936_));
  OAI21X1  g13500(.A0(new_n15936_), .A1(new_n15930_), .B0(pi0778), .Y(new_n15937_));
  OR2X1    g13501(.A(new_n15916_), .B(pi0778), .Y(new_n15938_));
  AOI21X1  g13502(.A0(new_n15938_), .A1(new_n15937_), .B0(pi0609), .Y(new_n15939_));
  OR2X1    g13503(.A(new_n15926_), .B(pi0778), .Y(new_n15940_));
  NOR2X1   g13504(.A(new_n15934_), .B(new_n15928_), .Y(new_n15941_));
  OAI21X1  g13505(.A0(new_n15941_), .A1(new_n11769_), .B0(new_n15940_), .Y(new_n15942_));
  OAI21X1  g13506(.A0(new_n15942_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n15943_));
  NOR2X1   g13507(.A(new_n15921_), .B(new_n12474_), .Y(new_n15944_));
  AOI21X1  g13508(.A0(new_n15919_), .A1(new_n12474_), .B0(new_n15944_), .Y(new_n15945_));
  INVX1    g13509(.A(new_n15921_), .Y(new_n15946_));
  AOI21X1  g13510(.A0(new_n15946_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n15947_));
  OAI21X1  g13511(.A0(new_n15945_), .A1(new_n12462_), .B0(new_n15947_), .Y(new_n15948_));
  AND2X1   g13512(.A(new_n15948_), .B(new_n12468_), .Y(new_n15949_));
  OAI21X1  g13513(.A0(new_n15943_), .A1(new_n15939_), .B0(new_n15949_), .Y(new_n15950_));
  AOI21X1  g13514(.A0(new_n15938_), .A1(new_n15937_), .B0(new_n12462_), .Y(new_n15951_));
  OAI21X1  g13515(.A0(new_n15942_), .A1(pi0609), .B0(pi1155), .Y(new_n15952_));
  AOI21X1  g13516(.A0(new_n15946_), .A1(pi0609), .B0(pi1155), .Y(new_n15953_));
  OAI21X1  g13517(.A0(new_n15945_), .A1(pi0609), .B0(new_n15953_), .Y(new_n15954_));
  AND2X1   g13518(.A(new_n15954_), .B(pi0660), .Y(new_n15955_));
  OAI21X1  g13519(.A0(new_n15952_), .A1(new_n15951_), .B0(new_n15955_), .Y(new_n15956_));
  AOI21X1  g13520(.A0(new_n15956_), .A1(new_n15950_), .B0(new_n11768_), .Y(new_n15957_));
  AOI21X1  g13521(.A0(new_n15938_), .A1(new_n15937_), .B0(pi0785), .Y(new_n15958_));
  OAI21X1  g13522(.A0(new_n15958_), .A1(new_n15957_), .B0(new_n12486_), .Y(new_n15959_));
  OR2X1    g13523(.A(new_n15921_), .B(new_n13910_), .Y(new_n15960_));
  OAI21X1  g13524(.A0(new_n15942_), .A1(new_n12490_), .B0(new_n15960_), .Y(new_n15961_));
  AOI21X1  g13525(.A0(new_n15961_), .A1(pi0618), .B0(pi1154), .Y(new_n15962_));
  AOI21X1  g13526(.A0(new_n15954_), .A1(new_n15948_), .B0(new_n11768_), .Y(new_n15963_));
  AOI21X1  g13527(.A0(new_n15945_), .A1(new_n11768_), .B0(new_n15963_), .Y(new_n15964_));
  OAI21X1  g13528(.A0(new_n15921_), .A1(pi0618), .B0(pi1154), .Y(new_n15965_));
  AOI21X1  g13529(.A0(new_n15964_), .A1(pi0618), .B0(new_n15965_), .Y(new_n15966_));
  OR2X1    g13530(.A(new_n15966_), .B(pi0627), .Y(new_n15967_));
  AOI21X1  g13531(.A0(new_n15962_), .A1(new_n15959_), .B0(new_n15967_), .Y(new_n15968_));
  OAI21X1  g13532(.A0(new_n15958_), .A1(new_n15957_), .B0(pi0618), .Y(new_n15969_));
  AOI21X1  g13533(.A0(new_n15961_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n15970_));
  OAI21X1  g13534(.A0(new_n15921_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n15971_));
  AOI21X1  g13535(.A0(new_n15964_), .A1(new_n12486_), .B0(new_n15971_), .Y(new_n15972_));
  OR2X1    g13536(.A(new_n15972_), .B(new_n12494_), .Y(new_n15973_));
  AOI21X1  g13537(.A0(new_n15970_), .A1(new_n15969_), .B0(new_n15973_), .Y(new_n15974_));
  OAI21X1  g13538(.A0(new_n15974_), .A1(new_n15968_), .B0(pi0781), .Y(new_n15975_));
  OAI21X1  g13539(.A0(new_n15958_), .A1(new_n15957_), .B0(new_n11767_), .Y(new_n15976_));
  AOI21X1  g13540(.A0(new_n15976_), .A1(new_n15975_), .B0(pi0619), .Y(new_n15977_));
  MX2X1    g13541(.A(new_n15961_), .B(new_n15946_), .S0(new_n12513_), .Y(new_n15978_));
  INVX1    g13542(.A(new_n15978_), .Y(new_n15979_));
  OAI21X1  g13543(.A0(new_n15979_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n15980_));
  OAI21X1  g13544(.A0(new_n15972_), .A1(new_n15966_), .B0(pi0781), .Y(new_n15981_));
  OAI21X1  g13545(.A0(new_n15964_), .A1(pi0781), .B0(new_n15981_), .Y(new_n15982_));
  AOI21X1  g13546(.A0(new_n15946_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n15983_));
  OAI21X1  g13547(.A0(new_n15982_), .A1(new_n12509_), .B0(new_n15983_), .Y(new_n15984_));
  AND2X1   g13548(.A(new_n15984_), .B(new_n12517_), .Y(new_n15985_));
  OAI21X1  g13549(.A0(new_n15980_), .A1(new_n15977_), .B0(new_n15985_), .Y(new_n15986_));
  AOI21X1  g13550(.A0(new_n15976_), .A1(new_n15975_), .B0(new_n12509_), .Y(new_n15987_));
  OAI21X1  g13551(.A0(new_n15979_), .A1(pi0619), .B0(pi1159), .Y(new_n15988_));
  AOI21X1  g13552(.A0(new_n15946_), .A1(pi0619), .B0(pi1159), .Y(new_n15989_));
  OAI21X1  g13553(.A0(new_n15982_), .A1(pi0619), .B0(new_n15989_), .Y(new_n15990_));
  AND2X1   g13554(.A(new_n15990_), .B(pi0648), .Y(new_n15991_));
  OAI21X1  g13555(.A0(new_n15988_), .A1(new_n15987_), .B0(new_n15991_), .Y(new_n15992_));
  AOI21X1  g13556(.A0(new_n15992_), .A1(new_n15986_), .B0(new_n11766_), .Y(new_n15993_));
  AOI21X1  g13557(.A0(new_n15976_), .A1(new_n15975_), .B0(pi0789), .Y(new_n15994_));
  OR3X1    g13558(.A(new_n15994_), .B(new_n15993_), .C(pi0788), .Y(new_n15995_));
  OR3X1    g13559(.A(new_n15994_), .B(new_n15993_), .C(pi0626), .Y(new_n15996_));
  MX2X1    g13560(.A(new_n15979_), .B(new_n15921_), .S0(new_n12531_), .Y(new_n15997_));
  AOI21X1  g13561(.A0(new_n15997_), .A1(pi0626), .B0(pi0641), .Y(new_n15998_));
  NAND2X1  g13562(.A(new_n15990_), .B(new_n15984_), .Y(new_n15999_));
  MX2X1    g13563(.A(new_n15999_), .B(new_n15982_), .S0(new_n11766_), .Y(new_n16000_));
  OAI21X1  g13564(.A0(new_n15946_), .A1(new_n12542_), .B0(pi0641), .Y(new_n16001_));
  AOI21X1  g13565(.A0(new_n16000_), .A1(new_n12542_), .B0(new_n16001_), .Y(new_n16002_));
  OR2X1    g13566(.A(new_n16002_), .B(pi1158), .Y(new_n16003_));
  AOI21X1  g13567(.A0(new_n15998_), .A1(new_n15996_), .B0(new_n16003_), .Y(new_n16004_));
  OR3X1    g13568(.A(new_n15994_), .B(new_n15993_), .C(new_n12542_), .Y(new_n16005_));
  AOI21X1  g13569(.A0(new_n15997_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n16006_));
  OAI21X1  g13570(.A0(new_n15946_), .A1(pi0626), .B0(new_n12543_), .Y(new_n16007_));
  AOI21X1  g13571(.A0(new_n16000_), .A1(pi0626), .B0(new_n16007_), .Y(new_n16008_));
  OR2X1    g13572(.A(new_n16008_), .B(new_n12548_), .Y(new_n16009_));
  AOI21X1  g13573(.A0(new_n16006_), .A1(new_n16005_), .B0(new_n16009_), .Y(new_n16010_));
  OAI21X1  g13574(.A0(new_n16010_), .A1(new_n16004_), .B0(pi0788), .Y(new_n16011_));
  AND3X1   g13575(.A(new_n16011_), .B(new_n15995_), .C(new_n12554_), .Y(new_n16012_));
  MX2X1    g13576(.A(new_n16000_), .B(new_n15921_), .S0(new_n12708_), .Y(new_n16013_));
  OAI21X1  g13577(.A0(new_n16013_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n16014_));
  AND2X1   g13578(.A(new_n15921_), .B(new_n12563_), .Y(new_n16015_));
  AOI21X1  g13579(.A0(new_n15997_), .A1(new_n13356_), .B0(new_n16015_), .Y(new_n16016_));
  OAI21X1  g13580(.A0(new_n15921_), .A1(pi0628), .B0(pi1156), .Y(new_n16017_));
  AOI21X1  g13581(.A0(new_n16016_), .A1(pi0628), .B0(new_n16017_), .Y(new_n16018_));
  NOR2X1   g13582(.A(new_n16018_), .B(pi0629), .Y(new_n16019_));
  OAI21X1  g13583(.A0(new_n16014_), .A1(new_n16012_), .B0(new_n16019_), .Y(new_n16020_));
  AND3X1   g13584(.A(new_n16011_), .B(new_n15995_), .C(pi0628), .Y(new_n16021_));
  OAI21X1  g13585(.A0(new_n16013_), .A1(pi0628), .B0(pi1156), .Y(new_n16022_));
  OAI21X1  g13586(.A0(new_n15921_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n16023_));
  AOI21X1  g13587(.A0(new_n16016_), .A1(new_n12554_), .B0(new_n16023_), .Y(new_n16024_));
  NOR2X1   g13588(.A(new_n16024_), .B(new_n12561_), .Y(new_n16025_));
  OAI21X1  g13589(.A0(new_n16022_), .A1(new_n16021_), .B0(new_n16025_), .Y(new_n16026_));
  AOI21X1  g13590(.A0(new_n16026_), .A1(new_n16020_), .B0(new_n11764_), .Y(new_n16027_));
  AND3X1   g13591(.A(new_n16011_), .B(new_n15995_), .C(new_n11764_), .Y(new_n16028_));
  OAI21X1  g13592(.A0(new_n16028_), .A1(new_n16027_), .B0(new_n12577_), .Y(new_n16029_));
  MX2X1    g13593(.A(new_n16013_), .B(new_n15921_), .S0(new_n12580_), .Y(new_n16030_));
  INVX1    g13594(.A(new_n16030_), .Y(new_n16031_));
  AOI21X1  g13595(.A0(new_n16031_), .A1(pi0647), .B0(pi1157), .Y(new_n16032_));
  NOR2X1   g13596(.A(new_n16024_), .B(new_n16018_), .Y(new_n16033_));
  MX2X1    g13597(.A(new_n16033_), .B(new_n16016_), .S0(new_n11764_), .Y(new_n16034_));
  OAI21X1  g13598(.A0(new_n15921_), .A1(pi0647), .B0(pi1157), .Y(new_n16035_));
  AOI21X1  g13599(.A0(new_n16034_), .A1(pi0647), .B0(new_n16035_), .Y(new_n16036_));
  OR2X1    g13600(.A(new_n16036_), .B(pi0630), .Y(new_n16037_));
  AOI21X1  g13601(.A0(new_n16032_), .A1(new_n16029_), .B0(new_n16037_), .Y(new_n16038_));
  OAI21X1  g13602(.A0(new_n16028_), .A1(new_n16027_), .B0(pi0647), .Y(new_n16039_));
  AOI21X1  g13603(.A0(new_n16031_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n16040_));
  OAI21X1  g13604(.A0(new_n15921_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n16041_));
  AOI21X1  g13605(.A0(new_n16034_), .A1(new_n12577_), .B0(new_n16041_), .Y(new_n16042_));
  OR2X1    g13606(.A(new_n16042_), .B(new_n12592_), .Y(new_n16043_));
  AOI21X1  g13607(.A0(new_n16040_), .A1(new_n16039_), .B0(new_n16043_), .Y(new_n16044_));
  OAI21X1  g13608(.A0(new_n16044_), .A1(new_n16038_), .B0(pi0787), .Y(new_n16045_));
  OAI21X1  g13609(.A0(new_n16028_), .A1(new_n16027_), .B0(new_n11763_), .Y(new_n16046_));
  AOI21X1  g13610(.A0(new_n16046_), .A1(new_n16045_), .B0(new_n12612_), .Y(new_n16047_));
  OAI21X1  g13611(.A0(new_n16042_), .A1(new_n16036_), .B0(pi0787), .Y(new_n16048_));
  OAI21X1  g13612(.A0(new_n16034_), .A1(pi0787), .B0(new_n16048_), .Y(new_n16049_));
  OAI21X1  g13613(.A0(new_n16049_), .A1(pi0644), .B0(pi0715), .Y(new_n16050_));
  MX2X1    g13614(.A(new_n16030_), .B(new_n15921_), .S0(new_n12604_), .Y(new_n16051_));
  AOI21X1  g13615(.A0(new_n15946_), .A1(new_n12612_), .B0(pi0715), .Y(new_n16052_));
  OAI21X1  g13616(.A0(new_n16051_), .A1(new_n12612_), .B0(new_n16052_), .Y(new_n16053_));
  AND2X1   g13617(.A(new_n16053_), .B(pi1160), .Y(new_n16054_));
  OAI21X1  g13618(.A0(new_n16050_), .A1(new_n16047_), .B0(new_n16054_), .Y(new_n16055_));
  AOI21X1  g13619(.A0(new_n16046_), .A1(new_n16045_), .B0(pi0644), .Y(new_n16056_));
  OAI21X1  g13620(.A0(new_n16049_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n16057_));
  AOI21X1  g13621(.A0(new_n15946_), .A1(pi0644), .B0(new_n12608_), .Y(new_n16058_));
  OAI21X1  g13622(.A0(new_n16051_), .A1(pi0644), .B0(new_n16058_), .Y(new_n16059_));
  AND2X1   g13623(.A(new_n16059_), .B(new_n11762_), .Y(new_n16060_));
  OAI21X1  g13624(.A0(new_n16057_), .A1(new_n16056_), .B0(new_n16060_), .Y(new_n16061_));
  AND3X1   g13625(.A(new_n16061_), .B(new_n16055_), .C(pi0790), .Y(new_n16062_));
  AND3X1   g13626(.A(new_n16046_), .B(new_n16045_), .C(new_n12766_), .Y(new_n16063_));
  OR2X1    g13627(.A(new_n16063_), .B(new_n5103_), .Y(new_n16064_));
  AOI21X1  g13628(.A0(new_n5103_), .A1(new_n6851_), .B0(pi0057), .Y(new_n16065_));
  OAI21X1  g13629(.A0(new_n16064_), .A1(new_n16062_), .B0(new_n16065_), .Y(new_n16066_));
  AOI21X1  g13630(.A0(pi0174), .A1(pi0057), .B0(pi0832), .Y(new_n16067_));
  NOR2X1   g13631(.A(new_n2720_), .B(new_n6851_), .Y(new_n16068_));
  AOI21X1  g13632(.A0(new_n12056_), .A1(pi0759), .B0(new_n16068_), .Y(new_n16069_));
  OAI21X1  g13633(.A0(new_n14068_), .A1(new_n14807_), .B0(new_n16069_), .Y(new_n16070_));
  AND3X1   g13634(.A(new_n13443_), .B(pi0696), .C(pi0625), .Y(new_n16071_));
  INVX1    g13635(.A(new_n16071_), .Y(new_n16072_));
  AOI21X1  g13636(.A0(new_n16072_), .A1(new_n16070_), .B0(pi1153), .Y(new_n16073_));
  AND3X1   g13637(.A(new_n12439_), .B(pi0696), .C(pi0625), .Y(new_n16074_));
  NOR3X1   g13638(.A(new_n16074_), .B(new_n16068_), .C(new_n12364_), .Y(new_n16075_));
  NOR3X1   g13639(.A(new_n16075_), .B(new_n16073_), .C(pi0608), .Y(new_n16076_));
  AOI21X1  g13640(.A0(new_n12439_), .A1(pi0696), .B0(new_n16068_), .Y(new_n16077_));
  OAI21X1  g13641(.A0(new_n16077_), .A1(new_n16074_), .B0(new_n12364_), .Y(new_n16078_));
  NAND3X1  g13642(.A(new_n16072_), .B(new_n16069_), .C(pi1153), .Y(new_n16079_));
  AND3X1   g13643(.A(new_n16079_), .B(new_n16078_), .C(pi0608), .Y(new_n16080_));
  OR2X1    g13644(.A(new_n16080_), .B(new_n16076_), .Y(new_n16081_));
  MX2X1    g13645(.A(new_n16081_), .B(new_n16070_), .S0(new_n11769_), .Y(new_n16082_));
  OAI21X1  g13646(.A0(new_n2720_), .A1(new_n6851_), .B0(pi1153), .Y(new_n16083_));
  OAI21X1  g13647(.A0(new_n16083_), .A1(new_n16074_), .B0(new_n16078_), .Y(new_n16084_));
  MX2X1    g13648(.A(new_n16084_), .B(new_n16077_), .S0(new_n11769_), .Y(new_n16085_));
  OAI21X1  g13649(.A0(new_n16085_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n16086_));
  AOI21X1  g13650(.A0(new_n16082_), .A1(new_n12462_), .B0(new_n16086_), .Y(new_n16087_));
  AND3X1   g13651(.A(new_n12471_), .B(new_n12056_), .C(pi0759), .Y(new_n16088_));
  OAI21X1  g13652(.A0(new_n2720_), .A1(new_n6851_), .B0(pi1155), .Y(new_n16089_));
  OAI21X1  g13653(.A0(new_n16089_), .A1(new_n16088_), .B0(new_n12468_), .Y(new_n16090_));
  OAI21X1  g13654(.A0(new_n16085_), .A1(pi0609), .B0(pi1155), .Y(new_n16091_));
  AOI21X1  g13655(.A0(new_n16082_), .A1(pi0609), .B0(new_n16091_), .Y(new_n16092_));
  AND3X1   g13656(.A(new_n12480_), .B(new_n12056_), .C(pi0759), .Y(new_n16093_));
  OAI21X1  g13657(.A0(new_n2720_), .A1(new_n6851_), .B0(new_n12463_), .Y(new_n16094_));
  OAI21X1  g13658(.A0(new_n16094_), .A1(new_n16093_), .B0(pi0660), .Y(new_n16095_));
  OAI22X1  g13659(.A0(new_n16095_), .A1(new_n16092_), .B0(new_n16090_), .B1(new_n16087_), .Y(new_n16096_));
  MX2X1    g13660(.A(new_n16096_), .B(new_n16082_), .S0(new_n11768_), .Y(new_n16097_));
  NAND2X1  g13661(.A(new_n16097_), .B(new_n12486_), .Y(new_n16098_));
  OAI22X1  g13662(.A0(new_n16085_), .A1(new_n12490_), .B0(new_n2720_), .B1(new_n6851_), .Y(new_n16099_));
  AOI21X1  g13663(.A0(new_n16099_), .A1(pi0618), .B0(pi1154), .Y(new_n16100_));
  OR3X1    g13664(.A(new_n14034_), .B(new_n12057_), .C(new_n14767_), .Y(new_n16101_));
  NOR3X1   g13665(.A(new_n16101_), .B(new_n12473_), .C(new_n12486_), .Y(new_n16102_));
  OAI21X1  g13666(.A0(new_n2720_), .A1(new_n6851_), .B0(pi1154), .Y(new_n16103_));
  OAI21X1  g13667(.A0(new_n16103_), .A1(new_n16102_), .B0(new_n12494_), .Y(new_n16104_));
  AOI21X1  g13668(.A0(new_n16100_), .A1(new_n16098_), .B0(new_n16104_), .Y(new_n16105_));
  NAND2X1  g13669(.A(new_n16097_), .B(pi0618), .Y(new_n16106_));
  AOI21X1  g13670(.A0(new_n16099_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n16107_));
  NOR3X1   g13671(.A(new_n16101_), .B(new_n12473_), .C(pi0618), .Y(new_n16108_));
  OAI21X1  g13672(.A0(new_n2720_), .A1(new_n6851_), .B0(new_n12487_), .Y(new_n16109_));
  OAI21X1  g13673(.A0(new_n16109_), .A1(new_n16108_), .B0(pi0627), .Y(new_n16110_));
  AOI21X1  g13674(.A0(new_n16107_), .A1(new_n16106_), .B0(new_n16110_), .Y(new_n16111_));
  OAI21X1  g13675(.A0(new_n16111_), .A1(new_n16105_), .B0(pi0781), .Y(new_n16112_));
  INVX1    g13676(.A(new_n12530_), .Y(new_n16113_));
  AND3X1   g13677(.A(pi1159), .B(pi0648), .C(new_n12509_), .Y(new_n16114_));
  AND3X1   g13678(.A(new_n12510_), .B(new_n12517_), .C(pi0619), .Y(new_n16115_));
  OR2X1    g13679(.A(new_n16115_), .B(new_n16114_), .Y(new_n16116_));
  NOR2X1   g13680(.A(new_n16116_), .B(new_n16113_), .Y(new_n16117_));
  NOR2X1   g13681(.A(new_n16117_), .B(new_n11766_), .Y(new_n16118_));
  AOI21X1  g13682(.A0(new_n16097_), .A1(new_n11767_), .B0(new_n16118_), .Y(new_n16119_));
  OR3X1    g13683(.A(new_n16085_), .B(new_n12513_), .C(new_n12490_), .Y(new_n16120_));
  OR2X1    g13684(.A(new_n12510_), .B(pi0648), .Y(new_n16121_));
  OR2X1    g13685(.A(pi1159), .B(new_n12517_), .Y(new_n16122_));
  NOR4X1   g13686(.A(new_n16101_), .B(new_n14039_), .C(new_n12473_), .D(pi0619), .Y(new_n16123_));
  NOR4X1   g13687(.A(new_n16101_), .B(new_n14039_), .C(new_n12473_), .D(new_n12509_), .Y(new_n16124_));
  OAI22X1  g13688(.A0(new_n16124_), .A1(new_n16121_), .B0(new_n16123_), .B1(new_n16122_), .Y(new_n16125_));
  AOI21X1  g13689(.A0(new_n16120_), .A1(new_n16116_), .B0(new_n16125_), .Y(new_n16126_));
  OAI21X1  g13690(.A0(new_n2720_), .A1(new_n6851_), .B0(pi0789), .Y(new_n16127_));
  OAI21X1  g13691(.A0(new_n16127_), .A1(new_n16126_), .B0(new_n12709_), .Y(new_n16128_));
  AOI21X1  g13692(.A0(new_n16119_), .A1(new_n16112_), .B0(new_n16128_), .Y(new_n16129_));
  OAI22X1  g13693(.A0(new_n16120_), .A1(new_n12531_), .B0(new_n2720_), .B1(new_n6851_), .Y(new_n16130_));
  NOR4X1   g13694(.A(new_n14040_), .B(new_n14034_), .C(new_n12057_), .D(new_n14767_), .Y(new_n16131_));
  AOI21X1  g13695(.A0(new_n16131_), .A1(new_n12542_), .B0(new_n16068_), .Y(new_n16132_));
  OAI21X1  g13696(.A0(new_n16132_), .A1(pi1158), .B0(pi0641), .Y(new_n16133_));
  AOI21X1  g13697(.A0(new_n16130_), .A1(new_n14049_), .B0(new_n16133_), .Y(new_n16134_));
  AOI21X1  g13698(.A0(new_n16131_), .A1(pi0626), .B0(new_n16068_), .Y(new_n16135_));
  OAI21X1  g13699(.A0(new_n16135_), .A1(new_n12548_), .B0(new_n12543_), .Y(new_n16136_));
  AOI21X1  g13700(.A0(new_n16130_), .A1(new_n14061_), .B0(new_n16136_), .Y(new_n16137_));
  NOR3X1   g13701(.A(new_n16137_), .B(new_n16134_), .C(new_n11765_), .Y(new_n16138_));
  OR2X1    g13702(.A(new_n16138_), .B(new_n14125_), .Y(new_n16139_));
  INVX1    g13703(.A(new_n12708_), .Y(new_n16140_));
  NAND2X1  g13704(.A(new_n16131_), .B(new_n16140_), .Y(new_n16141_));
  OAI21X1  g13705(.A0(new_n16141_), .A1(pi0629), .B0(pi0628), .Y(new_n16142_));
  NOR2X1   g13706(.A(new_n16085_), .B(new_n13489_), .Y(new_n16143_));
  OAI21X1  g13707(.A0(new_n16143_), .A1(new_n12561_), .B0(new_n16142_), .Y(new_n16144_));
  AOI21X1  g13708(.A0(new_n16131_), .A1(new_n16140_), .B0(pi0628), .Y(new_n16145_));
  OAI21X1  g13709(.A0(new_n16145_), .A1(new_n12561_), .B0(pi1156), .Y(new_n16146_));
  AOI21X1  g13710(.A0(new_n16143_), .A1(pi0628), .B0(new_n16146_), .Y(new_n16147_));
  AOI21X1  g13711(.A0(new_n16144_), .A1(new_n12555_), .B0(new_n16147_), .Y(new_n16148_));
  OAI21X1  g13712(.A0(new_n2720_), .A1(new_n6851_), .B0(pi0792), .Y(new_n16149_));
  OAI22X1  g13713(.A0(new_n16149_), .A1(new_n16148_), .B0(new_n16139_), .B1(new_n16129_), .Y(new_n16150_));
  NAND4X1  g13714(.A(new_n16131_), .B(new_n16140_), .C(new_n14327_), .D(new_n12592_), .Y(new_n16151_));
  NOR3X1   g13715(.A(new_n16085_), .B(new_n13508_), .C(new_n13489_), .Y(new_n16152_));
  INVX1    g13716(.A(new_n16152_), .Y(new_n16153_));
  AOI22X1  g13717(.A0(new_n16153_), .A1(pi0630), .B0(new_n16151_), .B1(pi0647), .Y(new_n16154_));
  AOI21X1  g13718(.A0(new_n16153_), .A1(new_n12592_), .B0(new_n12577_), .Y(new_n16155_));
  NAND4X1  g13719(.A(new_n16131_), .B(new_n16140_), .C(new_n14327_), .D(pi0630), .Y(new_n16156_));
  NAND2X1  g13720(.A(new_n16156_), .B(pi1157), .Y(new_n16157_));
  OAI22X1  g13721(.A0(new_n16157_), .A1(new_n16155_), .B0(new_n16154_), .B1(pi1157), .Y(new_n16158_));
  NOR2X1   g13722(.A(new_n16068_), .B(new_n11763_), .Y(new_n16159_));
  AOI22X1  g13723(.A0(new_n16159_), .A1(new_n16158_), .B0(new_n16150_), .B1(new_n14122_), .Y(new_n16160_));
  AOI21X1  g13724(.A0(new_n16152_), .A1(new_n14140_), .B0(new_n16068_), .Y(new_n16161_));
  OAI21X1  g13725(.A0(new_n16161_), .A1(pi0644), .B0(pi0715), .Y(new_n16162_));
  AOI21X1  g13726(.A0(new_n16160_), .A1(pi0644), .B0(new_n16162_), .Y(new_n16163_));
  OR2X1    g13727(.A(new_n12604_), .B(new_n12580_), .Y(new_n16164_));
  NOR3X1   g13728(.A(new_n16164_), .B(new_n16141_), .C(new_n12612_), .Y(new_n16165_));
  OAI21X1  g13729(.A0(new_n2720_), .A1(new_n6851_), .B0(new_n12608_), .Y(new_n16166_));
  OAI21X1  g13730(.A0(new_n16166_), .A1(new_n16165_), .B0(pi1160), .Y(new_n16167_));
  OAI21X1  g13731(.A0(new_n16161_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n16168_));
  AOI21X1  g13732(.A0(new_n16160_), .A1(new_n12612_), .B0(new_n16168_), .Y(new_n16169_));
  NOR3X1   g13733(.A(new_n16164_), .B(new_n16141_), .C(pi0644), .Y(new_n16170_));
  OAI21X1  g13734(.A0(new_n2720_), .A1(new_n6851_), .B0(pi0715), .Y(new_n16171_));
  OAI21X1  g13735(.A0(new_n16171_), .A1(new_n16170_), .B0(new_n11762_), .Y(new_n16172_));
  OAI22X1  g13736(.A0(new_n16172_), .A1(new_n16169_), .B0(new_n16167_), .B1(new_n16163_), .Y(new_n16173_));
  NAND2X1  g13737(.A(new_n16173_), .B(pi0790), .Y(new_n16174_));
  AOI21X1  g13738(.A0(new_n16160_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n16175_));
  AOI22X1  g13739(.A0(new_n16175_), .A1(new_n16174_), .B0(new_n16067_), .B1(new_n16066_), .Y(po0331));
  AOI21X1  g13740(.A0(pi1093), .A1(pi1092), .B0(pi0175), .Y(new_n16177_));
  INVX1    g13741(.A(new_n16177_), .Y(new_n16178_));
  AND2X1   g13742(.A(new_n12056_), .B(pi0766), .Y(new_n16179_));
  OAI21X1  g13743(.A0(new_n16179_), .A1(new_n16177_), .B0(new_n15771_), .Y(new_n16180_));
  AND3X1   g13744(.A(new_n12480_), .B(new_n12056_), .C(pi0766), .Y(new_n16181_));
  OAI21X1  g13745(.A0(new_n16181_), .A1(new_n16180_), .B0(pi1155), .Y(new_n16182_));
  NOR3X1   g13746(.A(new_n16181_), .B(new_n16177_), .C(pi1155), .Y(new_n16183_));
  INVX1    g13747(.A(new_n16183_), .Y(new_n16184_));
  AOI21X1  g13748(.A0(new_n16184_), .A1(new_n16182_), .B0(new_n11768_), .Y(new_n16185_));
  AOI21X1  g13749(.A0(new_n16180_), .A1(new_n11768_), .B0(new_n16185_), .Y(new_n16186_));
  AOI21X1  g13750(.A0(new_n16186_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n16187_));
  AOI21X1  g13751(.A0(new_n16186_), .A1(new_n12655_), .B0(pi1154), .Y(new_n16188_));
  NOR2X1   g13752(.A(new_n16188_), .B(new_n16187_), .Y(new_n16189_));
  MX2X1    g13753(.A(new_n16189_), .B(new_n16186_), .S0(new_n11767_), .Y(new_n16190_));
  NOR2X1   g13754(.A(new_n16190_), .B(pi0789), .Y(new_n16191_));
  AOI21X1  g13755(.A0(new_n16190_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n16192_));
  AOI21X1  g13756(.A0(new_n16190_), .A1(new_n15790_), .B0(pi1159), .Y(new_n16193_));
  OR2X1    g13757(.A(new_n16193_), .B(new_n16192_), .Y(new_n16194_));
  AOI21X1  g13758(.A0(new_n16194_), .A1(pi0789), .B0(new_n16191_), .Y(new_n16195_));
  INVX1    g13759(.A(new_n16195_), .Y(new_n16196_));
  MX2X1    g13760(.A(new_n16196_), .B(new_n16178_), .S0(new_n12708_), .Y(new_n16197_));
  MX2X1    g13761(.A(new_n16197_), .B(new_n16178_), .S0(new_n12580_), .Y(new_n16198_));
  AOI21X1  g13762(.A0(new_n12439_), .A1(pi0700), .B0(new_n16177_), .Y(new_n16199_));
  OR2X1    g13763(.A(new_n16199_), .B(pi0778), .Y(new_n16200_));
  INVX1    g13764(.A(new_n16199_), .Y(new_n16201_));
  AND3X1   g13765(.A(new_n12439_), .B(pi0700), .C(new_n12363_), .Y(new_n16202_));
  INVX1    g13766(.A(new_n16202_), .Y(new_n16203_));
  AOI21X1  g13767(.A0(new_n16203_), .A1(new_n16201_), .B0(new_n12364_), .Y(new_n16204_));
  NOR3X1   g13768(.A(new_n16202_), .B(new_n16177_), .C(pi1153), .Y(new_n16205_));
  OR3X1    g13769(.A(new_n16205_), .B(new_n16204_), .C(new_n11769_), .Y(new_n16206_));
  AND2X1   g13770(.A(new_n16206_), .B(new_n16200_), .Y(new_n16207_));
  NOR4X1   g13771(.A(new_n16207_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n16208_));
  AND3X1   g13772(.A(new_n16208_), .B(new_n12739_), .C(new_n12718_), .Y(new_n16209_));
  INVX1    g13773(.A(new_n16209_), .Y(new_n16210_));
  AOI21X1  g13774(.A0(new_n16177_), .A1(pi0647), .B0(pi1157), .Y(new_n16211_));
  OAI21X1  g13775(.A0(new_n16210_), .A1(pi0647), .B0(new_n16211_), .Y(new_n16212_));
  MX2X1    g13776(.A(new_n16209_), .B(new_n16177_), .S0(new_n12577_), .Y(new_n16213_));
  OAI22X1  g13777(.A0(new_n16213_), .A1(new_n14242_), .B0(new_n16212_), .B1(new_n12592_), .Y(new_n16214_));
  AOI21X1  g13778(.A0(new_n16198_), .A1(new_n14326_), .B0(new_n16214_), .Y(new_n16215_));
  OR2X1    g13779(.A(new_n16215_), .B(new_n11763_), .Y(new_n16216_));
  AND2X1   g13780(.A(new_n12548_), .B(pi0641), .Y(new_n16217_));
  INVX1    g13781(.A(new_n16217_), .Y(new_n16218_));
  AOI21X1  g13782(.A0(new_n16178_), .A1(pi0626), .B0(new_n16218_), .Y(new_n16219_));
  OAI21X1  g13783(.A0(new_n16195_), .A1(pi0626), .B0(new_n16219_), .Y(new_n16220_));
  AND2X1   g13784(.A(pi1158), .B(new_n12543_), .Y(new_n16221_));
  INVX1    g13785(.A(new_n16221_), .Y(new_n16222_));
  AOI21X1  g13786(.A0(new_n16178_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n16223_));
  OAI21X1  g13787(.A0(new_n16195_), .A1(new_n12542_), .B0(new_n16223_), .Y(new_n16224_));
  NAND2X1  g13788(.A(new_n16208_), .B(new_n12637_), .Y(new_n16225_));
  AND3X1   g13789(.A(new_n16225_), .B(new_n16224_), .C(new_n16220_), .Y(new_n16226_));
  NOR2X1   g13790(.A(new_n16226_), .B(new_n11765_), .Y(new_n16227_));
  NOR2X1   g13791(.A(new_n16177_), .B(pi1153), .Y(new_n16228_));
  NOR3X1   g13792(.A(new_n16199_), .B(new_n11991_), .C(new_n12363_), .Y(new_n16229_));
  AOI21X1  g13793(.A0(new_n12056_), .A1(pi0766), .B0(new_n16177_), .Y(new_n16230_));
  INVX1    g13794(.A(new_n16230_), .Y(new_n16231_));
  AOI21X1  g13795(.A0(new_n16201_), .A1(new_n12048_), .B0(new_n16231_), .Y(new_n16232_));
  OAI21X1  g13796(.A0(new_n16232_), .A1(new_n16229_), .B0(new_n16228_), .Y(new_n16233_));
  NOR2X1   g13797(.A(new_n16204_), .B(pi0608), .Y(new_n16234_));
  NOR3X1   g13798(.A(new_n16229_), .B(new_n16231_), .C(new_n12364_), .Y(new_n16235_));
  NOR3X1   g13799(.A(new_n16235_), .B(new_n16205_), .C(new_n12368_), .Y(new_n16236_));
  AOI21X1  g13800(.A0(new_n16234_), .A1(new_n16233_), .B0(new_n16236_), .Y(new_n16237_));
  OR2X1    g13801(.A(new_n16232_), .B(pi0778), .Y(new_n16238_));
  OAI21X1  g13802(.A0(new_n16237_), .A1(new_n11769_), .B0(new_n16238_), .Y(new_n16239_));
  INVX1    g13803(.A(new_n16239_), .Y(new_n16240_));
  AND2X1   g13804(.A(new_n16239_), .B(new_n12462_), .Y(new_n16241_));
  OAI21X1  g13805(.A0(new_n16207_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n16242_));
  OR2X1    g13806(.A(new_n16242_), .B(new_n16241_), .Y(new_n16243_));
  AND3X1   g13807(.A(new_n16243_), .B(new_n16182_), .C(new_n12468_), .Y(new_n16244_));
  OAI21X1  g13808(.A0(new_n16207_), .A1(pi0609), .B0(pi1155), .Y(new_n16245_));
  AOI21X1  g13809(.A0(new_n16239_), .A1(pi0609), .B0(new_n16245_), .Y(new_n16246_));
  NOR3X1   g13810(.A(new_n16246_), .B(new_n16183_), .C(new_n12468_), .Y(new_n16247_));
  NOR2X1   g13811(.A(new_n16247_), .B(new_n16244_), .Y(new_n16248_));
  MX2X1    g13812(.A(new_n16248_), .B(new_n16240_), .S0(new_n11768_), .Y(new_n16249_));
  AOI21X1  g13813(.A0(new_n16206_), .A1(new_n16200_), .B0(new_n12630_), .Y(new_n16250_));
  AOI21X1  g13814(.A0(new_n16250_), .A1(pi0618), .B0(pi1154), .Y(new_n16251_));
  OAI21X1  g13815(.A0(new_n16249_), .A1(pi0618), .B0(new_n16251_), .Y(new_n16252_));
  NOR2X1   g13816(.A(new_n16187_), .B(pi0627), .Y(new_n16253_));
  AOI21X1  g13817(.A0(new_n16250_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n16254_));
  OAI21X1  g13818(.A0(new_n16249_), .A1(new_n12486_), .B0(new_n16254_), .Y(new_n16255_));
  NOR2X1   g13819(.A(new_n16188_), .B(new_n12494_), .Y(new_n16256_));
  AOI22X1  g13820(.A0(new_n16256_), .A1(new_n16255_), .B0(new_n16253_), .B1(new_n16252_), .Y(new_n16257_));
  MX2X1    g13821(.A(new_n16257_), .B(new_n16249_), .S0(new_n11767_), .Y(new_n16258_));
  OR4X1    g13822(.A(new_n16207_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n16259_));
  AND2X1   g13823(.A(new_n16259_), .B(new_n12510_), .Y(new_n16260_));
  OAI21X1  g13824(.A0(new_n16258_), .A1(pi0619), .B0(new_n16260_), .Y(new_n16261_));
  NOR2X1   g13825(.A(new_n16192_), .B(pi0648), .Y(new_n16262_));
  AND2X1   g13826(.A(new_n16262_), .B(new_n16261_), .Y(new_n16263_));
  NOR4X1   g13827(.A(new_n16207_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n16264_));
  NOR2X1   g13828(.A(new_n16264_), .B(new_n12510_), .Y(new_n16265_));
  OAI21X1  g13829(.A0(new_n16258_), .A1(new_n12509_), .B0(new_n16265_), .Y(new_n16266_));
  NOR2X1   g13830(.A(new_n16193_), .B(new_n12517_), .Y(new_n16267_));
  AND2X1   g13831(.A(new_n16267_), .B(new_n16266_), .Y(new_n16268_));
  OR3X1    g13832(.A(new_n16268_), .B(new_n16263_), .C(new_n11766_), .Y(new_n16269_));
  AOI21X1  g13833(.A0(new_n16258_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n16270_));
  AOI21X1  g13834(.A0(new_n16270_), .A1(new_n16269_), .B0(new_n16227_), .Y(new_n16271_));
  INVX1    g13835(.A(new_n16197_), .Y(new_n16272_));
  AND2X1   g13836(.A(new_n16208_), .B(new_n12718_), .Y(new_n16273_));
  AOI22X1  g13837(.A0(new_n16273_), .A1(new_n14426_), .B0(new_n16272_), .B1(new_n12735_), .Y(new_n16274_));
  AOI22X1  g13838(.A0(new_n16273_), .A1(new_n14428_), .B0(new_n16272_), .B1(new_n12733_), .Y(new_n16275_));
  MX2X1    g13839(.A(new_n16275_), .B(new_n16274_), .S0(new_n12561_), .Y(new_n16276_));
  OAI21X1  g13840(.A0(new_n16276_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n16277_));
  INVX1    g13841(.A(new_n16277_), .Y(new_n16278_));
  OAI21X1  g13842(.A0(new_n16271_), .A1(new_n14125_), .B0(new_n16278_), .Y(new_n16279_));
  AND2X1   g13843(.A(new_n16279_), .B(new_n16216_), .Y(new_n16280_));
  OAI21X1  g13844(.A0(new_n16213_), .A1(new_n12578_), .B0(new_n16212_), .Y(new_n16281_));
  MX2X1    g13845(.A(new_n16281_), .B(new_n16210_), .S0(new_n11763_), .Y(new_n16282_));
  OAI21X1  g13846(.A0(new_n16282_), .A1(pi0644), .B0(pi0715), .Y(new_n16283_));
  AOI21X1  g13847(.A0(new_n16280_), .A1(pi0644), .B0(new_n16283_), .Y(new_n16284_));
  OR3X1    g13848(.A(new_n16178_), .B(new_n12603_), .C(new_n11763_), .Y(new_n16285_));
  OAI21X1  g13849(.A0(new_n16198_), .A1(new_n12604_), .B0(new_n16285_), .Y(new_n16286_));
  OAI21X1  g13850(.A0(new_n16178_), .A1(pi0644), .B0(new_n12608_), .Y(new_n16287_));
  AOI21X1  g13851(.A0(new_n16286_), .A1(pi0644), .B0(new_n16287_), .Y(new_n16288_));
  OR2X1    g13852(.A(new_n16288_), .B(new_n11762_), .Y(new_n16289_));
  OAI21X1  g13853(.A0(new_n16282_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n16290_));
  AOI21X1  g13854(.A0(new_n16280_), .A1(new_n12612_), .B0(new_n16290_), .Y(new_n16291_));
  OAI21X1  g13855(.A0(new_n16178_), .A1(new_n12612_), .B0(pi0715), .Y(new_n16292_));
  AOI21X1  g13856(.A0(new_n16286_), .A1(new_n12612_), .B0(new_n16292_), .Y(new_n16293_));
  OR2X1    g13857(.A(new_n16293_), .B(pi1160), .Y(new_n16294_));
  OAI22X1  g13858(.A0(new_n16294_), .A1(new_n16291_), .B0(new_n16289_), .B1(new_n16284_), .Y(new_n16295_));
  NAND2X1  g13859(.A(new_n16295_), .B(pi0790), .Y(new_n16296_));
  AOI21X1  g13860(.A0(new_n16280_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n16297_));
  AOI21X1  g13861(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0175), .Y(new_n16298_));
  INVX1    g13862(.A(new_n16298_), .Y(new_n16299_));
  INVX1    g13863(.A(pi0175), .Y(new_n16300_));
  OAI21X1  g13864(.A0(new_n12826_), .A1(new_n16300_), .B0(new_n2979_), .Y(new_n16301_));
  AOI21X1  g13865(.A0(new_n12825_), .A1(new_n16300_), .B0(new_n16301_), .Y(new_n16302_));
  AOI21X1  g13866(.A0(new_n12771_), .A1(new_n16300_), .B0(new_n12441_), .Y(new_n16303_));
  NOR3X1   g13867(.A(new_n16303_), .B(new_n16302_), .C(new_n14840_), .Y(new_n16304_));
  OR2X1    g13868(.A(pi0700), .B(pi0175), .Y(new_n16305_));
  OAI21X1  g13869(.A0(new_n16305_), .A1(new_n12447_), .B0(new_n3103_), .Y(new_n16306_));
  OAI22X1  g13870(.A0(new_n16306_), .A1(new_n16304_), .B0(new_n3103_), .B1(new_n16300_), .Y(new_n16307_));
  AND2X1   g13871(.A(new_n16307_), .B(new_n11769_), .Y(new_n16308_));
  AOI21X1  g13872(.A0(new_n16298_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n16309_));
  OAI21X1  g13873(.A0(new_n16307_), .A1(new_n12363_), .B0(new_n16309_), .Y(new_n16310_));
  AOI21X1  g13874(.A0(new_n16298_), .A1(pi0625), .B0(pi1153), .Y(new_n16311_));
  OAI21X1  g13875(.A0(new_n16307_), .A1(pi0625), .B0(new_n16311_), .Y(new_n16312_));
  AOI21X1  g13876(.A0(new_n16312_), .A1(new_n16310_), .B0(new_n11769_), .Y(new_n16313_));
  NOR2X1   g13877(.A(new_n16313_), .B(new_n16308_), .Y(new_n16314_));
  MX2X1    g13878(.A(new_n16314_), .B(new_n16298_), .S0(new_n12490_), .Y(new_n16315_));
  AND2X1   g13879(.A(new_n16298_), .B(new_n12513_), .Y(new_n16316_));
  AOI21X1  g13880(.A0(new_n16315_), .A1(new_n14053_), .B0(new_n16316_), .Y(new_n16317_));
  MX2X1    g13881(.A(new_n16317_), .B(new_n16299_), .S0(new_n12531_), .Y(new_n16318_));
  MX2X1    g13882(.A(new_n16318_), .B(new_n16299_), .S0(new_n12563_), .Y(new_n16319_));
  MX2X1    g13883(.A(new_n16319_), .B(new_n16299_), .S0(pi0628), .Y(new_n16320_));
  MX2X1    g13884(.A(new_n16319_), .B(new_n16299_), .S0(new_n12554_), .Y(new_n16321_));
  MX2X1    g13885(.A(new_n16321_), .B(new_n16320_), .S0(new_n12555_), .Y(new_n16322_));
  MX2X1    g13886(.A(new_n16322_), .B(new_n16319_), .S0(new_n11764_), .Y(new_n16323_));
  MX2X1    g13887(.A(new_n16323_), .B(new_n16299_), .S0(pi0647), .Y(new_n16324_));
  MX2X1    g13888(.A(new_n16323_), .B(new_n16299_), .S0(new_n12577_), .Y(new_n16325_));
  MX2X1    g13889(.A(new_n16325_), .B(new_n16324_), .S0(new_n12578_), .Y(new_n16326_));
  MX2X1    g13890(.A(new_n16326_), .B(new_n16323_), .S0(new_n11763_), .Y(new_n16327_));
  OAI21X1  g13891(.A0(new_n16327_), .A1(pi0644), .B0(pi0715), .Y(new_n16328_));
  AOI22X1  g13892(.A0(new_n12073_), .A1(pi0175), .B0(new_n12444_), .B1(new_n14844_), .Y(new_n16329_));
  OR3X1    g13893(.A(new_n12776_), .B(new_n14844_), .C(pi0175), .Y(new_n16330_));
  OAI21X1  g13894(.A0(new_n12045_), .A1(pi0039), .B0(pi0766), .Y(new_n16331_));
  AOI21X1  g13895(.A0(new_n16331_), .A1(pi0175), .B0(new_n14845_), .Y(new_n16332_));
  AND2X1   g13896(.A(new_n16332_), .B(new_n16330_), .Y(new_n16333_));
  OAI21X1  g13897(.A0(new_n16329_), .A1(new_n2939_), .B0(new_n16333_), .Y(new_n16334_));
  OAI21X1  g13898(.A0(new_n12077_), .A1(pi0175), .B0(pi0038), .Y(new_n16335_));
  AOI21X1  g13899(.A0(new_n12079_), .A1(pi0766), .B0(new_n16335_), .Y(new_n16336_));
  AOI21X1  g13900(.A0(new_n16334_), .A1(new_n2979_), .B0(new_n16336_), .Y(new_n16337_));
  MX2X1    g13901(.A(new_n16337_), .B(new_n16300_), .S0(new_n11770_), .Y(new_n16338_));
  MX2X1    g13902(.A(new_n16338_), .B(new_n16298_), .S0(new_n12473_), .Y(new_n16339_));
  NOR2X1   g13903(.A(new_n16338_), .B(new_n12473_), .Y(new_n16340_));
  AOI22X1  g13904(.A0(new_n16340_), .A1(pi0609), .B0(new_n16299_), .B1(new_n12472_), .Y(new_n16341_));
  AOI22X1  g13905(.A0(new_n16340_), .A1(new_n12462_), .B0(new_n16299_), .B1(new_n12481_), .Y(new_n16342_));
  MX2X1    g13906(.A(new_n16342_), .B(new_n16341_), .S0(pi1155), .Y(new_n16343_));
  MX2X1    g13907(.A(new_n16343_), .B(new_n16339_), .S0(new_n11768_), .Y(new_n16344_));
  OAI21X1  g13908(.A0(new_n16299_), .A1(pi0618), .B0(pi1154), .Y(new_n16345_));
  AOI21X1  g13909(.A0(new_n16344_), .A1(pi0618), .B0(new_n16345_), .Y(new_n16346_));
  OAI21X1  g13910(.A0(new_n16299_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n16347_));
  AOI21X1  g13911(.A0(new_n16344_), .A1(new_n12486_), .B0(new_n16347_), .Y(new_n16348_));
  NOR2X1   g13912(.A(new_n16348_), .B(new_n16346_), .Y(new_n16349_));
  MX2X1    g13913(.A(new_n16349_), .B(new_n16344_), .S0(new_n11767_), .Y(new_n16350_));
  OAI21X1  g13914(.A0(new_n16299_), .A1(pi0619), .B0(pi1159), .Y(new_n16351_));
  AOI21X1  g13915(.A0(new_n16350_), .A1(pi0619), .B0(new_n16351_), .Y(new_n16352_));
  OAI21X1  g13916(.A0(new_n16299_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n16353_));
  AOI21X1  g13917(.A0(new_n16350_), .A1(new_n12509_), .B0(new_n16353_), .Y(new_n16354_));
  NOR2X1   g13918(.A(new_n16354_), .B(new_n16352_), .Y(new_n16355_));
  MX2X1    g13919(.A(new_n16355_), .B(new_n16350_), .S0(new_n11766_), .Y(new_n16356_));
  AND2X1   g13920(.A(new_n16298_), .B(new_n12708_), .Y(new_n16357_));
  AOI21X1  g13921(.A0(new_n16356_), .A1(new_n16140_), .B0(new_n16357_), .Y(new_n16358_));
  MX2X1    g13922(.A(new_n16358_), .B(new_n16299_), .S0(new_n12580_), .Y(new_n16359_));
  MX2X1    g13923(.A(new_n16359_), .B(new_n16299_), .S0(new_n12604_), .Y(new_n16360_));
  AOI21X1  g13924(.A0(new_n16298_), .A1(new_n12612_), .B0(pi0715), .Y(new_n16361_));
  OAI21X1  g13925(.A0(new_n16360_), .A1(new_n12612_), .B0(new_n16361_), .Y(new_n16362_));
  NAND3X1  g13926(.A(new_n16362_), .B(new_n16328_), .C(pi1160), .Y(new_n16363_));
  OAI21X1  g13927(.A0(new_n16327_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n16364_));
  AOI21X1  g13928(.A0(new_n16298_), .A1(pi0644), .B0(new_n12608_), .Y(new_n16365_));
  OAI21X1  g13929(.A0(new_n16360_), .A1(pi0644), .B0(new_n16365_), .Y(new_n16366_));
  NAND3X1  g13930(.A(new_n16366_), .B(new_n16364_), .C(new_n11762_), .Y(new_n16367_));
  AND2X1   g13931(.A(new_n16367_), .B(new_n16363_), .Y(new_n16368_));
  NAND3X1  g13932(.A(new_n16366_), .B(new_n11762_), .C(new_n12612_), .Y(new_n16369_));
  NAND3X1  g13933(.A(new_n16362_), .B(pi1160), .C(pi0644), .Y(new_n16370_));
  AND3X1   g13934(.A(new_n16370_), .B(new_n16369_), .C(pi0790), .Y(new_n16371_));
  NAND2X1  g13935(.A(new_n16358_), .B(new_n14249_), .Y(new_n16372_));
  AND2X1   g13936(.A(pi1156), .B(new_n12561_), .Y(new_n16373_));
  AND2X1   g13937(.A(new_n12555_), .B(pi0629), .Y(new_n16374_));
  AOI22X1  g13938(.A0(new_n16321_), .A1(new_n16373_), .B0(new_n16320_), .B1(new_n16374_), .Y(new_n16375_));
  AOI21X1  g13939(.A0(new_n16375_), .A1(new_n16372_), .B0(new_n11764_), .Y(new_n16376_));
  AND2X1   g13940(.A(new_n16337_), .B(new_n14840_), .Y(new_n16377_));
  INVX1    g13941(.A(new_n16377_), .Y(new_n16378_));
  NAND2X1  g13942(.A(new_n12145_), .B(new_n12116_), .Y(new_n16379_));
  MX2X1    g13943(.A(new_n12154_), .B(new_n16379_), .S0(new_n2933_), .Y(new_n16380_));
  INVX1    g13944(.A(new_n12213_), .Y(new_n16381_));
  AOI21X1  g13945(.A0(new_n16381_), .A1(pi0175), .B0(pi0766), .Y(new_n16382_));
  OAI21X1  g13946(.A0(new_n16380_), .A1(pi0175), .B0(new_n16382_), .Y(new_n16383_));
  AOI21X1  g13947(.A0(new_n12788_), .A1(new_n16300_), .B0(new_n14844_), .Y(new_n16384_));
  OAI21X1  g13948(.A0(new_n12787_), .A1(new_n16300_), .B0(new_n16384_), .Y(new_n16385_));
  AND2X1   g13949(.A(new_n16385_), .B(pi0039), .Y(new_n16386_));
  AND2X1   g13950(.A(new_n16386_), .B(new_n16383_), .Y(new_n16387_));
  AOI21X1  g13951(.A0(new_n12795_), .A1(pi0175), .B0(pi0766), .Y(new_n16388_));
  OAI21X1  g13952(.A0(new_n12792_), .A1(pi0175), .B0(new_n16388_), .Y(new_n16389_));
  NOR2X1   g13953(.A(new_n12798_), .B(pi0175), .Y(new_n16390_));
  INVX1    g13954(.A(new_n16390_), .Y(new_n16391_));
  AOI21X1  g13955(.A0(new_n12800_), .A1(pi0175), .B0(new_n14844_), .Y(new_n16392_));
  AOI21X1  g13956(.A0(new_n16392_), .A1(new_n16391_), .B0(pi0039), .Y(new_n16393_));
  AOI21X1  g13957(.A0(new_n16393_), .A1(new_n16389_), .B0(pi0038), .Y(new_n16394_));
  INVX1    g13958(.A(new_n16394_), .Y(new_n16395_));
  NOR4X1   g13959(.A(new_n12085_), .B(new_n2985_), .C(new_n2725_), .D(new_n2536_), .Y(new_n16396_));
  AOI21X1  g13960(.A0(new_n16396_), .A1(new_n14844_), .B0(new_n12276_), .Y(new_n16397_));
  OAI21X1  g13961(.A0(new_n16397_), .A1(pi0039), .B0(new_n16300_), .Y(new_n16398_));
  INVX1    g13962(.A(new_n5782_), .Y(new_n16399_));
  OAI21X1  g13963(.A0(new_n16179_), .A1(new_n13443_), .B0(pi0175), .Y(new_n16400_));
  OAI21X1  g13964(.A0(new_n16400_), .A1(new_n16399_), .B0(pi0038), .Y(new_n16401_));
  INVX1    g13965(.A(new_n16401_), .Y(new_n16402_));
  AOI21X1  g13966(.A0(new_n16402_), .A1(new_n16398_), .B0(new_n14840_), .Y(new_n16403_));
  OAI21X1  g13967(.A0(new_n16395_), .A1(new_n16387_), .B0(new_n16403_), .Y(new_n16404_));
  AND2X1   g13968(.A(new_n16404_), .B(new_n3103_), .Y(new_n16405_));
  AOI22X1  g13969(.A0(new_n16405_), .A1(new_n16378_), .B0(new_n11770_), .B1(pi0175), .Y(new_n16406_));
  INVX1    g13970(.A(new_n16406_), .Y(new_n16407_));
  AOI21X1  g13971(.A0(new_n16338_), .A1(pi0625), .B0(pi1153), .Y(new_n16408_));
  OAI21X1  g13972(.A0(new_n16407_), .A1(pi0625), .B0(new_n16408_), .Y(new_n16409_));
  AND2X1   g13973(.A(new_n16310_), .B(new_n12368_), .Y(new_n16410_));
  AOI21X1  g13974(.A0(new_n16338_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n16411_));
  OAI21X1  g13975(.A0(new_n16407_), .A1(new_n12363_), .B0(new_n16411_), .Y(new_n16412_));
  AND2X1   g13976(.A(new_n16312_), .B(pi0608), .Y(new_n16413_));
  AOI22X1  g13977(.A0(new_n16413_), .A1(new_n16412_), .B0(new_n16410_), .B1(new_n16409_), .Y(new_n16414_));
  MX2X1    g13978(.A(new_n16414_), .B(new_n16407_), .S0(new_n11769_), .Y(new_n16415_));
  AOI21X1  g13979(.A0(new_n16314_), .A1(pi0609), .B0(pi1155), .Y(new_n16416_));
  OAI21X1  g13980(.A0(new_n16415_), .A1(pi0609), .B0(new_n16416_), .Y(new_n16417_));
  OAI21X1  g13981(.A0(new_n16341_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n16418_));
  INVX1    g13982(.A(new_n16418_), .Y(new_n16419_));
  AOI21X1  g13983(.A0(new_n16314_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n16420_));
  OAI21X1  g13984(.A0(new_n16415_), .A1(new_n12462_), .B0(new_n16420_), .Y(new_n16421_));
  OAI21X1  g13985(.A0(new_n16342_), .A1(pi1155), .B0(pi0660), .Y(new_n16422_));
  INVX1    g13986(.A(new_n16422_), .Y(new_n16423_));
  AOI22X1  g13987(.A0(new_n16423_), .A1(new_n16421_), .B0(new_n16419_), .B1(new_n16417_), .Y(new_n16424_));
  MX2X1    g13988(.A(new_n16424_), .B(new_n16415_), .S0(new_n11768_), .Y(new_n16425_));
  AOI21X1  g13989(.A0(new_n16315_), .A1(pi0618), .B0(pi1154), .Y(new_n16426_));
  OAI21X1  g13990(.A0(new_n16425_), .A1(pi0618), .B0(new_n16426_), .Y(new_n16427_));
  NOR2X1   g13991(.A(new_n16346_), .B(pi0627), .Y(new_n16428_));
  AOI21X1  g13992(.A0(new_n16315_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n16429_));
  OAI21X1  g13993(.A0(new_n16425_), .A1(new_n12486_), .B0(new_n16429_), .Y(new_n16430_));
  NOR2X1   g13994(.A(new_n16348_), .B(new_n12494_), .Y(new_n16431_));
  AOI22X1  g13995(.A0(new_n16431_), .A1(new_n16430_), .B0(new_n16428_), .B1(new_n16427_), .Y(new_n16432_));
  MX2X1    g13996(.A(new_n16432_), .B(new_n16425_), .S0(new_n11767_), .Y(new_n16433_));
  INVX1    g13997(.A(new_n16433_), .Y(new_n16434_));
  OAI21X1  g13998(.A0(new_n16317_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n16435_));
  AOI21X1  g13999(.A0(new_n16434_), .A1(new_n12509_), .B0(new_n16435_), .Y(new_n16436_));
  NOR3X1   g14000(.A(new_n16436_), .B(new_n16352_), .C(pi0648), .Y(new_n16437_));
  OAI21X1  g14001(.A0(new_n16317_), .A1(pi0619), .B0(pi1159), .Y(new_n16438_));
  AOI21X1  g14002(.A0(new_n16434_), .A1(pi0619), .B0(new_n16438_), .Y(new_n16439_));
  OR2X1    g14003(.A(new_n16354_), .B(new_n12517_), .Y(new_n16440_));
  OAI21X1  g14004(.A0(new_n16440_), .A1(new_n16439_), .B0(pi0789), .Y(new_n16441_));
  AOI21X1  g14005(.A0(new_n16433_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n16442_));
  OAI21X1  g14006(.A0(new_n16441_), .A1(new_n16437_), .B0(new_n16442_), .Y(new_n16443_));
  AOI21X1  g14007(.A0(new_n16299_), .A1(pi0626), .B0(new_n16218_), .Y(new_n16444_));
  OAI21X1  g14008(.A0(new_n16356_), .A1(pi0626), .B0(new_n16444_), .Y(new_n16445_));
  AOI21X1  g14009(.A0(new_n16299_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n16446_));
  OAI21X1  g14010(.A0(new_n16356_), .A1(new_n12542_), .B0(new_n16446_), .Y(new_n16447_));
  OR2X1    g14011(.A(new_n16318_), .B(new_n13439_), .Y(new_n16448_));
  NAND3X1  g14012(.A(new_n16448_), .B(new_n16447_), .C(new_n16445_), .Y(new_n16449_));
  AOI21X1  g14013(.A0(new_n16449_), .A1(pi0788), .B0(new_n14125_), .Y(new_n16450_));
  AOI21X1  g14014(.A0(new_n16450_), .A1(new_n16443_), .B0(new_n16376_), .Y(new_n16451_));
  AND2X1   g14015(.A(new_n16359_), .B(new_n14326_), .Y(new_n16452_));
  AND2X1   g14016(.A(new_n16325_), .B(new_n14241_), .Y(new_n16453_));
  AND2X1   g14017(.A(new_n16324_), .B(new_n14243_), .Y(new_n16454_));
  OR2X1    g14018(.A(new_n16454_), .B(new_n16453_), .Y(new_n16455_));
  OAI21X1  g14019(.A0(new_n16455_), .A1(new_n16452_), .B0(pi0787), .Y(new_n16456_));
  OAI21X1  g14020(.A0(new_n16451_), .A1(new_n14121_), .B0(new_n16456_), .Y(new_n16457_));
  OAI22X1  g14021(.A0(new_n16457_), .A1(new_n16371_), .B0(new_n16368_), .B1(new_n12766_), .Y(new_n16458_));
  OAI21X1  g14022(.A0(new_n6489_), .A1(pi0175), .B0(new_n12767_), .Y(new_n16459_));
  AOI21X1  g14023(.A0(new_n16458_), .A1(new_n6489_), .B0(new_n16459_), .Y(new_n16460_));
  AOI21X1  g14024(.A0(new_n16297_), .A1(new_n16296_), .B0(new_n16460_), .Y(po0332));
  AOI21X1  g14025(.A0(pi1093), .A1(pi1092), .B0(pi0176), .Y(new_n16462_));
  INVX1    g14026(.A(new_n16462_), .Y(new_n16463_));
  AOI21X1  g14027(.A0(new_n12056_), .A1(new_n14897_), .B0(new_n16462_), .Y(new_n16464_));
  AOI21X1  g14028(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n16464_), .Y(new_n16465_));
  INVX1    g14029(.A(new_n16464_), .Y(new_n16466_));
  AOI21X1  g14030(.A0(new_n16466_), .A1(new_n14331_), .B0(new_n12463_), .Y(new_n16467_));
  AOI21X1  g14031(.A0(new_n16465_), .A1(new_n12646_), .B0(pi1155), .Y(new_n16468_));
  OAI21X1  g14032(.A0(new_n16468_), .A1(new_n16467_), .B0(pi0785), .Y(new_n16469_));
  OAI21X1  g14033(.A0(new_n16465_), .A1(pi0785), .B0(new_n16469_), .Y(new_n16470_));
  INVX1    g14034(.A(new_n16470_), .Y(new_n16471_));
  AOI21X1  g14035(.A0(new_n16471_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n16472_));
  AOI21X1  g14036(.A0(new_n16471_), .A1(new_n12655_), .B0(pi1154), .Y(new_n16473_));
  NOR2X1   g14037(.A(new_n16473_), .B(new_n16472_), .Y(new_n16474_));
  MX2X1    g14038(.A(new_n16474_), .B(new_n16471_), .S0(new_n11767_), .Y(new_n16475_));
  OR2X1    g14039(.A(new_n16475_), .B(pi0789), .Y(new_n16476_));
  OAI21X1  g14040(.A0(new_n16463_), .A1(pi0619), .B0(pi1159), .Y(new_n16477_));
  AOI21X1  g14041(.A0(new_n16475_), .A1(pi0619), .B0(new_n16477_), .Y(new_n16478_));
  OAI21X1  g14042(.A0(new_n16463_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n16479_));
  AOI21X1  g14043(.A0(new_n16475_), .A1(new_n12509_), .B0(new_n16479_), .Y(new_n16480_));
  OAI21X1  g14044(.A0(new_n16480_), .A1(new_n16478_), .B0(pi0789), .Y(new_n16481_));
  AND2X1   g14045(.A(new_n16481_), .B(new_n16476_), .Y(new_n16482_));
  INVX1    g14046(.A(new_n16482_), .Y(new_n16483_));
  MX2X1    g14047(.A(new_n16483_), .B(new_n16463_), .S0(new_n12708_), .Y(new_n16484_));
  MX2X1    g14048(.A(new_n16484_), .B(new_n16463_), .S0(new_n12580_), .Y(new_n16485_));
  AOI21X1  g14049(.A0(new_n12439_), .A1(new_n14896_), .B0(new_n16462_), .Y(new_n16486_));
  AND3X1   g14050(.A(new_n12439_), .B(new_n14896_), .C(new_n12363_), .Y(new_n16487_));
  NOR2X1   g14051(.A(new_n16487_), .B(new_n16486_), .Y(new_n16488_));
  OR3X1    g14052(.A(new_n16487_), .B(new_n16462_), .C(pi1153), .Y(new_n16489_));
  OAI21X1  g14053(.A0(new_n16488_), .A1(new_n12364_), .B0(new_n16489_), .Y(new_n16490_));
  MX2X1    g14054(.A(new_n16490_), .B(new_n16486_), .S0(new_n11769_), .Y(new_n16491_));
  NOR4X1   g14055(.A(new_n16491_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n16492_));
  NAND4X1  g14056(.A(new_n16492_), .B(new_n12739_), .C(new_n12718_), .D(new_n12577_), .Y(new_n16493_));
  AOI21X1  g14057(.A0(new_n16462_), .A1(pi0647), .B0(pi1157), .Y(new_n16494_));
  NAND2X1  g14058(.A(new_n16494_), .B(new_n16493_), .Y(new_n16495_));
  INVX1    g14059(.A(new_n16495_), .Y(new_n16496_));
  AND3X1   g14060(.A(new_n16492_), .B(new_n12739_), .C(new_n12718_), .Y(new_n16497_));
  MX2X1    g14061(.A(new_n16497_), .B(new_n16462_), .S0(new_n12577_), .Y(new_n16498_));
  INVX1    g14062(.A(new_n16498_), .Y(new_n16499_));
  AOI22X1  g14063(.A0(new_n16499_), .A1(new_n14241_), .B0(new_n16496_), .B1(pi0630), .Y(new_n16500_));
  INVX1    g14064(.A(new_n16500_), .Y(new_n16501_));
  AOI21X1  g14065(.A0(new_n16485_), .A1(new_n14326_), .B0(new_n16501_), .Y(new_n16502_));
  AOI21X1  g14066(.A0(new_n16463_), .A1(pi0626), .B0(new_n16218_), .Y(new_n16503_));
  OAI21X1  g14067(.A0(new_n16482_), .A1(pi0626), .B0(new_n16503_), .Y(new_n16504_));
  AOI21X1  g14068(.A0(new_n16463_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n16505_));
  OAI21X1  g14069(.A0(new_n16482_), .A1(new_n12542_), .B0(new_n16505_), .Y(new_n16506_));
  NAND2X1  g14070(.A(new_n16492_), .B(new_n12637_), .Y(new_n16507_));
  AND3X1   g14071(.A(new_n16507_), .B(new_n16506_), .C(new_n16504_), .Y(new_n16508_));
  NOR2X1   g14072(.A(new_n16508_), .B(new_n11765_), .Y(new_n16509_));
  INVX1    g14073(.A(new_n16509_), .Y(new_n16510_));
  NOR2X1   g14074(.A(new_n16462_), .B(pi1153), .Y(new_n16511_));
  NOR2X1   g14075(.A(new_n16486_), .B(new_n11991_), .Y(new_n16512_));
  MX2X1    g14076(.A(new_n16464_), .B(pi0625), .S0(new_n16512_), .Y(new_n16513_));
  OAI21X1  g14077(.A0(new_n16488_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n16514_));
  AOI21X1  g14078(.A0(new_n16513_), .A1(new_n16511_), .B0(new_n16514_), .Y(new_n16515_));
  NOR3X1   g14079(.A(new_n16486_), .B(new_n11991_), .C(new_n12363_), .Y(new_n16516_));
  OR3X1    g14080(.A(new_n16516_), .B(new_n16466_), .C(new_n12364_), .Y(new_n16517_));
  AND3X1   g14081(.A(new_n16517_), .B(new_n16489_), .C(pi0608), .Y(new_n16518_));
  OAI21X1  g14082(.A0(new_n16518_), .A1(new_n16515_), .B0(pi0778), .Y(new_n16519_));
  OAI21X1  g14083(.A0(new_n16512_), .A1(new_n16466_), .B0(new_n11769_), .Y(new_n16520_));
  AND2X1   g14084(.A(new_n16520_), .B(new_n16519_), .Y(new_n16521_));
  NAND2X1  g14085(.A(new_n16520_), .B(new_n16519_), .Y(new_n16522_));
  OAI21X1  g14086(.A0(new_n16491_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n16523_));
  AOI21X1  g14087(.A0(new_n16522_), .A1(new_n12462_), .B0(new_n16523_), .Y(new_n16524_));
  NOR3X1   g14088(.A(new_n16524_), .B(new_n16467_), .C(pi0660), .Y(new_n16525_));
  OAI21X1  g14089(.A0(new_n16491_), .A1(pi0609), .B0(pi1155), .Y(new_n16526_));
  AOI21X1  g14090(.A0(new_n16522_), .A1(pi0609), .B0(new_n16526_), .Y(new_n16527_));
  NOR3X1   g14091(.A(new_n16527_), .B(new_n16468_), .C(new_n12468_), .Y(new_n16528_));
  NOR2X1   g14092(.A(new_n16528_), .B(new_n16525_), .Y(new_n16529_));
  MX2X1    g14093(.A(new_n16529_), .B(new_n16521_), .S0(new_n11768_), .Y(new_n16530_));
  OR3X1    g14094(.A(new_n16491_), .B(new_n12630_), .C(new_n12486_), .Y(new_n16531_));
  AND2X1   g14095(.A(new_n16531_), .B(new_n12487_), .Y(new_n16532_));
  OAI21X1  g14096(.A0(new_n16530_), .A1(pi0618), .B0(new_n16532_), .Y(new_n16533_));
  NOR2X1   g14097(.A(new_n16472_), .B(pi0627), .Y(new_n16534_));
  NOR3X1   g14098(.A(new_n16491_), .B(new_n12630_), .C(pi0618), .Y(new_n16535_));
  NOR2X1   g14099(.A(new_n16535_), .B(new_n12487_), .Y(new_n16536_));
  OAI21X1  g14100(.A0(new_n16530_), .A1(new_n12486_), .B0(new_n16536_), .Y(new_n16537_));
  NOR2X1   g14101(.A(new_n16473_), .B(new_n12494_), .Y(new_n16538_));
  AOI22X1  g14102(.A0(new_n16538_), .A1(new_n16537_), .B0(new_n16534_), .B1(new_n16533_), .Y(new_n16539_));
  MX2X1    g14103(.A(new_n16539_), .B(new_n16530_), .S0(new_n11767_), .Y(new_n16540_));
  OR4X1    g14104(.A(new_n16491_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n16541_));
  AND2X1   g14105(.A(new_n16541_), .B(new_n12510_), .Y(new_n16542_));
  OAI21X1  g14106(.A0(new_n16540_), .A1(pi0619), .B0(new_n16542_), .Y(new_n16543_));
  NOR2X1   g14107(.A(new_n16478_), .B(pi0648), .Y(new_n16544_));
  AND2X1   g14108(.A(new_n16544_), .B(new_n16543_), .Y(new_n16545_));
  NOR4X1   g14109(.A(new_n16491_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n16546_));
  NOR2X1   g14110(.A(new_n16546_), .B(new_n12510_), .Y(new_n16547_));
  OAI21X1  g14111(.A0(new_n16540_), .A1(new_n12509_), .B0(new_n16547_), .Y(new_n16548_));
  NOR2X1   g14112(.A(new_n16480_), .B(new_n12517_), .Y(new_n16549_));
  AOI21X1  g14113(.A0(new_n16549_), .A1(new_n16548_), .B0(new_n11766_), .Y(new_n16550_));
  INVX1    g14114(.A(new_n16550_), .Y(new_n16551_));
  AOI21X1  g14115(.A0(new_n16540_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n16552_));
  OAI21X1  g14116(.A0(new_n16551_), .A1(new_n16545_), .B0(new_n16552_), .Y(new_n16553_));
  AOI21X1  g14117(.A0(new_n16553_), .A1(new_n16510_), .B0(new_n14125_), .Y(new_n16554_));
  INVX1    g14118(.A(new_n16484_), .Y(new_n16555_));
  AND2X1   g14119(.A(new_n16492_), .B(new_n12718_), .Y(new_n16556_));
  AOI22X1  g14120(.A0(new_n16556_), .A1(new_n14426_), .B0(new_n16555_), .B1(new_n12735_), .Y(new_n16557_));
  AOI22X1  g14121(.A0(new_n16556_), .A1(new_n14428_), .B0(new_n16555_), .B1(new_n12733_), .Y(new_n16558_));
  MX2X1    g14122(.A(new_n16558_), .B(new_n16557_), .S0(new_n12561_), .Y(new_n16559_));
  OAI21X1  g14123(.A0(new_n16559_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n16560_));
  OAI22X1  g14124(.A0(new_n16560_), .A1(new_n16554_), .B0(new_n16502_), .B1(new_n11763_), .Y(new_n16561_));
  AOI21X1  g14125(.A0(new_n16499_), .A1(pi1157), .B0(new_n16496_), .Y(new_n16562_));
  MX2X1    g14126(.A(new_n16562_), .B(new_n16497_), .S0(new_n11763_), .Y(new_n16563_));
  AOI21X1  g14127(.A0(new_n16563_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n16564_));
  OAI21X1  g14128(.A0(new_n16561_), .A1(new_n12612_), .B0(new_n16564_), .Y(new_n16565_));
  MX2X1    g14129(.A(new_n16485_), .B(new_n16463_), .S0(new_n12604_), .Y(new_n16566_));
  AOI21X1  g14130(.A0(new_n16462_), .A1(new_n12612_), .B0(pi0715), .Y(new_n16567_));
  OAI21X1  g14131(.A0(new_n16566_), .A1(new_n12612_), .B0(new_n16567_), .Y(new_n16568_));
  AND2X1   g14132(.A(new_n16568_), .B(pi1160), .Y(new_n16569_));
  AOI21X1  g14133(.A0(new_n16563_), .A1(pi0644), .B0(pi0715), .Y(new_n16570_));
  OAI21X1  g14134(.A0(new_n16561_), .A1(pi0644), .B0(new_n16570_), .Y(new_n16571_));
  AOI21X1  g14135(.A0(new_n16462_), .A1(pi0644), .B0(new_n12608_), .Y(new_n16572_));
  OAI21X1  g14136(.A0(new_n16566_), .A1(pi0644), .B0(new_n16572_), .Y(new_n16573_));
  AND2X1   g14137(.A(new_n16573_), .B(new_n11762_), .Y(new_n16574_));
  AOI22X1  g14138(.A0(new_n16574_), .A1(new_n16571_), .B0(new_n16569_), .B1(new_n16565_), .Y(new_n16575_));
  OR2X1    g14139(.A(new_n16561_), .B(pi0790), .Y(new_n16576_));
  AND2X1   g14140(.A(new_n16576_), .B(pi0832), .Y(new_n16577_));
  OAI21X1  g14141(.A0(new_n16575_), .A1(new_n12766_), .B0(new_n16577_), .Y(new_n16578_));
  AOI21X1  g14142(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0176), .Y(new_n16579_));
  INVX1    g14143(.A(new_n16579_), .Y(new_n16580_));
  NOR2X1   g14144(.A(new_n13870_), .B(pi0038), .Y(new_n16581_));
  OR3X1    g14145(.A(new_n16581_), .B(new_n12440_), .C(new_n11770_), .Y(new_n16582_));
  OAI21X1  g14146(.A0(new_n13868_), .A1(pi0038), .B0(new_n13874_), .Y(new_n16583_));
  INVX1    g14147(.A(new_n16583_), .Y(new_n16584_));
  AOI21X1  g14148(.A0(new_n16584_), .A1(new_n6832_), .B0(pi0704), .Y(new_n16585_));
  INVX1    g14149(.A(new_n16585_), .Y(new_n16586_));
  AND2X1   g14150(.A(new_n12832_), .B(new_n6832_), .Y(new_n16587_));
  AOI21X1  g14151(.A0(new_n16587_), .A1(pi0704), .B0(new_n11770_), .Y(new_n16588_));
  AOI22X1  g14152(.A0(new_n16588_), .A1(new_n16586_), .B0(new_n16582_), .B1(pi0176), .Y(new_n16589_));
  OAI21X1  g14153(.A0(new_n16580_), .A1(pi0625), .B0(pi1153), .Y(new_n16590_));
  AOI21X1  g14154(.A0(new_n16589_), .A1(pi0625), .B0(new_n16590_), .Y(new_n16591_));
  OAI21X1  g14155(.A0(new_n16580_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n16592_));
  AOI21X1  g14156(.A0(new_n16589_), .A1(new_n12363_), .B0(new_n16592_), .Y(new_n16593_));
  NOR2X1   g14157(.A(new_n16593_), .B(new_n16591_), .Y(new_n16594_));
  MX2X1    g14158(.A(new_n16594_), .B(new_n16589_), .S0(new_n11769_), .Y(new_n16595_));
  MX2X1    g14159(.A(new_n16595_), .B(new_n16579_), .S0(new_n12490_), .Y(new_n16596_));
  AND2X1   g14160(.A(new_n16579_), .B(new_n12513_), .Y(new_n16597_));
  AOI21X1  g14161(.A0(new_n16596_), .A1(new_n14053_), .B0(new_n16597_), .Y(new_n16598_));
  MX2X1    g14162(.A(new_n16598_), .B(new_n16580_), .S0(new_n12531_), .Y(new_n16599_));
  MX2X1    g14163(.A(new_n16599_), .B(new_n16580_), .S0(new_n12563_), .Y(new_n16600_));
  MX2X1    g14164(.A(new_n16600_), .B(new_n16580_), .S0(pi0628), .Y(new_n16601_));
  MX2X1    g14165(.A(new_n16600_), .B(new_n16580_), .S0(new_n12554_), .Y(new_n16602_));
  MX2X1    g14166(.A(new_n16602_), .B(new_n16601_), .S0(new_n12555_), .Y(new_n16603_));
  MX2X1    g14167(.A(new_n16603_), .B(new_n16600_), .S0(new_n11764_), .Y(new_n16604_));
  MX2X1    g14168(.A(new_n16604_), .B(new_n16580_), .S0(pi0647), .Y(new_n16605_));
  MX2X1    g14169(.A(new_n16604_), .B(new_n16580_), .S0(new_n12577_), .Y(new_n16606_));
  MX2X1    g14170(.A(new_n16606_), .B(new_n16605_), .S0(new_n12578_), .Y(new_n16607_));
  OR2X1    g14171(.A(new_n16604_), .B(pi0787), .Y(new_n16608_));
  OAI21X1  g14172(.A0(new_n16607_), .A1(new_n11763_), .B0(new_n16608_), .Y(new_n16609_));
  AOI21X1  g14173(.A0(new_n16609_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n16610_));
  INVX1    g14174(.A(new_n13568_), .Y(new_n16611_));
  OAI21X1  g14175(.A0(new_n11972_), .A1(new_n11970_), .B0(pi0603), .Y(new_n16612_));
  OR3X1    g14176(.A(new_n12043_), .B(new_n12042_), .C(new_n11881_), .Y(new_n16613_));
  MX2X1    g14177(.A(new_n16613_), .B(new_n16612_), .S0(new_n2933_), .Y(new_n16614_));
  MX2X1    g14178(.A(new_n12073_), .B(new_n16614_), .S0(new_n2939_), .Y(new_n16615_));
  INVX1    g14179(.A(new_n13565_), .Y(new_n16616_));
  OAI21X1  g14180(.A0(new_n16615_), .A1(pi0038), .B0(new_n16616_), .Y(new_n16617_));
  MX2X1    g14181(.A(new_n16617_), .B(new_n16611_), .S0(new_n6832_), .Y(new_n16618_));
  MX2X1    g14182(.A(new_n16618_), .B(new_n16587_), .S0(pi0742), .Y(new_n16619_));
  MX2X1    g14183(.A(new_n16619_), .B(new_n6832_), .S0(new_n11770_), .Y(new_n16620_));
  MX2X1    g14184(.A(new_n16620_), .B(new_n16579_), .S0(new_n12473_), .Y(new_n16621_));
  NOR2X1   g14185(.A(new_n16620_), .B(new_n12473_), .Y(new_n16622_));
  AOI22X1  g14186(.A0(new_n16622_), .A1(pi0609), .B0(new_n16580_), .B1(new_n12472_), .Y(new_n16623_));
  AOI22X1  g14187(.A0(new_n16622_), .A1(new_n12462_), .B0(new_n16580_), .B1(new_n12481_), .Y(new_n16624_));
  MX2X1    g14188(.A(new_n16624_), .B(new_n16623_), .S0(pi1155), .Y(new_n16625_));
  MX2X1    g14189(.A(new_n16625_), .B(new_n16621_), .S0(new_n11768_), .Y(new_n16626_));
  OAI21X1  g14190(.A0(new_n16580_), .A1(pi0618), .B0(pi1154), .Y(new_n16627_));
  AOI21X1  g14191(.A0(new_n16626_), .A1(pi0618), .B0(new_n16627_), .Y(new_n16628_));
  OAI21X1  g14192(.A0(new_n16580_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n16629_));
  AOI21X1  g14193(.A0(new_n16626_), .A1(new_n12486_), .B0(new_n16629_), .Y(new_n16630_));
  NOR2X1   g14194(.A(new_n16630_), .B(new_n16628_), .Y(new_n16631_));
  MX2X1    g14195(.A(new_n16631_), .B(new_n16626_), .S0(new_n11767_), .Y(new_n16632_));
  OR2X1    g14196(.A(new_n16632_), .B(pi0789), .Y(new_n16633_));
  OAI21X1  g14197(.A0(new_n16580_), .A1(pi0619), .B0(pi1159), .Y(new_n16634_));
  AOI21X1  g14198(.A0(new_n16632_), .A1(pi0619), .B0(new_n16634_), .Y(new_n16635_));
  OAI21X1  g14199(.A0(new_n16580_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n16636_));
  AOI21X1  g14200(.A0(new_n16632_), .A1(new_n12509_), .B0(new_n16636_), .Y(new_n16637_));
  OAI21X1  g14201(.A0(new_n16637_), .A1(new_n16635_), .B0(pi0789), .Y(new_n16638_));
  AND2X1   g14202(.A(new_n16638_), .B(new_n16633_), .Y(new_n16639_));
  MX2X1    g14203(.A(new_n16639_), .B(new_n16579_), .S0(new_n12708_), .Y(new_n16640_));
  MX2X1    g14204(.A(new_n16640_), .B(new_n16579_), .S0(new_n12580_), .Y(new_n16641_));
  MX2X1    g14205(.A(new_n16641_), .B(new_n16579_), .S0(new_n12604_), .Y(new_n16642_));
  AOI21X1  g14206(.A0(new_n16579_), .A1(new_n12612_), .B0(pi0715), .Y(new_n16643_));
  INVX1    g14207(.A(new_n16643_), .Y(new_n16644_));
  AOI21X1  g14208(.A0(new_n16642_), .A1(pi0644), .B0(new_n16644_), .Y(new_n16645_));
  OR3X1    g14209(.A(new_n16645_), .B(new_n16610_), .C(new_n11762_), .Y(new_n16646_));
  AOI21X1  g14210(.A0(new_n16609_), .A1(pi0644), .B0(pi0715), .Y(new_n16647_));
  OAI21X1  g14211(.A0(new_n16580_), .A1(new_n12612_), .B0(pi0715), .Y(new_n16648_));
  AOI21X1  g14212(.A0(new_n16642_), .A1(new_n12612_), .B0(new_n16648_), .Y(new_n16649_));
  OR2X1    g14213(.A(new_n16649_), .B(pi1160), .Y(new_n16650_));
  OAI21X1  g14214(.A0(new_n16650_), .A1(new_n16647_), .B0(new_n16646_), .Y(new_n16651_));
  AOI22X1  g14215(.A0(new_n16602_), .A1(new_n16373_), .B0(new_n16601_), .B1(new_n16374_), .Y(new_n16652_));
  OAI21X1  g14216(.A0(new_n16640_), .A1(new_n14250_), .B0(new_n16652_), .Y(new_n16653_));
  AOI21X1  g14217(.A0(new_n16638_), .A1(new_n16633_), .B0(pi0626), .Y(new_n16654_));
  OAI21X1  g14218(.A0(new_n16579_), .A1(new_n12542_), .B0(new_n16217_), .Y(new_n16655_));
  NOR2X1   g14219(.A(new_n16655_), .B(new_n16654_), .Y(new_n16656_));
  AOI21X1  g14220(.A0(new_n16638_), .A1(new_n16633_), .B0(new_n12542_), .Y(new_n16657_));
  OAI21X1  g14221(.A0(new_n16579_), .A1(pi0626), .B0(new_n16221_), .Y(new_n16658_));
  OAI22X1  g14222(.A0(new_n16658_), .A1(new_n16657_), .B0(new_n16599_), .B1(new_n13439_), .Y(new_n16659_));
  OAI21X1  g14223(.A0(new_n16659_), .A1(new_n16656_), .B0(pi0788), .Y(new_n16660_));
  MX2X1    g14224(.A(new_n12792_), .B(new_n16380_), .S0(pi0039), .Y(new_n16661_));
  MX2X1    g14225(.A(new_n16661_), .B(new_n13540_), .S0(pi0038), .Y(new_n16662_));
  INVX1    g14226(.A(new_n13547_), .Y(new_n16663_));
  OAI21X1  g14227(.A0(new_n13544_), .A1(pi0038), .B0(new_n16663_), .Y(new_n16664_));
  AOI21X1  g14228(.A0(new_n16664_), .A1(pi0176), .B0(new_n14897_), .Y(new_n16665_));
  OAI21X1  g14229(.A0(new_n16662_), .A1(pi0176), .B0(new_n16665_), .Y(new_n16666_));
  NOR2X1   g14230(.A(new_n13551_), .B(new_n2979_), .Y(new_n16667_));
  INVX1    g14231(.A(new_n16667_), .Y(new_n16668_));
  OAI21X1  g14232(.A0(new_n13553_), .A1(pi0038), .B0(new_n16668_), .Y(new_n16669_));
  OR3X1    g14233(.A(new_n13558_), .B(new_n13557_), .C(new_n13555_), .Y(new_n16670_));
  AOI21X1  g14234(.A0(new_n16670_), .A1(new_n6832_), .B0(pi0742), .Y(new_n16671_));
  OAI21X1  g14235(.A0(new_n16669_), .A1(new_n6832_), .B0(new_n16671_), .Y(new_n16672_));
  AND3X1   g14236(.A(new_n16672_), .B(new_n16666_), .C(new_n14896_), .Y(new_n16673_));
  INVX1    g14237(.A(new_n16673_), .Y(new_n16674_));
  AOI21X1  g14238(.A0(new_n16619_), .A1(pi0704), .B0(new_n11770_), .Y(new_n16675_));
  AOI22X1  g14239(.A0(new_n16675_), .A1(new_n16674_), .B0(new_n11770_), .B1(pi0176), .Y(new_n16676_));
  INVX1    g14240(.A(new_n16676_), .Y(new_n16677_));
  AOI21X1  g14241(.A0(new_n16620_), .A1(pi0625), .B0(pi1153), .Y(new_n16678_));
  OAI21X1  g14242(.A0(new_n16677_), .A1(pi0625), .B0(new_n16678_), .Y(new_n16679_));
  NOR2X1   g14243(.A(new_n16591_), .B(pi0608), .Y(new_n16680_));
  AOI21X1  g14244(.A0(new_n16620_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n16681_));
  OAI21X1  g14245(.A0(new_n16677_), .A1(new_n12363_), .B0(new_n16681_), .Y(new_n16682_));
  NOR2X1   g14246(.A(new_n16593_), .B(new_n12368_), .Y(new_n16683_));
  AOI22X1  g14247(.A0(new_n16683_), .A1(new_n16682_), .B0(new_n16680_), .B1(new_n16679_), .Y(new_n16684_));
  MX2X1    g14248(.A(new_n16684_), .B(new_n16677_), .S0(new_n11769_), .Y(new_n16685_));
  AOI21X1  g14249(.A0(new_n16595_), .A1(pi0609), .B0(pi1155), .Y(new_n16686_));
  OAI21X1  g14250(.A0(new_n16685_), .A1(pi0609), .B0(new_n16686_), .Y(new_n16687_));
  OAI21X1  g14251(.A0(new_n16623_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n16688_));
  INVX1    g14252(.A(new_n16688_), .Y(new_n16689_));
  AOI21X1  g14253(.A0(new_n16595_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n16690_));
  OAI21X1  g14254(.A0(new_n16685_), .A1(new_n12462_), .B0(new_n16690_), .Y(new_n16691_));
  OAI21X1  g14255(.A0(new_n16624_), .A1(pi1155), .B0(pi0660), .Y(new_n16692_));
  INVX1    g14256(.A(new_n16692_), .Y(new_n16693_));
  AOI22X1  g14257(.A0(new_n16693_), .A1(new_n16691_), .B0(new_n16689_), .B1(new_n16687_), .Y(new_n16694_));
  MX2X1    g14258(.A(new_n16694_), .B(new_n16685_), .S0(new_n11768_), .Y(new_n16695_));
  AOI21X1  g14259(.A0(new_n16596_), .A1(pi0618), .B0(pi1154), .Y(new_n16696_));
  OAI21X1  g14260(.A0(new_n16695_), .A1(pi0618), .B0(new_n16696_), .Y(new_n16697_));
  NOR2X1   g14261(.A(new_n16628_), .B(pi0627), .Y(new_n16698_));
  AOI21X1  g14262(.A0(new_n16596_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n16699_));
  OAI21X1  g14263(.A0(new_n16695_), .A1(new_n12486_), .B0(new_n16699_), .Y(new_n16700_));
  NOR2X1   g14264(.A(new_n16630_), .B(new_n12494_), .Y(new_n16701_));
  AOI22X1  g14265(.A0(new_n16701_), .A1(new_n16700_), .B0(new_n16698_), .B1(new_n16697_), .Y(new_n16702_));
  MX2X1    g14266(.A(new_n16702_), .B(new_n16695_), .S0(new_n11767_), .Y(new_n16703_));
  INVX1    g14267(.A(new_n16703_), .Y(new_n16704_));
  OAI21X1  g14268(.A0(new_n16598_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n16705_));
  AOI21X1  g14269(.A0(new_n16704_), .A1(new_n12509_), .B0(new_n16705_), .Y(new_n16706_));
  NOR3X1   g14270(.A(new_n16706_), .B(new_n16635_), .C(pi0648), .Y(new_n16707_));
  OAI21X1  g14271(.A0(new_n16598_), .A1(pi0619), .B0(pi1159), .Y(new_n16708_));
  AOI21X1  g14272(.A0(new_n16704_), .A1(pi0619), .B0(new_n16708_), .Y(new_n16709_));
  OR2X1    g14273(.A(new_n16637_), .B(new_n12517_), .Y(new_n16710_));
  OAI21X1  g14274(.A0(new_n16710_), .A1(new_n16709_), .B0(pi0789), .Y(new_n16711_));
  AOI21X1  g14275(.A0(new_n16703_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n16712_));
  OAI21X1  g14276(.A0(new_n16711_), .A1(new_n16707_), .B0(new_n16712_), .Y(new_n16713_));
  AOI22X1  g14277(.A0(new_n16713_), .A1(new_n16660_), .B0(new_n16653_), .B1(pi0792), .Y(new_n16714_));
  OAI21X1  g14278(.A0(new_n16653_), .A1(new_n14126_), .B0(new_n14122_), .Y(new_n16715_));
  OR2X1    g14279(.A(new_n16715_), .B(new_n16714_), .Y(new_n16716_));
  OR3X1    g14280(.A(new_n16649_), .B(pi1160), .C(pi0644), .Y(new_n16717_));
  OR3X1    g14281(.A(new_n16645_), .B(new_n11762_), .C(new_n12612_), .Y(new_n16718_));
  AND3X1   g14282(.A(new_n16718_), .B(new_n16717_), .C(pi0790), .Y(new_n16719_));
  OR2X1    g14283(.A(new_n16641_), .B(new_n14239_), .Y(new_n16720_));
  AOI22X1  g14284(.A0(new_n16606_), .A1(new_n14241_), .B0(new_n16605_), .B1(new_n14243_), .Y(new_n16721_));
  AOI21X1  g14285(.A0(new_n16721_), .A1(new_n16720_), .B0(new_n11763_), .Y(new_n16722_));
  NOR2X1   g14286(.A(new_n16722_), .B(new_n16719_), .Y(new_n16723_));
  AOI22X1  g14287(.A0(new_n16723_), .A1(new_n16716_), .B0(new_n16651_), .B1(pi0790), .Y(new_n16724_));
  AOI21X1  g14288(.A0(po1038), .A1(new_n6832_), .B0(pi0832), .Y(new_n16725_));
  OAI21X1  g14289(.A0(new_n16724_), .A1(po1038), .B0(new_n16725_), .Y(new_n16726_));
  AND2X1   g14290(.A(new_n16726_), .B(new_n16578_), .Y(po0333));
  OR2X1    g14291(.A(new_n3103_), .B(new_n7450_), .Y(new_n16728_));
  MX2X1    g14292(.A(new_n16611_), .B(new_n12832_), .S0(pi0757), .Y(new_n16729_));
  AOI21X1  g14293(.A0(new_n16616_), .A1(new_n7450_), .B0(pi0757), .Y(new_n16730_));
  AOI22X1  g14294(.A0(new_n16730_), .A1(new_n16617_), .B0(new_n16729_), .B1(new_n7450_), .Y(new_n16731_));
  OAI21X1  g14295(.A0(new_n13544_), .A1(new_n7450_), .B0(new_n2979_), .Y(new_n16732_));
  AOI21X1  g14296(.A0(new_n13542_), .A1(new_n7450_), .B0(new_n16732_), .Y(new_n16733_));
  OAI21X1  g14297(.A0(new_n12077_), .A1(pi0177), .B0(new_n12806_), .Y(new_n16734_));
  AND2X1   g14298(.A(new_n16734_), .B(pi0757), .Y(new_n16735_));
  INVX1    g14299(.A(new_n16735_), .Y(new_n16736_));
  AND2X1   g14300(.A(new_n13553_), .B(pi0177), .Y(new_n16737_));
  MX2X1    g14301(.A(new_n13556_), .B(new_n12788_), .S0(pi0039), .Y(new_n16738_));
  AND2X1   g14302(.A(new_n16738_), .B(new_n7450_), .Y(new_n16739_));
  OR2X1    g14303(.A(new_n16739_), .B(pi0038), .Y(new_n16740_));
  AOI21X1  g14304(.A0(new_n12276_), .A1(new_n2939_), .B0(pi0177), .Y(new_n16741_));
  AND2X1   g14305(.A(new_n13551_), .B(pi0177), .Y(new_n16742_));
  OR3X1    g14306(.A(new_n16742_), .B(new_n16741_), .C(new_n2979_), .Y(new_n16743_));
  AND2X1   g14307(.A(new_n16743_), .B(new_n14928_), .Y(new_n16744_));
  OAI21X1  g14308(.A0(new_n16740_), .A1(new_n16737_), .B0(new_n16744_), .Y(new_n16745_));
  OAI21X1  g14309(.A0(new_n16736_), .A1(new_n16733_), .B0(new_n16745_), .Y(new_n16746_));
  AOI21X1  g14310(.A0(new_n16746_), .A1(new_n14935_), .B0(new_n11770_), .Y(new_n16747_));
  OAI21X1  g14311(.A0(new_n16731_), .A1(new_n14935_), .B0(new_n16747_), .Y(new_n16748_));
  AND3X1   g14312(.A(new_n16748_), .B(new_n16728_), .C(new_n12363_), .Y(new_n16749_));
  MX2X1    g14313(.A(new_n16731_), .B(pi0177), .S0(new_n11770_), .Y(new_n16750_));
  OAI21X1  g14314(.A0(new_n16750_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n16751_));
  OAI21X1  g14315(.A0(new_n12826_), .A1(new_n7450_), .B0(new_n2979_), .Y(new_n16752_));
  AOI21X1  g14316(.A0(new_n12825_), .A1(new_n7450_), .B0(new_n16752_), .Y(new_n16753_));
  AOI21X1  g14317(.A0(new_n12771_), .A1(new_n7450_), .B0(new_n12441_), .Y(new_n16754_));
  NOR3X1   g14318(.A(new_n16754_), .B(new_n16753_), .C(pi0686), .Y(new_n16755_));
  AND2X1   g14319(.A(pi0686), .B(new_n7450_), .Y(new_n16756_));
  INVX1    g14320(.A(new_n16756_), .Y(new_n16757_));
  OAI21X1  g14321(.A0(new_n16757_), .A1(new_n12447_), .B0(new_n3103_), .Y(new_n16758_));
  OAI21X1  g14322(.A0(new_n16758_), .A1(new_n16755_), .B0(new_n16728_), .Y(new_n16759_));
  OR2X1    g14323(.A(new_n16759_), .B(new_n12363_), .Y(new_n16760_));
  AOI21X1  g14324(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0177), .Y(new_n16761_));
  AOI21X1  g14325(.A0(new_n16761_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n16762_));
  AOI21X1  g14326(.A0(new_n16762_), .A1(new_n16760_), .B0(pi0608), .Y(new_n16763_));
  OAI21X1  g14327(.A0(new_n16751_), .A1(new_n16749_), .B0(new_n16763_), .Y(new_n16764_));
  AND3X1   g14328(.A(new_n16748_), .B(new_n16728_), .C(pi0625), .Y(new_n16765_));
  OAI21X1  g14329(.A0(new_n16750_), .A1(pi0625), .B0(pi1153), .Y(new_n16766_));
  OR2X1    g14330(.A(new_n16759_), .B(pi0625), .Y(new_n16767_));
  AOI21X1  g14331(.A0(new_n16761_), .A1(pi0625), .B0(pi1153), .Y(new_n16768_));
  AOI21X1  g14332(.A0(new_n16768_), .A1(new_n16767_), .B0(new_n12368_), .Y(new_n16769_));
  OAI21X1  g14333(.A0(new_n16766_), .A1(new_n16765_), .B0(new_n16769_), .Y(new_n16770_));
  AOI21X1  g14334(.A0(new_n16770_), .A1(new_n16764_), .B0(new_n11769_), .Y(new_n16771_));
  AND3X1   g14335(.A(new_n16748_), .B(new_n16728_), .C(new_n11769_), .Y(new_n16772_));
  NOR2X1   g14336(.A(new_n16772_), .B(new_n16771_), .Y(new_n16773_));
  NAND2X1  g14337(.A(new_n16759_), .B(new_n11769_), .Y(new_n16774_));
  AOI22X1  g14338(.A0(new_n16768_), .A1(new_n16767_), .B0(new_n16762_), .B1(new_n16760_), .Y(new_n16775_));
  OR2X1    g14339(.A(new_n16775_), .B(new_n11769_), .Y(new_n16776_));
  AND2X1   g14340(.A(new_n16776_), .B(new_n16774_), .Y(new_n16777_));
  AOI21X1  g14341(.A0(new_n16777_), .A1(pi0609), .B0(pi1155), .Y(new_n16778_));
  OAI21X1  g14342(.A0(new_n16773_), .A1(pi0609), .B0(new_n16778_), .Y(new_n16779_));
  INVX1    g14343(.A(new_n16761_), .Y(new_n16780_));
  AND2X1   g14344(.A(new_n16750_), .B(new_n12474_), .Y(new_n16781_));
  AOI22X1  g14345(.A0(new_n16781_), .A1(pi0609), .B0(new_n16780_), .B1(new_n12472_), .Y(new_n16782_));
  OR2X1    g14346(.A(new_n16782_), .B(new_n12463_), .Y(new_n16783_));
  AND2X1   g14347(.A(new_n16783_), .B(new_n12468_), .Y(new_n16784_));
  AOI21X1  g14348(.A0(new_n16777_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n16785_));
  OAI21X1  g14349(.A0(new_n16773_), .A1(new_n12462_), .B0(new_n16785_), .Y(new_n16786_));
  AOI22X1  g14350(.A0(new_n16781_), .A1(new_n12462_), .B0(new_n16780_), .B1(new_n12481_), .Y(new_n16787_));
  OR2X1    g14351(.A(new_n16787_), .B(pi1155), .Y(new_n16788_));
  AND2X1   g14352(.A(new_n16788_), .B(pi0660), .Y(new_n16789_));
  AOI22X1  g14353(.A0(new_n16789_), .A1(new_n16786_), .B0(new_n16784_), .B1(new_n16779_), .Y(new_n16790_));
  OAI21X1  g14354(.A0(new_n16772_), .A1(new_n16771_), .B0(new_n11768_), .Y(new_n16791_));
  OAI21X1  g14355(.A0(new_n16790_), .A1(new_n11768_), .B0(new_n16791_), .Y(new_n16792_));
  OR2X1    g14356(.A(new_n16761_), .B(new_n13910_), .Y(new_n16793_));
  OAI21X1  g14357(.A0(new_n16777_), .A1(new_n12490_), .B0(new_n16793_), .Y(new_n16794_));
  OAI21X1  g14358(.A0(new_n16794_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n16795_));
  AOI21X1  g14359(.A0(new_n16792_), .A1(new_n12486_), .B0(new_n16795_), .Y(new_n16796_));
  AOI21X1  g14360(.A0(new_n16780_), .A1(new_n12473_), .B0(new_n16781_), .Y(new_n16797_));
  MX2X1    g14361(.A(new_n16787_), .B(new_n16782_), .S0(pi1155), .Y(new_n16798_));
  MX2X1    g14362(.A(new_n16798_), .B(new_n16797_), .S0(new_n11768_), .Y(new_n16799_));
  OAI21X1  g14363(.A0(new_n16780_), .A1(pi0618), .B0(pi1154), .Y(new_n16800_));
  AOI21X1  g14364(.A0(new_n16799_), .A1(pi0618), .B0(new_n16800_), .Y(new_n16801_));
  OR2X1    g14365(.A(new_n16801_), .B(pi0627), .Y(new_n16802_));
  OAI21X1  g14366(.A0(new_n16794_), .A1(pi0618), .B0(pi1154), .Y(new_n16803_));
  AOI21X1  g14367(.A0(new_n16792_), .A1(pi0618), .B0(new_n16803_), .Y(new_n16804_));
  OAI21X1  g14368(.A0(new_n16780_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n16805_));
  AOI21X1  g14369(.A0(new_n16799_), .A1(new_n12486_), .B0(new_n16805_), .Y(new_n16806_));
  OR2X1    g14370(.A(new_n16806_), .B(new_n12494_), .Y(new_n16807_));
  OAI22X1  g14371(.A0(new_n16807_), .A1(new_n16804_), .B0(new_n16802_), .B1(new_n16796_), .Y(new_n16808_));
  MX2X1    g14372(.A(new_n16808_), .B(new_n16792_), .S0(new_n11767_), .Y(new_n16809_));
  MX2X1    g14373(.A(new_n16794_), .B(new_n16780_), .S0(new_n12513_), .Y(new_n16810_));
  OAI21X1  g14374(.A0(new_n16810_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n16811_));
  AOI21X1  g14375(.A0(new_n16809_), .A1(new_n12509_), .B0(new_n16811_), .Y(new_n16812_));
  OR2X1    g14376(.A(new_n16799_), .B(pi0781), .Y(new_n16813_));
  OAI21X1  g14377(.A0(new_n16806_), .A1(new_n16801_), .B0(pi0781), .Y(new_n16814_));
  NAND3X1  g14378(.A(new_n16814_), .B(new_n16813_), .C(pi0619), .Y(new_n16815_));
  AOI21X1  g14379(.A0(new_n16761_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n16816_));
  AND2X1   g14380(.A(new_n16816_), .B(new_n16815_), .Y(new_n16817_));
  OR2X1    g14381(.A(new_n16817_), .B(pi0648), .Y(new_n16818_));
  OAI21X1  g14382(.A0(new_n16810_), .A1(pi0619), .B0(pi1159), .Y(new_n16819_));
  AOI21X1  g14383(.A0(new_n16809_), .A1(pi0619), .B0(new_n16819_), .Y(new_n16820_));
  NAND3X1  g14384(.A(new_n16814_), .B(new_n16813_), .C(new_n12509_), .Y(new_n16821_));
  AOI21X1  g14385(.A0(new_n16761_), .A1(pi0619), .B0(pi1159), .Y(new_n16822_));
  AND2X1   g14386(.A(new_n16822_), .B(new_n16821_), .Y(new_n16823_));
  OR2X1    g14387(.A(new_n16823_), .B(new_n12517_), .Y(new_n16824_));
  OAI22X1  g14388(.A0(new_n16824_), .A1(new_n16820_), .B0(new_n16818_), .B1(new_n16812_), .Y(new_n16825_));
  MX2X1    g14389(.A(new_n16825_), .B(new_n16809_), .S0(new_n11766_), .Y(new_n16826_));
  MX2X1    g14390(.A(new_n16810_), .B(new_n16780_), .S0(new_n12531_), .Y(new_n16827_));
  AOI21X1  g14391(.A0(new_n16827_), .A1(pi0626), .B0(pi0641), .Y(new_n16828_));
  OAI21X1  g14392(.A0(new_n16826_), .A1(pi0626), .B0(new_n16828_), .Y(new_n16829_));
  AND2X1   g14393(.A(new_n16814_), .B(new_n16813_), .Y(new_n16830_));
  AOI22X1  g14394(.A0(new_n16822_), .A1(new_n16821_), .B0(new_n16816_), .B1(new_n16815_), .Y(new_n16831_));
  MX2X1    g14395(.A(new_n16831_), .B(new_n16830_), .S0(new_n11766_), .Y(new_n16832_));
  AOI21X1  g14396(.A0(new_n16780_), .A1(pi0626), .B0(new_n12543_), .Y(new_n16833_));
  OAI21X1  g14397(.A0(new_n16832_), .A1(pi0626), .B0(new_n16833_), .Y(new_n16834_));
  AND2X1   g14398(.A(new_n16834_), .B(new_n12548_), .Y(new_n16835_));
  AOI21X1  g14399(.A0(new_n16827_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n16836_));
  OAI21X1  g14400(.A0(new_n16826_), .A1(new_n12542_), .B0(new_n16836_), .Y(new_n16837_));
  AOI21X1  g14401(.A0(new_n16780_), .A1(new_n12542_), .B0(pi0641), .Y(new_n16838_));
  OAI21X1  g14402(.A0(new_n16832_), .A1(new_n12542_), .B0(new_n16838_), .Y(new_n16839_));
  AND2X1   g14403(.A(new_n16839_), .B(pi1158), .Y(new_n16840_));
  AOI22X1  g14404(.A0(new_n16840_), .A1(new_n16837_), .B0(new_n16835_), .B1(new_n16829_), .Y(new_n16841_));
  MX2X1    g14405(.A(new_n16841_), .B(new_n16826_), .S0(new_n11765_), .Y(new_n16842_));
  MX2X1    g14406(.A(new_n16832_), .B(new_n16761_), .S0(new_n12708_), .Y(new_n16843_));
  INVX1    g14407(.A(new_n16843_), .Y(new_n16844_));
  OAI21X1  g14408(.A0(new_n16844_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n16845_));
  AOI21X1  g14409(.A0(new_n16842_), .A1(new_n12554_), .B0(new_n16845_), .Y(new_n16846_));
  MX2X1    g14410(.A(new_n16827_), .B(new_n16780_), .S0(new_n12563_), .Y(new_n16847_));
  AOI21X1  g14411(.A0(new_n16761_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n16848_));
  OAI21X1  g14412(.A0(new_n16847_), .A1(new_n12554_), .B0(new_n16848_), .Y(new_n16849_));
  NAND2X1  g14413(.A(new_n16849_), .B(new_n12561_), .Y(new_n16850_));
  OAI21X1  g14414(.A0(new_n16844_), .A1(pi0628), .B0(pi1156), .Y(new_n16851_));
  AOI21X1  g14415(.A0(new_n16842_), .A1(pi0628), .B0(new_n16851_), .Y(new_n16852_));
  AOI21X1  g14416(.A0(new_n16761_), .A1(pi0628), .B0(pi1156), .Y(new_n16853_));
  OAI21X1  g14417(.A0(new_n16847_), .A1(pi0628), .B0(new_n16853_), .Y(new_n16854_));
  NAND2X1  g14418(.A(new_n16854_), .B(pi0629), .Y(new_n16855_));
  OAI22X1  g14419(.A0(new_n16855_), .A1(new_n16852_), .B0(new_n16850_), .B1(new_n16846_), .Y(new_n16856_));
  AND2X1   g14420(.A(new_n16842_), .B(new_n11764_), .Y(new_n16857_));
  AOI21X1  g14421(.A0(new_n16856_), .A1(pi0792), .B0(new_n16857_), .Y(new_n16858_));
  MX2X1    g14422(.A(new_n16844_), .B(new_n16780_), .S0(new_n12580_), .Y(new_n16859_));
  INVX1    g14423(.A(new_n16859_), .Y(new_n16860_));
  AOI21X1  g14424(.A0(new_n16860_), .A1(pi0647), .B0(pi1157), .Y(new_n16861_));
  OAI21X1  g14425(.A0(new_n16858_), .A1(pi0647), .B0(new_n16861_), .Y(new_n16862_));
  INVX1    g14426(.A(new_n16847_), .Y(new_n16863_));
  AND2X1   g14427(.A(new_n16854_), .B(new_n16849_), .Y(new_n16864_));
  MX2X1    g14428(.A(new_n16864_), .B(new_n16863_), .S0(new_n11764_), .Y(new_n16865_));
  INVX1    g14429(.A(new_n16865_), .Y(new_n16866_));
  AOI21X1  g14430(.A0(new_n16761_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n16867_));
  OAI21X1  g14431(.A0(new_n16866_), .A1(new_n12577_), .B0(new_n16867_), .Y(new_n16868_));
  AND2X1   g14432(.A(new_n16868_), .B(new_n12592_), .Y(new_n16869_));
  AOI21X1  g14433(.A0(new_n16860_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n16870_));
  OAI21X1  g14434(.A0(new_n16858_), .A1(new_n12577_), .B0(new_n16870_), .Y(new_n16871_));
  AOI21X1  g14435(.A0(new_n16761_), .A1(pi0647), .B0(pi1157), .Y(new_n16872_));
  OAI21X1  g14436(.A0(new_n16866_), .A1(pi0647), .B0(new_n16872_), .Y(new_n16873_));
  AND2X1   g14437(.A(new_n16873_), .B(pi0630), .Y(new_n16874_));
  AOI22X1  g14438(.A0(new_n16874_), .A1(new_n16871_), .B0(new_n16869_), .B1(new_n16862_), .Y(new_n16875_));
  MX2X1    g14439(.A(new_n16875_), .B(new_n16858_), .S0(new_n11763_), .Y(new_n16876_));
  AND2X1   g14440(.A(new_n16873_), .B(new_n16868_), .Y(new_n16877_));
  MX2X1    g14441(.A(new_n16877_), .B(new_n16865_), .S0(new_n11763_), .Y(new_n16878_));
  AOI21X1  g14442(.A0(new_n16878_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n16879_));
  OAI21X1  g14443(.A0(new_n16876_), .A1(new_n12612_), .B0(new_n16879_), .Y(new_n16880_));
  MX2X1    g14444(.A(new_n16860_), .B(new_n16761_), .S0(new_n12604_), .Y(new_n16881_));
  OAI21X1  g14445(.A0(new_n16780_), .A1(pi0644), .B0(new_n12608_), .Y(new_n16882_));
  AOI21X1  g14446(.A0(new_n16881_), .A1(pi0644), .B0(new_n16882_), .Y(new_n16883_));
  NOR2X1   g14447(.A(new_n16883_), .B(new_n11762_), .Y(new_n16884_));
  AND2X1   g14448(.A(new_n16884_), .B(new_n16880_), .Y(new_n16885_));
  OR2X1    g14449(.A(new_n16858_), .B(pi0787), .Y(new_n16886_));
  OAI21X1  g14450(.A0(new_n16875_), .A1(new_n11763_), .B0(new_n16886_), .Y(new_n16887_));
  AND2X1   g14451(.A(new_n16878_), .B(pi0644), .Y(new_n16888_));
  OR2X1    g14452(.A(new_n16888_), .B(pi0715), .Y(new_n16889_));
  AOI21X1  g14453(.A0(new_n16887_), .A1(new_n12612_), .B0(new_n16889_), .Y(new_n16890_));
  OAI21X1  g14454(.A0(new_n16780_), .A1(new_n12612_), .B0(pi0715), .Y(new_n16891_));
  AOI21X1  g14455(.A0(new_n16881_), .A1(new_n12612_), .B0(new_n16891_), .Y(new_n16892_));
  OR2X1    g14456(.A(new_n16892_), .B(pi1160), .Y(new_n16893_));
  OAI21X1  g14457(.A0(new_n16893_), .A1(new_n16890_), .B0(pi0790), .Y(new_n16894_));
  AOI21X1  g14458(.A0(new_n16876_), .A1(new_n12766_), .B0(po1038), .Y(new_n16895_));
  OAI21X1  g14459(.A0(new_n16894_), .A1(new_n16885_), .B0(new_n16895_), .Y(new_n16896_));
  AOI21X1  g14460(.A0(po1038), .A1(new_n7450_), .B0(pi0832), .Y(new_n16897_));
  AOI21X1  g14461(.A0(pi1093), .A1(pi1092), .B0(pi0177), .Y(new_n16898_));
  INVX1    g14462(.A(new_n16898_), .Y(new_n16899_));
  AOI21X1  g14463(.A0(new_n12056_), .A1(new_n14928_), .B0(new_n16898_), .Y(new_n16900_));
  AOI21X1  g14464(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n16900_), .Y(new_n16901_));
  INVX1    g14465(.A(new_n16900_), .Y(new_n16902_));
  AOI21X1  g14466(.A0(new_n16902_), .A1(new_n14331_), .B0(new_n12463_), .Y(new_n16903_));
  AOI21X1  g14467(.A0(new_n16901_), .A1(new_n12646_), .B0(pi1155), .Y(new_n16904_));
  OAI21X1  g14468(.A0(new_n16904_), .A1(new_n16903_), .B0(pi0785), .Y(new_n16905_));
  OAI21X1  g14469(.A0(new_n16901_), .A1(pi0785), .B0(new_n16905_), .Y(new_n16906_));
  INVX1    g14470(.A(new_n16906_), .Y(new_n16907_));
  AOI21X1  g14471(.A0(new_n16907_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n16908_));
  AOI21X1  g14472(.A0(new_n16907_), .A1(new_n12655_), .B0(pi1154), .Y(new_n16909_));
  NOR2X1   g14473(.A(new_n16909_), .B(new_n16908_), .Y(new_n16910_));
  MX2X1    g14474(.A(new_n16910_), .B(new_n16907_), .S0(new_n11767_), .Y(new_n16911_));
  NOR2X1   g14475(.A(new_n16911_), .B(pi0789), .Y(new_n16912_));
  INVX1    g14476(.A(new_n16911_), .Y(new_n16913_));
  AOI21X1  g14477(.A0(new_n16898_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n16914_));
  OAI21X1  g14478(.A0(new_n16913_), .A1(new_n12509_), .B0(new_n16914_), .Y(new_n16915_));
  AOI21X1  g14479(.A0(new_n16898_), .A1(pi0619), .B0(pi1159), .Y(new_n16916_));
  OAI21X1  g14480(.A0(new_n16913_), .A1(pi0619), .B0(new_n16916_), .Y(new_n16917_));
  AOI21X1  g14481(.A0(new_n16917_), .A1(new_n16915_), .B0(new_n11766_), .Y(new_n16918_));
  NOR2X1   g14482(.A(new_n16918_), .B(new_n16912_), .Y(new_n16919_));
  INVX1    g14483(.A(new_n16919_), .Y(new_n16920_));
  MX2X1    g14484(.A(new_n16920_), .B(new_n16899_), .S0(new_n12708_), .Y(new_n16921_));
  MX2X1    g14485(.A(new_n16921_), .B(new_n16899_), .S0(new_n12580_), .Y(new_n16922_));
  AOI21X1  g14486(.A0(new_n12439_), .A1(new_n14935_), .B0(new_n16898_), .Y(new_n16923_));
  AND3X1   g14487(.A(new_n12439_), .B(new_n14935_), .C(new_n12363_), .Y(new_n16924_));
  NOR2X1   g14488(.A(new_n16924_), .B(new_n16923_), .Y(new_n16925_));
  NOR2X1   g14489(.A(new_n16898_), .B(pi1153), .Y(new_n16926_));
  INVX1    g14490(.A(new_n16926_), .Y(new_n16927_));
  OAI22X1  g14491(.A0(new_n16927_), .A1(new_n16924_), .B0(new_n16925_), .B1(new_n12364_), .Y(new_n16928_));
  MX2X1    g14492(.A(new_n16928_), .B(new_n16923_), .S0(new_n11769_), .Y(new_n16929_));
  NOR4X1   g14493(.A(new_n16929_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n16930_));
  AND3X1   g14494(.A(new_n16930_), .B(new_n12739_), .C(new_n12718_), .Y(new_n16931_));
  INVX1    g14495(.A(new_n16931_), .Y(new_n16932_));
  AOI21X1  g14496(.A0(new_n16898_), .A1(pi0647), .B0(pi1157), .Y(new_n16933_));
  OAI21X1  g14497(.A0(new_n16932_), .A1(pi0647), .B0(new_n16933_), .Y(new_n16934_));
  MX2X1    g14498(.A(new_n16931_), .B(new_n16898_), .S0(new_n12577_), .Y(new_n16935_));
  OAI22X1  g14499(.A0(new_n16935_), .A1(new_n14242_), .B0(new_n16934_), .B1(new_n12592_), .Y(new_n16936_));
  AOI21X1  g14500(.A0(new_n16922_), .A1(new_n14326_), .B0(new_n16936_), .Y(new_n16937_));
  AOI21X1  g14501(.A0(new_n16899_), .A1(pi0626), .B0(new_n16218_), .Y(new_n16938_));
  OAI21X1  g14502(.A0(new_n16919_), .A1(pi0626), .B0(new_n16938_), .Y(new_n16939_));
  AOI21X1  g14503(.A0(new_n16899_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n16940_));
  OAI21X1  g14504(.A0(new_n16919_), .A1(new_n12542_), .B0(new_n16940_), .Y(new_n16941_));
  NAND2X1  g14505(.A(new_n16930_), .B(new_n12637_), .Y(new_n16942_));
  AND3X1   g14506(.A(new_n16942_), .B(new_n16941_), .C(new_n16939_), .Y(new_n16943_));
  NOR2X1   g14507(.A(new_n16943_), .B(new_n11765_), .Y(new_n16944_));
  INVX1    g14508(.A(new_n16944_), .Y(new_n16945_));
  NOR2X1   g14509(.A(new_n16923_), .B(new_n11991_), .Y(new_n16946_));
  MX2X1    g14510(.A(new_n16902_), .B(new_n12363_), .S0(new_n16946_), .Y(new_n16947_));
  NOR2X1   g14511(.A(new_n16947_), .B(new_n16927_), .Y(new_n16948_));
  OAI21X1  g14512(.A0(new_n16925_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n16949_));
  NOR2X1   g14513(.A(new_n16949_), .B(new_n16948_), .Y(new_n16950_));
  OR3X1    g14514(.A(new_n16923_), .B(new_n11991_), .C(new_n12363_), .Y(new_n16951_));
  AND2X1   g14515(.A(new_n16900_), .B(pi1153), .Y(new_n16952_));
  OAI21X1  g14516(.A0(new_n16927_), .A1(new_n16924_), .B0(pi0608), .Y(new_n16953_));
  AOI21X1  g14517(.A0(new_n16952_), .A1(new_n16951_), .B0(new_n16953_), .Y(new_n16954_));
  OAI21X1  g14518(.A0(new_n16954_), .A1(new_n16950_), .B0(pi0778), .Y(new_n16955_));
  OAI21X1  g14519(.A0(new_n16946_), .A1(new_n16902_), .B0(new_n11769_), .Y(new_n16956_));
  NAND2X1  g14520(.A(new_n16956_), .B(new_n16955_), .Y(new_n16957_));
  INVX1    g14521(.A(new_n16957_), .Y(new_n16958_));
  OAI21X1  g14522(.A0(new_n16929_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n16959_));
  AOI21X1  g14523(.A0(new_n16957_), .A1(new_n12462_), .B0(new_n16959_), .Y(new_n16960_));
  NOR3X1   g14524(.A(new_n16960_), .B(new_n16903_), .C(pi0660), .Y(new_n16961_));
  OAI21X1  g14525(.A0(new_n16929_), .A1(pi0609), .B0(pi1155), .Y(new_n16962_));
  AOI21X1  g14526(.A0(new_n16957_), .A1(pi0609), .B0(new_n16962_), .Y(new_n16963_));
  NOR3X1   g14527(.A(new_n16963_), .B(new_n16904_), .C(new_n12468_), .Y(new_n16964_));
  NOR2X1   g14528(.A(new_n16964_), .B(new_n16961_), .Y(new_n16965_));
  MX2X1    g14529(.A(new_n16965_), .B(new_n16958_), .S0(new_n11768_), .Y(new_n16966_));
  OR3X1    g14530(.A(new_n16929_), .B(new_n12630_), .C(new_n12486_), .Y(new_n16967_));
  AND2X1   g14531(.A(new_n16967_), .B(new_n12487_), .Y(new_n16968_));
  OAI21X1  g14532(.A0(new_n16966_), .A1(pi0618), .B0(new_n16968_), .Y(new_n16969_));
  NOR2X1   g14533(.A(new_n16908_), .B(pi0627), .Y(new_n16970_));
  NOR3X1   g14534(.A(new_n16929_), .B(new_n12630_), .C(pi0618), .Y(new_n16971_));
  NOR2X1   g14535(.A(new_n16971_), .B(new_n12487_), .Y(new_n16972_));
  OAI21X1  g14536(.A0(new_n16966_), .A1(new_n12486_), .B0(new_n16972_), .Y(new_n16973_));
  NOR2X1   g14537(.A(new_n16909_), .B(new_n12494_), .Y(new_n16974_));
  AOI22X1  g14538(.A0(new_n16974_), .A1(new_n16973_), .B0(new_n16970_), .B1(new_n16969_), .Y(new_n16975_));
  MX2X1    g14539(.A(new_n16975_), .B(new_n16966_), .S0(new_n11767_), .Y(new_n16976_));
  OR4X1    g14540(.A(new_n16929_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n16977_));
  AND2X1   g14541(.A(new_n16977_), .B(new_n12510_), .Y(new_n16978_));
  OAI21X1  g14542(.A0(new_n16976_), .A1(pi0619), .B0(new_n16978_), .Y(new_n16979_));
  AND3X1   g14543(.A(new_n16979_), .B(new_n16915_), .C(new_n12517_), .Y(new_n16980_));
  NOR4X1   g14544(.A(new_n16929_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n16981_));
  NOR2X1   g14545(.A(new_n16981_), .B(new_n12510_), .Y(new_n16982_));
  OAI21X1  g14546(.A0(new_n16976_), .A1(new_n12509_), .B0(new_n16982_), .Y(new_n16983_));
  AND2X1   g14547(.A(new_n16917_), .B(pi0648), .Y(new_n16984_));
  AOI21X1  g14548(.A0(new_n16984_), .A1(new_n16983_), .B0(new_n11766_), .Y(new_n16985_));
  INVX1    g14549(.A(new_n16985_), .Y(new_n16986_));
  AOI21X1  g14550(.A0(new_n16976_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n16987_));
  OAI21X1  g14551(.A0(new_n16986_), .A1(new_n16980_), .B0(new_n16987_), .Y(new_n16988_));
  AOI21X1  g14552(.A0(new_n16988_), .A1(new_n16945_), .B0(new_n14125_), .Y(new_n16989_));
  INVX1    g14553(.A(new_n16921_), .Y(new_n16990_));
  AND2X1   g14554(.A(new_n16930_), .B(new_n12718_), .Y(new_n16991_));
  AOI22X1  g14555(.A0(new_n16991_), .A1(new_n14426_), .B0(new_n16990_), .B1(new_n12735_), .Y(new_n16992_));
  AOI22X1  g14556(.A0(new_n16991_), .A1(new_n14428_), .B0(new_n16990_), .B1(new_n12733_), .Y(new_n16993_));
  MX2X1    g14557(.A(new_n16993_), .B(new_n16992_), .S0(new_n12561_), .Y(new_n16994_));
  OAI21X1  g14558(.A0(new_n16994_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n16995_));
  OAI22X1  g14559(.A0(new_n16995_), .A1(new_n16989_), .B0(new_n16937_), .B1(new_n11763_), .Y(new_n16996_));
  INVX1    g14560(.A(new_n16996_), .Y(new_n16997_));
  OAI21X1  g14561(.A0(new_n16935_), .A1(new_n12578_), .B0(new_n16934_), .Y(new_n16998_));
  MX2X1    g14562(.A(new_n16998_), .B(new_n16932_), .S0(new_n11763_), .Y(new_n16999_));
  OAI21X1  g14563(.A0(new_n16999_), .A1(pi0644), .B0(pi0715), .Y(new_n17000_));
  AOI21X1  g14564(.A0(new_n16997_), .A1(pi0644), .B0(new_n17000_), .Y(new_n17001_));
  OR3X1    g14565(.A(new_n16899_), .B(new_n12603_), .C(new_n11763_), .Y(new_n17002_));
  OAI21X1  g14566(.A0(new_n16922_), .A1(new_n12604_), .B0(new_n17002_), .Y(new_n17003_));
  OAI21X1  g14567(.A0(new_n16899_), .A1(pi0644), .B0(new_n12608_), .Y(new_n17004_));
  AOI21X1  g14568(.A0(new_n17003_), .A1(pi0644), .B0(new_n17004_), .Y(new_n17005_));
  OR2X1    g14569(.A(new_n17005_), .B(new_n11762_), .Y(new_n17006_));
  OAI21X1  g14570(.A0(new_n16999_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17007_));
  AOI21X1  g14571(.A0(new_n16997_), .A1(new_n12612_), .B0(new_n17007_), .Y(new_n17008_));
  OAI21X1  g14572(.A0(new_n16899_), .A1(new_n12612_), .B0(pi0715), .Y(new_n17009_));
  AOI21X1  g14573(.A0(new_n17003_), .A1(new_n12612_), .B0(new_n17009_), .Y(new_n17010_));
  OR2X1    g14574(.A(new_n17010_), .B(pi1160), .Y(new_n17011_));
  OAI22X1  g14575(.A0(new_n17011_), .A1(new_n17008_), .B0(new_n17006_), .B1(new_n17001_), .Y(new_n17012_));
  OAI21X1  g14576(.A0(new_n16996_), .A1(pi0790), .B0(pi0832), .Y(new_n17013_));
  AOI21X1  g14577(.A0(new_n17012_), .A1(pi0790), .B0(new_n17013_), .Y(new_n17014_));
  AOI21X1  g14578(.A0(new_n16897_), .A1(new_n16896_), .B0(new_n17014_), .Y(po0334));
  AOI21X1  g14579(.A0(pi1093), .A1(pi1092), .B0(pi0178), .Y(new_n17016_));
  INVX1    g14580(.A(new_n17016_), .Y(new_n17017_));
  AOI21X1  g14581(.A0(new_n12056_), .A1(new_n14970_), .B0(new_n17016_), .Y(new_n17018_));
  INVX1    g14582(.A(new_n17018_), .Y(new_n17019_));
  NAND2X1  g14583(.A(new_n17019_), .B(new_n15771_), .Y(new_n17020_));
  AND3X1   g14584(.A(new_n12480_), .B(new_n12056_), .C(new_n14970_), .Y(new_n17021_));
  OAI21X1  g14585(.A0(new_n17021_), .A1(new_n17020_), .B0(pi1155), .Y(new_n17022_));
  NOR3X1   g14586(.A(new_n17021_), .B(new_n17016_), .C(pi1155), .Y(new_n17023_));
  INVX1    g14587(.A(new_n17023_), .Y(new_n17024_));
  AOI21X1  g14588(.A0(new_n17024_), .A1(new_n17022_), .B0(new_n11768_), .Y(new_n17025_));
  AOI21X1  g14589(.A0(new_n17020_), .A1(new_n11768_), .B0(new_n17025_), .Y(new_n17026_));
  AOI21X1  g14590(.A0(new_n17026_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n17027_));
  AOI21X1  g14591(.A0(new_n17026_), .A1(new_n12655_), .B0(pi1154), .Y(new_n17028_));
  NOR2X1   g14592(.A(new_n17028_), .B(new_n17027_), .Y(new_n17029_));
  MX2X1    g14593(.A(new_n17029_), .B(new_n17026_), .S0(new_n11767_), .Y(new_n17030_));
  NOR2X1   g14594(.A(new_n17030_), .B(pi0789), .Y(new_n17031_));
  AOI21X1  g14595(.A0(new_n17030_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n17032_));
  AOI21X1  g14596(.A0(new_n17030_), .A1(new_n15790_), .B0(pi1159), .Y(new_n17033_));
  OR2X1    g14597(.A(new_n17033_), .B(new_n17032_), .Y(new_n17034_));
  AOI21X1  g14598(.A0(new_n17034_), .A1(pi0789), .B0(new_n17031_), .Y(new_n17035_));
  INVX1    g14599(.A(new_n17035_), .Y(new_n17036_));
  MX2X1    g14600(.A(new_n17036_), .B(new_n17017_), .S0(new_n12708_), .Y(new_n17037_));
  MX2X1    g14601(.A(new_n17037_), .B(new_n17017_), .S0(new_n12580_), .Y(new_n17038_));
  AOI21X1  g14602(.A0(new_n12439_), .A1(new_n14997_), .B0(new_n17016_), .Y(new_n17039_));
  OR2X1    g14603(.A(new_n17039_), .B(pi0778), .Y(new_n17040_));
  INVX1    g14604(.A(new_n17039_), .Y(new_n17041_));
  AND3X1   g14605(.A(new_n12439_), .B(new_n14997_), .C(new_n12363_), .Y(new_n17042_));
  INVX1    g14606(.A(new_n17042_), .Y(new_n17043_));
  AOI21X1  g14607(.A0(new_n17043_), .A1(new_n17041_), .B0(new_n12364_), .Y(new_n17044_));
  NOR3X1   g14608(.A(new_n17042_), .B(new_n17016_), .C(pi1153), .Y(new_n17045_));
  OR3X1    g14609(.A(new_n17045_), .B(new_n17044_), .C(new_n11769_), .Y(new_n17046_));
  AND2X1   g14610(.A(new_n17046_), .B(new_n17040_), .Y(new_n17047_));
  NOR4X1   g14611(.A(new_n17047_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n17048_));
  AND3X1   g14612(.A(new_n17048_), .B(new_n12739_), .C(new_n12718_), .Y(new_n17049_));
  INVX1    g14613(.A(new_n17049_), .Y(new_n17050_));
  AOI21X1  g14614(.A0(new_n17016_), .A1(pi0647), .B0(pi1157), .Y(new_n17051_));
  OAI21X1  g14615(.A0(new_n17050_), .A1(pi0647), .B0(new_n17051_), .Y(new_n17052_));
  MX2X1    g14616(.A(new_n17049_), .B(new_n17016_), .S0(new_n12577_), .Y(new_n17053_));
  OAI22X1  g14617(.A0(new_n17053_), .A1(new_n14242_), .B0(new_n17052_), .B1(new_n12592_), .Y(new_n17054_));
  AOI21X1  g14618(.A0(new_n17038_), .A1(new_n14326_), .B0(new_n17054_), .Y(new_n17055_));
  NOR2X1   g14619(.A(new_n17055_), .B(new_n11763_), .Y(new_n17056_));
  AOI21X1  g14620(.A0(new_n17017_), .A1(pi0626), .B0(new_n16218_), .Y(new_n17057_));
  OAI21X1  g14621(.A0(new_n17035_), .A1(pi0626), .B0(new_n17057_), .Y(new_n17058_));
  AOI21X1  g14622(.A0(new_n17017_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n17059_));
  OAI21X1  g14623(.A0(new_n17035_), .A1(new_n12542_), .B0(new_n17059_), .Y(new_n17060_));
  NAND2X1  g14624(.A(new_n17048_), .B(new_n12637_), .Y(new_n17061_));
  AND3X1   g14625(.A(new_n17061_), .B(new_n17060_), .C(new_n17058_), .Y(new_n17062_));
  NOR2X1   g14626(.A(new_n17062_), .B(new_n11765_), .Y(new_n17063_));
  NOR2X1   g14627(.A(new_n17016_), .B(pi1153), .Y(new_n17064_));
  NOR3X1   g14628(.A(new_n17039_), .B(new_n11991_), .C(new_n12363_), .Y(new_n17065_));
  AOI21X1  g14629(.A0(new_n17041_), .A1(new_n12048_), .B0(new_n17019_), .Y(new_n17066_));
  OAI21X1  g14630(.A0(new_n17066_), .A1(new_n17065_), .B0(new_n17064_), .Y(new_n17067_));
  NOR2X1   g14631(.A(new_n17044_), .B(pi0608), .Y(new_n17068_));
  NOR3X1   g14632(.A(new_n17065_), .B(new_n17019_), .C(new_n12364_), .Y(new_n17069_));
  NOR3X1   g14633(.A(new_n17069_), .B(new_n17045_), .C(new_n12368_), .Y(new_n17070_));
  AOI21X1  g14634(.A0(new_n17068_), .A1(new_n17067_), .B0(new_n17070_), .Y(new_n17071_));
  OR2X1    g14635(.A(new_n17066_), .B(pi0778), .Y(new_n17072_));
  OAI21X1  g14636(.A0(new_n17071_), .A1(new_n11769_), .B0(new_n17072_), .Y(new_n17073_));
  INVX1    g14637(.A(new_n17073_), .Y(new_n17074_));
  AND2X1   g14638(.A(new_n17073_), .B(new_n12462_), .Y(new_n17075_));
  OAI21X1  g14639(.A0(new_n17047_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n17076_));
  OR2X1    g14640(.A(new_n17076_), .B(new_n17075_), .Y(new_n17077_));
  AND3X1   g14641(.A(new_n17077_), .B(new_n17022_), .C(new_n12468_), .Y(new_n17078_));
  OAI21X1  g14642(.A0(new_n17047_), .A1(pi0609), .B0(pi1155), .Y(new_n17079_));
  AOI21X1  g14643(.A0(new_n17073_), .A1(pi0609), .B0(new_n17079_), .Y(new_n17080_));
  NOR3X1   g14644(.A(new_n17080_), .B(new_n17023_), .C(new_n12468_), .Y(new_n17081_));
  NOR2X1   g14645(.A(new_n17081_), .B(new_n17078_), .Y(new_n17082_));
  MX2X1    g14646(.A(new_n17082_), .B(new_n17074_), .S0(new_n11768_), .Y(new_n17083_));
  AOI21X1  g14647(.A0(new_n17046_), .A1(new_n17040_), .B0(new_n12630_), .Y(new_n17084_));
  AOI21X1  g14648(.A0(new_n17084_), .A1(pi0618), .B0(pi1154), .Y(new_n17085_));
  OAI21X1  g14649(.A0(new_n17083_), .A1(pi0618), .B0(new_n17085_), .Y(new_n17086_));
  NOR2X1   g14650(.A(new_n17027_), .B(pi0627), .Y(new_n17087_));
  AOI21X1  g14651(.A0(new_n17084_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17088_));
  OAI21X1  g14652(.A0(new_n17083_), .A1(new_n12486_), .B0(new_n17088_), .Y(new_n17089_));
  NOR2X1   g14653(.A(new_n17028_), .B(new_n12494_), .Y(new_n17090_));
  AOI22X1  g14654(.A0(new_n17090_), .A1(new_n17089_), .B0(new_n17087_), .B1(new_n17086_), .Y(new_n17091_));
  MX2X1    g14655(.A(new_n17091_), .B(new_n17083_), .S0(new_n11767_), .Y(new_n17092_));
  OR4X1    g14656(.A(new_n17047_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n17093_));
  AND2X1   g14657(.A(new_n17093_), .B(new_n12510_), .Y(new_n17094_));
  OAI21X1  g14658(.A0(new_n17092_), .A1(pi0619), .B0(new_n17094_), .Y(new_n17095_));
  NOR2X1   g14659(.A(new_n17032_), .B(pi0648), .Y(new_n17096_));
  AND2X1   g14660(.A(new_n17096_), .B(new_n17095_), .Y(new_n17097_));
  NOR4X1   g14661(.A(new_n17047_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n17098_));
  NOR2X1   g14662(.A(new_n17098_), .B(new_n12510_), .Y(new_n17099_));
  OAI21X1  g14663(.A0(new_n17092_), .A1(new_n12509_), .B0(new_n17099_), .Y(new_n17100_));
  NOR2X1   g14664(.A(new_n17033_), .B(new_n12517_), .Y(new_n17101_));
  AND2X1   g14665(.A(new_n17101_), .B(new_n17100_), .Y(new_n17102_));
  OR3X1    g14666(.A(new_n17102_), .B(new_n17097_), .C(new_n11766_), .Y(new_n17103_));
  AOI21X1  g14667(.A0(new_n17092_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n17104_));
  AOI21X1  g14668(.A0(new_n17104_), .A1(new_n17103_), .B0(new_n17063_), .Y(new_n17105_));
  OR2X1    g14669(.A(new_n17105_), .B(new_n14125_), .Y(new_n17106_));
  INVX1    g14670(.A(new_n17037_), .Y(new_n17107_));
  AND2X1   g14671(.A(new_n17048_), .B(new_n12718_), .Y(new_n17108_));
  AOI22X1  g14672(.A0(new_n17108_), .A1(new_n14426_), .B0(new_n17107_), .B1(new_n12735_), .Y(new_n17109_));
  AOI22X1  g14673(.A0(new_n17108_), .A1(new_n14428_), .B0(new_n17107_), .B1(new_n12733_), .Y(new_n17110_));
  MX2X1    g14674(.A(new_n17110_), .B(new_n17109_), .S0(new_n12561_), .Y(new_n17111_));
  OAI21X1  g14675(.A0(new_n17111_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n17112_));
  INVX1    g14676(.A(new_n17112_), .Y(new_n17113_));
  AOI21X1  g14677(.A0(new_n17113_), .A1(new_n17106_), .B0(new_n17056_), .Y(new_n17114_));
  OAI21X1  g14678(.A0(new_n17053_), .A1(new_n12578_), .B0(new_n17052_), .Y(new_n17115_));
  MX2X1    g14679(.A(new_n17115_), .B(new_n17050_), .S0(new_n11763_), .Y(new_n17116_));
  OAI21X1  g14680(.A0(new_n17116_), .A1(pi0644), .B0(pi0715), .Y(new_n17117_));
  AOI21X1  g14681(.A0(new_n17114_), .A1(pi0644), .B0(new_n17117_), .Y(new_n17118_));
  OR3X1    g14682(.A(new_n17017_), .B(new_n12603_), .C(new_n11763_), .Y(new_n17119_));
  OAI21X1  g14683(.A0(new_n17038_), .A1(new_n12604_), .B0(new_n17119_), .Y(new_n17120_));
  OAI21X1  g14684(.A0(new_n17017_), .A1(pi0644), .B0(new_n12608_), .Y(new_n17121_));
  AOI21X1  g14685(.A0(new_n17120_), .A1(pi0644), .B0(new_n17121_), .Y(new_n17122_));
  OR2X1    g14686(.A(new_n17122_), .B(new_n11762_), .Y(new_n17123_));
  OAI21X1  g14687(.A0(new_n17116_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17124_));
  AOI21X1  g14688(.A0(new_n17114_), .A1(new_n12612_), .B0(new_n17124_), .Y(new_n17125_));
  OAI21X1  g14689(.A0(new_n17017_), .A1(new_n12612_), .B0(pi0715), .Y(new_n17126_));
  AOI21X1  g14690(.A0(new_n17120_), .A1(new_n12612_), .B0(new_n17126_), .Y(new_n17127_));
  OR2X1    g14691(.A(new_n17127_), .B(pi1160), .Y(new_n17128_));
  OAI22X1  g14692(.A0(new_n17128_), .A1(new_n17125_), .B0(new_n17123_), .B1(new_n17118_), .Y(new_n17129_));
  NAND2X1  g14693(.A(new_n17129_), .B(pi0790), .Y(new_n17130_));
  AOI21X1  g14694(.A0(new_n17114_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n17131_));
  AOI21X1  g14695(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0178), .Y(new_n17132_));
  INVX1    g14696(.A(new_n17132_), .Y(new_n17133_));
  AOI21X1  g14697(.A0(new_n3103_), .A1(new_n14997_), .B0(new_n17133_), .Y(new_n17134_));
  OAI21X1  g14698(.A0(new_n12826_), .A1(new_n6801_), .B0(new_n2979_), .Y(new_n17135_));
  AOI22X1  g14699(.A0(new_n17135_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n6801_), .Y(new_n17136_));
  AOI21X1  g14700(.A0(new_n12771_), .A1(new_n6801_), .B0(new_n12441_), .Y(new_n17137_));
  NOR3X1   g14701(.A(new_n17137_), .B(new_n17136_), .C(pi0688), .Y(new_n17138_));
  NOR2X1   g14702(.A(new_n17138_), .B(new_n17134_), .Y(new_n17139_));
  INVX1    g14703(.A(new_n17139_), .Y(new_n17140_));
  AOI21X1  g14704(.A0(new_n17132_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n17141_));
  OAI21X1  g14705(.A0(new_n17139_), .A1(new_n12363_), .B0(new_n17141_), .Y(new_n17142_));
  AOI21X1  g14706(.A0(new_n17132_), .A1(pi0625), .B0(pi1153), .Y(new_n17143_));
  OAI21X1  g14707(.A0(new_n17139_), .A1(pi0625), .B0(new_n17143_), .Y(new_n17144_));
  AND2X1   g14708(.A(new_n17144_), .B(new_n17142_), .Y(new_n17145_));
  MX2X1    g14709(.A(new_n17145_), .B(new_n17140_), .S0(new_n11769_), .Y(new_n17146_));
  MX2X1    g14710(.A(new_n17146_), .B(new_n17132_), .S0(new_n12490_), .Y(new_n17147_));
  INVX1    g14711(.A(new_n17147_), .Y(new_n17148_));
  MX2X1    g14712(.A(new_n17148_), .B(new_n17133_), .S0(new_n12513_), .Y(new_n17149_));
  INVX1    g14713(.A(new_n17149_), .Y(new_n17150_));
  MX2X1    g14714(.A(new_n17150_), .B(new_n17132_), .S0(new_n12531_), .Y(new_n17151_));
  MX2X1    g14715(.A(new_n17151_), .B(new_n17132_), .S0(new_n12563_), .Y(new_n17152_));
  INVX1    g14716(.A(new_n17152_), .Y(new_n17153_));
  AOI21X1  g14717(.A0(new_n17132_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n17154_));
  OAI21X1  g14718(.A0(new_n17153_), .A1(new_n12554_), .B0(new_n17154_), .Y(new_n17155_));
  AOI21X1  g14719(.A0(new_n17132_), .A1(pi0628), .B0(pi1156), .Y(new_n17156_));
  OAI21X1  g14720(.A0(new_n17153_), .A1(pi0628), .B0(new_n17156_), .Y(new_n17157_));
  AOI21X1  g14721(.A0(new_n17157_), .A1(new_n17155_), .B0(new_n11764_), .Y(new_n17158_));
  AOI21X1  g14722(.A0(new_n17153_), .A1(new_n11764_), .B0(new_n17158_), .Y(new_n17159_));
  MX2X1    g14723(.A(new_n17159_), .B(new_n17132_), .S0(pi0647), .Y(new_n17160_));
  MX2X1    g14724(.A(new_n17159_), .B(new_n17132_), .S0(new_n12577_), .Y(new_n17161_));
  MX2X1    g14725(.A(new_n17161_), .B(new_n17160_), .S0(new_n12578_), .Y(new_n17162_));
  MX2X1    g14726(.A(new_n17162_), .B(new_n17159_), .S0(new_n11763_), .Y(new_n17163_));
  AOI21X1  g14727(.A0(new_n17163_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17164_));
  OAI22X1  g14728(.A0(new_n14197_), .A1(pi0760), .B0(new_n12077_), .B1(pi0178), .Y(new_n17165_));
  AOI21X1  g14729(.A0(new_n16615_), .A1(pi0178), .B0(pi0760), .Y(new_n17166_));
  OAI21X1  g14730(.A0(new_n12776_), .A1(pi0178), .B0(new_n17166_), .Y(new_n17167_));
  OR3X1    g14731(.A(new_n12445_), .B(new_n14970_), .C(pi0178), .Y(new_n17168_));
  AOI21X1  g14732(.A0(new_n17168_), .A1(new_n17167_), .B0(pi0038), .Y(new_n17169_));
  AOI21X1  g14733(.A0(new_n17165_), .A1(pi0038), .B0(new_n17169_), .Y(new_n17170_));
  MX2X1    g14734(.A(new_n17170_), .B(pi0178), .S0(new_n11770_), .Y(new_n17171_));
  AND2X1   g14735(.A(new_n17171_), .B(new_n12474_), .Y(new_n17172_));
  AOI21X1  g14736(.A0(new_n17133_), .A1(new_n12473_), .B0(new_n17172_), .Y(new_n17173_));
  AOI22X1  g14737(.A0(new_n17172_), .A1(pi0609), .B0(new_n17133_), .B1(new_n12472_), .Y(new_n17174_));
  AOI22X1  g14738(.A0(new_n17172_), .A1(new_n12462_), .B0(new_n17133_), .B1(new_n12481_), .Y(new_n17175_));
  MX2X1    g14739(.A(new_n17175_), .B(new_n17174_), .S0(pi1155), .Y(new_n17176_));
  MX2X1    g14740(.A(new_n17176_), .B(new_n17173_), .S0(new_n11768_), .Y(new_n17177_));
  OAI21X1  g14741(.A0(new_n17133_), .A1(pi0618), .B0(pi1154), .Y(new_n17178_));
  AOI21X1  g14742(.A0(new_n17177_), .A1(pi0618), .B0(new_n17178_), .Y(new_n17179_));
  OAI21X1  g14743(.A0(new_n17133_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17180_));
  AOI21X1  g14744(.A0(new_n17177_), .A1(new_n12486_), .B0(new_n17180_), .Y(new_n17181_));
  NOR2X1   g14745(.A(new_n17181_), .B(new_n17179_), .Y(new_n17182_));
  MX2X1    g14746(.A(new_n17182_), .B(new_n17177_), .S0(new_n11767_), .Y(new_n17183_));
  OAI21X1  g14747(.A0(new_n17133_), .A1(pi0619), .B0(pi1159), .Y(new_n17184_));
  AOI21X1  g14748(.A0(new_n17183_), .A1(pi0619), .B0(new_n17184_), .Y(new_n17185_));
  OAI21X1  g14749(.A0(new_n17133_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n17186_));
  AOI21X1  g14750(.A0(new_n17183_), .A1(new_n12509_), .B0(new_n17186_), .Y(new_n17187_));
  NOR2X1   g14751(.A(new_n17187_), .B(new_n17185_), .Y(new_n17188_));
  MX2X1    g14752(.A(new_n17188_), .B(new_n17183_), .S0(new_n11766_), .Y(new_n17189_));
  AND2X1   g14753(.A(new_n17132_), .B(new_n12708_), .Y(new_n17190_));
  AOI21X1  g14754(.A0(new_n17189_), .A1(new_n16140_), .B0(new_n17190_), .Y(new_n17191_));
  NAND2X1  g14755(.A(new_n17132_), .B(new_n12580_), .Y(new_n17192_));
  OAI21X1  g14756(.A0(new_n17191_), .A1(new_n12580_), .B0(new_n17192_), .Y(new_n17193_));
  MX2X1    g14757(.A(new_n17193_), .B(new_n17132_), .S0(new_n12604_), .Y(new_n17194_));
  OAI21X1  g14758(.A0(new_n17133_), .A1(pi0644), .B0(new_n12608_), .Y(new_n17195_));
  AOI21X1  g14759(.A0(new_n17194_), .A1(pi0644), .B0(new_n17195_), .Y(new_n17196_));
  OR2X1    g14760(.A(new_n17196_), .B(new_n11762_), .Y(new_n17197_));
  AOI21X1  g14761(.A0(new_n17163_), .A1(pi0644), .B0(pi0715), .Y(new_n17198_));
  OAI21X1  g14762(.A0(new_n17133_), .A1(new_n12612_), .B0(pi0715), .Y(new_n17199_));
  AOI21X1  g14763(.A0(new_n17194_), .A1(new_n12612_), .B0(new_n17199_), .Y(new_n17200_));
  OR2X1    g14764(.A(new_n17200_), .B(pi1160), .Y(new_n17201_));
  OAI22X1  g14765(.A0(new_n17201_), .A1(new_n17198_), .B0(new_n17197_), .B1(new_n17164_), .Y(new_n17202_));
  OR3X1    g14766(.A(new_n17200_), .B(pi1160), .C(pi0644), .Y(new_n17203_));
  OR3X1    g14767(.A(new_n17196_), .B(new_n11762_), .C(new_n12612_), .Y(new_n17204_));
  NAND3X1  g14768(.A(new_n17204_), .B(new_n17203_), .C(pi0790), .Y(new_n17205_));
  NAND2X1  g14769(.A(new_n17191_), .B(new_n14249_), .Y(new_n17206_));
  MX2X1    g14770(.A(new_n17157_), .B(new_n17155_), .S0(new_n12561_), .Y(new_n17207_));
  AND2X1   g14771(.A(new_n17207_), .B(new_n17206_), .Y(new_n17208_));
  OR2X1    g14772(.A(new_n17208_), .B(new_n11764_), .Y(new_n17209_));
  OR2X1    g14773(.A(new_n17170_), .B(new_n14997_), .Y(new_n17210_));
  OAI21X1  g14774(.A0(new_n12213_), .A1(new_n6801_), .B0(pi0760), .Y(new_n17211_));
  AOI21X1  g14775(.A0(new_n12155_), .A1(new_n6801_), .B0(new_n17211_), .Y(new_n17212_));
  AOI21X1  g14776(.A0(new_n12788_), .A1(new_n6801_), .B0(pi0760), .Y(new_n17213_));
  OAI21X1  g14777(.A0(new_n12787_), .A1(new_n6801_), .B0(new_n17213_), .Y(new_n17214_));
  NAND2X1  g14778(.A(new_n17214_), .B(pi0039), .Y(new_n17215_));
  AND2X1   g14779(.A(new_n12332_), .B(pi0178), .Y(new_n17216_));
  OAI21X1  g14780(.A0(new_n12315_), .A1(pi0178), .B0(pi0760), .Y(new_n17217_));
  NOR4X1   g14781(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0178), .Y(new_n17218_));
  OAI21X1  g14782(.A0(new_n12800_), .A1(new_n6801_), .B0(new_n14970_), .Y(new_n17219_));
  OAI22X1  g14783(.A0(new_n17219_), .A1(new_n17218_), .B0(new_n17217_), .B1(new_n17216_), .Y(new_n17220_));
  AOI21X1  g14784(.A0(new_n17220_), .A1(new_n2939_), .B0(pi0038), .Y(new_n17221_));
  OAI21X1  g14785(.A0(new_n17215_), .A1(new_n17212_), .B0(new_n17221_), .Y(new_n17222_));
  OAI21X1  g14786(.A0(new_n12276_), .A1(pi0760), .B0(new_n13540_), .Y(new_n17223_));
  NAND2X1  g14787(.A(new_n17223_), .B(new_n6801_), .Y(new_n17224_));
  AOI21X1  g14788(.A0(new_n12056_), .A1(new_n14970_), .B0(new_n13443_), .Y(new_n17225_));
  NOR2X1   g14789(.A(new_n17225_), .B(new_n6801_), .Y(new_n17226_));
  AOI21X1  g14790(.A0(new_n17226_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n17227_));
  AOI21X1  g14791(.A0(new_n17227_), .A1(new_n17224_), .B0(pi0688), .Y(new_n17228_));
  AOI21X1  g14792(.A0(new_n17228_), .A1(new_n17222_), .B0(new_n11770_), .Y(new_n17229_));
  AOI22X1  g14793(.A0(new_n17229_), .A1(new_n17210_), .B0(new_n11770_), .B1(pi0178), .Y(new_n17230_));
  OAI21X1  g14794(.A0(new_n17171_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n17231_));
  AOI21X1  g14795(.A0(new_n17230_), .A1(new_n12363_), .B0(new_n17231_), .Y(new_n17232_));
  NAND2X1  g14796(.A(new_n17142_), .B(new_n12368_), .Y(new_n17233_));
  OAI21X1  g14797(.A0(new_n17171_), .A1(pi0625), .B0(pi1153), .Y(new_n17234_));
  AOI21X1  g14798(.A0(new_n17230_), .A1(pi0625), .B0(new_n17234_), .Y(new_n17235_));
  NAND2X1  g14799(.A(new_n17144_), .B(pi0608), .Y(new_n17236_));
  OAI22X1  g14800(.A0(new_n17236_), .A1(new_n17235_), .B0(new_n17233_), .B1(new_n17232_), .Y(new_n17237_));
  MX2X1    g14801(.A(new_n17237_), .B(new_n17230_), .S0(new_n11769_), .Y(new_n17238_));
  INVX1    g14802(.A(new_n17146_), .Y(new_n17239_));
  OAI21X1  g14803(.A0(new_n17239_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n17240_));
  AOI21X1  g14804(.A0(new_n17238_), .A1(new_n12462_), .B0(new_n17240_), .Y(new_n17241_));
  OAI21X1  g14805(.A0(new_n17174_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n17242_));
  OAI21X1  g14806(.A0(new_n17239_), .A1(pi0609), .B0(pi1155), .Y(new_n17243_));
  AOI21X1  g14807(.A0(new_n17238_), .A1(pi0609), .B0(new_n17243_), .Y(new_n17244_));
  OAI21X1  g14808(.A0(new_n17175_), .A1(pi1155), .B0(pi0660), .Y(new_n17245_));
  OAI22X1  g14809(.A0(new_n17245_), .A1(new_n17244_), .B0(new_n17242_), .B1(new_n17241_), .Y(new_n17246_));
  MX2X1    g14810(.A(new_n17246_), .B(new_n17238_), .S0(new_n11768_), .Y(new_n17247_));
  OAI21X1  g14811(.A0(new_n17148_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17248_));
  AOI21X1  g14812(.A0(new_n17247_), .A1(new_n12486_), .B0(new_n17248_), .Y(new_n17249_));
  OR2X1    g14813(.A(new_n17179_), .B(pi0627), .Y(new_n17250_));
  OAI21X1  g14814(.A0(new_n17148_), .A1(pi0618), .B0(pi1154), .Y(new_n17251_));
  AOI21X1  g14815(.A0(new_n17247_), .A1(pi0618), .B0(new_n17251_), .Y(new_n17252_));
  OR2X1    g14816(.A(new_n17181_), .B(new_n12494_), .Y(new_n17253_));
  OAI22X1  g14817(.A0(new_n17253_), .A1(new_n17252_), .B0(new_n17250_), .B1(new_n17249_), .Y(new_n17254_));
  MX2X1    g14818(.A(new_n17254_), .B(new_n17247_), .S0(new_n11767_), .Y(new_n17255_));
  NAND2X1  g14819(.A(new_n17255_), .B(new_n12509_), .Y(new_n17256_));
  AOI21X1  g14820(.A0(new_n17150_), .A1(pi0619), .B0(pi1159), .Y(new_n17257_));
  OR2X1    g14821(.A(new_n17185_), .B(pi0648), .Y(new_n17258_));
  AOI21X1  g14822(.A0(new_n17257_), .A1(new_n17256_), .B0(new_n17258_), .Y(new_n17259_));
  NAND2X1  g14823(.A(new_n17255_), .B(pi0619), .Y(new_n17260_));
  AOI21X1  g14824(.A0(new_n17150_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n17261_));
  OR2X1    g14825(.A(new_n17187_), .B(new_n12517_), .Y(new_n17262_));
  AOI21X1  g14826(.A0(new_n17261_), .A1(new_n17260_), .B0(new_n17262_), .Y(new_n17263_));
  NOR3X1   g14827(.A(new_n17263_), .B(new_n17259_), .C(new_n11766_), .Y(new_n17264_));
  OAI21X1  g14828(.A0(new_n17255_), .A1(pi0789), .B0(new_n12709_), .Y(new_n17265_));
  AOI21X1  g14829(.A0(new_n17133_), .A1(pi0626), .B0(new_n16218_), .Y(new_n17266_));
  OAI21X1  g14830(.A0(new_n17189_), .A1(pi0626), .B0(new_n17266_), .Y(new_n17267_));
  AOI21X1  g14831(.A0(new_n17133_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n17268_));
  OAI21X1  g14832(.A0(new_n17189_), .A1(new_n12542_), .B0(new_n17268_), .Y(new_n17269_));
  NAND2X1  g14833(.A(new_n17151_), .B(new_n12637_), .Y(new_n17270_));
  NAND3X1  g14834(.A(new_n17270_), .B(new_n17269_), .C(new_n17267_), .Y(new_n17271_));
  AOI21X1  g14835(.A0(new_n17271_), .A1(pi0788), .B0(new_n14125_), .Y(new_n17272_));
  OAI21X1  g14836(.A0(new_n17265_), .A1(new_n17264_), .B0(new_n17272_), .Y(new_n17273_));
  AOI21X1  g14837(.A0(new_n17273_), .A1(new_n17209_), .B0(new_n14121_), .Y(new_n17274_));
  OR2X1    g14838(.A(new_n17193_), .B(new_n14239_), .Y(new_n17275_));
  OR2X1    g14839(.A(new_n17160_), .B(new_n14244_), .Y(new_n17276_));
  OR2X1    g14840(.A(new_n17161_), .B(new_n14242_), .Y(new_n17277_));
  NAND3X1  g14841(.A(new_n17277_), .B(new_n17276_), .C(new_n17275_), .Y(new_n17278_));
  AOI21X1  g14842(.A0(new_n17278_), .A1(pi0787), .B0(new_n17274_), .Y(new_n17279_));
  AOI22X1  g14843(.A0(new_n17279_), .A1(new_n17205_), .B0(new_n17202_), .B1(pi0790), .Y(new_n17280_));
  OR2X1    g14844(.A(new_n17280_), .B(po1038), .Y(new_n17281_));
  AOI21X1  g14845(.A0(po1038), .A1(new_n6801_), .B0(pi0832), .Y(new_n17282_));
  AOI22X1  g14846(.A0(new_n17282_), .A1(new_n17281_), .B0(new_n17131_), .B1(new_n17130_), .Y(po0335));
  OAI21X1  g14847(.A0(new_n12077_), .A1(pi0179), .B0(new_n12806_), .Y(new_n17284_));
  INVX1    g14848(.A(pi0179), .Y(new_n17285_));
  OAI21X1  g14849(.A0(new_n12213_), .A1(new_n17285_), .B0(pi0039), .Y(new_n17286_));
  AOI21X1  g14850(.A0(new_n12155_), .A1(new_n17285_), .B0(new_n17286_), .Y(new_n17287_));
  OAI21X1  g14851(.A0(new_n12332_), .A1(new_n17285_), .B0(new_n2939_), .Y(new_n17288_));
  AOI21X1  g14852(.A0(new_n12315_), .A1(new_n17285_), .B0(new_n17288_), .Y(new_n17289_));
  OAI21X1  g14853(.A0(new_n17289_), .A1(new_n17287_), .B0(new_n2979_), .Y(new_n17290_));
  AOI21X1  g14854(.A0(new_n17290_), .A1(new_n17284_), .B0(new_n14955_), .Y(new_n17291_));
  OAI21X1  g14855(.A0(new_n13559_), .A1(pi0179), .B0(new_n14955_), .Y(new_n17292_));
  AOI21X1  g14856(.A0(new_n13554_), .A1(pi0179), .B0(new_n17292_), .Y(new_n17293_));
  OR3X1    g14857(.A(new_n17293_), .B(new_n17291_), .C(pi0724), .Y(new_n17294_));
  AOI21X1  g14858(.A0(new_n16617_), .A1(new_n14955_), .B0(new_n17285_), .Y(new_n17295_));
  NOR3X1   g14859(.A(new_n13565_), .B(pi0741), .C(pi0179), .Y(new_n17296_));
  AND2X1   g14860(.A(new_n17296_), .B(new_n13568_), .Y(new_n17297_));
  OR2X1    g14861(.A(new_n17297_), .B(new_n17295_), .Y(new_n17298_));
  AOI21X1  g14862(.A0(new_n12447_), .A1(pi0741), .B0(new_n17298_), .Y(new_n17299_));
  AOI21X1  g14863(.A0(new_n17299_), .A1(pi0724), .B0(new_n11770_), .Y(new_n17300_));
  AOI22X1  g14864(.A0(new_n17300_), .A1(new_n17294_), .B0(new_n11770_), .B1(pi0179), .Y(new_n17301_));
  OR2X1    g14865(.A(new_n3103_), .B(new_n17285_), .Y(new_n17302_));
  OAI21X1  g14866(.A0(new_n17299_), .A1(new_n11770_), .B0(new_n17302_), .Y(new_n17303_));
  OAI21X1  g14867(.A0(new_n17303_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n17304_));
  AOI21X1  g14868(.A0(new_n17301_), .A1(new_n12363_), .B0(new_n17304_), .Y(new_n17305_));
  AOI21X1  g14869(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0179), .Y(new_n17306_));
  OAI21X1  g14870(.A0(new_n11770_), .A1(pi0724), .B0(new_n17306_), .Y(new_n17307_));
  OAI21X1  g14871(.A0(new_n12826_), .A1(new_n17285_), .B0(new_n2979_), .Y(new_n17308_));
  AOI22X1  g14872(.A0(new_n17308_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n17285_), .Y(new_n17309_));
  AOI21X1  g14873(.A0(new_n12771_), .A1(new_n17285_), .B0(new_n12441_), .Y(new_n17310_));
  OR3X1    g14874(.A(new_n17310_), .B(new_n17309_), .C(pi0724), .Y(new_n17311_));
  AOI21X1  g14875(.A0(new_n17311_), .A1(new_n17307_), .B0(new_n12363_), .Y(new_n17312_));
  OAI21X1  g14876(.A0(new_n12832_), .A1(new_n11770_), .B0(new_n17285_), .Y(new_n17313_));
  OAI21X1  g14877(.A0(new_n17313_), .A1(pi0625), .B0(pi1153), .Y(new_n17314_));
  OAI21X1  g14878(.A0(new_n17314_), .A1(new_n17312_), .B0(new_n12368_), .Y(new_n17315_));
  OAI21X1  g14879(.A0(new_n17303_), .A1(pi0625), .B0(pi1153), .Y(new_n17316_));
  AOI21X1  g14880(.A0(new_n17301_), .A1(pi0625), .B0(new_n17316_), .Y(new_n17317_));
  AOI21X1  g14881(.A0(new_n17311_), .A1(new_n17307_), .B0(pi0625), .Y(new_n17318_));
  OAI21X1  g14882(.A0(new_n17313_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n17319_));
  OAI21X1  g14883(.A0(new_n17319_), .A1(new_n17318_), .B0(pi0608), .Y(new_n17320_));
  OAI22X1  g14884(.A0(new_n17320_), .A1(new_n17317_), .B0(new_n17315_), .B1(new_n17305_), .Y(new_n17321_));
  AND2X1   g14885(.A(new_n17301_), .B(new_n11769_), .Y(new_n17322_));
  AOI21X1  g14886(.A0(new_n17321_), .A1(pi0778), .B0(new_n17322_), .Y(new_n17323_));
  NOR2X1   g14887(.A(new_n17323_), .B(pi0609), .Y(new_n17324_));
  AND2X1   g14888(.A(new_n17311_), .B(new_n17307_), .Y(new_n17325_));
  OAI22X1  g14889(.A0(new_n17319_), .A1(new_n17318_), .B0(new_n17314_), .B1(new_n17312_), .Y(new_n17326_));
  MX2X1    g14890(.A(new_n17326_), .B(new_n17325_), .S0(new_n11769_), .Y(new_n17327_));
  OAI21X1  g14891(.A0(new_n17327_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n17328_));
  AND2X1   g14892(.A(new_n17303_), .B(new_n12474_), .Y(new_n17329_));
  AOI22X1  g14893(.A0(new_n17329_), .A1(pi0609), .B0(new_n17313_), .B1(new_n12472_), .Y(new_n17330_));
  OR2X1    g14894(.A(new_n17330_), .B(new_n12463_), .Y(new_n17331_));
  AND2X1   g14895(.A(new_n17331_), .B(new_n12468_), .Y(new_n17332_));
  OAI21X1  g14896(.A0(new_n17328_), .A1(new_n17324_), .B0(new_n17332_), .Y(new_n17333_));
  NOR2X1   g14897(.A(new_n17323_), .B(new_n12462_), .Y(new_n17334_));
  OAI21X1  g14898(.A0(new_n17327_), .A1(pi0609), .B0(pi1155), .Y(new_n17335_));
  AOI22X1  g14899(.A0(new_n17329_), .A1(new_n12462_), .B0(new_n17313_), .B1(new_n12481_), .Y(new_n17336_));
  OR2X1    g14900(.A(new_n17336_), .B(pi1155), .Y(new_n17337_));
  AND2X1   g14901(.A(new_n17337_), .B(pi0660), .Y(new_n17338_));
  OAI21X1  g14902(.A0(new_n17335_), .A1(new_n17334_), .B0(new_n17338_), .Y(new_n17339_));
  AND2X1   g14903(.A(new_n17339_), .B(new_n17333_), .Y(new_n17340_));
  MX2X1    g14904(.A(new_n17340_), .B(new_n17323_), .S0(new_n11768_), .Y(new_n17341_));
  MX2X1    g14905(.A(new_n17327_), .B(new_n17313_), .S0(new_n12490_), .Y(new_n17342_));
  INVX1    g14906(.A(new_n17342_), .Y(new_n17343_));
  AOI21X1  g14907(.A0(new_n17343_), .A1(pi0618), .B0(pi1154), .Y(new_n17344_));
  OAI21X1  g14908(.A0(new_n17341_), .A1(pi0618), .B0(new_n17344_), .Y(new_n17345_));
  AOI21X1  g14909(.A0(new_n17313_), .A1(new_n12473_), .B0(new_n17329_), .Y(new_n17346_));
  MX2X1    g14910(.A(new_n17336_), .B(new_n17330_), .S0(pi1155), .Y(new_n17347_));
  MX2X1    g14911(.A(new_n17347_), .B(new_n17346_), .S0(new_n11768_), .Y(new_n17348_));
  OAI21X1  g14912(.A0(new_n17313_), .A1(pi0618), .B0(pi1154), .Y(new_n17349_));
  AOI21X1  g14913(.A0(new_n17348_), .A1(pi0618), .B0(new_n17349_), .Y(new_n17350_));
  NOR2X1   g14914(.A(new_n17350_), .B(pi0627), .Y(new_n17351_));
  AOI21X1  g14915(.A0(new_n17343_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17352_));
  OAI21X1  g14916(.A0(new_n17341_), .A1(new_n12486_), .B0(new_n17352_), .Y(new_n17353_));
  OAI21X1  g14917(.A0(new_n17313_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17354_));
  AOI21X1  g14918(.A0(new_n17348_), .A1(new_n12486_), .B0(new_n17354_), .Y(new_n17355_));
  NOR2X1   g14919(.A(new_n17355_), .B(new_n12494_), .Y(new_n17356_));
  AOI22X1  g14920(.A0(new_n17356_), .A1(new_n17353_), .B0(new_n17351_), .B1(new_n17345_), .Y(new_n17357_));
  OR2X1    g14921(.A(new_n17341_), .B(pi0781), .Y(new_n17358_));
  OAI21X1  g14922(.A0(new_n17357_), .A1(new_n11767_), .B0(new_n17358_), .Y(new_n17359_));
  MX2X1    g14923(.A(new_n17342_), .B(new_n17313_), .S0(new_n12513_), .Y(new_n17360_));
  OAI21X1  g14924(.A0(new_n17360_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n17361_));
  AOI21X1  g14925(.A0(new_n17359_), .A1(new_n12509_), .B0(new_n17361_), .Y(new_n17362_));
  OR2X1    g14926(.A(new_n17348_), .B(pi0781), .Y(new_n17363_));
  OAI21X1  g14927(.A0(new_n17355_), .A1(new_n17350_), .B0(pi0781), .Y(new_n17364_));
  NAND3X1  g14928(.A(new_n17364_), .B(new_n17363_), .C(pi0619), .Y(new_n17365_));
  AOI21X1  g14929(.A0(new_n17306_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n17366_));
  AND2X1   g14930(.A(new_n17366_), .B(new_n17365_), .Y(new_n17367_));
  OR2X1    g14931(.A(new_n17367_), .B(pi0648), .Y(new_n17368_));
  OAI21X1  g14932(.A0(new_n17360_), .A1(pi0619), .B0(pi1159), .Y(new_n17369_));
  AOI21X1  g14933(.A0(new_n17359_), .A1(pi0619), .B0(new_n17369_), .Y(new_n17370_));
  NAND3X1  g14934(.A(new_n17364_), .B(new_n17363_), .C(new_n12509_), .Y(new_n17371_));
  AOI21X1  g14935(.A0(new_n17306_), .A1(pi0619), .B0(pi1159), .Y(new_n17372_));
  AND2X1   g14936(.A(new_n17372_), .B(new_n17371_), .Y(new_n17373_));
  OR2X1    g14937(.A(new_n17373_), .B(new_n12517_), .Y(new_n17374_));
  OAI22X1  g14938(.A0(new_n17374_), .A1(new_n17370_), .B0(new_n17368_), .B1(new_n17362_), .Y(new_n17375_));
  MX2X1    g14939(.A(new_n17375_), .B(new_n17359_), .S0(new_n11766_), .Y(new_n17376_));
  OR2X1    g14940(.A(new_n17376_), .B(pi0788), .Y(new_n17377_));
  MX2X1    g14941(.A(new_n17360_), .B(new_n17313_), .S0(new_n12531_), .Y(new_n17378_));
  AOI21X1  g14942(.A0(new_n17378_), .A1(pi0626), .B0(pi0641), .Y(new_n17379_));
  OAI21X1  g14943(.A0(new_n17376_), .A1(pi0626), .B0(new_n17379_), .Y(new_n17380_));
  AND2X1   g14944(.A(new_n17364_), .B(new_n17363_), .Y(new_n17381_));
  AOI22X1  g14945(.A0(new_n17372_), .A1(new_n17371_), .B0(new_n17366_), .B1(new_n17365_), .Y(new_n17382_));
  MX2X1    g14946(.A(new_n17382_), .B(new_n17381_), .S0(new_n11766_), .Y(new_n17383_));
  AOI21X1  g14947(.A0(new_n17313_), .A1(pi0626), .B0(new_n12543_), .Y(new_n17384_));
  OAI21X1  g14948(.A0(new_n17383_), .A1(pi0626), .B0(new_n17384_), .Y(new_n17385_));
  AND2X1   g14949(.A(new_n17385_), .B(new_n12548_), .Y(new_n17386_));
  AOI21X1  g14950(.A0(new_n17378_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n17387_));
  OAI21X1  g14951(.A0(new_n17376_), .A1(new_n12542_), .B0(new_n17387_), .Y(new_n17388_));
  AOI21X1  g14952(.A0(new_n17313_), .A1(new_n12542_), .B0(pi0641), .Y(new_n17389_));
  OAI21X1  g14953(.A0(new_n17383_), .A1(new_n12542_), .B0(new_n17389_), .Y(new_n17390_));
  AND2X1   g14954(.A(new_n17390_), .B(pi1158), .Y(new_n17391_));
  AOI22X1  g14955(.A0(new_n17391_), .A1(new_n17388_), .B0(new_n17386_), .B1(new_n17380_), .Y(new_n17392_));
  OAI21X1  g14956(.A0(new_n17392_), .A1(new_n11765_), .B0(new_n17377_), .Y(new_n17393_));
  MX2X1    g14957(.A(new_n17383_), .B(new_n17306_), .S0(new_n12708_), .Y(new_n17394_));
  AOI21X1  g14958(.A0(new_n17394_), .A1(pi0628), .B0(pi1156), .Y(new_n17395_));
  OAI21X1  g14959(.A0(new_n17393_), .A1(pi0628), .B0(new_n17395_), .Y(new_n17396_));
  MX2X1    g14960(.A(new_n17378_), .B(new_n17313_), .S0(new_n12563_), .Y(new_n17397_));
  AOI21X1  g14961(.A0(new_n17306_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n17398_));
  OAI21X1  g14962(.A0(new_n17397_), .A1(new_n12554_), .B0(new_n17398_), .Y(new_n17399_));
  AND2X1   g14963(.A(new_n17399_), .B(new_n12561_), .Y(new_n17400_));
  AOI21X1  g14964(.A0(new_n17394_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n17401_));
  OAI21X1  g14965(.A0(new_n17393_), .A1(new_n12554_), .B0(new_n17401_), .Y(new_n17402_));
  AOI21X1  g14966(.A0(new_n17306_), .A1(pi0628), .B0(pi1156), .Y(new_n17403_));
  OAI21X1  g14967(.A0(new_n17397_), .A1(pi0628), .B0(new_n17403_), .Y(new_n17404_));
  AND2X1   g14968(.A(new_n17404_), .B(pi0629), .Y(new_n17405_));
  AOI22X1  g14969(.A0(new_n17405_), .A1(new_n17402_), .B0(new_n17400_), .B1(new_n17396_), .Y(new_n17406_));
  MX2X1    g14970(.A(new_n17406_), .B(new_n17393_), .S0(new_n11764_), .Y(new_n17407_));
  MX2X1    g14971(.A(new_n17394_), .B(new_n17306_), .S0(new_n12580_), .Y(new_n17408_));
  AOI21X1  g14972(.A0(new_n17408_), .A1(pi0647), .B0(pi1157), .Y(new_n17409_));
  OAI21X1  g14973(.A0(new_n17407_), .A1(pi0647), .B0(new_n17409_), .Y(new_n17410_));
  AOI21X1  g14974(.A0(new_n17404_), .A1(new_n17399_), .B0(new_n11764_), .Y(new_n17411_));
  AOI21X1  g14975(.A0(new_n17397_), .A1(new_n11764_), .B0(new_n17411_), .Y(new_n17412_));
  INVX1    g14976(.A(new_n17412_), .Y(new_n17413_));
  AOI21X1  g14977(.A0(new_n17306_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n17414_));
  OAI21X1  g14978(.A0(new_n17413_), .A1(new_n12577_), .B0(new_n17414_), .Y(new_n17415_));
  AND2X1   g14979(.A(new_n17415_), .B(new_n12592_), .Y(new_n17416_));
  AOI21X1  g14980(.A0(new_n17408_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n17417_));
  OAI21X1  g14981(.A0(new_n17407_), .A1(new_n12577_), .B0(new_n17417_), .Y(new_n17418_));
  AOI21X1  g14982(.A0(new_n17306_), .A1(pi0647), .B0(pi1157), .Y(new_n17419_));
  OAI21X1  g14983(.A0(new_n17413_), .A1(pi0647), .B0(new_n17419_), .Y(new_n17420_));
  AND2X1   g14984(.A(new_n17420_), .B(pi0630), .Y(new_n17421_));
  AOI22X1  g14985(.A0(new_n17421_), .A1(new_n17418_), .B0(new_n17416_), .B1(new_n17410_), .Y(new_n17422_));
  OR2X1    g14986(.A(new_n17407_), .B(pi0787), .Y(new_n17423_));
  OAI21X1  g14987(.A0(new_n17422_), .A1(new_n11763_), .B0(new_n17423_), .Y(new_n17424_));
  NAND2X1  g14988(.A(new_n17420_), .B(new_n17415_), .Y(new_n17425_));
  MX2X1    g14989(.A(new_n17425_), .B(new_n17413_), .S0(new_n11763_), .Y(new_n17426_));
  OAI21X1  g14990(.A0(new_n17426_), .A1(pi0644), .B0(pi0715), .Y(new_n17427_));
  AOI21X1  g14991(.A0(new_n17424_), .A1(pi0644), .B0(new_n17427_), .Y(new_n17428_));
  MX2X1    g14992(.A(new_n17408_), .B(new_n17306_), .S0(new_n12604_), .Y(new_n17429_));
  OAI21X1  g14993(.A0(new_n17313_), .A1(pi0644), .B0(new_n12608_), .Y(new_n17430_));
  AOI21X1  g14994(.A0(new_n17429_), .A1(pi0644), .B0(new_n17430_), .Y(new_n17431_));
  NOR3X1   g14995(.A(new_n17431_), .B(new_n17428_), .C(new_n11762_), .Y(new_n17432_));
  OAI21X1  g14996(.A0(new_n17426_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17433_));
  AOI21X1  g14997(.A0(new_n17424_), .A1(new_n12612_), .B0(new_n17433_), .Y(new_n17434_));
  OAI21X1  g14998(.A0(new_n17313_), .A1(new_n12612_), .B0(pi0715), .Y(new_n17435_));
  AOI21X1  g14999(.A0(new_n17429_), .A1(new_n12612_), .B0(new_n17435_), .Y(new_n17436_));
  OR2X1    g15000(.A(new_n17436_), .B(pi1160), .Y(new_n17437_));
  OAI21X1  g15001(.A0(new_n17437_), .A1(new_n17434_), .B0(pi0790), .Y(new_n17438_));
  MX2X1    g15002(.A(new_n17422_), .B(new_n17407_), .S0(new_n11763_), .Y(new_n17439_));
  AOI21X1  g15003(.A0(new_n17439_), .A1(new_n12766_), .B0(po1038), .Y(new_n17440_));
  OAI21X1  g15004(.A0(new_n17438_), .A1(new_n17432_), .B0(new_n17440_), .Y(new_n17441_));
  AOI21X1  g15005(.A0(po1038), .A1(new_n17285_), .B0(pi0832), .Y(new_n17442_));
  AOI21X1  g15006(.A0(pi1093), .A1(pi1092), .B0(pi0179), .Y(new_n17443_));
  INVX1    g15007(.A(new_n17443_), .Y(new_n17444_));
  AOI21X1  g15008(.A0(new_n12056_), .A1(new_n14955_), .B0(new_n17443_), .Y(new_n17445_));
  AOI21X1  g15009(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n17445_), .Y(new_n17446_));
  INVX1    g15010(.A(new_n17445_), .Y(new_n17447_));
  AOI21X1  g15011(.A0(new_n17447_), .A1(new_n14331_), .B0(new_n12463_), .Y(new_n17448_));
  AOI21X1  g15012(.A0(new_n17446_), .A1(new_n12646_), .B0(pi1155), .Y(new_n17449_));
  OAI21X1  g15013(.A0(new_n17449_), .A1(new_n17448_), .B0(pi0785), .Y(new_n17450_));
  OAI21X1  g15014(.A0(new_n17446_), .A1(pi0785), .B0(new_n17450_), .Y(new_n17451_));
  INVX1    g15015(.A(new_n17451_), .Y(new_n17452_));
  AOI21X1  g15016(.A0(new_n17452_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n17453_));
  AOI21X1  g15017(.A0(new_n17452_), .A1(new_n12655_), .B0(pi1154), .Y(new_n17454_));
  NOR2X1   g15018(.A(new_n17454_), .B(new_n17453_), .Y(new_n17455_));
  MX2X1    g15019(.A(new_n17455_), .B(new_n17452_), .S0(new_n11767_), .Y(new_n17456_));
  NOR2X1   g15020(.A(new_n17456_), .B(pi0789), .Y(new_n17457_));
  INVX1    g15021(.A(new_n17456_), .Y(new_n17458_));
  AOI21X1  g15022(.A0(new_n17443_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n17459_));
  OAI21X1  g15023(.A0(new_n17458_), .A1(new_n12509_), .B0(new_n17459_), .Y(new_n17460_));
  AOI21X1  g15024(.A0(new_n17443_), .A1(pi0619), .B0(pi1159), .Y(new_n17461_));
  OAI21X1  g15025(.A0(new_n17458_), .A1(pi0619), .B0(new_n17461_), .Y(new_n17462_));
  AOI21X1  g15026(.A0(new_n17462_), .A1(new_n17460_), .B0(new_n11766_), .Y(new_n17463_));
  NOR2X1   g15027(.A(new_n17463_), .B(new_n17457_), .Y(new_n17464_));
  INVX1    g15028(.A(new_n17464_), .Y(new_n17465_));
  MX2X1    g15029(.A(new_n17465_), .B(new_n17444_), .S0(new_n12708_), .Y(new_n17466_));
  MX2X1    g15030(.A(new_n17466_), .B(new_n17444_), .S0(new_n12580_), .Y(new_n17467_));
  AOI21X1  g15031(.A0(new_n12439_), .A1(new_n14956_), .B0(new_n17443_), .Y(new_n17468_));
  AND3X1   g15032(.A(new_n12439_), .B(new_n14956_), .C(new_n12363_), .Y(new_n17469_));
  NOR2X1   g15033(.A(new_n17469_), .B(new_n17468_), .Y(new_n17470_));
  NOR2X1   g15034(.A(new_n17443_), .B(pi1153), .Y(new_n17471_));
  INVX1    g15035(.A(new_n17471_), .Y(new_n17472_));
  OAI22X1  g15036(.A0(new_n17472_), .A1(new_n17469_), .B0(new_n17470_), .B1(new_n12364_), .Y(new_n17473_));
  MX2X1    g15037(.A(new_n17473_), .B(new_n17468_), .S0(new_n11769_), .Y(new_n17474_));
  NOR4X1   g15038(.A(new_n17474_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n17475_));
  AND3X1   g15039(.A(new_n17475_), .B(new_n12739_), .C(new_n12718_), .Y(new_n17476_));
  INVX1    g15040(.A(new_n17476_), .Y(new_n17477_));
  AOI21X1  g15041(.A0(new_n17443_), .A1(pi0647), .B0(pi1157), .Y(new_n17478_));
  OAI21X1  g15042(.A0(new_n17477_), .A1(pi0647), .B0(new_n17478_), .Y(new_n17479_));
  MX2X1    g15043(.A(new_n17476_), .B(new_n17443_), .S0(new_n12577_), .Y(new_n17480_));
  OAI22X1  g15044(.A0(new_n17480_), .A1(new_n14242_), .B0(new_n17479_), .B1(new_n12592_), .Y(new_n17481_));
  AOI21X1  g15045(.A0(new_n17467_), .A1(new_n14326_), .B0(new_n17481_), .Y(new_n17482_));
  AOI21X1  g15046(.A0(new_n17444_), .A1(pi0626), .B0(new_n16218_), .Y(new_n17483_));
  OAI21X1  g15047(.A0(new_n17464_), .A1(pi0626), .B0(new_n17483_), .Y(new_n17484_));
  AOI21X1  g15048(.A0(new_n17444_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n17485_));
  OAI21X1  g15049(.A0(new_n17464_), .A1(new_n12542_), .B0(new_n17485_), .Y(new_n17486_));
  NAND2X1  g15050(.A(new_n17475_), .B(new_n12637_), .Y(new_n17487_));
  AND3X1   g15051(.A(new_n17487_), .B(new_n17486_), .C(new_n17484_), .Y(new_n17488_));
  NOR2X1   g15052(.A(new_n17488_), .B(new_n11765_), .Y(new_n17489_));
  INVX1    g15053(.A(new_n17489_), .Y(new_n17490_));
  NOR2X1   g15054(.A(new_n17468_), .B(new_n11991_), .Y(new_n17491_));
  MX2X1    g15055(.A(new_n17447_), .B(new_n12363_), .S0(new_n17491_), .Y(new_n17492_));
  NOR2X1   g15056(.A(new_n17492_), .B(new_n17472_), .Y(new_n17493_));
  OAI21X1  g15057(.A0(new_n17470_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n17494_));
  NOR2X1   g15058(.A(new_n17494_), .B(new_n17493_), .Y(new_n17495_));
  OR3X1    g15059(.A(new_n17468_), .B(new_n11991_), .C(new_n12363_), .Y(new_n17496_));
  AND2X1   g15060(.A(new_n17445_), .B(pi1153), .Y(new_n17497_));
  OAI21X1  g15061(.A0(new_n17472_), .A1(new_n17469_), .B0(pi0608), .Y(new_n17498_));
  AOI21X1  g15062(.A0(new_n17497_), .A1(new_n17496_), .B0(new_n17498_), .Y(new_n17499_));
  OAI21X1  g15063(.A0(new_n17499_), .A1(new_n17495_), .B0(pi0778), .Y(new_n17500_));
  OAI21X1  g15064(.A0(new_n17491_), .A1(new_n17447_), .B0(new_n11769_), .Y(new_n17501_));
  NAND2X1  g15065(.A(new_n17501_), .B(new_n17500_), .Y(new_n17502_));
  INVX1    g15066(.A(new_n17502_), .Y(new_n17503_));
  OAI21X1  g15067(.A0(new_n17474_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n17504_));
  AOI21X1  g15068(.A0(new_n17502_), .A1(new_n12462_), .B0(new_n17504_), .Y(new_n17505_));
  NOR3X1   g15069(.A(new_n17505_), .B(new_n17448_), .C(pi0660), .Y(new_n17506_));
  OAI21X1  g15070(.A0(new_n17474_), .A1(pi0609), .B0(pi1155), .Y(new_n17507_));
  AOI21X1  g15071(.A0(new_n17502_), .A1(pi0609), .B0(new_n17507_), .Y(new_n17508_));
  NOR3X1   g15072(.A(new_n17508_), .B(new_n17449_), .C(new_n12468_), .Y(new_n17509_));
  NOR2X1   g15073(.A(new_n17509_), .B(new_n17506_), .Y(new_n17510_));
  MX2X1    g15074(.A(new_n17510_), .B(new_n17503_), .S0(new_n11768_), .Y(new_n17511_));
  OR3X1    g15075(.A(new_n17474_), .B(new_n12630_), .C(new_n12486_), .Y(new_n17512_));
  AND2X1   g15076(.A(new_n17512_), .B(new_n12487_), .Y(new_n17513_));
  OAI21X1  g15077(.A0(new_n17511_), .A1(pi0618), .B0(new_n17513_), .Y(new_n17514_));
  NOR2X1   g15078(.A(new_n17453_), .B(pi0627), .Y(new_n17515_));
  NOR3X1   g15079(.A(new_n17474_), .B(new_n12630_), .C(pi0618), .Y(new_n17516_));
  NOR2X1   g15080(.A(new_n17516_), .B(new_n12487_), .Y(new_n17517_));
  OAI21X1  g15081(.A0(new_n17511_), .A1(new_n12486_), .B0(new_n17517_), .Y(new_n17518_));
  NOR2X1   g15082(.A(new_n17454_), .B(new_n12494_), .Y(new_n17519_));
  AOI22X1  g15083(.A0(new_n17519_), .A1(new_n17518_), .B0(new_n17515_), .B1(new_n17514_), .Y(new_n17520_));
  MX2X1    g15084(.A(new_n17520_), .B(new_n17511_), .S0(new_n11767_), .Y(new_n17521_));
  OR4X1    g15085(.A(new_n17474_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n17522_));
  AND2X1   g15086(.A(new_n17522_), .B(new_n12510_), .Y(new_n17523_));
  OAI21X1  g15087(.A0(new_n17521_), .A1(pi0619), .B0(new_n17523_), .Y(new_n17524_));
  AND3X1   g15088(.A(new_n17524_), .B(new_n17460_), .C(new_n12517_), .Y(new_n17525_));
  NOR4X1   g15089(.A(new_n17474_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n17526_));
  NOR2X1   g15090(.A(new_n17526_), .B(new_n12510_), .Y(new_n17527_));
  OAI21X1  g15091(.A0(new_n17521_), .A1(new_n12509_), .B0(new_n17527_), .Y(new_n17528_));
  AND2X1   g15092(.A(new_n17462_), .B(pi0648), .Y(new_n17529_));
  AOI21X1  g15093(.A0(new_n17529_), .A1(new_n17528_), .B0(new_n11766_), .Y(new_n17530_));
  INVX1    g15094(.A(new_n17530_), .Y(new_n17531_));
  AOI21X1  g15095(.A0(new_n17521_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n17532_));
  OAI21X1  g15096(.A0(new_n17531_), .A1(new_n17525_), .B0(new_n17532_), .Y(new_n17533_));
  AOI21X1  g15097(.A0(new_n17533_), .A1(new_n17490_), .B0(new_n14125_), .Y(new_n17534_));
  INVX1    g15098(.A(new_n17466_), .Y(new_n17535_));
  AND2X1   g15099(.A(new_n17475_), .B(new_n12718_), .Y(new_n17536_));
  AOI22X1  g15100(.A0(new_n17536_), .A1(new_n14426_), .B0(new_n17535_), .B1(new_n12735_), .Y(new_n17537_));
  AOI22X1  g15101(.A0(new_n17536_), .A1(new_n14428_), .B0(new_n17535_), .B1(new_n12733_), .Y(new_n17538_));
  MX2X1    g15102(.A(new_n17538_), .B(new_n17537_), .S0(new_n12561_), .Y(new_n17539_));
  OAI21X1  g15103(.A0(new_n17539_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n17540_));
  OAI22X1  g15104(.A0(new_n17540_), .A1(new_n17534_), .B0(new_n17482_), .B1(new_n11763_), .Y(new_n17541_));
  INVX1    g15105(.A(new_n17541_), .Y(new_n17542_));
  OAI21X1  g15106(.A0(new_n17480_), .A1(new_n12578_), .B0(new_n17479_), .Y(new_n17543_));
  MX2X1    g15107(.A(new_n17543_), .B(new_n17477_), .S0(new_n11763_), .Y(new_n17544_));
  OAI21X1  g15108(.A0(new_n17544_), .A1(pi0644), .B0(pi0715), .Y(new_n17545_));
  AOI21X1  g15109(.A0(new_n17542_), .A1(pi0644), .B0(new_n17545_), .Y(new_n17546_));
  OR3X1    g15110(.A(new_n17444_), .B(new_n12603_), .C(new_n11763_), .Y(new_n17547_));
  OAI21X1  g15111(.A0(new_n17467_), .A1(new_n12604_), .B0(new_n17547_), .Y(new_n17548_));
  OAI21X1  g15112(.A0(new_n17444_), .A1(pi0644), .B0(new_n12608_), .Y(new_n17549_));
  AOI21X1  g15113(.A0(new_n17548_), .A1(pi0644), .B0(new_n17549_), .Y(new_n17550_));
  OR2X1    g15114(.A(new_n17550_), .B(new_n11762_), .Y(new_n17551_));
  OAI21X1  g15115(.A0(new_n17544_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17552_));
  AOI21X1  g15116(.A0(new_n17542_), .A1(new_n12612_), .B0(new_n17552_), .Y(new_n17553_));
  OAI21X1  g15117(.A0(new_n17444_), .A1(new_n12612_), .B0(pi0715), .Y(new_n17554_));
  AOI21X1  g15118(.A0(new_n17548_), .A1(new_n12612_), .B0(new_n17554_), .Y(new_n17555_));
  OR2X1    g15119(.A(new_n17555_), .B(pi1160), .Y(new_n17556_));
  OAI22X1  g15120(.A0(new_n17556_), .A1(new_n17553_), .B0(new_n17551_), .B1(new_n17546_), .Y(new_n17557_));
  OAI21X1  g15121(.A0(new_n17541_), .A1(pi0790), .B0(pi0832), .Y(new_n17558_));
  AOI21X1  g15122(.A0(new_n17557_), .A1(pi0790), .B0(new_n17558_), .Y(new_n17559_));
  AOI21X1  g15123(.A0(new_n17442_), .A1(new_n17441_), .B0(new_n17559_), .Y(po0336));
  AOI21X1  g15124(.A0(pi1093), .A1(pi1092), .B0(pi0180), .Y(new_n17561_));
  INVX1    g15125(.A(new_n17561_), .Y(new_n17562_));
  AOI21X1  g15126(.A0(new_n12056_), .A1(new_n15006_), .B0(new_n17561_), .Y(new_n17563_));
  INVX1    g15127(.A(new_n17563_), .Y(new_n17564_));
  NAND2X1  g15128(.A(new_n17564_), .B(new_n15771_), .Y(new_n17565_));
  AND3X1   g15129(.A(new_n12480_), .B(new_n12056_), .C(new_n15006_), .Y(new_n17566_));
  OAI21X1  g15130(.A0(new_n17566_), .A1(new_n17565_), .B0(pi1155), .Y(new_n17567_));
  NOR3X1   g15131(.A(new_n17566_), .B(new_n17561_), .C(pi1155), .Y(new_n17568_));
  INVX1    g15132(.A(new_n17568_), .Y(new_n17569_));
  AOI21X1  g15133(.A0(new_n17569_), .A1(new_n17567_), .B0(new_n11768_), .Y(new_n17570_));
  AOI21X1  g15134(.A0(new_n17565_), .A1(new_n11768_), .B0(new_n17570_), .Y(new_n17571_));
  AOI21X1  g15135(.A0(new_n17571_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n17572_));
  AOI21X1  g15136(.A0(new_n17571_), .A1(new_n12655_), .B0(pi1154), .Y(new_n17573_));
  NOR2X1   g15137(.A(new_n17573_), .B(new_n17572_), .Y(new_n17574_));
  MX2X1    g15138(.A(new_n17574_), .B(new_n17571_), .S0(new_n11767_), .Y(new_n17575_));
  NOR2X1   g15139(.A(new_n17575_), .B(pi0789), .Y(new_n17576_));
  AOI21X1  g15140(.A0(new_n17575_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n17577_));
  AOI21X1  g15141(.A0(new_n17575_), .A1(new_n15790_), .B0(pi1159), .Y(new_n17578_));
  OR2X1    g15142(.A(new_n17578_), .B(new_n17577_), .Y(new_n17579_));
  AOI21X1  g15143(.A0(new_n17579_), .A1(pi0789), .B0(new_n17576_), .Y(new_n17580_));
  INVX1    g15144(.A(new_n17580_), .Y(new_n17581_));
  MX2X1    g15145(.A(new_n17581_), .B(new_n17562_), .S0(new_n12708_), .Y(new_n17582_));
  MX2X1    g15146(.A(new_n17582_), .B(new_n17562_), .S0(new_n12580_), .Y(new_n17583_));
  AOI21X1  g15147(.A0(new_n12439_), .A1(new_n15025_), .B0(new_n17561_), .Y(new_n17584_));
  OR2X1    g15148(.A(new_n17584_), .B(pi0778), .Y(new_n17585_));
  INVX1    g15149(.A(new_n17584_), .Y(new_n17586_));
  AND3X1   g15150(.A(new_n12439_), .B(new_n15025_), .C(new_n12363_), .Y(new_n17587_));
  INVX1    g15151(.A(new_n17587_), .Y(new_n17588_));
  AOI21X1  g15152(.A0(new_n17588_), .A1(new_n17586_), .B0(new_n12364_), .Y(new_n17589_));
  NOR3X1   g15153(.A(new_n17587_), .B(new_n17561_), .C(pi1153), .Y(new_n17590_));
  OR3X1    g15154(.A(new_n17590_), .B(new_n17589_), .C(new_n11769_), .Y(new_n17591_));
  AND2X1   g15155(.A(new_n17591_), .B(new_n17585_), .Y(new_n17592_));
  NOR4X1   g15156(.A(new_n17592_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n17593_));
  AND3X1   g15157(.A(new_n17593_), .B(new_n12739_), .C(new_n12718_), .Y(new_n17594_));
  INVX1    g15158(.A(new_n17594_), .Y(new_n17595_));
  AOI21X1  g15159(.A0(new_n17561_), .A1(pi0647), .B0(pi1157), .Y(new_n17596_));
  OAI21X1  g15160(.A0(new_n17595_), .A1(pi0647), .B0(new_n17596_), .Y(new_n17597_));
  MX2X1    g15161(.A(new_n17594_), .B(new_n17561_), .S0(new_n12577_), .Y(new_n17598_));
  OAI22X1  g15162(.A0(new_n17598_), .A1(new_n14242_), .B0(new_n17597_), .B1(new_n12592_), .Y(new_n17599_));
  AOI21X1  g15163(.A0(new_n17583_), .A1(new_n14326_), .B0(new_n17599_), .Y(new_n17600_));
  NOR2X1   g15164(.A(new_n17600_), .B(new_n11763_), .Y(new_n17601_));
  AOI21X1  g15165(.A0(new_n17562_), .A1(pi0626), .B0(new_n16218_), .Y(new_n17602_));
  OAI21X1  g15166(.A0(new_n17580_), .A1(pi0626), .B0(new_n17602_), .Y(new_n17603_));
  AOI21X1  g15167(.A0(new_n17562_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n17604_));
  OAI21X1  g15168(.A0(new_n17580_), .A1(new_n12542_), .B0(new_n17604_), .Y(new_n17605_));
  NAND2X1  g15169(.A(new_n17593_), .B(new_n12637_), .Y(new_n17606_));
  AND3X1   g15170(.A(new_n17606_), .B(new_n17605_), .C(new_n17603_), .Y(new_n17607_));
  NOR2X1   g15171(.A(new_n17607_), .B(new_n11765_), .Y(new_n17608_));
  NOR2X1   g15172(.A(new_n17561_), .B(pi1153), .Y(new_n17609_));
  NOR3X1   g15173(.A(new_n17584_), .B(new_n11991_), .C(new_n12363_), .Y(new_n17610_));
  AOI21X1  g15174(.A0(new_n17586_), .A1(new_n12048_), .B0(new_n17564_), .Y(new_n17611_));
  OAI21X1  g15175(.A0(new_n17611_), .A1(new_n17610_), .B0(new_n17609_), .Y(new_n17612_));
  NOR2X1   g15176(.A(new_n17589_), .B(pi0608), .Y(new_n17613_));
  NOR3X1   g15177(.A(new_n17610_), .B(new_n17564_), .C(new_n12364_), .Y(new_n17614_));
  NOR3X1   g15178(.A(new_n17614_), .B(new_n17590_), .C(new_n12368_), .Y(new_n17615_));
  AOI21X1  g15179(.A0(new_n17613_), .A1(new_n17612_), .B0(new_n17615_), .Y(new_n17616_));
  OR2X1    g15180(.A(new_n17611_), .B(pi0778), .Y(new_n17617_));
  OAI21X1  g15181(.A0(new_n17616_), .A1(new_n11769_), .B0(new_n17617_), .Y(new_n17618_));
  INVX1    g15182(.A(new_n17618_), .Y(new_n17619_));
  AND2X1   g15183(.A(new_n17618_), .B(new_n12462_), .Y(new_n17620_));
  OAI21X1  g15184(.A0(new_n17592_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n17621_));
  OR2X1    g15185(.A(new_n17621_), .B(new_n17620_), .Y(new_n17622_));
  AND3X1   g15186(.A(new_n17622_), .B(new_n17567_), .C(new_n12468_), .Y(new_n17623_));
  OAI21X1  g15187(.A0(new_n17592_), .A1(pi0609), .B0(pi1155), .Y(new_n17624_));
  AOI21X1  g15188(.A0(new_n17618_), .A1(pi0609), .B0(new_n17624_), .Y(new_n17625_));
  NOR3X1   g15189(.A(new_n17625_), .B(new_n17568_), .C(new_n12468_), .Y(new_n17626_));
  NOR2X1   g15190(.A(new_n17626_), .B(new_n17623_), .Y(new_n17627_));
  MX2X1    g15191(.A(new_n17627_), .B(new_n17619_), .S0(new_n11768_), .Y(new_n17628_));
  AOI21X1  g15192(.A0(new_n17591_), .A1(new_n17585_), .B0(new_n12630_), .Y(new_n17629_));
  AOI21X1  g15193(.A0(new_n17629_), .A1(pi0618), .B0(pi1154), .Y(new_n17630_));
  OAI21X1  g15194(.A0(new_n17628_), .A1(pi0618), .B0(new_n17630_), .Y(new_n17631_));
  NOR2X1   g15195(.A(new_n17572_), .B(pi0627), .Y(new_n17632_));
  AOI21X1  g15196(.A0(new_n17629_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17633_));
  OAI21X1  g15197(.A0(new_n17628_), .A1(new_n12486_), .B0(new_n17633_), .Y(new_n17634_));
  NOR2X1   g15198(.A(new_n17573_), .B(new_n12494_), .Y(new_n17635_));
  AOI22X1  g15199(.A0(new_n17635_), .A1(new_n17634_), .B0(new_n17632_), .B1(new_n17631_), .Y(new_n17636_));
  MX2X1    g15200(.A(new_n17636_), .B(new_n17628_), .S0(new_n11767_), .Y(new_n17637_));
  OR4X1    g15201(.A(new_n17592_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n17638_));
  AND2X1   g15202(.A(new_n17638_), .B(new_n12510_), .Y(new_n17639_));
  OAI21X1  g15203(.A0(new_n17637_), .A1(pi0619), .B0(new_n17639_), .Y(new_n17640_));
  NOR2X1   g15204(.A(new_n17577_), .B(pi0648), .Y(new_n17641_));
  AND2X1   g15205(.A(new_n17641_), .B(new_n17640_), .Y(new_n17642_));
  NOR4X1   g15206(.A(new_n17592_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n17643_));
  NOR2X1   g15207(.A(new_n17643_), .B(new_n12510_), .Y(new_n17644_));
  OAI21X1  g15208(.A0(new_n17637_), .A1(new_n12509_), .B0(new_n17644_), .Y(new_n17645_));
  NOR2X1   g15209(.A(new_n17578_), .B(new_n12517_), .Y(new_n17646_));
  AND2X1   g15210(.A(new_n17646_), .B(new_n17645_), .Y(new_n17647_));
  OR3X1    g15211(.A(new_n17647_), .B(new_n17642_), .C(new_n11766_), .Y(new_n17648_));
  AOI21X1  g15212(.A0(new_n17637_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n17649_));
  AOI21X1  g15213(.A0(new_n17649_), .A1(new_n17648_), .B0(new_n17608_), .Y(new_n17650_));
  OR2X1    g15214(.A(new_n17650_), .B(new_n14125_), .Y(new_n17651_));
  INVX1    g15215(.A(new_n17582_), .Y(new_n17652_));
  AND2X1   g15216(.A(new_n17593_), .B(new_n12718_), .Y(new_n17653_));
  AOI22X1  g15217(.A0(new_n17653_), .A1(new_n14426_), .B0(new_n17652_), .B1(new_n12735_), .Y(new_n17654_));
  AOI22X1  g15218(.A0(new_n17653_), .A1(new_n14428_), .B0(new_n17652_), .B1(new_n12733_), .Y(new_n17655_));
  MX2X1    g15219(.A(new_n17655_), .B(new_n17654_), .S0(new_n12561_), .Y(new_n17656_));
  OAI21X1  g15220(.A0(new_n17656_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n17657_));
  INVX1    g15221(.A(new_n17657_), .Y(new_n17658_));
  AOI21X1  g15222(.A0(new_n17658_), .A1(new_n17651_), .B0(new_n17601_), .Y(new_n17659_));
  OAI21X1  g15223(.A0(new_n17598_), .A1(new_n12578_), .B0(new_n17597_), .Y(new_n17660_));
  MX2X1    g15224(.A(new_n17660_), .B(new_n17595_), .S0(new_n11763_), .Y(new_n17661_));
  OAI21X1  g15225(.A0(new_n17661_), .A1(pi0644), .B0(pi0715), .Y(new_n17662_));
  AOI21X1  g15226(.A0(new_n17659_), .A1(pi0644), .B0(new_n17662_), .Y(new_n17663_));
  OR3X1    g15227(.A(new_n17562_), .B(new_n12603_), .C(new_n11763_), .Y(new_n17664_));
  OAI21X1  g15228(.A0(new_n17583_), .A1(new_n12604_), .B0(new_n17664_), .Y(new_n17665_));
  OAI21X1  g15229(.A0(new_n17562_), .A1(pi0644), .B0(new_n12608_), .Y(new_n17666_));
  AOI21X1  g15230(.A0(new_n17665_), .A1(pi0644), .B0(new_n17666_), .Y(new_n17667_));
  OR2X1    g15231(.A(new_n17667_), .B(new_n11762_), .Y(new_n17668_));
  OAI21X1  g15232(.A0(new_n17661_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17669_));
  AOI21X1  g15233(.A0(new_n17659_), .A1(new_n12612_), .B0(new_n17669_), .Y(new_n17670_));
  OAI21X1  g15234(.A0(new_n17562_), .A1(new_n12612_), .B0(pi0715), .Y(new_n17671_));
  AOI21X1  g15235(.A0(new_n17665_), .A1(new_n12612_), .B0(new_n17671_), .Y(new_n17672_));
  OR2X1    g15236(.A(new_n17672_), .B(pi1160), .Y(new_n17673_));
  OAI22X1  g15237(.A0(new_n17673_), .A1(new_n17670_), .B0(new_n17668_), .B1(new_n17663_), .Y(new_n17674_));
  NAND2X1  g15238(.A(new_n17674_), .B(pi0790), .Y(new_n17675_));
  AOI21X1  g15239(.A0(new_n17659_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n17676_));
  AOI21X1  g15240(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0180), .Y(new_n17677_));
  INVX1    g15241(.A(new_n17677_), .Y(new_n17678_));
  AOI21X1  g15242(.A0(new_n3103_), .A1(new_n15025_), .B0(new_n17678_), .Y(new_n17679_));
  OAI21X1  g15243(.A0(new_n12826_), .A1(new_n5203_), .B0(new_n2979_), .Y(new_n17680_));
  AOI22X1  g15244(.A0(new_n17680_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n5203_), .Y(new_n17681_));
  AOI21X1  g15245(.A0(new_n12771_), .A1(new_n5203_), .B0(new_n12441_), .Y(new_n17682_));
  NOR3X1   g15246(.A(new_n17682_), .B(new_n17681_), .C(pi0702), .Y(new_n17683_));
  NOR2X1   g15247(.A(new_n17683_), .B(new_n17679_), .Y(new_n17684_));
  INVX1    g15248(.A(new_n17684_), .Y(new_n17685_));
  AOI21X1  g15249(.A0(new_n17677_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n17686_));
  OAI21X1  g15250(.A0(new_n17684_), .A1(new_n12363_), .B0(new_n17686_), .Y(new_n17687_));
  AOI21X1  g15251(.A0(new_n17677_), .A1(pi0625), .B0(pi1153), .Y(new_n17688_));
  OAI21X1  g15252(.A0(new_n17684_), .A1(pi0625), .B0(new_n17688_), .Y(new_n17689_));
  AND2X1   g15253(.A(new_n17689_), .B(new_n17687_), .Y(new_n17690_));
  MX2X1    g15254(.A(new_n17690_), .B(new_n17685_), .S0(new_n11769_), .Y(new_n17691_));
  MX2X1    g15255(.A(new_n17691_), .B(new_n17677_), .S0(new_n12490_), .Y(new_n17692_));
  INVX1    g15256(.A(new_n17692_), .Y(new_n17693_));
  MX2X1    g15257(.A(new_n17693_), .B(new_n17678_), .S0(new_n12513_), .Y(new_n17694_));
  INVX1    g15258(.A(new_n17694_), .Y(new_n17695_));
  MX2X1    g15259(.A(new_n17695_), .B(new_n17677_), .S0(new_n12531_), .Y(new_n17696_));
  MX2X1    g15260(.A(new_n17696_), .B(new_n17677_), .S0(new_n12563_), .Y(new_n17697_));
  INVX1    g15261(.A(new_n17697_), .Y(new_n17698_));
  AOI21X1  g15262(.A0(new_n17677_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n17699_));
  OAI21X1  g15263(.A0(new_n17698_), .A1(new_n12554_), .B0(new_n17699_), .Y(new_n17700_));
  AOI21X1  g15264(.A0(new_n17677_), .A1(pi0628), .B0(pi1156), .Y(new_n17701_));
  OAI21X1  g15265(.A0(new_n17698_), .A1(pi0628), .B0(new_n17701_), .Y(new_n17702_));
  AOI21X1  g15266(.A0(new_n17702_), .A1(new_n17700_), .B0(new_n11764_), .Y(new_n17703_));
  AOI21X1  g15267(.A0(new_n17698_), .A1(new_n11764_), .B0(new_n17703_), .Y(new_n17704_));
  MX2X1    g15268(.A(new_n17704_), .B(new_n17677_), .S0(pi0647), .Y(new_n17705_));
  MX2X1    g15269(.A(new_n17704_), .B(new_n17677_), .S0(new_n12577_), .Y(new_n17706_));
  MX2X1    g15270(.A(new_n17706_), .B(new_n17705_), .S0(new_n12578_), .Y(new_n17707_));
  MX2X1    g15271(.A(new_n17707_), .B(new_n17704_), .S0(new_n11763_), .Y(new_n17708_));
  AOI21X1  g15272(.A0(new_n17708_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17709_));
  AOI22X1  g15273(.A0(new_n12073_), .A1(pi0180), .B0(new_n12444_), .B1(pi0753), .Y(new_n17710_));
  OR3X1    g15274(.A(new_n12776_), .B(pi0753), .C(pi0180), .Y(new_n17711_));
  OAI22X1  g15275(.A0(new_n12045_), .A1(new_n5203_), .B0(new_n11822_), .B1(new_n15006_), .Y(new_n17712_));
  AOI22X1  g15276(.A0(new_n17712_), .A1(new_n2939_), .B0(pi0753), .B1(pi0180), .Y(new_n17713_));
  AND2X1   g15277(.A(new_n17713_), .B(new_n17711_), .Y(new_n17714_));
  OAI21X1  g15278(.A0(new_n17710_), .A1(new_n2939_), .B0(new_n17714_), .Y(new_n17715_));
  AND2X1   g15279(.A(new_n17715_), .B(new_n2979_), .Y(new_n17716_));
  OAI21X1  g15280(.A0(new_n12077_), .A1(pi0180), .B0(pi0038), .Y(new_n17717_));
  AOI21X1  g15281(.A0(new_n12079_), .A1(new_n15006_), .B0(new_n17717_), .Y(new_n17718_));
  OR2X1    g15282(.A(new_n17718_), .B(new_n17716_), .Y(new_n17719_));
  MX2X1    g15283(.A(new_n17719_), .B(pi0180), .S0(new_n11770_), .Y(new_n17720_));
  AND2X1   g15284(.A(new_n17720_), .B(new_n12474_), .Y(new_n17721_));
  AOI21X1  g15285(.A0(new_n17678_), .A1(new_n12473_), .B0(new_n17721_), .Y(new_n17722_));
  AOI22X1  g15286(.A0(new_n17721_), .A1(pi0609), .B0(new_n17678_), .B1(new_n12472_), .Y(new_n17723_));
  AOI22X1  g15287(.A0(new_n17721_), .A1(new_n12462_), .B0(new_n17678_), .B1(new_n12481_), .Y(new_n17724_));
  MX2X1    g15288(.A(new_n17724_), .B(new_n17723_), .S0(pi1155), .Y(new_n17725_));
  MX2X1    g15289(.A(new_n17725_), .B(new_n17722_), .S0(new_n11768_), .Y(new_n17726_));
  OAI21X1  g15290(.A0(new_n17678_), .A1(pi0618), .B0(pi1154), .Y(new_n17727_));
  AOI21X1  g15291(.A0(new_n17726_), .A1(pi0618), .B0(new_n17727_), .Y(new_n17728_));
  OAI21X1  g15292(.A0(new_n17678_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17729_));
  AOI21X1  g15293(.A0(new_n17726_), .A1(new_n12486_), .B0(new_n17729_), .Y(new_n17730_));
  NOR2X1   g15294(.A(new_n17730_), .B(new_n17728_), .Y(new_n17731_));
  MX2X1    g15295(.A(new_n17731_), .B(new_n17726_), .S0(new_n11767_), .Y(new_n17732_));
  OAI21X1  g15296(.A0(new_n17678_), .A1(pi0619), .B0(pi1159), .Y(new_n17733_));
  AOI21X1  g15297(.A0(new_n17732_), .A1(pi0619), .B0(new_n17733_), .Y(new_n17734_));
  OAI21X1  g15298(.A0(new_n17678_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n17735_));
  AOI21X1  g15299(.A0(new_n17732_), .A1(new_n12509_), .B0(new_n17735_), .Y(new_n17736_));
  NOR2X1   g15300(.A(new_n17736_), .B(new_n17734_), .Y(new_n17737_));
  MX2X1    g15301(.A(new_n17737_), .B(new_n17732_), .S0(new_n11766_), .Y(new_n17738_));
  AND2X1   g15302(.A(new_n17677_), .B(new_n12708_), .Y(new_n17739_));
  AOI21X1  g15303(.A0(new_n17738_), .A1(new_n16140_), .B0(new_n17739_), .Y(new_n17740_));
  NAND2X1  g15304(.A(new_n17677_), .B(new_n12580_), .Y(new_n17741_));
  OAI21X1  g15305(.A0(new_n17740_), .A1(new_n12580_), .B0(new_n17741_), .Y(new_n17742_));
  MX2X1    g15306(.A(new_n17742_), .B(new_n17677_), .S0(new_n12604_), .Y(new_n17743_));
  OAI21X1  g15307(.A0(new_n17678_), .A1(pi0644), .B0(new_n12608_), .Y(new_n17744_));
  AOI21X1  g15308(.A0(new_n17743_), .A1(pi0644), .B0(new_n17744_), .Y(new_n17745_));
  OR2X1    g15309(.A(new_n17745_), .B(new_n11762_), .Y(new_n17746_));
  AOI21X1  g15310(.A0(new_n17708_), .A1(pi0644), .B0(pi0715), .Y(new_n17747_));
  OAI21X1  g15311(.A0(new_n17678_), .A1(new_n12612_), .B0(pi0715), .Y(new_n17748_));
  AOI21X1  g15312(.A0(new_n17743_), .A1(new_n12612_), .B0(new_n17748_), .Y(new_n17749_));
  OR2X1    g15313(.A(new_n17749_), .B(pi1160), .Y(new_n17750_));
  OAI22X1  g15314(.A0(new_n17750_), .A1(new_n17747_), .B0(new_n17746_), .B1(new_n17709_), .Y(new_n17751_));
  OR3X1    g15315(.A(new_n17749_), .B(pi1160), .C(pi0644), .Y(new_n17752_));
  OR3X1    g15316(.A(new_n17745_), .B(new_n11762_), .C(new_n12612_), .Y(new_n17753_));
  NAND3X1  g15317(.A(new_n17753_), .B(new_n17752_), .C(pi0790), .Y(new_n17754_));
  NAND2X1  g15318(.A(new_n17740_), .B(new_n14249_), .Y(new_n17755_));
  MX2X1    g15319(.A(new_n17702_), .B(new_n17700_), .S0(new_n12561_), .Y(new_n17756_));
  AND2X1   g15320(.A(new_n17756_), .B(new_n17755_), .Y(new_n17757_));
  OR2X1    g15321(.A(new_n17757_), .B(new_n11764_), .Y(new_n17758_));
  OR3X1    g15322(.A(new_n17718_), .B(new_n17716_), .C(new_n15025_), .Y(new_n17759_));
  OAI21X1  g15323(.A0(new_n12213_), .A1(new_n5203_), .B0(pi0753), .Y(new_n17760_));
  AOI21X1  g15324(.A0(new_n12155_), .A1(new_n5203_), .B0(new_n17760_), .Y(new_n17761_));
  AOI21X1  g15325(.A0(new_n12788_), .A1(new_n5203_), .B0(pi0753), .Y(new_n17762_));
  OAI21X1  g15326(.A0(new_n12787_), .A1(new_n5203_), .B0(new_n17762_), .Y(new_n17763_));
  NAND2X1  g15327(.A(new_n17763_), .B(pi0039), .Y(new_n17764_));
  AND2X1   g15328(.A(new_n12332_), .B(pi0180), .Y(new_n17765_));
  OAI21X1  g15329(.A0(new_n12315_), .A1(pi0180), .B0(pi0753), .Y(new_n17766_));
  NOR4X1   g15330(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0180), .Y(new_n17767_));
  OAI21X1  g15331(.A0(new_n12800_), .A1(new_n5203_), .B0(new_n15006_), .Y(new_n17768_));
  OAI22X1  g15332(.A0(new_n17768_), .A1(new_n17767_), .B0(new_n17766_), .B1(new_n17765_), .Y(new_n17769_));
  AOI21X1  g15333(.A0(new_n17769_), .A1(new_n2939_), .B0(pi0038), .Y(new_n17770_));
  OAI21X1  g15334(.A0(new_n17764_), .A1(new_n17761_), .B0(new_n17770_), .Y(new_n17771_));
  OAI21X1  g15335(.A0(new_n12276_), .A1(pi0753), .B0(new_n13540_), .Y(new_n17772_));
  NAND2X1  g15336(.A(new_n17772_), .B(new_n5203_), .Y(new_n17773_));
  AOI21X1  g15337(.A0(new_n12056_), .A1(new_n15006_), .B0(new_n13443_), .Y(new_n17774_));
  NOR2X1   g15338(.A(new_n17774_), .B(new_n5203_), .Y(new_n17775_));
  AOI21X1  g15339(.A0(new_n17775_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n17776_));
  AOI21X1  g15340(.A0(new_n17776_), .A1(new_n17773_), .B0(pi0702), .Y(new_n17777_));
  AOI21X1  g15341(.A0(new_n17777_), .A1(new_n17771_), .B0(new_n11770_), .Y(new_n17778_));
  AOI22X1  g15342(.A0(new_n17778_), .A1(new_n17759_), .B0(new_n11770_), .B1(pi0180), .Y(new_n17779_));
  AND2X1   g15343(.A(new_n17779_), .B(new_n12363_), .Y(new_n17780_));
  OAI21X1  g15344(.A0(new_n17720_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n17781_));
  OR2X1    g15345(.A(new_n17781_), .B(new_n17780_), .Y(new_n17782_));
  NAND3X1  g15346(.A(new_n17782_), .B(new_n17687_), .C(new_n12368_), .Y(new_n17783_));
  AND2X1   g15347(.A(new_n17779_), .B(pi0625), .Y(new_n17784_));
  OAI21X1  g15348(.A0(new_n17720_), .A1(pi0625), .B0(pi1153), .Y(new_n17785_));
  OR2X1    g15349(.A(new_n17785_), .B(new_n17784_), .Y(new_n17786_));
  NAND3X1  g15350(.A(new_n17786_), .B(new_n17689_), .C(pi0608), .Y(new_n17787_));
  NAND2X1  g15351(.A(new_n17787_), .B(new_n17783_), .Y(new_n17788_));
  MX2X1    g15352(.A(new_n17788_), .B(new_n17779_), .S0(new_n11769_), .Y(new_n17789_));
  INVX1    g15353(.A(new_n17691_), .Y(new_n17790_));
  OAI21X1  g15354(.A0(new_n17790_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n17791_));
  AOI21X1  g15355(.A0(new_n17789_), .A1(new_n12462_), .B0(new_n17791_), .Y(new_n17792_));
  OAI21X1  g15356(.A0(new_n17723_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n17793_));
  OAI21X1  g15357(.A0(new_n17790_), .A1(pi0609), .B0(pi1155), .Y(new_n17794_));
  AOI21X1  g15358(.A0(new_n17789_), .A1(pi0609), .B0(new_n17794_), .Y(new_n17795_));
  OAI21X1  g15359(.A0(new_n17724_), .A1(pi1155), .B0(pi0660), .Y(new_n17796_));
  OAI22X1  g15360(.A0(new_n17796_), .A1(new_n17795_), .B0(new_n17793_), .B1(new_n17792_), .Y(new_n17797_));
  MX2X1    g15361(.A(new_n17797_), .B(new_n17789_), .S0(new_n11768_), .Y(new_n17798_));
  OAI21X1  g15362(.A0(new_n17693_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17799_));
  AOI21X1  g15363(.A0(new_n17798_), .A1(new_n12486_), .B0(new_n17799_), .Y(new_n17800_));
  OR2X1    g15364(.A(new_n17728_), .B(pi0627), .Y(new_n17801_));
  OAI21X1  g15365(.A0(new_n17693_), .A1(pi0618), .B0(pi1154), .Y(new_n17802_));
  AOI21X1  g15366(.A0(new_n17798_), .A1(pi0618), .B0(new_n17802_), .Y(new_n17803_));
  OR2X1    g15367(.A(new_n17730_), .B(new_n12494_), .Y(new_n17804_));
  OAI22X1  g15368(.A0(new_n17804_), .A1(new_n17803_), .B0(new_n17801_), .B1(new_n17800_), .Y(new_n17805_));
  MX2X1    g15369(.A(new_n17805_), .B(new_n17798_), .S0(new_n11767_), .Y(new_n17806_));
  NAND2X1  g15370(.A(new_n17806_), .B(new_n12509_), .Y(new_n17807_));
  AOI21X1  g15371(.A0(new_n17695_), .A1(pi0619), .B0(pi1159), .Y(new_n17808_));
  OR2X1    g15372(.A(new_n17734_), .B(pi0648), .Y(new_n17809_));
  AOI21X1  g15373(.A0(new_n17808_), .A1(new_n17807_), .B0(new_n17809_), .Y(new_n17810_));
  NAND2X1  g15374(.A(new_n17806_), .B(pi0619), .Y(new_n17811_));
  AOI21X1  g15375(.A0(new_n17695_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n17812_));
  OR2X1    g15376(.A(new_n17736_), .B(new_n12517_), .Y(new_n17813_));
  AOI21X1  g15377(.A0(new_n17812_), .A1(new_n17811_), .B0(new_n17813_), .Y(new_n17814_));
  NOR3X1   g15378(.A(new_n17814_), .B(new_n17810_), .C(new_n11766_), .Y(new_n17815_));
  OAI21X1  g15379(.A0(new_n17806_), .A1(pi0789), .B0(new_n12709_), .Y(new_n17816_));
  AOI21X1  g15380(.A0(new_n17678_), .A1(pi0626), .B0(new_n16218_), .Y(new_n17817_));
  OAI21X1  g15381(.A0(new_n17738_), .A1(pi0626), .B0(new_n17817_), .Y(new_n17818_));
  AOI21X1  g15382(.A0(new_n17678_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n17819_));
  OAI21X1  g15383(.A0(new_n17738_), .A1(new_n12542_), .B0(new_n17819_), .Y(new_n17820_));
  NAND2X1  g15384(.A(new_n17696_), .B(new_n12637_), .Y(new_n17821_));
  NAND3X1  g15385(.A(new_n17821_), .B(new_n17820_), .C(new_n17818_), .Y(new_n17822_));
  AOI21X1  g15386(.A0(new_n17822_), .A1(pi0788), .B0(new_n14125_), .Y(new_n17823_));
  OAI21X1  g15387(.A0(new_n17816_), .A1(new_n17815_), .B0(new_n17823_), .Y(new_n17824_));
  AOI21X1  g15388(.A0(new_n17824_), .A1(new_n17758_), .B0(new_n14121_), .Y(new_n17825_));
  OR2X1    g15389(.A(new_n17742_), .B(new_n14239_), .Y(new_n17826_));
  OR2X1    g15390(.A(new_n17705_), .B(new_n14244_), .Y(new_n17827_));
  OR2X1    g15391(.A(new_n17706_), .B(new_n14242_), .Y(new_n17828_));
  NAND3X1  g15392(.A(new_n17828_), .B(new_n17827_), .C(new_n17826_), .Y(new_n17829_));
  AOI21X1  g15393(.A0(new_n17829_), .A1(pi0787), .B0(new_n17825_), .Y(new_n17830_));
  AOI22X1  g15394(.A0(new_n17830_), .A1(new_n17754_), .B0(new_n17751_), .B1(pi0790), .Y(new_n17831_));
  OR2X1    g15395(.A(new_n17831_), .B(po1038), .Y(new_n17832_));
  AOI21X1  g15396(.A0(po1038), .A1(new_n5203_), .B0(pi0832), .Y(new_n17833_));
  AOI22X1  g15397(.A0(new_n17833_), .A1(new_n17832_), .B0(new_n17676_), .B1(new_n17675_), .Y(po0337));
  AOI21X1  g15398(.A0(pi1093), .A1(pi1092), .B0(pi0181), .Y(new_n17835_));
  INVX1    g15399(.A(new_n17835_), .Y(new_n17836_));
  AOI21X1  g15400(.A0(new_n12056_), .A1(new_n15037_), .B0(new_n17835_), .Y(new_n17837_));
  INVX1    g15401(.A(new_n17837_), .Y(new_n17838_));
  NAND2X1  g15402(.A(new_n17838_), .B(new_n15771_), .Y(new_n17839_));
  AND3X1   g15403(.A(new_n12480_), .B(new_n12056_), .C(new_n15037_), .Y(new_n17840_));
  OAI21X1  g15404(.A0(new_n17840_), .A1(new_n17839_), .B0(pi1155), .Y(new_n17841_));
  NOR3X1   g15405(.A(new_n17840_), .B(new_n17835_), .C(pi1155), .Y(new_n17842_));
  INVX1    g15406(.A(new_n17842_), .Y(new_n17843_));
  AOI21X1  g15407(.A0(new_n17843_), .A1(new_n17841_), .B0(new_n11768_), .Y(new_n17844_));
  AOI21X1  g15408(.A0(new_n17839_), .A1(new_n11768_), .B0(new_n17844_), .Y(new_n17845_));
  AOI21X1  g15409(.A0(new_n17845_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n17846_));
  AOI21X1  g15410(.A0(new_n17845_), .A1(new_n12655_), .B0(pi1154), .Y(new_n17847_));
  NOR2X1   g15411(.A(new_n17847_), .B(new_n17846_), .Y(new_n17848_));
  MX2X1    g15412(.A(new_n17848_), .B(new_n17845_), .S0(new_n11767_), .Y(new_n17849_));
  NOR2X1   g15413(.A(new_n17849_), .B(pi0789), .Y(new_n17850_));
  AOI21X1  g15414(.A0(new_n17849_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n17851_));
  AOI21X1  g15415(.A0(new_n17849_), .A1(new_n15790_), .B0(pi1159), .Y(new_n17852_));
  OR2X1    g15416(.A(new_n17852_), .B(new_n17851_), .Y(new_n17853_));
  AOI21X1  g15417(.A0(new_n17853_), .A1(pi0789), .B0(new_n17850_), .Y(new_n17854_));
  INVX1    g15418(.A(new_n17854_), .Y(new_n17855_));
  MX2X1    g15419(.A(new_n17855_), .B(new_n17836_), .S0(new_n12708_), .Y(new_n17856_));
  MX2X1    g15420(.A(new_n17856_), .B(new_n17836_), .S0(new_n12580_), .Y(new_n17857_));
  AOI21X1  g15421(.A0(new_n12439_), .A1(new_n15056_), .B0(new_n17835_), .Y(new_n17858_));
  OR2X1    g15422(.A(new_n17858_), .B(pi0778), .Y(new_n17859_));
  INVX1    g15423(.A(new_n17858_), .Y(new_n17860_));
  AND3X1   g15424(.A(new_n12439_), .B(new_n15056_), .C(new_n12363_), .Y(new_n17861_));
  INVX1    g15425(.A(new_n17861_), .Y(new_n17862_));
  AOI21X1  g15426(.A0(new_n17862_), .A1(new_n17860_), .B0(new_n12364_), .Y(new_n17863_));
  NOR3X1   g15427(.A(new_n17861_), .B(new_n17835_), .C(pi1153), .Y(new_n17864_));
  OR3X1    g15428(.A(new_n17864_), .B(new_n17863_), .C(new_n11769_), .Y(new_n17865_));
  AND2X1   g15429(.A(new_n17865_), .B(new_n17859_), .Y(new_n17866_));
  NOR4X1   g15430(.A(new_n17866_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n17867_));
  AND3X1   g15431(.A(new_n17867_), .B(new_n12739_), .C(new_n12718_), .Y(new_n17868_));
  INVX1    g15432(.A(new_n17868_), .Y(new_n17869_));
  AOI21X1  g15433(.A0(new_n17835_), .A1(pi0647), .B0(pi1157), .Y(new_n17870_));
  OAI21X1  g15434(.A0(new_n17869_), .A1(pi0647), .B0(new_n17870_), .Y(new_n17871_));
  MX2X1    g15435(.A(new_n17868_), .B(new_n17835_), .S0(new_n12577_), .Y(new_n17872_));
  OAI22X1  g15436(.A0(new_n17872_), .A1(new_n14242_), .B0(new_n17871_), .B1(new_n12592_), .Y(new_n17873_));
  AOI21X1  g15437(.A0(new_n17857_), .A1(new_n14326_), .B0(new_n17873_), .Y(new_n17874_));
  NOR2X1   g15438(.A(new_n17874_), .B(new_n11763_), .Y(new_n17875_));
  AOI21X1  g15439(.A0(new_n17836_), .A1(pi0626), .B0(new_n16218_), .Y(new_n17876_));
  OAI21X1  g15440(.A0(new_n17854_), .A1(pi0626), .B0(new_n17876_), .Y(new_n17877_));
  AOI21X1  g15441(.A0(new_n17836_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n17878_));
  OAI21X1  g15442(.A0(new_n17854_), .A1(new_n12542_), .B0(new_n17878_), .Y(new_n17879_));
  NAND2X1  g15443(.A(new_n17867_), .B(new_n12637_), .Y(new_n17880_));
  AND3X1   g15444(.A(new_n17880_), .B(new_n17879_), .C(new_n17877_), .Y(new_n17881_));
  NOR2X1   g15445(.A(new_n17881_), .B(new_n11765_), .Y(new_n17882_));
  NOR2X1   g15446(.A(new_n17835_), .B(pi1153), .Y(new_n17883_));
  NOR3X1   g15447(.A(new_n17858_), .B(new_n11991_), .C(new_n12363_), .Y(new_n17884_));
  AOI21X1  g15448(.A0(new_n17860_), .A1(new_n12048_), .B0(new_n17838_), .Y(new_n17885_));
  OAI21X1  g15449(.A0(new_n17885_), .A1(new_n17884_), .B0(new_n17883_), .Y(new_n17886_));
  NOR2X1   g15450(.A(new_n17863_), .B(pi0608), .Y(new_n17887_));
  NOR3X1   g15451(.A(new_n17884_), .B(new_n17838_), .C(new_n12364_), .Y(new_n17888_));
  NOR3X1   g15452(.A(new_n17888_), .B(new_n17864_), .C(new_n12368_), .Y(new_n17889_));
  AOI21X1  g15453(.A0(new_n17887_), .A1(new_n17886_), .B0(new_n17889_), .Y(new_n17890_));
  OR2X1    g15454(.A(new_n17885_), .B(pi0778), .Y(new_n17891_));
  OAI21X1  g15455(.A0(new_n17890_), .A1(new_n11769_), .B0(new_n17891_), .Y(new_n17892_));
  INVX1    g15456(.A(new_n17892_), .Y(new_n17893_));
  AND2X1   g15457(.A(new_n17892_), .B(new_n12462_), .Y(new_n17894_));
  OAI21X1  g15458(.A0(new_n17866_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n17895_));
  OR2X1    g15459(.A(new_n17895_), .B(new_n17894_), .Y(new_n17896_));
  AND3X1   g15460(.A(new_n17896_), .B(new_n17841_), .C(new_n12468_), .Y(new_n17897_));
  OAI21X1  g15461(.A0(new_n17866_), .A1(pi0609), .B0(pi1155), .Y(new_n17898_));
  AOI21X1  g15462(.A0(new_n17892_), .A1(pi0609), .B0(new_n17898_), .Y(new_n17899_));
  NOR3X1   g15463(.A(new_n17899_), .B(new_n17842_), .C(new_n12468_), .Y(new_n17900_));
  NOR2X1   g15464(.A(new_n17900_), .B(new_n17897_), .Y(new_n17901_));
  MX2X1    g15465(.A(new_n17901_), .B(new_n17893_), .S0(new_n11768_), .Y(new_n17902_));
  AOI21X1  g15466(.A0(new_n17865_), .A1(new_n17859_), .B0(new_n12630_), .Y(new_n17903_));
  AOI21X1  g15467(.A0(new_n17903_), .A1(pi0618), .B0(pi1154), .Y(new_n17904_));
  OAI21X1  g15468(.A0(new_n17902_), .A1(pi0618), .B0(new_n17904_), .Y(new_n17905_));
  NOR2X1   g15469(.A(new_n17846_), .B(pi0627), .Y(new_n17906_));
  AOI21X1  g15470(.A0(new_n17903_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n17907_));
  OAI21X1  g15471(.A0(new_n17902_), .A1(new_n12486_), .B0(new_n17907_), .Y(new_n17908_));
  NOR2X1   g15472(.A(new_n17847_), .B(new_n12494_), .Y(new_n17909_));
  AOI22X1  g15473(.A0(new_n17909_), .A1(new_n17908_), .B0(new_n17906_), .B1(new_n17905_), .Y(new_n17910_));
  MX2X1    g15474(.A(new_n17910_), .B(new_n17902_), .S0(new_n11767_), .Y(new_n17911_));
  OR4X1    g15475(.A(new_n17866_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n17912_));
  AND2X1   g15476(.A(new_n17912_), .B(new_n12510_), .Y(new_n17913_));
  OAI21X1  g15477(.A0(new_n17911_), .A1(pi0619), .B0(new_n17913_), .Y(new_n17914_));
  NOR2X1   g15478(.A(new_n17851_), .B(pi0648), .Y(new_n17915_));
  AND2X1   g15479(.A(new_n17915_), .B(new_n17914_), .Y(new_n17916_));
  NOR4X1   g15480(.A(new_n17866_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n17917_));
  NOR2X1   g15481(.A(new_n17917_), .B(new_n12510_), .Y(new_n17918_));
  OAI21X1  g15482(.A0(new_n17911_), .A1(new_n12509_), .B0(new_n17918_), .Y(new_n17919_));
  NOR2X1   g15483(.A(new_n17852_), .B(new_n12517_), .Y(new_n17920_));
  AND2X1   g15484(.A(new_n17920_), .B(new_n17919_), .Y(new_n17921_));
  OR3X1    g15485(.A(new_n17921_), .B(new_n17916_), .C(new_n11766_), .Y(new_n17922_));
  AOI21X1  g15486(.A0(new_n17911_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n17923_));
  AOI21X1  g15487(.A0(new_n17923_), .A1(new_n17922_), .B0(new_n17882_), .Y(new_n17924_));
  OR2X1    g15488(.A(new_n17924_), .B(new_n14125_), .Y(new_n17925_));
  INVX1    g15489(.A(new_n17856_), .Y(new_n17926_));
  AND2X1   g15490(.A(new_n17867_), .B(new_n12718_), .Y(new_n17927_));
  AOI22X1  g15491(.A0(new_n17927_), .A1(new_n14426_), .B0(new_n17926_), .B1(new_n12735_), .Y(new_n17928_));
  AOI22X1  g15492(.A0(new_n17927_), .A1(new_n14428_), .B0(new_n17926_), .B1(new_n12733_), .Y(new_n17929_));
  MX2X1    g15493(.A(new_n17929_), .B(new_n17928_), .S0(new_n12561_), .Y(new_n17930_));
  OAI21X1  g15494(.A0(new_n17930_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n17931_));
  INVX1    g15495(.A(new_n17931_), .Y(new_n17932_));
  AOI21X1  g15496(.A0(new_n17932_), .A1(new_n17925_), .B0(new_n17875_), .Y(new_n17933_));
  OAI21X1  g15497(.A0(new_n17872_), .A1(new_n12578_), .B0(new_n17871_), .Y(new_n17934_));
  MX2X1    g15498(.A(new_n17934_), .B(new_n17869_), .S0(new_n11763_), .Y(new_n17935_));
  OAI21X1  g15499(.A0(new_n17935_), .A1(pi0644), .B0(pi0715), .Y(new_n17936_));
  AOI21X1  g15500(.A0(new_n17933_), .A1(pi0644), .B0(new_n17936_), .Y(new_n17937_));
  OR3X1    g15501(.A(new_n17836_), .B(new_n12603_), .C(new_n11763_), .Y(new_n17938_));
  OAI21X1  g15502(.A0(new_n17857_), .A1(new_n12604_), .B0(new_n17938_), .Y(new_n17939_));
  OAI21X1  g15503(.A0(new_n17836_), .A1(pi0644), .B0(new_n12608_), .Y(new_n17940_));
  AOI21X1  g15504(.A0(new_n17939_), .A1(pi0644), .B0(new_n17940_), .Y(new_n17941_));
  OR2X1    g15505(.A(new_n17941_), .B(new_n11762_), .Y(new_n17942_));
  OAI21X1  g15506(.A0(new_n17935_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17943_));
  AOI21X1  g15507(.A0(new_n17933_), .A1(new_n12612_), .B0(new_n17943_), .Y(new_n17944_));
  OAI21X1  g15508(.A0(new_n17836_), .A1(new_n12612_), .B0(pi0715), .Y(new_n17945_));
  AOI21X1  g15509(.A0(new_n17939_), .A1(new_n12612_), .B0(new_n17945_), .Y(new_n17946_));
  OR2X1    g15510(.A(new_n17946_), .B(pi1160), .Y(new_n17947_));
  OAI22X1  g15511(.A0(new_n17947_), .A1(new_n17944_), .B0(new_n17942_), .B1(new_n17937_), .Y(new_n17948_));
  NAND2X1  g15512(.A(new_n17948_), .B(pi0790), .Y(new_n17949_));
  AOI21X1  g15513(.A0(new_n17933_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n17950_));
  AOI21X1  g15514(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0181), .Y(new_n17951_));
  INVX1    g15515(.A(new_n17951_), .Y(new_n17952_));
  AOI21X1  g15516(.A0(new_n3103_), .A1(new_n15056_), .B0(new_n17952_), .Y(new_n17953_));
  OAI21X1  g15517(.A0(new_n12826_), .A1(new_n5204_), .B0(new_n2979_), .Y(new_n17954_));
  AOI22X1  g15518(.A0(new_n17954_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n5204_), .Y(new_n17955_));
  AOI21X1  g15519(.A0(new_n12771_), .A1(new_n5204_), .B0(new_n12441_), .Y(new_n17956_));
  NOR3X1   g15520(.A(new_n17956_), .B(new_n17955_), .C(pi0709), .Y(new_n17957_));
  NOR2X1   g15521(.A(new_n17957_), .B(new_n17953_), .Y(new_n17958_));
  INVX1    g15522(.A(new_n17958_), .Y(new_n17959_));
  AOI21X1  g15523(.A0(new_n17951_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n17960_));
  OAI21X1  g15524(.A0(new_n17958_), .A1(new_n12363_), .B0(new_n17960_), .Y(new_n17961_));
  AOI21X1  g15525(.A0(new_n17951_), .A1(pi0625), .B0(pi1153), .Y(new_n17962_));
  OAI21X1  g15526(.A0(new_n17958_), .A1(pi0625), .B0(new_n17962_), .Y(new_n17963_));
  AND2X1   g15527(.A(new_n17963_), .B(new_n17961_), .Y(new_n17964_));
  MX2X1    g15528(.A(new_n17964_), .B(new_n17959_), .S0(new_n11769_), .Y(new_n17965_));
  MX2X1    g15529(.A(new_n17965_), .B(new_n17951_), .S0(new_n12490_), .Y(new_n17966_));
  INVX1    g15530(.A(new_n17966_), .Y(new_n17967_));
  MX2X1    g15531(.A(new_n17967_), .B(new_n17952_), .S0(new_n12513_), .Y(new_n17968_));
  INVX1    g15532(.A(new_n17968_), .Y(new_n17969_));
  MX2X1    g15533(.A(new_n17969_), .B(new_n17951_), .S0(new_n12531_), .Y(new_n17970_));
  MX2X1    g15534(.A(new_n17970_), .B(new_n17951_), .S0(new_n12563_), .Y(new_n17971_));
  INVX1    g15535(.A(new_n17971_), .Y(new_n17972_));
  AOI21X1  g15536(.A0(new_n17951_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n17973_));
  OAI21X1  g15537(.A0(new_n17972_), .A1(new_n12554_), .B0(new_n17973_), .Y(new_n17974_));
  AOI21X1  g15538(.A0(new_n17951_), .A1(pi0628), .B0(pi1156), .Y(new_n17975_));
  OAI21X1  g15539(.A0(new_n17972_), .A1(pi0628), .B0(new_n17975_), .Y(new_n17976_));
  AOI21X1  g15540(.A0(new_n17976_), .A1(new_n17974_), .B0(new_n11764_), .Y(new_n17977_));
  AOI21X1  g15541(.A0(new_n17972_), .A1(new_n11764_), .B0(new_n17977_), .Y(new_n17978_));
  MX2X1    g15542(.A(new_n17978_), .B(new_n17951_), .S0(pi0647), .Y(new_n17979_));
  MX2X1    g15543(.A(new_n17978_), .B(new_n17951_), .S0(new_n12577_), .Y(new_n17980_));
  MX2X1    g15544(.A(new_n17980_), .B(new_n17979_), .S0(new_n12578_), .Y(new_n17981_));
  MX2X1    g15545(.A(new_n17981_), .B(new_n17978_), .S0(new_n11763_), .Y(new_n17982_));
  AOI21X1  g15546(.A0(new_n17982_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n17983_));
  AOI22X1  g15547(.A0(new_n12073_), .A1(pi0181), .B0(new_n12444_), .B1(pi0754), .Y(new_n17984_));
  OR3X1    g15548(.A(new_n12776_), .B(pi0754), .C(pi0181), .Y(new_n17985_));
  OAI22X1  g15549(.A0(new_n12045_), .A1(new_n5204_), .B0(new_n11822_), .B1(new_n15037_), .Y(new_n17986_));
  AOI22X1  g15550(.A0(new_n17986_), .A1(new_n2939_), .B0(pi0754), .B1(pi0181), .Y(new_n17987_));
  AND2X1   g15551(.A(new_n17987_), .B(new_n17985_), .Y(new_n17988_));
  OAI21X1  g15552(.A0(new_n17984_), .A1(new_n2939_), .B0(new_n17988_), .Y(new_n17989_));
  AND2X1   g15553(.A(new_n17989_), .B(new_n2979_), .Y(new_n17990_));
  OAI21X1  g15554(.A0(new_n12077_), .A1(pi0181), .B0(pi0038), .Y(new_n17991_));
  AOI21X1  g15555(.A0(new_n12079_), .A1(new_n15037_), .B0(new_n17991_), .Y(new_n17992_));
  OR2X1    g15556(.A(new_n17992_), .B(new_n17990_), .Y(new_n17993_));
  MX2X1    g15557(.A(new_n17993_), .B(pi0181), .S0(new_n11770_), .Y(new_n17994_));
  AND2X1   g15558(.A(new_n17994_), .B(new_n12474_), .Y(new_n17995_));
  AOI21X1  g15559(.A0(new_n17952_), .A1(new_n12473_), .B0(new_n17995_), .Y(new_n17996_));
  AOI22X1  g15560(.A0(new_n17995_), .A1(pi0609), .B0(new_n17952_), .B1(new_n12472_), .Y(new_n17997_));
  AOI22X1  g15561(.A0(new_n17995_), .A1(new_n12462_), .B0(new_n17952_), .B1(new_n12481_), .Y(new_n17998_));
  MX2X1    g15562(.A(new_n17998_), .B(new_n17997_), .S0(pi1155), .Y(new_n17999_));
  MX2X1    g15563(.A(new_n17999_), .B(new_n17996_), .S0(new_n11768_), .Y(new_n18000_));
  OAI21X1  g15564(.A0(new_n17952_), .A1(pi0618), .B0(pi1154), .Y(new_n18001_));
  AOI21X1  g15565(.A0(new_n18000_), .A1(pi0618), .B0(new_n18001_), .Y(new_n18002_));
  OAI21X1  g15566(.A0(new_n17952_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18003_));
  AOI21X1  g15567(.A0(new_n18000_), .A1(new_n12486_), .B0(new_n18003_), .Y(new_n18004_));
  NOR2X1   g15568(.A(new_n18004_), .B(new_n18002_), .Y(new_n18005_));
  MX2X1    g15569(.A(new_n18005_), .B(new_n18000_), .S0(new_n11767_), .Y(new_n18006_));
  OAI21X1  g15570(.A0(new_n17952_), .A1(pi0619), .B0(pi1159), .Y(new_n18007_));
  AOI21X1  g15571(.A0(new_n18006_), .A1(pi0619), .B0(new_n18007_), .Y(new_n18008_));
  OAI21X1  g15572(.A0(new_n17952_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n18009_));
  AOI21X1  g15573(.A0(new_n18006_), .A1(new_n12509_), .B0(new_n18009_), .Y(new_n18010_));
  NOR2X1   g15574(.A(new_n18010_), .B(new_n18008_), .Y(new_n18011_));
  MX2X1    g15575(.A(new_n18011_), .B(new_n18006_), .S0(new_n11766_), .Y(new_n18012_));
  AND2X1   g15576(.A(new_n17951_), .B(new_n12708_), .Y(new_n18013_));
  AOI21X1  g15577(.A0(new_n18012_), .A1(new_n16140_), .B0(new_n18013_), .Y(new_n18014_));
  NAND2X1  g15578(.A(new_n17951_), .B(new_n12580_), .Y(new_n18015_));
  OAI21X1  g15579(.A0(new_n18014_), .A1(new_n12580_), .B0(new_n18015_), .Y(new_n18016_));
  MX2X1    g15580(.A(new_n18016_), .B(new_n17951_), .S0(new_n12604_), .Y(new_n18017_));
  OAI21X1  g15581(.A0(new_n17952_), .A1(pi0644), .B0(new_n12608_), .Y(new_n18018_));
  AOI21X1  g15582(.A0(new_n18017_), .A1(pi0644), .B0(new_n18018_), .Y(new_n18019_));
  OR2X1    g15583(.A(new_n18019_), .B(new_n11762_), .Y(new_n18020_));
  AOI21X1  g15584(.A0(new_n17982_), .A1(pi0644), .B0(pi0715), .Y(new_n18021_));
  OAI21X1  g15585(.A0(new_n17952_), .A1(new_n12612_), .B0(pi0715), .Y(new_n18022_));
  AOI21X1  g15586(.A0(new_n18017_), .A1(new_n12612_), .B0(new_n18022_), .Y(new_n18023_));
  OR2X1    g15587(.A(new_n18023_), .B(pi1160), .Y(new_n18024_));
  OAI22X1  g15588(.A0(new_n18024_), .A1(new_n18021_), .B0(new_n18020_), .B1(new_n17983_), .Y(new_n18025_));
  OR3X1    g15589(.A(new_n18023_), .B(pi1160), .C(pi0644), .Y(new_n18026_));
  OR3X1    g15590(.A(new_n18019_), .B(new_n11762_), .C(new_n12612_), .Y(new_n18027_));
  NAND3X1  g15591(.A(new_n18027_), .B(new_n18026_), .C(pi0790), .Y(new_n18028_));
  NAND2X1  g15592(.A(new_n18014_), .B(new_n14249_), .Y(new_n18029_));
  MX2X1    g15593(.A(new_n17976_), .B(new_n17974_), .S0(new_n12561_), .Y(new_n18030_));
  AND2X1   g15594(.A(new_n18030_), .B(new_n18029_), .Y(new_n18031_));
  OR2X1    g15595(.A(new_n18031_), .B(new_n11764_), .Y(new_n18032_));
  OR3X1    g15596(.A(new_n17992_), .B(new_n17990_), .C(new_n15056_), .Y(new_n18033_));
  OAI21X1  g15597(.A0(new_n12213_), .A1(new_n5204_), .B0(pi0754), .Y(new_n18034_));
  AOI21X1  g15598(.A0(new_n12155_), .A1(new_n5204_), .B0(new_n18034_), .Y(new_n18035_));
  AOI21X1  g15599(.A0(new_n12788_), .A1(new_n5204_), .B0(pi0754), .Y(new_n18036_));
  OAI21X1  g15600(.A0(new_n12787_), .A1(new_n5204_), .B0(new_n18036_), .Y(new_n18037_));
  NAND2X1  g15601(.A(new_n18037_), .B(pi0039), .Y(new_n18038_));
  AND2X1   g15602(.A(new_n12332_), .B(pi0181), .Y(new_n18039_));
  OAI21X1  g15603(.A0(new_n12315_), .A1(pi0181), .B0(pi0754), .Y(new_n18040_));
  NOR4X1   g15604(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0181), .Y(new_n18041_));
  OAI21X1  g15605(.A0(new_n12800_), .A1(new_n5204_), .B0(new_n15037_), .Y(new_n18042_));
  OAI22X1  g15606(.A0(new_n18042_), .A1(new_n18041_), .B0(new_n18040_), .B1(new_n18039_), .Y(new_n18043_));
  AOI21X1  g15607(.A0(new_n18043_), .A1(new_n2939_), .B0(pi0038), .Y(new_n18044_));
  OAI21X1  g15608(.A0(new_n18038_), .A1(new_n18035_), .B0(new_n18044_), .Y(new_n18045_));
  OAI21X1  g15609(.A0(new_n12276_), .A1(pi0754), .B0(new_n13540_), .Y(new_n18046_));
  NAND2X1  g15610(.A(new_n18046_), .B(new_n5204_), .Y(new_n18047_));
  AOI21X1  g15611(.A0(new_n12056_), .A1(new_n15037_), .B0(new_n13443_), .Y(new_n18048_));
  NOR2X1   g15612(.A(new_n18048_), .B(new_n5204_), .Y(new_n18049_));
  AOI21X1  g15613(.A0(new_n18049_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n18050_));
  AOI21X1  g15614(.A0(new_n18050_), .A1(new_n18047_), .B0(pi0709), .Y(new_n18051_));
  AOI21X1  g15615(.A0(new_n18051_), .A1(new_n18045_), .B0(new_n11770_), .Y(new_n18052_));
  AOI22X1  g15616(.A0(new_n18052_), .A1(new_n18033_), .B0(new_n11770_), .B1(pi0181), .Y(new_n18053_));
  AND2X1   g15617(.A(new_n18053_), .B(new_n12363_), .Y(new_n18054_));
  OAI21X1  g15618(.A0(new_n17994_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n18055_));
  OR2X1    g15619(.A(new_n18055_), .B(new_n18054_), .Y(new_n18056_));
  NAND3X1  g15620(.A(new_n18056_), .B(new_n17961_), .C(new_n12368_), .Y(new_n18057_));
  AND2X1   g15621(.A(new_n18053_), .B(pi0625), .Y(new_n18058_));
  OAI21X1  g15622(.A0(new_n17994_), .A1(pi0625), .B0(pi1153), .Y(new_n18059_));
  OR2X1    g15623(.A(new_n18059_), .B(new_n18058_), .Y(new_n18060_));
  NAND3X1  g15624(.A(new_n18060_), .B(new_n17963_), .C(pi0608), .Y(new_n18061_));
  NAND2X1  g15625(.A(new_n18061_), .B(new_n18057_), .Y(new_n18062_));
  MX2X1    g15626(.A(new_n18062_), .B(new_n18053_), .S0(new_n11769_), .Y(new_n18063_));
  INVX1    g15627(.A(new_n17965_), .Y(new_n18064_));
  OAI21X1  g15628(.A0(new_n18064_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n18065_));
  AOI21X1  g15629(.A0(new_n18063_), .A1(new_n12462_), .B0(new_n18065_), .Y(new_n18066_));
  OAI21X1  g15630(.A0(new_n17997_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n18067_));
  OAI21X1  g15631(.A0(new_n18064_), .A1(pi0609), .B0(pi1155), .Y(new_n18068_));
  AOI21X1  g15632(.A0(new_n18063_), .A1(pi0609), .B0(new_n18068_), .Y(new_n18069_));
  OAI21X1  g15633(.A0(new_n17998_), .A1(pi1155), .B0(pi0660), .Y(new_n18070_));
  OAI22X1  g15634(.A0(new_n18070_), .A1(new_n18069_), .B0(new_n18067_), .B1(new_n18066_), .Y(new_n18071_));
  MX2X1    g15635(.A(new_n18071_), .B(new_n18063_), .S0(new_n11768_), .Y(new_n18072_));
  OAI21X1  g15636(.A0(new_n17967_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18073_));
  AOI21X1  g15637(.A0(new_n18072_), .A1(new_n12486_), .B0(new_n18073_), .Y(new_n18074_));
  OR2X1    g15638(.A(new_n18002_), .B(pi0627), .Y(new_n18075_));
  OAI21X1  g15639(.A0(new_n17967_), .A1(pi0618), .B0(pi1154), .Y(new_n18076_));
  AOI21X1  g15640(.A0(new_n18072_), .A1(pi0618), .B0(new_n18076_), .Y(new_n18077_));
  OR2X1    g15641(.A(new_n18004_), .B(new_n12494_), .Y(new_n18078_));
  OAI22X1  g15642(.A0(new_n18078_), .A1(new_n18077_), .B0(new_n18075_), .B1(new_n18074_), .Y(new_n18079_));
  MX2X1    g15643(.A(new_n18079_), .B(new_n18072_), .S0(new_n11767_), .Y(new_n18080_));
  NAND2X1  g15644(.A(new_n18080_), .B(new_n12509_), .Y(new_n18081_));
  AOI21X1  g15645(.A0(new_n17969_), .A1(pi0619), .B0(pi1159), .Y(new_n18082_));
  OR2X1    g15646(.A(new_n18008_), .B(pi0648), .Y(new_n18083_));
  AOI21X1  g15647(.A0(new_n18082_), .A1(new_n18081_), .B0(new_n18083_), .Y(new_n18084_));
  NAND2X1  g15648(.A(new_n18080_), .B(pi0619), .Y(new_n18085_));
  AOI21X1  g15649(.A0(new_n17969_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n18086_));
  OR2X1    g15650(.A(new_n18010_), .B(new_n12517_), .Y(new_n18087_));
  AOI21X1  g15651(.A0(new_n18086_), .A1(new_n18085_), .B0(new_n18087_), .Y(new_n18088_));
  NOR3X1   g15652(.A(new_n18088_), .B(new_n18084_), .C(new_n11766_), .Y(new_n18089_));
  OAI21X1  g15653(.A0(new_n18080_), .A1(pi0789), .B0(new_n12709_), .Y(new_n18090_));
  AOI21X1  g15654(.A0(new_n17952_), .A1(pi0626), .B0(new_n16218_), .Y(new_n18091_));
  OAI21X1  g15655(.A0(new_n18012_), .A1(pi0626), .B0(new_n18091_), .Y(new_n18092_));
  AOI21X1  g15656(.A0(new_n17952_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n18093_));
  OAI21X1  g15657(.A0(new_n18012_), .A1(new_n12542_), .B0(new_n18093_), .Y(new_n18094_));
  NAND2X1  g15658(.A(new_n17970_), .B(new_n12637_), .Y(new_n18095_));
  NAND3X1  g15659(.A(new_n18095_), .B(new_n18094_), .C(new_n18092_), .Y(new_n18096_));
  AOI21X1  g15660(.A0(new_n18096_), .A1(pi0788), .B0(new_n14125_), .Y(new_n18097_));
  OAI21X1  g15661(.A0(new_n18090_), .A1(new_n18089_), .B0(new_n18097_), .Y(new_n18098_));
  AOI21X1  g15662(.A0(new_n18098_), .A1(new_n18032_), .B0(new_n14121_), .Y(new_n18099_));
  OR2X1    g15663(.A(new_n18016_), .B(new_n14239_), .Y(new_n18100_));
  OR2X1    g15664(.A(new_n17979_), .B(new_n14244_), .Y(new_n18101_));
  OR2X1    g15665(.A(new_n17980_), .B(new_n14242_), .Y(new_n18102_));
  NAND3X1  g15666(.A(new_n18102_), .B(new_n18101_), .C(new_n18100_), .Y(new_n18103_));
  AOI21X1  g15667(.A0(new_n18103_), .A1(pi0787), .B0(new_n18099_), .Y(new_n18104_));
  AOI22X1  g15668(.A0(new_n18104_), .A1(new_n18028_), .B0(new_n18025_), .B1(pi0790), .Y(new_n18105_));
  OR2X1    g15669(.A(new_n18105_), .B(po1038), .Y(new_n18106_));
  AOI21X1  g15670(.A0(po1038), .A1(new_n5204_), .B0(pi0832), .Y(new_n18107_));
  AOI22X1  g15671(.A0(new_n18107_), .A1(new_n18106_), .B0(new_n17950_), .B1(new_n17949_), .Y(po0338));
  AOI21X1  g15672(.A0(pi1093), .A1(pi1092), .B0(pi0182), .Y(new_n18109_));
  INVX1    g15673(.A(new_n18109_), .Y(new_n18110_));
  AOI21X1  g15674(.A0(new_n12056_), .A1(new_n15068_), .B0(new_n18109_), .Y(new_n18111_));
  INVX1    g15675(.A(new_n18111_), .Y(new_n18112_));
  NAND2X1  g15676(.A(new_n18112_), .B(new_n15771_), .Y(new_n18113_));
  AND3X1   g15677(.A(new_n12480_), .B(new_n12056_), .C(new_n15068_), .Y(new_n18114_));
  OAI21X1  g15678(.A0(new_n18114_), .A1(new_n18113_), .B0(pi1155), .Y(new_n18115_));
  NOR3X1   g15679(.A(new_n18114_), .B(new_n18109_), .C(pi1155), .Y(new_n18116_));
  INVX1    g15680(.A(new_n18116_), .Y(new_n18117_));
  AOI21X1  g15681(.A0(new_n18117_), .A1(new_n18115_), .B0(new_n11768_), .Y(new_n18118_));
  AOI21X1  g15682(.A0(new_n18113_), .A1(new_n11768_), .B0(new_n18118_), .Y(new_n18119_));
  AOI21X1  g15683(.A0(new_n18119_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n18120_));
  AOI21X1  g15684(.A0(new_n18119_), .A1(new_n12655_), .B0(pi1154), .Y(new_n18121_));
  NOR2X1   g15685(.A(new_n18121_), .B(new_n18120_), .Y(new_n18122_));
  MX2X1    g15686(.A(new_n18122_), .B(new_n18119_), .S0(new_n11767_), .Y(new_n18123_));
  NOR2X1   g15687(.A(new_n18123_), .B(pi0789), .Y(new_n18124_));
  AOI21X1  g15688(.A0(new_n18123_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n18125_));
  AOI21X1  g15689(.A0(new_n18123_), .A1(new_n15790_), .B0(pi1159), .Y(new_n18126_));
  OR2X1    g15690(.A(new_n18126_), .B(new_n18125_), .Y(new_n18127_));
  AOI21X1  g15691(.A0(new_n18127_), .A1(pi0789), .B0(new_n18124_), .Y(new_n18128_));
  INVX1    g15692(.A(new_n18128_), .Y(new_n18129_));
  MX2X1    g15693(.A(new_n18129_), .B(new_n18110_), .S0(new_n12708_), .Y(new_n18130_));
  MX2X1    g15694(.A(new_n18130_), .B(new_n18110_), .S0(new_n12580_), .Y(new_n18131_));
  AOI21X1  g15695(.A0(new_n12439_), .A1(new_n15095_), .B0(new_n18109_), .Y(new_n18132_));
  OR2X1    g15696(.A(new_n18132_), .B(pi0778), .Y(new_n18133_));
  INVX1    g15697(.A(new_n18132_), .Y(new_n18134_));
  AND3X1   g15698(.A(new_n12439_), .B(new_n15095_), .C(new_n12363_), .Y(new_n18135_));
  INVX1    g15699(.A(new_n18135_), .Y(new_n18136_));
  AOI21X1  g15700(.A0(new_n18136_), .A1(new_n18134_), .B0(new_n12364_), .Y(new_n18137_));
  NOR3X1   g15701(.A(new_n18135_), .B(new_n18109_), .C(pi1153), .Y(new_n18138_));
  OR3X1    g15702(.A(new_n18138_), .B(new_n18137_), .C(new_n11769_), .Y(new_n18139_));
  AND2X1   g15703(.A(new_n18139_), .B(new_n18133_), .Y(new_n18140_));
  NOR4X1   g15704(.A(new_n18140_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n18141_));
  AND3X1   g15705(.A(new_n18141_), .B(new_n12739_), .C(new_n12718_), .Y(new_n18142_));
  INVX1    g15706(.A(new_n18142_), .Y(new_n18143_));
  AOI21X1  g15707(.A0(new_n18109_), .A1(pi0647), .B0(pi1157), .Y(new_n18144_));
  OAI21X1  g15708(.A0(new_n18143_), .A1(pi0647), .B0(new_n18144_), .Y(new_n18145_));
  MX2X1    g15709(.A(new_n18142_), .B(new_n18109_), .S0(new_n12577_), .Y(new_n18146_));
  OAI22X1  g15710(.A0(new_n18146_), .A1(new_n14242_), .B0(new_n18145_), .B1(new_n12592_), .Y(new_n18147_));
  AOI21X1  g15711(.A0(new_n18131_), .A1(new_n14326_), .B0(new_n18147_), .Y(new_n18148_));
  NOR2X1   g15712(.A(new_n18148_), .B(new_n11763_), .Y(new_n18149_));
  AOI21X1  g15713(.A0(new_n18110_), .A1(pi0626), .B0(new_n16218_), .Y(new_n18150_));
  OAI21X1  g15714(.A0(new_n18128_), .A1(pi0626), .B0(new_n18150_), .Y(new_n18151_));
  AOI21X1  g15715(.A0(new_n18110_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n18152_));
  OAI21X1  g15716(.A0(new_n18128_), .A1(new_n12542_), .B0(new_n18152_), .Y(new_n18153_));
  NAND2X1  g15717(.A(new_n18141_), .B(new_n12637_), .Y(new_n18154_));
  AND3X1   g15718(.A(new_n18154_), .B(new_n18153_), .C(new_n18151_), .Y(new_n18155_));
  NOR2X1   g15719(.A(new_n18155_), .B(new_n11765_), .Y(new_n18156_));
  NOR2X1   g15720(.A(new_n18109_), .B(pi1153), .Y(new_n18157_));
  NOR3X1   g15721(.A(new_n18132_), .B(new_n11991_), .C(new_n12363_), .Y(new_n18158_));
  AOI21X1  g15722(.A0(new_n18134_), .A1(new_n12048_), .B0(new_n18112_), .Y(new_n18159_));
  OAI21X1  g15723(.A0(new_n18159_), .A1(new_n18158_), .B0(new_n18157_), .Y(new_n18160_));
  NOR2X1   g15724(.A(new_n18137_), .B(pi0608), .Y(new_n18161_));
  NOR3X1   g15725(.A(new_n18158_), .B(new_n18112_), .C(new_n12364_), .Y(new_n18162_));
  NOR3X1   g15726(.A(new_n18162_), .B(new_n18138_), .C(new_n12368_), .Y(new_n18163_));
  AOI21X1  g15727(.A0(new_n18161_), .A1(new_n18160_), .B0(new_n18163_), .Y(new_n18164_));
  OR2X1    g15728(.A(new_n18159_), .B(pi0778), .Y(new_n18165_));
  OAI21X1  g15729(.A0(new_n18164_), .A1(new_n11769_), .B0(new_n18165_), .Y(new_n18166_));
  INVX1    g15730(.A(new_n18166_), .Y(new_n18167_));
  AND2X1   g15731(.A(new_n18166_), .B(new_n12462_), .Y(new_n18168_));
  OAI21X1  g15732(.A0(new_n18140_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n18169_));
  OR2X1    g15733(.A(new_n18169_), .B(new_n18168_), .Y(new_n18170_));
  AND3X1   g15734(.A(new_n18170_), .B(new_n18115_), .C(new_n12468_), .Y(new_n18171_));
  OAI21X1  g15735(.A0(new_n18140_), .A1(pi0609), .B0(pi1155), .Y(new_n18172_));
  AOI21X1  g15736(.A0(new_n18166_), .A1(pi0609), .B0(new_n18172_), .Y(new_n18173_));
  NOR3X1   g15737(.A(new_n18173_), .B(new_n18116_), .C(new_n12468_), .Y(new_n18174_));
  NOR2X1   g15738(.A(new_n18174_), .B(new_n18171_), .Y(new_n18175_));
  MX2X1    g15739(.A(new_n18175_), .B(new_n18167_), .S0(new_n11768_), .Y(new_n18176_));
  AOI21X1  g15740(.A0(new_n18139_), .A1(new_n18133_), .B0(new_n12630_), .Y(new_n18177_));
  AOI21X1  g15741(.A0(new_n18177_), .A1(pi0618), .B0(pi1154), .Y(new_n18178_));
  OAI21X1  g15742(.A0(new_n18176_), .A1(pi0618), .B0(new_n18178_), .Y(new_n18179_));
  NOR2X1   g15743(.A(new_n18120_), .B(pi0627), .Y(new_n18180_));
  AOI21X1  g15744(.A0(new_n18177_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18181_));
  OAI21X1  g15745(.A0(new_n18176_), .A1(new_n12486_), .B0(new_n18181_), .Y(new_n18182_));
  NOR2X1   g15746(.A(new_n18121_), .B(new_n12494_), .Y(new_n18183_));
  AOI22X1  g15747(.A0(new_n18183_), .A1(new_n18182_), .B0(new_n18180_), .B1(new_n18179_), .Y(new_n18184_));
  MX2X1    g15748(.A(new_n18184_), .B(new_n18176_), .S0(new_n11767_), .Y(new_n18185_));
  OR4X1    g15749(.A(new_n18140_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n18186_));
  AND2X1   g15750(.A(new_n18186_), .B(new_n12510_), .Y(new_n18187_));
  OAI21X1  g15751(.A0(new_n18185_), .A1(pi0619), .B0(new_n18187_), .Y(new_n18188_));
  NOR2X1   g15752(.A(new_n18125_), .B(pi0648), .Y(new_n18189_));
  AND2X1   g15753(.A(new_n18189_), .B(new_n18188_), .Y(new_n18190_));
  NOR4X1   g15754(.A(new_n18140_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n18191_));
  NOR2X1   g15755(.A(new_n18191_), .B(new_n12510_), .Y(new_n18192_));
  OAI21X1  g15756(.A0(new_n18185_), .A1(new_n12509_), .B0(new_n18192_), .Y(new_n18193_));
  NOR2X1   g15757(.A(new_n18126_), .B(new_n12517_), .Y(new_n18194_));
  AND2X1   g15758(.A(new_n18194_), .B(new_n18193_), .Y(new_n18195_));
  OR3X1    g15759(.A(new_n18195_), .B(new_n18190_), .C(new_n11766_), .Y(new_n18196_));
  AOI21X1  g15760(.A0(new_n18185_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n18197_));
  AOI21X1  g15761(.A0(new_n18197_), .A1(new_n18196_), .B0(new_n18156_), .Y(new_n18198_));
  OR2X1    g15762(.A(new_n18198_), .B(new_n14125_), .Y(new_n18199_));
  INVX1    g15763(.A(new_n18130_), .Y(new_n18200_));
  AND2X1   g15764(.A(new_n18141_), .B(new_n12718_), .Y(new_n18201_));
  AOI22X1  g15765(.A0(new_n18201_), .A1(new_n14426_), .B0(new_n18200_), .B1(new_n12735_), .Y(new_n18202_));
  AOI22X1  g15766(.A0(new_n18201_), .A1(new_n14428_), .B0(new_n18200_), .B1(new_n12733_), .Y(new_n18203_));
  MX2X1    g15767(.A(new_n18203_), .B(new_n18202_), .S0(new_n12561_), .Y(new_n18204_));
  OAI21X1  g15768(.A0(new_n18204_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n18205_));
  INVX1    g15769(.A(new_n18205_), .Y(new_n18206_));
  AOI21X1  g15770(.A0(new_n18206_), .A1(new_n18199_), .B0(new_n18149_), .Y(new_n18207_));
  OAI21X1  g15771(.A0(new_n18146_), .A1(new_n12578_), .B0(new_n18145_), .Y(new_n18208_));
  MX2X1    g15772(.A(new_n18208_), .B(new_n18143_), .S0(new_n11763_), .Y(new_n18209_));
  OAI21X1  g15773(.A0(new_n18209_), .A1(pi0644), .B0(pi0715), .Y(new_n18210_));
  AOI21X1  g15774(.A0(new_n18207_), .A1(pi0644), .B0(new_n18210_), .Y(new_n18211_));
  OR3X1    g15775(.A(new_n18110_), .B(new_n12603_), .C(new_n11763_), .Y(new_n18212_));
  OAI21X1  g15776(.A0(new_n18131_), .A1(new_n12604_), .B0(new_n18212_), .Y(new_n18213_));
  OAI21X1  g15777(.A0(new_n18110_), .A1(pi0644), .B0(new_n12608_), .Y(new_n18214_));
  AOI21X1  g15778(.A0(new_n18213_), .A1(pi0644), .B0(new_n18214_), .Y(new_n18215_));
  OR2X1    g15779(.A(new_n18215_), .B(new_n11762_), .Y(new_n18216_));
  OAI21X1  g15780(.A0(new_n18209_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n18217_));
  AOI21X1  g15781(.A0(new_n18207_), .A1(new_n12612_), .B0(new_n18217_), .Y(new_n18218_));
  OAI21X1  g15782(.A0(new_n18110_), .A1(new_n12612_), .B0(pi0715), .Y(new_n18219_));
  AOI21X1  g15783(.A0(new_n18213_), .A1(new_n12612_), .B0(new_n18219_), .Y(new_n18220_));
  OR2X1    g15784(.A(new_n18220_), .B(pi1160), .Y(new_n18221_));
  OAI22X1  g15785(.A0(new_n18221_), .A1(new_n18218_), .B0(new_n18216_), .B1(new_n18211_), .Y(new_n18222_));
  NAND2X1  g15786(.A(new_n18222_), .B(pi0790), .Y(new_n18223_));
  AOI21X1  g15787(.A0(new_n18207_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n18224_));
  AOI21X1  g15788(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0182), .Y(new_n18225_));
  INVX1    g15789(.A(new_n18225_), .Y(new_n18226_));
  AOI21X1  g15790(.A0(new_n3103_), .A1(new_n15095_), .B0(new_n18226_), .Y(new_n18227_));
  OAI21X1  g15791(.A0(new_n12826_), .A1(new_n5205_), .B0(new_n2979_), .Y(new_n18228_));
  AOI22X1  g15792(.A0(new_n18228_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n5205_), .Y(new_n18229_));
  AOI21X1  g15793(.A0(new_n12771_), .A1(new_n5205_), .B0(new_n12441_), .Y(new_n18230_));
  NOR3X1   g15794(.A(new_n18230_), .B(new_n18229_), .C(pi0734), .Y(new_n18231_));
  NOR2X1   g15795(.A(new_n18231_), .B(new_n18227_), .Y(new_n18232_));
  INVX1    g15796(.A(new_n18232_), .Y(new_n18233_));
  AOI21X1  g15797(.A0(new_n18225_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n18234_));
  OAI21X1  g15798(.A0(new_n18232_), .A1(new_n12363_), .B0(new_n18234_), .Y(new_n18235_));
  AOI21X1  g15799(.A0(new_n18225_), .A1(pi0625), .B0(pi1153), .Y(new_n18236_));
  OAI21X1  g15800(.A0(new_n18232_), .A1(pi0625), .B0(new_n18236_), .Y(new_n18237_));
  AND2X1   g15801(.A(new_n18237_), .B(new_n18235_), .Y(new_n18238_));
  MX2X1    g15802(.A(new_n18238_), .B(new_n18233_), .S0(new_n11769_), .Y(new_n18239_));
  MX2X1    g15803(.A(new_n18239_), .B(new_n18225_), .S0(new_n12490_), .Y(new_n18240_));
  INVX1    g15804(.A(new_n18240_), .Y(new_n18241_));
  MX2X1    g15805(.A(new_n18241_), .B(new_n18226_), .S0(new_n12513_), .Y(new_n18242_));
  INVX1    g15806(.A(new_n18242_), .Y(new_n18243_));
  MX2X1    g15807(.A(new_n18243_), .B(new_n18225_), .S0(new_n12531_), .Y(new_n18244_));
  MX2X1    g15808(.A(new_n18244_), .B(new_n18225_), .S0(new_n12563_), .Y(new_n18245_));
  INVX1    g15809(.A(new_n18245_), .Y(new_n18246_));
  AOI21X1  g15810(.A0(new_n18225_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n18247_));
  OAI21X1  g15811(.A0(new_n18246_), .A1(new_n12554_), .B0(new_n18247_), .Y(new_n18248_));
  AOI21X1  g15812(.A0(new_n18225_), .A1(pi0628), .B0(pi1156), .Y(new_n18249_));
  OAI21X1  g15813(.A0(new_n18246_), .A1(pi0628), .B0(new_n18249_), .Y(new_n18250_));
  AOI21X1  g15814(.A0(new_n18250_), .A1(new_n18248_), .B0(new_n11764_), .Y(new_n18251_));
  AOI21X1  g15815(.A0(new_n18246_), .A1(new_n11764_), .B0(new_n18251_), .Y(new_n18252_));
  MX2X1    g15816(.A(new_n18252_), .B(new_n18225_), .S0(pi0647), .Y(new_n18253_));
  MX2X1    g15817(.A(new_n18252_), .B(new_n18225_), .S0(new_n12577_), .Y(new_n18254_));
  MX2X1    g15818(.A(new_n18254_), .B(new_n18253_), .S0(new_n12578_), .Y(new_n18255_));
  MX2X1    g15819(.A(new_n18255_), .B(new_n18252_), .S0(new_n11763_), .Y(new_n18256_));
  AOI21X1  g15820(.A0(new_n18256_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n18257_));
  OAI22X1  g15821(.A0(new_n14197_), .A1(pi0756), .B0(new_n12077_), .B1(pi0182), .Y(new_n18258_));
  AOI21X1  g15822(.A0(new_n16615_), .A1(pi0182), .B0(pi0756), .Y(new_n18259_));
  OAI21X1  g15823(.A0(new_n12776_), .A1(pi0182), .B0(new_n18259_), .Y(new_n18260_));
  OR3X1    g15824(.A(new_n12445_), .B(new_n15068_), .C(pi0182), .Y(new_n18261_));
  AOI21X1  g15825(.A0(new_n18261_), .A1(new_n18260_), .B0(pi0038), .Y(new_n18262_));
  AOI21X1  g15826(.A0(new_n18258_), .A1(pi0038), .B0(new_n18262_), .Y(new_n18263_));
  MX2X1    g15827(.A(new_n18263_), .B(pi0182), .S0(new_n11770_), .Y(new_n18264_));
  AND2X1   g15828(.A(new_n18264_), .B(new_n12474_), .Y(new_n18265_));
  AOI21X1  g15829(.A0(new_n18226_), .A1(new_n12473_), .B0(new_n18265_), .Y(new_n18266_));
  AOI22X1  g15830(.A0(new_n18265_), .A1(pi0609), .B0(new_n18226_), .B1(new_n12472_), .Y(new_n18267_));
  AOI22X1  g15831(.A0(new_n18265_), .A1(new_n12462_), .B0(new_n18226_), .B1(new_n12481_), .Y(new_n18268_));
  MX2X1    g15832(.A(new_n18268_), .B(new_n18267_), .S0(pi1155), .Y(new_n18269_));
  MX2X1    g15833(.A(new_n18269_), .B(new_n18266_), .S0(new_n11768_), .Y(new_n18270_));
  OAI21X1  g15834(.A0(new_n18226_), .A1(pi0618), .B0(pi1154), .Y(new_n18271_));
  AOI21X1  g15835(.A0(new_n18270_), .A1(pi0618), .B0(new_n18271_), .Y(new_n18272_));
  OAI21X1  g15836(.A0(new_n18226_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18273_));
  AOI21X1  g15837(.A0(new_n18270_), .A1(new_n12486_), .B0(new_n18273_), .Y(new_n18274_));
  NOR2X1   g15838(.A(new_n18274_), .B(new_n18272_), .Y(new_n18275_));
  MX2X1    g15839(.A(new_n18275_), .B(new_n18270_), .S0(new_n11767_), .Y(new_n18276_));
  OAI21X1  g15840(.A0(new_n18226_), .A1(pi0619), .B0(pi1159), .Y(new_n18277_));
  AOI21X1  g15841(.A0(new_n18276_), .A1(pi0619), .B0(new_n18277_), .Y(new_n18278_));
  OAI21X1  g15842(.A0(new_n18226_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n18279_));
  AOI21X1  g15843(.A0(new_n18276_), .A1(new_n12509_), .B0(new_n18279_), .Y(new_n18280_));
  NOR2X1   g15844(.A(new_n18280_), .B(new_n18278_), .Y(new_n18281_));
  MX2X1    g15845(.A(new_n18281_), .B(new_n18276_), .S0(new_n11766_), .Y(new_n18282_));
  AND2X1   g15846(.A(new_n18225_), .B(new_n12708_), .Y(new_n18283_));
  AOI21X1  g15847(.A0(new_n18282_), .A1(new_n16140_), .B0(new_n18283_), .Y(new_n18284_));
  NAND2X1  g15848(.A(new_n18225_), .B(new_n12580_), .Y(new_n18285_));
  OAI21X1  g15849(.A0(new_n18284_), .A1(new_n12580_), .B0(new_n18285_), .Y(new_n18286_));
  MX2X1    g15850(.A(new_n18286_), .B(new_n18225_), .S0(new_n12604_), .Y(new_n18287_));
  OAI21X1  g15851(.A0(new_n18226_), .A1(pi0644), .B0(new_n12608_), .Y(new_n18288_));
  AOI21X1  g15852(.A0(new_n18287_), .A1(pi0644), .B0(new_n18288_), .Y(new_n18289_));
  OR2X1    g15853(.A(new_n18289_), .B(new_n11762_), .Y(new_n18290_));
  AOI21X1  g15854(.A0(new_n18256_), .A1(pi0644), .B0(pi0715), .Y(new_n18291_));
  OAI21X1  g15855(.A0(new_n18226_), .A1(new_n12612_), .B0(pi0715), .Y(new_n18292_));
  AOI21X1  g15856(.A0(new_n18287_), .A1(new_n12612_), .B0(new_n18292_), .Y(new_n18293_));
  OR2X1    g15857(.A(new_n18293_), .B(pi1160), .Y(new_n18294_));
  OAI22X1  g15858(.A0(new_n18294_), .A1(new_n18291_), .B0(new_n18290_), .B1(new_n18257_), .Y(new_n18295_));
  OR3X1    g15859(.A(new_n18293_), .B(pi1160), .C(pi0644), .Y(new_n18296_));
  OR3X1    g15860(.A(new_n18289_), .B(new_n11762_), .C(new_n12612_), .Y(new_n18297_));
  NAND3X1  g15861(.A(new_n18297_), .B(new_n18296_), .C(pi0790), .Y(new_n18298_));
  NAND2X1  g15862(.A(new_n18284_), .B(new_n14249_), .Y(new_n18299_));
  MX2X1    g15863(.A(new_n18250_), .B(new_n18248_), .S0(new_n12561_), .Y(new_n18300_));
  AND2X1   g15864(.A(new_n18300_), .B(new_n18299_), .Y(new_n18301_));
  OR2X1    g15865(.A(new_n18301_), .B(new_n11764_), .Y(new_n18302_));
  OR2X1    g15866(.A(new_n18263_), .B(new_n15095_), .Y(new_n18303_));
  OAI21X1  g15867(.A0(new_n12213_), .A1(new_n5205_), .B0(pi0756), .Y(new_n18304_));
  AOI21X1  g15868(.A0(new_n12155_), .A1(new_n5205_), .B0(new_n18304_), .Y(new_n18305_));
  AOI21X1  g15869(.A0(new_n12788_), .A1(new_n5205_), .B0(pi0756), .Y(new_n18306_));
  OAI21X1  g15870(.A0(new_n12787_), .A1(new_n5205_), .B0(new_n18306_), .Y(new_n18307_));
  NAND2X1  g15871(.A(new_n18307_), .B(pi0039), .Y(new_n18308_));
  AND2X1   g15872(.A(new_n12332_), .B(pi0182), .Y(new_n18309_));
  OAI21X1  g15873(.A0(new_n12315_), .A1(pi0182), .B0(pi0756), .Y(new_n18310_));
  NOR4X1   g15874(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0182), .Y(new_n18311_));
  OAI21X1  g15875(.A0(new_n12800_), .A1(new_n5205_), .B0(new_n15068_), .Y(new_n18312_));
  OAI22X1  g15876(.A0(new_n18312_), .A1(new_n18311_), .B0(new_n18310_), .B1(new_n18309_), .Y(new_n18313_));
  AOI21X1  g15877(.A0(new_n18313_), .A1(new_n2939_), .B0(pi0038), .Y(new_n18314_));
  OAI21X1  g15878(.A0(new_n18308_), .A1(new_n18305_), .B0(new_n18314_), .Y(new_n18315_));
  OAI21X1  g15879(.A0(new_n12276_), .A1(pi0756), .B0(new_n13540_), .Y(new_n18316_));
  NAND2X1  g15880(.A(new_n18316_), .B(new_n5205_), .Y(new_n18317_));
  AOI21X1  g15881(.A0(new_n12056_), .A1(new_n15068_), .B0(new_n13443_), .Y(new_n18318_));
  NOR2X1   g15882(.A(new_n18318_), .B(new_n5205_), .Y(new_n18319_));
  AOI21X1  g15883(.A0(new_n18319_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n18320_));
  AOI21X1  g15884(.A0(new_n18320_), .A1(new_n18317_), .B0(pi0734), .Y(new_n18321_));
  AOI21X1  g15885(.A0(new_n18321_), .A1(new_n18315_), .B0(new_n11770_), .Y(new_n18322_));
  AOI22X1  g15886(.A0(new_n18322_), .A1(new_n18303_), .B0(new_n11770_), .B1(pi0182), .Y(new_n18323_));
  OAI21X1  g15887(.A0(new_n18264_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n18324_));
  AOI21X1  g15888(.A0(new_n18323_), .A1(new_n12363_), .B0(new_n18324_), .Y(new_n18325_));
  NAND2X1  g15889(.A(new_n18235_), .B(new_n12368_), .Y(new_n18326_));
  OAI21X1  g15890(.A0(new_n18264_), .A1(pi0625), .B0(pi1153), .Y(new_n18327_));
  AOI21X1  g15891(.A0(new_n18323_), .A1(pi0625), .B0(new_n18327_), .Y(new_n18328_));
  NAND2X1  g15892(.A(new_n18237_), .B(pi0608), .Y(new_n18329_));
  OAI22X1  g15893(.A0(new_n18329_), .A1(new_n18328_), .B0(new_n18326_), .B1(new_n18325_), .Y(new_n18330_));
  MX2X1    g15894(.A(new_n18330_), .B(new_n18323_), .S0(new_n11769_), .Y(new_n18331_));
  INVX1    g15895(.A(new_n18239_), .Y(new_n18332_));
  OAI21X1  g15896(.A0(new_n18332_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n18333_));
  AOI21X1  g15897(.A0(new_n18331_), .A1(new_n12462_), .B0(new_n18333_), .Y(new_n18334_));
  OAI21X1  g15898(.A0(new_n18267_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n18335_));
  OAI21X1  g15899(.A0(new_n18332_), .A1(pi0609), .B0(pi1155), .Y(new_n18336_));
  AOI21X1  g15900(.A0(new_n18331_), .A1(pi0609), .B0(new_n18336_), .Y(new_n18337_));
  OAI21X1  g15901(.A0(new_n18268_), .A1(pi1155), .B0(pi0660), .Y(new_n18338_));
  OAI22X1  g15902(.A0(new_n18338_), .A1(new_n18337_), .B0(new_n18335_), .B1(new_n18334_), .Y(new_n18339_));
  MX2X1    g15903(.A(new_n18339_), .B(new_n18331_), .S0(new_n11768_), .Y(new_n18340_));
  OAI21X1  g15904(.A0(new_n18241_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18341_));
  AOI21X1  g15905(.A0(new_n18340_), .A1(new_n12486_), .B0(new_n18341_), .Y(new_n18342_));
  OR2X1    g15906(.A(new_n18272_), .B(pi0627), .Y(new_n18343_));
  OAI21X1  g15907(.A0(new_n18241_), .A1(pi0618), .B0(pi1154), .Y(new_n18344_));
  AOI21X1  g15908(.A0(new_n18340_), .A1(pi0618), .B0(new_n18344_), .Y(new_n18345_));
  OR2X1    g15909(.A(new_n18274_), .B(new_n12494_), .Y(new_n18346_));
  OAI22X1  g15910(.A0(new_n18346_), .A1(new_n18345_), .B0(new_n18343_), .B1(new_n18342_), .Y(new_n18347_));
  MX2X1    g15911(.A(new_n18347_), .B(new_n18340_), .S0(new_n11767_), .Y(new_n18348_));
  NAND2X1  g15912(.A(new_n18348_), .B(new_n12509_), .Y(new_n18349_));
  AOI21X1  g15913(.A0(new_n18243_), .A1(pi0619), .B0(pi1159), .Y(new_n18350_));
  OR2X1    g15914(.A(new_n18278_), .B(pi0648), .Y(new_n18351_));
  AOI21X1  g15915(.A0(new_n18350_), .A1(new_n18349_), .B0(new_n18351_), .Y(new_n18352_));
  NAND2X1  g15916(.A(new_n18348_), .B(pi0619), .Y(new_n18353_));
  AOI21X1  g15917(.A0(new_n18243_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n18354_));
  OR2X1    g15918(.A(new_n18280_), .B(new_n12517_), .Y(new_n18355_));
  AOI21X1  g15919(.A0(new_n18354_), .A1(new_n18353_), .B0(new_n18355_), .Y(new_n18356_));
  NOR3X1   g15920(.A(new_n18356_), .B(new_n18352_), .C(new_n11766_), .Y(new_n18357_));
  OAI21X1  g15921(.A0(new_n18348_), .A1(pi0789), .B0(new_n12709_), .Y(new_n18358_));
  AOI21X1  g15922(.A0(new_n18226_), .A1(pi0626), .B0(new_n16218_), .Y(new_n18359_));
  OAI21X1  g15923(.A0(new_n18282_), .A1(pi0626), .B0(new_n18359_), .Y(new_n18360_));
  AOI21X1  g15924(.A0(new_n18226_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n18361_));
  OAI21X1  g15925(.A0(new_n18282_), .A1(new_n12542_), .B0(new_n18361_), .Y(new_n18362_));
  NAND2X1  g15926(.A(new_n18244_), .B(new_n12637_), .Y(new_n18363_));
  NAND3X1  g15927(.A(new_n18363_), .B(new_n18362_), .C(new_n18360_), .Y(new_n18364_));
  AOI21X1  g15928(.A0(new_n18364_), .A1(pi0788), .B0(new_n14125_), .Y(new_n18365_));
  OAI21X1  g15929(.A0(new_n18358_), .A1(new_n18357_), .B0(new_n18365_), .Y(new_n18366_));
  AOI21X1  g15930(.A0(new_n18366_), .A1(new_n18302_), .B0(new_n14121_), .Y(new_n18367_));
  OR2X1    g15931(.A(new_n18286_), .B(new_n14239_), .Y(new_n18368_));
  OR2X1    g15932(.A(new_n18253_), .B(new_n14244_), .Y(new_n18369_));
  OR2X1    g15933(.A(new_n18254_), .B(new_n14242_), .Y(new_n18370_));
  NAND3X1  g15934(.A(new_n18370_), .B(new_n18369_), .C(new_n18368_), .Y(new_n18371_));
  AOI21X1  g15935(.A0(new_n18371_), .A1(pi0787), .B0(new_n18367_), .Y(new_n18372_));
  AOI22X1  g15936(.A0(new_n18372_), .A1(new_n18298_), .B0(new_n18295_), .B1(pi0790), .Y(new_n18373_));
  OR2X1    g15937(.A(new_n18373_), .B(po1038), .Y(new_n18374_));
  AOI21X1  g15938(.A0(po1038), .A1(new_n5205_), .B0(pi0832), .Y(new_n18375_));
  AOI22X1  g15939(.A0(new_n18375_), .A1(new_n18374_), .B0(new_n18224_), .B1(new_n18223_), .Y(po0339));
  AOI21X1  g15940(.A0(pi1093), .A1(pi1092), .B0(pi0183), .Y(new_n18377_));
  INVX1    g15941(.A(new_n18377_), .Y(new_n18378_));
  AOI21X1  g15942(.A0(new_n12056_), .A1(new_n14640_), .B0(new_n18377_), .Y(new_n18379_));
  INVX1    g15943(.A(new_n18379_), .Y(new_n18380_));
  NAND2X1  g15944(.A(new_n18380_), .B(new_n15771_), .Y(new_n18381_));
  AND3X1   g15945(.A(new_n12480_), .B(new_n12056_), .C(new_n14640_), .Y(new_n18382_));
  OAI21X1  g15946(.A0(new_n18382_), .A1(new_n18381_), .B0(pi1155), .Y(new_n18383_));
  NOR3X1   g15947(.A(new_n18382_), .B(new_n18377_), .C(pi1155), .Y(new_n18384_));
  INVX1    g15948(.A(new_n18384_), .Y(new_n18385_));
  AOI21X1  g15949(.A0(new_n18385_), .A1(new_n18383_), .B0(new_n11768_), .Y(new_n18386_));
  AOI21X1  g15950(.A0(new_n18381_), .A1(new_n11768_), .B0(new_n18386_), .Y(new_n18387_));
  AOI21X1  g15951(.A0(new_n18387_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n18388_));
  AOI21X1  g15952(.A0(new_n18387_), .A1(new_n12655_), .B0(pi1154), .Y(new_n18389_));
  NOR2X1   g15953(.A(new_n18389_), .B(new_n18388_), .Y(new_n18390_));
  MX2X1    g15954(.A(new_n18390_), .B(new_n18387_), .S0(new_n11767_), .Y(new_n18391_));
  NOR2X1   g15955(.A(new_n18391_), .B(pi0789), .Y(new_n18392_));
  AOI21X1  g15956(.A0(new_n18391_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n18393_));
  AOI21X1  g15957(.A0(new_n18391_), .A1(new_n15790_), .B0(pi1159), .Y(new_n18394_));
  OR2X1    g15958(.A(new_n18394_), .B(new_n18393_), .Y(new_n18395_));
  AOI21X1  g15959(.A0(new_n18395_), .A1(pi0789), .B0(new_n18392_), .Y(new_n18396_));
  INVX1    g15960(.A(new_n18396_), .Y(new_n18397_));
  MX2X1    g15961(.A(new_n18397_), .B(new_n18378_), .S0(new_n12708_), .Y(new_n18398_));
  MX2X1    g15962(.A(new_n18398_), .B(new_n18378_), .S0(new_n12580_), .Y(new_n18399_));
  AOI21X1  g15963(.A0(new_n12439_), .A1(new_n14667_), .B0(new_n18377_), .Y(new_n18400_));
  OR2X1    g15964(.A(new_n18400_), .B(pi0778), .Y(new_n18401_));
  INVX1    g15965(.A(new_n18400_), .Y(new_n18402_));
  AND3X1   g15966(.A(new_n12439_), .B(new_n14667_), .C(new_n12363_), .Y(new_n18403_));
  INVX1    g15967(.A(new_n18403_), .Y(new_n18404_));
  AOI21X1  g15968(.A0(new_n18404_), .A1(new_n18402_), .B0(new_n12364_), .Y(new_n18405_));
  NOR3X1   g15969(.A(new_n18403_), .B(new_n18377_), .C(pi1153), .Y(new_n18406_));
  OR3X1    g15970(.A(new_n18406_), .B(new_n18405_), .C(new_n11769_), .Y(new_n18407_));
  AND2X1   g15971(.A(new_n18407_), .B(new_n18401_), .Y(new_n18408_));
  NOR4X1   g15972(.A(new_n18408_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n18409_));
  AND3X1   g15973(.A(new_n18409_), .B(new_n12739_), .C(new_n12718_), .Y(new_n18410_));
  INVX1    g15974(.A(new_n18410_), .Y(new_n18411_));
  AOI21X1  g15975(.A0(new_n18377_), .A1(pi0647), .B0(pi1157), .Y(new_n18412_));
  OAI21X1  g15976(.A0(new_n18411_), .A1(pi0647), .B0(new_n18412_), .Y(new_n18413_));
  MX2X1    g15977(.A(new_n18410_), .B(new_n18377_), .S0(new_n12577_), .Y(new_n18414_));
  OAI22X1  g15978(.A0(new_n18414_), .A1(new_n14242_), .B0(new_n18413_), .B1(new_n12592_), .Y(new_n18415_));
  AOI21X1  g15979(.A0(new_n18399_), .A1(new_n14326_), .B0(new_n18415_), .Y(new_n18416_));
  NOR2X1   g15980(.A(new_n18416_), .B(new_n11763_), .Y(new_n18417_));
  AOI21X1  g15981(.A0(new_n18378_), .A1(pi0626), .B0(new_n16218_), .Y(new_n18418_));
  OAI21X1  g15982(.A0(new_n18396_), .A1(pi0626), .B0(new_n18418_), .Y(new_n18419_));
  AOI21X1  g15983(.A0(new_n18378_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n18420_));
  OAI21X1  g15984(.A0(new_n18396_), .A1(new_n12542_), .B0(new_n18420_), .Y(new_n18421_));
  NAND2X1  g15985(.A(new_n18409_), .B(new_n12637_), .Y(new_n18422_));
  AND3X1   g15986(.A(new_n18422_), .B(new_n18421_), .C(new_n18419_), .Y(new_n18423_));
  NOR2X1   g15987(.A(new_n18423_), .B(new_n11765_), .Y(new_n18424_));
  NOR2X1   g15988(.A(new_n18377_), .B(pi1153), .Y(new_n18425_));
  NOR3X1   g15989(.A(new_n18400_), .B(new_n11991_), .C(new_n12363_), .Y(new_n18426_));
  AOI21X1  g15990(.A0(new_n18402_), .A1(new_n12048_), .B0(new_n18380_), .Y(new_n18427_));
  OAI21X1  g15991(.A0(new_n18427_), .A1(new_n18426_), .B0(new_n18425_), .Y(new_n18428_));
  NOR2X1   g15992(.A(new_n18405_), .B(pi0608), .Y(new_n18429_));
  NOR3X1   g15993(.A(new_n18426_), .B(new_n18380_), .C(new_n12364_), .Y(new_n18430_));
  NOR3X1   g15994(.A(new_n18430_), .B(new_n18406_), .C(new_n12368_), .Y(new_n18431_));
  AOI21X1  g15995(.A0(new_n18429_), .A1(new_n18428_), .B0(new_n18431_), .Y(new_n18432_));
  OR2X1    g15996(.A(new_n18427_), .B(pi0778), .Y(new_n18433_));
  OAI21X1  g15997(.A0(new_n18432_), .A1(new_n11769_), .B0(new_n18433_), .Y(new_n18434_));
  INVX1    g15998(.A(new_n18434_), .Y(new_n18435_));
  AND2X1   g15999(.A(new_n18434_), .B(new_n12462_), .Y(new_n18436_));
  OAI21X1  g16000(.A0(new_n18408_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n18437_));
  OR2X1    g16001(.A(new_n18437_), .B(new_n18436_), .Y(new_n18438_));
  AND3X1   g16002(.A(new_n18438_), .B(new_n18383_), .C(new_n12468_), .Y(new_n18439_));
  OAI21X1  g16003(.A0(new_n18408_), .A1(pi0609), .B0(pi1155), .Y(new_n18440_));
  AOI21X1  g16004(.A0(new_n18434_), .A1(pi0609), .B0(new_n18440_), .Y(new_n18441_));
  NOR3X1   g16005(.A(new_n18441_), .B(new_n18384_), .C(new_n12468_), .Y(new_n18442_));
  NOR2X1   g16006(.A(new_n18442_), .B(new_n18439_), .Y(new_n18443_));
  MX2X1    g16007(.A(new_n18443_), .B(new_n18435_), .S0(new_n11768_), .Y(new_n18444_));
  AOI21X1  g16008(.A0(new_n18407_), .A1(new_n18401_), .B0(new_n12630_), .Y(new_n18445_));
  AOI21X1  g16009(.A0(new_n18445_), .A1(pi0618), .B0(pi1154), .Y(new_n18446_));
  OAI21X1  g16010(.A0(new_n18444_), .A1(pi0618), .B0(new_n18446_), .Y(new_n18447_));
  NOR2X1   g16011(.A(new_n18388_), .B(pi0627), .Y(new_n18448_));
  AOI21X1  g16012(.A0(new_n18445_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18449_));
  OAI21X1  g16013(.A0(new_n18444_), .A1(new_n12486_), .B0(new_n18449_), .Y(new_n18450_));
  NOR2X1   g16014(.A(new_n18389_), .B(new_n12494_), .Y(new_n18451_));
  AOI22X1  g16015(.A0(new_n18451_), .A1(new_n18450_), .B0(new_n18448_), .B1(new_n18447_), .Y(new_n18452_));
  MX2X1    g16016(.A(new_n18452_), .B(new_n18444_), .S0(new_n11767_), .Y(new_n18453_));
  OR4X1    g16017(.A(new_n18408_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n18454_));
  AND2X1   g16018(.A(new_n18454_), .B(new_n12510_), .Y(new_n18455_));
  OAI21X1  g16019(.A0(new_n18453_), .A1(pi0619), .B0(new_n18455_), .Y(new_n18456_));
  NOR2X1   g16020(.A(new_n18393_), .B(pi0648), .Y(new_n18457_));
  AND2X1   g16021(.A(new_n18457_), .B(new_n18456_), .Y(new_n18458_));
  NOR4X1   g16022(.A(new_n18408_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n18459_));
  NOR2X1   g16023(.A(new_n18459_), .B(new_n12510_), .Y(new_n18460_));
  OAI21X1  g16024(.A0(new_n18453_), .A1(new_n12509_), .B0(new_n18460_), .Y(new_n18461_));
  NOR2X1   g16025(.A(new_n18394_), .B(new_n12517_), .Y(new_n18462_));
  AND2X1   g16026(.A(new_n18462_), .B(new_n18461_), .Y(new_n18463_));
  OR3X1    g16027(.A(new_n18463_), .B(new_n18458_), .C(new_n11766_), .Y(new_n18464_));
  AOI21X1  g16028(.A0(new_n18453_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n18465_));
  AOI21X1  g16029(.A0(new_n18465_), .A1(new_n18464_), .B0(new_n18424_), .Y(new_n18466_));
  OR2X1    g16030(.A(new_n18466_), .B(new_n14125_), .Y(new_n18467_));
  INVX1    g16031(.A(new_n18398_), .Y(new_n18468_));
  AND2X1   g16032(.A(new_n18409_), .B(new_n12718_), .Y(new_n18469_));
  AOI22X1  g16033(.A0(new_n18469_), .A1(new_n14426_), .B0(new_n18468_), .B1(new_n12735_), .Y(new_n18470_));
  AOI22X1  g16034(.A0(new_n18469_), .A1(new_n14428_), .B0(new_n18468_), .B1(new_n12733_), .Y(new_n18471_));
  MX2X1    g16035(.A(new_n18471_), .B(new_n18470_), .S0(new_n12561_), .Y(new_n18472_));
  OAI21X1  g16036(.A0(new_n18472_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n18473_));
  INVX1    g16037(.A(new_n18473_), .Y(new_n18474_));
  AOI21X1  g16038(.A0(new_n18474_), .A1(new_n18467_), .B0(new_n18417_), .Y(new_n18475_));
  OAI21X1  g16039(.A0(new_n18414_), .A1(new_n12578_), .B0(new_n18413_), .Y(new_n18476_));
  MX2X1    g16040(.A(new_n18476_), .B(new_n18411_), .S0(new_n11763_), .Y(new_n18477_));
  OAI21X1  g16041(.A0(new_n18477_), .A1(pi0644), .B0(pi0715), .Y(new_n18478_));
  AOI21X1  g16042(.A0(new_n18475_), .A1(pi0644), .B0(new_n18478_), .Y(new_n18479_));
  OR3X1    g16043(.A(new_n18378_), .B(new_n12603_), .C(new_n11763_), .Y(new_n18480_));
  OAI21X1  g16044(.A0(new_n18399_), .A1(new_n12604_), .B0(new_n18480_), .Y(new_n18481_));
  OAI21X1  g16045(.A0(new_n18378_), .A1(pi0644), .B0(new_n12608_), .Y(new_n18482_));
  AOI21X1  g16046(.A0(new_n18481_), .A1(pi0644), .B0(new_n18482_), .Y(new_n18483_));
  OR2X1    g16047(.A(new_n18483_), .B(new_n11762_), .Y(new_n18484_));
  OAI21X1  g16048(.A0(new_n18477_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n18485_));
  AOI21X1  g16049(.A0(new_n18475_), .A1(new_n12612_), .B0(new_n18485_), .Y(new_n18486_));
  OAI21X1  g16050(.A0(new_n18378_), .A1(new_n12612_), .B0(pi0715), .Y(new_n18487_));
  AOI21X1  g16051(.A0(new_n18481_), .A1(new_n12612_), .B0(new_n18487_), .Y(new_n18488_));
  OR2X1    g16052(.A(new_n18488_), .B(pi1160), .Y(new_n18489_));
  OAI22X1  g16053(.A0(new_n18489_), .A1(new_n18486_), .B0(new_n18484_), .B1(new_n18479_), .Y(new_n18490_));
  NAND2X1  g16054(.A(new_n18490_), .B(pi0790), .Y(new_n18491_));
  AOI21X1  g16055(.A0(new_n18475_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n18492_));
  AOI21X1  g16056(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0183), .Y(new_n18493_));
  INVX1    g16057(.A(new_n18493_), .Y(new_n18494_));
  AOI21X1  g16058(.A0(new_n3103_), .A1(new_n14667_), .B0(new_n18494_), .Y(new_n18495_));
  OAI21X1  g16059(.A0(new_n12826_), .A1(new_n6802_), .B0(new_n2979_), .Y(new_n18496_));
  AOI22X1  g16060(.A0(new_n18496_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n6802_), .Y(new_n18497_));
  AOI21X1  g16061(.A0(new_n12771_), .A1(new_n6802_), .B0(new_n12441_), .Y(new_n18498_));
  NOR3X1   g16062(.A(new_n18498_), .B(new_n18497_), .C(pi0725), .Y(new_n18499_));
  NOR2X1   g16063(.A(new_n18499_), .B(new_n18495_), .Y(new_n18500_));
  INVX1    g16064(.A(new_n18500_), .Y(new_n18501_));
  AOI21X1  g16065(.A0(new_n18493_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n18502_));
  OAI21X1  g16066(.A0(new_n18500_), .A1(new_n12363_), .B0(new_n18502_), .Y(new_n18503_));
  AOI21X1  g16067(.A0(new_n18493_), .A1(pi0625), .B0(pi1153), .Y(new_n18504_));
  OAI21X1  g16068(.A0(new_n18500_), .A1(pi0625), .B0(new_n18504_), .Y(new_n18505_));
  AND2X1   g16069(.A(new_n18505_), .B(new_n18503_), .Y(new_n18506_));
  MX2X1    g16070(.A(new_n18506_), .B(new_n18501_), .S0(new_n11769_), .Y(new_n18507_));
  MX2X1    g16071(.A(new_n18507_), .B(new_n18493_), .S0(new_n12490_), .Y(new_n18508_));
  INVX1    g16072(.A(new_n18508_), .Y(new_n18509_));
  MX2X1    g16073(.A(new_n18509_), .B(new_n18494_), .S0(new_n12513_), .Y(new_n18510_));
  INVX1    g16074(.A(new_n18510_), .Y(new_n18511_));
  MX2X1    g16075(.A(new_n18511_), .B(new_n18493_), .S0(new_n12531_), .Y(new_n18512_));
  MX2X1    g16076(.A(new_n18512_), .B(new_n18493_), .S0(new_n12563_), .Y(new_n18513_));
  INVX1    g16077(.A(new_n18513_), .Y(new_n18514_));
  AOI21X1  g16078(.A0(new_n18493_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n18515_));
  OAI21X1  g16079(.A0(new_n18514_), .A1(new_n12554_), .B0(new_n18515_), .Y(new_n18516_));
  AOI21X1  g16080(.A0(new_n18493_), .A1(pi0628), .B0(pi1156), .Y(new_n18517_));
  OAI21X1  g16081(.A0(new_n18514_), .A1(pi0628), .B0(new_n18517_), .Y(new_n18518_));
  AOI21X1  g16082(.A0(new_n18518_), .A1(new_n18516_), .B0(new_n11764_), .Y(new_n18519_));
  AOI21X1  g16083(.A0(new_n18514_), .A1(new_n11764_), .B0(new_n18519_), .Y(new_n18520_));
  MX2X1    g16084(.A(new_n18520_), .B(new_n18493_), .S0(pi0647), .Y(new_n18521_));
  MX2X1    g16085(.A(new_n18520_), .B(new_n18493_), .S0(new_n12577_), .Y(new_n18522_));
  MX2X1    g16086(.A(new_n18522_), .B(new_n18521_), .S0(new_n12578_), .Y(new_n18523_));
  MX2X1    g16087(.A(new_n18523_), .B(new_n18520_), .S0(new_n11763_), .Y(new_n18524_));
  AOI21X1  g16088(.A0(new_n18524_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n18525_));
  OAI22X1  g16089(.A0(new_n14197_), .A1(pi0755), .B0(new_n12077_), .B1(pi0183), .Y(new_n18526_));
  AOI21X1  g16090(.A0(new_n16615_), .A1(pi0183), .B0(pi0755), .Y(new_n18527_));
  OAI21X1  g16091(.A0(new_n12776_), .A1(pi0183), .B0(new_n18527_), .Y(new_n18528_));
  OR3X1    g16092(.A(new_n12445_), .B(new_n14640_), .C(pi0183), .Y(new_n18529_));
  AOI21X1  g16093(.A0(new_n18529_), .A1(new_n18528_), .B0(pi0038), .Y(new_n18530_));
  AOI21X1  g16094(.A0(new_n18526_), .A1(pi0038), .B0(new_n18530_), .Y(new_n18531_));
  MX2X1    g16095(.A(new_n18531_), .B(pi0183), .S0(new_n11770_), .Y(new_n18532_));
  AND2X1   g16096(.A(new_n18532_), .B(new_n12474_), .Y(new_n18533_));
  AOI21X1  g16097(.A0(new_n18494_), .A1(new_n12473_), .B0(new_n18533_), .Y(new_n18534_));
  AOI22X1  g16098(.A0(new_n18533_), .A1(pi0609), .B0(new_n18494_), .B1(new_n12472_), .Y(new_n18535_));
  AOI22X1  g16099(.A0(new_n18533_), .A1(new_n12462_), .B0(new_n18494_), .B1(new_n12481_), .Y(new_n18536_));
  MX2X1    g16100(.A(new_n18536_), .B(new_n18535_), .S0(pi1155), .Y(new_n18537_));
  MX2X1    g16101(.A(new_n18537_), .B(new_n18534_), .S0(new_n11768_), .Y(new_n18538_));
  OAI21X1  g16102(.A0(new_n18494_), .A1(pi0618), .B0(pi1154), .Y(new_n18539_));
  AOI21X1  g16103(.A0(new_n18538_), .A1(pi0618), .B0(new_n18539_), .Y(new_n18540_));
  OAI21X1  g16104(.A0(new_n18494_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18541_));
  AOI21X1  g16105(.A0(new_n18538_), .A1(new_n12486_), .B0(new_n18541_), .Y(new_n18542_));
  NOR2X1   g16106(.A(new_n18542_), .B(new_n18540_), .Y(new_n18543_));
  MX2X1    g16107(.A(new_n18543_), .B(new_n18538_), .S0(new_n11767_), .Y(new_n18544_));
  OAI21X1  g16108(.A0(new_n18494_), .A1(pi0619), .B0(pi1159), .Y(new_n18545_));
  AOI21X1  g16109(.A0(new_n18544_), .A1(pi0619), .B0(new_n18545_), .Y(new_n18546_));
  OAI21X1  g16110(.A0(new_n18494_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n18547_));
  AOI21X1  g16111(.A0(new_n18544_), .A1(new_n12509_), .B0(new_n18547_), .Y(new_n18548_));
  NOR2X1   g16112(.A(new_n18548_), .B(new_n18546_), .Y(new_n18549_));
  MX2X1    g16113(.A(new_n18549_), .B(new_n18544_), .S0(new_n11766_), .Y(new_n18550_));
  AND2X1   g16114(.A(new_n18493_), .B(new_n12708_), .Y(new_n18551_));
  AOI21X1  g16115(.A0(new_n18550_), .A1(new_n16140_), .B0(new_n18551_), .Y(new_n18552_));
  NAND2X1  g16116(.A(new_n18493_), .B(new_n12580_), .Y(new_n18553_));
  OAI21X1  g16117(.A0(new_n18552_), .A1(new_n12580_), .B0(new_n18553_), .Y(new_n18554_));
  MX2X1    g16118(.A(new_n18554_), .B(new_n18493_), .S0(new_n12604_), .Y(new_n18555_));
  OAI21X1  g16119(.A0(new_n18494_), .A1(pi0644), .B0(new_n12608_), .Y(new_n18556_));
  AOI21X1  g16120(.A0(new_n18555_), .A1(pi0644), .B0(new_n18556_), .Y(new_n18557_));
  OR2X1    g16121(.A(new_n18557_), .B(new_n11762_), .Y(new_n18558_));
  AOI21X1  g16122(.A0(new_n18524_), .A1(pi0644), .B0(pi0715), .Y(new_n18559_));
  OAI21X1  g16123(.A0(new_n18494_), .A1(new_n12612_), .B0(pi0715), .Y(new_n18560_));
  AOI21X1  g16124(.A0(new_n18555_), .A1(new_n12612_), .B0(new_n18560_), .Y(new_n18561_));
  OR2X1    g16125(.A(new_n18561_), .B(pi1160), .Y(new_n18562_));
  OAI22X1  g16126(.A0(new_n18562_), .A1(new_n18559_), .B0(new_n18558_), .B1(new_n18525_), .Y(new_n18563_));
  OR3X1    g16127(.A(new_n18561_), .B(pi1160), .C(pi0644), .Y(new_n18564_));
  OR3X1    g16128(.A(new_n18557_), .B(new_n11762_), .C(new_n12612_), .Y(new_n18565_));
  NAND3X1  g16129(.A(new_n18565_), .B(new_n18564_), .C(pi0790), .Y(new_n18566_));
  NAND2X1  g16130(.A(new_n18552_), .B(new_n14249_), .Y(new_n18567_));
  MX2X1    g16131(.A(new_n18518_), .B(new_n18516_), .S0(new_n12561_), .Y(new_n18568_));
  AND2X1   g16132(.A(new_n18568_), .B(new_n18567_), .Y(new_n18569_));
  OR2X1    g16133(.A(new_n18569_), .B(new_n11764_), .Y(new_n18570_));
  OR2X1    g16134(.A(new_n18531_), .B(new_n14667_), .Y(new_n18571_));
  OAI21X1  g16135(.A0(new_n12213_), .A1(new_n6802_), .B0(pi0755), .Y(new_n18572_));
  AOI21X1  g16136(.A0(new_n12155_), .A1(new_n6802_), .B0(new_n18572_), .Y(new_n18573_));
  AOI21X1  g16137(.A0(new_n12788_), .A1(new_n6802_), .B0(pi0755), .Y(new_n18574_));
  OAI21X1  g16138(.A0(new_n12787_), .A1(new_n6802_), .B0(new_n18574_), .Y(new_n18575_));
  NAND2X1  g16139(.A(new_n18575_), .B(pi0039), .Y(new_n18576_));
  AND2X1   g16140(.A(new_n12332_), .B(pi0183), .Y(new_n18577_));
  OAI21X1  g16141(.A0(new_n12315_), .A1(pi0183), .B0(pi0755), .Y(new_n18578_));
  NOR4X1   g16142(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0183), .Y(new_n18579_));
  OAI21X1  g16143(.A0(new_n12800_), .A1(new_n6802_), .B0(new_n14640_), .Y(new_n18580_));
  OAI22X1  g16144(.A0(new_n18580_), .A1(new_n18579_), .B0(new_n18578_), .B1(new_n18577_), .Y(new_n18581_));
  AOI21X1  g16145(.A0(new_n18581_), .A1(new_n2939_), .B0(pi0038), .Y(new_n18582_));
  OAI21X1  g16146(.A0(new_n18576_), .A1(new_n18573_), .B0(new_n18582_), .Y(new_n18583_));
  OAI21X1  g16147(.A0(new_n12276_), .A1(pi0755), .B0(new_n13540_), .Y(new_n18584_));
  NAND2X1  g16148(.A(new_n18584_), .B(new_n6802_), .Y(new_n18585_));
  AOI21X1  g16149(.A0(new_n12056_), .A1(new_n14640_), .B0(new_n13443_), .Y(new_n18586_));
  NOR2X1   g16150(.A(new_n18586_), .B(new_n6802_), .Y(new_n18587_));
  AOI21X1  g16151(.A0(new_n18587_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n18588_));
  AOI21X1  g16152(.A0(new_n18588_), .A1(new_n18585_), .B0(pi0725), .Y(new_n18589_));
  AOI21X1  g16153(.A0(new_n18589_), .A1(new_n18583_), .B0(new_n11770_), .Y(new_n18590_));
  AOI22X1  g16154(.A0(new_n18590_), .A1(new_n18571_), .B0(new_n11770_), .B1(pi0183), .Y(new_n18591_));
  OAI21X1  g16155(.A0(new_n18532_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n18592_));
  AOI21X1  g16156(.A0(new_n18591_), .A1(new_n12363_), .B0(new_n18592_), .Y(new_n18593_));
  NAND2X1  g16157(.A(new_n18503_), .B(new_n12368_), .Y(new_n18594_));
  OAI21X1  g16158(.A0(new_n18532_), .A1(pi0625), .B0(pi1153), .Y(new_n18595_));
  AOI21X1  g16159(.A0(new_n18591_), .A1(pi0625), .B0(new_n18595_), .Y(new_n18596_));
  NAND2X1  g16160(.A(new_n18505_), .B(pi0608), .Y(new_n18597_));
  OAI22X1  g16161(.A0(new_n18597_), .A1(new_n18596_), .B0(new_n18594_), .B1(new_n18593_), .Y(new_n18598_));
  MX2X1    g16162(.A(new_n18598_), .B(new_n18591_), .S0(new_n11769_), .Y(new_n18599_));
  INVX1    g16163(.A(new_n18507_), .Y(new_n18600_));
  OAI21X1  g16164(.A0(new_n18600_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n18601_));
  AOI21X1  g16165(.A0(new_n18599_), .A1(new_n12462_), .B0(new_n18601_), .Y(new_n18602_));
  OAI21X1  g16166(.A0(new_n18535_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n18603_));
  OAI21X1  g16167(.A0(new_n18600_), .A1(pi0609), .B0(pi1155), .Y(new_n18604_));
  AOI21X1  g16168(.A0(new_n18599_), .A1(pi0609), .B0(new_n18604_), .Y(new_n18605_));
  OAI21X1  g16169(.A0(new_n18536_), .A1(pi1155), .B0(pi0660), .Y(new_n18606_));
  OAI22X1  g16170(.A0(new_n18606_), .A1(new_n18605_), .B0(new_n18603_), .B1(new_n18602_), .Y(new_n18607_));
  MX2X1    g16171(.A(new_n18607_), .B(new_n18599_), .S0(new_n11768_), .Y(new_n18608_));
  OAI21X1  g16172(.A0(new_n18509_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18609_));
  AOI21X1  g16173(.A0(new_n18608_), .A1(new_n12486_), .B0(new_n18609_), .Y(new_n18610_));
  OR2X1    g16174(.A(new_n18540_), .B(pi0627), .Y(new_n18611_));
  OAI21X1  g16175(.A0(new_n18509_), .A1(pi0618), .B0(pi1154), .Y(new_n18612_));
  AOI21X1  g16176(.A0(new_n18608_), .A1(pi0618), .B0(new_n18612_), .Y(new_n18613_));
  OR2X1    g16177(.A(new_n18542_), .B(new_n12494_), .Y(new_n18614_));
  OAI22X1  g16178(.A0(new_n18614_), .A1(new_n18613_), .B0(new_n18611_), .B1(new_n18610_), .Y(new_n18615_));
  MX2X1    g16179(.A(new_n18615_), .B(new_n18608_), .S0(new_n11767_), .Y(new_n18616_));
  NAND2X1  g16180(.A(new_n18616_), .B(new_n12509_), .Y(new_n18617_));
  AOI21X1  g16181(.A0(new_n18511_), .A1(pi0619), .B0(pi1159), .Y(new_n18618_));
  OR2X1    g16182(.A(new_n18546_), .B(pi0648), .Y(new_n18619_));
  AOI21X1  g16183(.A0(new_n18618_), .A1(new_n18617_), .B0(new_n18619_), .Y(new_n18620_));
  NAND2X1  g16184(.A(new_n18616_), .B(pi0619), .Y(new_n18621_));
  AOI21X1  g16185(.A0(new_n18511_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n18622_));
  OR2X1    g16186(.A(new_n18548_), .B(new_n12517_), .Y(new_n18623_));
  AOI21X1  g16187(.A0(new_n18622_), .A1(new_n18621_), .B0(new_n18623_), .Y(new_n18624_));
  NOR3X1   g16188(.A(new_n18624_), .B(new_n18620_), .C(new_n11766_), .Y(new_n18625_));
  OAI21X1  g16189(.A0(new_n18616_), .A1(pi0789), .B0(new_n12709_), .Y(new_n18626_));
  AOI21X1  g16190(.A0(new_n18494_), .A1(pi0626), .B0(new_n16218_), .Y(new_n18627_));
  OAI21X1  g16191(.A0(new_n18550_), .A1(pi0626), .B0(new_n18627_), .Y(new_n18628_));
  AOI21X1  g16192(.A0(new_n18494_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n18629_));
  OAI21X1  g16193(.A0(new_n18550_), .A1(new_n12542_), .B0(new_n18629_), .Y(new_n18630_));
  NAND2X1  g16194(.A(new_n18512_), .B(new_n12637_), .Y(new_n18631_));
  NAND3X1  g16195(.A(new_n18631_), .B(new_n18630_), .C(new_n18628_), .Y(new_n18632_));
  AOI21X1  g16196(.A0(new_n18632_), .A1(pi0788), .B0(new_n14125_), .Y(new_n18633_));
  OAI21X1  g16197(.A0(new_n18626_), .A1(new_n18625_), .B0(new_n18633_), .Y(new_n18634_));
  AOI21X1  g16198(.A0(new_n18634_), .A1(new_n18570_), .B0(new_n14121_), .Y(new_n18635_));
  OR2X1    g16199(.A(new_n18554_), .B(new_n14239_), .Y(new_n18636_));
  OR2X1    g16200(.A(new_n18521_), .B(new_n14244_), .Y(new_n18637_));
  OR2X1    g16201(.A(new_n18522_), .B(new_n14242_), .Y(new_n18638_));
  NAND3X1  g16202(.A(new_n18638_), .B(new_n18637_), .C(new_n18636_), .Y(new_n18639_));
  AOI21X1  g16203(.A0(new_n18639_), .A1(pi0787), .B0(new_n18635_), .Y(new_n18640_));
  AOI22X1  g16204(.A0(new_n18640_), .A1(new_n18566_), .B0(new_n18563_), .B1(pi0790), .Y(new_n18641_));
  OR2X1    g16205(.A(new_n18641_), .B(po1038), .Y(new_n18642_));
  AOI21X1  g16206(.A0(po1038), .A1(new_n6802_), .B0(pi0832), .Y(new_n18643_));
  AOI22X1  g16207(.A0(new_n18643_), .A1(new_n18642_), .B0(new_n18492_), .B1(new_n18491_), .Y(po0340));
  AOI21X1  g16208(.A0(pi1093), .A1(pi1092), .B0(pi0184), .Y(new_n18645_));
  INVX1    g16209(.A(new_n18645_), .Y(new_n18646_));
  AOI21X1  g16210(.A0(new_n12056_), .A1(new_n15193_), .B0(new_n18645_), .Y(new_n18647_));
  INVX1    g16211(.A(new_n18647_), .Y(new_n18648_));
  NAND2X1  g16212(.A(new_n18648_), .B(new_n15771_), .Y(new_n18649_));
  AND3X1   g16213(.A(new_n12480_), .B(new_n12056_), .C(new_n15193_), .Y(new_n18650_));
  OAI21X1  g16214(.A0(new_n18650_), .A1(new_n18649_), .B0(pi1155), .Y(new_n18651_));
  NOR3X1   g16215(.A(new_n18650_), .B(new_n18645_), .C(pi1155), .Y(new_n18652_));
  INVX1    g16216(.A(new_n18652_), .Y(new_n18653_));
  AOI21X1  g16217(.A0(new_n18653_), .A1(new_n18651_), .B0(new_n11768_), .Y(new_n18654_));
  AOI21X1  g16218(.A0(new_n18649_), .A1(new_n11768_), .B0(new_n18654_), .Y(new_n18655_));
  AOI21X1  g16219(.A0(new_n18655_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n18656_));
  AOI21X1  g16220(.A0(new_n18655_), .A1(new_n12655_), .B0(pi1154), .Y(new_n18657_));
  NOR2X1   g16221(.A(new_n18657_), .B(new_n18656_), .Y(new_n18658_));
  MX2X1    g16222(.A(new_n18658_), .B(new_n18655_), .S0(new_n11767_), .Y(new_n18659_));
  NOR2X1   g16223(.A(new_n18659_), .B(pi0789), .Y(new_n18660_));
  AOI21X1  g16224(.A0(new_n18659_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n18661_));
  AOI21X1  g16225(.A0(new_n18659_), .A1(new_n15790_), .B0(pi1159), .Y(new_n18662_));
  OR2X1    g16226(.A(new_n18662_), .B(new_n18661_), .Y(new_n18663_));
  AOI21X1  g16227(.A0(new_n18663_), .A1(pi0789), .B0(new_n18660_), .Y(new_n18664_));
  INVX1    g16228(.A(new_n18664_), .Y(new_n18665_));
  MX2X1    g16229(.A(new_n18665_), .B(new_n18646_), .S0(new_n12708_), .Y(new_n18666_));
  MX2X1    g16230(.A(new_n18666_), .B(new_n18646_), .S0(new_n12580_), .Y(new_n18667_));
  AOI21X1  g16231(.A0(new_n12439_), .A1(new_n15220_), .B0(new_n18645_), .Y(new_n18668_));
  OR2X1    g16232(.A(new_n18668_), .B(pi0778), .Y(new_n18669_));
  INVX1    g16233(.A(new_n18668_), .Y(new_n18670_));
  AND3X1   g16234(.A(new_n12439_), .B(new_n15220_), .C(new_n12363_), .Y(new_n18671_));
  INVX1    g16235(.A(new_n18671_), .Y(new_n18672_));
  AOI21X1  g16236(.A0(new_n18672_), .A1(new_n18670_), .B0(new_n12364_), .Y(new_n18673_));
  NOR3X1   g16237(.A(new_n18671_), .B(new_n18645_), .C(pi1153), .Y(new_n18674_));
  OR3X1    g16238(.A(new_n18674_), .B(new_n18673_), .C(new_n11769_), .Y(new_n18675_));
  AND2X1   g16239(.A(new_n18675_), .B(new_n18669_), .Y(new_n18676_));
  NOR4X1   g16240(.A(new_n18676_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n18677_));
  AND3X1   g16241(.A(new_n18677_), .B(new_n12739_), .C(new_n12718_), .Y(new_n18678_));
  INVX1    g16242(.A(new_n18678_), .Y(new_n18679_));
  AOI21X1  g16243(.A0(new_n18645_), .A1(pi0647), .B0(pi1157), .Y(new_n18680_));
  OAI21X1  g16244(.A0(new_n18679_), .A1(pi0647), .B0(new_n18680_), .Y(new_n18681_));
  MX2X1    g16245(.A(new_n18678_), .B(new_n18645_), .S0(new_n12577_), .Y(new_n18682_));
  OAI22X1  g16246(.A0(new_n18682_), .A1(new_n14242_), .B0(new_n18681_), .B1(new_n12592_), .Y(new_n18683_));
  AOI21X1  g16247(.A0(new_n18667_), .A1(new_n14326_), .B0(new_n18683_), .Y(new_n18684_));
  NOR2X1   g16248(.A(new_n18684_), .B(new_n11763_), .Y(new_n18685_));
  AOI21X1  g16249(.A0(new_n18646_), .A1(pi0626), .B0(new_n16218_), .Y(new_n18686_));
  OAI21X1  g16250(.A0(new_n18664_), .A1(pi0626), .B0(new_n18686_), .Y(new_n18687_));
  AOI21X1  g16251(.A0(new_n18646_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n18688_));
  OAI21X1  g16252(.A0(new_n18664_), .A1(new_n12542_), .B0(new_n18688_), .Y(new_n18689_));
  NAND2X1  g16253(.A(new_n18677_), .B(new_n12637_), .Y(new_n18690_));
  AND3X1   g16254(.A(new_n18690_), .B(new_n18689_), .C(new_n18687_), .Y(new_n18691_));
  NOR2X1   g16255(.A(new_n18691_), .B(new_n11765_), .Y(new_n18692_));
  NOR2X1   g16256(.A(new_n18645_), .B(pi1153), .Y(new_n18693_));
  NOR3X1   g16257(.A(new_n18668_), .B(new_n11991_), .C(new_n12363_), .Y(new_n18694_));
  AOI21X1  g16258(.A0(new_n18670_), .A1(new_n12048_), .B0(new_n18648_), .Y(new_n18695_));
  OAI21X1  g16259(.A0(new_n18695_), .A1(new_n18694_), .B0(new_n18693_), .Y(new_n18696_));
  NOR2X1   g16260(.A(new_n18673_), .B(pi0608), .Y(new_n18697_));
  NOR3X1   g16261(.A(new_n18694_), .B(new_n18648_), .C(new_n12364_), .Y(new_n18698_));
  NOR3X1   g16262(.A(new_n18698_), .B(new_n18674_), .C(new_n12368_), .Y(new_n18699_));
  AOI21X1  g16263(.A0(new_n18697_), .A1(new_n18696_), .B0(new_n18699_), .Y(new_n18700_));
  OR2X1    g16264(.A(new_n18695_), .B(pi0778), .Y(new_n18701_));
  OAI21X1  g16265(.A0(new_n18700_), .A1(new_n11769_), .B0(new_n18701_), .Y(new_n18702_));
  INVX1    g16266(.A(new_n18702_), .Y(new_n18703_));
  AND2X1   g16267(.A(new_n18702_), .B(new_n12462_), .Y(new_n18704_));
  OAI21X1  g16268(.A0(new_n18676_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n18705_));
  OR2X1    g16269(.A(new_n18705_), .B(new_n18704_), .Y(new_n18706_));
  AND3X1   g16270(.A(new_n18706_), .B(new_n18651_), .C(new_n12468_), .Y(new_n18707_));
  OAI21X1  g16271(.A0(new_n18676_), .A1(pi0609), .B0(pi1155), .Y(new_n18708_));
  AOI21X1  g16272(.A0(new_n18702_), .A1(pi0609), .B0(new_n18708_), .Y(new_n18709_));
  NOR3X1   g16273(.A(new_n18709_), .B(new_n18652_), .C(new_n12468_), .Y(new_n18710_));
  NOR2X1   g16274(.A(new_n18710_), .B(new_n18707_), .Y(new_n18711_));
  MX2X1    g16275(.A(new_n18711_), .B(new_n18703_), .S0(new_n11768_), .Y(new_n18712_));
  AOI21X1  g16276(.A0(new_n18675_), .A1(new_n18669_), .B0(new_n12630_), .Y(new_n18713_));
  AOI21X1  g16277(.A0(new_n18713_), .A1(pi0618), .B0(pi1154), .Y(new_n18714_));
  OAI21X1  g16278(.A0(new_n18712_), .A1(pi0618), .B0(new_n18714_), .Y(new_n18715_));
  NOR2X1   g16279(.A(new_n18656_), .B(pi0627), .Y(new_n18716_));
  AOI21X1  g16280(.A0(new_n18713_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18717_));
  OAI21X1  g16281(.A0(new_n18712_), .A1(new_n12486_), .B0(new_n18717_), .Y(new_n18718_));
  NOR2X1   g16282(.A(new_n18657_), .B(new_n12494_), .Y(new_n18719_));
  AOI22X1  g16283(.A0(new_n18719_), .A1(new_n18718_), .B0(new_n18716_), .B1(new_n18715_), .Y(new_n18720_));
  MX2X1    g16284(.A(new_n18720_), .B(new_n18712_), .S0(new_n11767_), .Y(new_n18721_));
  OR4X1    g16285(.A(new_n18676_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n18722_));
  AND2X1   g16286(.A(new_n18722_), .B(new_n12510_), .Y(new_n18723_));
  OAI21X1  g16287(.A0(new_n18721_), .A1(pi0619), .B0(new_n18723_), .Y(new_n18724_));
  NOR2X1   g16288(.A(new_n18661_), .B(pi0648), .Y(new_n18725_));
  AND2X1   g16289(.A(new_n18725_), .B(new_n18724_), .Y(new_n18726_));
  NOR4X1   g16290(.A(new_n18676_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n18727_));
  NOR2X1   g16291(.A(new_n18727_), .B(new_n12510_), .Y(new_n18728_));
  OAI21X1  g16292(.A0(new_n18721_), .A1(new_n12509_), .B0(new_n18728_), .Y(new_n18729_));
  NOR2X1   g16293(.A(new_n18662_), .B(new_n12517_), .Y(new_n18730_));
  AND2X1   g16294(.A(new_n18730_), .B(new_n18729_), .Y(new_n18731_));
  OR3X1    g16295(.A(new_n18731_), .B(new_n18726_), .C(new_n11766_), .Y(new_n18732_));
  AOI21X1  g16296(.A0(new_n18721_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n18733_));
  AOI21X1  g16297(.A0(new_n18733_), .A1(new_n18732_), .B0(new_n18692_), .Y(new_n18734_));
  OR2X1    g16298(.A(new_n18734_), .B(new_n14125_), .Y(new_n18735_));
  INVX1    g16299(.A(new_n18666_), .Y(new_n18736_));
  AND2X1   g16300(.A(new_n18677_), .B(new_n12718_), .Y(new_n18737_));
  AOI22X1  g16301(.A0(new_n18737_), .A1(new_n14426_), .B0(new_n18736_), .B1(new_n12735_), .Y(new_n18738_));
  AOI22X1  g16302(.A0(new_n18737_), .A1(new_n14428_), .B0(new_n18736_), .B1(new_n12733_), .Y(new_n18739_));
  MX2X1    g16303(.A(new_n18739_), .B(new_n18738_), .S0(new_n12561_), .Y(new_n18740_));
  OAI21X1  g16304(.A0(new_n18740_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n18741_));
  INVX1    g16305(.A(new_n18741_), .Y(new_n18742_));
  AOI21X1  g16306(.A0(new_n18742_), .A1(new_n18735_), .B0(new_n18685_), .Y(new_n18743_));
  OAI21X1  g16307(.A0(new_n18682_), .A1(new_n12578_), .B0(new_n18681_), .Y(new_n18744_));
  MX2X1    g16308(.A(new_n18744_), .B(new_n18679_), .S0(new_n11763_), .Y(new_n18745_));
  OAI21X1  g16309(.A0(new_n18745_), .A1(pi0644), .B0(pi0715), .Y(new_n18746_));
  AOI21X1  g16310(.A0(new_n18743_), .A1(pi0644), .B0(new_n18746_), .Y(new_n18747_));
  OR3X1    g16311(.A(new_n18646_), .B(new_n12603_), .C(new_n11763_), .Y(new_n18748_));
  OAI21X1  g16312(.A0(new_n18667_), .A1(new_n12604_), .B0(new_n18748_), .Y(new_n18749_));
  OAI21X1  g16313(.A0(new_n18646_), .A1(pi0644), .B0(new_n12608_), .Y(new_n18750_));
  AOI21X1  g16314(.A0(new_n18749_), .A1(pi0644), .B0(new_n18750_), .Y(new_n18751_));
  OR2X1    g16315(.A(new_n18751_), .B(new_n11762_), .Y(new_n18752_));
  OAI21X1  g16316(.A0(new_n18745_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n18753_));
  AOI21X1  g16317(.A0(new_n18743_), .A1(new_n12612_), .B0(new_n18753_), .Y(new_n18754_));
  OAI21X1  g16318(.A0(new_n18646_), .A1(new_n12612_), .B0(pi0715), .Y(new_n18755_));
  AOI21X1  g16319(.A0(new_n18749_), .A1(new_n12612_), .B0(new_n18755_), .Y(new_n18756_));
  OR2X1    g16320(.A(new_n18756_), .B(pi1160), .Y(new_n18757_));
  OAI22X1  g16321(.A0(new_n18757_), .A1(new_n18754_), .B0(new_n18752_), .B1(new_n18747_), .Y(new_n18758_));
  NAND2X1  g16322(.A(new_n18758_), .B(pi0790), .Y(new_n18759_));
  AOI21X1  g16323(.A0(new_n18743_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n18760_));
  AOI21X1  g16324(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0184), .Y(new_n18761_));
  INVX1    g16325(.A(new_n18761_), .Y(new_n18762_));
  AOI21X1  g16326(.A0(new_n3103_), .A1(new_n15220_), .B0(new_n18762_), .Y(new_n18763_));
  OAI21X1  g16327(.A0(new_n12826_), .A1(new_n8634_), .B0(new_n2979_), .Y(new_n18764_));
  AOI22X1  g16328(.A0(new_n18764_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n8634_), .Y(new_n18765_));
  AOI21X1  g16329(.A0(new_n12771_), .A1(new_n8634_), .B0(new_n12441_), .Y(new_n18766_));
  NOR3X1   g16330(.A(new_n18766_), .B(new_n18765_), .C(pi0737), .Y(new_n18767_));
  NOR2X1   g16331(.A(new_n18767_), .B(new_n18763_), .Y(new_n18768_));
  INVX1    g16332(.A(new_n18768_), .Y(new_n18769_));
  AOI21X1  g16333(.A0(new_n18761_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n18770_));
  OAI21X1  g16334(.A0(new_n18768_), .A1(new_n12363_), .B0(new_n18770_), .Y(new_n18771_));
  AOI21X1  g16335(.A0(new_n18761_), .A1(pi0625), .B0(pi1153), .Y(new_n18772_));
  OAI21X1  g16336(.A0(new_n18768_), .A1(pi0625), .B0(new_n18772_), .Y(new_n18773_));
  AND2X1   g16337(.A(new_n18773_), .B(new_n18771_), .Y(new_n18774_));
  MX2X1    g16338(.A(new_n18774_), .B(new_n18769_), .S0(new_n11769_), .Y(new_n18775_));
  MX2X1    g16339(.A(new_n18775_), .B(new_n18761_), .S0(new_n12490_), .Y(new_n18776_));
  INVX1    g16340(.A(new_n18776_), .Y(new_n18777_));
  MX2X1    g16341(.A(new_n18777_), .B(new_n18762_), .S0(new_n12513_), .Y(new_n18778_));
  INVX1    g16342(.A(new_n18778_), .Y(new_n18779_));
  MX2X1    g16343(.A(new_n18779_), .B(new_n18761_), .S0(new_n12531_), .Y(new_n18780_));
  MX2X1    g16344(.A(new_n18780_), .B(new_n18761_), .S0(new_n12563_), .Y(new_n18781_));
  INVX1    g16345(.A(new_n18781_), .Y(new_n18782_));
  AOI21X1  g16346(.A0(new_n18761_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n18783_));
  OAI21X1  g16347(.A0(new_n18782_), .A1(new_n12554_), .B0(new_n18783_), .Y(new_n18784_));
  AOI21X1  g16348(.A0(new_n18761_), .A1(pi0628), .B0(pi1156), .Y(new_n18785_));
  OAI21X1  g16349(.A0(new_n18782_), .A1(pi0628), .B0(new_n18785_), .Y(new_n18786_));
  AOI21X1  g16350(.A0(new_n18786_), .A1(new_n18784_), .B0(new_n11764_), .Y(new_n18787_));
  AOI21X1  g16351(.A0(new_n18782_), .A1(new_n11764_), .B0(new_n18787_), .Y(new_n18788_));
  MX2X1    g16352(.A(new_n18788_), .B(new_n18761_), .S0(pi0647), .Y(new_n18789_));
  MX2X1    g16353(.A(new_n18788_), .B(new_n18761_), .S0(new_n12577_), .Y(new_n18790_));
  MX2X1    g16354(.A(new_n18790_), .B(new_n18789_), .S0(new_n12578_), .Y(new_n18791_));
  MX2X1    g16355(.A(new_n18791_), .B(new_n18788_), .S0(new_n11763_), .Y(new_n18792_));
  AOI21X1  g16356(.A0(new_n18792_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n18793_));
  OAI22X1  g16357(.A0(new_n14197_), .A1(pi0777), .B0(new_n12077_), .B1(pi0184), .Y(new_n18794_));
  AOI21X1  g16358(.A0(new_n16615_), .A1(pi0184), .B0(pi0777), .Y(new_n18795_));
  OAI21X1  g16359(.A0(new_n12776_), .A1(pi0184), .B0(new_n18795_), .Y(new_n18796_));
  OR3X1    g16360(.A(new_n12445_), .B(new_n15193_), .C(pi0184), .Y(new_n18797_));
  AOI21X1  g16361(.A0(new_n18797_), .A1(new_n18796_), .B0(pi0038), .Y(new_n18798_));
  AOI21X1  g16362(.A0(new_n18794_), .A1(pi0038), .B0(new_n18798_), .Y(new_n18799_));
  MX2X1    g16363(.A(new_n18799_), .B(pi0184), .S0(new_n11770_), .Y(new_n18800_));
  AND2X1   g16364(.A(new_n18800_), .B(new_n12474_), .Y(new_n18801_));
  AOI21X1  g16365(.A0(new_n18762_), .A1(new_n12473_), .B0(new_n18801_), .Y(new_n18802_));
  AOI22X1  g16366(.A0(new_n18801_), .A1(pi0609), .B0(new_n18762_), .B1(new_n12472_), .Y(new_n18803_));
  AOI22X1  g16367(.A0(new_n18801_), .A1(new_n12462_), .B0(new_n18762_), .B1(new_n12481_), .Y(new_n18804_));
  MX2X1    g16368(.A(new_n18804_), .B(new_n18803_), .S0(pi1155), .Y(new_n18805_));
  MX2X1    g16369(.A(new_n18805_), .B(new_n18802_), .S0(new_n11768_), .Y(new_n18806_));
  OAI21X1  g16370(.A0(new_n18762_), .A1(pi0618), .B0(pi1154), .Y(new_n18807_));
  AOI21X1  g16371(.A0(new_n18806_), .A1(pi0618), .B0(new_n18807_), .Y(new_n18808_));
  OAI21X1  g16372(.A0(new_n18762_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18809_));
  AOI21X1  g16373(.A0(new_n18806_), .A1(new_n12486_), .B0(new_n18809_), .Y(new_n18810_));
  NOR2X1   g16374(.A(new_n18810_), .B(new_n18808_), .Y(new_n18811_));
  MX2X1    g16375(.A(new_n18811_), .B(new_n18806_), .S0(new_n11767_), .Y(new_n18812_));
  OAI21X1  g16376(.A0(new_n18762_), .A1(pi0619), .B0(pi1159), .Y(new_n18813_));
  AOI21X1  g16377(.A0(new_n18812_), .A1(pi0619), .B0(new_n18813_), .Y(new_n18814_));
  OAI21X1  g16378(.A0(new_n18762_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n18815_));
  AOI21X1  g16379(.A0(new_n18812_), .A1(new_n12509_), .B0(new_n18815_), .Y(new_n18816_));
  NOR2X1   g16380(.A(new_n18816_), .B(new_n18814_), .Y(new_n18817_));
  MX2X1    g16381(.A(new_n18817_), .B(new_n18812_), .S0(new_n11766_), .Y(new_n18818_));
  AND2X1   g16382(.A(new_n18761_), .B(new_n12708_), .Y(new_n18819_));
  AOI21X1  g16383(.A0(new_n18818_), .A1(new_n16140_), .B0(new_n18819_), .Y(new_n18820_));
  NAND2X1  g16384(.A(new_n18761_), .B(new_n12580_), .Y(new_n18821_));
  OAI21X1  g16385(.A0(new_n18820_), .A1(new_n12580_), .B0(new_n18821_), .Y(new_n18822_));
  MX2X1    g16386(.A(new_n18822_), .B(new_n18761_), .S0(new_n12604_), .Y(new_n18823_));
  OAI21X1  g16387(.A0(new_n18762_), .A1(pi0644), .B0(new_n12608_), .Y(new_n18824_));
  AOI21X1  g16388(.A0(new_n18823_), .A1(pi0644), .B0(new_n18824_), .Y(new_n18825_));
  OR2X1    g16389(.A(new_n18825_), .B(new_n11762_), .Y(new_n18826_));
  AOI21X1  g16390(.A0(new_n18792_), .A1(pi0644), .B0(pi0715), .Y(new_n18827_));
  OAI21X1  g16391(.A0(new_n18762_), .A1(new_n12612_), .B0(pi0715), .Y(new_n18828_));
  AOI21X1  g16392(.A0(new_n18823_), .A1(new_n12612_), .B0(new_n18828_), .Y(new_n18829_));
  OR2X1    g16393(.A(new_n18829_), .B(pi1160), .Y(new_n18830_));
  OAI22X1  g16394(.A0(new_n18830_), .A1(new_n18827_), .B0(new_n18826_), .B1(new_n18793_), .Y(new_n18831_));
  OR3X1    g16395(.A(new_n18829_), .B(pi1160), .C(pi0644), .Y(new_n18832_));
  OR3X1    g16396(.A(new_n18825_), .B(new_n11762_), .C(new_n12612_), .Y(new_n18833_));
  NAND3X1  g16397(.A(new_n18833_), .B(new_n18832_), .C(pi0790), .Y(new_n18834_));
  NAND2X1  g16398(.A(new_n18820_), .B(new_n14249_), .Y(new_n18835_));
  MX2X1    g16399(.A(new_n18786_), .B(new_n18784_), .S0(new_n12561_), .Y(new_n18836_));
  AND2X1   g16400(.A(new_n18836_), .B(new_n18835_), .Y(new_n18837_));
  OR2X1    g16401(.A(new_n18837_), .B(new_n11764_), .Y(new_n18838_));
  OR2X1    g16402(.A(new_n18799_), .B(new_n15220_), .Y(new_n18839_));
  OAI21X1  g16403(.A0(new_n12213_), .A1(new_n8634_), .B0(pi0777), .Y(new_n18840_));
  AOI21X1  g16404(.A0(new_n12155_), .A1(new_n8634_), .B0(new_n18840_), .Y(new_n18841_));
  AOI21X1  g16405(.A0(new_n12788_), .A1(new_n8634_), .B0(pi0777), .Y(new_n18842_));
  OAI21X1  g16406(.A0(new_n12787_), .A1(new_n8634_), .B0(new_n18842_), .Y(new_n18843_));
  NAND2X1  g16407(.A(new_n18843_), .B(pi0039), .Y(new_n18844_));
  AND2X1   g16408(.A(new_n12332_), .B(pi0184), .Y(new_n18845_));
  OAI21X1  g16409(.A0(new_n12315_), .A1(pi0184), .B0(pi0777), .Y(new_n18846_));
  NOR4X1   g16410(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0184), .Y(new_n18847_));
  OAI21X1  g16411(.A0(new_n12800_), .A1(new_n8634_), .B0(new_n15193_), .Y(new_n18848_));
  OAI22X1  g16412(.A0(new_n18848_), .A1(new_n18847_), .B0(new_n18846_), .B1(new_n18845_), .Y(new_n18849_));
  AOI21X1  g16413(.A0(new_n18849_), .A1(new_n2939_), .B0(pi0038), .Y(new_n18850_));
  OAI21X1  g16414(.A0(new_n18844_), .A1(new_n18841_), .B0(new_n18850_), .Y(new_n18851_));
  OAI21X1  g16415(.A0(new_n12276_), .A1(pi0777), .B0(new_n13540_), .Y(new_n18852_));
  NAND2X1  g16416(.A(new_n18852_), .B(new_n8634_), .Y(new_n18853_));
  AOI21X1  g16417(.A0(new_n12056_), .A1(new_n15193_), .B0(new_n13443_), .Y(new_n18854_));
  NOR2X1   g16418(.A(new_n18854_), .B(new_n8634_), .Y(new_n18855_));
  AOI21X1  g16419(.A0(new_n18855_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n18856_));
  AOI21X1  g16420(.A0(new_n18856_), .A1(new_n18853_), .B0(pi0737), .Y(new_n18857_));
  AOI21X1  g16421(.A0(new_n18857_), .A1(new_n18851_), .B0(new_n11770_), .Y(new_n18858_));
  AOI22X1  g16422(.A0(new_n18858_), .A1(new_n18839_), .B0(new_n11770_), .B1(pi0184), .Y(new_n18859_));
  OAI21X1  g16423(.A0(new_n18800_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n18860_));
  AOI21X1  g16424(.A0(new_n18859_), .A1(new_n12363_), .B0(new_n18860_), .Y(new_n18861_));
  NAND2X1  g16425(.A(new_n18771_), .B(new_n12368_), .Y(new_n18862_));
  OAI21X1  g16426(.A0(new_n18800_), .A1(pi0625), .B0(pi1153), .Y(new_n18863_));
  AOI21X1  g16427(.A0(new_n18859_), .A1(pi0625), .B0(new_n18863_), .Y(new_n18864_));
  NAND2X1  g16428(.A(new_n18773_), .B(pi0608), .Y(new_n18865_));
  OAI22X1  g16429(.A0(new_n18865_), .A1(new_n18864_), .B0(new_n18862_), .B1(new_n18861_), .Y(new_n18866_));
  MX2X1    g16430(.A(new_n18866_), .B(new_n18859_), .S0(new_n11769_), .Y(new_n18867_));
  INVX1    g16431(.A(new_n18775_), .Y(new_n18868_));
  OAI21X1  g16432(.A0(new_n18868_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n18869_));
  AOI21X1  g16433(.A0(new_n18867_), .A1(new_n12462_), .B0(new_n18869_), .Y(new_n18870_));
  OAI21X1  g16434(.A0(new_n18803_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n18871_));
  OAI21X1  g16435(.A0(new_n18868_), .A1(pi0609), .B0(pi1155), .Y(new_n18872_));
  AOI21X1  g16436(.A0(new_n18867_), .A1(pi0609), .B0(new_n18872_), .Y(new_n18873_));
  OAI21X1  g16437(.A0(new_n18804_), .A1(pi1155), .B0(pi0660), .Y(new_n18874_));
  OAI22X1  g16438(.A0(new_n18874_), .A1(new_n18873_), .B0(new_n18871_), .B1(new_n18870_), .Y(new_n18875_));
  MX2X1    g16439(.A(new_n18875_), .B(new_n18867_), .S0(new_n11768_), .Y(new_n18876_));
  OAI21X1  g16440(.A0(new_n18777_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18877_));
  AOI21X1  g16441(.A0(new_n18876_), .A1(new_n12486_), .B0(new_n18877_), .Y(new_n18878_));
  OR2X1    g16442(.A(new_n18808_), .B(pi0627), .Y(new_n18879_));
  OAI21X1  g16443(.A0(new_n18777_), .A1(pi0618), .B0(pi1154), .Y(new_n18880_));
  AOI21X1  g16444(.A0(new_n18876_), .A1(pi0618), .B0(new_n18880_), .Y(new_n18881_));
  OR2X1    g16445(.A(new_n18810_), .B(new_n12494_), .Y(new_n18882_));
  OAI22X1  g16446(.A0(new_n18882_), .A1(new_n18881_), .B0(new_n18879_), .B1(new_n18878_), .Y(new_n18883_));
  MX2X1    g16447(.A(new_n18883_), .B(new_n18876_), .S0(new_n11767_), .Y(new_n18884_));
  NAND2X1  g16448(.A(new_n18884_), .B(new_n12509_), .Y(new_n18885_));
  AOI21X1  g16449(.A0(new_n18779_), .A1(pi0619), .B0(pi1159), .Y(new_n18886_));
  OR2X1    g16450(.A(new_n18814_), .B(pi0648), .Y(new_n18887_));
  AOI21X1  g16451(.A0(new_n18886_), .A1(new_n18885_), .B0(new_n18887_), .Y(new_n18888_));
  NAND2X1  g16452(.A(new_n18884_), .B(pi0619), .Y(new_n18889_));
  AOI21X1  g16453(.A0(new_n18779_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n18890_));
  OR2X1    g16454(.A(new_n18816_), .B(new_n12517_), .Y(new_n18891_));
  AOI21X1  g16455(.A0(new_n18890_), .A1(new_n18889_), .B0(new_n18891_), .Y(new_n18892_));
  NOR3X1   g16456(.A(new_n18892_), .B(new_n18888_), .C(new_n11766_), .Y(new_n18893_));
  OAI21X1  g16457(.A0(new_n18884_), .A1(pi0789), .B0(new_n12709_), .Y(new_n18894_));
  AOI21X1  g16458(.A0(new_n18762_), .A1(pi0626), .B0(new_n16218_), .Y(new_n18895_));
  OAI21X1  g16459(.A0(new_n18818_), .A1(pi0626), .B0(new_n18895_), .Y(new_n18896_));
  AOI21X1  g16460(.A0(new_n18762_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n18897_));
  OAI21X1  g16461(.A0(new_n18818_), .A1(new_n12542_), .B0(new_n18897_), .Y(new_n18898_));
  NAND2X1  g16462(.A(new_n18780_), .B(new_n12637_), .Y(new_n18899_));
  NAND3X1  g16463(.A(new_n18899_), .B(new_n18898_), .C(new_n18896_), .Y(new_n18900_));
  AOI21X1  g16464(.A0(new_n18900_), .A1(pi0788), .B0(new_n14125_), .Y(new_n18901_));
  OAI21X1  g16465(.A0(new_n18894_), .A1(new_n18893_), .B0(new_n18901_), .Y(new_n18902_));
  AOI21X1  g16466(.A0(new_n18902_), .A1(new_n18838_), .B0(new_n14121_), .Y(new_n18903_));
  OR2X1    g16467(.A(new_n18822_), .B(new_n14239_), .Y(new_n18904_));
  OR2X1    g16468(.A(new_n18789_), .B(new_n14244_), .Y(new_n18905_));
  OR2X1    g16469(.A(new_n18790_), .B(new_n14242_), .Y(new_n18906_));
  NAND3X1  g16470(.A(new_n18906_), .B(new_n18905_), .C(new_n18904_), .Y(new_n18907_));
  AOI21X1  g16471(.A0(new_n18907_), .A1(pi0787), .B0(new_n18903_), .Y(new_n18908_));
  AOI22X1  g16472(.A0(new_n18908_), .A1(new_n18834_), .B0(new_n18831_), .B1(pi0790), .Y(new_n18909_));
  OR2X1    g16473(.A(new_n18909_), .B(po1038), .Y(new_n18910_));
  AOI21X1  g16474(.A0(po1038), .A1(new_n8634_), .B0(pi0832), .Y(new_n18911_));
  AOI22X1  g16475(.A0(new_n18911_), .A1(new_n18910_), .B0(new_n18760_), .B1(new_n18759_), .Y(po0341));
  AOI21X1  g16476(.A0(pi1093), .A1(pi1092), .B0(pi0185), .Y(new_n18913_));
  INVX1    g16477(.A(new_n18913_), .Y(new_n18914_));
  AOI21X1  g16478(.A0(new_n12056_), .A1(new_n14678_), .B0(new_n18913_), .Y(new_n18915_));
  INVX1    g16479(.A(new_n18915_), .Y(new_n18916_));
  NAND2X1  g16480(.A(new_n18916_), .B(new_n15771_), .Y(new_n18917_));
  AND3X1   g16481(.A(new_n12480_), .B(new_n12056_), .C(new_n14678_), .Y(new_n18918_));
  OAI21X1  g16482(.A0(new_n18918_), .A1(new_n18917_), .B0(pi1155), .Y(new_n18919_));
  NOR3X1   g16483(.A(new_n18918_), .B(new_n18913_), .C(pi1155), .Y(new_n18920_));
  INVX1    g16484(.A(new_n18920_), .Y(new_n18921_));
  AOI21X1  g16485(.A0(new_n18921_), .A1(new_n18919_), .B0(new_n11768_), .Y(new_n18922_));
  AOI21X1  g16486(.A0(new_n18917_), .A1(new_n11768_), .B0(new_n18922_), .Y(new_n18923_));
  AOI21X1  g16487(.A0(new_n18923_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n18924_));
  AOI21X1  g16488(.A0(new_n18923_), .A1(new_n12655_), .B0(pi1154), .Y(new_n18925_));
  NOR2X1   g16489(.A(new_n18925_), .B(new_n18924_), .Y(new_n18926_));
  MX2X1    g16490(.A(new_n18926_), .B(new_n18923_), .S0(new_n11767_), .Y(new_n18927_));
  NOR2X1   g16491(.A(new_n18927_), .B(pi0789), .Y(new_n18928_));
  AOI21X1  g16492(.A0(new_n18927_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n18929_));
  AOI21X1  g16493(.A0(new_n18927_), .A1(new_n15790_), .B0(pi1159), .Y(new_n18930_));
  OR2X1    g16494(.A(new_n18930_), .B(new_n18929_), .Y(new_n18931_));
  AOI21X1  g16495(.A0(new_n18931_), .A1(pi0789), .B0(new_n18928_), .Y(new_n18932_));
  INVX1    g16496(.A(new_n18932_), .Y(new_n18933_));
  MX2X1    g16497(.A(new_n18933_), .B(new_n18914_), .S0(new_n12708_), .Y(new_n18934_));
  MX2X1    g16498(.A(new_n18934_), .B(new_n18914_), .S0(new_n12580_), .Y(new_n18935_));
  AOI21X1  g16499(.A0(new_n12439_), .A1(new_n14697_), .B0(new_n18913_), .Y(new_n18936_));
  OR2X1    g16500(.A(new_n18936_), .B(pi0778), .Y(new_n18937_));
  INVX1    g16501(.A(new_n18936_), .Y(new_n18938_));
  AND3X1   g16502(.A(new_n12439_), .B(new_n14697_), .C(new_n12363_), .Y(new_n18939_));
  INVX1    g16503(.A(new_n18939_), .Y(new_n18940_));
  AOI21X1  g16504(.A0(new_n18940_), .A1(new_n18938_), .B0(new_n12364_), .Y(new_n18941_));
  NOR3X1   g16505(.A(new_n18939_), .B(new_n18913_), .C(pi1153), .Y(new_n18942_));
  OR3X1    g16506(.A(new_n18942_), .B(new_n18941_), .C(new_n11769_), .Y(new_n18943_));
  AND2X1   g16507(.A(new_n18943_), .B(new_n18937_), .Y(new_n18944_));
  NOR4X1   g16508(.A(new_n18944_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n18945_));
  AND3X1   g16509(.A(new_n18945_), .B(new_n12739_), .C(new_n12718_), .Y(new_n18946_));
  INVX1    g16510(.A(new_n18946_), .Y(new_n18947_));
  AOI21X1  g16511(.A0(new_n18913_), .A1(pi0647), .B0(pi1157), .Y(new_n18948_));
  OAI21X1  g16512(.A0(new_n18947_), .A1(pi0647), .B0(new_n18948_), .Y(new_n18949_));
  MX2X1    g16513(.A(new_n18946_), .B(new_n18913_), .S0(new_n12577_), .Y(new_n18950_));
  OAI22X1  g16514(.A0(new_n18950_), .A1(new_n14242_), .B0(new_n18949_), .B1(new_n12592_), .Y(new_n18951_));
  AOI21X1  g16515(.A0(new_n18935_), .A1(new_n14326_), .B0(new_n18951_), .Y(new_n18952_));
  NOR2X1   g16516(.A(new_n18952_), .B(new_n11763_), .Y(new_n18953_));
  AOI21X1  g16517(.A0(new_n18914_), .A1(pi0626), .B0(new_n16218_), .Y(new_n18954_));
  OAI21X1  g16518(.A0(new_n18932_), .A1(pi0626), .B0(new_n18954_), .Y(new_n18955_));
  AOI21X1  g16519(.A0(new_n18914_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n18956_));
  OAI21X1  g16520(.A0(new_n18932_), .A1(new_n12542_), .B0(new_n18956_), .Y(new_n18957_));
  NAND2X1  g16521(.A(new_n18945_), .B(new_n12637_), .Y(new_n18958_));
  AND3X1   g16522(.A(new_n18958_), .B(new_n18957_), .C(new_n18955_), .Y(new_n18959_));
  NOR2X1   g16523(.A(new_n18959_), .B(new_n11765_), .Y(new_n18960_));
  NOR2X1   g16524(.A(new_n18913_), .B(pi1153), .Y(new_n18961_));
  NOR3X1   g16525(.A(new_n18936_), .B(new_n11991_), .C(new_n12363_), .Y(new_n18962_));
  AOI21X1  g16526(.A0(new_n18938_), .A1(new_n12048_), .B0(new_n18916_), .Y(new_n18963_));
  OAI21X1  g16527(.A0(new_n18963_), .A1(new_n18962_), .B0(new_n18961_), .Y(new_n18964_));
  NOR2X1   g16528(.A(new_n18941_), .B(pi0608), .Y(new_n18965_));
  NOR3X1   g16529(.A(new_n18962_), .B(new_n18916_), .C(new_n12364_), .Y(new_n18966_));
  NOR3X1   g16530(.A(new_n18966_), .B(new_n18942_), .C(new_n12368_), .Y(new_n18967_));
  AOI21X1  g16531(.A0(new_n18965_), .A1(new_n18964_), .B0(new_n18967_), .Y(new_n18968_));
  OR2X1    g16532(.A(new_n18963_), .B(pi0778), .Y(new_n18969_));
  OAI21X1  g16533(.A0(new_n18968_), .A1(new_n11769_), .B0(new_n18969_), .Y(new_n18970_));
  INVX1    g16534(.A(new_n18970_), .Y(new_n18971_));
  AND2X1   g16535(.A(new_n18970_), .B(new_n12462_), .Y(new_n18972_));
  OAI21X1  g16536(.A0(new_n18944_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n18973_));
  OR2X1    g16537(.A(new_n18973_), .B(new_n18972_), .Y(new_n18974_));
  AND3X1   g16538(.A(new_n18974_), .B(new_n18919_), .C(new_n12468_), .Y(new_n18975_));
  OAI21X1  g16539(.A0(new_n18944_), .A1(pi0609), .B0(pi1155), .Y(new_n18976_));
  AOI21X1  g16540(.A0(new_n18970_), .A1(pi0609), .B0(new_n18976_), .Y(new_n18977_));
  NOR3X1   g16541(.A(new_n18977_), .B(new_n18920_), .C(new_n12468_), .Y(new_n18978_));
  NOR2X1   g16542(.A(new_n18978_), .B(new_n18975_), .Y(new_n18979_));
  MX2X1    g16543(.A(new_n18979_), .B(new_n18971_), .S0(new_n11768_), .Y(new_n18980_));
  AOI21X1  g16544(.A0(new_n18943_), .A1(new_n18937_), .B0(new_n12630_), .Y(new_n18981_));
  AOI21X1  g16545(.A0(new_n18981_), .A1(pi0618), .B0(pi1154), .Y(new_n18982_));
  OAI21X1  g16546(.A0(new_n18980_), .A1(pi0618), .B0(new_n18982_), .Y(new_n18983_));
  NOR2X1   g16547(.A(new_n18924_), .B(pi0627), .Y(new_n18984_));
  AOI21X1  g16548(.A0(new_n18981_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n18985_));
  OAI21X1  g16549(.A0(new_n18980_), .A1(new_n12486_), .B0(new_n18985_), .Y(new_n18986_));
  NOR2X1   g16550(.A(new_n18925_), .B(new_n12494_), .Y(new_n18987_));
  AOI22X1  g16551(.A0(new_n18987_), .A1(new_n18986_), .B0(new_n18984_), .B1(new_n18983_), .Y(new_n18988_));
  MX2X1    g16552(.A(new_n18988_), .B(new_n18980_), .S0(new_n11767_), .Y(new_n18989_));
  OR4X1    g16553(.A(new_n18944_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n18990_));
  AND2X1   g16554(.A(new_n18990_), .B(new_n12510_), .Y(new_n18991_));
  OAI21X1  g16555(.A0(new_n18989_), .A1(pi0619), .B0(new_n18991_), .Y(new_n18992_));
  NOR2X1   g16556(.A(new_n18929_), .B(pi0648), .Y(new_n18993_));
  AND2X1   g16557(.A(new_n18993_), .B(new_n18992_), .Y(new_n18994_));
  NOR4X1   g16558(.A(new_n18944_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n18995_));
  NOR2X1   g16559(.A(new_n18995_), .B(new_n12510_), .Y(new_n18996_));
  OAI21X1  g16560(.A0(new_n18989_), .A1(new_n12509_), .B0(new_n18996_), .Y(new_n18997_));
  NOR2X1   g16561(.A(new_n18930_), .B(new_n12517_), .Y(new_n18998_));
  AND2X1   g16562(.A(new_n18998_), .B(new_n18997_), .Y(new_n18999_));
  OR3X1    g16563(.A(new_n18999_), .B(new_n18994_), .C(new_n11766_), .Y(new_n19000_));
  AOI21X1  g16564(.A0(new_n18989_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n19001_));
  AOI21X1  g16565(.A0(new_n19001_), .A1(new_n19000_), .B0(new_n18960_), .Y(new_n19002_));
  OR2X1    g16566(.A(new_n19002_), .B(new_n14125_), .Y(new_n19003_));
  INVX1    g16567(.A(new_n18934_), .Y(new_n19004_));
  AND2X1   g16568(.A(new_n18945_), .B(new_n12718_), .Y(new_n19005_));
  AOI22X1  g16569(.A0(new_n19005_), .A1(new_n14426_), .B0(new_n19004_), .B1(new_n12735_), .Y(new_n19006_));
  AOI22X1  g16570(.A0(new_n19005_), .A1(new_n14428_), .B0(new_n19004_), .B1(new_n12733_), .Y(new_n19007_));
  MX2X1    g16571(.A(new_n19007_), .B(new_n19006_), .S0(new_n12561_), .Y(new_n19008_));
  OAI21X1  g16572(.A0(new_n19008_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n19009_));
  INVX1    g16573(.A(new_n19009_), .Y(new_n19010_));
  AOI21X1  g16574(.A0(new_n19010_), .A1(new_n19003_), .B0(new_n18953_), .Y(new_n19011_));
  OAI21X1  g16575(.A0(new_n18950_), .A1(new_n12578_), .B0(new_n18949_), .Y(new_n19012_));
  MX2X1    g16576(.A(new_n19012_), .B(new_n18947_), .S0(new_n11763_), .Y(new_n19013_));
  OAI21X1  g16577(.A0(new_n19013_), .A1(pi0644), .B0(pi0715), .Y(new_n19014_));
  AOI21X1  g16578(.A0(new_n19011_), .A1(pi0644), .B0(new_n19014_), .Y(new_n19015_));
  OR3X1    g16579(.A(new_n18914_), .B(new_n12603_), .C(new_n11763_), .Y(new_n19016_));
  OAI21X1  g16580(.A0(new_n18935_), .A1(new_n12604_), .B0(new_n19016_), .Y(new_n19017_));
  OAI21X1  g16581(.A0(new_n18914_), .A1(pi0644), .B0(new_n12608_), .Y(new_n19018_));
  AOI21X1  g16582(.A0(new_n19017_), .A1(pi0644), .B0(new_n19018_), .Y(new_n19019_));
  OR2X1    g16583(.A(new_n19019_), .B(new_n11762_), .Y(new_n19020_));
  OAI21X1  g16584(.A0(new_n19013_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n19021_));
  AOI21X1  g16585(.A0(new_n19011_), .A1(new_n12612_), .B0(new_n19021_), .Y(new_n19022_));
  OAI21X1  g16586(.A0(new_n18914_), .A1(new_n12612_), .B0(pi0715), .Y(new_n19023_));
  AOI21X1  g16587(.A0(new_n19017_), .A1(new_n12612_), .B0(new_n19023_), .Y(new_n19024_));
  OR2X1    g16588(.A(new_n19024_), .B(pi1160), .Y(new_n19025_));
  OAI22X1  g16589(.A0(new_n19025_), .A1(new_n19022_), .B0(new_n19020_), .B1(new_n19015_), .Y(new_n19026_));
  NAND2X1  g16590(.A(new_n19026_), .B(pi0790), .Y(new_n19027_));
  AOI21X1  g16591(.A0(new_n19011_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n19028_));
  AOI21X1  g16592(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0185), .Y(new_n19029_));
  INVX1    g16593(.A(new_n19029_), .Y(new_n19030_));
  AOI21X1  g16594(.A0(new_n3103_), .A1(new_n14697_), .B0(new_n19030_), .Y(new_n19031_));
  OAI21X1  g16595(.A0(new_n12826_), .A1(new_n9902_), .B0(new_n2979_), .Y(new_n19032_));
  AOI22X1  g16596(.A0(new_n19032_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n9902_), .Y(new_n19033_));
  AOI21X1  g16597(.A0(new_n12771_), .A1(new_n9902_), .B0(new_n12441_), .Y(new_n19034_));
  NOR3X1   g16598(.A(new_n19034_), .B(new_n19033_), .C(pi0701), .Y(new_n19035_));
  NOR2X1   g16599(.A(new_n19035_), .B(new_n19031_), .Y(new_n19036_));
  INVX1    g16600(.A(new_n19036_), .Y(new_n19037_));
  AOI21X1  g16601(.A0(new_n19029_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n19038_));
  OAI21X1  g16602(.A0(new_n19036_), .A1(new_n12363_), .B0(new_n19038_), .Y(new_n19039_));
  AOI21X1  g16603(.A0(new_n19029_), .A1(pi0625), .B0(pi1153), .Y(new_n19040_));
  OAI21X1  g16604(.A0(new_n19036_), .A1(pi0625), .B0(new_n19040_), .Y(new_n19041_));
  AND2X1   g16605(.A(new_n19041_), .B(new_n19039_), .Y(new_n19042_));
  MX2X1    g16606(.A(new_n19042_), .B(new_n19037_), .S0(new_n11769_), .Y(new_n19043_));
  MX2X1    g16607(.A(new_n19043_), .B(new_n19029_), .S0(new_n12490_), .Y(new_n19044_));
  INVX1    g16608(.A(new_n19044_), .Y(new_n19045_));
  MX2X1    g16609(.A(new_n19045_), .B(new_n19030_), .S0(new_n12513_), .Y(new_n19046_));
  INVX1    g16610(.A(new_n19046_), .Y(new_n19047_));
  MX2X1    g16611(.A(new_n19047_), .B(new_n19029_), .S0(new_n12531_), .Y(new_n19048_));
  MX2X1    g16612(.A(new_n19048_), .B(new_n19029_), .S0(new_n12563_), .Y(new_n19049_));
  INVX1    g16613(.A(new_n19049_), .Y(new_n19050_));
  AOI21X1  g16614(.A0(new_n19029_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n19051_));
  OAI21X1  g16615(.A0(new_n19050_), .A1(new_n12554_), .B0(new_n19051_), .Y(new_n19052_));
  AOI21X1  g16616(.A0(new_n19029_), .A1(pi0628), .B0(pi1156), .Y(new_n19053_));
  OAI21X1  g16617(.A0(new_n19050_), .A1(pi0628), .B0(new_n19053_), .Y(new_n19054_));
  AOI21X1  g16618(.A0(new_n19054_), .A1(new_n19052_), .B0(new_n11764_), .Y(new_n19055_));
  AOI21X1  g16619(.A0(new_n19050_), .A1(new_n11764_), .B0(new_n19055_), .Y(new_n19056_));
  MX2X1    g16620(.A(new_n19056_), .B(new_n19029_), .S0(pi0647), .Y(new_n19057_));
  MX2X1    g16621(.A(new_n19056_), .B(new_n19029_), .S0(new_n12577_), .Y(new_n19058_));
  MX2X1    g16622(.A(new_n19058_), .B(new_n19057_), .S0(new_n12578_), .Y(new_n19059_));
  MX2X1    g16623(.A(new_n19059_), .B(new_n19056_), .S0(new_n11763_), .Y(new_n19060_));
  AOI21X1  g16624(.A0(new_n19060_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n19061_));
  AOI22X1  g16625(.A0(new_n12073_), .A1(pi0185), .B0(new_n12444_), .B1(pi0751), .Y(new_n19062_));
  OR3X1    g16626(.A(new_n12776_), .B(pi0751), .C(pi0185), .Y(new_n19063_));
  OAI22X1  g16627(.A0(new_n12045_), .A1(new_n9902_), .B0(new_n11822_), .B1(new_n14678_), .Y(new_n19064_));
  AOI22X1  g16628(.A0(new_n19064_), .A1(new_n2939_), .B0(pi0751), .B1(pi0185), .Y(new_n19065_));
  AND2X1   g16629(.A(new_n19065_), .B(new_n19063_), .Y(new_n19066_));
  OAI21X1  g16630(.A0(new_n19062_), .A1(new_n2939_), .B0(new_n19066_), .Y(new_n19067_));
  AND2X1   g16631(.A(new_n19067_), .B(new_n2979_), .Y(new_n19068_));
  OAI21X1  g16632(.A0(new_n12077_), .A1(pi0185), .B0(pi0038), .Y(new_n19069_));
  AOI21X1  g16633(.A0(new_n12079_), .A1(new_n14678_), .B0(new_n19069_), .Y(new_n19070_));
  OR2X1    g16634(.A(new_n19070_), .B(new_n19068_), .Y(new_n19071_));
  MX2X1    g16635(.A(new_n19071_), .B(pi0185), .S0(new_n11770_), .Y(new_n19072_));
  AND2X1   g16636(.A(new_n19072_), .B(new_n12474_), .Y(new_n19073_));
  AOI21X1  g16637(.A0(new_n19030_), .A1(new_n12473_), .B0(new_n19073_), .Y(new_n19074_));
  AOI22X1  g16638(.A0(new_n19073_), .A1(pi0609), .B0(new_n19030_), .B1(new_n12472_), .Y(new_n19075_));
  AOI22X1  g16639(.A0(new_n19073_), .A1(new_n12462_), .B0(new_n19030_), .B1(new_n12481_), .Y(new_n19076_));
  MX2X1    g16640(.A(new_n19076_), .B(new_n19075_), .S0(pi1155), .Y(new_n19077_));
  MX2X1    g16641(.A(new_n19077_), .B(new_n19074_), .S0(new_n11768_), .Y(new_n19078_));
  OAI21X1  g16642(.A0(new_n19030_), .A1(pi0618), .B0(pi1154), .Y(new_n19079_));
  AOI21X1  g16643(.A0(new_n19078_), .A1(pi0618), .B0(new_n19079_), .Y(new_n19080_));
  OAI21X1  g16644(.A0(new_n19030_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n19081_));
  AOI21X1  g16645(.A0(new_n19078_), .A1(new_n12486_), .B0(new_n19081_), .Y(new_n19082_));
  NOR2X1   g16646(.A(new_n19082_), .B(new_n19080_), .Y(new_n19083_));
  MX2X1    g16647(.A(new_n19083_), .B(new_n19078_), .S0(new_n11767_), .Y(new_n19084_));
  OAI21X1  g16648(.A0(new_n19030_), .A1(pi0619), .B0(pi1159), .Y(new_n19085_));
  AOI21X1  g16649(.A0(new_n19084_), .A1(pi0619), .B0(new_n19085_), .Y(new_n19086_));
  OAI21X1  g16650(.A0(new_n19030_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19087_));
  AOI21X1  g16651(.A0(new_n19084_), .A1(new_n12509_), .B0(new_n19087_), .Y(new_n19088_));
  NOR2X1   g16652(.A(new_n19088_), .B(new_n19086_), .Y(new_n19089_));
  MX2X1    g16653(.A(new_n19089_), .B(new_n19084_), .S0(new_n11766_), .Y(new_n19090_));
  AND2X1   g16654(.A(new_n19029_), .B(new_n12708_), .Y(new_n19091_));
  AOI21X1  g16655(.A0(new_n19090_), .A1(new_n16140_), .B0(new_n19091_), .Y(new_n19092_));
  NAND2X1  g16656(.A(new_n19029_), .B(new_n12580_), .Y(new_n19093_));
  OAI21X1  g16657(.A0(new_n19092_), .A1(new_n12580_), .B0(new_n19093_), .Y(new_n19094_));
  MX2X1    g16658(.A(new_n19094_), .B(new_n19029_), .S0(new_n12604_), .Y(new_n19095_));
  OAI21X1  g16659(.A0(new_n19030_), .A1(pi0644), .B0(new_n12608_), .Y(new_n19096_));
  AOI21X1  g16660(.A0(new_n19095_), .A1(pi0644), .B0(new_n19096_), .Y(new_n19097_));
  OR2X1    g16661(.A(new_n19097_), .B(new_n11762_), .Y(new_n19098_));
  AOI21X1  g16662(.A0(new_n19060_), .A1(pi0644), .B0(pi0715), .Y(new_n19099_));
  OAI21X1  g16663(.A0(new_n19030_), .A1(new_n12612_), .B0(pi0715), .Y(new_n19100_));
  AOI21X1  g16664(.A0(new_n19095_), .A1(new_n12612_), .B0(new_n19100_), .Y(new_n19101_));
  OR2X1    g16665(.A(new_n19101_), .B(pi1160), .Y(new_n19102_));
  OAI22X1  g16666(.A0(new_n19102_), .A1(new_n19099_), .B0(new_n19098_), .B1(new_n19061_), .Y(new_n19103_));
  OR3X1    g16667(.A(new_n19101_), .B(pi1160), .C(pi0644), .Y(new_n19104_));
  OR3X1    g16668(.A(new_n19097_), .B(new_n11762_), .C(new_n12612_), .Y(new_n19105_));
  NAND3X1  g16669(.A(new_n19105_), .B(new_n19104_), .C(pi0790), .Y(new_n19106_));
  NAND2X1  g16670(.A(new_n19092_), .B(new_n14249_), .Y(new_n19107_));
  MX2X1    g16671(.A(new_n19054_), .B(new_n19052_), .S0(new_n12561_), .Y(new_n19108_));
  AND2X1   g16672(.A(new_n19108_), .B(new_n19107_), .Y(new_n19109_));
  OR2X1    g16673(.A(new_n19109_), .B(new_n11764_), .Y(new_n19110_));
  OR3X1    g16674(.A(new_n19070_), .B(new_n19068_), .C(new_n14697_), .Y(new_n19111_));
  OAI21X1  g16675(.A0(new_n12213_), .A1(new_n9902_), .B0(pi0751), .Y(new_n19112_));
  AOI21X1  g16676(.A0(new_n12155_), .A1(new_n9902_), .B0(new_n19112_), .Y(new_n19113_));
  AOI21X1  g16677(.A0(new_n12788_), .A1(new_n9902_), .B0(pi0751), .Y(new_n19114_));
  OAI21X1  g16678(.A0(new_n12787_), .A1(new_n9902_), .B0(new_n19114_), .Y(new_n19115_));
  NAND2X1  g16679(.A(new_n19115_), .B(pi0039), .Y(new_n19116_));
  AND2X1   g16680(.A(new_n12332_), .B(pi0185), .Y(new_n19117_));
  OAI21X1  g16681(.A0(new_n12315_), .A1(pi0185), .B0(pi0751), .Y(new_n19118_));
  NOR4X1   g16682(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0185), .Y(new_n19119_));
  OAI21X1  g16683(.A0(new_n12800_), .A1(new_n9902_), .B0(new_n14678_), .Y(new_n19120_));
  OAI22X1  g16684(.A0(new_n19120_), .A1(new_n19119_), .B0(new_n19118_), .B1(new_n19117_), .Y(new_n19121_));
  AOI21X1  g16685(.A0(new_n19121_), .A1(new_n2939_), .B0(pi0038), .Y(new_n19122_));
  OAI21X1  g16686(.A0(new_n19116_), .A1(new_n19113_), .B0(new_n19122_), .Y(new_n19123_));
  OAI21X1  g16687(.A0(new_n12276_), .A1(pi0751), .B0(new_n13540_), .Y(new_n19124_));
  NAND2X1  g16688(.A(new_n19124_), .B(new_n9902_), .Y(new_n19125_));
  AOI21X1  g16689(.A0(new_n12056_), .A1(new_n14678_), .B0(new_n13443_), .Y(new_n19126_));
  NOR2X1   g16690(.A(new_n19126_), .B(new_n9902_), .Y(new_n19127_));
  AOI21X1  g16691(.A0(new_n19127_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n19128_));
  AOI21X1  g16692(.A0(new_n19128_), .A1(new_n19125_), .B0(pi0701), .Y(new_n19129_));
  AOI21X1  g16693(.A0(new_n19129_), .A1(new_n19123_), .B0(new_n11770_), .Y(new_n19130_));
  AOI22X1  g16694(.A0(new_n19130_), .A1(new_n19111_), .B0(new_n11770_), .B1(pi0185), .Y(new_n19131_));
  AND2X1   g16695(.A(new_n19131_), .B(new_n12363_), .Y(new_n19132_));
  OAI21X1  g16696(.A0(new_n19072_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n19133_));
  OR2X1    g16697(.A(new_n19133_), .B(new_n19132_), .Y(new_n19134_));
  NAND3X1  g16698(.A(new_n19134_), .B(new_n19039_), .C(new_n12368_), .Y(new_n19135_));
  AND2X1   g16699(.A(new_n19131_), .B(pi0625), .Y(new_n19136_));
  OAI21X1  g16700(.A0(new_n19072_), .A1(pi0625), .B0(pi1153), .Y(new_n19137_));
  OR2X1    g16701(.A(new_n19137_), .B(new_n19136_), .Y(new_n19138_));
  NAND3X1  g16702(.A(new_n19138_), .B(new_n19041_), .C(pi0608), .Y(new_n19139_));
  NAND2X1  g16703(.A(new_n19139_), .B(new_n19135_), .Y(new_n19140_));
  MX2X1    g16704(.A(new_n19140_), .B(new_n19131_), .S0(new_n11769_), .Y(new_n19141_));
  INVX1    g16705(.A(new_n19043_), .Y(new_n19142_));
  OAI21X1  g16706(.A0(new_n19142_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n19143_));
  AOI21X1  g16707(.A0(new_n19141_), .A1(new_n12462_), .B0(new_n19143_), .Y(new_n19144_));
  OAI21X1  g16708(.A0(new_n19075_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n19145_));
  OAI21X1  g16709(.A0(new_n19142_), .A1(pi0609), .B0(pi1155), .Y(new_n19146_));
  AOI21X1  g16710(.A0(new_n19141_), .A1(pi0609), .B0(new_n19146_), .Y(new_n19147_));
  OAI21X1  g16711(.A0(new_n19076_), .A1(pi1155), .B0(pi0660), .Y(new_n19148_));
  OAI22X1  g16712(.A0(new_n19148_), .A1(new_n19147_), .B0(new_n19145_), .B1(new_n19144_), .Y(new_n19149_));
  MX2X1    g16713(.A(new_n19149_), .B(new_n19141_), .S0(new_n11768_), .Y(new_n19150_));
  OAI21X1  g16714(.A0(new_n19045_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n19151_));
  AOI21X1  g16715(.A0(new_n19150_), .A1(new_n12486_), .B0(new_n19151_), .Y(new_n19152_));
  OR2X1    g16716(.A(new_n19080_), .B(pi0627), .Y(new_n19153_));
  OAI21X1  g16717(.A0(new_n19045_), .A1(pi0618), .B0(pi1154), .Y(new_n19154_));
  AOI21X1  g16718(.A0(new_n19150_), .A1(pi0618), .B0(new_n19154_), .Y(new_n19155_));
  OR2X1    g16719(.A(new_n19082_), .B(new_n12494_), .Y(new_n19156_));
  OAI22X1  g16720(.A0(new_n19156_), .A1(new_n19155_), .B0(new_n19153_), .B1(new_n19152_), .Y(new_n19157_));
  MX2X1    g16721(.A(new_n19157_), .B(new_n19150_), .S0(new_n11767_), .Y(new_n19158_));
  NAND2X1  g16722(.A(new_n19158_), .B(new_n12509_), .Y(new_n19159_));
  AOI21X1  g16723(.A0(new_n19047_), .A1(pi0619), .B0(pi1159), .Y(new_n19160_));
  OR2X1    g16724(.A(new_n19086_), .B(pi0648), .Y(new_n19161_));
  AOI21X1  g16725(.A0(new_n19160_), .A1(new_n19159_), .B0(new_n19161_), .Y(new_n19162_));
  NAND2X1  g16726(.A(new_n19158_), .B(pi0619), .Y(new_n19163_));
  AOI21X1  g16727(.A0(new_n19047_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19164_));
  OR2X1    g16728(.A(new_n19088_), .B(new_n12517_), .Y(new_n19165_));
  AOI21X1  g16729(.A0(new_n19164_), .A1(new_n19163_), .B0(new_n19165_), .Y(new_n19166_));
  NOR3X1   g16730(.A(new_n19166_), .B(new_n19162_), .C(new_n11766_), .Y(new_n19167_));
  OAI21X1  g16731(.A0(new_n19158_), .A1(pi0789), .B0(new_n12709_), .Y(new_n19168_));
  AOI21X1  g16732(.A0(new_n19030_), .A1(pi0626), .B0(new_n16218_), .Y(new_n19169_));
  OAI21X1  g16733(.A0(new_n19090_), .A1(pi0626), .B0(new_n19169_), .Y(new_n19170_));
  AOI21X1  g16734(.A0(new_n19030_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n19171_));
  OAI21X1  g16735(.A0(new_n19090_), .A1(new_n12542_), .B0(new_n19171_), .Y(new_n19172_));
  NAND2X1  g16736(.A(new_n19048_), .B(new_n12637_), .Y(new_n19173_));
  NAND3X1  g16737(.A(new_n19173_), .B(new_n19172_), .C(new_n19170_), .Y(new_n19174_));
  AOI21X1  g16738(.A0(new_n19174_), .A1(pi0788), .B0(new_n14125_), .Y(new_n19175_));
  OAI21X1  g16739(.A0(new_n19168_), .A1(new_n19167_), .B0(new_n19175_), .Y(new_n19176_));
  AOI21X1  g16740(.A0(new_n19176_), .A1(new_n19110_), .B0(new_n14121_), .Y(new_n19177_));
  OR2X1    g16741(.A(new_n19094_), .B(new_n14239_), .Y(new_n19178_));
  OR2X1    g16742(.A(new_n19057_), .B(new_n14244_), .Y(new_n19179_));
  OR2X1    g16743(.A(new_n19058_), .B(new_n14242_), .Y(new_n19180_));
  NAND3X1  g16744(.A(new_n19180_), .B(new_n19179_), .C(new_n19178_), .Y(new_n19181_));
  AOI21X1  g16745(.A0(new_n19181_), .A1(pi0787), .B0(new_n19177_), .Y(new_n19182_));
  AOI22X1  g16746(.A0(new_n19182_), .A1(new_n19106_), .B0(new_n19103_), .B1(pi0790), .Y(new_n19183_));
  OR2X1    g16747(.A(new_n19183_), .B(po1038), .Y(new_n19184_));
  AOI21X1  g16748(.A0(po1038), .A1(new_n9902_), .B0(pi0832), .Y(new_n19185_));
  AOI22X1  g16749(.A0(new_n19185_), .A1(new_n19184_), .B0(new_n19028_), .B1(new_n19027_), .Y(po0342));
  NOR2X1   g16750(.A(new_n13547_), .B(new_n15235_), .Y(new_n19187_));
  OAI21X1  g16751(.A0(new_n13545_), .A1(new_n6818_), .B0(new_n19187_), .Y(new_n19188_));
  AOI21X1  g16752(.A0(new_n13543_), .A1(new_n6818_), .B0(new_n19188_), .Y(new_n19189_));
  OAI21X1  g16753(.A0(new_n13559_), .A1(pi0186), .B0(new_n15235_), .Y(new_n19190_));
  AOI21X1  g16754(.A0(new_n13554_), .A1(pi0186), .B0(new_n19190_), .Y(new_n19191_));
  OR3X1    g16755(.A(new_n19191_), .B(new_n19189_), .C(new_n15229_), .Y(new_n19192_));
  OAI21X1  g16756(.A0(new_n12447_), .A1(pi0186), .B0(pi0752), .Y(new_n19193_));
  AOI21X1  g16757(.A0(new_n12074_), .A1(new_n2979_), .B0(new_n6818_), .Y(new_n19194_));
  NOR2X1   g16758(.A(pi0752), .B(pi0186), .Y(new_n19195_));
  AOI21X1  g16759(.A0(new_n19195_), .A1(new_n13568_), .B0(new_n19194_), .Y(new_n19196_));
  OR2X1    g16760(.A(new_n19196_), .B(new_n13565_), .Y(new_n19197_));
  AND2X1   g16761(.A(new_n19197_), .B(new_n19193_), .Y(new_n19198_));
  AOI21X1  g16762(.A0(new_n19198_), .A1(new_n15229_), .B0(new_n11770_), .Y(new_n19199_));
  AOI22X1  g16763(.A0(new_n19199_), .A1(new_n19192_), .B0(new_n11770_), .B1(pi0186), .Y(new_n19200_));
  NAND2X1  g16764(.A(new_n19197_), .B(new_n19193_), .Y(new_n19201_));
  MX2X1    g16765(.A(new_n19201_), .B(pi0186), .S0(new_n11770_), .Y(new_n19202_));
  OAI21X1  g16766(.A0(new_n19202_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n19203_));
  AOI21X1  g16767(.A0(new_n19200_), .A1(new_n12363_), .B0(new_n19203_), .Y(new_n19204_));
  AND3X1   g16768(.A(new_n12832_), .B(new_n15229_), .C(new_n6818_), .Y(new_n19205_));
  OAI21X1  g16769(.A0(new_n12826_), .A1(new_n6818_), .B0(new_n2979_), .Y(new_n19206_));
  AOI21X1  g16770(.A0(new_n12825_), .A1(new_n6818_), .B0(new_n19206_), .Y(new_n19207_));
  OAI21X1  g16771(.A0(new_n12077_), .A1(pi0186), .B0(new_n12440_), .Y(new_n19208_));
  NAND2X1  g16772(.A(new_n19208_), .B(pi0703), .Y(new_n19209_));
  OAI21X1  g16773(.A0(new_n19209_), .A1(new_n19207_), .B0(new_n3103_), .Y(new_n19210_));
  OAI22X1  g16774(.A0(new_n19210_), .A1(new_n19205_), .B0(new_n3103_), .B1(new_n6818_), .Y(new_n19211_));
  AOI21X1  g16775(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0186), .Y(new_n19212_));
  AOI21X1  g16776(.A0(new_n19212_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n19213_));
  OAI21X1  g16777(.A0(new_n19211_), .A1(new_n12363_), .B0(new_n19213_), .Y(new_n19214_));
  NAND2X1  g16778(.A(new_n19214_), .B(new_n12368_), .Y(new_n19215_));
  OAI21X1  g16779(.A0(new_n19202_), .A1(pi0625), .B0(pi1153), .Y(new_n19216_));
  AOI21X1  g16780(.A0(new_n19200_), .A1(pi0625), .B0(new_n19216_), .Y(new_n19217_));
  AOI21X1  g16781(.A0(new_n19212_), .A1(pi0625), .B0(pi1153), .Y(new_n19218_));
  OAI21X1  g16782(.A0(new_n19211_), .A1(pi0625), .B0(new_n19218_), .Y(new_n19219_));
  NAND2X1  g16783(.A(new_n19219_), .B(pi0608), .Y(new_n19220_));
  OAI22X1  g16784(.A0(new_n19220_), .A1(new_n19217_), .B0(new_n19215_), .B1(new_n19204_), .Y(new_n19221_));
  MX2X1    g16785(.A(new_n19221_), .B(new_n19200_), .S0(new_n11769_), .Y(new_n19222_));
  NAND2X1  g16786(.A(new_n19219_), .B(new_n19214_), .Y(new_n19223_));
  MX2X1    g16787(.A(new_n19223_), .B(new_n19211_), .S0(new_n11769_), .Y(new_n19224_));
  OAI21X1  g16788(.A0(new_n19224_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n19225_));
  AOI21X1  g16789(.A0(new_n19222_), .A1(new_n12462_), .B0(new_n19225_), .Y(new_n19226_));
  NOR2X1   g16790(.A(new_n19212_), .B(new_n12471_), .Y(new_n19227_));
  AND3X1   g16791(.A(new_n19202_), .B(new_n12474_), .C(pi0609), .Y(new_n19228_));
  OAI21X1  g16792(.A0(new_n19228_), .A1(new_n19227_), .B0(pi1155), .Y(new_n19229_));
  NAND2X1  g16793(.A(new_n19229_), .B(new_n12468_), .Y(new_n19230_));
  OAI21X1  g16794(.A0(new_n19224_), .A1(pi0609), .B0(pi1155), .Y(new_n19231_));
  AOI21X1  g16795(.A0(new_n19222_), .A1(pi0609), .B0(new_n19231_), .Y(new_n19232_));
  INVX1    g16796(.A(new_n19212_), .Y(new_n19233_));
  AND3X1   g16797(.A(new_n19202_), .B(new_n12474_), .C(new_n12462_), .Y(new_n19234_));
  AOI21X1  g16798(.A0(new_n19233_), .A1(new_n12481_), .B0(new_n19234_), .Y(new_n19235_));
  OAI21X1  g16799(.A0(new_n19235_), .A1(pi1155), .B0(pi0660), .Y(new_n19236_));
  OAI22X1  g16800(.A0(new_n19236_), .A1(new_n19232_), .B0(new_n19230_), .B1(new_n19226_), .Y(new_n19237_));
  MX2X1    g16801(.A(new_n19237_), .B(new_n19222_), .S0(new_n11768_), .Y(new_n19238_));
  MX2X1    g16802(.A(new_n19224_), .B(new_n19233_), .S0(new_n12490_), .Y(new_n19239_));
  OAI21X1  g16803(.A0(new_n19239_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n19240_));
  AOI21X1  g16804(.A0(new_n19238_), .A1(new_n12486_), .B0(new_n19240_), .Y(new_n19241_));
  MX2X1    g16805(.A(new_n19233_), .B(new_n19202_), .S0(new_n12474_), .Y(new_n19242_));
  AND2X1   g16806(.A(new_n19242_), .B(new_n11768_), .Y(new_n19243_));
  OAI21X1  g16807(.A0(new_n19235_), .A1(pi1155), .B0(new_n19229_), .Y(new_n19244_));
  AOI21X1  g16808(.A0(new_n19244_), .A1(pi0785), .B0(new_n19243_), .Y(new_n19245_));
  OAI21X1  g16809(.A0(new_n19233_), .A1(pi0618), .B0(pi1154), .Y(new_n19246_));
  AOI21X1  g16810(.A0(new_n19245_), .A1(pi0618), .B0(new_n19246_), .Y(new_n19247_));
  OR2X1    g16811(.A(new_n19247_), .B(pi0627), .Y(new_n19248_));
  OAI21X1  g16812(.A0(new_n19239_), .A1(pi0618), .B0(pi1154), .Y(new_n19249_));
  AOI21X1  g16813(.A0(new_n19238_), .A1(pi0618), .B0(new_n19249_), .Y(new_n19250_));
  OAI21X1  g16814(.A0(new_n19233_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n19251_));
  AOI21X1  g16815(.A0(new_n19245_), .A1(new_n12486_), .B0(new_n19251_), .Y(new_n19252_));
  OR2X1    g16816(.A(new_n19252_), .B(new_n12494_), .Y(new_n19253_));
  OAI22X1  g16817(.A0(new_n19253_), .A1(new_n19250_), .B0(new_n19248_), .B1(new_n19241_), .Y(new_n19254_));
  MX2X1    g16818(.A(new_n19254_), .B(new_n19238_), .S0(new_n11767_), .Y(new_n19255_));
  MX2X1    g16819(.A(new_n19239_), .B(new_n19233_), .S0(new_n12513_), .Y(new_n19256_));
  OAI21X1  g16820(.A0(new_n19256_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19257_));
  AOI21X1  g16821(.A0(new_n19255_), .A1(new_n12509_), .B0(new_n19257_), .Y(new_n19258_));
  NOR2X1   g16822(.A(new_n19252_), .B(new_n19247_), .Y(new_n19259_));
  MX2X1    g16823(.A(new_n19259_), .B(new_n19245_), .S0(new_n11767_), .Y(new_n19260_));
  OAI21X1  g16824(.A0(new_n19233_), .A1(pi0619), .B0(pi1159), .Y(new_n19261_));
  AOI21X1  g16825(.A0(new_n19260_), .A1(pi0619), .B0(new_n19261_), .Y(new_n19262_));
  OR2X1    g16826(.A(new_n19262_), .B(pi0648), .Y(new_n19263_));
  OAI21X1  g16827(.A0(new_n19256_), .A1(pi0619), .B0(pi1159), .Y(new_n19264_));
  AOI21X1  g16828(.A0(new_n19255_), .A1(pi0619), .B0(new_n19264_), .Y(new_n19265_));
  OAI21X1  g16829(.A0(new_n19233_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19266_));
  AOI21X1  g16830(.A0(new_n19260_), .A1(new_n12509_), .B0(new_n19266_), .Y(new_n19267_));
  OR2X1    g16831(.A(new_n19267_), .B(new_n12517_), .Y(new_n19268_));
  OAI22X1  g16832(.A0(new_n19268_), .A1(new_n19265_), .B0(new_n19263_), .B1(new_n19258_), .Y(new_n19269_));
  MX2X1    g16833(.A(new_n19269_), .B(new_n19255_), .S0(new_n11766_), .Y(new_n19270_));
  MX2X1    g16834(.A(new_n19256_), .B(new_n19233_), .S0(new_n12531_), .Y(new_n19271_));
  AOI21X1  g16835(.A0(new_n19271_), .A1(pi0626), .B0(pi0641), .Y(new_n19272_));
  OAI21X1  g16836(.A0(new_n19270_), .A1(pi0626), .B0(new_n19272_), .Y(new_n19273_));
  OR2X1    g16837(.A(new_n19260_), .B(pi0789), .Y(new_n19274_));
  OAI21X1  g16838(.A0(new_n19267_), .A1(new_n19262_), .B0(pi0789), .Y(new_n19275_));
  NAND2X1  g16839(.A(new_n19275_), .B(new_n19274_), .Y(new_n19276_));
  NAND2X1  g16840(.A(new_n19276_), .B(new_n12542_), .Y(new_n19277_));
  AOI21X1  g16841(.A0(new_n19233_), .A1(pi0626), .B0(new_n12543_), .Y(new_n19278_));
  AOI21X1  g16842(.A0(new_n19278_), .A1(new_n19277_), .B0(pi1158), .Y(new_n19279_));
  AOI21X1  g16843(.A0(new_n19271_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n19280_));
  OAI21X1  g16844(.A0(new_n19270_), .A1(new_n12542_), .B0(new_n19280_), .Y(new_n19281_));
  NAND2X1  g16845(.A(new_n19276_), .B(pi0626), .Y(new_n19282_));
  AOI21X1  g16846(.A0(new_n19233_), .A1(new_n12542_), .B0(pi0641), .Y(new_n19283_));
  AOI21X1  g16847(.A0(new_n19283_), .A1(new_n19282_), .B0(new_n12548_), .Y(new_n19284_));
  AOI22X1  g16848(.A0(new_n19284_), .A1(new_n19281_), .B0(new_n19279_), .B1(new_n19273_), .Y(new_n19285_));
  MX2X1    g16849(.A(new_n19285_), .B(new_n19270_), .S0(new_n11765_), .Y(new_n19286_));
  MX2X1    g16850(.A(new_n19276_), .B(new_n19233_), .S0(new_n12708_), .Y(new_n19287_));
  OAI21X1  g16851(.A0(new_n19287_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n19288_));
  AOI21X1  g16852(.A0(new_n19286_), .A1(new_n12554_), .B0(new_n19288_), .Y(new_n19289_));
  MX2X1    g16853(.A(new_n19271_), .B(new_n19233_), .S0(new_n12563_), .Y(new_n19290_));
  AOI21X1  g16854(.A0(new_n19212_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n19291_));
  OAI21X1  g16855(.A0(new_n19290_), .A1(new_n12554_), .B0(new_n19291_), .Y(new_n19292_));
  AND2X1   g16856(.A(new_n19292_), .B(new_n12561_), .Y(new_n19293_));
  INVX1    g16857(.A(new_n19293_), .Y(new_n19294_));
  OAI21X1  g16858(.A0(new_n19287_), .A1(pi0628), .B0(pi1156), .Y(new_n19295_));
  AOI21X1  g16859(.A0(new_n19286_), .A1(pi0628), .B0(new_n19295_), .Y(new_n19296_));
  AOI21X1  g16860(.A0(new_n19212_), .A1(pi0628), .B0(pi1156), .Y(new_n19297_));
  OAI21X1  g16861(.A0(new_n19290_), .A1(pi0628), .B0(new_n19297_), .Y(new_n19298_));
  AND2X1   g16862(.A(new_n19298_), .B(pi0629), .Y(new_n19299_));
  INVX1    g16863(.A(new_n19299_), .Y(new_n19300_));
  OAI22X1  g16864(.A0(new_n19300_), .A1(new_n19296_), .B0(new_n19294_), .B1(new_n19289_), .Y(new_n19301_));
  MX2X1    g16865(.A(new_n19301_), .B(new_n19286_), .S0(new_n11764_), .Y(new_n19302_));
  MX2X1    g16866(.A(new_n19287_), .B(new_n19233_), .S0(new_n12580_), .Y(new_n19303_));
  OAI21X1  g16867(.A0(new_n19303_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n19304_));
  AOI21X1  g16868(.A0(new_n19302_), .A1(new_n12577_), .B0(new_n19304_), .Y(new_n19305_));
  AOI21X1  g16869(.A0(new_n19298_), .A1(new_n19292_), .B0(new_n11764_), .Y(new_n19306_));
  AOI21X1  g16870(.A0(new_n19290_), .A1(new_n11764_), .B0(new_n19306_), .Y(new_n19307_));
  OAI21X1  g16871(.A0(new_n19233_), .A1(pi0647), .B0(pi1157), .Y(new_n19308_));
  AOI21X1  g16872(.A0(new_n19307_), .A1(pi0647), .B0(new_n19308_), .Y(new_n19309_));
  NOR2X1   g16873(.A(new_n19309_), .B(pi0630), .Y(new_n19310_));
  INVX1    g16874(.A(new_n19310_), .Y(new_n19311_));
  OAI21X1  g16875(.A0(new_n19303_), .A1(pi0647), .B0(pi1157), .Y(new_n19312_));
  AOI21X1  g16876(.A0(new_n19302_), .A1(pi0647), .B0(new_n19312_), .Y(new_n19313_));
  OAI21X1  g16877(.A0(new_n19233_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n19314_));
  AOI21X1  g16878(.A0(new_n19307_), .A1(new_n12577_), .B0(new_n19314_), .Y(new_n19315_));
  NOR2X1   g16879(.A(new_n19315_), .B(new_n12592_), .Y(new_n19316_));
  INVX1    g16880(.A(new_n19316_), .Y(new_n19317_));
  OAI22X1  g16881(.A0(new_n19317_), .A1(new_n19313_), .B0(new_n19311_), .B1(new_n19305_), .Y(new_n19318_));
  MX2X1    g16882(.A(new_n19318_), .B(new_n19302_), .S0(new_n11763_), .Y(new_n19319_));
  OAI21X1  g16883(.A0(new_n19315_), .A1(new_n19309_), .B0(pi0787), .Y(new_n19320_));
  OAI21X1  g16884(.A0(new_n19307_), .A1(pi0787), .B0(new_n19320_), .Y(new_n19321_));
  OAI21X1  g16885(.A0(new_n19321_), .A1(pi0644), .B0(pi0715), .Y(new_n19322_));
  AOI21X1  g16886(.A0(new_n19319_), .A1(pi0644), .B0(new_n19322_), .Y(new_n19323_));
  NOR2X1   g16887(.A(new_n19212_), .B(new_n12605_), .Y(new_n19324_));
  AOI21X1  g16888(.A0(new_n19303_), .A1(new_n12605_), .B0(new_n19324_), .Y(new_n19325_));
  OAI21X1  g16889(.A0(new_n19233_), .A1(pi0644), .B0(new_n12608_), .Y(new_n19326_));
  AOI21X1  g16890(.A0(new_n19325_), .A1(pi0644), .B0(new_n19326_), .Y(new_n19327_));
  NOR3X1   g16891(.A(new_n19327_), .B(new_n19323_), .C(new_n11762_), .Y(new_n19328_));
  OAI21X1  g16892(.A0(new_n19321_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n19329_));
  AOI21X1  g16893(.A0(new_n19319_), .A1(new_n12612_), .B0(new_n19329_), .Y(new_n19330_));
  OAI21X1  g16894(.A0(new_n19233_), .A1(new_n12612_), .B0(pi0715), .Y(new_n19331_));
  AOI21X1  g16895(.A0(new_n19325_), .A1(new_n12612_), .B0(new_n19331_), .Y(new_n19332_));
  OR2X1    g16896(.A(new_n19332_), .B(pi1160), .Y(new_n19333_));
  OAI21X1  g16897(.A0(new_n19333_), .A1(new_n19330_), .B0(pi0790), .Y(new_n19334_));
  OR2X1    g16898(.A(new_n19319_), .B(pi0790), .Y(new_n19335_));
  AND2X1   g16899(.A(new_n19335_), .B(new_n6489_), .Y(new_n19336_));
  OAI21X1  g16900(.A0(new_n19334_), .A1(new_n19328_), .B0(new_n19336_), .Y(new_n19337_));
  AOI21X1  g16901(.A0(po1038), .A1(new_n6818_), .B0(pi0832), .Y(new_n19338_));
  AOI21X1  g16902(.A0(pi1093), .A1(pi1092), .B0(pi0186), .Y(new_n19339_));
  INVX1    g16903(.A(new_n19339_), .Y(new_n19340_));
  AOI21X1  g16904(.A0(new_n12056_), .A1(new_n15235_), .B0(new_n19339_), .Y(new_n19341_));
  AOI21X1  g16905(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n19341_), .Y(new_n19342_));
  INVX1    g16906(.A(new_n19341_), .Y(new_n19343_));
  AOI21X1  g16907(.A0(new_n19343_), .A1(new_n14331_), .B0(new_n12463_), .Y(new_n19344_));
  AOI21X1  g16908(.A0(new_n19342_), .A1(new_n12646_), .B0(pi1155), .Y(new_n19345_));
  OAI21X1  g16909(.A0(new_n19345_), .A1(new_n19344_), .B0(pi0785), .Y(new_n19346_));
  OAI21X1  g16910(.A0(new_n19342_), .A1(pi0785), .B0(new_n19346_), .Y(new_n19347_));
  INVX1    g16911(.A(new_n19347_), .Y(new_n19348_));
  AOI21X1  g16912(.A0(new_n19348_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n19349_));
  AOI21X1  g16913(.A0(new_n19348_), .A1(new_n12655_), .B0(pi1154), .Y(new_n19350_));
  NOR2X1   g16914(.A(new_n19350_), .B(new_n19349_), .Y(new_n19351_));
  MX2X1    g16915(.A(new_n19351_), .B(new_n19348_), .S0(new_n11767_), .Y(new_n19352_));
  NOR2X1   g16916(.A(new_n19352_), .B(pi0789), .Y(new_n19353_));
  INVX1    g16917(.A(new_n19352_), .Y(new_n19354_));
  AOI21X1  g16918(.A0(new_n19339_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19355_));
  OAI21X1  g16919(.A0(new_n19354_), .A1(new_n12509_), .B0(new_n19355_), .Y(new_n19356_));
  AOI21X1  g16920(.A0(new_n19339_), .A1(pi0619), .B0(pi1159), .Y(new_n19357_));
  OAI21X1  g16921(.A0(new_n19354_), .A1(pi0619), .B0(new_n19357_), .Y(new_n19358_));
  AOI21X1  g16922(.A0(new_n19358_), .A1(new_n19356_), .B0(new_n11766_), .Y(new_n19359_));
  NOR2X1   g16923(.A(new_n19359_), .B(new_n19353_), .Y(new_n19360_));
  INVX1    g16924(.A(new_n19360_), .Y(new_n19361_));
  MX2X1    g16925(.A(new_n19361_), .B(new_n19340_), .S0(new_n12708_), .Y(new_n19362_));
  MX2X1    g16926(.A(new_n19362_), .B(new_n19340_), .S0(new_n12580_), .Y(new_n19363_));
  AOI21X1  g16927(.A0(new_n12439_), .A1(pi0703), .B0(new_n19339_), .Y(new_n19364_));
  AND3X1   g16928(.A(new_n12439_), .B(pi0703), .C(new_n12363_), .Y(new_n19365_));
  NOR2X1   g16929(.A(new_n19365_), .B(new_n19364_), .Y(new_n19366_));
  NOR2X1   g16930(.A(new_n19339_), .B(pi1153), .Y(new_n19367_));
  INVX1    g16931(.A(new_n19367_), .Y(new_n19368_));
  OAI22X1  g16932(.A0(new_n19368_), .A1(new_n19365_), .B0(new_n19366_), .B1(new_n12364_), .Y(new_n19369_));
  MX2X1    g16933(.A(new_n19369_), .B(new_n19364_), .S0(new_n11769_), .Y(new_n19370_));
  NOR4X1   g16934(.A(new_n19370_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n19371_));
  AND3X1   g16935(.A(new_n19371_), .B(new_n12739_), .C(new_n12718_), .Y(new_n19372_));
  INVX1    g16936(.A(new_n19372_), .Y(new_n19373_));
  AOI21X1  g16937(.A0(new_n19339_), .A1(pi0647), .B0(pi1157), .Y(new_n19374_));
  OAI21X1  g16938(.A0(new_n19373_), .A1(pi0647), .B0(new_n19374_), .Y(new_n19375_));
  MX2X1    g16939(.A(new_n19372_), .B(new_n19339_), .S0(new_n12577_), .Y(new_n19376_));
  OAI22X1  g16940(.A0(new_n19376_), .A1(new_n14242_), .B0(new_n19375_), .B1(new_n12592_), .Y(new_n19377_));
  AOI21X1  g16941(.A0(new_n19363_), .A1(new_n14326_), .B0(new_n19377_), .Y(new_n19378_));
  AOI21X1  g16942(.A0(new_n19340_), .A1(pi0626), .B0(new_n16218_), .Y(new_n19379_));
  OAI21X1  g16943(.A0(new_n19360_), .A1(pi0626), .B0(new_n19379_), .Y(new_n19380_));
  AOI21X1  g16944(.A0(new_n19340_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n19381_));
  OAI21X1  g16945(.A0(new_n19360_), .A1(new_n12542_), .B0(new_n19381_), .Y(new_n19382_));
  NAND2X1  g16946(.A(new_n19371_), .B(new_n12637_), .Y(new_n19383_));
  AND3X1   g16947(.A(new_n19383_), .B(new_n19382_), .C(new_n19380_), .Y(new_n19384_));
  NOR2X1   g16948(.A(new_n19384_), .B(new_n11765_), .Y(new_n19385_));
  INVX1    g16949(.A(new_n19385_), .Y(new_n19386_));
  NOR2X1   g16950(.A(new_n19364_), .B(new_n11991_), .Y(new_n19387_));
  MX2X1    g16951(.A(new_n19343_), .B(new_n12363_), .S0(new_n19387_), .Y(new_n19388_));
  NOR2X1   g16952(.A(new_n19388_), .B(new_n19368_), .Y(new_n19389_));
  OAI21X1  g16953(.A0(new_n19366_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n19390_));
  NOR2X1   g16954(.A(new_n19390_), .B(new_n19389_), .Y(new_n19391_));
  OR3X1    g16955(.A(new_n19364_), .B(new_n11991_), .C(new_n12363_), .Y(new_n19392_));
  AND2X1   g16956(.A(new_n19341_), .B(pi1153), .Y(new_n19393_));
  OAI21X1  g16957(.A0(new_n19368_), .A1(new_n19365_), .B0(pi0608), .Y(new_n19394_));
  AOI21X1  g16958(.A0(new_n19393_), .A1(new_n19392_), .B0(new_n19394_), .Y(new_n19395_));
  OAI21X1  g16959(.A0(new_n19395_), .A1(new_n19391_), .B0(pi0778), .Y(new_n19396_));
  OAI21X1  g16960(.A0(new_n19387_), .A1(new_n19343_), .B0(new_n11769_), .Y(new_n19397_));
  NAND2X1  g16961(.A(new_n19397_), .B(new_n19396_), .Y(new_n19398_));
  INVX1    g16962(.A(new_n19398_), .Y(new_n19399_));
  OAI21X1  g16963(.A0(new_n19370_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n19400_));
  AOI21X1  g16964(.A0(new_n19398_), .A1(new_n12462_), .B0(new_n19400_), .Y(new_n19401_));
  NOR3X1   g16965(.A(new_n19401_), .B(new_n19344_), .C(pi0660), .Y(new_n19402_));
  OAI21X1  g16966(.A0(new_n19370_), .A1(pi0609), .B0(pi1155), .Y(new_n19403_));
  AOI21X1  g16967(.A0(new_n19398_), .A1(pi0609), .B0(new_n19403_), .Y(new_n19404_));
  NOR3X1   g16968(.A(new_n19404_), .B(new_n19345_), .C(new_n12468_), .Y(new_n19405_));
  NOR2X1   g16969(.A(new_n19405_), .B(new_n19402_), .Y(new_n19406_));
  MX2X1    g16970(.A(new_n19406_), .B(new_n19399_), .S0(new_n11768_), .Y(new_n19407_));
  OR3X1    g16971(.A(new_n19370_), .B(new_n12630_), .C(new_n12486_), .Y(new_n19408_));
  AND2X1   g16972(.A(new_n19408_), .B(new_n12487_), .Y(new_n19409_));
  OAI21X1  g16973(.A0(new_n19407_), .A1(pi0618), .B0(new_n19409_), .Y(new_n19410_));
  NOR2X1   g16974(.A(new_n19349_), .B(pi0627), .Y(new_n19411_));
  NOR3X1   g16975(.A(new_n19370_), .B(new_n12630_), .C(pi0618), .Y(new_n19412_));
  NOR2X1   g16976(.A(new_n19412_), .B(new_n12487_), .Y(new_n19413_));
  OAI21X1  g16977(.A0(new_n19407_), .A1(new_n12486_), .B0(new_n19413_), .Y(new_n19414_));
  NOR2X1   g16978(.A(new_n19350_), .B(new_n12494_), .Y(new_n19415_));
  AOI22X1  g16979(.A0(new_n19415_), .A1(new_n19414_), .B0(new_n19411_), .B1(new_n19410_), .Y(new_n19416_));
  MX2X1    g16980(.A(new_n19416_), .B(new_n19407_), .S0(new_n11767_), .Y(new_n19417_));
  OR4X1    g16981(.A(new_n19370_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n19418_));
  AND2X1   g16982(.A(new_n19418_), .B(new_n12510_), .Y(new_n19419_));
  OAI21X1  g16983(.A0(new_n19417_), .A1(pi0619), .B0(new_n19419_), .Y(new_n19420_));
  AND3X1   g16984(.A(new_n19420_), .B(new_n19356_), .C(new_n12517_), .Y(new_n19421_));
  NOR4X1   g16985(.A(new_n19370_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n19422_));
  NOR2X1   g16986(.A(new_n19422_), .B(new_n12510_), .Y(new_n19423_));
  OAI21X1  g16987(.A0(new_n19417_), .A1(new_n12509_), .B0(new_n19423_), .Y(new_n19424_));
  AND2X1   g16988(.A(new_n19358_), .B(pi0648), .Y(new_n19425_));
  AOI21X1  g16989(.A0(new_n19425_), .A1(new_n19424_), .B0(new_n11766_), .Y(new_n19426_));
  INVX1    g16990(.A(new_n19426_), .Y(new_n19427_));
  AOI21X1  g16991(.A0(new_n19417_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n19428_));
  OAI21X1  g16992(.A0(new_n19427_), .A1(new_n19421_), .B0(new_n19428_), .Y(new_n19429_));
  AOI21X1  g16993(.A0(new_n19429_), .A1(new_n19386_), .B0(new_n14125_), .Y(new_n19430_));
  INVX1    g16994(.A(new_n19362_), .Y(new_n19431_));
  AND2X1   g16995(.A(new_n19371_), .B(new_n12718_), .Y(new_n19432_));
  AOI22X1  g16996(.A0(new_n19432_), .A1(new_n14426_), .B0(new_n19431_), .B1(new_n12735_), .Y(new_n19433_));
  AOI22X1  g16997(.A0(new_n19432_), .A1(new_n14428_), .B0(new_n19431_), .B1(new_n12733_), .Y(new_n19434_));
  MX2X1    g16998(.A(new_n19434_), .B(new_n19433_), .S0(new_n12561_), .Y(new_n19435_));
  OAI21X1  g16999(.A0(new_n19435_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n19436_));
  OAI22X1  g17000(.A0(new_n19436_), .A1(new_n19430_), .B0(new_n19378_), .B1(new_n11763_), .Y(new_n19437_));
  INVX1    g17001(.A(new_n19437_), .Y(new_n19438_));
  OAI21X1  g17002(.A0(new_n19376_), .A1(new_n12578_), .B0(new_n19375_), .Y(new_n19439_));
  MX2X1    g17003(.A(new_n19439_), .B(new_n19373_), .S0(new_n11763_), .Y(new_n19440_));
  OAI21X1  g17004(.A0(new_n19440_), .A1(pi0644), .B0(pi0715), .Y(new_n19441_));
  AOI21X1  g17005(.A0(new_n19438_), .A1(pi0644), .B0(new_n19441_), .Y(new_n19442_));
  OR3X1    g17006(.A(new_n19340_), .B(new_n12603_), .C(new_n11763_), .Y(new_n19443_));
  OAI21X1  g17007(.A0(new_n19363_), .A1(new_n12604_), .B0(new_n19443_), .Y(new_n19444_));
  OAI21X1  g17008(.A0(new_n19340_), .A1(pi0644), .B0(new_n12608_), .Y(new_n19445_));
  AOI21X1  g17009(.A0(new_n19444_), .A1(pi0644), .B0(new_n19445_), .Y(new_n19446_));
  OR2X1    g17010(.A(new_n19446_), .B(new_n11762_), .Y(new_n19447_));
  OAI21X1  g17011(.A0(new_n19440_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n19448_));
  AOI21X1  g17012(.A0(new_n19438_), .A1(new_n12612_), .B0(new_n19448_), .Y(new_n19449_));
  OAI21X1  g17013(.A0(new_n19340_), .A1(new_n12612_), .B0(pi0715), .Y(new_n19450_));
  AOI21X1  g17014(.A0(new_n19444_), .A1(new_n12612_), .B0(new_n19450_), .Y(new_n19451_));
  OR2X1    g17015(.A(new_n19451_), .B(pi1160), .Y(new_n19452_));
  OAI22X1  g17016(.A0(new_n19452_), .A1(new_n19449_), .B0(new_n19447_), .B1(new_n19442_), .Y(new_n19453_));
  OAI21X1  g17017(.A0(new_n19437_), .A1(pi0790), .B0(pi0832), .Y(new_n19454_));
  AOI21X1  g17018(.A0(new_n19453_), .A1(pi0790), .B0(new_n19454_), .Y(new_n19455_));
  AOI21X1  g17019(.A0(new_n19338_), .A1(new_n19337_), .B0(new_n19455_), .Y(po0343));
  OR2X1    g17020(.A(new_n3103_), .B(new_n8646_), .Y(new_n19457_));
  MX2X1    g17021(.A(new_n16611_), .B(new_n12832_), .S0(pi0770), .Y(new_n19458_));
  AOI21X1  g17022(.A0(new_n16616_), .A1(new_n8646_), .B0(pi0770), .Y(new_n19459_));
  AOI22X1  g17023(.A0(new_n19459_), .A1(new_n16617_), .B0(new_n19458_), .B1(new_n8646_), .Y(new_n19460_));
  OR3X1    g17024(.A(new_n13544_), .B(new_n8646_), .C(pi0038), .Y(new_n19461_));
  AND3X1   g17025(.A(new_n19461_), .B(new_n16663_), .C(pi0770), .Y(new_n19462_));
  OAI21X1  g17026(.A0(new_n16662_), .A1(pi0187), .B0(new_n19462_), .Y(new_n19463_));
  AOI21X1  g17027(.A0(new_n16670_), .A1(new_n8646_), .B0(pi0770), .Y(new_n19464_));
  OAI21X1  g17028(.A0(new_n16669_), .A1(new_n8646_), .B0(new_n19464_), .Y(new_n19465_));
  AND2X1   g17029(.A(new_n19465_), .B(pi0726), .Y(new_n19466_));
  AOI21X1  g17030(.A0(new_n19466_), .A1(new_n19463_), .B0(new_n11770_), .Y(new_n19467_));
  OAI21X1  g17031(.A0(new_n19460_), .A1(pi0726), .B0(new_n19467_), .Y(new_n19468_));
  AND3X1   g17032(.A(new_n19468_), .B(new_n19457_), .C(new_n12363_), .Y(new_n19469_));
  MX2X1    g17033(.A(new_n19460_), .B(pi0187), .S0(new_n11770_), .Y(new_n19470_));
  OAI21X1  g17034(.A0(new_n19470_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n19471_));
  OAI21X1  g17035(.A0(new_n12826_), .A1(new_n8646_), .B0(new_n2979_), .Y(new_n19472_));
  AOI21X1  g17036(.A0(new_n12825_), .A1(new_n8646_), .B0(new_n19472_), .Y(new_n19473_));
  AOI21X1  g17037(.A0(new_n12771_), .A1(new_n8646_), .B0(new_n12441_), .Y(new_n19474_));
  NOR3X1   g17038(.A(new_n19474_), .B(new_n19473_), .C(new_n14500_), .Y(new_n19475_));
  NOR2X1   g17039(.A(pi0726), .B(pi0187), .Y(new_n19476_));
  INVX1    g17040(.A(new_n19476_), .Y(new_n19477_));
  OAI21X1  g17041(.A0(new_n19477_), .A1(new_n12447_), .B0(new_n3103_), .Y(new_n19478_));
  OAI21X1  g17042(.A0(new_n19478_), .A1(new_n19475_), .B0(new_n19457_), .Y(new_n19479_));
  OR2X1    g17043(.A(new_n19479_), .B(new_n12363_), .Y(new_n19480_));
  AOI21X1  g17044(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0187), .Y(new_n19481_));
  AOI21X1  g17045(.A0(new_n19481_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n19482_));
  AOI21X1  g17046(.A0(new_n19482_), .A1(new_n19480_), .B0(pi0608), .Y(new_n19483_));
  OAI21X1  g17047(.A0(new_n19471_), .A1(new_n19469_), .B0(new_n19483_), .Y(new_n19484_));
  AND3X1   g17048(.A(new_n19468_), .B(new_n19457_), .C(pi0625), .Y(new_n19485_));
  OAI21X1  g17049(.A0(new_n19470_), .A1(pi0625), .B0(pi1153), .Y(new_n19486_));
  OR2X1    g17050(.A(new_n19479_), .B(pi0625), .Y(new_n19487_));
  AOI21X1  g17051(.A0(new_n19481_), .A1(pi0625), .B0(pi1153), .Y(new_n19488_));
  AOI21X1  g17052(.A0(new_n19488_), .A1(new_n19487_), .B0(new_n12368_), .Y(new_n19489_));
  OAI21X1  g17053(.A0(new_n19486_), .A1(new_n19485_), .B0(new_n19489_), .Y(new_n19490_));
  AOI21X1  g17054(.A0(new_n19490_), .A1(new_n19484_), .B0(new_n11769_), .Y(new_n19491_));
  AND3X1   g17055(.A(new_n19468_), .B(new_n19457_), .C(new_n11769_), .Y(new_n19492_));
  NOR2X1   g17056(.A(new_n19492_), .B(new_n19491_), .Y(new_n19493_));
  NAND2X1  g17057(.A(new_n19479_), .B(new_n11769_), .Y(new_n19494_));
  AOI22X1  g17058(.A0(new_n19488_), .A1(new_n19487_), .B0(new_n19482_), .B1(new_n19480_), .Y(new_n19495_));
  OR2X1    g17059(.A(new_n19495_), .B(new_n11769_), .Y(new_n19496_));
  AND2X1   g17060(.A(new_n19496_), .B(new_n19494_), .Y(new_n19497_));
  AOI21X1  g17061(.A0(new_n19497_), .A1(pi0609), .B0(pi1155), .Y(new_n19498_));
  OAI21X1  g17062(.A0(new_n19493_), .A1(pi0609), .B0(new_n19498_), .Y(new_n19499_));
  INVX1    g17063(.A(new_n19481_), .Y(new_n19500_));
  AND2X1   g17064(.A(new_n19470_), .B(new_n12474_), .Y(new_n19501_));
  AOI22X1  g17065(.A0(new_n19501_), .A1(pi0609), .B0(new_n19500_), .B1(new_n12472_), .Y(new_n19502_));
  OR2X1    g17066(.A(new_n19502_), .B(new_n12463_), .Y(new_n19503_));
  AND2X1   g17067(.A(new_n19503_), .B(new_n12468_), .Y(new_n19504_));
  AOI21X1  g17068(.A0(new_n19497_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n19505_));
  OAI21X1  g17069(.A0(new_n19493_), .A1(new_n12462_), .B0(new_n19505_), .Y(new_n19506_));
  AOI22X1  g17070(.A0(new_n19501_), .A1(new_n12462_), .B0(new_n19500_), .B1(new_n12481_), .Y(new_n19507_));
  OR2X1    g17071(.A(new_n19507_), .B(pi1155), .Y(new_n19508_));
  AND2X1   g17072(.A(new_n19508_), .B(pi0660), .Y(new_n19509_));
  AOI22X1  g17073(.A0(new_n19509_), .A1(new_n19506_), .B0(new_n19504_), .B1(new_n19499_), .Y(new_n19510_));
  OAI21X1  g17074(.A0(new_n19492_), .A1(new_n19491_), .B0(new_n11768_), .Y(new_n19511_));
  OAI21X1  g17075(.A0(new_n19510_), .A1(new_n11768_), .B0(new_n19511_), .Y(new_n19512_));
  OR2X1    g17076(.A(new_n19481_), .B(new_n13910_), .Y(new_n19513_));
  OAI21X1  g17077(.A0(new_n19497_), .A1(new_n12490_), .B0(new_n19513_), .Y(new_n19514_));
  OAI21X1  g17078(.A0(new_n19514_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n19515_));
  AOI21X1  g17079(.A0(new_n19512_), .A1(new_n12486_), .B0(new_n19515_), .Y(new_n19516_));
  AOI21X1  g17080(.A0(new_n19500_), .A1(new_n12473_), .B0(new_n19501_), .Y(new_n19517_));
  MX2X1    g17081(.A(new_n19507_), .B(new_n19502_), .S0(pi1155), .Y(new_n19518_));
  MX2X1    g17082(.A(new_n19518_), .B(new_n19517_), .S0(new_n11768_), .Y(new_n19519_));
  OAI21X1  g17083(.A0(new_n19500_), .A1(pi0618), .B0(pi1154), .Y(new_n19520_));
  AOI21X1  g17084(.A0(new_n19519_), .A1(pi0618), .B0(new_n19520_), .Y(new_n19521_));
  OR2X1    g17085(.A(new_n19521_), .B(pi0627), .Y(new_n19522_));
  OAI21X1  g17086(.A0(new_n19514_), .A1(pi0618), .B0(pi1154), .Y(new_n19523_));
  AOI21X1  g17087(.A0(new_n19512_), .A1(pi0618), .B0(new_n19523_), .Y(new_n19524_));
  OAI21X1  g17088(.A0(new_n19500_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n19525_));
  AOI21X1  g17089(.A0(new_n19519_), .A1(new_n12486_), .B0(new_n19525_), .Y(new_n19526_));
  OR2X1    g17090(.A(new_n19526_), .B(new_n12494_), .Y(new_n19527_));
  OAI22X1  g17091(.A0(new_n19527_), .A1(new_n19524_), .B0(new_n19522_), .B1(new_n19516_), .Y(new_n19528_));
  MX2X1    g17092(.A(new_n19528_), .B(new_n19512_), .S0(new_n11767_), .Y(new_n19529_));
  MX2X1    g17093(.A(new_n19514_), .B(new_n19500_), .S0(new_n12513_), .Y(new_n19530_));
  OAI21X1  g17094(.A0(new_n19530_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19531_));
  AOI21X1  g17095(.A0(new_n19529_), .A1(new_n12509_), .B0(new_n19531_), .Y(new_n19532_));
  OR2X1    g17096(.A(new_n19519_), .B(pi0781), .Y(new_n19533_));
  OAI21X1  g17097(.A0(new_n19526_), .A1(new_n19521_), .B0(pi0781), .Y(new_n19534_));
  NAND3X1  g17098(.A(new_n19534_), .B(new_n19533_), .C(pi0619), .Y(new_n19535_));
  AOI21X1  g17099(.A0(new_n19481_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19536_));
  AND2X1   g17100(.A(new_n19536_), .B(new_n19535_), .Y(new_n19537_));
  OR2X1    g17101(.A(new_n19537_), .B(pi0648), .Y(new_n19538_));
  OAI21X1  g17102(.A0(new_n19530_), .A1(pi0619), .B0(pi1159), .Y(new_n19539_));
  AOI21X1  g17103(.A0(new_n19529_), .A1(pi0619), .B0(new_n19539_), .Y(new_n19540_));
  NAND3X1  g17104(.A(new_n19534_), .B(new_n19533_), .C(new_n12509_), .Y(new_n19541_));
  AOI21X1  g17105(.A0(new_n19481_), .A1(pi0619), .B0(pi1159), .Y(new_n19542_));
  AND2X1   g17106(.A(new_n19542_), .B(new_n19541_), .Y(new_n19543_));
  OR2X1    g17107(.A(new_n19543_), .B(new_n12517_), .Y(new_n19544_));
  OAI22X1  g17108(.A0(new_n19544_), .A1(new_n19540_), .B0(new_n19538_), .B1(new_n19532_), .Y(new_n19545_));
  MX2X1    g17109(.A(new_n19545_), .B(new_n19529_), .S0(new_n11766_), .Y(new_n19546_));
  MX2X1    g17110(.A(new_n19530_), .B(new_n19500_), .S0(new_n12531_), .Y(new_n19547_));
  AOI21X1  g17111(.A0(new_n19547_), .A1(pi0626), .B0(pi0641), .Y(new_n19548_));
  OAI21X1  g17112(.A0(new_n19546_), .A1(pi0626), .B0(new_n19548_), .Y(new_n19549_));
  AND2X1   g17113(.A(new_n19534_), .B(new_n19533_), .Y(new_n19550_));
  AOI22X1  g17114(.A0(new_n19542_), .A1(new_n19541_), .B0(new_n19536_), .B1(new_n19535_), .Y(new_n19551_));
  MX2X1    g17115(.A(new_n19551_), .B(new_n19550_), .S0(new_n11766_), .Y(new_n19552_));
  AOI21X1  g17116(.A0(new_n19500_), .A1(pi0626), .B0(new_n12543_), .Y(new_n19553_));
  OAI21X1  g17117(.A0(new_n19552_), .A1(pi0626), .B0(new_n19553_), .Y(new_n19554_));
  AND2X1   g17118(.A(new_n19554_), .B(new_n12548_), .Y(new_n19555_));
  AOI21X1  g17119(.A0(new_n19547_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n19556_));
  OAI21X1  g17120(.A0(new_n19546_), .A1(new_n12542_), .B0(new_n19556_), .Y(new_n19557_));
  AOI21X1  g17121(.A0(new_n19500_), .A1(new_n12542_), .B0(pi0641), .Y(new_n19558_));
  OAI21X1  g17122(.A0(new_n19552_), .A1(new_n12542_), .B0(new_n19558_), .Y(new_n19559_));
  AND2X1   g17123(.A(new_n19559_), .B(pi1158), .Y(new_n19560_));
  AOI22X1  g17124(.A0(new_n19560_), .A1(new_n19557_), .B0(new_n19555_), .B1(new_n19549_), .Y(new_n19561_));
  MX2X1    g17125(.A(new_n19561_), .B(new_n19546_), .S0(new_n11765_), .Y(new_n19562_));
  MX2X1    g17126(.A(new_n19552_), .B(new_n19481_), .S0(new_n12708_), .Y(new_n19563_));
  INVX1    g17127(.A(new_n19563_), .Y(new_n19564_));
  OAI21X1  g17128(.A0(new_n19564_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n19565_));
  AOI21X1  g17129(.A0(new_n19562_), .A1(new_n12554_), .B0(new_n19565_), .Y(new_n19566_));
  MX2X1    g17130(.A(new_n19547_), .B(new_n19500_), .S0(new_n12563_), .Y(new_n19567_));
  AOI21X1  g17131(.A0(new_n19481_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n19568_));
  OAI21X1  g17132(.A0(new_n19567_), .A1(new_n12554_), .B0(new_n19568_), .Y(new_n19569_));
  NAND2X1  g17133(.A(new_n19569_), .B(new_n12561_), .Y(new_n19570_));
  OAI21X1  g17134(.A0(new_n19564_), .A1(pi0628), .B0(pi1156), .Y(new_n19571_));
  AOI21X1  g17135(.A0(new_n19562_), .A1(pi0628), .B0(new_n19571_), .Y(new_n19572_));
  AOI21X1  g17136(.A0(new_n19481_), .A1(pi0628), .B0(pi1156), .Y(new_n19573_));
  OAI21X1  g17137(.A0(new_n19567_), .A1(pi0628), .B0(new_n19573_), .Y(new_n19574_));
  NAND2X1  g17138(.A(new_n19574_), .B(pi0629), .Y(new_n19575_));
  OAI22X1  g17139(.A0(new_n19575_), .A1(new_n19572_), .B0(new_n19570_), .B1(new_n19566_), .Y(new_n19576_));
  AND2X1   g17140(.A(new_n19562_), .B(new_n11764_), .Y(new_n19577_));
  AOI21X1  g17141(.A0(new_n19576_), .A1(pi0792), .B0(new_n19577_), .Y(new_n19578_));
  MX2X1    g17142(.A(new_n19564_), .B(new_n19500_), .S0(new_n12580_), .Y(new_n19579_));
  INVX1    g17143(.A(new_n19579_), .Y(new_n19580_));
  AOI21X1  g17144(.A0(new_n19580_), .A1(pi0647), .B0(pi1157), .Y(new_n19581_));
  OAI21X1  g17145(.A0(new_n19578_), .A1(pi0647), .B0(new_n19581_), .Y(new_n19582_));
  INVX1    g17146(.A(new_n19567_), .Y(new_n19583_));
  AND2X1   g17147(.A(new_n19574_), .B(new_n19569_), .Y(new_n19584_));
  MX2X1    g17148(.A(new_n19584_), .B(new_n19583_), .S0(new_n11764_), .Y(new_n19585_));
  INVX1    g17149(.A(new_n19585_), .Y(new_n19586_));
  AOI21X1  g17150(.A0(new_n19481_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n19587_));
  OAI21X1  g17151(.A0(new_n19586_), .A1(new_n12577_), .B0(new_n19587_), .Y(new_n19588_));
  AND2X1   g17152(.A(new_n19588_), .B(new_n12592_), .Y(new_n19589_));
  AOI21X1  g17153(.A0(new_n19580_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n19590_));
  OAI21X1  g17154(.A0(new_n19578_), .A1(new_n12577_), .B0(new_n19590_), .Y(new_n19591_));
  AOI21X1  g17155(.A0(new_n19481_), .A1(pi0647), .B0(pi1157), .Y(new_n19592_));
  OAI21X1  g17156(.A0(new_n19586_), .A1(pi0647), .B0(new_n19592_), .Y(new_n19593_));
  AND2X1   g17157(.A(new_n19593_), .B(pi0630), .Y(new_n19594_));
  AOI22X1  g17158(.A0(new_n19594_), .A1(new_n19591_), .B0(new_n19589_), .B1(new_n19582_), .Y(new_n19595_));
  MX2X1    g17159(.A(new_n19595_), .B(new_n19578_), .S0(new_n11763_), .Y(new_n19596_));
  AND2X1   g17160(.A(new_n19593_), .B(new_n19588_), .Y(new_n19597_));
  MX2X1    g17161(.A(new_n19597_), .B(new_n19585_), .S0(new_n11763_), .Y(new_n19598_));
  AOI21X1  g17162(.A0(new_n19598_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n19599_));
  OAI21X1  g17163(.A0(new_n19596_), .A1(new_n12612_), .B0(new_n19599_), .Y(new_n19600_));
  MX2X1    g17164(.A(new_n19580_), .B(new_n19481_), .S0(new_n12604_), .Y(new_n19601_));
  OAI21X1  g17165(.A0(new_n19500_), .A1(pi0644), .B0(new_n12608_), .Y(new_n19602_));
  AOI21X1  g17166(.A0(new_n19601_), .A1(pi0644), .B0(new_n19602_), .Y(new_n19603_));
  NOR2X1   g17167(.A(new_n19603_), .B(new_n11762_), .Y(new_n19604_));
  AND2X1   g17168(.A(new_n19604_), .B(new_n19600_), .Y(new_n19605_));
  OR2X1    g17169(.A(new_n19578_), .B(pi0787), .Y(new_n19606_));
  OAI21X1  g17170(.A0(new_n19595_), .A1(new_n11763_), .B0(new_n19606_), .Y(new_n19607_));
  AND2X1   g17171(.A(new_n19598_), .B(pi0644), .Y(new_n19608_));
  OR2X1    g17172(.A(new_n19608_), .B(pi0715), .Y(new_n19609_));
  AOI21X1  g17173(.A0(new_n19607_), .A1(new_n12612_), .B0(new_n19609_), .Y(new_n19610_));
  OAI21X1  g17174(.A0(new_n19500_), .A1(new_n12612_), .B0(pi0715), .Y(new_n19611_));
  AOI21X1  g17175(.A0(new_n19601_), .A1(new_n12612_), .B0(new_n19611_), .Y(new_n19612_));
  OR2X1    g17176(.A(new_n19612_), .B(pi1160), .Y(new_n19613_));
  OAI21X1  g17177(.A0(new_n19613_), .A1(new_n19610_), .B0(pi0790), .Y(new_n19614_));
  AOI21X1  g17178(.A0(new_n19596_), .A1(new_n12766_), .B0(po1038), .Y(new_n19615_));
  OAI21X1  g17179(.A0(new_n19614_), .A1(new_n19605_), .B0(new_n19615_), .Y(new_n19616_));
  AOI21X1  g17180(.A0(po1038), .A1(new_n8646_), .B0(pi0832), .Y(new_n19617_));
  AOI21X1  g17181(.A0(pi1093), .A1(pi1092), .B0(pi0187), .Y(new_n19618_));
  INVX1    g17182(.A(new_n19618_), .Y(new_n19619_));
  AOI21X1  g17183(.A0(new_n12056_), .A1(new_n14522_), .B0(new_n19618_), .Y(new_n19620_));
  AOI21X1  g17184(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n19620_), .Y(new_n19621_));
  INVX1    g17185(.A(new_n19620_), .Y(new_n19622_));
  AOI21X1  g17186(.A0(new_n19622_), .A1(new_n14331_), .B0(new_n12463_), .Y(new_n19623_));
  AOI21X1  g17187(.A0(new_n19621_), .A1(new_n12646_), .B0(pi1155), .Y(new_n19624_));
  OAI21X1  g17188(.A0(new_n19624_), .A1(new_n19623_), .B0(pi0785), .Y(new_n19625_));
  OAI21X1  g17189(.A0(new_n19621_), .A1(pi0785), .B0(new_n19625_), .Y(new_n19626_));
  INVX1    g17190(.A(new_n19626_), .Y(new_n19627_));
  AOI21X1  g17191(.A0(new_n19627_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n19628_));
  AOI21X1  g17192(.A0(new_n19627_), .A1(new_n12655_), .B0(pi1154), .Y(new_n19629_));
  NOR2X1   g17193(.A(new_n19629_), .B(new_n19628_), .Y(new_n19630_));
  MX2X1    g17194(.A(new_n19630_), .B(new_n19627_), .S0(new_n11767_), .Y(new_n19631_));
  NOR2X1   g17195(.A(new_n19631_), .B(pi0789), .Y(new_n19632_));
  INVX1    g17196(.A(new_n19631_), .Y(new_n19633_));
  AOI21X1  g17197(.A0(new_n19618_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19634_));
  OAI21X1  g17198(.A0(new_n19633_), .A1(new_n12509_), .B0(new_n19634_), .Y(new_n19635_));
  AOI21X1  g17199(.A0(new_n19618_), .A1(pi0619), .B0(pi1159), .Y(new_n19636_));
  OAI21X1  g17200(.A0(new_n19633_), .A1(pi0619), .B0(new_n19636_), .Y(new_n19637_));
  AOI21X1  g17201(.A0(new_n19637_), .A1(new_n19635_), .B0(new_n11766_), .Y(new_n19638_));
  NOR2X1   g17202(.A(new_n19638_), .B(new_n19632_), .Y(new_n19639_));
  INVX1    g17203(.A(new_n19639_), .Y(new_n19640_));
  MX2X1    g17204(.A(new_n19640_), .B(new_n19619_), .S0(new_n12708_), .Y(new_n19641_));
  MX2X1    g17205(.A(new_n19641_), .B(new_n19619_), .S0(new_n12580_), .Y(new_n19642_));
  AOI21X1  g17206(.A0(new_n12439_), .A1(pi0726), .B0(new_n19618_), .Y(new_n19643_));
  AND3X1   g17207(.A(new_n12439_), .B(pi0726), .C(new_n12363_), .Y(new_n19644_));
  NOR2X1   g17208(.A(new_n19644_), .B(new_n19643_), .Y(new_n19645_));
  NOR2X1   g17209(.A(new_n19618_), .B(pi1153), .Y(new_n19646_));
  INVX1    g17210(.A(new_n19646_), .Y(new_n19647_));
  OAI22X1  g17211(.A0(new_n19647_), .A1(new_n19644_), .B0(new_n19645_), .B1(new_n12364_), .Y(new_n19648_));
  MX2X1    g17212(.A(new_n19648_), .B(new_n19643_), .S0(new_n11769_), .Y(new_n19649_));
  NOR4X1   g17213(.A(new_n19649_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n19650_));
  AND3X1   g17214(.A(new_n19650_), .B(new_n12739_), .C(new_n12718_), .Y(new_n19651_));
  INVX1    g17215(.A(new_n19651_), .Y(new_n19652_));
  AOI21X1  g17216(.A0(new_n19618_), .A1(pi0647), .B0(pi1157), .Y(new_n19653_));
  OAI21X1  g17217(.A0(new_n19652_), .A1(pi0647), .B0(new_n19653_), .Y(new_n19654_));
  MX2X1    g17218(.A(new_n19651_), .B(new_n19618_), .S0(new_n12577_), .Y(new_n19655_));
  OAI22X1  g17219(.A0(new_n19655_), .A1(new_n14242_), .B0(new_n19654_), .B1(new_n12592_), .Y(new_n19656_));
  AOI21X1  g17220(.A0(new_n19642_), .A1(new_n14326_), .B0(new_n19656_), .Y(new_n19657_));
  AOI21X1  g17221(.A0(new_n19619_), .A1(pi0626), .B0(new_n16218_), .Y(new_n19658_));
  OAI21X1  g17222(.A0(new_n19639_), .A1(pi0626), .B0(new_n19658_), .Y(new_n19659_));
  AOI21X1  g17223(.A0(new_n19619_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n19660_));
  OAI21X1  g17224(.A0(new_n19639_), .A1(new_n12542_), .B0(new_n19660_), .Y(new_n19661_));
  NAND2X1  g17225(.A(new_n19650_), .B(new_n12637_), .Y(new_n19662_));
  AND3X1   g17226(.A(new_n19662_), .B(new_n19661_), .C(new_n19659_), .Y(new_n19663_));
  NOR2X1   g17227(.A(new_n19663_), .B(new_n11765_), .Y(new_n19664_));
  INVX1    g17228(.A(new_n19664_), .Y(new_n19665_));
  NOR2X1   g17229(.A(new_n19643_), .B(new_n11991_), .Y(new_n19666_));
  MX2X1    g17230(.A(new_n19622_), .B(new_n12363_), .S0(new_n19666_), .Y(new_n19667_));
  NOR2X1   g17231(.A(new_n19667_), .B(new_n19647_), .Y(new_n19668_));
  OAI21X1  g17232(.A0(new_n19645_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n19669_));
  NOR2X1   g17233(.A(new_n19669_), .B(new_n19668_), .Y(new_n19670_));
  OR3X1    g17234(.A(new_n19643_), .B(new_n11991_), .C(new_n12363_), .Y(new_n19671_));
  AND2X1   g17235(.A(new_n19620_), .B(pi1153), .Y(new_n19672_));
  OAI21X1  g17236(.A0(new_n19647_), .A1(new_n19644_), .B0(pi0608), .Y(new_n19673_));
  AOI21X1  g17237(.A0(new_n19672_), .A1(new_n19671_), .B0(new_n19673_), .Y(new_n19674_));
  OAI21X1  g17238(.A0(new_n19674_), .A1(new_n19670_), .B0(pi0778), .Y(new_n19675_));
  OAI21X1  g17239(.A0(new_n19666_), .A1(new_n19622_), .B0(new_n11769_), .Y(new_n19676_));
  NAND2X1  g17240(.A(new_n19676_), .B(new_n19675_), .Y(new_n19677_));
  INVX1    g17241(.A(new_n19677_), .Y(new_n19678_));
  OAI21X1  g17242(.A0(new_n19649_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n19679_));
  AOI21X1  g17243(.A0(new_n19677_), .A1(new_n12462_), .B0(new_n19679_), .Y(new_n19680_));
  NOR3X1   g17244(.A(new_n19680_), .B(new_n19623_), .C(pi0660), .Y(new_n19681_));
  OAI21X1  g17245(.A0(new_n19649_), .A1(pi0609), .B0(pi1155), .Y(new_n19682_));
  AOI21X1  g17246(.A0(new_n19677_), .A1(pi0609), .B0(new_n19682_), .Y(new_n19683_));
  NOR3X1   g17247(.A(new_n19683_), .B(new_n19624_), .C(new_n12468_), .Y(new_n19684_));
  NOR2X1   g17248(.A(new_n19684_), .B(new_n19681_), .Y(new_n19685_));
  MX2X1    g17249(.A(new_n19685_), .B(new_n19678_), .S0(new_n11768_), .Y(new_n19686_));
  OR3X1    g17250(.A(new_n19649_), .B(new_n12630_), .C(new_n12486_), .Y(new_n19687_));
  AND2X1   g17251(.A(new_n19687_), .B(new_n12487_), .Y(new_n19688_));
  OAI21X1  g17252(.A0(new_n19686_), .A1(pi0618), .B0(new_n19688_), .Y(new_n19689_));
  NOR2X1   g17253(.A(new_n19628_), .B(pi0627), .Y(new_n19690_));
  NOR3X1   g17254(.A(new_n19649_), .B(new_n12630_), .C(pi0618), .Y(new_n19691_));
  NOR2X1   g17255(.A(new_n19691_), .B(new_n12487_), .Y(new_n19692_));
  OAI21X1  g17256(.A0(new_n19686_), .A1(new_n12486_), .B0(new_n19692_), .Y(new_n19693_));
  NOR2X1   g17257(.A(new_n19629_), .B(new_n12494_), .Y(new_n19694_));
  AOI22X1  g17258(.A0(new_n19694_), .A1(new_n19693_), .B0(new_n19690_), .B1(new_n19689_), .Y(new_n19695_));
  MX2X1    g17259(.A(new_n19695_), .B(new_n19686_), .S0(new_n11767_), .Y(new_n19696_));
  OR4X1    g17260(.A(new_n19649_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n19697_));
  AND2X1   g17261(.A(new_n19697_), .B(new_n12510_), .Y(new_n19698_));
  OAI21X1  g17262(.A0(new_n19696_), .A1(pi0619), .B0(new_n19698_), .Y(new_n19699_));
  AND3X1   g17263(.A(new_n19699_), .B(new_n19635_), .C(new_n12517_), .Y(new_n19700_));
  NOR4X1   g17264(.A(new_n19649_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n19701_));
  NOR2X1   g17265(.A(new_n19701_), .B(new_n12510_), .Y(new_n19702_));
  OAI21X1  g17266(.A0(new_n19696_), .A1(new_n12509_), .B0(new_n19702_), .Y(new_n19703_));
  AND2X1   g17267(.A(new_n19637_), .B(pi0648), .Y(new_n19704_));
  AOI21X1  g17268(.A0(new_n19704_), .A1(new_n19703_), .B0(new_n11766_), .Y(new_n19705_));
  INVX1    g17269(.A(new_n19705_), .Y(new_n19706_));
  AOI21X1  g17270(.A0(new_n19696_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n19707_));
  OAI21X1  g17271(.A0(new_n19706_), .A1(new_n19700_), .B0(new_n19707_), .Y(new_n19708_));
  AOI21X1  g17272(.A0(new_n19708_), .A1(new_n19665_), .B0(new_n14125_), .Y(new_n19709_));
  INVX1    g17273(.A(new_n19641_), .Y(new_n19710_));
  AND2X1   g17274(.A(new_n19650_), .B(new_n12718_), .Y(new_n19711_));
  AOI22X1  g17275(.A0(new_n19711_), .A1(new_n14426_), .B0(new_n19710_), .B1(new_n12735_), .Y(new_n19712_));
  AOI22X1  g17276(.A0(new_n19711_), .A1(new_n14428_), .B0(new_n19710_), .B1(new_n12733_), .Y(new_n19713_));
  MX2X1    g17277(.A(new_n19713_), .B(new_n19712_), .S0(new_n12561_), .Y(new_n19714_));
  OAI21X1  g17278(.A0(new_n19714_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n19715_));
  OAI22X1  g17279(.A0(new_n19715_), .A1(new_n19709_), .B0(new_n19657_), .B1(new_n11763_), .Y(new_n19716_));
  INVX1    g17280(.A(new_n19716_), .Y(new_n19717_));
  OAI21X1  g17281(.A0(new_n19655_), .A1(new_n12578_), .B0(new_n19654_), .Y(new_n19718_));
  MX2X1    g17282(.A(new_n19718_), .B(new_n19652_), .S0(new_n11763_), .Y(new_n19719_));
  OAI21X1  g17283(.A0(new_n19719_), .A1(pi0644), .B0(pi0715), .Y(new_n19720_));
  AOI21X1  g17284(.A0(new_n19717_), .A1(pi0644), .B0(new_n19720_), .Y(new_n19721_));
  OR3X1    g17285(.A(new_n19619_), .B(new_n12603_), .C(new_n11763_), .Y(new_n19722_));
  OAI21X1  g17286(.A0(new_n19642_), .A1(new_n12604_), .B0(new_n19722_), .Y(new_n19723_));
  OAI21X1  g17287(.A0(new_n19619_), .A1(pi0644), .B0(new_n12608_), .Y(new_n19724_));
  AOI21X1  g17288(.A0(new_n19723_), .A1(pi0644), .B0(new_n19724_), .Y(new_n19725_));
  OR2X1    g17289(.A(new_n19725_), .B(new_n11762_), .Y(new_n19726_));
  OAI21X1  g17290(.A0(new_n19719_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n19727_));
  AOI21X1  g17291(.A0(new_n19717_), .A1(new_n12612_), .B0(new_n19727_), .Y(new_n19728_));
  OAI21X1  g17292(.A0(new_n19619_), .A1(new_n12612_), .B0(pi0715), .Y(new_n19729_));
  AOI21X1  g17293(.A0(new_n19723_), .A1(new_n12612_), .B0(new_n19729_), .Y(new_n19730_));
  OR2X1    g17294(.A(new_n19730_), .B(pi1160), .Y(new_n19731_));
  OAI22X1  g17295(.A0(new_n19731_), .A1(new_n19728_), .B0(new_n19726_), .B1(new_n19721_), .Y(new_n19732_));
  OAI21X1  g17296(.A0(new_n19716_), .A1(pi0790), .B0(pi0832), .Y(new_n19733_));
  AOI21X1  g17297(.A0(new_n19732_), .A1(pi0790), .B0(new_n19733_), .Y(new_n19734_));
  AOI21X1  g17298(.A0(new_n19617_), .A1(new_n19616_), .B0(new_n19734_), .Y(po0344));
  OR2X1    g17299(.A(new_n3103_), .B(new_n7436_), .Y(new_n19736_));
  MX2X1    g17300(.A(new_n16611_), .B(new_n12832_), .S0(pi0768), .Y(new_n19737_));
  AOI21X1  g17301(.A0(new_n16616_), .A1(new_n7436_), .B0(pi0768), .Y(new_n19738_));
  AOI22X1  g17302(.A0(new_n19738_), .A1(new_n16617_), .B0(new_n19737_), .B1(new_n7436_), .Y(new_n19739_));
  OR3X1    g17303(.A(new_n13544_), .B(new_n7436_), .C(pi0038), .Y(new_n19740_));
  AND3X1   g17304(.A(new_n19740_), .B(new_n16663_), .C(pi0768), .Y(new_n19741_));
  OAI21X1  g17305(.A0(new_n16662_), .A1(pi0188), .B0(new_n19741_), .Y(new_n19742_));
  AOI21X1  g17306(.A0(new_n16670_), .A1(new_n7436_), .B0(pi0768), .Y(new_n19743_));
  OAI21X1  g17307(.A0(new_n16669_), .A1(new_n7436_), .B0(new_n19743_), .Y(new_n19744_));
  AND2X1   g17308(.A(new_n19744_), .B(pi0705), .Y(new_n19745_));
  AOI21X1  g17309(.A0(new_n19745_), .A1(new_n19742_), .B0(new_n11770_), .Y(new_n19746_));
  OAI21X1  g17310(.A0(new_n19739_), .A1(pi0705), .B0(new_n19746_), .Y(new_n19747_));
  AND3X1   g17311(.A(new_n19747_), .B(new_n19736_), .C(new_n12363_), .Y(new_n19748_));
  MX2X1    g17312(.A(new_n19739_), .B(pi0188), .S0(new_n11770_), .Y(new_n19749_));
  OAI21X1  g17313(.A0(new_n19749_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n19750_));
  OAI21X1  g17314(.A0(new_n12826_), .A1(new_n7436_), .B0(new_n2979_), .Y(new_n19751_));
  AOI21X1  g17315(.A0(new_n12825_), .A1(new_n7436_), .B0(new_n19751_), .Y(new_n19752_));
  AOI21X1  g17316(.A0(new_n12771_), .A1(new_n7436_), .B0(new_n12441_), .Y(new_n19753_));
  NOR3X1   g17317(.A(new_n19753_), .B(new_n19752_), .C(new_n15335_), .Y(new_n19754_));
  NOR2X1   g17318(.A(pi0705), .B(pi0188), .Y(new_n19755_));
  INVX1    g17319(.A(new_n19755_), .Y(new_n19756_));
  OAI21X1  g17320(.A0(new_n19756_), .A1(new_n12447_), .B0(new_n3103_), .Y(new_n19757_));
  OAI21X1  g17321(.A0(new_n19757_), .A1(new_n19754_), .B0(new_n19736_), .Y(new_n19758_));
  OR2X1    g17322(.A(new_n19758_), .B(new_n12363_), .Y(new_n19759_));
  AOI21X1  g17323(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0188), .Y(new_n19760_));
  AOI21X1  g17324(.A0(new_n19760_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n19761_));
  AOI21X1  g17325(.A0(new_n19761_), .A1(new_n19759_), .B0(pi0608), .Y(new_n19762_));
  OAI21X1  g17326(.A0(new_n19750_), .A1(new_n19748_), .B0(new_n19762_), .Y(new_n19763_));
  AND3X1   g17327(.A(new_n19747_), .B(new_n19736_), .C(pi0625), .Y(new_n19764_));
  OAI21X1  g17328(.A0(new_n19749_), .A1(pi0625), .B0(pi1153), .Y(new_n19765_));
  OR2X1    g17329(.A(new_n19758_), .B(pi0625), .Y(new_n19766_));
  AOI21X1  g17330(.A0(new_n19760_), .A1(pi0625), .B0(pi1153), .Y(new_n19767_));
  AOI21X1  g17331(.A0(new_n19767_), .A1(new_n19766_), .B0(new_n12368_), .Y(new_n19768_));
  OAI21X1  g17332(.A0(new_n19765_), .A1(new_n19764_), .B0(new_n19768_), .Y(new_n19769_));
  AOI21X1  g17333(.A0(new_n19769_), .A1(new_n19763_), .B0(new_n11769_), .Y(new_n19770_));
  AND3X1   g17334(.A(new_n19747_), .B(new_n19736_), .C(new_n11769_), .Y(new_n19771_));
  NOR2X1   g17335(.A(new_n19771_), .B(new_n19770_), .Y(new_n19772_));
  NAND2X1  g17336(.A(new_n19758_), .B(new_n11769_), .Y(new_n19773_));
  AOI22X1  g17337(.A0(new_n19767_), .A1(new_n19766_), .B0(new_n19761_), .B1(new_n19759_), .Y(new_n19774_));
  OR2X1    g17338(.A(new_n19774_), .B(new_n11769_), .Y(new_n19775_));
  AND2X1   g17339(.A(new_n19775_), .B(new_n19773_), .Y(new_n19776_));
  AOI21X1  g17340(.A0(new_n19776_), .A1(pi0609), .B0(pi1155), .Y(new_n19777_));
  OAI21X1  g17341(.A0(new_n19772_), .A1(pi0609), .B0(new_n19777_), .Y(new_n19778_));
  INVX1    g17342(.A(new_n19760_), .Y(new_n19779_));
  AND2X1   g17343(.A(new_n19749_), .B(new_n12474_), .Y(new_n19780_));
  AOI22X1  g17344(.A0(new_n19780_), .A1(pi0609), .B0(new_n19779_), .B1(new_n12472_), .Y(new_n19781_));
  OR2X1    g17345(.A(new_n19781_), .B(new_n12463_), .Y(new_n19782_));
  AND2X1   g17346(.A(new_n19782_), .B(new_n12468_), .Y(new_n19783_));
  AOI21X1  g17347(.A0(new_n19776_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n19784_));
  OAI21X1  g17348(.A0(new_n19772_), .A1(new_n12462_), .B0(new_n19784_), .Y(new_n19785_));
  AOI22X1  g17349(.A0(new_n19780_), .A1(new_n12462_), .B0(new_n19779_), .B1(new_n12481_), .Y(new_n19786_));
  OR2X1    g17350(.A(new_n19786_), .B(pi1155), .Y(new_n19787_));
  AND2X1   g17351(.A(new_n19787_), .B(pi0660), .Y(new_n19788_));
  AOI22X1  g17352(.A0(new_n19788_), .A1(new_n19785_), .B0(new_n19783_), .B1(new_n19778_), .Y(new_n19789_));
  OAI21X1  g17353(.A0(new_n19771_), .A1(new_n19770_), .B0(new_n11768_), .Y(new_n19790_));
  OAI21X1  g17354(.A0(new_n19789_), .A1(new_n11768_), .B0(new_n19790_), .Y(new_n19791_));
  OR2X1    g17355(.A(new_n19760_), .B(new_n13910_), .Y(new_n19792_));
  OAI21X1  g17356(.A0(new_n19776_), .A1(new_n12490_), .B0(new_n19792_), .Y(new_n19793_));
  OAI21X1  g17357(.A0(new_n19793_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n19794_));
  AOI21X1  g17358(.A0(new_n19791_), .A1(new_n12486_), .B0(new_n19794_), .Y(new_n19795_));
  AOI21X1  g17359(.A0(new_n19779_), .A1(new_n12473_), .B0(new_n19780_), .Y(new_n19796_));
  MX2X1    g17360(.A(new_n19786_), .B(new_n19781_), .S0(pi1155), .Y(new_n19797_));
  MX2X1    g17361(.A(new_n19797_), .B(new_n19796_), .S0(new_n11768_), .Y(new_n19798_));
  OAI21X1  g17362(.A0(new_n19779_), .A1(pi0618), .B0(pi1154), .Y(new_n19799_));
  AOI21X1  g17363(.A0(new_n19798_), .A1(pi0618), .B0(new_n19799_), .Y(new_n19800_));
  OR2X1    g17364(.A(new_n19800_), .B(pi0627), .Y(new_n19801_));
  OAI21X1  g17365(.A0(new_n19793_), .A1(pi0618), .B0(pi1154), .Y(new_n19802_));
  AOI21X1  g17366(.A0(new_n19791_), .A1(pi0618), .B0(new_n19802_), .Y(new_n19803_));
  OAI21X1  g17367(.A0(new_n19779_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n19804_));
  AOI21X1  g17368(.A0(new_n19798_), .A1(new_n12486_), .B0(new_n19804_), .Y(new_n19805_));
  OR2X1    g17369(.A(new_n19805_), .B(new_n12494_), .Y(new_n19806_));
  OAI22X1  g17370(.A0(new_n19806_), .A1(new_n19803_), .B0(new_n19801_), .B1(new_n19795_), .Y(new_n19807_));
  MX2X1    g17371(.A(new_n19807_), .B(new_n19791_), .S0(new_n11767_), .Y(new_n19808_));
  MX2X1    g17372(.A(new_n19793_), .B(new_n19779_), .S0(new_n12513_), .Y(new_n19809_));
  OAI21X1  g17373(.A0(new_n19809_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19810_));
  AOI21X1  g17374(.A0(new_n19808_), .A1(new_n12509_), .B0(new_n19810_), .Y(new_n19811_));
  OR2X1    g17375(.A(new_n19798_), .B(pi0781), .Y(new_n19812_));
  OAI21X1  g17376(.A0(new_n19805_), .A1(new_n19800_), .B0(pi0781), .Y(new_n19813_));
  NAND3X1  g17377(.A(new_n19813_), .B(new_n19812_), .C(pi0619), .Y(new_n19814_));
  AOI21X1  g17378(.A0(new_n19760_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19815_));
  AND2X1   g17379(.A(new_n19815_), .B(new_n19814_), .Y(new_n19816_));
  OR2X1    g17380(.A(new_n19816_), .B(pi0648), .Y(new_n19817_));
  OAI21X1  g17381(.A0(new_n19809_), .A1(pi0619), .B0(pi1159), .Y(new_n19818_));
  AOI21X1  g17382(.A0(new_n19808_), .A1(pi0619), .B0(new_n19818_), .Y(new_n19819_));
  NAND3X1  g17383(.A(new_n19813_), .B(new_n19812_), .C(new_n12509_), .Y(new_n19820_));
  AOI21X1  g17384(.A0(new_n19760_), .A1(pi0619), .B0(pi1159), .Y(new_n19821_));
  AND2X1   g17385(.A(new_n19821_), .B(new_n19820_), .Y(new_n19822_));
  OR2X1    g17386(.A(new_n19822_), .B(new_n12517_), .Y(new_n19823_));
  OAI22X1  g17387(.A0(new_n19823_), .A1(new_n19819_), .B0(new_n19817_), .B1(new_n19811_), .Y(new_n19824_));
  MX2X1    g17388(.A(new_n19824_), .B(new_n19808_), .S0(new_n11766_), .Y(new_n19825_));
  MX2X1    g17389(.A(new_n19809_), .B(new_n19779_), .S0(new_n12531_), .Y(new_n19826_));
  AOI21X1  g17390(.A0(new_n19826_), .A1(pi0626), .B0(pi0641), .Y(new_n19827_));
  OAI21X1  g17391(.A0(new_n19825_), .A1(pi0626), .B0(new_n19827_), .Y(new_n19828_));
  AND2X1   g17392(.A(new_n19813_), .B(new_n19812_), .Y(new_n19829_));
  AOI22X1  g17393(.A0(new_n19821_), .A1(new_n19820_), .B0(new_n19815_), .B1(new_n19814_), .Y(new_n19830_));
  MX2X1    g17394(.A(new_n19830_), .B(new_n19829_), .S0(new_n11766_), .Y(new_n19831_));
  AOI21X1  g17395(.A0(new_n19779_), .A1(pi0626), .B0(new_n12543_), .Y(new_n19832_));
  OAI21X1  g17396(.A0(new_n19831_), .A1(pi0626), .B0(new_n19832_), .Y(new_n19833_));
  AND2X1   g17397(.A(new_n19833_), .B(new_n12548_), .Y(new_n19834_));
  AOI21X1  g17398(.A0(new_n19826_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n19835_));
  OAI21X1  g17399(.A0(new_n19825_), .A1(new_n12542_), .B0(new_n19835_), .Y(new_n19836_));
  AOI21X1  g17400(.A0(new_n19779_), .A1(new_n12542_), .B0(pi0641), .Y(new_n19837_));
  OAI21X1  g17401(.A0(new_n19831_), .A1(new_n12542_), .B0(new_n19837_), .Y(new_n19838_));
  AND2X1   g17402(.A(new_n19838_), .B(pi1158), .Y(new_n19839_));
  AOI22X1  g17403(.A0(new_n19839_), .A1(new_n19836_), .B0(new_n19834_), .B1(new_n19828_), .Y(new_n19840_));
  MX2X1    g17404(.A(new_n19840_), .B(new_n19825_), .S0(new_n11765_), .Y(new_n19841_));
  MX2X1    g17405(.A(new_n19831_), .B(new_n19760_), .S0(new_n12708_), .Y(new_n19842_));
  INVX1    g17406(.A(new_n19842_), .Y(new_n19843_));
  OAI21X1  g17407(.A0(new_n19843_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n19844_));
  AOI21X1  g17408(.A0(new_n19841_), .A1(new_n12554_), .B0(new_n19844_), .Y(new_n19845_));
  MX2X1    g17409(.A(new_n19826_), .B(new_n19779_), .S0(new_n12563_), .Y(new_n19846_));
  AOI21X1  g17410(.A0(new_n19760_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n19847_));
  OAI21X1  g17411(.A0(new_n19846_), .A1(new_n12554_), .B0(new_n19847_), .Y(new_n19848_));
  NAND2X1  g17412(.A(new_n19848_), .B(new_n12561_), .Y(new_n19849_));
  OAI21X1  g17413(.A0(new_n19843_), .A1(pi0628), .B0(pi1156), .Y(new_n19850_));
  AOI21X1  g17414(.A0(new_n19841_), .A1(pi0628), .B0(new_n19850_), .Y(new_n19851_));
  AOI21X1  g17415(.A0(new_n19760_), .A1(pi0628), .B0(pi1156), .Y(new_n19852_));
  OAI21X1  g17416(.A0(new_n19846_), .A1(pi0628), .B0(new_n19852_), .Y(new_n19853_));
  NAND2X1  g17417(.A(new_n19853_), .B(pi0629), .Y(new_n19854_));
  OAI22X1  g17418(.A0(new_n19854_), .A1(new_n19851_), .B0(new_n19849_), .B1(new_n19845_), .Y(new_n19855_));
  AND2X1   g17419(.A(new_n19841_), .B(new_n11764_), .Y(new_n19856_));
  AOI21X1  g17420(.A0(new_n19855_), .A1(pi0792), .B0(new_n19856_), .Y(new_n19857_));
  MX2X1    g17421(.A(new_n19843_), .B(new_n19779_), .S0(new_n12580_), .Y(new_n19858_));
  INVX1    g17422(.A(new_n19858_), .Y(new_n19859_));
  AOI21X1  g17423(.A0(new_n19859_), .A1(pi0647), .B0(pi1157), .Y(new_n19860_));
  OAI21X1  g17424(.A0(new_n19857_), .A1(pi0647), .B0(new_n19860_), .Y(new_n19861_));
  INVX1    g17425(.A(new_n19846_), .Y(new_n19862_));
  AND2X1   g17426(.A(new_n19853_), .B(new_n19848_), .Y(new_n19863_));
  MX2X1    g17427(.A(new_n19863_), .B(new_n19862_), .S0(new_n11764_), .Y(new_n19864_));
  INVX1    g17428(.A(new_n19864_), .Y(new_n19865_));
  AOI21X1  g17429(.A0(new_n19760_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n19866_));
  OAI21X1  g17430(.A0(new_n19865_), .A1(new_n12577_), .B0(new_n19866_), .Y(new_n19867_));
  AND2X1   g17431(.A(new_n19867_), .B(new_n12592_), .Y(new_n19868_));
  AOI21X1  g17432(.A0(new_n19859_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n19869_));
  OAI21X1  g17433(.A0(new_n19857_), .A1(new_n12577_), .B0(new_n19869_), .Y(new_n19870_));
  AOI21X1  g17434(.A0(new_n19760_), .A1(pi0647), .B0(pi1157), .Y(new_n19871_));
  OAI21X1  g17435(.A0(new_n19865_), .A1(pi0647), .B0(new_n19871_), .Y(new_n19872_));
  AND2X1   g17436(.A(new_n19872_), .B(pi0630), .Y(new_n19873_));
  AOI22X1  g17437(.A0(new_n19873_), .A1(new_n19870_), .B0(new_n19868_), .B1(new_n19861_), .Y(new_n19874_));
  MX2X1    g17438(.A(new_n19874_), .B(new_n19857_), .S0(new_n11763_), .Y(new_n19875_));
  AND2X1   g17439(.A(new_n19872_), .B(new_n19867_), .Y(new_n19876_));
  MX2X1    g17440(.A(new_n19876_), .B(new_n19864_), .S0(new_n11763_), .Y(new_n19877_));
  AOI21X1  g17441(.A0(new_n19877_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n19878_));
  OAI21X1  g17442(.A0(new_n19875_), .A1(new_n12612_), .B0(new_n19878_), .Y(new_n19879_));
  MX2X1    g17443(.A(new_n19859_), .B(new_n19760_), .S0(new_n12604_), .Y(new_n19880_));
  OAI21X1  g17444(.A0(new_n19779_), .A1(pi0644), .B0(new_n12608_), .Y(new_n19881_));
  AOI21X1  g17445(.A0(new_n19880_), .A1(pi0644), .B0(new_n19881_), .Y(new_n19882_));
  NOR2X1   g17446(.A(new_n19882_), .B(new_n11762_), .Y(new_n19883_));
  AND2X1   g17447(.A(new_n19883_), .B(new_n19879_), .Y(new_n19884_));
  OR2X1    g17448(.A(new_n19857_), .B(pi0787), .Y(new_n19885_));
  OAI21X1  g17449(.A0(new_n19874_), .A1(new_n11763_), .B0(new_n19885_), .Y(new_n19886_));
  AND2X1   g17450(.A(new_n19877_), .B(pi0644), .Y(new_n19887_));
  OR2X1    g17451(.A(new_n19887_), .B(pi0715), .Y(new_n19888_));
  AOI21X1  g17452(.A0(new_n19886_), .A1(new_n12612_), .B0(new_n19888_), .Y(new_n19889_));
  OAI21X1  g17453(.A0(new_n19779_), .A1(new_n12612_), .B0(pi0715), .Y(new_n19890_));
  AOI21X1  g17454(.A0(new_n19880_), .A1(new_n12612_), .B0(new_n19890_), .Y(new_n19891_));
  OR2X1    g17455(.A(new_n19891_), .B(pi1160), .Y(new_n19892_));
  OAI21X1  g17456(.A0(new_n19892_), .A1(new_n19889_), .B0(pi0790), .Y(new_n19893_));
  AOI21X1  g17457(.A0(new_n19875_), .A1(new_n12766_), .B0(po1038), .Y(new_n19894_));
  OAI21X1  g17458(.A0(new_n19893_), .A1(new_n19884_), .B0(new_n19894_), .Y(new_n19895_));
  AOI21X1  g17459(.A0(po1038), .A1(new_n7436_), .B0(pi0832), .Y(new_n19896_));
  AOI21X1  g17460(.A0(pi1093), .A1(pi1092), .B0(pi0188), .Y(new_n19897_));
  INVX1    g17461(.A(new_n19897_), .Y(new_n19898_));
  AOI21X1  g17462(.A0(new_n12056_), .A1(new_n15345_), .B0(new_n19897_), .Y(new_n19899_));
  AOI21X1  g17463(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n19899_), .Y(new_n19900_));
  INVX1    g17464(.A(new_n19899_), .Y(new_n19901_));
  AOI21X1  g17465(.A0(new_n19901_), .A1(new_n14331_), .B0(new_n12463_), .Y(new_n19902_));
  AOI21X1  g17466(.A0(new_n19900_), .A1(new_n12646_), .B0(pi1155), .Y(new_n19903_));
  OAI21X1  g17467(.A0(new_n19903_), .A1(new_n19902_), .B0(pi0785), .Y(new_n19904_));
  OAI21X1  g17468(.A0(new_n19900_), .A1(pi0785), .B0(new_n19904_), .Y(new_n19905_));
  INVX1    g17469(.A(new_n19905_), .Y(new_n19906_));
  AOI21X1  g17470(.A0(new_n19906_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n19907_));
  AOI21X1  g17471(.A0(new_n19906_), .A1(new_n12655_), .B0(pi1154), .Y(new_n19908_));
  NOR2X1   g17472(.A(new_n19908_), .B(new_n19907_), .Y(new_n19909_));
  MX2X1    g17473(.A(new_n19909_), .B(new_n19906_), .S0(new_n11767_), .Y(new_n19910_));
  NOR2X1   g17474(.A(new_n19910_), .B(pi0789), .Y(new_n19911_));
  INVX1    g17475(.A(new_n19910_), .Y(new_n19912_));
  AOI21X1  g17476(.A0(new_n19897_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n19913_));
  OAI21X1  g17477(.A0(new_n19912_), .A1(new_n12509_), .B0(new_n19913_), .Y(new_n19914_));
  AOI21X1  g17478(.A0(new_n19897_), .A1(pi0619), .B0(pi1159), .Y(new_n19915_));
  OAI21X1  g17479(.A0(new_n19912_), .A1(pi0619), .B0(new_n19915_), .Y(new_n19916_));
  AOI21X1  g17480(.A0(new_n19916_), .A1(new_n19914_), .B0(new_n11766_), .Y(new_n19917_));
  NOR2X1   g17481(.A(new_n19917_), .B(new_n19911_), .Y(new_n19918_));
  INVX1    g17482(.A(new_n19918_), .Y(new_n19919_));
  MX2X1    g17483(.A(new_n19919_), .B(new_n19898_), .S0(new_n12708_), .Y(new_n19920_));
  MX2X1    g17484(.A(new_n19920_), .B(new_n19898_), .S0(new_n12580_), .Y(new_n19921_));
  AOI21X1  g17485(.A0(new_n12439_), .A1(pi0705), .B0(new_n19897_), .Y(new_n19922_));
  AND3X1   g17486(.A(new_n12439_), .B(pi0705), .C(new_n12363_), .Y(new_n19923_));
  NOR2X1   g17487(.A(new_n19923_), .B(new_n19922_), .Y(new_n19924_));
  NOR2X1   g17488(.A(new_n19897_), .B(pi1153), .Y(new_n19925_));
  INVX1    g17489(.A(new_n19925_), .Y(new_n19926_));
  OAI22X1  g17490(.A0(new_n19926_), .A1(new_n19923_), .B0(new_n19924_), .B1(new_n12364_), .Y(new_n19927_));
  MX2X1    g17491(.A(new_n19927_), .B(new_n19922_), .S0(new_n11769_), .Y(new_n19928_));
  NOR4X1   g17492(.A(new_n19928_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n19929_));
  AND3X1   g17493(.A(new_n19929_), .B(new_n12739_), .C(new_n12718_), .Y(new_n19930_));
  INVX1    g17494(.A(new_n19930_), .Y(new_n19931_));
  AOI21X1  g17495(.A0(new_n19897_), .A1(pi0647), .B0(pi1157), .Y(new_n19932_));
  OAI21X1  g17496(.A0(new_n19931_), .A1(pi0647), .B0(new_n19932_), .Y(new_n19933_));
  MX2X1    g17497(.A(new_n19930_), .B(new_n19897_), .S0(new_n12577_), .Y(new_n19934_));
  OAI22X1  g17498(.A0(new_n19934_), .A1(new_n14242_), .B0(new_n19933_), .B1(new_n12592_), .Y(new_n19935_));
  AOI21X1  g17499(.A0(new_n19921_), .A1(new_n14326_), .B0(new_n19935_), .Y(new_n19936_));
  AOI21X1  g17500(.A0(new_n19898_), .A1(pi0626), .B0(new_n16218_), .Y(new_n19937_));
  OAI21X1  g17501(.A0(new_n19918_), .A1(pi0626), .B0(new_n19937_), .Y(new_n19938_));
  AOI21X1  g17502(.A0(new_n19898_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n19939_));
  OAI21X1  g17503(.A0(new_n19918_), .A1(new_n12542_), .B0(new_n19939_), .Y(new_n19940_));
  NAND2X1  g17504(.A(new_n19929_), .B(new_n12637_), .Y(new_n19941_));
  AND3X1   g17505(.A(new_n19941_), .B(new_n19940_), .C(new_n19938_), .Y(new_n19942_));
  NOR2X1   g17506(.A(new_n19942_), .B(new_n11765_), .Y(new_n19943_));
  INVX1    g17507(.A(new_n19943_), .Y(new_n19944_));
  NOR2X1   g17508(.A(new_n19922_), .B(new_n11991_), .Y(new_n19945_));
  MX2X1    g17509(.A(new_n19901_), .B(new_n12363_), .S0(new_n19945_), .Y(new_n19946_));
  NOR2X1   g17510(.A(new_n19946_), .B(new_n19926_), .Y(new_n19947_));
  OAI21X1  g17511(.A0(new_n19924_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n19948_));
  NOR2X1   g17512(.A(new_n19948_), .B(new_n19947_), .Y(new_n19949_));
  OR3X1    g17513(.A(new_n19922_), .B(new_n11991_), .C(new_n12363_), .Y(new_n19950_));
  AND2X1   g17514(.A(new_n19899_), .B(pi1153), .Y(new_n19951_));
  OAI21X1  g17515(.A0(new_n19926_), .A1(new_n19923_), .B0(pi0608), .Y(new_n19952_));
  AOI21X1  g17516(.A0(new_n19951_), .A1(new_n19950_), .B0(new_n19952_), .Y(new_n19953_));
  OAI21X1  g17517(.A0(new_n19953_), .A1(new_n19949_), .B0(pi0778), .Y(new_n19954_));
  OAI21X1  g17518(.A0(new_n19945_), .A1(new_n19901_), .B0(new_n11769_), .Y(new_n19955_));
  NAND2X1  g17519(.A(new_n19955_), .B(new_n19954_), .Y(new_n19956_));
  INVX1    g17520(.A(new_n19956_), .Y(new_n19957_));
  OAI21X1  g17521(.A0(new_n19928_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n19958_));
  AOI21X1  g17522(.A0(new_n19956_), .A1(new_n12462_), .B0(new_n19958_), .Y(new_n19959_));
  NOR3X1   g17523(.A(new_n19959_), .B(new_n19902_), .C(pi0660), .Y(new_n19960_));
  OAI21X1  g17524(.A0(new_n19928_), .A1(pi0609), .B0(pi1155), .Y(new_n19961_));
  AOI21X1  g17525(.A0(new_n19956_), .A1(pi0609), .B0(new_n19961_), .Y(new_n19962_));
  NOR3X1   g17526(.A(new_n19962_), .B(new_n19903_), .C(new_n12468_), .Y(new_n19963_));
  NOR2X1   g17527(.A(new_n19963_), .B(new_n19960_), .Y(new_n19964_));
  MX2X1    g17528(.A(new_n19964_), .B(new_n19957_), .S0(new_n11768_), .Y(new_n19965_));
  OR3X1    g17529(.A(new_n19928_), .B(new_n12630_), .C(new_n12486_), .Y(new_n19966_));
  AND2X1   g17530(.A(new_n19966_), .B(new_n12487_), .Y(new_n19967_));
  OAI21X1  g17531(.A0(new_n19965_), .A1(pi0618), .B0(new_n19967_), .Y(new_n19968_));
  NOR2X1   g17532(.A(new_n19907_), .B(pi0627), .Y(new_n19969_));
  NOR3X1   g17533(.A(new_n19928_), .B(new_n12630_), .C(pi0618), .Y(new_n19970_));
  NOR2X1   g17534(.A(new_n19970_), .B(new_n12487_), .Y(new_n19971_));
  OAI21X1  g17535(.A0(new_n19965_), .A1(new_n12486_), .B0(new_n19971_), .Y(new_n19972_));
  NOR2X1   g17536(.A(new_n19908_), .B(new_n12494_), .Y(new_n19973_));
  AOI22X1  g17537(.A0(new_n19973_), .A1(new_n19972_), .B0(new_n19969_), .B1(new_n19968_), .Y(new_n19974_));
  MX2X1    g17538(.A(new_n19974_), .B(new_n19965_), .S0(new_n11767_), .Y(new_n19975_));
  OR4X1    g17539(.A(new_n19928_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n19976_));
  AND2X1   g17540(.A(new_n19976_), .B(new_n12510_), .Y(new_n19977_));
  OAI21X1  g17541(.A0(new_n19975_), .A1(pi0619), .B0(new_n19977_), .Y(new_n19978_));
  AND3X1   g17542(.A(new_n19978_), .B(new_n19914_), .C(new_n12517_), .Y(new_n19979_));
  NOR4X1   g17543(.A(new_n19928_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n19980_));
  NOR2X1   g17544(.A(new_n19980_), .B(new_n12510_), .Y(new_n19981_));
  OAI21X1  g17545(.A0(new_n19975_), .A1(new_n12509_), .B0(new_n19981_), .Y(new_n19982_));
  AND2X1   g17546(.A(new_n19916_), .B(pi0648), .Y(new_n19983_));
  AOI21X1  g17547(.A0(new_n19983_), .A1(new_n19982_), .B0(new_n11766_), .Y(new_n19984_));
  INVX1    g17548(.A(new_n19984_), .Y(new_n19985_));
  AOI21X1  g17549(.A0(new_n19975_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n19986_));
  OAI21X1  g17550(.A0(new_n19985_), .A1(new_n19979_), .B0(new_n19986_), .Y(new_n19987_));
  AOI21X1  g17551(.A0(new_n19987_), .A1(new_n19944_), .B0(new_n14125_), .Y(new_n19988_));
  INVX1    g17552(.A(new_n19920_), .Y(new_n19989_));
  AND2X1   g17553(.A(new_n19929_), .B(new_n12718_), .Y(new_n19990_));
  AOI22X1  g17554(.A0(new_n19990_), .A1(new_n14426_), .B0(new_n19989_), .B1(new_n12735_), .Y(new_n19991_));
  AOI22X1  g17555(.A0(new_n19990_), .A1(new_n14428_), .B0(new_n19989_), .B1(new_n12733_), .Y(new_n19992_));
  MX2X1    g17556(.A(new_n19992_), .B(new_n19991_), .S0(new_n12561_), .Y(new_n19993_));
  OAI21X1  g17557(.A0(new_n19993_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n19994_));
  OAI22X1  g17558(.A0(new_n19994_), .A1(new_n19988_), .B0(new_n19936_), .B1(new_n11763_), .Y(new_n19995_));
  INVX1    g17559(.A(new_n19995_), .Y(new_n19996_));
  OAI21X1  g17560(.A0(new_n19934_), .A1(new_n12578_), .B0(new_n19933_), .Y(new_n19997_));
  MX2X1    g17561(.A(new_n19997_), .B(new_n19931_), .S0(new_n11763_), .Y(new_n19998_));
  OAI21X1  g17562(.A0(new_n19998_), .A1(pi0644), .B0(pi0715), .Y(new_n19999_));
  AOI21X1  g17563(.A0(new_n19996_), .A1(pi0644), .B0(new_n19999_), .Y(new_n20000_));
  OR3X1    g17564(.A(new_n19898_), .B(new_n12603_), .C(new_n11763_), .Y(new_n20001_));
  OAI21X1  g17565(.A0(new_n19921_), .A1(new_n12604_), .B0(new_n20001_), .Y(new_n20002_));
  OAI21X1  g17566(.A0(new_n19898_), .A1(pi0644), .B0(new_n12608_), .Y(new_n20003_));
  AOI21X1  g17567(.A0(new_n20002_), .A1(pi0644), .B0(new_n20003_), .Y(new_n20004_));
  OR2X1    g17568(.A(new_n20004_), .B(new_n11762_), .Y(new_n20005_));
  OAI21X1  g17569(.A0(new_n19998_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n20006_));
  AOI21X1  g17570(.A0(new_n19996_), .A1(new_n12612_), .B0(new_n20006_), .Y(new_n20007_));
  OAI21X1  g17571(.A0(new_n19898_), .A1(new_n12612_), .B0(pi0715), .Y(new_n20008_));
  AOI21X1  g17572(.A0(new_n20002_), .A1(new_n12612_), .B0(new_n20008_), .Y(new_n20009_));
  OR2X1    g17573(.A(new_n20009_), .B(pi1160), .Y(new_n20010_));
  OAI22X1  g17574(.A0(new_n20010_), .A1(new_n20007_), .B0(new_n20005_), .B1(new_n20000_), .Y(new_n20011_));
  OAI21X1  g17575(.A0(new_n19995_), .A1(pi0790), .B0(pi0832), .Y(new_n20012_));
  AOI21X1  g17576(.A0(new_n20011_), .A1(pi0790), .B0(new_n20012_), .Y(new_n20013_));
  AOI21X1  g17577(.A0(new_n19896_), .A1(new_n19895_), .B0(new_n20013_), .Y(po0345));
  AND2X1   g17578(.A(new_n12034_), .B(pi0772), .Y(new_n20015_));
  OAI21X1  g17579(.A0(new_n20015_), .A1(new_n15285_), .B0(pi0039), .Y(new_n20016_));
  AOI21X1  g17580(.A0(new_n11821_), .A1(new_n15306_), .B0(pi0039), .Y(new_n20017_));
  OAI21X1  g17581(.A0(new_n11975_), .A1(new_n15306_), .B0(new_n20017_), .Y(new_n20018_));
  AOI21X1  g17582(.A0(new_n20018_), .A1(new_n20016_), .B0(new_n7872_), .Y(new_n20019_));
  AND3X1   g17583(.A(new_n12074_), .B(pi0772), .C(new_n7872_), .Y(new_n20020_));
  OAI21X1  g17584(.A0(new_n20020_), .A1(new_n20019_), .B0(new_n2979_), .Y(new_n20021_));
  NOR2X1   g17585(.A(new_n12077_), .B(pi0189), .Y(new_n20022_));
  AOI21X1  g17586(.A0(new_n11991_), .A1(pi0772), .B0(new_n12771_), .Y(new_n20023_));
  NOR3X1   g17587(.A(new_n20023_), .B(new_n20022_), .C(new_n2979_), .Y(new_n20024_));
  INVX1    g17588(.A(new_n20024_), .Y(new_n20025_));
  AND3X1   g17589(.A(new_n20025_), .B(new_n20021_), .C(new_n15292_), .Y(new_n20026_));
  AOI21X1  g17590(.A0(new_n12213_), .A1(new_n7872_), .B0(pi0772), .Y(new_n20027_));
  OAI21X1  g17591(.A0(new_n12155_), .A1(new_n7872_), .B0(new_n20027_), .Y(new_n20028_));
  AOI21X1  g17592(.A0(new_n12301_), .A1(pi0189), .B0(new_n15306_), .Y(new_n20029_));
  OAI21X1  g17593(.A0(new_n12260_), .A1(pi0189), .B0(new_n20029_), .Y(new_n20030_));
  AND3X1   g17594(.A(new_n20030_), .B(new_n20028_), .C(pi0039), .Y(new_n20031_));
  OAI21X1  g17595(.A0(new_n12315_), .A1(new_n7872_), .B0(new_n15306_), .Y(new_n20032_));
  AOI21X1  g17596(.A0(new_n12332_), .A1(new_n7872_), .B0(new_n20032_), .Y(new_n20033_));
  NOR4X1   g17597(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(new_n7872_), .Y(new_n20034_));
  OAI21X1  g17598(.A0(new_n12800_), .A1(pi0189), .B0(pi0772), .Y(new_n20035_));
  OAI21X1  g17599(.A0(new_n20035_), .A1(new_n20034_), .B0(new_n2939_), .Y(new_n20036_));
  OAI21X1  g17600(.A0(new_n20036_), .A1(new_n20033_), .B0(new_n2979_), .Y(new_n20037_));
  NOR3X1   g17601(.A(new_n20024_), .B(new_n13547_), .C(new_n15292_), .Y(new_n20038_));
  OAI21X1  g17602(.A0(new_n20037_), .A1(new_n20031_), .B0(new_n20038_), .Y(new_n20039_));
  NAND2X1  g17603(.A(new_n20039_), .B(new_n3103_), .Y(new_n20040_));
  OAI22X1  g17604(.A0(new_n20040_), .A1(new_n20026_), .B0(new_n3103_), .B1(new_n7872_), .Y(new_n20041_));
  OR2X1    g17605(.A(new_n20041_), .B(pi0625), .Y(new_n20042_));
  AND2X1   g17606(.A(new_n20025_), .B(new_n20021_), .Y(new_n20043_));
  MX2X1    g17607(.A(new_n20043_), .B(new_n7872_), .S0(new_n11770_), .Y(new_n20044_));
  AOI21X1  g17608(.A0(new_n20044_), .A1(pi0625), .B0(pi1153), .Y(new_n20045_));
  AOI21X1  g17609(.A0(new_n12447_), .A1(new_n3103_), .B0(new_n7872_), .Y(new_n20046_));
  NOR4X1   g17610(.A(new_n10543_), .B(new_n15292_), .C(pi0100), .D(pi0087), .Y(new_n20047_));
  OAI21X1  g17611(.A0(new_n13870_), .A1(pi0189), .B0(new_n2979_), .Y(new_n20048_));
  AOI21X1  g17612(.A0(new_n13868_), .A1(pi0189), .B0(new_n20048_), .Y(new_n20049_));
  OAI21X1  g17613(.A0(new_n20022_), .A1(new_n13874_), .B0(new_n20047_), .Y(new_n20050_));
  OAI22X1  g17614(.A0(new_n20050_), .A1(new_n20049_), .B0(new_n20047_), .B1(new_n20046_), .Y(new_n20051_));
  OAI21X1  g17615(.A0(new_n20046_), .A1(pi0625), .B0(pi1153), .Y(new_n20052_));
  AOI21X1  g17616(.A0(new_n20051_), .A1(pi0625), .B0(new_n20052_), .Y(new_n20053_));
  OR2X1    g17617(.A(new_n20053_), .B(pi0608), .Y(new_n20054_));
  AOI21X1  g17618(.A0(new_n20045_), .A1(new_n20042_), .B0(new_n20054_), .Y(new_n20055_));
  OR2X1    g17619(.A(new_n20041_), .B(new_n12363_), .Y(new_n20056_));
  AOI21X1  g17620(.A0(new_n20044_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n20057_));
  OAI21X1  g17621(.A0(new_n20046_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n20058_));
  AOI21X1  g17622(.A0(new_n20051_), .A1(new_n12363_), .B0(new_n20058_), .Y(new_n20059_));
  OR2X1    g17623(.A(new_n20059_), .B(new_n12368_), .Y(new_n20060_));
  AOI21X1  g17624(.A0(new_n20057_), .A1(new_n20056_), .B0(new_n20060_), .Y(new_n20061_));
  OAI21X1  g17625(.A0(new_n20061_), .A1(new_n20055_), .B0(pi0778), .Y(new_n20062_));
  OR2X1    g17626(.A(new_n20041_), .B(pi0778), .Y(new_n20063_));
  AOI21X1  g17627(.A0(new_n20063_), .A1(new_n20062_), .B0(pi0609), .Y(new_n20064_));
  OR2X1    g17628(.A(new_n20051_), .B(pi0778), .Y(new_n20065_));
  NOR2X1   g17629(.A(new_n20059_), .B(new_n20053_), .Y(new_n20066_));
  OAI21X1  g17630(.A0(new_n20066_), .A1(new_n11769_), .B0(new_n20065_), .Y(new_n20067_));
  OAI21X1  g17631(.A0(new_n20067_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n20068_));
  NOR2X1   g17632(.A(new_n20046_), .B(new_n12474_), .Y(new_n20069_));
  AOI21X1  g17633(.A0(new_n20044_), .A1(new_n12474_), .B0(new_n20069_), .Y(new_n20070_));
  INVX1    g17634(.A(new_n20046_), .Y(new_n20071_));
  AOI21X1  g17635(.A0(new_n20071_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n20072_));
  OAI21X1  g17636(.A0(new_n20070_), .A1(new_n12462_), .B0(new_n20072_), .Y(new_n20073_));
  AND2X1   g17637(.A(new_n20073_), .B(new_n12468_), .Y(new_n20074_));
  OAI21X1  g17638(.A0(new_n20068_), .A1(new_n20064_), .B0(new_n20074_), .Y(new_n20075_));
  AOI21X1  g17639(.A0(new_n20063_), .A1(new_n20062_), .B0(new_n12462_), .Y(new_n20076_));
  OAI21X1  g17640(.A0(new_n20067_), .A1(pi0609), .B0(pi1155), .Y(new_n20077_));
  AOI21X1  g17641(.A0(new_n20071_), .A1(pi0609), .B0(pi1155), .Y(new_n20078_));
  OAI21X1  g17642(.A0(new_n20070_), .A1(pi0609), .B0(new_n20078_), .Y(new_n20079_));
  AND2X1   g17643(.A(new_n20079_), .B(pi0660), .Y(new_n20080_));
  OAI21X1  g17644(.A0(new_n20077_), .A1(new_n20076_), .B0(new_n20080_), .Y(new_n20081_));
  AOI21X1  g17645(.A0(new_n20081_), .A1(new_n20075_), .B0(new_n11768_), .Y(new_n20082_));
  AOI21X1  g17646(.A0(new_n20063_), .A1(new_n20062_), .B0(pi0785), .Y(new_n20083_));
  OAI21X1  g17647(.A0(new_n20083_), .A1(new_n20082_), .B0(new_n12486_), .Y(new_n20084_));
  OR2X1    g17648(.A(new_n20046_), .B(new_n13910_), .Y(new_n20085_));
  OAI21X1  g17649(.A0(new_n20067_), .A1(new_n12490_), .B0(new_n20085_), .Y(new_n20086_));
  AOI21X1  g17650(.A0(new_n20086_), .A1(pi0618), .B0(pi1154), .Y(new_n20087_));
  AOI21X1  g17651(.A0(new_n20079_), .A1(new_n20073_), .B0(new_n11768_), .Y(new_n20088_));
  AOI21X1  g17652(.A0(new_n20070_), .A1(new_n11768_), .B0(new_n20088_), .Y(new_n20089_));
  OAI21X1  g17653(.A0(new_n20046_), .A1(pi0618), .B0(pi1154), .Y(new_n20090_));
  AOI21X1  g17654(.A0(new_n20089_), .A1(pi0618), .B0(new_n20090_), .Y(new_n20091_));
  OR2X1    g17655(.A(new_n20091_), .B(pi0627), .Y(new_n20092_));
  AOI21X1  g17656(.A0(new_n20087_), .A1(new_n20084_), .B0(new_n20092_), .Y(new_n20093_));
  OAI21X1  g17657(.A0(new_n20083_), .A1(new_n20082_), .B0(pi0618), .Y(new_n20094_));
  AOI21X1  g17658(.A0(new_n20086_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20095_));
  OAI21X1  g17659(.A0(new_n20046_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20096_));
  AOI21X1  g17660(.A0(new_n20089_), .A1(new_n12486_), .B0(new_n20096_), .Y(new_n20097_));
  OR2X1    g17661(.A(new_n20097_), .B(new_n12494_), .Y(new_n20098_));
  AOI21X1  g17662(.A0(new_n20095_), .A1(new_n20094_), .B0(new_n20098_), .Y(new_n20099_));
  OAI21X1  g17663(.A0(new_n20099_), .A1(new_n20093_), .B0(pi0781), .Y(new_n20100_));
  OAI21X1  g17664(.A0(new_n20083_), .A1(new_n20082_), .B0(new_n11767_), .Y(new_n20101_));
  AOI21X1  g17665(.A0(new_n20101_), .A1(new_n20100_), .B0(pi0619), .Y(new_n20102_));
  MX2X1    g17666(.A(new_n20086_), .B(new_n20071_), .S0(new_n12513_), .Y(new_n20103_));
  INVX1    g17667(.A(new_n20103_), .Y(new_n20104_));
  OAI21X1  g17668(.A0(new_n20104_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n20105_));
  OAI21X1  g17669(.A0(new_n20097_), .A1(new_n20091_), .B0(pi0781), .Y(new_n20106_));
  OAI21X1  g17670(.A0(new_n20089_), .A1(pi0781), .B0(new_n20106_), .Y(new_n20107_));
  AOI21X1  g17671(.A0(new_n20071_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n20108_));
  OAI21X1  g17672(.A0(new_n20107_), .A1(new_n12509_), .B0(new_n20108_), .Y(new_n20109_));
  AND2X1   g17673(.A(new_n20109_), .B(new_n12517_), .Y(new_n20110_));
  OAI21X1  g17674(.A0(new_n20105_), .A1(new_n20102_), .B0(new_n20110_), .Y(new_n20111_));
  AOI21X1  g17675(.A0(new_n20101_), .A1(new_n20100_), .B0(new_n12509_), .Y(new_n20112_));
  OAI21X1  g17676(.A0(new_n20104_), .A1(pi0619), .B0(pi1159), .Y(new_n20113_));
  AOI21X1  g17677(.A0(new_n20071_), .A1(pi0619), .B0(pi1159), .Y(new_n20114_));
  OAI21X1  g17678(.A0(new_n20107_), .A1(pi0619), .B0(new_n20114_), .Y(new_n20115_));
  AND2X1   g17679(.A(new_n20115_), .B(pi0648), .Y(new_n20116_));
  OAI21X1  g17680(.A0(new_n20113_), .A1(new_n20112_), .B0(new_n20116_), .Y(new_n20117_));
  AOI21X1  g17681(.A0(new_n20117_), .A1(new_n20111_), .B0(new_n11766_), .Y(new_n20118_));
  AOI21X1  g17682(.A0(new_n20101_), .A1(new_n20100_), .B0(pi0789), .Y(new_n20119_));
  OR3X1    g17683(.A(new_n20119_), .B(new_n20118_), .C(pi0788), .Y(new_n20120_));
  OR3X1    g17684(.A(new_n20119_), .B(new_n20118_), .C(pi0626), .Y(new_n20121_));
  MX2X1    g17685(.A(new_n20104_), .B(new_n20046_), .S0(new_n12531_), .Y(new_n20122_));
  AOI21X1  g17686(.A0(new_n20122_), .A1(pi0626), .B0(pi0641), .Y(new_n20123_));
  NAND2X1  g17687(.A(new_n20115_), .B(new_n20109_), .Y(new_n20124_));
  MX2X1    g17688(.A(new_n20124_), .B(new_n20107_), .S0(new_n11766_), .Y(new_n20125_));
  OAI21X1  g17689(.A0(new_n20071_), .A1(new_n12542_), .B0(pi0641), .Y(new_n20126_));
  AOI21X1  g17690(.A0(new_n20125_), .A1(new_n12542_), .B0(new_n20126_), .Y(new_n20127_));
  OR2X1    g17691(.A(new_n20127_), .B(pi1158), .Y(new_n20128_));
  AOI21X1  g17692(.A0(new_n20123_), .A1(new_n20121_), .B0(new_n20128_), .Y(new_n20129_));
  OR3X1    g17693(.A(new_n20119_), .B(new_n20118_), .C(new_n12542_), .Y(new_n20130_));
  AOI21X1  g17694(.A0(new_n20122_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n20131_));
  OAI21X1  g17695(.A0(new_n20071_), .A1(pi0626), .B0(new_n12543_), .Y(new_n20132_));
  AOI21X1  g17696(.A0(new_n20125_), .A1(pi0626), .B0(new_n20132_), .Y(new_n20133_));
  OR2X1    g17697(.A(new_n20133_), .B(new_n12548_), .Y(new_n20134_));
  AOI21X1  g17698(.A0(new_n20131_), .A1(new_n20130_), .B0(new_n20134_), .Y(new_n20135_));
  OAI21X1  g17699(.A0(new_n20135_), .A1(new_n20129_), .B0(pi0788), .Y(new_n20136_));
  AND3X1   g17700(.A(new_n20136_), .B(new_n20120_), .C(new_n12554_), .Y(new_n20137_));
  MX2X1    g17701(.A(new_n20125_), .B(new_n20046_), .S0(new_n12708_), .Y(new_n20138_));
  OAI21X1  g17702(.A0(new_n20138_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n20139_));
  AND2X1   g17703(.A(new_n20046_), .B(new_n12563_), .Y(new_n20140_));
  AOI21X1  g17704(.A0(new_n20122_), .A1(new_n13356_), .B0(new_n20140_), .Y(new_n20141_));
  OAI21X1  g17705(.A0(new_n20046_), .A1(pi0628), .B0(pi1156), .Y(new_n20142_));
  AOI21X1  g17706(.A0(new_n20141_), .A1(pi0628), .B0(new_n20142_), .Y(new_n20143_));
  NOR2X1   g17707(.A(new_n20143_), .B(pi0629), .Y(new_n20144_));
  OAI21X1  g17708(.A0(new_n20139_), .A1(new_n20137_), .B0(new_n20144_), .Y(new_n20145_));
  AND3X1   g17709(.A(new_n20136_), .B(new_n20120_), .C(pi0628), .Y(new_n20146_));
  OAI21X1  g17710(.A0(new_n20138_), .A1(pi0628), .B0(pi1156), .Y(new_n20147_));
  OAI21X1  g17711(.A0(new_n20046_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n20148_));
  AOI21X1  g17712(.A0(new_n20141_), .A1(new_n12554_), .B0(new_n20148_), .Y(new_n20149_));
  NOR2X1   g17713(.A(new_n20149_), .B(new_n12561_), .Y(new_n20150_));
  OAI21X1  g17714(.A0(new_n20147_), .A1(new_n20146_), .B0(new_n20150_), .Y(new_n20151_));
  AOI21X1  g17715(.A0(new_n20151_), .A1(new_n20145_), .B0(new_n11764_), .Y(new_n20152_));
  AND3X1   g17716(.A(new_n20136_), .B(new_n20120_), .C(new_n11764_), .Y(new_n20153_));
  OAI21X1  g17717(.A0(new_n20153_), .A1(new_n20152_), .B0(new_n12577_), .Y(new_n20154_));
  MX2X1    g17718(.A(new_n20138_), .B(new_n20046_), .S0(new_n12580_), .Y(new_n20155_));
  INVX1    g17719(.A(new_n20155_), .Y(new_n20156_));
  AOI21X1  g17720(.A0(new_n20156_), .A1(pi0647), .B0(pi1157), .Y(new_n20157_));
  NOR2X1   g17721(.A(new_n20149_), .B(new_n20143_), .Y(new_n20158_));
  MX2X1    g17722(.A(new_n20158_), .B(new_n20141_), .S0(new_n11764_), .Y(new_n20159_));
  OAI21X1  g17723(.A0(new_n20046_), .A1(pi0647), .B0(pi1157), .Y(new_n20160_));
  AOI21X1  g17724(.A0(new_n20159_), .A1(pi0647), .B0(new_n20160_), .Y(new_n20161_));
  OR2X1    g17725(.A(new_n20161_), .B(pi0630), .Y(new_n20162_));
  AOI21X1  g17726(.A0(new_n20157_), .A1(new_n20154_), .B0(new_n20162_), .Y(new_n20163_));
  OAI21X1  g17727(.A0(new_n20153_), .A1(new_n20152_), .B0(pi0647), .Y(new_n20164_));
  AOI21X1  g17728(.A0(new_n20156_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n20165_));
  OAI21X1  g17729(.A0(new_n20046_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n20166_));
  AOI21X1  g17730(.A0(new_n20159_), .A1(new_n12577_), .B0(new_n20166_), .Y(new_n20167_));
  OR2X1    g17731(.A(new_n20167_), .B(new_n12592_), .Y(new_n20168_));
  AOI21X1  g17732(.A0(new_n20165_), .A1(new_n20164_), .B0(new_n20168_), .Y(new_n20169_));
  OAI21X1  g17733(.A0(new_n20169_), .A1(new_n20163_), .B0(pi0787), .Y(new_n20170_));
  OAI21X1  g17734(.A0(new_n20153_), .A1(new_n20152_), .B0(new_n11763_), .Y(new_n20171_));
  AOI21X1  g17735(.A0(new_n20171_), .A1(new_n20170_), .B0(new_n12612_), .Y(new_n20172_));
  OAI21X1  g17736(.A0(new_n20167_), .A1(new_n20161_), .B0(pi0787), .Y(new_n20173_));
  OAI21X1  g17737(.A0(new_n20159_), .A1(pi0787), .B0(new_n20173_), .Y(new_n20174_));
  OAI21X1  g17738(.A0(new_n20174_), .A1(pi0644), .B0(pi0715), .Y(new_n20175_));
  MX2X1    g17739(.A(new_n20155_), .B(new_n20046_), .S0(new_n12604_), .Y(new_n20176_));
  AOI21X1  g17740(.A0(new_n20071_), .A1(new_n12612_), .B0(pi0715), .Y(new_n20177_));
  OAI21X1  g17741(.A0(new_n20176_), .A1(new_n12612_), .B0(new_n20177_), .Y(new_n20178_));
  AND2X1   g17742(.A(new_n20178_), .B(pi1160), .Y(new_n20179_));
  OAI21X1  g17743(.A0(new_n20175_), .A1(new_n20172_), .B0(new_n20179_), .Y(new_n20180_));
  AOI21X1  g17744(.A0(new_n20171_), .A1(new_n20170_), .B0(pi0644), .Y(new_n20181_));
  OAI21X1  g17745(.A0(new_n20174_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n20182_));
  AOI21X1  g17746(.A0(new_n20071_), .A1(pi0644), .B0(new_n12608_), .Y(new_n20183_));
  OAI21X1  g17747(.A0(new_n20176_), .A1(pi0644), .B0(new_n20183_), .Y(new_n20184_));
  AND2X1   g17748(.A(new_n20184_), .B(new_n11762_), .Y(new_n20185_));
  OAI21X1  g17749(.A0(new_n20182_), .A1(new_n20181_), .B0(new_n20185_), .Y(new_n20186_));
  AND3X1   g17750(.A(new_n20186_), .B(new_n20180_), .C(pi0790), .Y(new_n20187_));
  AND3X1   g17751(.A(new_n20171_), .B(new_n20170_), .C(new_n12766_), .Y(new_n20188_));
  OR2X1    g17752(.A(new_n20188_), .B(new_n5103_), .Y(new_n20189_));
  AOI21X1  g17753(.A0(new_n5103_), .A1(new_n7872_), .B0(pi0057), .Y(new_n20190_));
  OAI21X1  g17754(.A0(new_n20189_), .A1(new_n20187_), .B0(new_n20190_), .Y(new_n20191_));
  AOI21X1  g17755(.A0(pi0189), .A1(pi0057), .B0(pi0832), .Y(new_n20192_));
  NOR2X1   g17756(.A(new_n2720_), .B(new_n7872_), .Y(new_n20193_));
  AOI21X1  g17757(.A0(new_n12056_), .A1(pi0772), .B0(new_n20193_), .Y(new_n20194_));
  OAI21X1  g17758(.A0(new_n14068_), .A1(new_n15292_), .B0(new_n20194_), .Y(new_n20195_));
  AND3X1   g17759(.A(new_n13443_), .B(pi0727), .C(pi0625), .Y(new_n20196_));
  INVX1    g17760(.A(new_n20196_), .Y(new_n20197_));
  AOI21X1  g17761(.A0(new_n20197_), .A1(new_n20195_), .B0(pi1153), .Y(new_n20198_));
  AND3X1   g17762(.A(new_n12439_), .B(pi0727), .C(pi0625), .Y(new_n20199_));
  NOR3X1   g17763(.A(new_n20199_), .B(new_n20193_), .C(new_n12364_), .Y(new_n20200_));
  NOR3X1   g17764(.A(new_n20200_), .B(new_n20198_), .C(pi0608), .Y(new_n20201_));
  AOI21X1  g17765(.A0(new_n12439_), .A1(pi0727), .B0(new_n20193_), .Y(new_n20202_));
  OAI21X1  g17766(.A0(new_n20202_), .A1(new_n20199_), .B0(new_n12364_), .Y(new_n20203_));
  NAND3X1  g17767(.A(new_n20197_), .B(new_n20194_), .C(pi1153), .Y(new_n20204_));
  AND3X1   g17768(.A(new_n20204_), .B(new_n20203_), .C(pi0608), .Y(new_n20205_));
  OR2X1    g17769(.A(new_n20205_), .B(new_n20201_), .Y(new_n20206_));
  MX2X1    g17770(.A(new_n20206_), .B(new_n20195_), .S0(new_n11769_), .Y(new_n20207_));
  OAI21X1  g17771(.A0(new_n2720_), .A1(new_n7872_), .B0(pi1153), .Y(new_n20208_));
  OAI21X1  g17772(.A0(new_n20208_), .A1(new_n20199_), .B0(new_n20203_), .Y(new_n20209_));
  MX2X1    g17773(.A(new_n20209_), .B(new_n20202_), .S0(new_n11769_), .Y(new_n20210_));
  OAI21X1  g17774(.A0(new_n20210_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n20211_));
  AOI21X1  g17775(.A0(new_n20207_), .A1(new_n12462_), .B0(new_n20211_), .Y(new_n20212_));
  AND3X1   g17776(.A(new_n12471_), .B(new_n12056_), .C(pi0772), .Y(new_n20213_));
  OAI21X1  g17777(.A0(new_n2720_), .A1(new_n7872_), .B0(pi1155), .Y(new_n20214_));
  OAI21X1  g17778(.A0(new_n20214_), .A1(new_n20213_), .B0(new_n12468_), .Y(new_n20215_));
  OAI21X1  g17779(.A0(new_n20210_), .A1(pi0609), .B0(pi1155), .Y(new_n20216_));
  AOI21X1  g17780(.A0(new_n20207_), .A1(pi0609), .B0(new_n20216_), .Y(new_n20217_));
  AND3X1   g17781(.A(new_n12480_), .B(new_n12056_), .C(pi0772), .Y(new_n20218_));
  OAI21X1  g17782(.A0(new_n2720_), .A1(new_n7872_), .B0(new_n12463_), .Y(new_n20219_));
  OAI21X1  g17783(.A0(new_n20219_), .A1(new_n20218_), .B0(pi0660), .Y(new_n20220_));
  OAI22X1  g17784(.A0(new_n20220_), .A1(new_n20217_), .B0(new_n20215_), .B1(new_n20212_), .Y(new_n20221_));
  MX2X1    g17785(.A(new_n20221_), .B(new_n20207_), .S0(new_n11768_), .Y(new_n20222_));
  NAND2X1  g17786(.A(new_n20222_), .B(pi0618), .Y(new_n20223_));
  OAI22X1  g17787(.A0(new_n20210_), .A1(new_n12490_), .B0(new_n2720_), .B1(new_n7872_), .Y(new_n20224_));
  AOI21X1  g17788(.A0(new_n20224_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20225_));
  OR3X1    g17789(.A(new_n14034_), .B(new_n12057_), .C(new_n15306_), .Y(new_n20226_));
  NOR3X1   g17790(.A(new_n20226_), .B(new_n12473_), .C(pi0618), .Y(new_n20227_));
  OAI21X1  g17791(.A0(new_n2720_), .A1(new_n7872_), .B0(new_n12487_), .Y(new_n20228_));
  OAI21X1  g17792(.A0(new_n20228_), .A1(new_n20227_), .B0(pi0627), .Y(new_n20229_));
  AOI21X1  g17793(.A0(new_n20225_), .A1(new_n20223_), .B0(new_n20229_), .Y(new_n20230_));
  NAND2X1  g17794(.A(new_n20222_), .B(new_n12486_), .Y(new_n20231_));
  AOI21X1  g17795(.A0(new_n20224_), .A1(pi0618), .B0(pi1154), .Y(new_n20232_));
  NOR3X1   g17796(.A(new_n20226_), .B(new_n12473_), .C(new_n12486_), .Y(new_n20233_));
  OAI21X1  g17797(.A0(new_n2720_), .A1(new_n7872_), .B0(pi1154), .Y(new_n20234_));
  OAI21X1  g17798(.A0(new_n20234_), .A1(new_n20233_), .B0(new_n12494_), .Y(new_n20235_));
  AOI21X1  g17799(.A0(new_n20232_), .A1(new_n20231_), .B0(new_n20235_), .Y(new_n20236_));
  OAI21X1  g17800(.A0(new_n20236_), .A1(new_n20230_), .B0(pi0781), .Y(new_n20237_));
  AOI21X1  g17801(.A0(new_n20222_), .A1(new_n11767_), .B0(new_n16118_), .Y(new_n20238_));
  OR3X1    g17802(.A(new_n20210_), .B(new_n12513_), .C(new_n12490_), .Y(new_n20239_));
  NOR4X1   g17803(.A(new_n20226_), .B(new_n14039_), .C(new_n12473_), .D(pi0619), .Y(new_n20240_));
  NOR4X1   g17804(.A(new_n20226_), .B(new_n14039_), .C(new_n12473_), .D(new_n12509_), .Y(new_n20241_));
  OAI22X1  g17805(.A0(new_n20241_), .A1(new_n16121_), .B0(new_n20240_), .B1(new_n16122_), .Y(new_n20242_));
  AOI21X1  g17806(.A0(new_n20239_), .A1(new_n16116_), .B0(new_n20242_), .Y(new_n20243_));
  OAI21X1  g17807(.A0(new_n2720_), .A1(new_n7872_), .B0(pi0789), .Y(new_n20244_));
  OAI21X1  g17808(.A0(new_n20244_), .A1(new_n20243_), .B0(new_n12709_), .Y(new_n20245_));
  AOI21X1  g17809(.A0(new_n20238_), .A1(new_n20237_), .B0(new_n20245_), .Y(new_n20246_));
  OAI22X1  g17810(.A0(new_n20239_), .A1(new_n12531_), .B0(new_n2720_), .B1(new_n7872_), .Y(new_n20247_));
  NOR4X1   g17811(.A(new_n14040_), .B(new_n14034_), .C(new_n12057_), .D(new_n15306_), .Y(new_n20248_));
  AOI21X1  g17812(.A0(new_n20248_), .A1(new_n12542_), .B0(new_n20193_), .Y(new_n20249_));
  OAI21X1  g17813(.A0(new_n20249_), .A1(pi1158), .B0(pi0641), .Y(new_n20250_));
  AOI21X1  g17814(.A0(new_n20247_), .A1(new_n14049_), .B0(new_n20250_), .Y(new_n20251_));
  AOI21X1  g17815(.A0(new_n20248_), .A1(pi0626), .B0(new_n20193_), .Y(new_n20252_));
  OAI21X1  g17816(.A0(new_n20252_), .A1(new_n12548_), .B0(new_n12543_), .Y(new_n20253_));
  AOI21X1  g17817(.A0(new_n20247_), .A1(new_n14061_), .B0(new_n20253_), .Y(new_n20254_));
  NOR3X1   g17818(.A(new_n20254_), .B(new_n20251_), .C(new_n11765_), .Y(new_n20255_));
  OR2X1    g17819(.A(new_n20255_), .B(new_n14125_), .Y(new_n20256_));
  AND3X1   g17820(.A(new_n20248_), .B(new_n16140_), .C(new_n12561_), .Y(new_n20257_));
  NOR2X1   g17821(.A(new_n20210_), .B(new_n13489_), .Y(new_n20258_));
  OAI22X1  g17822(.A0(new_n20258_), .A1(new_n12561_), .B0(new_n20257_), .B1(new_n12554_), .Y(new_n20259_));
  AOI21X1  g17823(.A0(new_n20248_), .A1(new_n16140_), .B0(pi0628), .Y(new_n20260_));
  OAI21X1  g17824(.A0(new_n20260_), .A1(new_n12561_), .B0(pi1156), .Y(new_n20261_));
  AOI21X1  g17825(.A0(new_n20258_), .A1(pi0628), .B0(new_n20261_), .Y(new_n20262_));
  AOI21X1  g17826(.A0(new_n20259_), .A1(new_n12555_), .B0(new_n20262_), .Y(new_n20263_));
  OAI21X1  g17827(.A0(new_n2720_), .A1(new_n7872_), .B0(pi0792), .Y(new_n20264_));
  OAI22X1  g17828(.A0(new_n20264_), .A1(new_n20263_), .B0(new_n20256_), .B1(new_n20246_), .Y(new_n20265_));
  NAND4X1  g17829(.A(new_n20248_), .B(new_n16140_), .C(new_n14327_), .D(new_n12592_), .Y(new_n20266_));
  NOR3X1   g17830(.A(new_n20210_), .B(new_n13508_), .C(new_n13489_), .Y(new_n20267_));
  INVX1    g17831(.A(new_n20267_), .Y(new_n20268_));
  AOI22X1  g17832(.A0(new_n20268_), .A1(pi0630), .B0(new_n20266_), .B1(pi0647), .Y(new_n20269_));
  AOI21X1  g17833(.A0(new_n20268_), .A1(new_n12592_), .B0(new_n12577_), .Y(new_n20270_));
  NAND4X1  g17834(.A(new_n20248_), .B(new_n16140_), .C(new_n14327_), .D(pi0630), .Y(new_n20271_));
  NAND2X1  g17835(.A(new_n20271_), .B(pi1157), .Y(new_n20272_));
  OAI22X1  g17836(.A0(new_n20272_), .A1(new_n20270_), .B0(new_n20269_), .B1(pi1157), .Y(new_n20273_));
  NOR2X1   g17837(.A(new_n20193_), .B(new_n11763_), .Y(new_n20274_));
  AOI22X1  g17838(.A0(new_n20274_), .A1(new_n20273_), .B0(new_n20265_), .B1(new_n14122_), .Y(new_n20275_));
  AOI21X1  g17839(.A0(new_n20267_), .A1(new_n14140_), .B0(new_n20193_), .Y(new_n20276_));
  OAI21X1  g17840(.A0(new_n20276_), .A1(pi0644), .B0(pi0715), .Y(new_n20277_));
  AOI21X1  g17841(.A0(new_n20275_), .A1(pi0644), .B0(new_n20277_), .Y(new_n20278_));
  NOR4X1   g17842(.A(new_n20226_), .B(new_n16164_), .C(new_n14040_), .D(new_n12708_), .Y(new_n20279_));
  OAI21X1  g17843(.A0(new_n2720_), .A1(new_n7872_), .B0(new_n12608_), .Y(new_n20280_));
  AOI21X1  g17844(.A0(new_n20279_), .A1(pi0644), .B0(new_n20280_), .Y(new_n20281_));
  NOR3X1   g17845(.A(new_n20281_), .B(new_n20278_), .C(new_n11762_), .Y(new_n20282_));
  OAI21X1  g17846(.A0(new_n20276_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n20283_));
  AOI21X1  g17847(.A0(new_n20275_), .A1(new_n12612_), .B0(new_n20283_), .Y(new_n20284_));
  OAI21X1  g17848(.A0(new_n2720_), .A1(new_n7872_), .B0(pi0715), .Y(new_n20285_));
  AOI21X1  g17849(.A0(new_n20279_), .A1(new_n12612_), .B0(new_n20285_), .Y(new_n20286_));
  NOR3X1   g17850(.A(new_n20286_), .B(new_n20284_), .C(pi1160), .Y(new_n20287_));
  OAI21X1  g17851(.A0(new_n20287_), .A1(new_n20282_), .B0(pi0790), .Y(new_n20288_));
  AOI21X1  g17852(.A0(new_n20275_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n20289_));
  AOI22X1  g17853(.A0(new_n20289_), .A1(new_n20288_), .B0(new_n20192_), .B1(new_n20191_), .Y(po0346));
  AOI21X1  g17854(.A0(pi1093), .A1(pi1092), .B0(pi0190), .Y(new_n20291_));
  INVX1    g17855(.A(new_n20291_), .Y(new_n20292_));
  AND2X1   g17856(.A(new_n12056_), .B(pi0763), .Y(new_n20293_));
  OAI21X1  g17857(.A0(new_n20293_), .A1(new_n20291_), .B0(new_n15771_), .Y(new_n20294_));
  AND3X1   g17858(.A(new_n12480_), .B(new_n12056_), .C(pi0763), .Y(new_n20295_));
  OAI21X1  g17859(.A0(new_n20295_), .A1(new_n20294_), .B0(pi1155), .Y(new_n20296_));
  NOR3X1   g17860(.A(new_n20295_), .B(new_n20291_), .C(pi1155), .Y(new_n20297_));
  INVX1    g17861(.A(new_n20297_), .Y(new_n20298_));
  AOI21X1  g17862(.A0(new_n20298_), .A1(new_n20296_), .B0(new_n11768_), .Y(new_n20299_));
  AOI21X1  g17863(.A0(new_n20294_), .A1(new_n11768_), .B0(new_n20299_), .Y(new_n20300_));
  AOI21X1  g17864(.A0(new_n20300_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n20301_));
  AOI21X1  g17865(.A0(new_n20300_), .A1(new_n12655_), .B0(pi1154), .Y(new_n20302_));
  NOR2X1   g17866(.A(new_n20302_), .B(new_n20301_), .Y(new_n20303_));
  MX2X1    g17867(.A(new_n20303_), .B(new_n20300_), .S0(new_n11767_), .Y(new_n20304_));
  NOR2X1   g17868(.A(new_n20304_), .B(pi0789), .Y(new_n20305_));
  AOI21X1  g17869(.A0(new_n20304_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n20306_));
  AOI21X1  g17870(.A0(new_n20304_), .A1(new_n15790_), .B0(pi1159), .Y(new_n20307_));
  OR2X1    g17871(.A(new_n20307_), .B(new_n20306_), .Y(new_n20308_));
  AOI21X1  g17872(.A0(new_n20308_), .A1(pi0789), .B0(new_n20305_), .Y(new_n20309_));
  INVX1    g17873(.A(new_n20309_), .Y(new_n20310_));
  MX2X1    g17874(.A(new_n20310_), .B(new_n20292_), .S0(new_n12708_), .Y(new_n20311_));
  MX2X1    g17875(.A(new_n20311_), .B(new_n20292_), .S0(new_n12580_), .Y(new_n20312_));
  AOI21X1  g17876(.A0(new_n12439_), .A1(pi0699), .B0(new_n20291_), .Y(new_n20313_));
  OR2X1    g17877(.A(new_n20313_), .B(pi0778), .Y(new_n20314_));
  INVX1    g17878(.A(new_n20313_), .Y(new_n20315_));
  AND3X1   g17879(.A(new_n12439_), .B(pi0699), .C(new_n12363_), .Y(new_n20316_));
  INVX1    g17880(.A(new_n20316_), .Y(new_n20317_));
  AOI21X1  g17881(.A0(new_n20317_), .A1(new_n20315_), .B0(new_n12364_), .Y(new_n20318_));
  NOR3X1   g17882(.A(new_n20316_), .B(new_n20291_), .C(pi1153), .Y(new_n20319_));
  OR3X1    g17883(.A(new_n20319_), .B(new_n20318_), .C(new_n11769_), .Y(new_n20320_));
  AND2X1   g17884(.A(new_n20320_), .B(new_n20314_), .Y(new_n20321_));
  NOR4X1   g17885(.A(new_n20321_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n20322_));
  AND3X1   g17886(.A(new_n20322_), .B(new_n12739_), .C(new_n12718_), .Y(new_n20323_));
  INVX1    g17887(.A(new_n20323_), .Y(new_n20324_));
  AOI21X1  g17888(.A0(new_n20291_), .A1(pi0647), .B0(pi1157), .Y(new_n20325_));
  OAI21X1  g17889(.A0(new_n20324_), .A1(pi0647), .B0(new_n20325_), .Y(new_n20326_));
  MX2X1    g17890(.A(new_n20323_), .B(new_n20291_), .S0(new_n12577_), .Y(new_n20327_));
  OAI22X1  g17891(.A0(new_n20327_), .A1(new_n14242_), .B0(new_n20326_), .B1(new_n12592_), .Y(new_n20328_));
  AOI21X1  g17892(.A0(new_n20312_), .A1(new_n14326_), .B0(new_n20328_), .Y(new_n20329_));
  OR2X1    g17893(.A(new_n20329_), .B(new_n11763_), .Y(new_n20330_));
  AOI21X1  g17894(.A0(new_n20292_), .A1(pi0626), .B0(new_n16218_), .Y(new_n20331_));
  OAI21X1  g17895(.A0(new_n20309_), .A1(pi0626), .B0(new_n20331_), .Y(new_n20332_));
  AOI21X1  g17896(.A0(new_n20292_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n20333_));
  OAI21X1  g17897(.A0(new_n20309_), .A1(new_n12542_), .B0(new_n20333_), .Y(new_n20334_));
  NAND2X1  g17898(.A(new_n20322_), .B(new_n12637_), .Y(new_n20335_));
  AND3X1   g17899(.A(new_n20335_), .B(new_n20334_), .C(new_n20332_), .Y(new_n20336_));
  NOR2X1   g17900(.A(new_n20336_), .B(new_n11765_), .Y(new_n20337_));
  NOR2X1   g17901(.A(new_n20291_), .B(pi1153), .Y(new_n20338_));
  NOR3X1   g17902(.A(new_n20313_), .B(new_n11991_), .C(new_n12363_), .Y(new_n20339_));
  AOI21X1  g17903(.A0(new_n12056_), .A1(pi0763), .B0(new_n20291_), .Y(new_n20340_));
  INVX1    g17904(.A(new_n20340_), .Y(new_n20341_));
  AOI21X1  g17905(.A0(new_n20315_), .A1(new_n12048_), .B0(new_n20341_), .Y(new_n20342_));
  OAI21X1  g17906(.A0(new_n20342_), .A1(new_n20339_), .B0(new_n20338_), .Y(new_n20343_));
  NOR2X1   g17907(.A(new_n20318_), .B(pi0608), .Y(new_n20344_));
  NOR3X1   g17908(.A(new_n20339_), .B(new_n20341_), .C(new_n12364_), .Y(new_n20345_));
  NOR3X1   g17909(.A(new_n20345_), .B(new_n20319_), .C(new_n12368_), .Y(new_n20346_));
  AOI21X1  g17910(.A0(new_n20344_), .A1(new_n20343_), .B0(new_n20346_), .Y(new_n20347_));
  OR2X1    g17911(.A(new_n20342_), .B(pi0778), .Y(new_n20348_));
  OAI21X1  g17912(.A0(new_n20347_), .A1(new_n11769_), .B0(new_n20348_), .Y(new_n20349_));
  INVX1    g17913(.A(new_n20349_), .Y(new_n20350_));
  AND2X1   g17914(.A(new_n20349_), .B(new_n12462_), .Y(new_n20351_));
  OAI21X1  g17915(.A0(new_n20321_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n20352_));
  OR2X1    g17916(.A(new_n20352_), .B(new_n20351_), .Y(new_n20353_));
  AND3X1   g17917(.A(new_n20353_), .B(new_n20296_), .C(new_n12468_), .Y(new_n20354_));
  OAI21X1  g17918(.A0(new_n20321_), .A1(pi0609), .B0(pi1155), .Y(new_n20355_));
  AOI21X1  g17919(.A0(new_n20349_), .A1(pi0609), .B0(new_n20355_), .Y(new_n20356_));
  NOR3X1   g17920(.A(new_n20356_), .B(new_n20297_), .C(new_n12468_), .Y(new_n20357_));
  NOR2X1   g17921(.A(new_n20357_), .B(new_n20354_), .Y(new_n20358_));
  MX2X1    g17922(.A(new_n20358_), .B(new_n20350_), .S0(new_n11768_), .Y(new_n20359_));
  AOI21X1  g17923(.A0(new_n20320_), .A1(new_n20314_), .B0(new_n12630_), .Y(new_n20360_));
  AOI21X1  g17924(.A0(new_n20360_), .A1(pi0618), .B0(pi1154), .Y(new_n20361_));
  OAI21X1  g17925(.A0(new_n20359_), .A1(pi0618), .B0(new_n20361_), .Y(new_n20362_));
  NOR2X1   g17926(.A(new_n20301_), .B(pi0627), .Y(new_n20363_));
  AOI21X1  g17927(.A0(new_n20360_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20364_));
  OAI21X1  g17928(.A0(new_n20359_), .A1(new_n12486_), .B0(new_n20364_), .Y(new_n20365_));
  NOR2X1   g17929(.A(new_n20302_), .B(new_n12494_), .Y(new_n20366_));
  AOI22X1  g17930(.A0(new_n20366_), .A1(new_n20365_), .B0(new_n20363_), .B1(new_n20362_), .Y(new_n20367_));
  MX2X1    g17931(.A(new_n20367_), .B(new_n20359_), .S0(new_n11767_), .Y(new_n20368_));
  OR4X1    g17932(.A(new_n20321_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n20369_));
  AND2X1   g17933(.A(new_n20369_), .B(new_n12510_), .Y(new_n20370_));
  OAI21X1  g17934(.A0(new_n20368_), .A1(pi0619), .B0(new_n20370_), .Y(new_n20371_));
  NOR2X1   g17935(.A(new_n20306_), .B(pi0648), .Y(new_n20372_));
  AND2X1   g17936(.A(new_n20372_), .B(new_n20371_), .Y(new_n20373_));
  NOR4X1   g17937(.A(new_n20321_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n20374_));
  NOR2X1   g17938(.A(new_n20374_), .B(new_n12510_), .Y(new_n20375_));
  OAI21X1  g17939(.A0(new_n20368_), .A1(new_n12509_), .B0(new_n20375_), .Y(new_n20376_));
  NOR2X1   g17940(.A(new_n20307_), .B(new_n12517_), .Y(new_n20377_));
  AND2X1   g17941(.A(new_n20377_), .B(new_n20376_), .Y(new_n20378_));
  OR3X1    g17942(.A(new_n20378_), .B(new_n20373_), .C(new_n11766_), .Y(new_n20379_));
  AOI21X1  g17943(.A0(new_n20368_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n20380_));
  AOI21X1  g17944(.A0(new_n20380_), .A1(new_n20379_), .B0(new_n20337_), .Y(new_n20381_));
  INVX1    g17945(.A(new_n20311_), .Y(new_n20382_));
  AND2X1   g17946(.A(new_n20322_), .B(new_n12718_), .Y(new_n20383_));
  AOI22X1  g17947(.A0(new_n20383_), .A1(new_n14426_), .B0(new_n20382_), .B1(new_n12735_), .Y(new_n20384_));
  AOI22X1  g17948(.A0(new_n20383_), .A1(new_n14428_), .B0(new_n20382_), .B1(new_n12733_), .Y(new_n20385_));
  MX2X1    g17949(.A(new_n20385_), .B(new_n20384_), .S0(new_n12561_), .Y(new_n20386_));
  OAI21X1  g17950(.A0(new_n20386_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n20387_));
  INVX1    g17951(.A(new_n20387_), .Y(new_n20388_));
  OAI21X1  g17952(.A0(new_n20381_), .A1(new_n14125_), .B0(new_n20388_), .Y(new_n20389_));
  AND2X1   g17953(.A(new_n20389_), .B(new_n20330_), .Y(new_n20390_));
  OAI21X1  g17954(.A0(new_n20327_), .A1(new_n12578_), .B0(new_n20326_), .Y(new_n20391_));
  MX2X1    g17955(.A(new_n20391_), .B(new_n20324_), .S0(new_n11763_), .Y(new_n20392_));
  OAI21X1  g17956(.A0(new_n20392_), .A1(pi0644), .B0(pi0715), .Y(new_n20393_));
  AOI21X1  g17957(.A0(new_n20390_), .A1(pi0644), .B0(new_n20393_), .Y(new_n20394_));
  OR3X1    g17958(.A(new_n20292_), .B(new_n12603_), .C(new_n11763_), .Y(new_n20395_));
  OAI21X1  g17959(.A0(new_n20312_), .A1(new_n12604_), .B0(new_n20395_), .Y(new_n20396_));
  OAI21X1  g17960(.A0(new_n20292_), .A1(pi0644), .B0(new_n12608_), .Y(new_n20397_));
  AOI21X1  g17961(.A0(new_n20396_), .A1(pi0644), .B0(new_n20397_), .Y(new_n20398_));
  OR2X1    g17962(.A(new_n20398_), .B(new_n11762_), .Y(new_n20399_));
  OAI21X1  g17963(.A0(new_n20392_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n20400_));
  AOI21X1  g17964(.A0(new_n20390_), .A1(new_n12612_), .B0(new_n20400_), .Y(new_n20401_));
  OAI21X1  g17965(.A0(new_n20292_), .A1(new_n12612_), .B0(pi0715), .Y(new_n20402_));
  AOI21X1  g17966(.A0(new_n20396_), .A1(new_n12612_), .B0(new_n20402_), .Y(new_n20403_));
  OR2X1    g17967(.A(new_n20403_), .B(pi1160), .Y(new_n20404_));
  OAI22X1  g17968(.A0(new_n20404_), .A1(new_n20401_), .B0(new_n20399_), .B1(new_n20394_), .Y(new_n20405_));
  NAND2X1  g17969(.A(new_n20405_), .B(pi0790), .Y(new_n20406_));
  AOI21X1  g17970(.A0(new_n20390_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n20407_));
  AOI21X1  g17971(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0190), .Y(new_n20408_));
  INVX1    g17972(.A(new_n20408_), .Y(new_n20409_));
  OAI21X1  g17973(.A0(new_n12826_), .A1(new_n9900_), .B0(new_n2979_), .Y(new_n20410_));
  AOI21X1  g17974(.A0(new_n12825_), .A1(new_n9900_), .B0(new_n20410_), .Y(new_n20411_));
  AOI21X1  g17975(.A0(new_n12771_), .A1(new_n9900_), .B0(new_n12441_), .Y(new_n20412_));
  NOR3X1   g17976(.A(new_n20412_), .B(new_n20411_), .C(new_n15361_), .Y(new_n20413_));
  OR2X1    g17977(.A(pi0699), .B(pi0190), .Y(new_n20414_));
  OAI21X1  g17978(.A0(new_n20414_), .A1(new_n12447_), .B0(new_n3103_), .Y(new_n20415_));
  OAI22X1  g17979(.A0(new_n20415_), .A1(new_n20413_), .B0(new_n3103_), .B1(new_n9900_), .Y(new_n20416_));
  AND2X1   g17980(.A(new_n20416_), .B(new_n11769_), .Y(new_n20417_));
  AOI21X1  g17981(.A0(new_n20408_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n20418_));
  OAI21X1  g17982(.A0(new_n20416_), .A1(new_n12363_), .B0(new_n20418_), .Y(new_n20419_));
  AOI21X1  g17983(.A0(new_n20408_), .A1(pi0625), .B0(pi1153), .Y(new_n20420_));
  OAI21X1  g17984(.A0(new_n20416_), .A1(pi0625), .B0(new_n20420_), .Y(new_n20421_));
  AOI21X1  g17985(.A0(new_n20421_), .A1(new_n20419_), .B0(new_n11769_), .Y(new_n20422_));
  NOR2X1   g17986(.A(new_n20422_), .B(new_n20417_), .Y(new_n20423_));
  MX2X1    g17987(.A(new_n20423_), .B(new_n20408_), .S0(new_n12490_), .Y(new_n20424_));
  AND2X1   g17988(.A(new_n20408_), .B(new_n12513_), .Y(new_n20425_));
  AOI21X1  g17989(.A0(new_n20424_), .A1(new_n14053_), .B0(new_n20425_), .Y(new_n20426_));
  MX2X1    g17990(.A(new_n20426_), .B(new_n20409_), .S0(new_n12531_), .Y(new_n20427_));
  MX2X1    g17991(.A(new_n20427_), .B(new_n20409_), .S0(new_n12563_), .Y(new_n20428_));
  MX2X1    g17992(.A(new_n20428_), .B(new_n20409_), .S0(pi0628), .Y(new_n20429_));
  MX2X1    g17993(.A(new_n20428_), .B(new_n20409_), .S0(new_n12554_), .Y(new_n20430_));
  MX2X1    g17994(.A(new_n20430_), .B(new_n20429_), .S0(new_n12555_), .Y(new_n20431_));
  MX2X1    g17995(.A(new_n20431_), .B(new_n20428_), .S0(new_n11764_), .Y(new_n20432_));
  MX2X1    g17996(.A(new_n20432_), .B(new_n20409_), .S0(pi0647), .Y(new_n20433_));
  MX2X1    g17997(.A(new_n20432_), .B(new_n20409_), .S0(new_n12577_), .Y(new_n20434_));
  MX2X1    g17998(.A(new_n20434_), .B(new_n20433_), .S0(new_n12578_), .Y(new_n20435_));
  MX2X1    g17999(.A(new_n20435_), .B(new_n20432_), .S0(new_n11763_), .Y(new_n20436_));
  OAI21X1  g18000(.A0(new_n20436_), .A1(pi0644), .B0(pi0715), .Y(new_n20437_));
  AOI22X1  g18001(.A0(new_n12073_), .A1(pi0190), .B0(new_n12444_), .B1(new_n15365_), .Y(new_n20438_));
  OR3X1    g18002(.A(new_n12776_), .B(new_n15365_), .C(pi0190), .Y(new_n20439_));
  OAI21X1  g18003(.A0(new_n12045_), .A1(pi0039), .B0(pi0763), .Y(new_n20440_));
  AOI21X1  g18004(.A0(new_n20440_), .A1(pi0190), .B0(new_n15366_), .Y(new_n20441_));
  AND2X1   g18005(.A(new_n20441_), .B(new_n20439_), .Y(new_n20442_));
  OAI21X1  g18006(.A0(new_n20438_), .A1(new_n2939_), .B0(new_n20442_), .Y(new_n20443_));
  OAI21X1  g18007(.A0(new_n12077_), .A1(pi0190), .B0(pi0038), .Y(new_n20444_));
  AOI21X1  g18008(.A0(new_n12079_), .A1(pi0763), .B0(new_n20444_), .Y(new_n20445_));
  AOI21X1  g18009(.A0(new_n20443_), .A1(new_n2979_), .B0(new_n20445_), .Y(new_n20446_));
  MX2X1    g18010(.A(new_n20446_), .B(new_n9900_), .S0(new_n11770_), .Y(new_n20447_));
  MX2X1    g18011(.A(new_n20447_), .B(new_n20408_), .S0(new_n12473_), .Y(new_n20448_));
  NOR2X1   g18012(.A(new_n20447_), .B(new_n12473_), .Y(new_n20449_));
  AOI22X1  g18013(.A0(new_n20449_), .A1(pi0609), .B0(new_n20409_), .B1(new_n12472_), .Y(new_n20450_));
  AOI22X1  g18014(.A0(new_n20449_), .A1(new_n12462_), .B0(new_n20409_), .B1(new_n12481_), .Y(new_n20451_));
  MX2X1    g18015(.A(new_n20451_), .B(new_n20450_), .S0(pi1155), .Y(new_n20452_));
  MX2X1    g18016(.A(new_n20452_), .B(new_n20448_), .S0(new_n11768_), .Y(new_n20453_));
  OAI21X1  g18017(.A0(new_n20409_), .A1(pi0618), .B0(pi1154), .Y(new_n20454_));
  AOI21X1  g18018(.A0(new_n20453_), .A1(pi0618), .B0(new_n20454_), .Y(new_n20455_));
  OAI21X1  g18019(.A0(new_n20409_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20456_));
  AOI21X1  g18020(.A0(new_n20453_), .A1(new_n12486_), .B0(new_n20456_), .Y(new_n20457_));
  NOR2X1   g18021(.A(new_n20457_), .B(new_n20455_), .Y(new_n20458_));
  MX2X1    g18022(.A(new_n20458_), .B(new_n20453_), .S0(new_n11767_), .Y(new_n20459_));
  OAI21X1  g18023(.A0(new_n20409_), .A1(pi0619), .B0(pi1159), .Y(new_n20460_));
  AOI21X1  g18024(.A0(new_n20459_), .A1(pi0619), .B0(new_n20460_), .Y(new_n20461_));
  OAI21X1  g18025(.A0(new_n20409_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n20462_));
  AOI21X1  g18026(.A0(new_n20459_), .A1(new_n12509_), .B0(new_n20462_), .Y(new_n20463_));
  NOR2X1   g18027(.A(new_n20463_), .B(new_n20461_), .Y(new_n20464_));
  MX2X1    g18028(.A(new_n20464_), .B(new_n20459_), .S0(new_n11766_), .Y(new_n20465_));
  AND2X1   g18029(.A(new_n20408_), .B(new_n12708_), .Y(new_n20466_));
  AOI21X1  g18030(.A0(new_n20465_), .A1(new_n16140_), .B0(new_n20466_), .Y(new_n20467_));
  MX2X1    g18031(.A(new_n20467_), .B(new_n20409_), .S0(new_n12580_), .Y(new_n20468_));
  MX2X1    g18032(.A(new_n20468_), .B(new_n20409_), .S0(new_n12604_), .Y(new_n20469_));
  AOI21X1  g18033(.A0(new_n20408_), .A1(new_n12612_), .B0(pi0715), .Y(new_n20470_));
  OAI21X1  g18034(.A0(new_n20469_), .A1(new_n12612_), .B0(new_n20470_), .Y(new_n20471_));
  NAND3X1  g18035(.A(new_n20471_), .B(new_n20437_), .C(pi1160), .Y(new_n20472_));
  OAI21X1  g18036(.A0(new_n20436_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n20473_));
  AOI21X1  g18037(.A0(new_n20408_), .A1(pi0644), .B0(new_n12608_), .Y(new_n20474_));
  OAI21X1  g18038(.A0(new_n20469_), .A1(pi0644), .B0(new_n20474_), .Y(new_n20475_));
  NAND3X1  g18039(.A(new_n20475_), .B(new_n20473_), .C(new_n11762_), .Y(new_n20476_));
  AND2X1   g18040(.A(new_n20476_), .B(new_n20472_), .Y(new_n20477_));
  NAND3X1  g18041(.A(new_n20475_), .B(new_n11762_), .C(new_n12612_), .Y(new_n20478_));
  NAND3X1  g18042(.A(new_n20471_), .B(pi1160), .C(pi0644), .Y(new_n20479_));
  AND3X1   g18043(.A(new_n20479_), .B(new_n20478_), .C(pi0790), .Y(new_n20480_));
  NAND2X1  g18044(.A(new_n20467_), .B(new_n14249_), .Y(new_n20481_));
  AOI22X1  g18045(.A0(new_n20430_), .A1(new_n16373_), .B0(new_n20429_), .B1(new_n16374_), .Y(new_n20482_));
  AOI21X1  g18046(.A0(new_n20482_), .A1(new_n20481_), .B0(new_n11764_), .Y(new_n20483_));
  AND2X1   g18047(.A(new_n20446_), .B(new_n15361_), .Y(new_n20484_));
  INVX1    g18048(.A(new_n20484_), .Y(new_n20485_));
  AOI21X1  g18049(.A0(new_n16381_), .A1(pi0190), .B0(pi0763), .Y(new_n20486_));
  OAI21X1  g18050(.A0(new_n16380_), .A1(pi0190), .B0(new_n20486_), .Y(new_n20487_));
  AOI21X1  g18051(.A0(new_n12788_), .A1(new_n9900_), .B0(new_n15365_), .Y(new_n20488_));
  OAI21X1  g18052(.A0(new_n12787_), .A1(new_n9900_), .B0(new_n20488_), .Y(new_n20489_));
  AND2X1   g18053(.A(new_n20489_), .B(pi0039), .Y(new_n20490_));
  AND2X1   g18054(.A(new_n20490_), .B(new_n20487_), .Y(new_n20491_));
  AOI21X1  g18055(.A0(new_n12795_), .A1(pi0190), .B0(pi0763), .Y(new_n20492_));
  OAI21X1  g18056(.A0(new_n12792_), .A1(pi0190), .B0(new_n20492_), .Y(new_n20493_));
  NOR2X1   g18057(.A(new_n12798_), .B(pi0190), .Y(new_n20494_));
  INVX1    g18058(.A(new_n20494_), .Y(new_n20495_));
  AOI21X1  g18059(.A0(new_n12800_), .A1(pi0190), .B0(new_n15365_), .Y(new_n20496_));
  AOI21X1  g18060(.A0(new_n20496_), .A1(new_n20495_), .B0(pi0039), .Y(new_n20497_));
  AOI21X1  g18061(.A0(new_n20497_), .A1(new_n20493_), .B0(pi0038), .Y(new_n20498_));
  INVX1    g18062(.A(new_n20498_), .Y(new_n20499_));
  AOI21X1  g18063(.A0(new_n16396_), .A1(new_n15365_), .B0(new_n12276_), .Y(new_n20500_));
  OAI21X1  g18064(.A0(new_n20500_), .A1(pi0039), .B0(new_n9900_), .Y(new_n20501_));
  OAI21X1  g18065(.A0(new_n20293_), .A1(new_n13443_), .B0(pi0190), .Y(new_n20502_));
  OAI21X1  g18066(.A0(new_n20502_), .A1(new_n16399_), .B0(pi0038), .Y(new_n20503_));
  INVX1    g18067(.A(new_n20503_), .Y(new_n20504_));
  AOI21X1  g18068(.A0(new_n20504_), .A1(new_n20501_), .B0(new_n15361_), .Y(new_n20505_));
  OAI21X1  g18069(.A0(new_n20499_), .A1(new_n20491_), .B0(new_n20505_), .Y(new_n20506_));
  AND2X1   g18070(.A(new_n20506_), .B(new_n3103_), .Y(new_n20507_));
  AOI22X1  g18071(.A0(new_n20507_), .A1(new_n20485_), .B0(new_n11770_), .B1(pi0190), .Y(new_n20508_));
  INVX1    g18072(.A(new_n20508_), .Y(new_n20509_));
  AOI21X1  g18073(.A0(new_n20447_), .A1(pi0625), .B0(pi1153), .Y(new_n20510_));
  OAI21X1  g18074(.A0(new_n20509_), .A1(pi0625), .B0(new_n20510_), .Y(new_n20511_));
  AND2X1   g18075(.A(new_n20419_), .B(new_n12368_), .Y(new_n20512_));
  AOI21X1  g18076(.A0(new_n20447_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n20513_));
  OAI21X1  g18077(.A0(new_n20509_), .A1(new_n12363_), .B0(new_n20513_), .Y(new_n20514_));
  AND2X1   g18078(.A(new_n20421_), .B(pi0608), .Y(new_n20515_));
  AOI22X1  g18079(.A0(new_n20515_), .A1(new_n20514_), .B0(new_n20512_), .B1(new_n20511_), .Y(new_n20516_));
  MX2X1    g18080(.A(new_n20516_), .B(new_n20509_), .S0(new_n11769_), .Y(new_n20517_));
  AOI21X1  g18081(.A0(new_n20423_), .A1(pi0609), .B0(pi1155), .Y(new_n20518_));
  OAI21X1  g18082(.A0(new_n20517_), .A1(pi0609), .B0(new_n20518_), .Y(new_n20519_));
  OAI21X1  g18083(.A0(new_n20450_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n20520_));
  INVX1    g18084(.A(new_n20520_), .Y(new_n20521_));
  AOI21X1  g18085(.A0(new_n20423_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n20522_));
  OAI21X1  g18086(.A0(new_n20517_), .A1(new_n12462_), .B0(new_n20522_), .Y(new_n20523_));
  OAI21X1  g18087(.A0(new_n20451_), .A1(pi1155), .B0(pi0660), .Y(new_n20524_));
  INVX1    g18088(.A(new_n20524_), .Y(new_n20525_));
  AOI22X1  g18089(.A0(new_n20525_), .A1(new_n20523_), .B0(new_n20521_), .B1(new_n20519_), .Y(new_n20526_));
  MX2X1    g18090(.A(new_n20526_), .B(new_n20517_), .S0(new_n11768_), .Y(new_n20527_));
  AOI21X1  g18091(.A0(new_n20424_), .A1(pi0618), .B0(pi1154), .Y(new_n20528_));
  OAI21X1  g18092(.A0(new_n20527_), .A1(pi0618), .B0(new_n20528_), .Y(new_n20529_));
  NOR2X1   g18093(.A(new_n20455_), .B(pi0627), .Y(new_n20530_));
  AOI21X1  g18094(.A0(new_n20424_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20531_));
  OAI21X1  g18095(.A0(new_n20527_), .A1(new_n12486_), .B0(new_n20531_), .Y(new_n20532_));
  NOR2X1   g18096(.A(new_n20457_), .B(new_n12494_), .Y(new_n20533_));
  AOI22X1  g18097(.A0(new_n20533_), .A1(new_n20532_), .B0(new_n20530_), .B1(new_n20529_), .Y(new_n20534_));
  MX2X1    g18098(.A(new_n20534_), .B(new_n20527_), .S0(new_n11767_), .Y(new_n20535_));
  INVX1    g18099(.A(new_n20535_), .Y(new_n20536_));
  OAI21X1  g18100(.A0(new_n20426_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n20537_));
  AOI21X1  g18101(.A0(new_n20536_), .A1(new_n12509_), .B0(new_n20537_), .Y(new_n20538_));
  NOR3X1   g18102(.A(new_n20538_), .B(new_n20461_), .C(pi0648), .Y(new_n20539_));
  OAI21X1  g18103(.A0(new_n20426_), .A1(pi0619), .B0(pi1159), .Y(new_n20540_));
  AOI21X1  g18104(.A0(new_n20536_), .A1(pi0619), .B0(new_n20540_), .Y(new_n20541_));
  OR2X1    g18105(.A(new_n20463_), .B(new_n12517_), .Y(new_n20542_));
  OAI21X1  g18106(.A0(new_n20542_), .A1(new_n20541_), .B0(pi0789), .Y(new_n20543_));
  AOI21X1  g18107(.A0(new_n20535_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n20544_));
  OAI21X1  g18108(.A0(new_n20543_), .A1(new_n20539_), .B0(new_n20544_), .Y(new_n20545_));
  AOI21X1  g18109(.A0(new_n20409_), .A1(pi0626), .B0(new_n16218_), .Y(new_n20546_));
  OAI21X1  g18110(.A0(new_n20465_), .A1(pi0626), .B0(new_n20546_), .Y(new_n20547_));
  AOI21X1  g18111(.A0(new_n20409_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n20548_));
  OAI21X1  g18112(.A0(new_n20465_), .A1(new_n12542_), .B0(new_n20548_), .Y(new_n20549_));
  OR2X1    g18113(.A(new_n20427_), .B(new_n13439_), .Y(new_n20550_));
  NAND3X1  g18114(.A(new_n20550_), .B(new_n20549_), .C(new_n20547_), .Y(new_n20551_));
  AOI21X1  g18115(.A0(new_n20551_), .A1(pi0788), .B0(new_n14125_), .Y(new_n20552_));
  AOI21X1  g18116(.A0(new_n20552_), .A1(new_n20545_), .B0(new_n20483_), .Y(new_n20553_));
  AND2X1   g18117(.A(new_n20468_), .B(new_n14326_), .Y(new_n20554_));
  AND2X1   g18118(.A(new_n20434_), .B(new_n14241_), .Y(new_n20555_));
  AND2X1   g18119(.A(new_n20433_), .B(new_n14243_), .Y(new_n20556_));
  OR2X1    g18120(.A(new_n20556_), .B(new_n20555_), .Y(new_n20557_));
  OAI21X1  g18121(.A0(new_n20557_), .A1(new_n20554_), .B0(pi0787), .Y(new_n20558_));
  OAI21X1  g18122(.A0(new_n20553_), .A1(new_n14121_), .B0(new_n20558_), .Y(new_n20559_));
  OAI22X1  g18123(.A0(new_n20559_), .A1(new_n20480_), .B0(new_n20477_), .B1(new_n12766_), .Y(new_n20560_));
  OAI21X1  g18124(.A0(new_n6489_), .A1(pi0190), .B0(new_n12767_), .Y(new_n20561_));
  AOI21X1  g18125(.A0(new_n20560_), .A1(new_n6489_), .B0(new_n20561_), .Y(new_n20562_));
  AOI21X1  g18126(.A0(new_n20407_), .A1(new_n20406_), .B0(new_n20562_), .Y(po0347));
  AOI21X1  g18127(.A0(pi1093), .A1(pi1092), .B0(pi0191), .Y(new_n20564_));
  INVX1    g18128(.A(new_n20564_), .Y(new_n20565_));
  AND2X1   g18129(.A(new_n12056_), .B(pi0746), .Y(new_n20566_));
  OAI21X1  g18130(.A0(new_n20566_), .A1(new_n20564_), .B0(new_n15771_), .Y(new_n20567_));
  AND3X1   g18131(.A(new_n12480_), .B(new_n12056_), .C(pi0746), .Y(new_n20568_));
  OAI21X1  g18132(.A0(new_n20568_), .A1(new_n20567_), .B0(pi1155), .Y(new_n20569_));
  NOR3X1   g18133(.A(new_n20568_), .B(new_n20564_), .C(pi1155), .Y(new_n20570_));
  INVX1    g18134(.A(new_n20570_), .Y(new_n20571_));
  AOI21X1  g18135(.A0(new_n20571_), .A1(new_n20569_), .B0(new_n11768_), .Y(new_n20572_));
  AOI21X1  g18136(.A0(new_n20567_), .A1(new_n11768_), .B0(new_n20572_), .Y(new_n20573_));
  AOI21X1  g18137(.A0(new_n20573_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n20574_));
  AOI21X1  g18138(.A0(new_n20573_), .A1(new_n12655_), .B0(pi1154), .Y(new_n20575_));
  NOR2X1   g18139(.A(new_n20575_), .B(new_n20574_), .Y(new_n20576_));
  MX2X1    g18140(.A(new_n20576_), .B(new_n20573_), .S0(new_n11767_), .Y(new_n20577_));
  NOR2X1   g18141(.A(new_n20577_), .B(pi0789), .Y(new_n20578_));
  AOI21X1  g18142(.A0(new_n20577_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n20579_));
  AOI21X1  g18143(.A0(new_n20577_), .A1(new_n15790_), .B0(pi1159), .Y(new_n20580_));
  OR2X1    g18144(.A(new_n20580_), .B(new_n20579_), .Y(new_n20581_));
  AOI21X1  g18145(.A0(new_n20581_), .A1(pi0789), .B0(new_n20578_), .Y(new_n20582_));
  INVX1    g18146(.A(new_n20582_), .Y(new_n20583_));
  MX2X1    g18147(.A(new_n20583_), .B(new_n20565_), .S0(new_n12708_), .Y(new_n20584_));
  MX2X1    g18148(.A(new_n20584_), .B(new_n20565_), .S0(new_n12580_), .Y(new_n20585_));
  AOI21X1  g18149(.A0(new_n12439_), .A1(pi0729), .B0(new_n20564_), .Y(new_n20586_));
  OR2X1    g18150(.A(new_n20586_), .B(pi0778), .Y(new_n20587_));
  INVX1    g18151(.A(new_n20586_), .Y(new_n20588_));
  AND3X1   g18152(.A(new_n12439_), .B(pi0729), .C(new_n12363_), .Y(new_n20589_));
  INVX1    g18153(.A(new_n20589_), .Y(new_n20590_));
  AOI21X1  g18154(.A0(new_n20590_), .A1(new_n20588_), .B0(new_n12364_), .Y(new_n20591_));
  NOR3X1   g18155(.A(new_n20589_), .B(new_n20564_), .C(pi1153), .Y(new_n20592_));
  OR3X1    g18156(.A(new_n20592_), .B(new_n20591_), .C(new_n11769_), .Y(new_n20593_));
  AND2X1   g18157(.A(new_n20593_), .B(new_n20587_), .Y(new_n20594_));
  NOR4X1   g18158(.A(new_n20594_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n20595_));
  AND3X1   g18159(.A(new_n20595_), .B(new_n12739_), .C(new_n12718_), .Y(new_n20596_));
  INVX1    g18160(.A(new_n20596_), .Y(new_n20597_));
  AOI21X1  g18161(.A0(new_n20564_), .A1(pi0647), .B0(pi1157), .Y(new_n20598_));
  OAI21X1  g18162(.A0(new_n20597_), .A1(pi0647), .B0(new_n20598_), .Y(new_n20599_));
  MX2X1    g18163(.A(new_n20596_), .B(new_n20564_), .S0(new_n12577_), .Y(new_n20600_));
  OAI22X1  g18164(.A0(new_n20600_), .A1(new_n14242_), .B0(new_n20599_), .B1(new_n12592_), .Y(new_n20601_));
  AOI21X1  g18165(.A0(new_n20585_), .A1(new_n14326_), .B0(new_n20601_), .Y(new_n20602_));
  OR2X1    g18166(.A(new_n20602_), .B(new_n11763_), .Y(new_n20603_));
  AOI21X1  g18167(.A0(new_n20565_), .A1(pi0626), .B0(new_n16218_), .Y(new_n20604_));
  OAI21X1  g18168(.A0(new_n20582_), .A1(pi0626), .B0(new_n20604_), .Y(new_n20605_));
  AOI21X1  g18169(.A0(new_n20565_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n20606_));
  OAI21X1  g18170(.A0(new_n20582_), .A1(new_n12542_), .B0(new_n20606_), .Y(new_n20607_));
  NAND2X1  g18171(.A(new_n20595_), .B(new_n12637_), .Y(new_n20608_));
  AND3X1   g18172(.A(new_n20608_), .B(new_n20607_), .C(new_n20605_), .Y(new_n20609_));
  NOR2X1   g18173(.A(new_n20609_), .B(new_n11765_), .Y(new_n20610_));
  NOR2X1   g18174(.A(new_n20564_), .B(pi1153), .Y(new_n20611_));
  NOR3X1   g18175(.A(new_n20586_), .B(new_n11991_), .C(new_n12363_), .Y(new_n20612_));
  AOI21X1  g18176(.A0(new_n12056_), .A1(pi0746), .B0(new_n20564_), .Y(new_n20613_));
  INVX1    g18177(.A(new_n20613_), .Y(new_n20614_));
  AOI21X1  g18178(.A0(new_n20588_), .A1(new_n12048_), .B0(new_n20614_), .Y(new_n20615_));
  OAI21X1  g18179(.A0(new_n20615_), .A1(new_n20612_), .B0(new_n20611_), .Y(new_n20616_));
  NOR2X1   g18180(.A(new_n20591_), .B(pi0608), .Y(new_n20617_));
  NOR3X1   g18181(.A(new_n20612_), .B(new_n20614_), .C(new_n12364_), .Y(new_n20618_));
  NOR3X1   g18182(.A(new_n20618_), .B(new_n20592_), .C(new_n12368_), .Y(new_n20619_));
  AOI21X1  g18183(.A0(new_n20617_), .A1(new_n20616_), .B0(new_n20619_), .Y(new_n20620_));
  OR2X1    g18184(.A(new_n20615_), .B(pi0778), .Y(new_n20621_));
  OAI21X1  g18185(.A0(new_n20620_), .A1(new_n11769_), .B0(new_n20621_), .Y(new_n20622_));
  INVX1    g18186(.A(new_n20622_), .Y(new_n20623_));
  AND2X1   g18187(.A(new_n20622_), .B(new_n12462_), .Y(new_n20624_));
  OAI21X1  g18188(.A0(new_n20594_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n20625_));
  OR2X1    g18189(.A(new_n20625_), .B(new_n20624_), .Y(new_n20626_));
  AND3X1   g18190(.A(new_n20626_), .B(new_n20569_), .C(new_n12468_), .Y(new_n20627_));
  OAI21X1  g18191(.A0(new_n20594_), .A1(pi0609), .B0(pi1155), .Y(new_n20628_));
  AOI21X1  g18192(.A0(new_n20622_), .A1(pi0609), .B0(new_n20628_), .Y(new_n20629_));
  NOR3X1   g18193(.A(new_n20629_), .B(new_n20570_), .C(new_n12468_), .Y(new_n20630_));
  NOR2X1   g18194(.A(new_n20630_), .B(new_n20627_), .Y(new_n20631_));
  MX2X1    g18195(.A(new_n20631_), .B(new_n20623_), .S0(new_n11768_), .Y(new_n20632_));
  AOI21X1  g18196(.A0(new_n20593_), .A1(new_n20587_), .B0(new_n12630_), .Y(new_n20633_));
  AOI21X1  g18197(.A0(new_n20633_), .A1(pi0618), .B0(pi1154), .Y(new_n20634_));
  OAI21X1  g18198(.A0(new_n20632_), .A1(pi0618), .B0(new_n20634_), .Y(new_n20635_));
  NOR2X1   g18199(.A(new_n20574_), .B(pi0627), .Y(new_n20636_));
  AOI21X1  g18200(.A0(new_n20633_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20637_));
  OAI21X1  g18201(.A0(new_n20632_), .A1(new_n12486_), .B0(new_n20637_), .Y(new_n20638_));
  NOR2X1   g18202(.A(new_n20575_), .B(new_n12494_), .Y(new_n20639_));
  AOI22X1  g18203(.A0(new_n20639_), .A1(new_n20638_), .B0(new_n20636_), .B1(new_n20635_), .Y(new_n20640_));
  MX2X1    g18204(.A(new_n20640_), .B(new_n20632_), .S0(new_n11767_), .Y(new_n20641_));
  OR4X1    g18205(.A(new_n20594_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n20642_));
  AND2X1   g18206(.A(new_n20642_), .B(new_n12510_), .Y(new_n20643_));
  OAI21X1  g18207(.A0(new_n20641_), .A1(pi0619), .B0(new_n20643_), .Y(new_n20644_));
  NOR2X1   g18208(.A(new_n20579_), .B(pi0648), .Y(new_n20645_));
  AND2X1   g18209(.A(new_n20645_), .B(new_n20644_), .Y(new_n20646_));
  NOR4X1   g18210(.A(new_n20594_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n20647_));
  NOR2X1   g18211(.A(new_n20647_), .B(new_n12510_), .Y(new_n20648_));
  OAI21X1  g18212(.A0(new_n20641_), .A1(new_n12509_), .B0(new_n20648_), .Y(new_n20649_));
  NOR2X1   g18213(.A(new_n20580_), .B(new_n12517_), .Y(new_n20650_));
  AND2X1   g18214(.A(new_n20650_), .B(new_n20649_), .Y(new_n20651_));
  OR3X1    g18215(.A(new_n20651_), .B(new_n20646_), .C(new_n11766_), .Y(new_n20652_));
  AOI21X1  g18216(.A0(new_n20641_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n20653_));
  AOI21X1  g18217(.A0(new_n20653_), .A1(new_n20652_), .B0(new_n20610_), .Y(new_n20654_));
  INVX1    g18218(.A(new_n20584_), .Y(new_n20655_));
  AND2X1   g18219(.A(new_n20595_), .B(new_n12718_), .Y(new_n20656_));
  AOI22X1  g18220(.A0(new_n20656_), .A1(new_n14426_), .B0(new_n20655_), .B1(new_n12735_), .Y(new_n20657_));
  AOI22X1  g18221(.A0(new_n20656_), .A1(new_n14428_), .B0(new_n20655_), .B1(new_n12733_), .Y(new_n20658_));
  MX2X1    g18222(.A(new_n20658_), .B(new_n20657_), .S0(new_n12561_), .Y(new_n20659_));
  OAI21X1  g18223(.A0(new_n20659_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n20660_));
  INVX1    g18224(.A(new_n20660_), .Y(new_n20661_));
  OAI21X1  g18225(.A0(new_n20654_), .A1(new_n14125_), .B0(new_n20661_), .Y(new_n20662_));
  AND2X1   g18226(.A(new_n20662_), .B(new_n20603_), .Y(new_n20663_));
  OAI21X1  g18227(.A0(new_n20600_), .A1(new_n12578_), .B0(new_n20599_), .Y(new_n20664_));
  MX2X1    g18228(.A(new_n20664_), .B(new_n20597_), .S0(new_n11763_), .Y(new_n20665_));
  OAI21X1  g18229(.A0(new_n20665_), .A1(pi0644), .B0(pi0715), .Y(new_n20666_));
  AOI21X1  g18230(.A0(new_n20663_), .A1(pi0644), .B0(new_n20666_), .Y(new_n20667_));
  OR3X1    g18231(.A(new_n20565_), .B(new_n12603_), .C(new_n11763_), .Y(new_n20668_));
  OAI21X1  g18232(.A0(new_n20585_), .A1(new_n12604_), .B0(new_n20668_), .Y(new_n20669_));
  OAI21X1  g18233(.A0(new_n20565_), .A1(pi0644), .B0(new_n12608_), .Y(new_n20670_));
  AOI21X1  g18234(.A0(new_n20669_), .A1(pi0644), .B0(new_n20670_), .Y(new_n20671_));
  OR2X1    g18235(.A(new_n20671_), .B(new_n11762_), .Y(new_n20672_));
  OAI21X1  g18236(.A0(new_n20665_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n20673_));
  AOI21X1  g18237(.A0(new_n20663_), .A1(new_n12612_), .B0(new_n20673_), .Y(new_n20674_));
  OAI21X1  g18238(.A0(new_n20565_), .A1(new_n12612_), .B0(pi0715), .Y(new_n20675_));
  AOI21X1  g18239(.A0(new_n20669_), .A1(new_n12612_), .B0(new_n20675_), .Y(new_n20676_));
  OR2X1    g18240(.A(new_n20676_), .B(pi1160), .Y(new_n20677_));
  OAI22X1  g18241(.A0(new_n20677_), .A1(new_n20674_), .B0(new_n20672_), .B1(new_n20667_), .Y(new_n20678_));
  NAND2X1  g18242(.A(new_n20678_), .B(pi0790), .Y(new_n20679_));
  AOI21X1  g18243(.A0(new_n20663_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n20680_));
  AOI21X1  g18244(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0191), .Y(new_n20681_));
  INVX1    g18245(.A(new_n20681_), .Y(new_n20682_));
  OAI21X1  g18246(.A0(new_n12826_), .A1(new_n6810_), .B0(new_n2979_), .Y(new_n20683_));
  AOI21X1  g18247(.A0(new_n12825_), .A1(new_n6810_), .B0(new_n20683_), .Y(new_n20684_));
  AOI21X1  g18248(.A0(new_n12771_), .A1(new_n6810_), .B0(new_n12441_), .Y(new_n20685_));
  NOR3X1   g18249(.A(new_n20685_), .B(new_n20684_), .C(new_n15412_), .Y(new_n20686_));
  OR2X1    g18250(.A(pi0729), .B(pi0191), .Y(new_n20687_));
  OAI21X1  g18251(.A0(new_n20687_), .A1(new_n12447_), .B0(new_n3103_), .Y(new_n20688_));
  OAI22X1  g18252(.A0(new_n20688_), .A1(new_n20686_), .B0(new_n3103_), .B1(new_n6810_), .Y(new_n20689_));
  AND2X1   g18253(.A(new_n20689_), .B(new_n11769_), .Y(new_n20690_));
  AOI21X1  g18254(.A0(new_n20681_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n20691_));
  OAI21X1  g18255(.A0(new_n20689_), .A1(new_n12363_), .B0(new_n20691_), .Y(new_n20692_));
  AOI21X1  g18256(.A0(new_n20681_), .A1(pi0625), .B0(pi1153), .Y(new_n20693_));
  OAI21X1  g18257(.A0(new_n20689_), .A1(pi0625), .B0(new_n20693_), .Y(new_n20694_));
  AOI21X1  g18258(.A0(new_n20694_), .A1(new_n20692_), .B0(new_n11769_), .Y(new_n20695_));
  NOR2X1   g18259(.A(new_n20695_), .B(new_n20690_), .Y(new_n20696_));
  MX2X1    g18260(.A(new_n20696_), .B(new_n20681_), .S0(new_n12490_), .Y(new_n20697_));
  AND2X1   g18261(.A(new_n20681_), .B(new_n12513_), .Y(new_n20698_));
  AOI21X1  g18262(.A0(new_n20697_), .A1(new_n14053_), .B0(new_n20698_), .Y(new_n20699_));
  MX2X1    g18263(.A(new_n20699_), .B(new_n20682_), .S0(new_n12531_), .Y(new_n20700_));
  MX2X1    g18264(.A(new_n20700_), .B(new_n20682_), .S0(new_n12563_), .Y(new_n20701_));
  MX2X1    g18265(.A(new_n20701_), .B(new_n20682_), .S0(pi0628), .Y(new_n20702_));
  MX2X1    g18266(.A(new_n20701_), .B(new_n20682_), .S0(new_n12554_), .Y(new_n20703_));
  MX2X1    g18267(.A(new_n20703_), .B(new_n20702_), .S0(new_n12555_), .Y(new_n20704_));
  MX2X1    g18268(.A(new_n20704_), .B(new_n20701_), .S0(new_n11764_), .Y(new_n20705_));
  MX2X1    g18269(.A(new_n20705_), .B(new_n20682_), .S0(pi0647), .Y(new_n20706_));
  MX2X1    g18270(.A(new_n20705_), .B(new_n20682_), .S0(new_n12577_), .Y(new_n20707_));
  MX2X1    g18271(.A(new_n20707_), .B(new_n20706_), .S0(new_n12578_), .Y(new_n20708_));
  MX2X1    g18272(.A(new_n20708_), .B(new_n20705_), .S0(new_n11763_), .Y(new_n20709_));
  OAI21X1  g18273(.A0(new_n20709_), .A1(pi0644), .B0(pi0715), .Y(new_n20710_));
  AOI22X1  g18274(.A0(new_n12073_), .A1(pi0191), .B0(new_n12444_), .B1(new_n15416_), .Y(new_n20711_));
  OR3X1    g18275(.A(new_n12776_), .B(new_n15416_), .C(pi0191), .Y(new_n20712_));
  OAI21X1  g18276(.A0(new_n12045_), .A1(pi0039), .B0(pi0746), .Y(new_n20713_));
  AOI21X1  g18277(.A0(new_n20713_), .A1(pi0191), .B0(new_n15417_), .Y(new_n20714_));
  AND2X1   g18278(.A(new_n20714_), .B(new_n20712_), .Y(new_n20715_));
  OAI21X1  g18279(.A0(new_n20711_), .A1(new_n2939_), .B0(new_n20715_), .Y(new_n20716_));
  OAI21X1  g18280(.A0(new_n12077_), .A1(pi0191), .B0(pi0038), .Y(new_n20717_));
  AOI21X1  g18281(.A0(new_n12079_), .A1(pi0746), .B0(new_n20717_), .Y(new_n20718_));
  AOI21X1  g18282(.A0(new_n20716_), .A1(new_n2979_), .B0(new_n20718_), .Y(new_n20719_));
  MX2X1    g18283(.A(new_n20719_), .B(new_n6810_), .S0(new_n11770_), .Y(new_n20720_));
  MX2X1    g18284(.A(new_n20720_), .B(new_n20681_), .S0(new_n12473_), .Y(new_n20721_));
  NOR2X1   g18285(.A(new_n20720_), .B(new_n12473_), .Y(new_n20722_));
  AOI22X1  g18286(.A0(new_n20722_), .A1(pi0609), .B0(new_n20682_), .B1(new_n12472_), .Y(new_n20723_));
  AOI22X1  g18287(.A0(new_n20722_), .A1(new_n12462_), .B0(new_n20682_), .B1(new_n12481_), .Y(new_n20724_));
  MX2X1    g18288(.A(new_n20724_), .B(new_n20723_), .S0(pi1155), .Y(new_n20725_));
  MX2X1    g18289(.A(new_n20725_), .B(new_n20721_), .S0(new_n11768_), .Y(new_n20726_));
  OAI21X1  g18290(.A0(new_n20682_), .A1(pi0618), .B0(pi1154), .Y(new_n20727_));
  AOI21X1  g18291(.A0(new_n20726_), .A1(pi0618), .B0(new_n20727_), .Y(new_n20728_));
  OAI21X1  g18292(.A0(new_n20682_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20729_));
  AOI21X1  g18293(.A0(new_n20726_), .A1(new_n12486_), .B0(new_n20729_), .Y(new_n20730_));
  NOR2X1   g18294(.A(new_n20730_), .B(new_n20728_), .Y(new_n20731_));
  MX2X1    g18295(.A(new_n20731_), .B(new_n20726_), .S0(new_n11767_), .Y(new_n20732_));
  OAI21X1  g18296(.A0(new_n20682_), .A1(pi0619), .B0(pi1159), .Y(new_n20733_));
  AOI21X1  g18297(.A0(new_n20732_), .A1(pi0619), .B0(new_n20733_), .Y(new_n20734_));
  OAI21X1  g18298(.A0(new_n20682_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n20735_));
  AOI21X1  g18299(.A0(new_n20732_), .A1(new_n12509_), .B0(new_n20735_), .Y(new_n20736_));
  NOR2X1   g18300(.A(new_n20736_), .B(new_n20734_), .Y(new_n20737_));
  MX2X1    g18301(.A(new_n20737_), .B(new_n20732_), .S0(new_n11766_), .Y(new_n20738_));
  AND2X1   g18302(.A(new_n20681_), .B(new_n12708_), .Y(new_n20739_));
  AOI21X1  g18303(.A0(new_n20738_), .A1(new_n16140_), .B0(new_n20739_), .Y(new_n20740_));
  MX2X1    g18304(.A(new_n20740_), .B(new_n20682_), .S0(new_n12580_), .Y(new_n20741_));
  MX2X1    g18305(.A(new_n20741_), .B(new_n20682_), .S0(new_n12604_), .Y(new_n20742_));
  AOI21X1  g18306(.A0(new_n20681_), .A1(new_n12612_), .B0(pi0715), .Y(new_n20743_));
  OAI21X1  g18307(.A0(new_n20742_), .A1(new_n12612_), .B0(new_n20743_), .Y(new_n20744_));
  NAND3X1  g18308(.A(new_n20744_), .B(new_n20710_), .C(pi1160), .Y(new_n20745_));
  OAI21X1  g18309(.A0(new_n20709_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n20746_));
  AOI21X1  g18310(.A0(new_n20681_), .A1(pi0644), .B0(new_n12608_), .Y(new_n20747_));
  OAI21X1  g18311(.A0(new_n20742_), .A1(pi0644), .B0(new_n20747_), .Y(new_n20748_));
  NAND3X1  g18312(.A(new_n20748_), .B(new_n20746_), .C(new_n11762_), .Y(new_n20749_));
  AND2X1   g18313(.A(new_n20749_), .B(new_n20745_), .Y(new_n20750_));
  NAND3X1  g18314(.A(new_n20748_), .B(new_n11762_), .C(new_n12612_), .Y(new_n20751_));
  NAND3X1  g18315(.A(new_n20744_), .B(pi1160), .C(pi0644), .Y(new_n20752_));
  AND3X1   g18316(.A(new_n20752_), .B(new_n20751_), .C(pi0790), .Y(new_n20753_));
  NAND2X1  g18317(.A(new_n20740_), .B(new_n14249_), .Y(new_n20754_));
  AOI22X1  g18318(.A0(new_n20703_), .A1(new_n16373_), .B0(new_n20702_), .B1(new_n16374_), .Y(new_n20755_));
  AOI21X1  g18319(.A0(new_n20755_), .A1(new_n20754_), .B0(new_n11764_), .Y(new_n20756_));
  AND2X1   g18320(.A(new_n20719_), .B(new_n15412_), .Y(new_n20757_));
  INVX1    g18321(.A(new_n20757_), .Y(new_n20758_));
  AOI21X1  g18322(.A0(new_n16381_), .A1(pi0191), .B0(pi0746), .Y(new_n20759_));
  OAI21X1  g18323(.A0(new_n16380_), .A1(pi0191), .B0(new_n20759_), .Y(new_n20760_));
  AOI21X1  g18324(.A0(new_n12788_), .A1(new_n6810_), .B0(new_n15416_), .Y(new_n20761_));
  OAI21X1  g18325(.A0(new_n12787_), .A1(new_n6810_), .B0(new_n20761_), .Y(new_n20762_));
  AND2X1   g18326(.A(new_n20762_), .B(pi0039), .Y(new_n20763_));
  AND2X1   g18327(.A(new_n20763_), .B(new_n20760_), .Y(new_n20764_));
  AOI21X1  g18328(.A0(new_n12795_), .A1(pi0191), .B0(pi0746), .Y(new_n20765_));
  OAI21X1  g18329(.A0(new_n12792_), .A1(pi0191), .B0(new_n20765_), .Y(new_n20766_));
  NOR2X1   g18330(.A(new_n12798_), .B(pi0191), .Y(new_n20767_));
  INVX1    g18331(.A(new_n20767_), .Y(new_n20768_));
  AOI21X1  g18332(.A0(new_n12800_), .A1(pi0191), .B0(new_n15416_), .Y(new_n20769_));
  AOI21X1  g18333(.A0(new_n20769_), .A1(new_n20768_), .B0(pi0039), .Y(new_n20770_));
  AOI21X1  g18334(.A0(new_n20770_), .A1(new_n20766_), .B0(pi0038), .Y(new_n20771_));
  INVX1    g18335(.A(new_n20771_), .Y(new_n20772_));
  AOI21X1  g18336(.A0(new_n16396_), .A1(new_n15416_), .B0(new_n12276_), .Y(new_n20773_));
  OAI21X1  g18337(.A0(new_n20773_), .A1(pi0039), .B0(new_n6810_), .Y(new_n20774_));
  OAI21X1  g18338(.A0(new_n20566_), .A1(new_n13443_), .B0(pi0191), .Y(new_n20775_));
  OAI21X1  g18339(.A0(new_n20775_), .A1(new_n16399_), .B0(pi0038), .Y(new_n20776_));
  INVX1    g18340(.A(new_n20776_), .Y(new_n20777_));
  AOI21X1  g18341(.A0(new_n20777_), .A1(new_n20774_), .B0(new_n15412_), .Y(new_n20778_));
  OAI21X1  g18342(.A0(new_n20772_), .A1(new_n20764_), .B0(new_n20778_), .Y(new_n20779_));
  AND2X1   g18343(.A(new_n20779_), .B(new_n3103_), .Y(new_n20780_));
  AOI22X1  g18344(.A0(new_n20780_), .A1(new_n20758_), .B0(new_n11770_), .B1(pi0191), .Y(new_n20781_));
  INVX1    g18345(.A(new_n20781_), .Y(new_n20782_));
  AOI21X1  g18346(.A0(new_n20720_), .A1(pi0625), .B0(pi1153), .Y(new_n20783_));
  OAI21X1  g18347(.A0(new_n20782_), .A1(pi0625), .B0(new_n20783_), .Y(new_n20784_));
  AND2X1   g18348(.A(new_n20692_), .B(new_n12368_), .Y(new_n20785_));
  AOI21X1  g18349(.A0(new_n20720_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n20786_));
  OAI21X1  g18350(.A0(new_n20782_), .A1(new_n12363_), .B0(new_n20786_), .Y(new_n20787_));
  AND2X1   g18351(.A(new_n20694_), .B(pi0608), .Y(new_n20788_));
  AOI22X1  g18352(.A0(new_n20788_), .A1(new_n20787_), .B0(new_n20785_), .B1(new_n20784_), .Y(new_n20789_));
  MX2X1    g18353(.A(new_n20789_), .B(new_n20782_), .S0(new_n11769_), .Y(new_n20790_));
  AOI21X1  g18354(.A0(new_n20696_), .A1(pi0609), .B0(pi1155), .Y(new_n20791_));
  OAI21X1  g18355(.A0(new_n20790_), .A1(pi0609), .B0(new_n20791_), .Y(new_n20792_));
  OAI21X1  g18356(.A0(new_n20723_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n20793_));
  INVX1    g18357(.A(new_n20793_), .Y(new_n20794_));
  AOI21X1  g18358(.A0(new_n20696_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n20795_));
  OAI21X1  g18359(.A0(new_n20790_), .A1(new_n12462_), .B0(new_n20795_), .Y(new_n20796_));
  OAI21X1  g18360(.A0(new_n20724_), .A1(pi1155), .B0(pi0660), .Y(new_n20797_));
  INVX1    g18361(.A(new_n20797_), .Y(new_n20798_));
  AOI22X1  g18362(.A0(new_n20798_), .A1(new_n20796_), .B0(new_n20794_), .B1(new_n20792_), .Y(new_n20799_));
  MX2X1    g18363(.A(new_n20799_), .B(new_n20790_), .S0(new_n11768_), .Y(new_n20800_));
  AOI21X1  g18364(.A0(new_n20697_), .A1(pi0618), .B0(pi1154), .Y(new_n20801_));
  OAI21X1  g18365(.A0(new_n20800_), .A1(pi0618), .B0(new_n20801_), .Y(new_n20802_));
  NOR2X1   g18366(.A(new_n20728_), .B(pi0627), .Y(new_n20803_));
  AOI21X1  g18367(.A0(new_n20697_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20804_));
  OAI21X1  g18368(.A0(new_n20800_), .A1(new_n12486_), .B0(new_n20804_), .Y(new_n20805_));
  NOR2X1   g18369(.A(new_n20730_), .B(new_n12494_), .Y(new_n20806_));
  AOI22X1  g18370(.A0(new_n20806_), .A1(new_n20805_), .B0(new_n20803_), .B1(new_n20802_), .Y(new_n20807_));
  MX2X1    g18371(.A(new_n20807_), .B(new_n20800_), .S0(new_n11767_), .Y(new_n20808_));
  INVX1    g18372(.A(new_n20808_), .Y(new_n20809_));
  OAI21X1  g18373(.A0(new_n20699_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n20810_));
  AOI21X1  g18374(.A0(new_n20809_), .A1(new_n12509_), .B0(new_n20810_), .Y(new_n20811_));
  NOR3X1   g18375(.A(new_n20811_), .B(new_n20734_), .C(pi0648), .Y(new_n20812_));
  OAI21X1  g18376(.A0(new_n20699_), .A1(pi0619), .B0(pi1159), .Y(new_n20813_));
  AOI21X1  g18377(.A0(new_n20809_), .A1(pi0619), .B0(new_n20813_), .Y(new_n20814_));
  OR2X1    g18378(.A(new_n20736_), .B(new_n12517_), .Y(new_n20815_));
  OAI21X1  g18379(.A0(new_n20815_), .A1(new_n20814_), .B0(pi0789), .Y(new_n20816_));
  AOI21X1  g18380(.A0(new_n20808_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n20817_));
  OAI21X1  g18381(.A0(new_n20816_), .A1(new_n20812_), .B0(new_n20817_), .Y(new_n20818_));
  AOI21X1  g18382(.A0(new_n20682_), .A1(pi0626), .B0(new_n16218_), .Y(new_n20819_));
  OAI21X1  g18383(.A0(new_n20738_), .A1(pi0626), .B0(new_n20819_), .Y(new_n20820_));
  AOI21X1  g18384(.A0(new_n20682_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n20821_));
  OAI21X1  g18385(.A0(new_n20738_), .A1(new_n12542_), .B0(new_n20821_), .Y(new_n20822_));
  OR2X1    g18386(.A(new_n20700_), .B(new_n13439_), .Y(new_n20823_));
  NAND3X1  g18387(.A(new_n20823_), .B(new_n20822_), .C(new_n20820_), .Y(new_n20824_));
  AOI21X1  g18388(.A0(new_n20824_), .A1(pi0788), .B0(new_n14125_), .Y(new_n20825_));
  AOI21X1  g18389(.A0(new_n20825_), .A1(new_n20818_), .B0(new_n20756_), .Y(new_n20826_));
  AND2X1   g18390(.A(new_n20741_), .B(new_n14326_), .Y(new_n20827_));
  AND2X1   g18391(.A(new_n20707_), .B(new_n14241_), .Y(new_n20828_));
  AND2X1   g18392(.A(new_n20706_), .B(new_n14243_), .Y(new_n20829_));
  OR2X1    g18393(.A(new_n20829_), .B(new_n20828_), .Y(new_n20830_));
  OAI21X1  g18394(.A0(new_n20830_), .A1(new_n20827_), .B0(pi0787), .Y(new_n20831_));
  OAI21X1  g18395(.A0(new_n20826_), .A1(new_n14121_), .B0(new_n20831_), .Y(new_n20832_));
  OAI22X1  g18396(.A0(new_n20832_), .A1(new_n20753_), .B0(new_n20750_), .B1(new_n12766_), .Y(new_n20833_));
  OAI21X1  g18397(.A0(new_n6489_), .A1(pi0191), .B0(new_n12767_), .Y(new_n20834_));
  AOI21X1  g18398(.A0(new_n20833_), .A1(new_n6489_), .B0(new_n20834_), .Y(new_n20835_));
  AOI21X1  g18399(.A0(new_n20680_), .A1(new_n20679_), .B0(new_n20835_), .Y(po0348));
  AOI21X1  g18400(.A0(pi1093), .A1(pi1092), .B0(pi0192), .Y(new_n20837_));
  INVX1    g18401(.A(new_n20837_), .Y(new_n20838_));
  AND2X1   g18402(.A(new_n12056_), .B(pi0764), .Y(new_n20839_));
  OAI21X1  g18403(.A0(new_n20839_), .A1(new_n20837_), .B0(new_n15771_), .Y(new_n20840_));
  AND3X1   g18404(.A(new_n12480_), .B(new_n12056_), .C(pi0764), .Y(new_n20841_));
  OAI21X1  g18405(.A0(new_n20841_), .A1(new_n20840_), .B0(pi1155), .Y(new_n20842_));
  NOR3X1   g18406(.A(new_n20841_), .B(new_n20837_), .C(pi1155), .Y(new_n20843_));
  INVX1    g18407(.A(new_n20843_), .Y(new_n20844_));
  AOI21X1  g18408(.A0(new_n20844_), .A1(new_n20842_), .B0(new_n11768_), .Y(new_n20845_));
  AOI21X1  g18409(.A0(new_n20840_), .A1(new_n11768_), .B0(new_n20845_), .Y(new_n20846_));
  AOI21X1  g18410(.A0(new_n20846_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n20847_));
  AOI21X1  g18411(.A0(new_n20846_), .A1(new_n12655_), .B0(pi1154), .Y(new_n20848_));
  NOR2X1   g18412(.A(new_n20848_), .B(new_n20847_), .Y(new_n20849_));
  MX2X1    g18413(.A(new_n20849_), .B(new_n20846_), .S0(new_n11767_), .Y(new_n20850_));
  NOR2X1   g18414(.A(new_n20850_), .B(pi0789), .Y(new_n20851_));
  AOI21X1  g18415(.A0(new_n20850_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n20852_));
  AOI21X1  g18416(.A0(new_n20850_), .A1(new_n15790_), .B0(pi1159), .Y(new_n20853_));
  OR2X1    g18417(.A(new_n20853_), .B(new_n20852_), .Y(new_n20854_));
  AOI21X1  g18418(.A0(new_n20854_), .A1(pi0789), .B0(new_n20851_), .Y(new_n20855_));
  INVX1    g18419(.A(new_n20855_), .Y(new_n20856_));
  MX2X1    g18420(.A(new_n20856_), .B(new_n20838_), .S0(new_n12708_), .Y(new_n20857_));
  MX2X1    g18421(.A(new_n20857_), .B(new_n20838_), .S0(new_n12580_), .Y(new_n20858_));
  AOI21X1  g18422(.A0(new_n12439_), .A1(pi0691), .B0(new_n20837_), .Y(new_n20859_));
  OR2X1    g18423(.A(new_n20859_), .B(pi0778), .Y(new_n20860_));
  INVX1    g18424(.A(new_n20859_), .Y(new_n20861_));
  AND3X1   g18425(.A(new_n12439_), .B(pi0691), .C(new_n12363_), .Y(new_n20862_));
  INVX1    g18426(.A(new_n20862_), .Y(new_n20863_));
  AOI21X1  g18427(.A0(new_n20863_), .A1(new_n20861_), .B0(new_n12364_), .Y(new_n20864_));
  NOR3X1   g18428(.A(new_n20862_), .B(new_n20837_), .C(pi1153), .Y(new_n20865_));
  OR3X1    g18429(.A(new_n20865_), .B(new_n20864_), .C(new_n11769_), .Y(new_n20866_));
  AND2X1   g18430(.A(new_n20866_), .B(new_n20860_), .Y(new_n20867_));
  NOR4X1   g18431(.A(new_n20867_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n20868_));
  AND3X1   g18432(.A(new_n20868_), .B(new_n12739_), .C(new_n12718_), .Y(new_n20869_));
  INVX1    g18433(.A(new_n20869_), .Y(new_n20870_));
  AOI21X1  g18434(.A0(new_n20837_), .A1(pi0647), .B0(pi1157), .Y(new_n20871_));
  OAI21X1  g18435(.A0(new_n20870_), .A1(pi0647), .B0(new_n20871_), .Y(new_n20872_));
  MX2X1    g18436(.A(new_n20869_), .B(new_n20837_), .S0(new_n12577_), .Y(new_n20873_));
  OAI22X1  g18437(.A0(new_n20873_), .A1(new_n14242_), .B0(new_n20872_), .B1(new_n12592_), .Y(new_n20874_));
  AOI21X1  g18438(.A0(new_n20858_), .A1(new_n14326_), .B0(new_n20874_), .Y(new_n20875_));
  OR2X1    g18439(.A(new_n20875_), .B(new_n11763_), .Y(new_n20876_));
  AOI21X1  g18440(.A0(new_n20838_), .A1(pi0626), .B0(new_n16218_), .Y(new_n20877_));
  OAI21X1  g18441(.A0(new_n20855_), .A1(pi0626), .B0(new_n20877_), .Y(new_n20878_));
  AOI21X1  g18442(.A0(new_n20838_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n20879_));
  OAI21X1  g18443(.A0(new_n20855_), .A1(new_n12542_), .B0(new_n20879_), .Y(new_n20880_));
  NAND2X1  g18444(.A(new_n20868_), .B(new_n12637_), .Y(new_n20881_));
  AND3X1   g18445(.A(new_n20881_), .B(new_n20880_), .C(new_n20878_), .Y(new_n20882_));
  NOR2X1   g18446(.A(new_n20882_), .B(new_n11765_), .Y(new_n20883_));
  NOR2X1   g18447(.A(new_n20837_), .B(pi1153), .Y(new_n20884_));
  NOR3X1   g18448(.A(new_n20859_), .B(new_n11991_), .C(new_n12363_), .Y(new_n20885_));
  AOI21X1  g18449(.A0(new_n12056_), .A1(pi0764), .B0(new_n20837_), .Y(new_n20886_));
  INVX1    g18450(.A(new_n20886_), .Y(new_n20887_));
  AOI21X1  g18451(.A0(new_n20861_), .A1(new_n12048_), .B0(new_n20887_), .Y(new_n20888_));
  OAI21X1  g18452(.A0(new_n20888_), .A1(new_n20885_), .B0(new_n20884_), .Y(new_n20889_));
  NOR2X1   g18453(.A(new_n20864_), .B(pi0608), .Y(new_n20890_));
  NOR3X1   g18454(.A(new_n20885_), .B(new_n20887_), .C(new_n12364_), .Y(new_n20891_));
  NOR3X1   g18455(.A(new_n20891_), .B(new_n20865_), .C(new_n12368_), .Y(new_n20892_));
  AOI21X1  g18456(.A0(new_n20890_), .A1(new_n20889_), .B0(new_n20892_), .Y(new_n20893_));
  OR2X1    g18457(.A(new_n20888_), .B(pi0778), .Y(new_n20894_));
  OAI21X1  g18458(.A0(new_n20893_), .A1(new_n11769_), .B0(new_n20894_), .Y(new_n20895_));
  INVX1    g18459(.A(new_n20895_), .Y(new_n20896_));
  AND2X1   g18460(.A(new_n20895_), .B(new_n12462_), .Y(new_n20897_));
  OAI21X1  g18461(.A0(new_n20867_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n20898_));
  OR2X1    g18462(.A(new_n20898_), .B(new_n20897_), .Y(new_n20899_));
  AND3X1   g18463(.A(new_n20899_), .B(new_n20842_), .C(new_n12468_), .Y(new_n20900_));
  OAI21X1  g18464(.A0(new_n20867_), .A1(pi0609), .B0(pi1155), .Y(new_n20901_));
  AOI21X1  g18465(.A0(new_n20895_), .A1(pi0609), .B0(new_n20901_), .Y(new_n20902_));
  NOR3X1   g18466(.A(new_n20902_), .B(new_n20843_), .C(new_n12468_), .Y(new_n20903_));
  NOR2X1   g18467(.A(new_n20903_), .B(new_n20900_), .Y(new_n20904_));
  MX2X1    g18468(.A(new_n20904_), .B(new_n20896_), .S0(new_n11768_), .Y(new_n20905_));
  AOI21X1  g18469(.A0(new_n20866_), .A1(new_n20860_), .B0(new_n12630_), .Y(new_n20906_));
  AOI21X1  g18470(.A0(new_n20906_), .A1(pi0618), .B0(pi1154), .Y(new_n20907_));
  OAI21X1  g18471(.A0(new_n20905_), .A1(pi0618), .B0(new_n20907_), .Y(new_n20908_));
  NOR2X1   g18472(.A(new_n20847_), .B(pi0627), .Y(new_n20909_));
  AOI21X1  g18473(.A0(new_n20906_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n20910_));
  OAI21X1  g18474(.A0(new_n20905_), .A1(new_n12486_), .B0(new_n20910_), .Y(new_n20911_));
  NOR2X1   g18475(.A(new_n20848_), .B(new_n12494_), .Y(new_n20912_));
  AOI22X1  g18476(.A0(new_n20912_), .A1(new_n20911_), .B0(new_n20909_), .B1(new_n20908_), .Y(new_n20913_));
  MX2X1    g18477(.A(new_n20913_), .B(new_n20905_), .S0(new_n11767_), .Y(new_n20914_));
  OR4X1    g18478(.A(new_n20867_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n20915_));
  AND2X1   g18479(.A(new_n20915_), .B(new_n12510_), .Y(new_n20916_));
  OAI21X1  g18480(.A0(new_n20914_), .A1(pi0619), .B0(new_n20916_), .Y(new_n20917_));
  NOR2X1   g18481(.A(new_n20852_), .B(pi0648), .Y(new_n20918_));
  AND2X1   g18482(.A(new_n20918_), .B(new_n20917_), .Y(new_n20919_));
  NOR4X1   g18483(.A(new_n20867_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n20920_));
  NOR2X1   g18484(.A(new_n20920_), .B(new_n12510_), .Y(new_n20921_));
  OAI21X1  g18485(.A0(new_n20914_), .A1(new_n12509_), .B0(new_n20921_), .Y(new_n20922_));
  NOR2X1   g18486(.A(new_n20853_), .B(new_n12517_), .Y(new_n20923_));
  AND2X1   g18487(.A(new_n20923_), .B(new_n20922_), .Y(new_n20924_));
  OR3X1    g18488(.A(new_n20924_), .B(new_n20919_), .C(new_n11766_), .Y(new_n20925_));
  AOI21X1  g18489(.A0(new_n20914_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n20926_));
  AOI21X1  g18490(.A0(new_n20926_), .A1(new_n20925_), .B0(new_n20883_), .Y(new_n20927_));
  INVX1    g18491(.A(new_n20857_), .Y(new_n20928_));
  AND2X1   g18492(.A(new_n20868_), .B(new_n12718_), .Y(new_n20929_));
  AOI22X1  g18493(.A0(new_n20929_), .A1(new_n14426_), .B0(new_n20928_), .B1(new_n12735_), .Y(new_n20930_));
  AOI22X1  g18494(.A0(new_n20929_), .A1(new_n14428_), .B0(new_n20928_), .B1(new_n12733_), .Y(new_n20931_));
  MX2X1    g18495(.A(new_n20931_), .B(new_n20930_), .S0(new_n12561_), .Y(new_n20932_));
  OAI21X1  g18496(.A0(new_n20932_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n20933_));
  INVX1    g18497(.A(new_n20933_), .Y(new_n20934_));
  OAI21X1  g18498(.A0(new_n20927_), .A1(new_n14125_), .B0(new_n20934_), .Y(new_n20935_));
  AND2X1   g18499(.A(new_n20935_), .B(new_n20876_), .Y(new_n20936_));
  OAI21X1  g18500(.A0(new_n20873_), .A1(new_n12578_), .B0(new_n20872_), .Y(new_n20937_));
  MX2X1    g18501(.A(new_n20937_), .B(new_n20870_), .S0(new_n11763_), .Y(new_n20938_));
  OAI21X1  g18502(.A0(new_n20938_), .A1(pi0644), .B0(pi0715), .Y(new_n20939_));
  AOI21X1  g18503(.A0(new_n20936_), .A1(pi0644), .B0(new_n20939_), .Y(new_n20940_));
  OR3X1    g18504(.A(new_n20838_), .B(new_n12603_), .C(new_n11763_), .Y(new_n20941_));
  OAI21X1  g18505(.A0(new_n20858_), .A1(new_n12604_), .B0(new_n20941_), .Y(new_n20942_));
  OAI21X1  g18506(.A0(new_n20838_), .A1(pi0644), .B0(new_n12608_), .Y(new_n20943_));
  AOI21X1  g18507(.A0(new_n20942_), .A1(pi0644), .B0(new_n20943_), .Y(new_n20944_));
  OR2X1    g18508(.A(new_n20944_), .B(new_n11762_), .Y(new_n20945_));
  OAI21X1  g18509(.A0(new_n20938_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n20946_));
  AOI21X1  g18510(.A0(new_n20936_), .A1(new_n12612_), .B0(new_n20946_), .Y(new_n20947_));
  OAI21X1  g18511(.A0(new_n20838_), .A1(new_n12612_), .B0(pi0715), .Y(new_n20948_));
  AOI21X1  g18512(.A0(new_n20942_), .A1(new_n12612_), .B0(new_n20948_), .Y(new_n20949_));
  OR2X1    g18513(.A(new_n20949_), .B(pi1160), .Y(new_n20950_));
  OAI22X1  g18514(.A0(new_n20950_), .A1(new_n20947_), .B0(new_n20945_), .B1(new_n20940_), .Y(new_n20951_));
  NAND2X1  g18515(.A(new_n20951_), .B(pi0790), .Y(new_n20952_));
  AOI21X1  g18516(.A0(new_n20936_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n20953_));
  AOI21X1  g18517(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0192), .Y(new_n20954_));
  INVX1    g18518(.A(new_n20954_), .Y(new_n20955_));
  OAI21X1  g18519(.A0(new_n12826_), .A1(new_n11458_), .B0(new_n2979_), .Y(new_n20956_));
  AOI21X1  g18520(.A0(new_n12825_), .A1(new_n11458_), .B0(new_n20956_), .Y(new_n20957_));
  AOI21X1  g18521(.A0(new_n12771_), .A1(new_n11458_), .B0(new_n12441_), .Y(new_n20958_));
  NOR3X1   g18522(.A(new_n20958_), .B(new_n20957_), .C(new_n15513_), .Y(new_n20959_));
  OR2X1    g18523(.A(pi0691), .B(pi0192), .Y(new_n20960_));
  OAI21X1  g18524(.A0(new_n20960_), .A1(new_n12447_), .B0(new_n3103_), .Y(new_n20961_));
  OAI22X1  g18525(.A0(new_n20961_), .A1(new_n20959_), .B0(new_n3103_), .B1(new_n11458_), .Y(new_n20962_));
  AND2X1   g18526(.A(new_n20962_), .B(new_n11769_), .Y(new_n20963_));
  AOI21X1  g18527(.A0(new_n20954_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n20964_));
  OAI21X1  g18528(.A0(new_n20962_), .A1(new_n12363_), .B0(new_n20964_), .Y(new_n20965_));
  AOI21X1  g18529(.A0(new_n20954_), .A1(pi0625), .B0(pi1153), .Y(new_n20966_));
  OAI21X1  g18530(.A0(new_n20962_), .A1(pi0625), .B0(new_n20966_), .Y(new_n20967_));
  AOI21X1  g18531(.A0(new_n20967_), .A1(new_n20965_), .B0(new_n11769_), .Y(new_n20968_));
  NOR2X1   g18532(.A(new_n20968_), .B(new_n20963_), .Y(new_n20969_));
  MX2X1    g18533(.A(new_n20969_), .B(new_n20954_), .S0(new_n12490_), .Y(new_n20970_));
  AND2X1   g18534(.A(new_n20954_), .B(new_n12513_), .Y(new_n20971_));
  AOI21X1  g18535(.A0(new_n20970_), .A1(new_n14053_), .B0(new_n20971_), .Y(new_n20972_));
  MX2X1    g18536(.A(new_n20972_), .B(new_n20955_), .S0(new_n12531_), .Y(new_n20973_));
  MX2X1    g18537(.A(new_n20973_), .B(new_n20955_), .S0(new_n12563_), .Y(new_n20974_));
  MX2X1    g18538(.A(new_n20974_), .B(new_n20955_), .S0(pi0628), .Y(new_n20975_));
  MX2X1    g18539(.A(new_n20974_), .B(new_n20955_), .S0(new_n12554_), .Y(new_n20976_));
  MX2X1    g18540(.A(new_n20976_), .B(new_n20975_), .S0(new_n12555_), .Y(new_n20977_));
  MX2X1    g18541(.A(new_n20977_), .B(new_n20974_), .S0(new_n11764_), .Y(new_n20978_));
  MX2X1    g18542(.A(new_n20978_), .B(new_n20955_), .S0(pi0647), .Y(new_n20979_));
  MX2X1    g18543(.A(new_n20978_), .B(new_n20955_), .S0(new_n12577_), .Y(new_n20980_));
  MX2X1    g18544(.A(new_n20980_), .B(new_n20979_), .S0(new_n12578_), .Y(new_n20981_));
  MX2X1    g18545(.A(new_n20981_), .B(new_n20978_), .S0(new_n11763_), .Y(new_n20982_));
  OAI21X1  g18546(.A0(new_n20982_), .A1(pi0644), .B0(pi0715), .Y(new_n20983_));
  AOI22X1  g18547(.A0(new_n12073_), .A1(pi0192), .B0(new_n12444_), .B1(new_n15517_), .Y(new_n20984_));
  OR3X1    g18548(.A(new_n12776_), .B(new_n15517_), .C(pi0192), .Y(new_n20985_));
  OAI21X1  g18549(.A0(new_n12045_), .A1(pi0039), .B0(pi0764), .Y(new_n20986_));
  AOI21X1  g18550(.A0(new_n20986_), .A1(pi0192), .B0(new_n15518_), .Y(new_n20987_));
  AND2X1   g18551(.A(new_n20987_), .B(new_n20985_), .Y(new_n20988_));
  OAI21X1  g18552(.A0(new_n20984_), .A1(new_n2939_), .B0(new_n20988_), .Y(new_n20989_));
  OAI21X1  g18553(.A0(new_n12077_), .A1(pi0192), .B0(pi0038), .Y(new_n20990_));
  AOI21X1  g18554(.A0(new_n12079_), .A1(pi0764), .B0(new_n20990_), .Y(new_n20991_));
  AOI21X1  g18555(.A0(new_n20989_), .A1(new_n2979_), .B0(new_n20991_), .Y(new_n20992_));
  MX2X1    g18556(.A(new_n20992_), .B(new_n11458_), .S0(new_n11770_), .Y(new_n20993_));
  MX2X1    g18557(.A(new_n20993_), .B(new_n20954_), .S0(new_n12473_), .Y(new_n20994_));
  NOR2X1   g18558(.A(new_n20993_), .B(new_n12473_), .Y(new_n20995_));
  AOI22X1  g18559(.A0(new_n20995_), .A1(pi0609), .B0(new_n20955_), .B1(new_n12472_), .Y(new_n20996_));
  AOI22X1  g18560(.A0(new_n20995_), .A1(new_n12462_), .B0(new_n20955_), .B1(new_n12481_), .Y(new_n20997_));
  MX2X1    g18561(.A(new_n20997_), .B(new_n20996_), .S0(pi1155), .Y(new_n20998_));
  MX2X1    g18562(.A(new_n20998_), .B(new_n20994_), .S0(new_n11768_), .Y(new_n20999_));
  OAI21X1  g18563(.A0(new_n20955_), .A1(pi0618), .B0(pi1154), .Y(new_n21000_));
  AOI21X1  g18564(.A0(new_n20999_), .A1(pi0618), .B0(new_n21000_), .Y(new_n21001_));
  OAI21X1  g18565(.A0(new_n20955_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n21002_));
  AOI21X1  g18566(.A0(new_n20999_), .A1(new_n12486_), .B0(new_n21002_), .Y(new_n21003_));
  NOR2X1   g18567(.A(new_n21003_), .B(new_n21001_), .Y(new_n21004_));
  MX2X1    g18568(.A(new_n21004_), .B(new_n20999_), .S0(new_n11767_), .Y(new_n21005_));
  OAI21X1  g18569(.A0(new_n20955_), .A1(pi0619), .B0(pi1159), .Y(new_n21006_));
  AOI21X1  g18570(.A0(new_n21005_), .A1(pi0619), .B0(new_n21006_), .Y(new_n21007_));
  OAI21X1  g18571(.A0(new_n20955_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n21008_));
  AOI21X1  g18572(.A0(new_n21005_), .A1(new_n12509_), .B0(new_n21008_), .Y(new_n21009_));
  NOR2X1   g18573(.A(new_n21009_), .B(new_n21007_), .Y(new_n21010_));
  MX2X1    g18574(.A(new_n21010_), .B(new_n21005_), .S0(new_n11766_), .Y(new_n21011_));
  AND2X1   g18575(.A(new_n20954_), .B(new_n12708_), .Y(new_n21012_));
  AOI21X1  g18576(.A0(new_n21011_), .A1(new_n16140_), .B0(new_n21012_), .Y(new_n21013_));
  MX2X1    g18577(.A(new_n21013_), .B(new_n20955_), .S0(new_n12580_), .Y(new_n21014_));
  MX2X1    g18578(.A(new_n21014_), .B(new_n20955_), .S0(new_n12604_), .Y(new_n21015_));
  AOI21X1  g18579(.A0(new_n20954_), .A1(new_n12612_), .B0(pi0715), .Y(new_n21016_));
  OAI21X1  g18580(.A0(new_n21015_), .A1(new_n12612_), .B0(new_n21016_), .Y(new_n21017_));
  NAND3X1  g18581(.A(new_n21017_), .B(new_n20983_), .C(pi1160), .Y(new_n21018_));
  OAI21X1  g18582(.A0(new_n20982_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n21019_));
  AOI21X1  g18583(.A0(new_n20954_), .A1(pi0644), .B0(new_n12608_), .Y(new_n21020_));
  OAI21X1  g18584(.A0(new_n21015_), .A1(pi0644), .B0(new_n21020_), .Y(new_n21021_));
  NAND3X1  g18585(.A(new_n21021_), .B(new_n21019_), .C(new_n11762_), .Y(new_n21022_));
  AND2X1   g18586(.A(new_n21022_), .B(new_n21018_), .Y(new_n21023_));
  NAND3X1  g18587(.A(new_n21021_), .B(new_n11762_), .C(new_n12612_), .Y(new_n21024_));
  NAND3X1  g18588(.A(new_n21017_), .B(pi1160), .C(pi0644), .Y(new_n21025_));
  AND3X1   g18589(.A(new_n21025_), .B(new_n21024_), .C(pi0790), .Y(new_n21026_));
  NAND2X1  g18590(.A(new_n21013_), .B(new_n14249_), .Y(new_n21027_));
  AOI22X1  g18591(.A0(new_n20976_), .A1(new_n16373_), .B0(new_n20975_), .B1(new_n16374_), .Y(new_n21028_));
  AOI21X1  g18592(.A0(new_n21028_), .A1(new_n21027_), .B0(new_n11764_), .Y(new_n21029_));
  AND2X1   g18593(.A(new_n20992_), .B(new_n15513_), .Y(new_n21030_));
  INVX1    g18594(.A(new_n21030_), .Y(new_n21031_));
  AOI21X1  g18595(.A0(new_n16381_), .A1(pi0192), .B0(pi0764), .Y(new_n21032_));
  OAI21X1  g18596(.A0(new_n16380_), .A1(pi0192), .B0(new_n21032_), .Y(new_n21033_));
  AOI21X1  g18597(.A0(new_n12788_), .A1(new_n11458_), .B0(new_n15517_), .Y(new_n21034_));
  OAI21X1  g18598(.A0(new_n12787_), .A1(new_n11458_), .B0(new_n21034_), .Y(new_n21035_));
  AND2X1   g18599(.A(new_n21035_), .B(pi0039), .Y(new_n21036_));
  AND2X1   g18600(.A(new_n21036_), .B(new_n21033_), .Y(new_n21037_));
  AOI21X1  g18601(.A0(new_n12795_), .A1(pi0192), .B0(pi0764), .Y(new_n21038_));
  OAI21X1  g18602(.A0(new_n12792_), .A1(pi0192), .B0(new_n21038_), .Y(new_n21039_));
  NOR2X1   g18603(.A(new_n12798_), .B(pi0192), .Y(new_n21040_));
  INVX1    g18604(.A(new_n21040_), .Y(new_n21041_));
  AOI21X1  g18605(.A0(new_n12800_), .A1(pi0192), .B0(new_n15517_), .Y(new_n21042_));
  AOI21X1  g18606(.A0(new_n21042_), .A1(new_n21041_), .B0(pi0039), .Y(new_n21043_));
  AOI21X1  g18607(.A0(new_n21043_), .A1(new_n21039_), .B0(pi0038), .Y(new_n21044_));
  INVX1    g18608(.A(new_n21044_), .Y(new_n21045_));
  AOI21X1  g18609(.A0(new_n16396_), .A1(new_n15517_), .B0(new_n12276_), .Y(new_n21046_));
  OAI21X1  g18610(.A0(new_n21046_), .A1(pi0039), .B0(new_n11458_), .Y(new_n21047_));
  OAI21X1  g18611(.A0(new_n20839_), .A1(new_n13443_), .B0(pi0192), .Y(new_n21048_));
  OAI21X1  g18612(.A0(new_n21048_), .A1(new_n16399_), .B0(pi0038), .Y(new_n21049_));
  INVX1    g18613(.A(new_n21049_), .Y(new_n21050_));
  AOI21X1  g18614(.A0(new_n21050_), .A1(new_n21047_), .B0(new_n15513_), .Y(new_n21051_));
  OAI21X1  g18615(.A0(new_n21045_), .A1(new_n21037_), .B0(new_n21051_), .Y(new_n21052_));
  AND2X1   g18616(.A(new_n21052_), .B(new_n3103_), .Y(new_n21053_));
  AOI22X1  g18617(.A0(new_n21053_), .A1(new_n21031_), .B0(new_n11770_), .B1(pi0192), .Y(new_n21054_));
  INVX1    g18618(.A(new_n21054_), .Y(new_n21055_));
  AOI21X1  g18619(.A0(new_n20993_), .A1(pi0625), .B0(pi1153), .Y(new_n21056_));
  OAI21X1  g18620(.A0(new_n21055_), .A1(pi0625), .B0(new_n21056_), .Y(new_n21057_));
  AND2X1   g18621(.A(new_n20965_), .B(new_n12368_), .Y(new_n21058_));
  AOI21X1  g18622(.A0(new_n20993_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n21059_));
  OAI21X1  g18623(.A0(new_n21055_), .A1(new_n12363_), .B0(new_n21059_), .Y(new_n21060_));
  AND2X1   g18624(.A(new_n20967_), .B(pi0608), .Y(new_n21061_));
  AOI22X1  g18625(.A0(new_n21061_), .A1(new_n21060_), .B0(new_n21058_), .B1(new_n21057_), .Y(new_n21062_));
  MX2X1    g18626(.A(new_n21062_), .B(new_n21055_), .S0(new_n11769_), .Y(new_n21063_));
  AOI21X1  g18627(.A0(new_n20969_), .A1(pi0609), .B0(pi1155), .Y(new_n21064_));
  OAI21X1  g18628(.A0(new_n21063_), .A1(pi0609), .B0(new_n21064_), .Y(new_n21065_));
  OAI21X1  g18629(.A0(new_n20996_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n21066_));
  INVX1    g18630(.A(new_n21066_), .Y(new_n21067_));
  AOI21X1  g18631(.A0(new_n20969_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n21068_));
  OAI21X1  g18632(.A0(new_n21063_), .A1(new_n12462_), .B0(new_n21068_), .Y(new_n21069_));
  OAI21X1  g18633(.A0(new_n20997_), .A1(pi1155), .B0(pi0660), .Y(new_n21070_));
  INVX1    g18634(.A(new_n21070_), .Y(new_n21071_));
  AOI22X1  g18635(.A0(new_n21071_), .A1(new_n21069_), .B0(new_n21067_), .B1(new_n21065_), .Y(new_n21072_));
  MX2X1    g18636(.A(new_n21072_), .B(new_n21063_), .S0(new_n11768_), .Y(new_n21073_));
  AOI21X1  g18637(.A0(new_n20970_), .A1(pi0618), .B0(pi1154), .Y(new_n21074_));
  OAI21X1  g18638(.A0(new_n21073_), .A1(pi0618), .B0(new_n21074_), .Y(new_n21075_));
  NOR2X1   g18639(.A(new_n21001_), .B(pi0627), .Y(new_n21076_));
  AOI21X1  g18640(.A0(new_n20970_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n21077_));
  OAI21X1  g18641(.A0(new_n21073_), .A1(new_n12486_), .B0(new_n21077_), .Y(new_n21078_));
  NOR2X1   g18642(.A(new_n21003_), .B(new_n12494_), .Y(new_n21079_));
  AOI22X1  g18643(.A0(new_n21079_), .A1(new_n21078_), .B0(new_n21076_), .B1(new_n21075_), .Y(new_n21080_));
  MX2X1    g18644(.A(new_n21080_), .B(new_n21073_), .S0(new_n11767_), .Y(new_n21081_));
  INVX1    g18645(.A(new_n21081_), .Y(new_n21082_));
  OAI21X1  g18646(.A0(new_n20972_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n21083_));
  AOI21X1  g18647(.A0(new_n21082_), .A1(new_n12509_), .B0(new_n21083_), .Y(new_n21084_));
  NOR3X1   g18648(.A(new_n21084_), .B(new_n21007_), .C(pi0648), .Y(new_n21085_));
  OAI21X1  g18649(.A0(new_n20972_), .A1(pi0619), .B0(pi1159), .Y(new_n21086_));
  AOI21X1  g18650(.A0(new_n21082_), .A1(pi0619), .B0(new_n21086_), .Y(new_n21087_));
  OR2X1    g18651(.A(new_n21009_), .B(new_n12517_), .Y(new_n21088_));
  OAI21X1  g18652(.A0(new_n21088_), .A1(new_n21087_), .B0(pi0789), .Y(new_n21089_));
  AOI21X1  g18653(.A0(new_n21081_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n21090_));
  OAI21X1  g18654(.A0(new_n21089_), .A1(new_n21085_), .B0(new_n21090_), .Y(new_n21091_));
  AOI21X1  g18655(.A0(new_n20955_), .A1(pi0626), .B0(new_n16218_), .Y(new_n21092_));
  OAI21X1  g18656(.A0(new_n21011_), .A1(pi0626), .B0(new_n21092_), .Y(new_n21093_));
  AOI21X1  g18657(.A0(new_n20955_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n21094_));
  OAI21X1  g18658(.A0(new_n21011_), .A1(new_n12542_), .B0(new_n21094_), .Y(new_n21095_));
  OR2X1    g18659(.A(new_n20973_), .B(new_n13439_), .Y(new_n21096_));
  NAND3X1  g18660(.A(new_n21096_), .B(new_n21095_), .C(new_n21093_), .Y(new_n21097_));
  AOI21X1  g18661(.A0(new_n21097_), .A1(pi0788), .B0(new_n14125_), .Y(new_n21098_));
  AOI21X1  g18662(.A0(new_n21098_), .A1(new_n21091_), .B0(new_n21029_), .Y(new_n21099_));
  AND2X1   g18663(.A(new_n21014_), .B(new_n14326_), .Y(new_n21100_));
  AND2X1   g18664(.A(new_n20980_), .B(new_n14241_), .Y(new_n21101_));
  AND2X1   g18665(.A(new_n20979_), .B(new_n14243_), .Y(new_n21102_));
  OR2X1    g18666(.A(new_n21102_), .B(new_n21101_), .Y(new_n21103_));
  OAI21X1  g18667(.A0(new_n21103_), .A1(new_n21100_), .B0(pi0787), .Y(new_n21104_));
  OAI21X1  g18668(.A0(new_n21099_), .A1(new_n14121_), .B0(new_n21104_), .Y(new_n21105_));
  OAI22X1  g18669(.A0(new_n21105_), .A1(new_n21026_), .B0(new_n21023_), .B1(new_n12766_), .Y(new_n21106_));
  OAI21X1  g18670(.A0(new_n6489_), .A1(pi0192), .B0(new_n12767_), .Y(new_n21107_));
  AOI21X1  g18671(.A0(new_n21106_), .A1(new_n6489_), .B0(new_n21107_), .Y(new_n21108_));
  AOI21X1  g18672(.A0(new_n20953_), .A1(new_n20952_), .B0(new_n21108_), .Y(po0349));
  AOI21X1  g18673(.A0(pi1093), .A1(pi1092), .B0(pi0193), .Y(new_n21110_));
  INVX1    g18674(.A(new_n21110_), .Y(new_n21111_));
  AOI21X1  g18675(.A0(new_n12056_), .A1(pi0739), .B0(new_n21110_), .Y(new_n21112_));
  INVX1    g18676(.A(new_n21112_), .Y(new_n21113_));
  NAND2X1  g18677(.A(new_n21113_), .B(new_n15771_), .Y(new_n21114_));
  AND3X1   g18678(.A(new_n12480_), .B(new_n12056_), .C(pi0739), .Y(new_n21115_));
  OAI21X1  g18679(.A0(new_n21115_), .A1(new_n21114_), .B0(pi1155), .Y(new_n21116_));
  NOR3X1   g18680(.A(new_n21115_), .B(new_n21110_), .C(pi1155), .Y(new_n21117_));
  INVX1    g18681(.A(new_n21117_), .Y(new_n21118_));
  AOI21X1  g18682(.A0(new_n21118_), .A1(new_n21116_), .B0(new_n11768_), .Y(new_n21119_));
  AOI21X1  g18683(.A0(new_n21114_), .A1(new_n11768_), .B0(new_n21119_), .Y(new_n21120_));
  AOI21X1  g18684(.A0(new_n21120_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n21121_));
  AOI21X1  g18685(.A0(new_n21120_), .A1(new_n12655_), .B0(pi1154), .Y(new_n21122_));
  NOR2X1   g18686(.A(new_n21122_), .B(new_n21121_), .Y(new_n21123_));
  MX2X1    g18687(.A(new_n21123_), .B(new_n21120_), .S0(new_n11767_), .Y(new_n21124_));
  NOR2X1   g18688(.A(new_n21124_), .B(pi0789), .Y(new_n21125_));
  AOI21X1  g18689(.A0(new_n21124_), .A1(new_n15787_), .B0(new_n12510_), .Y(new_n21126_));
  AOI21X1  g18690(.A0(new_n21124_), .A1(new_n15790_), .B0(pi1159), .Y(new_n21127_));
  OR2X1    g18691(.A(new_n21127_), .B(new_n21126_), .Y(new_n21128_));
  AOI21X1  g18692(.A0(new_n21128_), .A1(pi0789), .B0(new_n21125_), .Y(new_n21129_));
  INVX1    g18693(.A(new_n21129_), .Y(new_n21130_));
  MX2X1    g18694(.A(new_n21130_), .B(new_n21111_), .S0(new_n12708_), .Y(new_n21131_));
  MX2X1    g18695(.A(new_n21131_), .B(new_n21111_), .S0(new_n12580_), .Y(new_n21132_));
  AOI21X1  g18696(.A0(new_n12439_), .A1(pi0690), .B0(new_n21110_), .Y(new_n21133_));
  OR2X1    g18697(.A(new_n21133_), .B(pi0778), .Y(new_n21134_));
  INVX1    g18698(.A(new_n21133_), .Y(new_n21135_));
  AND3X1   g18699(.A(new_n12439_), .B(pi0690), .C(new_n12363_), .Y(new_n21136_));
  INVX1    g18700(.A(new_n21136_), .Y(new_n21137_));
  AOI21X1  g18701(.A0(new_n21137_), .A1(new_n21135_), .B0(new_n12364_), .Y(new_n21138_));
  NOR3X1   g18702(.A(new_n21136_), .B(new_n21110_), .C(pi1153), .Y(new_n21139_));
  OR3X1    g18703(.A(new_n21139_), .B(new_n21138_), .C(new_n11769_), .Y(new_n21140_));
  AND2X1   g18704(.A(new_n21140_), .B(new_n21134_), .Y(new_n21141_));
  NOR4X1   g18705(.A(new_n21141_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n21142_));
  AND3X1   g18706(.A(new_n21142_), .B(new_n12739_), .C(new_n12718_), .Y(new_n21143_));
  INVX1    g18707(.A(new_n21143_), .Y(new_n21144_));
  AOI21X1  g18708(.A0(new_n21110_), .A1(pi0647), .B0(pi1157), .Y(new_n21145_));
  OAI21X1  g18709(.A0(new_n21144_), .A1(pi0647), .B0(new_n21145_), .Y(new_n21146_));
  MX2X1    g18710(.A(new_n21143_), .B(new_n21110_), .S0(new_n12577_), .Y(new_n21147_));
  OAI22X1  g18711(.A0(new_n21147_), .A1(new_n14242_), .B0(new_n21146_), .B1(new_n12592_), .Y(new_n21148_));
  AOI21X1  g18712(.A0(new_n21132_), .A1(new_n14326_), .B0(new_n21148_), .Y(new_n21149_));
  NOR2X1   g18713(.A(new_n21149_), .B(new_n11763_), .Y(new_n21150_));
  AOI21X1  g18714(.A0(new_n21111_), .A1(pi0626), .B0(new_n16218_), .Y(new_n21151_));
  OAI21X1  g18715(.A0(new_n21129_), .A1(pi0626), .B0(new_n21151_), .Y(new_n21152_));
  AOI21X1  g18716(.A0(new_n21111_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n21153_));
  OAI21X1  g18717(.A0(new_n21129_), .A1(new_n12542_), .B0(new_n21153_), .Y(new_n21154_));
  NAND2X1  g18718(.A(new_n21142_), .B(new_n12637_), .Y(new_n21155_));
  AND3X1   g18719(.A(new_n21155_), .B(new_n21154_), .C(new_n21152_), .Y(new_n21156_));
  NOR2X1   g18720(.A(new_n21156_), .B(new_n11765_), .Y(new_n21157_));
  NOR2X1   g18721(.A(new_n21110_), .B(pi1153), .Y(new_n21158_));
  NOR3X1   g18722(.A(new_n21133_), .B(new_n11991_), .C(new_n12363_), .Y(new_n21159_));
  AOI21X1  g18723(.A0(new_n21135_), .A1(new_n12048_), .B0(new_n21113_), .Y(new_n21160_));
  OAI21X1  g18724(.A0(new_n21160_), .A1(new_n21159_), .B0(new_n21158_), .Y(new_n21161_));
  NOR2X1   g18725(.A(new_n21138_), .B(pi0608), .Y(new_n21162_));
  NOR3X1   g18726(.A(new_n21159_), .B(new_n21113_), .C(new_n12364_), .Y(new_n21163_));
  NOR3X1   g18727(.A(new_n21163_), .B(new_n21139_), .C(new_n12368_), .Y(new_n21164_));
  AOI21X1  g18728(.A0(new_n21162_), .A1(new_n21161_), .B0(new_n21164_), .Y(new_n21165_));
  OR2X1    g18729(.A(new_n21160_), .B(pi0778), .Y(new_n21166_));
  OAI21X1  g18730(.A0(new_n21165_), .A1(new_n11769_), .B0(new_n21166_), .Y(new_n21167_));
  INVX1    g18731(.A(new_n21167_), .Y(new_n21168_));
  AND2X1   g18732(.A(new_n21167_), .B(new_n12462_), .Y(new_n21169_));
  OAI21X1  g18733(.A0(new_n21141_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n21170_));
  OR2X1    g18734(.A(new_n21170_), .B(new_n21169_), .Y(new_n21171_));
  AND3X1   g18735(.A(new_n21171_), .B(new_n21116_), .C(new_n12468_), .Y(new_n21172_));
  OAI21X1  g18736(.A0(new_n21141_), .A1(pi0609), .B0(pi1155), .Y(new_n21173_));
  AOI21X1  g18737(.A0(new_n21167_), .A1(pi0609), .B0(new_n21173_), .Y(new_n21174_));
  NOR3X1   g18738(.A(new_n21174_), .B(new_n21117_), .C(new_n12468_), .Y(new_n21175_));
  NOR2X1   g18739(.A(new_n21175_), .B(new_n21172_), .Y(new_n21176_));
  MX2X1    g18740(.A(new_n21176_), .B(new_n21168_), .S0(new_n11768_), .Y(new_n21177_));
  AOI21X1  g18741(.A0(new_n21140_), .A1(new_n21134_), .B0(new_n12630_), .Y(new_n21178_));
  AOI21X1  g18742(.A0(new_n21178_), .A1(pi0618), .B0(pi1154), .Y(new_n21179_));
  OAI21X1  g18743(.A0(new_n21177_), .A1(pi0618), .B0(new_n21179_), .Y(new_n21180_));
  NOR2X1   g18744(.A(new_n21121_), .B(pi0627), .Y(new_n21181_));
  AOI21X1  g18745(.A0(new_n21178_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n21182_));
  OAI21X1  g18746(.A0(new_n21177_), .A1(new_n12486_), .B0(new_n21182_), .Y(new_n21183_));
  NOR2X1   g18747(.A(new_n21122_), .B(new_n12494_), .Y(new_n21184_));
  AOI22X1  g18748(.A0(new_n21184_), .A1(new_n21183_), .B0(new_n21181_), .B1(new_n21180_), .Y(new_n21185_));
  MX2X1    g18749(.A(new_n21185_), .B(new_n21177_), .S0(new_n11767_), .Y(new_n21186_));
  OR4X1    g18750(.A(new_n21141_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n21187_));
  AND2X1   g18751(.A(new_n21187_), .B(new_n12510_), .Y(new_n21188_));
  OAI21X1  g18752(.A0(new_n21186_), .A1(pi0619), .B0(new_n21188_), .Y(new_n21189_));
  NOR2X1   g18753(.A(new_n21126_), .B(pi0648), .Y(new_n21190_));
  AND2X1   g18754(.A(new_n21190_), .B(new_n21189_), .Y(new_n21191_));
  NOR4X1   g18755(.A(new_n21141_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n21192_));
  NOR2X1   g18756(.A(new_n21192_), .B(new_n12510_), .Y(new_n21193_));
  OAI21X1  g18757(.A0(new_n21186_), .A1(new_n12509_), .B0(new_n21193_), .Y(new_n21194_));
  NOR2X1   g18758(.A(new_n21127_), .B(new_n12517_), .Y(new_n21195_));
  AND2X1   g18759(.A(new_n21195_), .B(new_n21194_), .Y(new_n21196_));
  OR3X1    g18760(.A(new_n21196_), .B(new_n21191_), .C(new_n11766_), .Y(new_n21197_));
  AOI21X1  g18761(.A0(new_n21186_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n21198_));
  AOI21X1  g18762(.A0(new_n21198_), .A1(new_n21197_), .B0(new_n21157_), .Y(new_n21199_));
  OR2X1    g18763(.A(new_n21199_), .B(new_n14125_), .Y(new_n21200_));
  INVX1    g18764(.A(new_n21131_), .Y(new_n21201_));
  AND2X1   g18765(.A(new_n21142_), .B(new_n12718_), .Y(new_n21202_));
  AOI22X1  g18766(.A0(new_n21202_), .A1(new_n14426_), .B0(new_n21201_), .B1(new_n12735_), .Y(new_n21203_));
  AOI22X1  g18767(.A0(new_n21202_), .A1(new_n14428_), .B0(new_n21201_), .B1(new_n12733_), .Y(new_n21204_));
  MX2X1    g18768(.A(new_n21204_), .B(new_n21203_), .S0(new_n12561_), .Y(new_n21205_));
  OAI21X1  g18769(.A0(new_n21205_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n21206_));
  INVX1    g18770(.A(new_n21206_), .Y(new_n21207_));
  AOI21X1  g18771(.A0(new_n21207_), .A1(new_n21200_), .B0(new_n21150_), .Y(new_n21208_));
  OAI21X1  g18772(.A0(new_n21147_), .A1(new_n12578_), .B0(new_n21146_), .Y(new_n21209_));
  MX2X1    g18773(.A(new_n21209_), .B(new_n21144_), .S0(new_n11763_), .Y(new_n21210_));
  OAI21X1  g18774(.A0(new_n21210_), .A1(pi0644), .B0(pi0715), .Y(new_n21211_));
  AOI21X1  g18775(.A0(new_n21208_), .A1(pi0644), .B0(new_n21211_), .Y(new_n21212_));
  OR3X1    g18776(.A(new_n21111_), .B(new_n12603_), .C(new_n11763_), .Y(new_n21213_));
  OAI21X1  g18777(.A0(new_n21132_), .A1(new_n12604_), .B0(new_n21213_), .Y(new_n21214_));
  OAI21X1  g18778(.A0(new_n21111_), .A1(pi0644), .B0(new_n12608_), .Y(new_n21215_));
  AOI21X1  g18779(.A0(new_n21214_), .A1(pi0644), .B0(new_n21215_), .Y(new_n21216_));
  OR2X1    g18780(.A(new_n21216_), .B(new_n11762_), .Y(new_n21217_));
  OAI21X1  g18781(.A0(new_n21210_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n21218_));
  AOI21X1  g18782(.A0(new_n21208_), .A1(new_n12612_), .B0(new_n21218_), .Y(new_n21219_));
  OAI21X1  g18783(.A0(new_n21111_), .A1(new_n12612_), .B0(pi0715), .Y(new_n21220_));
  AOI21X1  g18784(.A0(new_n21214_), .A1(new_n12612_), .B0(new_n21220_), .Y(new_n21221_));
  OR2X1    g18785(.A(new_n21221_), .B(pi1160), .Y(new_n21222_));
  OAI22X1  g18786(.A0(new_n21222_), .A1(new_n21219_), .B0(new_n21217_), .B1(new_n21212_), .Y(new_n21223_));
  NAND2X1  g18787(.A(new_n21223_), .B(pi0790), .Y(new_n21224_));
  AOI21X1  g18788(.A0(new_n21208_), .A1(new_n12766_), .B0(new_n12767_), .Y(new_n21225_));
  AOI21X1  g18789(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0193), .Y(new_n21226_));
  INVX1    g18790(.A(new_n21226_), .Y(new_n21227_));
  AOI21X1  g18791(.A0(new_n3103_), .A1(pi0690), .B0(new_n21227_), .Y(new_n21228_));
  OAI21X1  g18792(.A0(new_n12826_), .A1(new_n6885_), .B0(new_n2979_), .Y(new_n21229_));
  AOI22X1  g18793(.A0(new_n21229_), .A1(new_n3103_), .B0(new_n12825_), .B1(new_n6885_), .Y(new_n21230_));
  AOI21X1  g18794(.A0(new_n12771_), .A1(new_n6885_), .B0(new_n12441_), .Y(new_n21231_));
  NOR3X1   g18795(.A(new_n21231_), .B(new_n21230_), .C(new_n15565_), .Y(new_n21232_));
  NOR2X1   g18796(.A(new_n21232_), .B(new_n21228_), .Y(new_n21233_));
  INVX1    g18797(.A(new_n21233_), .Y(new_n21234_));
  AOI21X1  g18798(.A0(new_n21226_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n21235_));
  OAI21X1  g18799(.A0(new_n21233_), .A1(new_n12363_), .B0(new_n21235_), .Y(new_n21236_));
  AOI21X1  g18800(.A0(new_n21226_), .A1(pi0625), .B0(pi1153), .Y(new_n21237_));
  OAI21X1  g18801(.A0(new_n21233_), .A1(pi0625), .B0(new_n21237_), .Y(new_n21238_));
  AND2X1   g18802(.A(new_n21238_), .B(new_n21236_), .Y(new_n21239_));
  MX2X1    g18803(.A(new_n21239_), .B(new_n21234_), .S0(new_n11769_), .Y(new_n21240_));
  MX2X1    g18804(.A(new_n21240_), .B(new_n21226_), .S0(new_n12490_), .Y(new_n21241_));
  INVX1    g18805(.A(new_n21241_), .Y(new_n21242_));
  MX2X1    g18806(.A(new_n21242_), .B(new_n21227_), .S0(new_n12513_), .Y(new_n21243_));
  INVX1    g18807(.A(new_n21243_), .Y(new_n21244_));
  MX2X1    g18808(.A(new_n21244_), .B(new_n21226_), .S0(new_n12531_), .Y(new_n21245_));
  MX2X1    g18809(.A(new_n21245_), .B(new_n21226_), .S0(new_n12563_), .Y(new_n21246_));
  INVX1    g18810(.A(new_n21246_), .Y(new_n21247_));
  AOI21X1  g18811(.A0(new_n21226_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n21248_));
  OAI21X1  g18812(.A0(new_n21247_), .A1(new_n12554_), .B0(new_n21248_), .Y(new_n21249_));
  AOI21X1  g18813(.A0(new_n21226_), .A1(pi0628), .B0(pi1156), .Y(new_n21250_));
  OAI21X1  g18814(.A0(new_n21247_), .A1(pi0628), .B0(new_n21250_), .Y(new_n21251_));
  AOI21X1  g18815(.A0(new_n21251_), .A1(new_n21249_), .B0(new_n11764_), .Y(new_n21252_));
  AOI21X1  g18816(.A0(new_n21247_), .A1(new_n11764_), .B0(new_n21252_), .Y(new_n21253_));
  MX2X1    g18817(.A(new_n21253_), .B(new_n21226_), .S0(pi0647), .Y(new_n21254_));
  MX2X1    g18818(.A(new_n21253_), .B(new_n21226_), .S0(new_n12577_), .Y(new_n21255_));
  MX2X1    g18819(.A(new_n21255_), .B(new_n21254_), .S0(new_n12578_), .Y(new_n21256_));
  MX2X1    g18820(.A(new_n21256_), .B(new_n21253_), .S0(new_n11763_), .Y(new_n21257_));
  AOI21X1  g18821(.A0(new_n21257_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n21258_));
  OAI22X1  g18822(.A0(new_n14197_), .A1(new_n15571_), .B0(new_n12077_), .B1(pi0193), .Y(new_n21259_));
  AOI21X1  g18823(.A0(new_n16615_), .A1(pi0193), .B0(new_n15571_), .Y(new_n21260_));
  OAI21X1  g18824(.A0(new_n12776_), .A1(pi0193), .B0(new_n21260_), .Y(new_n21261_));
  OR3X1    g18825(.A(new_n12445_), .B(pi0739), .C(pi0193), .Y(new_n21262_));
  AOI21X1  g18826(.A0(new_n21262_), .A1(new_n21261_), .B0(pi0038), .Y(new_n21263_));
  AOI21X1  g18827(.A0(new_n21259_), .A1(pi0038), .B0(new_n21263_), .Y(new_n21264_));
  MX2X1    g18828(.A(new_n21264_), .B(pi0193), .S0(new_n11770_), .Y(new_n21265_));
  AND2X1   g18829(.A(new_n21265_), .B(new_n12474_), .Y(new_n21266_));
  AOI21X1  g18830(.A0(new_n21227_), .A1(new_n12473_), .B0(new_n21266_), .Y(new_n21267_));
  AOI22X1  g18831(.A0(new_n21266_), .A1(pi0609), .B0(new_n21227_), .B1(new_n12472_), .Y(new_n21268_));
  AOI22X1  g18832(.A0(new_n21266_), .A1(new_n12462_), .B0(new_n21227_), .B1(new_n12481_), .Y(new_n21269_));
  MX2X1    g18833(.A(new_n21269_), .B(new_n21268_), .S0(pi1155), .Y(new_n21270_));
  MX2X1    g18834(.A(new_n21270_), .B(new_n21267_), .S0(new_n11768_), .Y(new_n21271_));
  OAI21X1  g18835(.A0(new_n21227_), .A1(pi0618), .B0(pi1154), .Y(new_n21272_));
  AOI21X1  g18836(.A0(new_n21271_), .A1(pi0618), .B0(new_n21272_), .Y(new_n21273_));
  OAI21X1  g18837(.A0(new_n21227_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n21274_));
  AOI21X1  g18838(.A0(new_n21271_), .A1(new_n12486_), .B0(new_n21274_), .Y(new_n21275_));
  NOR2X1   g18839(.A(new_n21275_), .B(new_n21273_), .Y(new_n21276_));
  MX2X1    g18840(.A(new_n21276_), .B(new_n21271_), .S0(new_n11767_), .Y(new_n21277_));
  OAI21X1  g18841(.A0(new_n21227_), .A1(pi0619), .B0(pi1159), .Y(new_n21278_));
  AOI21X1  g18842(.A0(new_n21277_), .A1(pi0619), .B0(new_n21278_), .Y(new_n21279_));
  OAI21X1  g18843(.A0(new_n21227_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n21280_));
  AOI21X1  g18844(.A0(new_n21277_), .A1(new_n12509_), .B0(new_n21280_), .Y(new_n21281_));
  NOR2X1   g18845(.A(new_n21281_), .B(new_n21279_), .Y(new_n21282_));
  MX2X1    g18846(.A(new_n21282_), .B(new_n21277_), .S0(new_n11766_), .Y(new_n21283_));
  AND2X1   g18847(.A(new_n21226_), .B(new_n12708_), .Y(new_n21284_));
  AOI21X1  g18848(.A0(new_n21283_), .A1(new_n16140_), .B0(new_n21284_), .Y(new_n21285_));
  NAND2X1  g18849(.A(new_n21226_), .B(new_n12580_), .Y(new_n21286_));
  OAI21X1  g18850(.A0(new_n21285_), .A1(new_n12580_), .B0(new_n21286_), .Y(new_n21287_));
  MX2X1    g18851(.A(new_n21287_), .B(new_n21226_), .S0(new_n12604_), .Y(new_n21288_));
  OAI21X1  g18852(.A0(new_n21227_), .A1(pi0644), .B0(new_n12608_), .Y(new_n21289_));
  AOI21X1  g18853(.A0(new_n21288_), .A1(pi0644), .B0(new_n21289_), .Y(new_n21290_));
  OR2X1    g18854(.A(new_n21290_), .B(new_n11762_), .Y(new_n21291_));
  AOI21X1  g18855(.A0(new_n21257_), .A1(pi0644), .B0(pi0715), .Y(new_n21292_));
  OAI21X1  g18856(.A0(new_n21227_), .A1(new_n12612_), .B0(pi0715), .Y(new_n21293_));
  AOI21X1  g18857(.A0(new_n21288_), .A1(new_n12612_), .B0(new_n21293_), .Y(new_n21294_));
  OR2X1    g18858(.A(new_n21294_), .B(pi1160), .Y(new_n21295_));
  OAI22X1  g18859(.A0(new_n21295_), .A1(new_n21292_), .B0(new_n21291_), .B1(new_n21258_), .Y(new_n21296_));
  OR3X1    g18860(.A(new_n21294_), .B(pi1160), .C(pi0644), .Y(new_n21297_));
  OR3X1    g18861(.A(new_n21290_), .B(new_n11762_), .C(new_n12612_), .Y(new_n21298_));
  NAND3X1  g18862(.A(new_n21298_), .B(new_n21297_), .C(pi0790), .Y(new_n21299_));
  NAND2X1  g18863(.A(new_n21285_), .B(new_n14249_), .Y(new_n21300_));
  MX2X1    g18864(.A(new_n21251_), .B(new_n21249_), .S0(new_n12561_), .Y(new_n21301_));
  AND2X1   g18865(.A(new_n21301_), .B(new_n21300_), .Y(new_n21302_));
  OR2X1    g18866(.A(new_n21302_), .B(new_n11764_), .Y(new_n21303_));
  OR2X1    g18867(.A(new_n21264_), .B(pi0690), .Y(new_n21304_));
  OAI21X1  g18868(.A0(new_n12213_), .A1(new_n6885_), .B0(new_n15571_), .Y(new_n21305_));
  AOI21X1  g18869(.A0(new_n12155_), .A1(new_n6885_), .B0(new_n21305_), .Y(new_n21306_));
  AOI21X1  g18870(.A0(new_n12788_), .A1(new_n6885_), .B0(new_n15571_), .Y(new_n21307_));
  OAI21X1  g18871(.A0(new_n12787_), .A1(new_n6885_), .B0(new_n21307_), .Y(new_n21308_));
  NAND2X1  g18872(.A(new_n21308_), .B(pi0039), .Y(new_n21309_));
  NOR4X1   g18873(.A(new_n12340_), .B(new_n11974_), .C(new_n11967_), .D(pi0193), .Y(new_n21310_));
  OAI21X1  g18874(.A0(new_n12800_), .A1(new_n6885_), .B0(pi0739), .Y(new_n21311_));
  AND2X1   g18875(.A(new_n12332_), .B(pi0193), .Y(new_n21312_));
  OAI21X1  g18876(.A0(new_n12315_), .A1(pi0193), .B0(new_n15571_), .Y(new_n21313_));
  OAI22X1  g18877(.A0(new_n21313_), .A1(new_n21312_), .B0(new_n21311_), .B1(new_n21310_), .Y(new_n21314_));
  AOI21X1  g18878(.A0(new_n21314_), .A1(new_n2939_), .B0(pi0038), .Y(new_n21315_));
  OAI21X1  g18879(.A0(new_n21309_), .A1(new_n21306_), .B0(new_n21315_), .Y(new_n21316_));
  AOI21X1  g18880(.A0(new_n16396_), .A1(new_n15571_), .B0(new_n12276_), .Y(new_n21317_));
  OAI21X1  g18881(.A0(new_n21317_), .A1(pi0039), .B0(new_n6885_), .Y(new_n21318_));
  AOI21X1  g18882(.A0(new_n12056_), .A1(pi0739), .B0(new_n13443_), .Y(new_n21319_));
  NOR2X1   g18883(.A(new_n21319_), .B(new_n6885_), .Y(new_n21320_));
  AOI21X1  g18884(.A0(new_n21320_), .A1(new_n5782_), .B0(new_n2979_), .Y(new_n21321_));
  AOI21X1  g18885(.A0(new_n21321_), .A1(new_n21318_), .B0(new_n15565_), .Y(new_n21322_));
  AOI21X1  g18886(.A0(new_n21322_), .A1(new_n21316_), .B0(new_n11770_), .Y(new_n21323_));
  AOI22X1  g18887(.A0(new_n21323_), .A1(new_n21304_), .B0(new_n11770_), .B1(pi0193), .Y(new_n21324_));
  OAI21X1  g18888(.A0(new_n21265_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n21325_));
  AOI21X1  g18889(.A0(new_n21324_), .A1(new_n12363_), .B0(new_n21325_), .Y(new_n21326_));
  NAND2X1  g18890(.A(new_n21236_), .B(new_n12368_), .Y(new_n21327_));
  OAI21X1  g18891(.A0(new_n21265_), .A1(pi0625), .B0(pi1153), .Y(new_n21328_));
  AOI21X1  g18892(.A0(new_n21324_), .A1(pi0625), .B0(new_n21328_), .Y(new_n21329_));
  NAND2X1  g18893(.A(new_n21238_), .B(pi0608), .Y(new_n21330_));
  OAI22X1  g18894(.A0(new_n21330_), .A1(new_n21329_), .B0(new_n21327_), .B1(new_n21326_), .Y(new_n21331_));
  MX2X1    g18895(.A(new_n21331_), .B(new_n21324_), .S0(new_n11769_), .Y(new_n21332_));
  INVX1    g18896(.A(new_n21240_), .Y(new_n21333_));
  OAI21X1  g18897(.A0(new_n21333_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n21334_));
  AOI21X1  g18898(.A0(new_n21332_), .A1(new_n12462_), .B0(new_n21334_), .Y(new_n21335_));
  OAI21X1  g18899(.A0(new_n21268_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n21336_));
  OAI21X1  g18900(.A0(new_n21333_), .A1(pi0609), .B0(pi1155), .Y(new_n21337_));
  AOI21X1  g18901(.A0(new_n21332_), .A1(pi0609), .B0(new_n21337_), .Y(new_n21338_));
  OAI21X1  g18902(.A0(new_n21269_), .A1(pi1155), .B0(pi0660), .Y(new_n21339_));
  OAI22X1  g18903(.A0(new_n21339_), .A1(new_n21338_), .B0(new_n21336_), .B1(new_n21335_), .Y(new_n21340_));
  MX2X1    g18904(.A(new_n21340_), .B(new_n21332_), .S0(new_n11768_), .Y(new_n21341_));
  OAI21X1  g18905(.A0(new_n21242_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n21342_));
  AOI21X1  g18906(.A0(new_n21341_), .A1(new_n12486_), .B0(new_n21342_), .Y(new_n21343_));
  OR2X1    g18907(.A(new_n21273_), .B(pi0627), .Y(new_n21344_));
  OAI21X1  g18908(.A0(new_n21242_), .A1(pi0618), .B0(pi1154), .Y(new_n21345_));
  AOI21X1  g18909(.A0(new_n21341_), .A1(pi0618), .B0(new_n21345_), .Y(new_n21346_));
  OR2X1    g18910(.A(new_n21275_), .B(new_n12494_), .Y(new_n21347_));
  OAI22X1  g18911(.A0(new_n21347_), .A1(new_n21346_), .B0(new_n21344_), .B1(new_n21343_), .Y(new_n21348_));
  MX2X1    g18912(.A(new_n21348_), .B(new_n21341_), .S0(new_n11767_), .Y(new_n21349_));
  NAND2X1  g18913(.A(new_n21349_), .B(new_n12509_), .Y(new_n21350_));
  AOI21X1  g18914(.A0(new_n21244_), .A1(pi0619), .B0(pi1159), .Y(new_n21351_));
  OR2X1    g18915(.A(new_n21279_), .B(pi0648), .Y(new_n21352_));
  AOI21X1  g18916(.A0(new_n21351_), .A1(new_n21350_), .B0(new_n21352_), .Y(new_n21353_));
  NAND2X1  g18917(.A(new_n21349_), .B(pi0619), .Y(new_n21354_));
  AOI21X1  g18918(.A0(new_n21244_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n21355_));
  OR2X1    g18919(.A(new_n21281_), .B(new_n12517_), .Y(new_n21356_));
  AOI21X1  g18920(.A0(new_n21355_), .A1(new_n21354_), .B0(new_n21356_), .Y(new_n21357_));
  NOR3X1   g18921(.A(new_n21357_), .B(new_n21353_), .C(new_n11766_), .Y(new_n21358_));
  OAI21X1  g18922(.A0(new_n21349_), .A1(pi0789), .B0(new_n12709_), .Y(new_n21359_));
  AOI21X1  g18923(.A0(new_n21227_), .A1(pi0626), .B0(new_n16218_), .Y(new_n21360_));
  OAI21X1  g18924(.A0(new_n21283_), .A1(pi0626), .B0(new_n21360_), .Y(new_n21361_));
  AOI21X1  g18925(.A0(new_n21227_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n21362_));
  OAI21X1  g18926(.A0(new_n21283_), .A1(new_n12542_), .B0(new_n21362_), .Y(new_n21363_));
  NAND2X1  g18927(.A(new_n21245_), .B(new_n12637_), .Y(new_n21364_));
  NAND3X1  g18928(.A(new_n21364_), .B(new_n21363_), .C(new_n21361_), .Y(new_n21365_));
  AOI21X1  g18929(.A0(new_n21365_), .A1(pi0788), .B0(new_n14125_), .Y(new_n21366_));
  OAI21X1  g18930(.A0(new_n21359_), .A1(new_n21358_), .B0(new_n21366_), .Y(new_n21367_));
  AOI21X1  g18931(.A0(new_n21367_), .A1(new_n21303_), .B0(new_n14121_), .Y(new_n21368_));
  OR2X1    g18932(.A(new_n21287_), .B(new_n14239_), .Y(new_n21369_));
  OR2X1    g18933(.A(new_n21254_), .B(new_n14244_), .Y(new_n21370_));
  OR2X1    g18934(.A(new_n21255_), .B(new_n14242_), .Y(new_n21371_));
  NAND3X1  g18935(.A(new_n21371_), .B(new_n21370_), .C(new_n21369_), .Y(new_n21372_));
  AOI21X1  g18936(.A0(new_n21372_), .A1(pi0787), .B0(new_n21368_), .Y(new_n21373_));
  AOI22X1  g18937(.A0(new_n21373_), .A1(new_n21299_), .B0(new_n21296_), .B1(pi0790), .Y(new_n21374_));
  OR2X1    g18938(.A(new_n21374_), .B(po1038), .Y(new_n21375_));
  AOI21X1  g18939(.A0(po1038), .A1(new_n6885_), .B0(pi0832), .Y(new_n21376_));
  AOI22X1  g18940(.A0(new_n21376_), .A1(new_n21375_), .B0(new_n21225_), .B1(new_n21224_), .Y(po0350));
  OR2X1    g18941(.A(new_n3103_), .B(new_n11554_), .Y(new_n21378_));
  MX2X1    g18942(.A(new_n16617_), .B(new_n16611_), .S0(new_n11554_), .Y(new_n21379_));
  OAI21X1  g18943(.A0(new_n12447_), .A1(pi0194), .B0(new_n15462_), .Y(new_n21380_));
  OAI21X1  g18944(.A0(new_n21379_), .A1(new_n15462_), .B0(new_n21380_), .Y(new_n21381_));
  AOI21X1  g18945(.A0(new_n16664_), .A1(pi0194), .B0(pi0748), .Y(new_n21382_));
  OAI21X1  g18946(.A0(new_n16662_), .A1(pi0194), .B0(new_n21382_), .Y(new_n21383_));
  OAI21X1  g18947(.A0(new_n13559_), .A1(pi0194), .B0(pi0748), .Y(new_n21384_));
  AOI21X1  g18948(.A0(new_n13554_), .A1(pi0194), .B0(new_n21384_), .Y(new_n21385_));
  NOR2X1   g18949(.A(new_n21385_), .B(new_n15466_), .Y(new_n21386_));
  AOI21X1  g18950(.A0(new_n21386_), .A1(new_n21383_), .B0(new_n11770_), .Y(new_n21387_));
  OAI21X1  g18951(.A0(new_n21381_), .A1(pi0730), .B0(new_n21387_), .Y(new_n21388_));
  AND2X1   g18952(.A(new_n21388_), .B(new_n21378_), .Y(new_n21389_));
  MX2X1    g18953(.A(new_n21381_), .B(pi0194), .S0(new_n11770_), .Y(new_n21390_));
  OAI21X1  g18954(.A0(new_n21390_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n21391_));
  AOI21X1  g18955(.A0(new_n21389_), .A1(new_n12363_), .B0(new_n21391_), .Y(new_n21392_));
  OAI21X1  g18956(.A0(new_n16583_), .A1(pi0194), .B0(pi0730), .Y(new_n21393_));
  OR3X1    g18957(.A(new_n12447_), .B(pi0730), .C(pi0194), .Y(new_n21394_));
  AND3X1   g18958(.A(new_n21394_), .B(new_n21393_), .C(new_n3103_), .Y(new_n21395_));
  AOI21X1  g18959(.A0(new_n16582_), .A1(pi0194), .B0(new_n21395_), .Y(new_n21396_));
  OAI21X1  g18960(.A0(new_n12832_), .A1(new_n11770_), .B0(new_n11554_), .Y(new_n21397_));
  OAI21X1  g18961(.A0(new_n21397_), .A1(pi0625), .B0(pi1153), .Y(new_n21398_));
  AOI21X1  g18962(.A0(new_n21396_), .A1(pi0625), .B0(new_n21398_), .Y(new_n21399_));
  OR2X1    g18963(.A(new_n21399_), .B(pi0608), .Y(new_n21400_));
  OAI21X1  g18964(.A0(new_n21390_), .A1(pi0625), .B0(pi1153), .Y(new_n21401_));
  AOI21X1  g18965(.A0(new_n21389_), .A1(pi0625), .B0(new_n21401_), .Y(new_n21402_));
  OAI21X1  g18966(.A0(new_n21397_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n21403_));
  AOI21X1  g18967(.A0(new_n21396_), .A1(new_n12363_), .B0(new_n21403_), .Y(new_n21404_));
  OR2X1    g18968(.A(new_n21404_), .B(new_n12368_), .Y(new_n21405_));
  OAI22X1  g18969(.A0(new_n21405_), .A1(new_n21402_), .B0(new_n21400_), .B1(new_n21392_), .Y(new_n21406_));
  MX2X1    g18970(.A(new_n21406_), .B(new_n21389_), .S0(new_n11769_), .Y(new_n21407_));
  OAI21X1  g18971(.A0(new_n21404_), .A1(new_n21399_), .B0(pi0778), .Y(new_n21408_));
  OAI21X1  g18972(.A0(new_n21396_), .A1(pi0778), .B0(new_n21408_), .Y(new_n21409_));
  OAI21X1  g18973(.A0(new_n21409_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n21410_));
  AOI21X1  g18974(.A0(new_n21407_), .A1(new_n12462_), .B0(new_n21410_), .Y(new_n21411_));
  AND2X1   g18975(.A(new_n21390_), .B(new_n12474_), .Y(new_n21412_));
  AOI22X1  g18976(.A0(new_n21412_), .A1(pi0609), .B0(new_n21397_), .B1(new_n12472_), .Y(new_n21413_));
  OAI21X1  g18977(.A0(new_n21413_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n21414_));
  OAI21X1  g18978(.A0(new_n21409_), .A1(pi0609), .B0(pi1155), .Y(new_n21415_));
  AOI21X1  g18979(.A0(new_n21407_), .A1(pi0609), .B0(new_n21415_), .Y(new_n21416_));
  AOI22X1  g18980(.A0(new_n21412_), .A1(new_n12462_), .B0(new_n21397_), .B1(new_n12481_), .Y(new_n21417_));
  OAI21X1  g18981(.A0(new_n21417_), .A1(pi1155), .B0(pi0660), .Y(new_n21418_));
  OAI22X1  g18982(.A0(new_n21418_), .A1(new_n21416_), .B0(new_n21414_), .B1(new_n21411_), .Y(new_n21419_));
  MX2X1    g18983(.A(new_n21419_), .B(new_n21407_), .S0(new_n11768_), .Y(new_n21420_));
  MX2X1    g18984(.A(new_n21409_), .B(new_n21397_), .S0(new_n12490_), .Y(new_n21421_));
  OAI21X1  g18985(.A0(new_n21421_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n21422_));
  AOI21X1  g18986(.A0(new_n21420_), .A1(new_n12486_), .B0(new_n21422_), .Y(new_n21423_));
  AOI21X1  g18987(.A0(new_n21397_), .A1(new_n12473_), .B0(new_n21412_), .Y(new_n21424_));
  MX2X1    g18988(.A(new_n21417_), .B(new_n21413_), .S0(pi1155), .Y(new_n21425_));
  MX2X1    g18989(.A(new_n21425_), .B(new_n21424_), .S0(new_n11768_), .Y(new_n21426_));
  OAI21X1  g18990(.A0(new_n21397_), .A1(pi0618), .B0(pi1154), .Y(new_n21427_));
  AOI21X1  g18991(.A0(new_n21426_), .A1(pi0618), .B0(new_n21427_), .Y(new_n21428_));
  OR2X1    g18992(.A(new_n21428_), .B(pi0627), .Y(new_n21429_));
  OAI21X1  g18993(.A0(new_n21421_), .A1(pi0618), .B0(pi1154), .Y(new_n21430_));
  AOI21X1  g18994(.A0(new_n21420_), .A1(pi0618), .B0(new_n21430_), .Y(new_n21431_));
  OAI21X1  g18995(.A0(new_n21397_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n21432_));
  AOI21X1  g18996(.A0(new_n21426_), .A1(new_n12486_), .B0(new_n21432_), .Y(new_n21433_));
  OR2X1    g18997(.A(new_n21433_), .B(new_n12494_), .Y(new_n21434_));
  OAI22X1  g18998(.A0(new_n21434_), .A1(new_n21431_), .B0(new_n21429_), .B1(new_n21423_), .Y(new_n21435_));
  MX2X1    g18999(.A(new_n21435_), .B(new_n21420_), .S0(new_n11767_), .Y(new_n21436_));
  MX2X1    g19000(.A(new_n21421_), .B(new_n21397_), .S0(new_n12513_), .Y(new_n21437_));
  OAI21X1  g19001(.A0(new_n21437_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n21438_));
  AOI21X1  g19002(.A0(new_n21436_), .A1(new_n12509_), .B0(new_n21438_), .Y(new_n21439_));
  NOR2X1   g19003(.A(new_n21433_), .B(new_n21428_), .Y(new_n21440_));
  MX2X1    g19004(.A(new_n21440_), .B(new_n21426_), .S0(new_n11767_), .Y(new_n21441_));
  OAI21X1  g19005(.A0(new_n21397_), .A1(pi0619), .B0(pi1159), .Y(new_n21442_));
  AOI21X1  g19006(.A0(new_n21441_), .A1(pi0619), .B0(new_n21442_), .Y(new_n21443_));
  OR2X1    g19007(.A(new_n21443_), .B(pi0648), .Y(new_n21444_));
  OAI21X1  g19008(.A0(new_n21437_), .A1(pi0619), .B0(pi1159), .Y(new_n21445_));
  AOI21X1  g19009(.A0(new_n21436_), .A1(pi0619), .B0(new_n21445_), .Y(new_n21446_));
  OAI21X1  g19010(.A0(new_n21397_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n21447_));
  AOI21X1  g19011(.A0(new_n21441_), .A1(new_n12509_), .B0(new_n21447_), .Y(new_n21448_));
  OR2X1    g19012(.A(new_n21448_), .B(new_n12517_), .Y(new_n21449_));
  OAI22X1  g19013(.A0(new_n21449_), .A1(new_n21446_), .B0(new_n21444_), .B1(new_n21439_), .Y(new_n21450_));
  MX2X1    g19014(.A(new_n21450_), .B(new_n21436_), .S0(new_n11766_), .Y(new_n21451_));
  MX2X1    g19015(.A(new_n21437_), .B(new_n21397_), .S0(new_n12531_), .Y(new_n21452_));
  AOI21X1  g19016(.A0(new_n21452_), .A1(pi0626), .B0(pi0641), .Y(new_n21453_));
  OAI21X1  g19017(.A0(new_n21451_), .A1(pi0626), .B0(new_n21453_), .Y(new_n21454_));
  OR2X1    g19018(.A(new_n21441_), .B(pi0789), .Y(new_n21455_));
  OAI21X1  g19019(.A0(new_n21448_), .A1(new_n21443_), .B0(pi0789), .Y(new_n21456_));
  NAND2X1  g19020(.A(new_n21456_), .B(new_n21455_), .Y(new_n21457_));
  NAND2X1  g19021(.A(new_n21457_), .B(new_n12542_), .Y(new_n21458_));
  AOI21X1  g19022(.A0(new_n21397_), .A1(pi0626), .B0(new_n12543_), .Y(new_n21459_));
  AOI21X1  g19023(.A0(new_n21459_), .A1(new_n21458_), .B0(pi1158), .Y(new_n21460_));
  AOI21X1  g19024(.A0(new_n21452_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n21461_));
  OAI21X1  g19025(.A0(new_n21451_), .A1(new_n12542_), .B0(new_n21461_), .Y(new_n21462_));
  NAND2X1  g19026(.A(new_n21457_), .B(pi0626), .Y(new_n21463_));
  AOI21X1  g19027(.A0(new_n21397_), .A1(new_n12542_), .B0(pi0641), .Y(new_n21464_));
  AOI21X1  g19028(.A0(new_n21464_), .A1(new_n21463_), .B0(new_n12548_), .Y(new_n21465_));
  AOI22X1  g19029(.A0(new_n21465_), .A1(new_n21462_), .B0(new_n21460_), .B1(new_n21454_), .Y(new_n21466_));
  MX2X1    g19030(.A(new_n21466_), .B(new_n21451_), .S0(new_n11765_), .Y(new_n21467_));
  MX2X1    g19031(.A(new_n21457_), .B(new_n21397_), .S0(new_n12708_), .Y(new_n21468_));
  OAI21X1  g19032(.A0(new_n21468_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n21469_));
  AOI21X1  g19033(.A0(new_n21467_), .A1(new_n12554_), .B0(new_n21469_), .Y(new_n21470_));
  MX2X1    g19034(.A(new_n21452_), .B(new_n21397_), .S0(new_n12563_), .Y(new_n21471_));
  INVX1    g19035(.A(new_n21397_), .Y(new_n21472_));
  AOI21X1  g19036(.A0(new_n21472_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n21473_));
  OAI21X1  g19037(.A0(new_n21471_), .A1(new_n12554_), .B0(new_n21473_), .Y(new_n21474_));
  AND2X1   g19038(.A(new_n21474_), .B(new_n12561_), .Y(new_n21475_));
  INVX1    g19039(.A(new_n21475_), .Y(new_n21476_));
  OAI21X1  g19040(.A0(new_n21468_), .A1(pi0628), .B0(pi1156), .Y(new_n21477_));
  AOI21X1  g19041(.A0(new_n21467_), .A1(pi0628), .B0(new_n21477_), .Y(new_n21478_));
  AOI21X1  g19042(.A0(new_n21472_), .A1(pi0628), .B0(pi1156), .Y(new_n21479_));
  OAI21X1  g19043(.A0(new_n21471_), .A1(pi0628), .B0(new_n21479_), .Y(new_n21480_));
  AND2X1   g19044(.A(new_n21480_), .B(pi0629), .Y(new_n21481_));
  INVX1    g19045(.A(new_n21481_), .Y(new_n21482_));
  OAI22X1  g19046(.A0(new_n21482_), .A1(new_n21478_), .B0(new_n21476_), .B1(new_n21470_), .Y(new_n21483_));
  AND2X1   g19047(.A(new_n21467_), .B(new_n11764_), .Y(new_n21484_));
  AOI21X1  g19048(.A0(new_n21483_), .A1(pi0792), .B0(new_n21484_), .Y(new_n21485_));
  MX2X1    g19049(.A(new_n21468_), .B(new_n21397_), .S0(new_n12580_), .Y(new_n21486_));
  INVX1    g19050(.A(new_n21486_), .Y(new_n21487_));
  AOI21X1  g19051(.A0(new_n21487_), .A1(pi0647), .B0(pi1157), .Y(new_n21488_));
  OAI21X1  g19052(.A0(new_n21485_), .A1(pi0647), .B0(new_n21488_), .Y(new_n21489_));
  AOI21X1  g19053(.A0(new_n21480_), .A1(new_n21474_), .B0(new_n11764_), .Y(new_n21490_));
  AOI21X1  g19054(.A0(new_n21471_), .A1(new_n11764_), .B0(new_n21490_), .Y(new_n21491_));
  OAI21X1  g19055(.A0(new_n21397_), .A1(pi0647), .B0(pi1157), .Y(new_n21492_));
  AOI21X1  g19056(.A0(new_n21491_), .A1(pi0647), .B0(new_n21492_), .Y(new_n21493_));
  NOR2X1   g19057(.A(new_n21493_), .B(pi0630), .Y(new_n21494_));
  AOI21X1  g19058(.A0(new_n21487_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n21495_));
  OAI21X1  g19059(.A0(new_n21485_), .A1(new_n12577_), .B0(new_n21495_), .Y(new_n21496_));
  OAI21X1  g19060(.A0(new_n21397_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n21497_));
  AOI21X1  g19061(.A0(new_n21491_), .A1(new_n12577_), .B0(new_n21497_), .Y(new_n21498_));
  NOR2X1   g19062(.A(new_n21498_), .B(new_n12592_), .Y(new_n21499_));
  AOI22X1  g19063(.A0(new_n21499_), .A1(new_n21496_), .B0(new_n21494_), .B1(new_n21489_), .Y(new_n21500_));
  OR2X1    g19064(.A(new_n21485_), .B(pi0787), .Y(new_n21501_));
  OAI21X1  g19065(.A0(new_n21500_), .A1(new_n11763_), .B0(new_n21501_), .Y(new_n21502_));
  OAI21X1  g19066(.A0(new_n21498_), .A1(new_n21493_), .B0(pi0787), .Y(new_n21503_));
  OAI21X1  g19067(.A0(new_n21491_), .A1(pi0787), .B0(new_n21503_), .Y(new_n21504_));
  OAI21X1  g19068(.A0(new_n21504_), .A1(pi0644), .B0(pi0715), .Y(new_n21505_));
  AOI21X1  g19069(.A0(new_n21502_), .A1(pi0644), .B0(new_n21505_), .Y(new_n21506_));
  MX2X1    g19070(.A(new_n21487_), .B(new_n21472_), .S0(new_n12604_), .Y(new_n21507_));
  OAI21X1  g19071(.A0(new_n21397_), .A1(pi0644), .B0(new_n12608_), .Y(new_n21508_));
  AOI21X1  g19072(.A0(new_n21507_), .A1(pi0644), .B0(new_n21508_), .Y(new_n21509_));
  NOR3X1   g19073(.A(new_n21509_), .B(new_n21506_), .C(new_n11762_), .Y(new_n21510_));
  OAI21X1  g19074(.A0(new_n21504_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n21511_));
  AOI21X1  g19075(.A0(new_n21502_), .A1(new_n12612_), .B0(new_n21511_), .Y(new_n21512_));
  OAI21X1  g19076(.A0(new_n21397_), .A1(new_n12612_), .B0(pi0715), .Y(new_n21513_));
  AOI21X1  g19077(.A0(new_n21507_), .A1(new_n12612_), .B0(new_n21513_), .Y(new_n21514_));
  OR2X1    g19078(.A(new_n21514_), .B(pi1160), .Y(new_n21515_));
  OAI21X1  g19079(.A0(new_n21515_), .A1(new_n21512_), .B0(pi0790), .Y(new_n21516_));
  MX2X1    g19080(.A(new_n21500_), .B(new_n21485_), .S0(new_n11763_), .Y(new_n21517_));
  AOI21X1  g19081(.A0(new_n21517_), .A1(new_n12766_), .B0(po1038), .Y(new_n21518_));
  OAI21X1  g19082(.A0(new_n21516_), .A1(new_n21510_), .B0(new_n21518_), .Y(new_n21519_));
  AOI21X1  g19083(.A0(po1038), .A1(new_n11554_), .B0(pi0832), .Y(new_n21520_));
  AOI21X1  g19084(.A0(pi1093), .A1(pi1092), .B0(pi0194), .Y(new_n21521_));
  INVX1    g19085(.A(new_n21521_), .Y(new_n21522_));
  AOI21X1  g19086(.A0(new_n12056_), .A1(pi0748), .B0(new_n21521_), .Y(new_n21523_));
  AOI21X1  g19087(.A0(new_n12473_), .A1(new_n2720_), .B0(new_n21523_), .Y(new_n21524_));
  INVX1    g19088(.A(new_n21523_), .Y(new_n21525_));
  AOI21X1  g19089(.A0(new_n21525_), .A1(new_n14331_), .B0(new_n12463_), .Y(new_n21526_));
  AOI21X1  g19090(.A0(new_n21524_), .A1(new_n12646_), .B0(pi1155), .Y(new_n21527_));
  OAI21X1  g19091(.A0(new_n21527_), .A1(new_n21526_), .B0(pi0785), .Y(new_n21528_));
  OAI21X1  g19092(.A0(new_n21524_), .A1(pi0785), .B0(new_n21528_), .Y(new_n21529_));
  INVX1    g19093(.A(new_n21529_), .Y(new_n21530_));
  AOI21X1  g19094(.A0(new_n21530_), .A1(new_n12652_), .B0(new_n12487_), .Y(new_n21531_));
  AOI21X1  g19095(.A0(new_n21530_), .A1(new_n12655_), .B0(pi1154), .Y(new_n21532_));
  NOR2X1   g19096(.A(new_n21532_), .B(new_n21531_), .Y(new_n21533_));
  MX2X1    g19097(.A(new_n21533_), .B(new_n21530_), .S0(new_n11767_), .Y(new_n21534_));
  NOR2X1   g19098(.A(new_n21534_), .B(pi0789), .Y(new_n21535_));
  INVX1    g19099(.A(new_n21534_), .Y(new_n21536_));
  AOI21X1  g19100(.A0(new_n21521_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n21537_));
  OAI21X1  g19101(.A0(new_n21536_), .A1(new_n12509_), .B0(new_n21537_), .Y(new_n21538_));
  AOI21X1  g19102(.A0(new_n21521_), .A1(pi0619), .B0(pi1159), .Y(new_n21539_));
  OAI21X1  g19103(.A0(new_n21536_), .A1(pi0619), .B0(new_n21539_), .Y(new_n21540_));
  AOI21X1  g19104(.A0(new_n21540_), .A1(new_n21538_), .B0(new_n11766_), .Y(new_n21541_));
  NOR2X1   g19105(.A(new_n21541_), .B(new_n21535_), .Y(new_n21542_));
  INVX1    g19106(.A(new_n21542_), .Y(new_n21543_));
  MX2X1    g19107(.A(new_n21543_), .B(new_n21522_), .S0(new_n12708_), .Y(new_n21544_));
  MX2X1    g19108(.A(new_n21544_), .B(new_n21522_), .S0(new_n12580_), .Y(new_n21545_));
  AOI21X1  g19109(.A0(new_n12439_), .A1(pi0730), .B0(new_n21521_), .Y(new_n21546_));
  AND3X1   g19110(.A(new_n12439_), .B(pi0730), .C(new_n12363_), .Y(new_n21547_));
  NOR2X1   g19111(.A(new_n21547_), .B(new_n21546_), .Y(new_n21548_));
  NOR2X1   g19112(.A(new_n21521_), .B(pi1153), .Y(new_n21549_));
  INVX1    g19113(.A(new_n21549_), .Y(new_n21550_));
  OAI22X1  g19114(.A0(new_n21550_), .A1(new_n21547_), .B0(new_n21548_), .B1(new_n12364_), .Y(new_n21551_));
  MX2X1    g19115(.A(new_n21551_), .B(new_n21546_), .S0(new_n11769_), .Y(new_n21552_));
  NOR4X1   g19116(.A(new_n21552_), .B(new_n12633_), .C(new_n12631_), .D(new_n12630_), .Y(new_n21553_));
  AND3X1   g19117(.A(new_n21553_), .B(new_n12739_), .C(new_n12718_), .Y(new_n21554_));
  INVX1    g19118(.A(new_n21554_), .Y(new_n21555_));
  AOI21X1  g19119(.A0(new_n21521_), .A1(pi0647), .B0(pi1157), .Y(new_n21556_));
  OAI21X1  g19120(.A0(new_n21555_), .A1(pi0647), .B0(new_n21556_), .Y(new_n21557_));
  MX2X1    g19121(.A(new_n21554_), .B(new_n21521_), .S0(new_n12577_), .Y(new_n21558_));
  OAI22X1  g19122(.A0(new_n21558_), .A1(new_n14242_), .B0(new_n21557_), .B1(new_n12592_), .Y(new_n21559_));
  AOI21X1  g19123(.A0(new_n21545_), .A1(new_n14326_), .B0(new_n21559_), .Y(new_n21560_));
  AOI21X1  g19124(.A0(new_n21522_), .A1(pi0626), .B0(new_n16218_), .Y(new_n21561_));
  OAI21X1  g19125(.A0(new_n21542_), .A1(pi0626), .B0(new_n21561_), .Y(new_n21562_));
  AOI21X1  g19126(.A0(new_n21522_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n21563_));
  OAI21X1  g19127(.A0(new_n21542_), .A1(new_n12542_), .B0(new_n21563_), .Y(new_n21564_));
  NAND2X1  g19128(.A(new_n21553_), .B(new_n12637_), .Y(new_n21565_));
  AND3X1   g19129(.A(new_n21565_), .B(new_n21564_), .C(new_n21562_), .Y(new_n21566_));
  NOR2X1   g19130(.A(new_n21566_), .B(new_n11765_), .Y(new_n21567_));
  INVX1    g19131(.A(new_n21567_), .Y(new_n21568_));
  NOR2X1   g19132(.A(new_n21546_), .B(new_n11991_), .Y(new_n21569_));
  MX2X1    g19133(.A(new_n21525_), .B(new_n12363_), .S0(new_n21569_), .Y(new_n21570_));
  NOR2X1   g19134(.A(new_n21570_), .B(new_n21550_), .Y(new_n21571_));
  OAI21X1  g19135(.A0(new_n21548_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n21572_));
  NOR2X1   g19136(.A(new_n21572_), .B(new_n21571_), .Y(new_n21573_));
  OR3X1    g19137(.A(new_n21546_), .B(new_n11991_), .C(new_n12363_), .Y(new_n21574_));
  AND2X1   g19138(.A(new_n21523_), .B(pi1153), .Y(new_n21575_));
  OAI21X1  g19139(.A0(new_n21550_), .A1(new_n21547_), .B0(pi0608), .Y(new_n21576_));
  AOI21X1  g19140(.A0(new_n21575_), .A1(new_n21574_), .B0(new_n21576_), .Y(new_n21577_));
  OAI21X1  g19141(.A0(new_n21577_), .A1(new_n21573_), .B0(pi0778), .Y(new_n21578_));
  OAI21X1  g19142(.A0(new_n21569_), .A1(new_n21525_), .B0(new_n11769_), .Y(new_n21579_));
  NAND2X1  g19143(.A(new_n21579_), .B(new_n21578_), .Y(new_n21580_));
  INVX1    g19144(.A(new_n21580_), .Y(new_n21581_));
  OAI21X1  g19145(.A0(new_n21552_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n21582_));
  AOI21X1  g19146(.A0(new_n21580_), .A1(new_n12462_), .B0(new_n21582_), .Y(new_n21583_));
  NOR3X1   g19147(.A(new_n21583_), .B(new_n21526_), .C(pi0660), .Y(new_n21584_));
  OAI21X1  g19148(.A0(new_n21552_), .A1(pi0609), .B0(pi1155), .Y(new_n21585_));
  AOI21X1  g19149(.A0(new_n21580_), .A1(pi0609), .B0(new_n21585_), .Y(new_n21586_));
  NOR3X1   g19150(.A(new_n21586_), .B(new_n21527_), .C(new_n12468_), .Y(new_n21587_));
  NOR2X1   g19151(.A(new_n21587_), .B(new_n21584_), .Y(new_n21588_));
  MX2X1    g19152(.A(new_n21588_), .B(new_n21581_), .S0(new_n11768_), .Y(new_n21589_));
  OR3X1    g19153(.A(new_n21552_), .B(new_n12630_), .C(new_n12486_), .Y(new_n21590_));
  AND2X1   g19154(.A(new_n21590_), .B(new_n12487_), .Y(new_n21591_));
  OAI21X1  g19155(.A0(new_n21589_), .A1(pi0618), .B0(new_n21591_), .Y(new_n21592_));
  NOR2X1   g19156(.A(new_n21531_), .B(pi0627), .Y(new_n21593_));
  NOR3X1   g19157(.A(new_n21552_), .B(new_n12630_), .C(pi0618), .Y(new_n21594_));
  NOR2X1   g19158(.A(new_n21594_), .B(new_n12487_), .Y(new_n21595_));
  OAI21X1  g19159(.A0(new_n21589_), .A1(new_n12486_), .B0(new_n21595_), .Y(new_n21596_));
  NOR2X1   g19160(.A(new_n21532_), .B(new_n12494_), .Y(new_n21597_));
  AOI22X1  g19161(.A0(new_n21597_), .A1(new_n21596_), .B0(new_n21593_), .B1(new_n21592_), .Y(new_n21598_));
  MX2X1    g19162(.A(new_n21598_), .B(new_n21589_), .S0(new_n11767_), .Y(new_n21599_));
  OR4X1    g19163(.A(new_n21552_), .B(new_n12631_), .C(new_n12630_), .D(new_n12509_), .Y(new_n21600_));
  AND2X1   g19164(.A(new_n21600_), .B(new_n12510_), .Y(new_n21601_));
  OAI21X1  g19165(.A0(new_n21599_), .A1(pi0619), .B0(new_n21601_), .Y(new_n21602_));
  AND3X1   g19166(.A(new_n21602_), .B(new_n21538_), .C(new_n12517_), .Y(new_n21603_));
  NOR4X1   g19167(.A(new_n21552_), .B(new_n12631_), .C(new_n12630_), .D(pi0619), .Y(new_n21604_));
  NOR2X1   g19168(.A(new_n21604_), .B(new_n12510_), .Y(new_n21605_));
  OAI21X1  g19169(.A0(new_n21599_), .A1(new_n12509_), .B0(new_n21605_), .Y(new_n21606_));
  AND2X1   g19170(.A(new_n21540_), .B(pi0648), .Y(new_n21607_));
  AOI21X1  g19171(.A0(new_n21607_), .A1(new_n21606_), .B0(new_n11766_), .Y(new_n21608_));
  INVX1    g19172(.A(new_n21608_), .Y(new_n21609_));
  AOI21X1  g19173(.A0(new_n21599_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n21610_));
  OAI21X1  g19174(.A0(new_n21609_), .A1(new_n21603_), .B0(new_n21610_), .Y(new_n21611_));
  AOI21X1  g19175(.A0(new_n21611_), .A1(new_n21568_), .B0(new_n14125_), .Y(new_n21612_));
  INVX1    g19176(.A(new_n21544_), .Y(new_n21613_));
  AND2X1   g19177(.A(new_n21553_), .B(new_n12718_), .Y(new_n21614_));
  AOI22X1  g19178(.A0(new_n21614_), .A1(new_n14426_), .B0(new_n21613_), .B1(new_n12735_), .Y(new_n21615_));
  AOI22X1  g19179(.A0(new_n21614_), .A1(new_n14428_), .B0(new_n21613_), .B1(new_n12733_), .Y(new_n21616_));
  MX2X1    g19180(.A(new_n21616_), .B(new_n21615_), .S0(new_n12561_), .Y(new_n21617_));
  OAI21X1  g19181(.A0(new_n21617_), .A1(new_n11764_), .B0(new_n14122_), .Y(new_n21618_));
  OAI22X1  g19182(.A0(new_n21618_), .A1(new_n21612_), .B0(new_n21560_), .B1(new_n11763_), .Y(new_n21619_));
  INVX1    g19183(.A(new_n21619_), .Y(new_n21620_));
  OAI21X1  g19184(.A0(new_n21558_), .A1(new_n12578_), .B0(new_n21557_), .Y(new_n21621_));
  MX2X1    g19185(.A(new_n21621_), .B(new_n21555_), .S0(new_n11763_), .Y(new_n21622_));
  OAI21X1  g19186(.A0(new_n21622_), .A1(pi0644), .B0(pi0715), .Y(new_n21623_));
  AOI21X1  g19187(.A0(new_n21620_), .A1(pi0644), .B0(new_n21623_), .Y(new_n21624_));
  OR3X1    g19188(.A(new_n21522_), .B(new_n12603_), .C(new_n11763_), .Y(new_n21625_));
  OAI21X1  g19189(.A0(new_n21545_), .A1(new_n12604_), .B0(new_n21625_), .Y(new_n21626_));
  OAI21X1  g19190(.A0(new_n21522_), .A1(pi0644), .B0(new_n12608_), .Y(new_n21627_));
  AOI21X1  g19191(.A0(new_n21626_), .A1(pi0644), .B0(new_n21627_), .Y(new_n21628_));
  OR2X1    g19192(.A(new_n21628_), .B(new_n11762_), .Y(new_n21629_));
  OAI21X1  g19193(.A0(new_n21622_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n21630_));
  AOI21X1  g19194(.A0(new_n21620_), .A1(new_n12612_), .B0(new_n21630_), .Y(new_n21631_));
  OAI21X1  g19195(.A0(new_n21522_), .A1(new_n12612_), .B0(pi0715), .Y(new_n21632_));
  AOI21X1  g19196(.A0(new_n21626_), .A1(new_n12612_), .B0(new_n21632_), .Y(new_n21633_));
  OR2X1    g19197(.A(new_n21633_), .B(pi1160), .Y(new_n21634_));
  OAI22X1  g19198(.A0(new_n21634_), .A1(new_n21631_), .B0(new_n21629_), .B1(new_n21624_), .Y(new_n21635_));
  OAI21X1  g19199(.A0(new_n21619_), .A1(pi0790), .B0(pi0832), .Y(new_n21636_));
  AOI21X1  g19200(.A0(new_n21635_), .A1(pi0790), .B0(new_n21636_), .Y(new_n21637_));
  AOI21X1  g19201(.A0(new_n21520_), .A1(new_n21519_), .B0(new_n21637_), .Y(po0351));
  NAND2X1  g19202(.A(pi0299), .B(pi0171), .Y(new_n21639_));
  OAI21X1  g19203(.A0(new_n21639_), .A1(new_n6255_), .B0(new_n8491_), .Y(new_n21640_));
  OAI22X1  g19204(.A0(new_n11716_), .A1(new_n11459_), .B0(new_n11475_), .B1(new_n8489_), .Y(new_n21641_));
  OAI21X1  g19205(.A0(new_n21641_), .A1(new_n21640_), .B0(pi0232), .Y(new_n21642_));
  AOI21X1  g19206(.A0(new_n21642_), .A1(new_n11714_), .B0(new_n2939_), .Y(new_n21643_));
  AOI21X1  g19207(.A0(new_n11514_), .A1(new_n6819_), .B0(new_n9999_), .Y(new_n21644_));
  AND2X1   g19208(.A(new_n11724_), .B(new_n11666_), .Y(new_n21645_));
  INVX1    g19209(.A(new_n21645_), .Y(new_n21646_));
  OAI21X1  g19210(.A0(new_n21646_), .A1(pi0196), .B0(pi0195), .Y(new_n21647_));
  AND2X1   g19211(.A(new_n21647_), .B(new_n7628_), .Y(new_n21648_));
  OAI21X1  g19212(.A0(new_n21644_), .A1(pi0039), .B0(new_n21648_), .Y(new_n21649_));
  OR3X1    g19213(.A(new_n11678_), .B(pi0299), .C(new_n11458_), .Y(new_n21650_));
  OAI22X1  g19214(.A0(new_n11465_), .A1(new_n11680_), .B0(new_n11682_), .B1(new_n3715_), .Y(new_n21651_));
  OAI21X1  g19215(.A0(new_n11685_), .A1(pi0192), .B0(pi0232), .Y(new_n21652_));
  AOI21X1  g19216(.A0(new_n21651_), .A1(pi0299), .B0(new_n21652_), .Y(new_n21653_));
  AOI21X1  g19217(.A0(new_n21653_), .A1(new_n21650_), .B0(new_n11675_), .Y(new_n21654_));
  OAI22X1  g19218(.A0(new_n11692_), .A1(new_n11697_), .B0(new_n11689_), .B1(pi0171), .Y(new_n21655_));
  AOI21X1  g19219(.A0(new_n21655_), .A1(new_n6856_), .B0(new_n8800_), .Y(new_n21656_));
  MX2X1    g19220(.A(new_n11701_), .B(new_n11691_), .S0(new_n11458_), .Y(new_n21657_));
  OAI21X1  g19221(.A0(new_n21657_), .A1(new_n21656_), .B0(pi0232), .Y(new_n21658_));
  AOI21X1  g19222(.A0(new_n21658_), .A1(new_n11696_), .B0(new_n2939_), .Y(new_n21659_));
  OR2X1    g19223(.A(new_n21659_), .B(new_n3252_), .Y(new_n21660_));
  OAI21X1  g19224(.A0(new_n21660_), .A1(new_n21654_), .B0(new_n3131_), .Y(new_n21661_));
  AOI21X1  g19225(.A0(new_n21661_), .A1(new_n11670_), .B0(pi0092), .Y(new_n21662_));
  OAI21X1  g19226(.A0(new_n21662_), .A1(new_n11669_), .B0(new_n3107_), .Y(new_n21663_));
  AOI21X1  g19227(.A0(new_n21663_), .A1(new_n11710_), .B0(new_n4975_), .Y(new_n21664_));
  OR2X1    g19228(.A(new_n21647_), .B(new_n9836_), .Y(new_n21665_));
  OAI22X1  g19229(.A0(new_n21665_), .A1(new_n21664_), .B0(new_n21649_), .B1(new_n21643_), .Y(po0352));
  INVX1    g19230(.A(pi0196), .Y(new_n21667_));
  INVX1    g19231(.A(new_n11710_), .Y(new_n21668_));
  INVX1    g19232(.A(new_n11669_), .Y(new_n21669_));
  INVX1    g19233(.A(new_n11670_), .Y(new_n21670_));
  OAI22X1  g19234(.A0(new_n11692_), .A1(new_n11697_), .B0(new_n11689_), .B1(pi0170), .Y(new_n21671_));
  AOI21X1  g19235(.A0(new_n21671_), .A1(new_n6856_), .B0(new_n8800_), .Y(new_n21672_));
  OAI21X1  g19236(.A0(new_n21672_), .A1(new_n11691_), .B0(pi0232), .Y(new_n21673_));
  NAND2X1  g19237(.A(new_n21673_), .B(new_n11696_), .Y(new_n21674_));
  AOI21X1  g19238(.A0(new_n11701_), .A1(pi0232), .B0(new_n21674_), .Y(new_n21675_));
  AND2X1   g19239(.A(pi0194), .B(new_n2979_), .Y(new_n21676_));
  OAI21X1  g19240(.A0(new_n21675_), .A1(new_n2939_), .B0(new_n21676_), .Y(new_n21677_));
  INVX1    g19241(.A(new_n21677_), .Y(new_n21678_));
  AOI21X1  g19242(.A0(new_n21673_), .A1(new_n11696_), .B0(new_n2939_), .Y(new_n21679_));
  NOR3X1   g19243(.A(new_n21679_), .B(pi0194), .C(pi0038), .Y(new_n21680_));
  OAI22X1  g19244(.A0(new_n21680_), .A1(new_n21678_), .B0(new_n11673_), .B1(pi0039), .Y(new_n21681_));
  OR2X1    g19245(.A(new_n11678_), .B(pi0299), .Y(new_n21682_));
  AOI22X1  g19246(.A0(new_n21680_), .A1(new_n11685_), .B0(new_n21678_), .B1(new_n21682_), .Y(new_n21683_));
  AOI21X1  g19247(.A0(new_n7089_), .A1(new_n7063_), .B0(new_n11531_), .Y(new_n21684_));
  AOI21X1  g19248(.A0(new_n11681_), .A1(pi0170), .B0(new_n21684_), .Y(new_n21685_));
  OAI21X1  g19249(.A0(new_n21685_), .A1(new_n2933_), .B0(pi0232), .Y(new_n21686_));
  OAI21X1  g19250(.A0(new_n21686_), .A1(new_n21683_), .B0(new_n21681_), .Y(new_n21687_));
  AOI21X1  g19251(.A0(new_n21687_), .A1(new_n3007_), .B0(pi0087), .Y(new_n21688_));
  OAI21X1  g19252(.A0(new_n21688_), .A1(new_n21670_), .B0(new_n3079_), .Y(new_n21689_));
  AOI21X1  g19253(.A0(new_n21689_), .A1(new_n21669_), .B0(pi0055), .Y(new_n21690_));
  OAI21X1  g19254(.A0(new_n21690_), .A1(new_n21668_), .B0(new_n3123_), .Y(new_n21691_));
  AOI21X1  g19255(.A0(new_n21691_), .A1(new_n7323_), .B0(new_n21667_), .Y(new_n21692_));
  AOI21X1  g19256(.A0(new_n7189_), .A1(new_n3865_), .B0(new_n11715_), .Y(new_n21693_));
  NOR4X1   g19257(.A(new_n21693_), .B(new_n4890_), .C(new_n2437_), .D(new_n2438_), .Y(new_n21694_));
  AND2X1   g19258(.A(new_n11715_), .B(new_n9494_), .Y(new_n21695_));
  NOR3X1   g19259(.A(new_n21695_), .B(new_n21694_), .C(new_n5215_), .Y(new_n21696_));
  AOI21X1  g19260(.A0(new_n8492_), .A1(new_n5215_), .B0(new_n21696_), .Y(new_n21697_));
  MX2X1    g19261(.A(new_n21697_), .B(new_n8489_), .S0(new_n2933_), .Y(new_n21698_));
  OR3X1    g19262(.A(new_n11525_), .B(new_n7251_), .C(new_n7619_), .Y(new_n21699_));
  AOI21X1  g19263(.A0(new_n21699_), .A1(new_n2939_), .B0(pi0038), .Y(new_n21700_));
  OAI21X1  g19264(.A0(new_n21698_), .A1(new_n2939_), .B0(new_n21700_), .Y(new_n21701_));
  NOR2X1   g19265(.A(new_n21697_), .B(new_n2939_), .Y(new_n21702_));
  NOR4X1   g19266(.A(new_n11564_), .B(new_n7251_), .C(new_n6827_), .D(new_n7619_), .Y(new_n21703_));
  OAI21X1  g19267(.A0(new_n21703_), .A1(pi0039), .B0(new_n2979_), .Y(new_n21704_));
  OAI21X1  g19268(.A0(new_n21704_), .A1(new_n21702_), .B0(pi0194), .Y(new_n21705_));
  NAND2X1  g19269(.A(new_n21705_), .B(new_n7625_), .Y(new_n21706_));
  AOI21X1  g19270(.A0(new_n21701_), .A1(new_n11554_), .B0(new_n21706_), .Y(new_n21707_));
  OAI21X1  g19271(.A0(new_n21707_), .A1(pi0196), .B0(new_n21646_), .Y(new_n21708_));
  AND2X1   g19272(.A(new_n21667_), .B(pi0195), .Y(new_n21709_));
  INVX1    g19273(.A(new_n21709_), .Y(new_n21710_));
  AOI21X1  g19274(.A0(new_n21691_), .A1(new_n7323_), .B0(new_n21710_), .Y(new_n21711_));
  OAI21X1  g19275(.A0(new_n21709_), .A1(new_n21707_), .B0(new_n21645_), .Y(new_n21712_));
  OAI22X1  g19276(.A0(new_n21712_), .A1(new_n21711_), .B0(new_n21708_), .B1(new_n21692_), .Y(po0353));
  AND2X1   g19277(.A(pi0947), .B(new_n14191_), .Y(new_n21714_));
  INVX1    g19278(.A(new_n21714_), .Y(new_n21715_));
  OAI21X1  g19279(.A0(new_n14501_), .A1(pi0698), .B0(new_n21715_), .Y(new_n21716_));
  OAI21X1  g19280(.A0(new_n2720_), .A1(pi0197), .B0(pi0832), .Y(new_n21717_));
  AOI21X1  g19281(.A0(new_n21716_), .A1(new_n2720_), .B0(new_n21717_), .Y(new_n21718_));
  AOI21X1  g19282(.A0(new_n21715_), .A1(new_n12077_), .B0(new_n2979_), .Y(new_n21719_));
  OAI21X1  g19283(.A0(new_n12446_), .A1(new_n7307_), .B0(new_n21719_), .Y(new_n21720_));
  AOI21X1  g19284(.A0(new_n14617_), .A1(pi0197), .B0(new_n2933_), .Y(new_n21721_));
  OAI21X1  g19285(.A0(new_n14515_), .A1(pi0197), .B0(new_n21721_), .Y(new_n21722_));
  OAI21X1  g19286(.A0(new_n14508_), .A1(pi0197), .B0(new_n14526_), .Y(new_n21723_));
  AND2X1   g19287(.A(new_n21723_), .B(new_n14191_), .Y(new_n21724_));
  OR2X1    g19288(.A(new_n14191_), .B(pi0197), .Y(new_n21725_));
  OAI21X1  g19289(.A0(new_n21725_), .A1(new_n12444_), .B0(pi0039), .Y(new_n21726_));
  AOI21X1  g19290(.A0(new_n21724_), .A1(new_n21722_), .B0(new_n21726_), .Y(new_n21727_));
  AOI21X1  g19291(.A0(new_n21714_), .A1(new_n11821_), .B0(pi0039), .Y(new_n21728_));
  OAI21X1  g19292(.A0(new_n11821_), .A1(pi0197), .B0(new_n21728_), .Y(new_n21729_));
  NAND2X1  g19293(.A(new_n21729_), .B(new_n2979_), .Y(new_n21730_));
  OAI21X1  g19294(.A0(new_n21730_), .A1(new_n21727_), .B0(new_n21720_), .Y(new_n21731_));
  AND2X1   g19295(.A(new_n21731_), .B(pi0698), .Y(new_n21732_));
  OAI21X1  g19296(.A0(new_n14603_), .A1(new_n7307_), .B0(new_n14191_), .Y(new_n21733_));
  AOI21X1  g19297(.A0(new_n14555_), .A1(new_n7307_), .B0(new_n21733_), .Y(new_n21734_));
  OAI21X1  g19298(.A0(new_n14582_), .A1(new_n7307_), .B0(pi0299), .Y(new_n21735_));
  AOI21X1  g19299(.A0(new_n14572_), .A1(new_n7307_), .B0(new_n21735_), .Y(new_n21736_));
  NOR2X1   g19300(.A(new_n14508_), .B(pi0197), .Y(new_n21737_));
  OAI21X1  g19301(.A0(new_n21737_), .A1(new_n14737_), .B0(pi0767), .Y(new_n21738_));
  OAI21X1  g19302(.A0(new_n21738_), .A1(new_n21736_), .B0(pi0039), .Y(new_n21739_));
  OAI22X1  g19303(.A0(new_n21739_), .A1(new_n21734_), .B0(new_n21729_), .B1(new_n14586_), .Y(new_n21740_));
  NOR2X1   g19304(.A(new_n12077_), .B(pi0197), .Y(new_n21741_));
  OAI21X1  g19305(.A0(new_n5362_), .A1(new_n14191_), .B0(new_n2939_), .Y(new_n21742_));
  OAI21X1  g19306(.A0(new_n21742_), .A1(new_n14669_), .B0(pi0038), .Y(new_n21743_));
  OAI21X1  g19307(.A0(new_n21743_), .A1(new_n21741_), .B0(new_n14359_), .Y(new_n21744_));
  AOI21X1  g19308(.A0(new_n21740_), .A1(new_n2979_), .B0(new_n21744_), .Y(new_n21745_));
  OAI21X1  g19309(.A0(new_n21745_), .A1(new_n21732_), .B0(new_n7625_), .Y(new_n21746_));
  AOI21X1  g19310(.A0(new_n9483_), .A1(new_n7307_), .B0(pi0832), .Y(new_n21747_));
  AOI21X1  g19311(.A0(new_n21747_), .A1(new_n21746_), .B0(new_n21718_), .Y(po0354));
  INVX1    g19312(.A(new_n13266_), .Y(new_n21749_));
  AOI21X1  g19313(.A0(new_n11822_), .A1(new_n3047_), .B0(new_n21749_), .Y(new_n21750_));
  OR3X1    g19314(.A(new_n11976_), .B(new_n5058_), .C(new_n2954_), .Y(new_n21751_));
  AND2X1   g19315(.A(new_n11825_), .B(pi0198), .Y(new_n21752_));
  NOR2X1   g19316(.A(new_n11900_), .B(new_n2954_), .Y(new_n21753_));
  MX2X1    g19317(.A(new_n21753_), .B(new_n21752_), .S0(new_n5021_), .Y(new_n21754_));
  AOI21X1  g19318(.A0(new_n21754_), .A1(new_n5058_), .B0(new_n10044_), .Y(new_n21755_));
  INVX1    g19319(.A(new_n21752_), .Y(new_n21756_));
  AOI21X1  g19320(.A0(new_n21756_), .A1(new_n10044_), .B0(pi0215), .Y(new_n21757_));
  INVX1    g19321(.A(new_n21757_), .Y(new_n21758_));
  AOI21X1  g19322(.A0(new_n21755_), .A1(new_n21751_), .B0(new_n21758_), .Y(new_n21759_));
  AOI21X1  g19323(.A0(new_n11843_), .A1(new_n11842_), .B0(new_n2954_), .Y(new_n21760_));
  INVX1    g19324(.A(new_n21760_), .Y(new_n21761_));
  AOI21X1  g19325(.A0(new_n21756_), .A1(new_n5021_), .B0(new_n21761_), .Y(new_n21762_));
  AOI21X1  g19326(.A0(new_n12195_), .A1(new_n5018_), .B0(new_n2954_), .Y(new_n21763_));
  OAI21X1  g19327(.A0(new_n11836_), .A1(new_n5018_), .B0(new_n21763_), .Y(new_n21764_));
  INVX1    g19328(.A(new_n21764_), .Y(new_n21765_));
  AOI21X1  g19329(.A0(new_n21765_), .A1(new_n5059_), .B0(new_n21762_), .Y(new_n21766_));
  OAI21X1  g19330(.A0(new_n21766_), .A1(new_n2934_), .B0(pi0299), .Y(new_n21767_));
  NOR2X1   g19331(.A(new_n21767_), .B(new_n21759_), .Y(new_n21768_));
  NOR3X1   g19332(.A(new_n11976_), .B(new_n5041_), .C(new_n2954_), .Y(new_n21769_));
  AND2X1   g19333(.A(new_n21754_), .B(new_n5041_), .Y(new_n21770_));
  OR3X1    g19334(.A(new_n21770_), .B(new_n21769_), .C(new_n2951_), .Y(new_n21771_));
  AOI21X1  g19335(.A0(new_n21756_), .A1(new_n2951_), .B0(pi0223), .Y(new_n21772_));
  AOI21X1  g19336(.A0(new_n21765_), .A1(new_n5042_), .B0(new_n21762_), .Y(new_n21773_));
  OAI21X1  g19337(.A0(new_n21773_), .A1(new_n2940_), .B0(new_n2933_), .Y(new_n21774_));
  AOI21X1  g19338(.A0(new_n21772_), .A1(new_n21771_), .B0(new_n21774_), .Y(new_n21775_));
  OR3X1    g19339(.A(new_n21775_), .B(new_n11576_), .C(new_n11770_), .Y(new_n21776_));
  OAI22X1  g19340(.A0(new_n21776_), .A1(new_n21768_), .B0(new_n21750_), .B1(new_n2954_), .Y(new_n21777_));
  INVX1    g19341(.A(new_n21777_), .Y(new_n21778_));
  AND2X1   g19342(.A(new_n11961_), .B(pi0198), .Y(new_n21779_));
  NAND2X1  g19343(.A(pi0633), .B(pi0603), .Y(new_n21780_));
  NOR2X1   g19344(.A(new_n12043_), .B(new_n12042_), .Y(new_n21781_));
  MX2X1    g19345(.A(new_n21781_), .B(new_n11965_), .S0(pi0198), .Y(new_n21782_));
  MX2X1    g19346(.A(new_n21782_), .B(new_n21779_), .S0(new_n21780_), .Y(new_n21783_));
  INVX1    g19347(.A(pi0633), .Y(new_n21784_));
  AOI21X1  g19348(.A0(new_n11964_), .A1(pi0198), .B0(new_n11970_), .Y(new_n21785_));
  OAI22X1  g19349(.A0(new_n21785_), .A1(new_n21784_), .B0(new_n11818_), .B1(new_n2954_), .Y(new_n21786_));
  NAND2X1  g19350(.A(new_n21786_), .B(new_n11973_), .Y(new_n21787_));
  OAI21X1  g19351(.A0(new_n21787_), .A1(pi0299), .B0(new_n2939_), .Y(new_n21788_));
  AOI21X1  g19352(.A0(new_n21783_), .A1(pi0299), .B0(new_n21788_), .Y(new_n21789_));
  NOR4X1   g19353(.A(new_n11979_), .B(new_n11824_), .C(new_n2725_), .D(new_n21784_), .Y(new_n21790_));
  AOI22X1  g19354(.A0(new_n21790_), .A1(pi0603), .B0(new_n11825_), .B1(pi0198), .Y(new_n21791_));
  AOI21X1  g19355(.A0(new_n11825_), .A1(pi0198), .B0(new_n21790_), .Y(new_n21792_));
  NOR2X1   g19356(.A(new_n21792_), .B(new_n5048_), .Y(new_n21793_));
  INVX1    g19357(.A(new_n21793_), .Y(new_n21794_));
  AOI21X1  g19358(.A0(new_n21790_), .A1(new_n12195_), .B0(new_n21760_), .Y(new_n21795_));
  AOI21X1  g19359(.A0(new_n21795_), .A1(new_n21794_), .B0(new_n11881_), .Y(new_n21796_));
  INVX1    g19360(.A(new_n21796_), .Y(new_n21797_));
  AOI21X1  g19361(.A0(new_n21752_), .A1(new_n11881_), .B0(new_n12001_), .Y(new_n21798_));
  AOI22X1  g19362(.A0(new_n21798_), .A1(new_n21797_), .B0(new_n21791_), .B1(new_n12001_), .Y(new_n21799_));
  AOI21X1  g19363(.A0(new_n21797_), .A1(new_n21761_), .B0(new_n5262_), .Y(new_n21800_));
  AOI21X1  g19364(.A0(new_n21799_), .A1(new_n5262_), .B0(new_n21800_), .Y(new_n21801_));
  INVX1    g19365(.A(new_n12023_), .Y(new_n21802_));
  OR4X1    g19366(.A(new_n12061_), .B(new_n12050_), .C(new_n11836_), .D(new_n21784_), .Y(new_n21803_));
  AND2X1   g19367(.A(new_n21803_), .B(new_n21764_), .Y(new_n21804_));
  NOR3X1   g19368(.A(new_n11834_), .B(new_n11831_), .C(new_n2954_), .Y(new_n21805_));
  AOI21X1  g19369(.A0(new_n21790_), .A1(new_n12195_), .B0(new_n21805_), .Y(new_n21806_));
  OAI22X1  g19370(.A0(new_n21806_), .A1(new_n21802_), .B0(new_n21804_), .B1(new_n5020_), .Y(new_n21807_));
  OAI21X1  g19371(.A0(new_n21807_), .A1(new_n5041_), .B0(pi0223), .Y(new_n21808_));
  AOI21X1  g19372(.A0(new_n21801_), .A1(new_n5041_), .B0(new_n21808_), .Y(new_n21809_));
  INVX1    g19373(.A(new_n11987_), .Y(new_n21810_));
  NOR2X1   g19374(.A(new_n11899_), .B(new_n2954_), .Y(new_n21811_));
  AOI21X1  g19375(.A0(new_n21810_), .A1(pi0633), .B0(new_n21811_), .Y(new_n21812_));
  MX2X1    g19376(.A(new_n21812_), .B(new_n21792_), .S0(new_n5023_), .Y(new_n21813_));
  NOR2X1   g19377(.A(new_n21813_), .B(new_n11881_), .Y(new_n21814_));
  OAI21X1  g19378(.A0(new_n21813_), .A1(new_n11881_), .B0(new_n5016_), .Y(new_n21815_));
  INVX1    g19379(.A(new_n5017_), .Y(new_n21816_));
  NOR2X1   g19380(.A(new_n21792_), .B(new_n11881_), .Y(new_n21817_));
  INVX1    g19381(.A(new_n21817_), .Y(new_n21818_));
  AOI21X1  g19382(.A0(new_n21818_), .A1(pi0642), .B0(new_n21816_), .Y(new_n21819_));
  OAI22X1  g19383(.A0(new_n21818_), .A1(new_n5017_), .B0(new_n21756_), .B1(pi0603), .Y(new_n21820_));
  AOI21X1  g19384(.A0(new_n21819_), .A1(new_n21815_), .B0(new_n21820_), .Y(new_n21821_));
  INVX1    g19385(.A(new_n21821_), .Y(new_n21822_));
  NOR3X1   g19386(.A(new_n11900_), .B(pi0603), .C(new_n2954_), .Y(new_n21823_));
  OR2X1    g19387(.A(new_n21823_), .B(new_n5262_), .Y(new_n21824_));
  OAI22X1  g19388(.A0(new_n21824_), .A1(new_n21814_), .B0(new_n21822_), .B1(new_n5020_), .Y(new_n21825_));
  OR3X1    g19389(.A(new_n21812_), .B(new_n12001_), .C(new_n11881_), .Y(new_n21826_));
  INVX1    g19390(.A(new_n21812_), .Y(new_n21827_));
  AND2X1   g19391(.A(new_n21792_), .B(new_n5048_), .Y(new_n21828_));
  NOR3X1   g19392(.A(new_n21828_), .B(new_n11999_), .C(new_n11881_), .Y(new_n21829_));
  OAI21X1  g19393(.A0(new_n21827_), .A1(new_n5048_), .B0(new_n21829_), .Y(new_n21830_));
  OR3X1    g19394(.A(new_n11925_), .B(pi0603), .C(new_n2954_), .Y(new_n21831_));
  AND3X1   g19395(.A(new_n21831_), .B(new_n21830_), .C(new_n21826_), .Y(new_n21832_));
  NOR2X1   g19396(.A(new_n21812_), .B(new_n11881_), .Y(new_n21833_));
  NOR3X1   g19397(.A(new_n21833_), .B(new_n21811_), .C(new_n5262_), .Y(new_n21834_));
  AOI21X1  g19398(.A0(new_n21832_), .A1(new_n5262_), .B0(new_n21834_), .Y(new_n21835_));
  AOI21X1  g19399(.A0(new_n21835_), .A1(new_n5042_), .B0(new_n2951_), .Y(new_n21836_));
  OAI21X1  g19400(.A0(new_n21825_), .A1(new_n5042_), .B0(new_n21836_), .Y(new_n21837_));
  AOI21X1  g19401(.A0(new_n21791_), .A1(new_n2951_), .B0(pi0223), .Y(new_n21838_));
  AOI21X1  g19402(.A0(new_n21838_), .A1(new_n21837_), .B0(new_n21809_), .Y(new_n21839_));
  NOR2X1   g19403(.A(new_n21839_), .B(pi0299), .Y(new_n21840_));
  OAI21X1  g19404(.A0(new_n21807_), .A1(new_n5058_), .B0(pi0215), .Y(new_n21841_));
  AOI21X1  g19405(.A0(new_n21801_), .A1(new_n5058_), .B0(new_n21841_), .Y(new_n21842_));
  AOI21X1  g19406(.A0(new_n21835_), .A1(new_n5059_), .B0(new_n10044_), .Y(new_n21843_));
  OAI21X1  g19407(.A0(new_n21825_), .A1(new_n5059_), .B0(new_n21843_), .Y(new_n21844_));
  AOI21X1  g19408(.A0(new_n21791_), .A1(new_n10044_), .B0(pi0215), .Y(new_n21845_));
  AOI21X1  g19409(.A0(new_n21845_), .A1(new_n21844_), .B0(new_n21842_), .Y(new_n21846_));
  OAI21X1  g19410(.A0(new_n21846_), .A1(new_n2933_), .B0(pi0039), .Y(new_n21847_));
  NOR2X1   g19411(.A(new_n21847_), .B(new_n21840_), .Y(new_n21848_));
  OAI21X1  g19412(.A0(new_n21848_), .A1(new_n21789_), .B0(new_n2979_), .Y(new_n21849_));
  AOI21X1  g19413(.A0(pi0198), .A1(pi0039), .B0(new_n2979_), .Y(new_n21850_));
  NOR3X1   g19414(.A(new_n11979_), .B(new_n21784_), .C(new_n11881_), .Y(new_n21851_));
  MX2X1    g19415(.A(pi0198), .B(new_n21851_), .S0(new_n11828_), .Y(new_n21852_));
  NAND2X1  g19416(.A(new_n21852_), .B(new_n2939_), .Y(new_n21853_));
  AOI21X1  g19417(.A0(new_n21853_), .A1(new_n21850_), .B0(new_n11770_), .Y(new_n21854_));
  AOI22X1  g19418(.A0(new_n21854_), .A1(new_n21849_), .B0(new_n11770_), .B1(pi0198), .Y(new_n21855_));
  MX2X1    g19419(.A(new_n21855_), .B(new_n21778_), .S0(new_n12473_), .Y(new_n21856_));
  OR2X1    g19420(.A(new_n21856_), .B(pi0785), .Y(new_n21857_));
  NOR2X1   g19421(.A(new_n21855_), .B(new_n12473_), .Y(new_n21858_));
  AOI22X1  g19422(.A0(new_n21858_), .A1(pi0609), .B0(new_n21777_), .B1(new_n12472_), .Y(new_n21859_));
  AOI22X1  g19423(.A0(new_n21858_), .A1(new_n12462_), .B0(new_n21777_), .B1(new_n12481_), .Y(new_n21860_));
  MX2X1    g19424(.A(new_n21860_), .B(new_n21859_), .S0(pi1155), .Y(new_n21861_));
  OAI21X1  g19425(.A0(new_n21861_), .A1(new_n11768_), .B0(new_n21857_), .Y(new_n21862_));
  NOR2X1   g19426(.A(new_n21862_), .B(new_n12486_), .Y(new_n21863_));
  OAI21X1  g19427(.A0(new_n21777_), .A1(pi0618), .B0(pi1154), .Y(new_n21864_));
  NOR2X1   g19428(.A(new_n21862_), .B(pi0618), .Y(new_n21865_));
  OAI21X1  g19429(.A0(new_n21777_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n21866_));
  OAI22X1  g19430(.A0(new_n21866_), .A1(new_n21865_), .B0(new_n21864_), .B1(new_n21863_), .Y(new_n21867_));
  MX2X1    g19431(.A(new_n21867_), .B(new_n21862_), .S0(new_n11767_), .Y(new_n21868_));
  AOI21X1  g19432(.A0(new_n21778_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n21869_));
  OAI21X1  g19433(.A0(new_n21868_), .A1(new_n12509_), .B0(new_n21869_), .Y(new_n21870_));
  AOI21X1  g19434(.A0(new_n21778_), .A1(pi0619), .B0(pi1159), .Y(new_n21871_));
  OAI21X1  g19435(.A0(new_n21868_), .A1(pi0619), .B0(new_n21871_), .Y(new_n21872_));
  AOI21X1  g19436(.A0(new_n21872_), .A1(new_n21870_), .B0(new_n11766_), .Y(new_n21873_));
  AOI21X1  g19437(.A0(new_n21868_), .A1(new_n11766_), .B0(new_n21873_), .Y(new_n21874_));
  MX2X1    g19438(.A(new_n21874_), .B(new_n21778_), .S0(new_n12708_), .Y(new_n21875_));
  MX2X1    g19439(.A(new_n21875_), .B(new_n21778_), .S0(new_n12580_), .Y(new_n21876_));
  NOR2X1   g19440(.A(new_n12563_), .B(new_n12531_), .Y(new_n21877_));
  INVX1    g19441(.A(new_n21877_), .Y(new_n21878_));
  AND2X1   g19442(.A(new_n21777_), .B(new_n12513_), .Y(new_n21879_));
  AOI22X1  g19443(.A0(new_n12157_), .A1(pi0634), .B0(new_n11825_), .B1(pi0198), .Y(new_n21880_));
  AOI21X1  g19444(.A0(new_n21880_), .A1(new_n5348_), .B0(new_n12108_), .Y(new_n21881_));
  AND3X1   g19445(.A(new_n12158_), .B(new_n11899_), .C(pi0634), .Y(new_n21882_));
  NOR2X1   g19446(.A(new_n21882_), .B(new_n21811_), .Y(new_n21883_));
  MX2X1    g19447(.A(new_n21883_), .B(new_n21880_), .S0(new_n5023_), .Y(new_n21884_));
  INVX1    g19448(.A(new_n21884_), .Y(new_n21885_));
  OAI21X1  g19449(.A0(new_n21885_), .A1(new_n5348_), .B0(new_n21881_), .Y(new_n21886_));
  OAI21X1  g19450(.A0(new_n11900_), .A1(new_n2954_), .B0(new_n5018_), .Y(new_n21887_));
  AOI21X1  g19451(.A0(new_n21756_), .A1(new_n5348_), .B0(pi0680), .Y(new_n21888_));
  AOI22X1  g19452(.A0(new_n21888_), .A1(new_n21887_), .B0(new_n21885_), .B1(new_n5020_), .Y(new_n21889_));
  AOI21X1  g19453(.A0(new_n21889_), .A1(new_n21886_), .B0(new_n5042_), .Y(new_n21890_));
  MX2X1    g19454(.A(new_n21883_), .B(new_n21880_), .S0(new_n5048_), .Y(new_n21891_));
  NOR3X1   g19455(.A(new_n21882_), .B(new_n21811_), .C(new_n5348_), .Y(new_n21892_));
  OR2X1    g19456(.A(new_n21892_), .B(new_n12108_), .Y(new_n21893_));
  AOI21X1  g19457(.A0(new_n21891_), .A1(new_n5348_), .B0(new_n21893_), .Y(new_n21894_));
  OR3X1    g19458(.A(new_n11926_), .B(pi0680), .C(new_n2954_), .Y(new_n21895_));
  OAI21X1  g19459(.A0(new_n21883_), .A1(new_n5262_), .B0(new_n21895_), .Y(new_n21896_));
  NOR2X1   g19460(.A(new_n21896_), .B(new_n21894_), .Y(new_n21897_));
  OAI21X1  g19461(.A0(new_n21897_), .A1(new_n5041_), .B0(new_n2952_), .Y(new_n21898_));
  NOR2X1   g19462(.A(new_n21898_), .B(new_n21890_), .Y(new_n21899_));
  OAI21X1  g19463(.A0(new_n21752_), .A1(new_n12157_), .B0(pi0634), .Y(new_n21900_));
  OAI21X1  g19464(.A0(new_n21900_), .A1(new_n5019_), .B0(new_n21756_), .Y(new_n21901_));
  OAI21X1  g19465(.A0(new_n21901_), .A1(new_n2952_), .B0(new_n2940_), .Y(new_n21902_));
  INVX1    g19466(.A(new_n21880_), .Y(new_n21903_));
  INVX1    g19467(.A(pi0634), .Y(new_n21904_));
  NOR3X1   g19468(.A(new_n12177_), .B(new_n11835_), .C(new_n21904_), .Y(new_n21905_));
  NOR2X1   g19469(.A(new_n21905_), .B(new_n21805_), .Y(new_n21906_));
  INVX1    g19470(.A(new_n21906_), .Y(new_n21907_));
  MX2X1    g19471(.A(new_n21907_), .B(new_n21903_), .S0(new_n5048_), .Y(new_n21908_));
  AOI21X1  g19472(.A0(new_n21906_), .A1(new_n5018_), .B0(new_n12108_), .Y(new_n21909_));
  OAI21X1  g19473(.A0(new_n21908_), .A1(new_n5018_), .B0(new_n21909_), .Y(new_n21910_));
  AOI22X1  g19474(.A0(new_n21907_), .A1(new_n5020_), .B0(new_n21765_), .B1(new_n5019_), .Y(new_n21911_));
  NAND3X1  g19475(.A(new_n21911_), .B(new_n21910_), .C(new_n5042_), .Y(new_n21912_));
  MX2X1    g19476(.A(new_n21906_), .B(new_n21880_), .S0(new_n5023_), .Y(new_n21913_));
  NAND2X1  g19477(.A(new_n21913_), .B(new_n5018_), .Y(new_n21914_));
  OR3X1    g19478(.A(new_n21764_), .B(new_n21761_), .C(pi0680), .Y(new_n21915_));
  OAI21X1  g19479(.A0(new_n21913_), .A1(new_n5262_), .B0(new_n21915_), .Y(new_n21916_));
  AOI21X1  g19480(.A0(new_n21914_), .A1(new_n21881_), .B0(new_n21916_), .Y(new_n21917_));
  AOI21X1  g19481(.A0(new_n21917_), .A1(new_n5041_), .B0(new_n2940_), .Y(new_n21918_));
  AOI21X1  g19482(.A0(new_n21918_), .A1(new_n21912_), .B0(pi0299), .Y(new_n21919_));
  OAI21X1  g19483(.A0(new_n21902_), .A1(new_n21899_), .B0(new_n21919_), .Y(new_n21920_));
  NOR2X1   g19484(.A(new_n21897_), .B(new_n5058_), .Y(new_n21921_));
  AOI21X1  g19485(.A0(new_n21889_), .A1(new_n21886_), .B0(new_n5059_), .Y(new_n21922_));
  NOR3X1   g19486(.A(new_n21922_), .B(new_n21921_), .C(new_n10044_), .Y(new_n21923_));
  OAI21X1  g19487(.A0(new_n21901_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n21924_));
  NAND3X1  g19488(.A(new_n21911_), .B(new_n21910_), .C(new_n5059_), .Y(new_n21925_));
  AOI21X1  g19489(.A0(new_n21917_), .A1(new_n5058_), .B0(new_n2934_), .Y(new_n21926_));
  AOI21X1  g19490(.A0(new_n21926_), .A1(new_n21925_), .B0(new_n2933_), .Y(new_n21927_));
  OAI21X1  g19491(.A0(new_n21924_), .A1(new_n21923_), .B0(new_n21927_), .Y(new_n21928_));
  AOI21X1  g19492(.A0(new_n21928_), .A1(new_n21920_), .B0(new_n2939_), .Y(new_n21929_));
  NAND2X1  g19493(.A(pi0680), .B(pi0634), .Y(new_n21930_));
  AND3X1   g19494(.A(new_n12327_), .B(new_n12326_), .C(new_n2954_), .Y(new_n21931_));
  AND2X1   g19495(.A(new_n12312_), .B(pi0198), .Y(new_n21932_));
  OR2X1    g19496(.A(new_n21932_), .B(new_n21931_), .Y(new_n21933_));
  MX2X1    g19497(.A(new_n21933_), .B(new_n21779_), .S0(new_n21930_), .Y(new_n21934_));
  NOR2X1   g19498(.A(new_n11818_), .B(new_n2954_), .Y(new_n21935_));
  OR4X1    g19499(.A(new_n11817_), .B(new_n11805_), .C(new_n12091_), .D(new_n2954_), .Y(new_n21936_));
  AOI21X1  g19500(.A0(new_n12317_), .A1(new_n2954_), .B0(new_n21930_), .Y(new_n21937_));
  AOI21X1  g19501(.A0(new_n21937_), .A1(new_n21936_), .B0(new_n21935_), .Y(new_n21938_));
  OAI21X1  g19502(.A0(new_n21938_), .A1(pi0299), .B0(new_n2939_), .Y(new_n21939_));
  AOI21X1  g19503(.A0(new_n21934_), .A1(pi0299), .B0(new_n21939_), .Y(new_n21940_));
  OAI21X1  g19504(.A0(new_n21940_), .A1(new_n21929_), .B0(new_n2979_), .Y(new_n21941_));
  OR3X1    g19505(.A(new_n12084_), .B(new_n5019_), .C(new_n21904_), .Y(new_n21942_));
  MX2X1    g19506(.A(new_n2954_), .B(new_n21942_), .S0(new_n11828_), .Y(new_n21943_));
  OAI21X1  g19507(.A0(new_n21943_), .A1(pi0039), .B0(new_n21850_), .Y(new_n21944_));
  AND2X1   g19508(.A(new_n21944_), .B(new_n3103_), .Y(new_n21945_));
  AOI22X1  g19509(.A0(new_n21945_), .A1(new_n21941_), .B0(new_n11770_), .B1(pi0198), .Y(new_n21946_));
  OAI21X1  g19510(.A0(new_n21777_), .A1(pi0625), .B0(pi1153), .Y(new_n21947_));
  AOI21X1  g19511(.A0(new_n21946_), .A1(pi0625), .B0(new_n21947_), .Y(new_n21948_));
  OAI21X1  g19512(.A0(new_n21777_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n21949_));
  AOI21X1  g19513(.A0(new_n21946_), .A1(new_n12363_), .B0(new_n21949_), .Y(new_n21950_));
  NOR2X1   g19514(.A(new_n21950_), .B(new_n21948_), .Y(new_n21951_));
  MX2X1    g19515(.A(new_n21951_), .B(new_n21946_), .S0(new_n11769_), .Y(new_n21952_));
  INVX1    g19516(.A(new_n21952_), .Y(new_n21953_));
  MX2X1    g19517(.A(new_n21953_), .B(new_n21777_), .S0(new_n12490_), .Y(new_n21954_));
  AOI21X1  g19518(.A0(new_n21954_), .A1(new_n14053_), .B0(new_n21879_), .Y(new_n21955_));
  AND3X1   g19519(.A(new_n21955_), .B(new_n13356_), .C(new_n14051_), .Y(new_n21956_));
  AOI21X1  g19520(.A0(new_n21778_), .A1(new_n21878_), .B0(new_n21956_), .Y(new_n21957_));
  MX2X1    g19521(.A(new_n21957_), .B(new_n21777_), .S0(new_n12554_), .Y(new_n21958_));
  INVX1    g19522(.A(new_n21958_), .Y(new_n21959_));
  AOI21X1  g19523(.A0(new_n21778_), .A1(pi0628), .B0(pi1156), .Y(new_n21960_));
  OAI21X1  g19524(.A0(new_n21957_), .A1(pi0628), .B0(new_n21960_), .Y(new_n21961_));
  OAI21X1  g19525(.A0(new_n21959_), .A1(new_n12555_), .B0(new_n21961_), .Y(new_n21962_));
  MX2X1    g19526(.A(new_n21962_), .B(new_n21957_), .S0(new_n11764_), .Y(new_n21963_));
  AOI21X1  g19527(.A0(new_n21778_), .A1(pi0647), .B0(pi1157), .Y(new_n21964_));
  OAI21X1  g19528(.A0(new_n21963_), .A1(pi0647), .B0(new_n21964_), .Y(new_n21965_));
  INVX1    g19529(.A(new_n21965_), .Y(new_n21966_));
  INVX1    g19530(.A(new_n21963_), .Y(new_n21967_));
  MX2X1    g19531(.A(new_n21967_), .B(new_n21778_), .S0(new_n12577_), .Y(new_n21968_));
  INVX1    g19532(.A(new_n21968_), .Y(new_n21969_));
  AOI22X1  g19533(.A0(new_n21969_), .A1(new_n14241_), .B0(new_n21966_), .B1(pi0630), .Y(new_n21970_));
  OAI21X1  g19534(.A0(new_n21876_), .A1(new_n14239_), .B0(new_n21970_), .Y(new_n21971_));
  NOR2X1   g19535(.A(new_n21875_), .B(new_n14250_), .Y(new_n21972_));
  INVX1    g19536(.A(new_n16373_), .Y(new_n21973_));
  OAI22X1  g19537(.A0(new_n21961_), .A1(new_n12561_), .B0(new_n21959_), .B1(new_n21973_), .Y(new_n21974_));
  NOR2X1   g19538(.A(new_n21974_), .B(new_n21972_), .Y(new_n21975_));
  AOI21X1  g19539(.A0(new_n21777_), .A1(pi0626), .B0(new_n16218_), .Y(new_n21976_));
  OAI21X1  g19540(.A0(new_n21874_), .A1(pi0626), .B0(new_n21976_), .Y(new_n21977_));
  AOI21X1  g19541(.A0(new_n21777_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n21978_));
  OAI21X1  g19542(.A0(new_n21874_), .A1(new_n12542_), .B0(new_n21978_), .Y(new_n21979_));
  MX2X1    g19543(.A(new_n21955_), .B(new_n21778_), .S0(new_n12531_), .Y(new_n21980_));
  NAND2X1  g19544(.A(new_n21980_), .B(new_n12637_), .Y(new_n21981_));
  AND3X1   g19545(.A(new_n21981_), .B(new_n21979_), .C(new_n21977_), .Y(new_n21982_));
  OAI21X1  g19546(.A0(pi0665), .A1(new_n2954_), .B0(pi0633), .Y(new_n21983_));
  NOR3X1   g19547(.A(new_n21983_), .B(new_n21931_), .C(new_n21782_), .Y(new_n21984_));
  NOR3X1   g19548(.A(new_n12338_), .B(new_n21781_), .C(new_n2954_), .Y(new_n21985_));
  OR2X1    g19549(.A(pi0665), .B(pi0198), .Y(new_n21986_));
  OAI21X1  g19550(.A0(new_n21986_), .A1(new_n11965_), .B0(new_n21784_), .Y(new_n21987_));
  OAI21X1  g19551(.A0(new_n21987_), .A1(new_n21985_), .B0(pi0603), .Y(new_n21988_));
  NOR2X1   g19552(.A(new_n21988_), .B(new_n21984_), .Y(new_n21989_));
  AOI21X1  g19553(.A0(new_n21933_), .A1(new_n11881_), .B0(new_n21989_), .Y(new_n21990_));
  AOI21X1  g19554(.A0(new_n21930_), .A1(new_n21783_), .B0(new_n2933_), .Y(new_n21991_));
  OAI21X1  g19555(.A0(new_n21990_), .A1(new_n21930_), .B0(new_n21991_), .Y(new_n21992_));
  AND2X1   g19556(.A(new_n11971_), .B(new_n11818_), .Y(new_n21993_));
  OR3X1    g19557(.A(new_n11818_), .B(pi0634), .C(new_n2954_), .Y(new_n21994_));
  NAND3X1  g19558(.A(new_n12307_), .B(pi0634), .C(pi0198), .Y(new_n21995_));
  OAI21X1  g19559(.A0(new_n21995_), .A1(new_n21993_), .B0(new_n21994_), .Y(new_n21996_));
  AOI21X1  g19560(.A0(new_n11806_), .A1(pi0621), .B0(pi0198), .Y(new_n21997_));
  INVX1    g19561(.A(new_n21997_), .Y(new_n21998_));
  OR2X1    g19562(.A(pi0665), .B(new_n21904_), .Y(new_n21999_));
  AOI21X1  g19563(.A0(new_n21784_), .A1(pi0198), .B0(new_n21999_), .Y(new_n22000_));
  AOI21X1  g19564(.A0(new_n22000_), .A1(new_n21998_), .B0(new_n11881_), .Y(new_n22001_));
  OAI21X1  g19565(.A0(new_n21785_), .A1(new_n21784_), .B0(new_n22001_), .Y(new_n22002_));
  AOI21X1  g19566(.A0(new_n21996_), .A1(new_n21784_), .B0(new_n22002_), .Y(new_n22003_));
  AND2X1   g19567(.A(new_n21938_), .B(new_n11881_), .Y(new_n22004_));
  NOR3X1   g19568(.A(new_n22004_), .B(new_n22003_), .C(new_n5019_), .Y(new_n22005_));
  OAI21X1  g19569(.A0(new_n21787_), .A1(pi0680), .B0(new_n2933_), .Y(new_n22006_));
  OR2X1    g19570(.A(new_n22006_), .B(new_n22005_), .Y(new_n22007_));
  AOI21X1  g19571(.A0(new_n22007_), .A1(new_n21992_), .B0(pi0039), .Y(new_n22008_));
  OAI21X1  g19572(.A0(new_n21999_), .A1(new_n11994_), .B0(new_n21792_), .Y(new_n22009_));
  OAI21X1  g19573(.A0(new_n12163_), .A1(new_n21904_), .B0(new_n21812_), .Y(new_n22010_));
  MX2X1    g19574(.A(new_n22010_), .B(new_n22009_), .S0(new_n5023_), .Y(new_n22011_));
  NAND2X1  g19575(.A(new_n22011_), .B(pi0603), .Y(new_n22012_));
  AND3X1   g19576(.A(new_n22011_), .B(new_n5016_), .C(pi0603), .Y(new_n22013_));
  AND2X1   g19577(.A(new_n22009_), .B(pi0603), .Y(new_n22014_));
  AOI22X1  g19578(.A0(new_n22014_), .A1(pi0642), .B0(new_n21903_), .B1(new_n11881_), .Y(new_n22015_));
  INVX1    g19579(.A(new_n22015_), .Y(new_n22016_));
  OAI21X1  g19580(.A0(new_n22016_), .A1(new_n22013_), .B0(new_n5017_), .Y(new_n22017_));
  AOI21X1  g19581(.A0(new_n21903_), .A1(new_n11881_), .B0(new_n22014_), .Y(new_n22018_));
  INVX1    g19582(.A(new_n22018_), .Y(new_n22019_));
  AOI21X1  g19583(.A0(new_n22019_), .A1(new_n21816_), .B0(new_n11863_), .Y(new_n22020_));
  AOI21X1  g19584(.A0(new_n21885_), .A1(new_n11881_), .B0(new_n11867_), .Y(new_n22021_));
  AOI22X1  g19585(.A0(new_n22021_), .A1(new_n22012_), .B0(new_n22020_), .B1(new_n22017_), .Y(new_n22022_));
  MX2X1    g19586(.A(new_n22022_), .B(new_n21822_), .S0(new_n5019_), .Y(new_n22023_));
  OR2X1    g19587(.A(new_n21832_), .B(pi0680), .Y(new_n22024_));
  NOR2X1   g19588(.A(new_n21891_), .B(pi0603), .Y(new_n22025_));
  AOI21X1  g19589(.A0(new_n12162_), .A1(pi0634), .B0(new_n21827_), .Y(new_n22026_));
  AND3X1   g19590(.A(new_n22009_), .B(new_n12001_), .C(pi0603), .Y(new_n22027_));
  NOR2X1   g19591(.A(new_n22027_), .B(new_n21829_), .Y(new_n22028_));
  OAI21X1  g19592(.A0(new_n22027_), .A1(new_n21829_), .B0(new_n5048_), .Y(new_n22029_));
  AOI22X1  g19593(.A0(new_n22029_), .A1(new_n22026_), .B0(new_n22028_), .B1(new_n5348_), .Y(new_n22030_));
  OAI21X1  g19594(.A0(new_n22030_), .A1(new_n22025_), .B0(new_n12083_), .Y(new_n22031_));
  OAI22X1  g19595(.A0(new_n21883_), .A1(new_n11991_), .B0(new_n21812_), .B1(new_n11881_), .Y(new_n22032_));
  NAND2X1  g19596(.A(new_n22032_), .B(new_n5020_), .Y(new_n22033_));
  AND3X1   g19597(.A(new_n22033_), .B(new_n22031_), .C(new_n22024_), .Y(new_n22034_));
  OAI21X1  g19598(.A0(new_n22034_), .A1(new_n5041_), .B0(new_n2952_), .Y(new_n22035_));
  AOI21X1  g19599(.A0(new_n22023_), .A1(new_n5041_), .B0(new_n22035_), .Y(new_n22036_));
  OAI21X1  g19600(.A0(new_n21900_), .A1(new_n12352_), .B0(new_n21791_), .Y(new_n22037_));
  OAI21X1  g19601(.A0(new_n22037_), .A1(new_n2952_), .B0(new_n2940_), .Y(new_n22038_));
  NOR2X1   g19602(.A(new_n22038_), .B(new_n22036_), .Y(new_n22039_));
  NOR2X1   g19603(.A(new_n21986_), .B(new_n12009_), .Y(new_n22040_));
  AND3X1   g19604(.A(new_n11979_), .B(new_n12091_), .C(pi0198), .Y(new_n22041_));
  NOR3X1   g19605(.A(new_n22041_), .B(new_n22040_), .C(new_n21805_), .Y(new_n22042_));
  AOI22X1  g19606(.A0(new_n21805_), .A1(new_n21904_), .B0(new_n21790_), .B1(new_n12195_), .Y(new_n22043_));
  OAI21X1  g19607(.A0(new_n22042_), .A1(new_n21904_), .B0(new_n22043_), .Y(new_n22044_));
  MX2X1    g19608(.A(new_n22044_), .B(new_n22009_), .S0(new_n5023_), .Y(new_n22045_));
  NOR2X1   g19609(.A(new_n21913_), .B(pi0603), .Y(new_n22046_));
  AOI21X1  g19610(.A0(new_n22045_), .A1(pi0603), .B0(new_n22046_), .Y(new_n22047_));
  NOR2X1   g19611(.A(new_n22047_), .B(new_n5262_), .Y(new_n22048_));
  OAI21X1  g19612(.A0(new_n21880_), .A1(pi0603), .B0(new_n11999_), .Y(new_n22049_));
  AOI21X1  g19613(.A0(new_n22045_), .A1(pi0603), .B0(new_n22049_), .Y(new_n22050_));
  OAI21X1  g19614(.A0(new_n22019_), .A1(new_n11999_), .B0(new_n12083_), .Y(new_n22051_));
  NAND2X1  g19615(.A(new_n21799_), .B(new_n5019_), .Y(new_n22052_));
  OAI21X1  g19616(.A0(new_n22051_), .A1(new_n22050_), .B0(new_n22052_), .Y(new_n22053_));
  OR3X1    g19617(.A(new_n22053_), .B(new_n22048_), .C(new_n5042_), .Y(new_n22054_));
  NOR2X1   g19618(.A(new_n22028_), .B(new_n5023_), .Y(new_n22055_));
  AND2X1   g19619(.A(new_n21908_), .B(new_n11881_), .Y(new_n22056_));
  AND3X1   g19620(.A(new_n22044_), .B(new_n11999_), .C(pi0603), .Y(new_n22057_));
  INVX1    g19621(.A(new_n22044_), .Y(new_n22058_));
  NOR2X1   g19622(.A(new_n22058_), .B(new_n22028_), .Y(new_n22059_));
  NOR4X1   g19623(.A(new_n22059_), .B(new_n22057_), .C(new_n22056_), .D(new_n22055_), .Y(new_n22060_));
  OR2X1    g19624(.A(new_n22060_), .B(new_n12108_), .Y(new_n22061_));
  MX2X1    g19625(.A(new_n22058_), .B(new_n21906_), .S0(new_n11881_), .Y(new_n22062_));
  OAI22X1  g19626(.A0(new_n22062_), .A1(new_n5262_), .B0(new_n21804_), .B1(pi0680), .Y(new_n22063_));
  INVX1    g19627(.A(new_n22063_), .Y(new_n22064_));
  NAND3X1  g19628(.A(new_n22064_), .B(new_n22061_), .C(new_n5042_), .Y(new_n22065_));
  AND3X1   g19629(.A(new_n22065_), .B(new_n22054_), .C(pi0223), .Y(new_n22066_));
  OAI21X1  g19630(.A0(new_n22066_), .A1(new_n22039_), .B0(new_n2933_), .Y(new_n22067_));
  OAI21X1  g19631(.A0(new_n22034_), .A1(new_n5058_), .B0(new_n10045_), .Y(new_n22068_));
  AOI21X1  g19632(.A0(new_n22023_), .A1(new_n5058_), .B0(new_n22068_), .Y(new_n22069_));
  OAI21X1  g19633(.A0(new_n22037_), .A1(new_n10045_), .B0(new_n2934_), .Y(new_n22070_));
  NOR3X1   g19634(.A(new_n22053_), .B(new_n22048_), .C(new_n5059_), .Y(new_n22071_));
  AND3X1   g19635(.A(new_n22064_), .B(new_n22061_), .C(new_n5059_), .Y(new_n22072_));
  OR3X1    g19636(.A(new_n22072_), .B(new_n22071_), .C(new_n2934_), .Y(new_n22073_));
  OAI21X1  g19637(.A0(new_n22070_), .A1(new_n22069_), .B0(new_n22073_), .Y(new_n22074_));
  AOI21X1  g19638(.A0(new_n22074_), .A1(pi0299), .B0(new_n2939_), .Y(new_n22075_));
  AOI21X1  g19639(.A0(new_n22075_), .A1(new_n22067_), .B0(new_n22008_), .Y(new_n22076_));
  AND2X1   g19640(.A(new_n12353_), .B(pi0634), .Y(new_n22077_));
  OAI21X1  g19641(.A0(new_n22077_), .A1(new_n21852_), .B0(new_n2939_), .Y(new_n22078_));
  AOI21X1  g19642(.A0(new_n22078_), .A1(new_n21850_), .B0(new_n11770_), .Y(new_n22079_));
  OAI21X1  g19643(.A0(new_n22076_), .A1(pi0038), .B0(new_n22079_), .Y(new_n22080_));
  OAI21X1  g19644(.A0(new_n3103_), .A1(new_n2954_), .B0(new_n22080_), .Y(new_n22081_));
  AOI21X1  g19645(.A0(new_n21855_), .A1(pi0625), .B0(pi1153), .Y(new_n22082_));
  OAI21X1  g19646(.A0(new_n22081_), .A1(pi0625), .B0(new_n22082_), .Y(new_n22083_));
  NOR2X1   g19647(.A(new_n21948_), .B(pi0608), .Y(new_n22084_));
  AOI21X1  g19648(.A0(new_n21855_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n22085_));
  OAI21X1  g19649(.A0(new_n22081_), .A1(new_n12363_), .B0(new_n22085_), .Y(new_n22086_));
  NOR2X1   g19650(.A(new_n21950_), .B(new_n12368_), .Y(new_n22087_));
  AOI22X1  g19651(.A0(new_n22087_), .A1(new_n22086_), .B0(new_n22084_), .B1(new_n22083_), .Y(new_n22088_));
  OR2X1    g19652(.A(new_n22081_), .B(pi0778), .Y(new_n22089_));
  OAI21X1  g19653(.A0(new_n22088_), .A1(new_n11769_), .B0(new_n22089_), .Y(new_n22090_));
  OAI21X1  g19654(.A0(new_n21953_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n22091_));
  AOI21X1  g19655(.A0(new_n22090_), .A1(new_n12462_), .B0(new_n22091_), .Y(new_n22092_));
  OAI21X1  g19656(.A0(new_n21859_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n22093_));
  OAI21X1  g19657(.A0(new_n21953_), .A1(pi0609), .B0(pi1155), .Y(new_n22094_));
  AOI21X1  g19658(.A0(new_n22090_), .A1(pi0609), .B0(new_n22094_), .Y(new_n22095_));
  OAI21X1  g19659(.A0(new_n21860_), .A1(pi1155), .B0(pi0660), .Y(new_n22096_));
  OAI22X1  g19660(.A0(new_n22096_), .A1(new_n22095_), .B0(new_n22093_), .B1(new_n22092_), .Y(new_n22097_));
  MX2X1    g19661(.A(new_n22097_), .B(new_n22090_), .S0(new_n11768_), .Y(new_n22098_));
  OAI21X1  g19662(.A0(new_n21954_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n22099_));
  AOI21X1  g19663(.A0(new_n22098_), .A1(new_n12486_), .B0(new_n22099_), .Y(new_n22100_));
  OAI21X1  g19664(.A0(new_n21864_), .A1(new_n21863_), .B0(new_n12494_), .Y(new_n22101_));
  OAI21X1  g19665(.A0(new_n21954_), .A1(pi0618), .B0(pi1154), .Y(new_n22102_));
  AOI21X1  g19666(.A0(new_n22098_), .A1(pi0618), .B0(new_n22102_), .Y(new_n22103_));
  OAI21X1  g19667(.A0(new_n21866_), .A1(new_n21865_), .B0(pi0627), .Y(new_n22104_));
  OAI22X1  g19668(.A0(new_n22104_), .A1(new_n22103_), .B0(new_n22101_), .B1(new_n22100_), .Y(new_n22105_));
  MX2X1    g19669(.A(new_n22105_), .B(new_n22098_), .S0(new_n11767_), .Y(new_n22106_));
  NAND2X1  g19670(.A(new_n22106_), .B(new_n12509_), .Y(new_n22107_));
  AOI21X1  g19671(.A0(new_n21955_), .A1(pi0619), .B0(pi1159), .Y(new_n22108_));
  NAND2X1  g19672(.A(new_n21870_), .B(new_n12517_), .Y(new_n22109_));
  AOI21X1  g19673(.A0(new_n22108_), .A1(new_n22107_), .B0(new_n22109_), .Y(new_n22110_));
  NAND2X1  g19674(.A(new_n22106_), .B(pi0619), .Y(new_n22111_));
  AOI21X1  g19675(.A0(new_n21955_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n22112_));
  NAND2X1  g19676(.A(new_n21872_), .B(pi0648), .Y(new_n22113_));
  AOI21X1  g19677(.A0(new_n22112_), .A1(new_n22111_), .B0(new_n22113_), .Y(new_n22114_));
  NOR3X1   g19678(.A(new_n22114_), .B(new_n22110_), .C(new_n11766_), .Y(new_n22115_));
  OAI21X1  g19679(.A0(new_n22106_), .A1(pi0789), .B0(new_n12709_), .Y(new_n22116_));
  OAI22X1  g19680(.A0(new_n22116_), .A1(new_n22115_), .B0(new_n21982_), .B1(new_n11765_), .Y(new_n22117_));
  OAI21X1  g19681(.A0(new_n21975_), .A1(new_n11764_), .B0(new_n22117_), .Y(new_n22118_));
  AOI21X1  g19682(.A0(new_n21975_), .A1(new_n14125_), .B0(new_n14121_), .Y(new_n22119_));
  AOI22X1  g19683(.A0(new_n22119_), .A1(new_n22118_), .B0(new_n21971_), .B1(pi0787), .Y(new_n22120_));
  NAND2X1  g19684(.A(new_n22120_), .B(pi0644), .Y(new_n22121_));
  AOI21X1  g19685(.A0(new_n21969_), .A1(pi1157), .B0(new_n21966_), .Y(new_n22122_));
  MX2X1    g19686(.A(new_n22122_), .B(new_n21967_), .S0(new_n11763_), .Y(new_n22123_));
  AOI21X1  g19687(.A0(new_n22123_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n22124_));
  MX2X1    g19688(.A(new_n21876_), .B(new_n21778_), .S0(new_n12604_), .Y(new_n22125_));
  OAI21X1  g19689(.A0(new_n21777_), .A1(pi0644), .B0(new_n12608_), .Y(new_n22126_));
  AOI21X1  g19690(.A0(new_n22125_), .A1(pi0644), .B0(new_n22126_), .Y(new_n22127_));
  OR2X1    g19691(.A(new_n22127_), .B(new_n11762_), .Y(new_n22128_));
  AOI21X1  g19692(.A0(new_n22124_), .A1(new_n22121_), .B0(new_n22128_), .Y(new_n22129_));
  NAND2X1  g19693(.A(new_n22120_), .B(new_n12612_), .Y(new_n22130_));
  AOI21X1  g19694(.A0(new_n22123_), .A1(pi0644), .B0(pi0715), .Y(new_n22131_));
  OAI21X1  g19695(.A0(new_n21777_), .A1(new_n12612_), .B0(pi0715), .Y(new_n22132_));
  AOI21X1  g19696(.A0(new_n22125_), .A1(new_n12612_), .B0(new_n22132_), .Y(new_n22133_));
  OR2X1    g19697(.A(new_n22133_), .B(pi1160), .Y(new_n22134_));
  AOI21X1  g19698(.A0(new_n22131_), .A1(new_n22130_), .B0(new_n22134_), .Y(new_n22135_));
  OR3X1    g19699(.A(new_n22135_), .B(new_n22129_), .C(new_n12766_), .Y(new_n22136_));
  OAI21X1  g19700(.A0(new_n22120_), .A1(pi0790), .B0(new_n22136_), .Y(new_n22137_));
  MX2X1    g19701(.A(new_n22137_), .B(pi0198), .S0(po1038), .Y(po0355));
  INVX1    g19702(.A(pi0637), .Y(new_n22139_));
  AOI21X1  g19703(.A0(new_n12447_), .A1(new_n3103_), .B0(new_n7871_), .Y(new_n22140_));
  INVX1    g19704(.A(new_n13567_), .Y(new_n22141_));
  NOR2X1   g19705(.A(new_n13564_), .B(pi0199), .Y(new_n22142_));
  NOR2X1   g19706(.A(new_n12776_), .B(new_n7871_), .Y(new_n22143_));
  OAI21X1  g19707(.A0(new_n12074_), .A1(pi0199), .B0(new_n2979_), .Y(new_n22144_));
  OAI22X1  g19708(.A0(new_n22144_), .A1(new_n22143_), .B0(new_n22142_), .B1(new_n22141_), .Y(new_n22145_));
  AND2X1   g19709(.A(new_n22145_), .B(new_n3103_), .Y(new_n22146_));
  OAI21X1  g19710(.A0(new_n3103_), .A1(new_n7871_), .B0(pi0617), .Y(new_n22147_));
  OAI22X1  g19711(.A0(new_n22147_), .A1(new_n22146_), .B0(new_n22140_), .B1(pi0617), .Y(new_n22148_));
  OR3X1    g19712(.A(new_n13542_), .B(new_n7871_), .C(pi0038), .Y(new_n22149_));
  NAND2X1  g19713(.A(new_n16664_), .B(new_n3103_), .Y(new_n22150_));
  INVX1    g19714(.A(pi0617), .Y(new_n22151_));
  OAI21X1  g19715(.A0(new_n13541_), .A1(new_n2979_), .B0(new_n22151_), .Y(new_n22152_));
  AOI21X1  g19716(.A0(new_n22150_), .A1(new_n7871_), .B0(new_n22152_), .Y(new_n22153_));
  OR2X1    g19717(.A(new_n3103_), .B(new_n7871_), .Y(new_n22154_));
  AOI21X1  g19718(.A0(new_n13554_), .A1(new_n3103_), .B0(pi0199), .Y(new_n22155_));
  OAI21X1  g19719(.A0(new_n16670_), .A1(new_n7871_), .B0(pi0617), .Y(new_n22156_));
  OAI21X1  g19720(.A0(new_n22156_), .A1(new_n22155_), .B0(new_n22154_), .Y(new_n22157_));
  AOI21X1  g19721(.A0(new_n22153_), .A1(new_n22149_), .B0(new_n22157_), .Y(new_n22158_));
  MX2X1    g19722(.A(new_n22158_), .B(new_n22148_), .S0(new_n22139_), .Y(new_n22159_));
  OAI21X1  g19723(.A0(new_n12832_), .A1(new_n11770_), .B0(pi0199), .Y(new_n22160_));
  AOI21X1  g19724(.A0(new_n22145_), .A1(new_n3103_), .B0(new_n22147_), .Y(new_n22161_));
  AOI21X1  g19725(.A0(new_n22160_), .A1(new_n22151_), .B0(new_n22161_), .Y(new_n22162_));
  OAI21X1  g19726(.A0(new_n22162_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n22163_));
  AOI21X1  g19727(.A0(new_n22159_), .A1(new_n12363_), .B0(new_n22163_), .Y(new_n22164_));
  AND2X1   g19728(.A(new_n22160_), .B(new_n22139_), .Y(new_n22165_));
  AOI21X1  g19729(.A0(new_n12771_), .A1(new_n7871_), .B0(new_n13874_), .Y(new_n22166_));
  OAI21X1  g19730(.A0(new_n12394_), .A1(pi0199), .B0(pi0039), .Y(new_n22167_));
  AOI21X1  g19731(.A0(new_n12824_), .A1(pi0199), .B0(new_n22167_), .Y(new_n22168_));
  OAI21X1  g19732(.A0(new_n12435_), .A1(pi0199), .B0(new_n2939_), .Y(new_n22169_));
  AOI21X1  g19733(.A0(new_n12340_), .A1(pi0199), .B0(new_n22169_), .Y(new_n22170_));
  NOR3X1   g19734(.A(new_n22170_), .B(new_n22168_), .C(pi0038), .Y(new_n22171_));
  OAI21X1  g19735(.A0(new_n22171_), .A1(new_n22166_), .B0(new_n3103_), .Y(new_n22172_));
  AND3X1   g19736(.A(new_n22172_), .B(new_n22154_), .C(pi0637), .Y(new_n22173_));
  OR2X1    g19737(.A(new_n22173_), .B(new_n22165_), .Y(new_n22174_));
  AND2X1   g19738(.A(new_n22174_), .B(pi0625), .Y(new_n22175_));
  OAI21X1  g19739(.A0(new_n22140_), .A1(pi0625), .B0(pi1153), .Y(new_n22176_));
  OAI21X1  g19740(.A0(new_n22176_), .A1(new_n22175_), .B0(new_n12368_), .Y(new_n22177_));
  OAI21X1  g19741(.A0(new_n22162_), .A1(pi0625), .B0(pi1153), .Y(new_n22178_));
  AOI21X1  g19742(.A0(new_n22159_), .A1(pi0625), .B0(new_n22178_), .Y(new_n22179_));
  AND2X1   g19743(.A(new_n22174_), .B(new_n12363_), .Y(new_n22180_));
  OAI21X1  g19744(.A0(new_n22140_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n22181_));
  OAI21X1  g19745(.A0(new_n22181_), .A1(new_n22180_), .B0(pi0608), .Y(new_n22182_));
  OAI22X1  g19746(.A0(new_n22182_), .A1(new_n22179_), .B0(new_n22177_), .B1(new_n22164_), .Y(new_n22183_));
  MX2X1    g19747(.A(new_n22183_), .B(new_n22159_), .S0(new_n11769_), .Y(new_n22184_));
  INVX1    g19748(.A(new_n22174_), .Y(new_n22185_));
  OAI22X1  g19749(.A0(new_n22181_), .A1(new_n22180_), .B0(new_n22176_), .B1(new_n22175_), .Y(new_n22186_));
  MX2X1    g19750(.A(new_n22186_), .B(new_n22185_), .S0(new_n11769_), .Y(new_n22187_));
  OAI21X1  g19751(.A0(new_n22187_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n22188_));
  AOI21X1  g19752(.A0(new_n22184_), .A1(new_n12462_), .B0(new_n22188_), .Y(new_n22189_));
  MX2X1    g19753(.A(new_n22148_), .B(new_n22160_), .S0(new_n12473_), .Y(new_n22190_));
  OAI21X1  g19754(.A0(new_n22140_), .A1(pi0609), .B0(pi1155), .Y(new_n22191_));
  AOI21X1  g19755(.A0(new_n22190_), .A1(pi0609), .B0(new_n22191_), .Y(new_n22192_));
  OR2X1    g19756(.A(new_n22192_), .B(pi0660), .Y(new_n22193_));
  OAI21X1  g19757(.A0(new_n22187_), .A1(pi0609), .B0(pi1155), .Y(new_n22194_));
  AOI21X1  g19758(.A0(new_n22184_), .A1(pi0609), .B0(new_n22194_), .Y(new_n22195_));
  OAI21X1  g19759(.A0(new_n22140_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n22196_));
  AOI21X1  g19760(.A0(new_n22190_), .A1(new_n12462_), .B0(new_n22196_), .Y(new_n22197_));
  OR2X1    g19761(.A(new_n22197_), .B(new_n12468_), .Y(new_n22198_));
  OAI22X1  g19762(.A0(new_n22198_), .A1(new_n22195_), .B0(new_n22193_), .B1(new_n22189_), .Y(new_n22199_));
  MX2X1    g19763(.A(new_n22199_), .B(new_n22184_), .S0(new_n11768_), .Y(new_n22200_));
  MX2X1    g19764(.A(new_n22187_), .B(new_n22140_), .S0(new_n12490_), .Y(new_n22201_));
  OAI21X1  g19765(.A0(new_n22201_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n22202_));
  AOI21X1  g19766(.A0(new_n22200_), .A1(new_n12486_), .B0(new_n22202_), .Y(new_n22203_));
  OAI21X1  g19767(.A0(new_n22197_), .A1(new_n22192_), .B0(pi0785), .Y(new_n22204_));
  OAI21X1  g19768(.A0(new_n22190_), .A1(pi0785), .B0(new_n22204_), .Y(new_n22205_));
  AOI21X1  g19769(.A0(new_n22160_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n22206_));
  OAI21X1  g19770(.A0(new_n22205_), .A1(new_n12486_), .B0(new_n22206_), .Y(new_n22207_));
  NAND2X1  g19771(.A(new_n22207_), .B(new_n12494_), .Y(new_n22208_));
  OAI21X1  g19772(.A0(new_n22201_), .A1(pi0618), .B0(pi1154), .Y(new_n22209_));
  AOI21X1  g19773(.A0(new_n22200_), .A1(pi0618), .B0(new_n22209_), .Y(new_n22210_));
  AOI21X1  g19774(.A0(new_n22160_), .A1(pi0618), .B0(pi1154), .Y(new_n22211_));
  OAI21X1  g19775(.A0(new_n22205_), .A1(pi0618), .B0(new_n22211_), .Y(new_n22212_));
  NAND2X1  g19776(.A(new_n22212_), .B(pi0627), .Y(new_n22213_));
  OAI22X1  g19777(.A0(new_n22213_), .A1(new_n22210_), .B0(new_n22208_), .B1(new_n22203_), .Y(new_n22214_));
  MX2X1    g19778(.A(new_n22214_), .B(new_n22200_), .S0(new_n11767_), .Y(new_n22215_));
  MX2X1    g19779(.A(new_n22201_), .B(new_n22140_), .S0(new_n12513_), .Y(new_n22216_));
  OAI21X1  g19780(.A0(new_n22216_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n22217_));
  AOI21X1  g19781(.A0(new_n22215_), .A1(new_n12509_), .B0(new_n22217_), .Y(new_n22218_));
  AOI21X1  g19782(.A0(new_n22212_), .A1(new_n22207_), .B0(new_n11767_), .Y(new_n22219_));
  AOI21X1  g19783(.A0(new_n22205_), .A1(new_n11767_), .B0(new_n22219_), .Y(new_n22220_));
  OAI21X1  g19784(.A0(new_n22140_), .A1(pi0619), .B0(pi1159), .Y(new_n22221_));
  AOI21X1  g19785(.A0(new_n22220_), .A1(pi0619), .B0(new_n22221_), .Y(new_n22222_));
  OR2X1    g19786(.A(new_n22222_), .B(pi0648), .Y(new_n22223_));
  OAI21X1  g19787(.A0(new_n22216_), .A1(pi0619), .B0(pi1159), .Y(new_n22224_));
  AOI21X1  g19788(.A0(new_n22215_), .A1(pi0619), .B0(new_n22224_), .Y(new_n22225_));
  OAI21X1  g19789(.A0(new_n22140_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n22226_));
  AOI21X1  g19790(.A0(new_n22220_), .A1(new_n12509_), .B0(new_n22226_), .Y(new_n22227_));
  OR2X1    g19791(.A(new_n22227_), .B(new_n12517_), .Y(new_n22228_));
  OAI22X1  g19792(.A0(new_n22228_), .A1(new_n22225_), .B0(new_n22223_), .B1(new_n22218_), .Y(new_n22229_));
  MX2X1    g19793(.A(new_n22229_), .B(new_n22215_), .S0(new_n11766_), .Y(new_n22230_));
  MX2X1    g19794(.A(new_n22216_), .B(new_n22140_), .S0(new_n12531_), .Y(new_n22231_));
  AOI21X1  g19795(.A0(new_n22231_), .A1(pi0626), .B0(pi0641), .Y(new_n22232_));
  OAI21X1  g19796(.A0(new_n22230_), .A1(pi0626), .B0(new_n22232_), .Y(new_n22233_));
  NOR2X1   g19797(.A(new_n22227_), .B(new_n22222_), .Y(new_n22234_));
  MX2X1    g19798(.A(new_n22234_), .B(new_n22220_), .S0(new_n11766_), .Y(new_n22235_));
  AOI21X1  g19799(.A0(new_n22140_), .A1(pi0626), .B0(new_n12543_), .Y(new_n22236_));
  OAI21X1  g19800(.A0(new_n22235_), .A1(pi0626), .B0(new_n22236_), .Y(new_n22237_));
  AND2X1   g19801(.A(new_n22237_), .B(new_n12548_), .Y(new_n22238_));
  AOI21X1  g19802(.A0(new_n22231_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n22239_));
  OAI21X1  g19803(.A0(new_n22230_), .A1(new_n12542_), .B0(new_n22239_), .Y(new_n22240_));
  AOI21X1  g19804(.A0(new_n22140_), .A1(new_n12542_), .B0(pi0641), .Y(new_n22241_));
  OAI21X1  g19805(.A0(new_n22235_), .A1(new_n12542_), .B0(new_n22241_), .Y(new_n22242_));
  AND2X1   g19806(.A(new_n22242_), .B(pi1158), .Y(new_n22243_));
  AOI22X1  g19807(.A0(new_n22243_), .A1(new_n22240_), .B0(new_n22238_), .B1(new_n22233_), .Y(new_n22244_));
  MX2X1    g19808(.A(new_n22244_), .B(new_n22230_), .S0(new_n11765_), .Y(new_n22245_));
  MX2X1    g19809(.A(new_n22235_), .B(new_n22160_), .S0(new_n12708_), .Y(new_n22246_));
  INVX1    g19810(.A(new_n22246_), .Y(new_n22247_));
  OAI21X1  g19811(.A0(new_n22247_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n22248_));
  AOI21X1  g19812(.A0(new_n22245_), .A1(new_n12554_), .B0(new_n22248_), .Y(new_n22249_));
  MX2X1    g19813(.A(new_n22231_), .B(new_n22140_), .S0(new_n12563_), .Y(new_n22250_));
  AOI21X1  g19814(.A0(new_n22160_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n22251_));
  OAI21X1  g19815(.A0(new_n22250_), .A1(new_n12554_), .B0(new_n22251_), .Y(new_n22252_));
  NAND2X1  g19816(.A(new_n22252_), .B(new_n12561_), .Y(new_n22253_));
  OAI21X1  g19817(.A0(new_n22247_), .A1(pi0628), .B0(pi1156), .Y(new_n22254_));
  AOI21X1  g19818(.A0(new_n22245_), .A1(pi0628), .B0(new_n22254_), .Y(new_n22255_));
  AOI21X1  g19819(.A0(new_n22160_), .A1(pi0628), .B0(pi1156), .Y(new_n22256_));
  OAI21X1  g19820(.A0(new_n22250_), .A1(pi0628), .B0(new_n22256_), .Y(new_n22257_));
  NAND2X1  g19821(.A(new_n22257_), .B(pi0629), .Y(new_n22258_));
  OAI22X1  g19822(.A0(new_n22258_), .A1(new_n22255_), .B0(new_n22253_), .B1(new_n22249_), .Y(new_n22259_));
  MX2X1    g19823(.A(new_n22259_), .B(new_n22245_), .S0(new_n11764_), .Y(new_n22260_));
  MX2X1    g19824(.A(new_n22246_), .B(new_n22160_), .S0(new_n12580_), .Y(new_n22261_));
  INVX1    g19825(.A(new_n22261_), .Y(new_n22262_));
  OAI21X1  g19826(.A0(new_n22262_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n22263_));
  AOI21X1  g19827(.A0(new_n22260_), .A1(new_n12577_), .B0(new_n22263_), .Y(new_n22264_));
  AND2X1   g19828(.A(new_n22250_), .B(new_n11764_), .Y(new_n22265_));
  AOI21X1  g19829(.A0(new_n22257_), .A1(new_n22252_), .B0(new_n11764_), .Y(new_n22266_));
  NOR2X1   g19830(.A(new_n22266_), .B(new_n22265_), .Y(new_n22267_));
  INVX1    g19831(.A(new_n22267_), .Y(new_n22268_));
  AOI21X1  g19832(.A0(new_n22160_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n22269_));
  OAI21X1  g19833(.A0(new_n22268_), .A1(new_n12577_), .B0(new_n22269_), .Y(new_n22270_));
  NAND2X1  g19834(.A(new_n22270_), .B(new_n12592_), .Y(new_n22271_));
  OAI21X1  g19835(.A0(new_n22262_), .A1(pi0647), .B0(pi1157), .Y(new_n22272_));
  AOI21X1  g19836(.A0(new_n22260_), .A1(pi0647), .B0(new_n22272_), .Y(new_n22273_));
  AOI21X1  g19837(.A0(new_n22160_), .A1(pi0647), .B0(pi1157), .Y(new_n22274_));
  OAI21X1  g19838(.A0(new_n22268_), .A1(pi0647), .B0(new_n22274_), .Y(new_n22275_));
  NAND2X1  g19839(.A(new_n22275_), .B(pi0630), .Y(new_n22276_));
  OAI22X1  g19840(.A0(new_n22276_), .A1(new_n22273_), .B0(new_n22271_), .B1(new_n22264_), .Y(new_n22277_));
  MX2X1    g19841(.A(new_n22277_), .B(new_n22260_), .S0(new_n11763_), .Y(new_n22278_));
  NAND2X1  g19842(.A(new_n22278_), .B(pi0644), .Y(new_n22279_));
  AND2X1   g19843(.A(new_n22275_), .B(new_n22270_), .Y(new_n22280_));
  MX2X1    g19844(.A(new_n22280_), .B(new_n22267_), .S0(new_n11763_), .Y(new_n22281_));
  AOI21X1  g19845(.A0(new_n22281_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n22282_));
  MX2X1    g19846(.A(new_n22261_), .B(new_n22160_), .S0(new_n12604_), .Y(new_n22283_));
  OAI21X1  g19847(.A0(new_n22140_), .A1(pi0644), .B0(new_n12608_), .Y(new_n22284_));
  AOI21X1  g19848(.A0(new_n22283_), .A1(pi0644), .B0(new_n22284_), .Y(new_n22285_));
  OR2X1    g19849(.A(new_n22285_), .B(new_n11762_), .Y(new_n22286_));
  AOI21X1  g19850(.A0(new_n22282_), .A1(new_n22279_), .B0(new_n22286_), .Y(new_n22287_));
  AND2X1   g19851(.A(new_n22281_), .B(pi0644), .Y(new_n22288_));
  OR2X1    g19852(.A(new_n22288_), .B(pi0715), .Y(new_n22289_));
  AOI21X1  g19853(.A0(new_n22278_), .A1(new_n12612_), .B0(new_n22289_), .Y(new_n22290_));
  OAI21X1  g19854(.A0(new_n22140_), .A1(new_n12612_), .B0(pi0715), .Y(new_n22291_));
  AOI21X1  g19855(.A0(new_n22283_), .A1(new_n12612_), .B0(new_n22291_), .Y(new_n22292_));
  OR2X1    g19856(.A(new_n22292_), .B(pi1160), .Y(new_n22293_));
  OAI21X1  g19857(.A0(new_n22293_), .A1(new_n22290_), .B0(pi0790), .Y(new_n22294_));
  OAI22X1  g19858(.A0(new_n22294_), .A1(new_n22287_), .B0(new_n22278_), .B1(pi0790), .Y(new_n22295_));
  MX2X1    g19859(.A(new_n22295_), .B(pi0199), .S0(po1038), .Y(po0356));
  AOI21X1  g19860(.A0(new_n12447_), .A1(new_n3103_), .B0(new_n7937_), .Y(new_n22297_));
  INVX1    g19861(.A(new_n22297_), .Y(new_n22298_));
  INVX1    g19862(.A(pi0606), .Y(new_n22299_));
  OR2X1    g19863(.A(new_n13564_), .B(pi0200), .Y(new_n22300_));
  AND2X1   g19864(.A(new_n22300_), .B(new_n13567_), .Y(new_n22301_));
  INVX1    g19865(.A(new_n22301_), .Y(new_n22302_));
  AOI21X1  g19866(.A0(new_n16615_), .A1(new_n7937_), .B0(pi0038), .Y(new_n22303_));
  OAI21X1  g19867(.A0(new_n12776_), .A1(new_n7937_), .B0(new_n22303_), .Y(new_n22304_));
  AOI21X1  g19868(.A0(new_n22304_), .A1(new_n22302_), .B0(new_n11770_), .Y(new_n22305_));
  NOR2X1   g19869(.A(new_n3103_), .B(new_n7937_), .Y(new_n22306_));
  NOR3X1   g19870(.A(new_n22306_), .B(new_n22305_), .C(new_n22299_), .Y(new_n22307_));
  AOI21X1  g19871(.A0(new_n22298_), .A1(new_n22299_), .B0(new_n22307_), .Y(new_n22308_));
  MX2X1    g19872(.A(new_n22308_), .B(new_n22297_), .S0(new_n12473_), .Y(new_n22309_));
  INVX1    g19873(.A(new_n22309_), .Y(new_n22310_));
  AOI21X1  g19874(.A0(new_n22298_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n22311_));
  OAI21X1  g19875(.A0(new_n22309_), .A1(new_n12462_), .B0(new_n22311_), .Y(new_n22312_));
  AOI21X1  g19876(.A0(new_n22298_), .A1(pi0609), .B0(pi1155), .Y(new_n22313_));
  OAI21X1  g19877(.A0(new_n22309_), .A1(pi0609), .B0(new_n22313_), .Y(new_n22314_));
  AND2X1   g19878(.A(new_n22314_), .B(new_n22312_), .Y(new_n22315_));
  MX2X1    g19879(.A(new_n22315_), .B(new_n22310_), .S0(new_n11768_), .Y(new_n22316_));
  NOR2X1   g19880(.A(new_n22316_), .B(pi0781), .Y(new_n22317_));
  INVX1    g19881(.A(new_n22316_), .Y(new_n22318_));
  AOI21X1  g19882(.A0(new_n22298_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n22319_));
  OAI21X1  g19883(.A0(new_n22318_), .A1(new_n12486_), .B0(new_n22319_), .Y(new_n22320_));
  AOI21X1  g19884(.A0(new_n22298_), .A1(pi0618), .B0(pi1154), .Y(new_n22321_));
  OAI21X1  g19885(.A0(new_n22318_), .A1(pi0618), .B0(new_n22321_), .Y(new_n22322_));
  AOI21X1  g19886(.A0(new_n22322_), .A1(new_n22320_), .B0(new_n11767_), .Y(new_n22323_));
  NOR2X1   g19887(.A(new_n22323_), .B(new_n22317_), .Y(new_n22324_));
  INVX1    g19888(.A(new_n22324_), .Y(new_n22325_));
  AOI21X1  g19889(.A0(new_n22298_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n22326_));
  OAI21X1  g19890(.A0(new_n22325_), .A1(new_n12509_), .B0(new_n22326_), .Y(new_n22327_));
  AOI21X1  g19891(.A0(new_n22298_), .A1(pi0619), .B0(pi1159), .Y(new_n22328_));
  OAI21X1  g19892(.A0(new_n22325_), .A1(pi0619), .B0(new_n22328_), .Y(new_n22329_));
  AND2X1   g19893(.A(new_n22329_), .B(new_n22327_), .Y(new_n22330_));
  MX2X1    g19894(.A(new_n22330_), .B(new_n22324_), .S0(new_n11766_), .Y(new_n22331_));
  MX2X1    g19895(.A(new_n22331_), .B(new_n22298_), .S0(new_n12708_), .Y(new_n22332_));
  OAI21X1  g19896(.A0(new_n12077_), .A1(pi0200), .B0(new_n13873_), .Y(new_n22333_));
  AOI21X1  g19897(.A0(new_n12384_), .A1(new_n7937_), .B0(pi0299), .Y(new_n22334_));
  OAI21X1  g19898(.A0(new_n12819_), .A1(new_n7937_), .B0(new_n22334_), .Y(new_n22335_));
  AOI21X1  g19899(.A0(new_n12393_), .A1(new_n7937_), .B0(new_n2933_), .Y(new_n22336_));
  OAI21X1  g19900(.A0(new_n12823_), .A1(new_n7937_), .B0(new_n22336_), .Y(new_n22337_));
  AOI21X1  g19901(.A0(new_n22337_), .A1(new_n22335_), .B0(new_n2939_), .Y(new_n22338_));
  OAI21X1  g19902(.A0(new_n12340_), .A1(new_n7937_), .B0(new_n2939_), .Y(new_n22339_));
  AOI21X1  g19903(.A0(new_n12435_), .A1(new_n7937_), .B0(new_n22339_), .Y(new_n22340_));
  OAI21X1  g19904(.A0(new_n22340_), .A1(new_n22338_), .B0(new_n2979_), .Y(new_n22341_));
  AOI21X1  g19905(.A0(new_n22341_), .A1(new_n22333_), .B0(new_n11770_), .Y(new_n22342_));
  OAI21X1  g19906(.A0(new_n3103_), .A1(new_n7937_), .B0(pi0643), .Y(new_n22343_));
  OAI22X1  g19907(.A0(new_n22343_), .A1(new_n22342_), .B0(new_n22297_), .B1(pi0643), .Y(new_n22344_));
  OAI21X1  g19908(.A0(new_n22297_), .A1(pi0625), .B0(pi1153), .Y(new_n22345_));
  AOI21X1  g19909(.A0(new_n22344_), .A1(pi0625), .B0(new_n22345_), .Y(new_n22346_));
  OAI21X1  g19910(.A0(new_n22297_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n22347_));
  AOI21X1  g19911(.A0(new_n22344_), .A1(new_n12363_), .B0(new_n22347_), .Y(new_n22348_));
  NOR2X1   g19912(.A(new_n22348_), .B(new_n22346_), .Y(new_n22349_));
  MX2X1    g19913(.A(new_n22349_), .B(new_n22344_), .S0(new_n11769_), .Y(new_n22350_));
  INVX1    g19914(.A(new_n22350_), .Y(new_n22351_));
  MX2X1    g19915(.A(new_n22351_), .B(new_n22297_), .S0(new_n12490_), .Y(new_n22352_));
  INVX1    g19916(.A(new_n22352_), .Y(new_n22353_));
  MX2X1    g19917(.A(new_n22353_), .B(new_n22298_), .S0(new_n12513_), .Y(new_n22354_));
  INVX1    g19918(.A(new_n22354_), .Y(new_n22355_));
  MX2X1    g19919(.A(new_n22355_), .B(new_n22297_), .S0(new_n12531_), .Y(new_n22356_));
  AND2X1   g19920(.A(new_n22297_), .B(new_n12563_), .Y(new_n22357_));
  AOI21X1  g19921(.A0(new_n22356_), .A1(new_n13356_), .B0(new_n22357_), .Y(new_n22358_));
  AOI21X1  g19922(.A0(new_n22298_), .A1(new_n12554_), .B0(new_n12555_), .Y(new_n22359_));
  INVX1    g19923(.A(new_n22359_), .Y(new_n22360_));
  AOI21X1  g19924(.A0(new_n22358_), .A1(pi0628), .B0(new_n22360_), .Y(new_n22361_));
  AND2X1   g19925(.A(new_n22361_), .B(new_n12561_), .Y(new_n22362_));
  AOI21X1  g19926(.A0(new_n22298_), .A1(pi0628), .B0(pi1156), .Y(new_n22363_));
  INVX1    g19927(.A(new_n22363_), .Y(new_n22364_));
  AOI21X1  g19928(.A0(new_n22358_), .A1(new_n12554_), .B0(new_n22364_), .Y(new_n22365_));
  AOI21X1  g19929(.A0(new_n22365_), .A1(pi0629), .B0(new_n22362_), .Y(new_n22366_));
  OAI21X1  g19930(.A0(new_n22332_), .A1(new_n14250_), .B0(new_n22366_), .Y(new_n22367_));
  INVX1    g19931(.A(pi0643), .Y(new_n22368_));
  NOR2X1   g19932(.A(new_n12440_), .B(new_n12141_), .Y(new_n22369_));
  AOI21X1  g19933(.A0(new_n13544_), .A1(new_n7937_), .B0(pi0038), .Y(new_n22370_));
  OAI21X1  g19934(.A0(new_n13542_), .A1(new_n7937_), .B0(new_n22370_), .Y(new_n22371_));
  OAI21X1  g19935(.A0(new_n22369_), .A1(new_n22333_), .B0(new_n22371_), .Y(new_n22372_));
  NOR4X1   g19936(.A(new_n10543_), .B(pi0606), .C(pi0100), .D(pi0087), .Y(new_n22373_));
  AOI21X1  g19937(.A0(new_n12787_), .A1(pi0039), .B0(new_n16667_), .Y(new_n22374_));
  NOR2X1   g19938(.A(new_n22374_), .B(pi0200), .Y(new_n22375_));
  OAI21X1  g19939(.A0(new_n13552_), .A1(pi0200), .B0(new_n2979_), .Y(new_n22376_));
  AOI21X1  g19940(.A0(new_n16738_), .A1(pi0200), .B0(new_n22376_), .Y(new_n22377_));
  AND2X1   g19941(.A(pi0200), .B(pi0038), .Y(new_n22378_));
  AND3X1   g19942(.A(new_n22378_), .B(new_n12276_), .C(new_n2939_), .Y(new_n22379_));
  OR4X1    g19943(.A(new_n22379_), .B(new_n22377_), .C(new_n11770_), .D(new_n22299_), .Y(new_n22380_));
  OAI22X1  g19944(.A0(new_n22380_), .A1(new_n22375_), .B0(new_n3103_), .B1(new_n7937_), .Y(new_n22381_));
  AOI21X1  g19945(.A0(new_n22373_), .A1(new_n22372_), .B0(new_n22381_), .Y(new_n22382_));
  NOR2X1   g19946(.A(new_n22382_), .B(new_n22368_), .Y(new_n22383_));
  AOI21X1  g19947(.A0(new_n22308_), .A1(new_n22368_), .B0(new_n22383_), .Y(new_n22384_));
  OAI21X1  g19948(.A0(new_n22308_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n22385_));
  AOI21X1  g19949(.A0(new_n22384_), .A1(new_n12363_), .B0(new_n22385_), .Y(new_n22386_));
  OR2X1    g19950(.A(new_n22346_), .B(pi0608), .Y(new_n22387_));
  OAI21X1  g19951(.A0(new_n22308_), .A1(pi0625), .B0(pi1153), .Y(new_n22388_));
  AOI21X1  g19952(.A0(new_n22384_), .A1(pi0625), .B0(new_n22388_), .Y(new_n22389_));
  OR2X1    g19953(.A(new_n22348_), .B(new_n12368_), .Y(new_n22390_));
  OAI22X1  g19954(.A0(new_n22390_), .A1(new_n22389_), .B0(new_n22387_), .B1(new_n22386_), .Y(new_n22391_));
  MX2X1    g19955(.A(new_n22391_), .B(new_n22384_), .S0(new_n11769_), .Y(new_n22392_));
  OAI21X1  g19956(.A0(new_n22351_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n22393_));
  AOI21X1  g19957(.A0(new_n22392_), .A1(new_n12462_), .B0(new_n22393_), .Y(new_n22394_));
  NAND2X1  g19958(.A(new_n22312_), .B(new_n12468_), .Y(new_n22395_));
  OAI21X1  g19959(.A0(new_n22351_), .A1(pi0609), .B0(pi1155), .Y(new_n22396_));
  AOI21X1  g19960(.A0(new_n22392_), .A1(pi0609), .B0(new_n22396_), .Y(new_n22397_));
  NAND2X1  g19961(.A(new_n22314_), .B(pi0660), .Y(new_n22398_));
  OAI22X1  g19962(.A0(new_n22398_), .A1(new_n22397_), .B0(new_n22395_), .B1(new_n22394_), .Y(new_n22399_));
  MX2X1    g19963(.A(new_n22399_), .B(new_n22392_), .S0(new_n11768_), .Y(new_n22400_));
  INVX1    g19964(.A(new_n22400_), .Y(new_n22401_));
  AOI21X1  g19965(.A0(new_n22353_), .A1(pi0618), .B0(pi1154), .Y(new_n22402_));
  OAI21X1  g19966(.A0(new_n22401_), .A1(pi0618), .B0(new_n22402_), .Y(new_n22403_));
  AND2X1   g19967(.A(new_n22320_), .B(new_n12494_), .Y(new_n22404_));
  AOI21X1  g19968(.A0(new_n22353_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n22405_));
  OAI21X1  g19969(.A0(new_n22401_), .A1(new_n12486_), .B0(new_n22405_), .Y(new_n22406_));
  AND2X1   g19970(.A(new_n22322_), .B(pi0627), .Y(new_n22407_));
  AOI22X1  g19971(.A0(new_n22407_), .A1(new_n22406_), .B0(new_n22404_), .B1(new_n22403_), .Y(new_n22408_));
  MX2X1    g19972(.A(new_n22408_), .B(new_n22401_), .S0(new_n11767_), .Y(new_n22409_));
  AOI21X1  g19973(.A0(new_n22354_), .A1(pi0619), .B0(pi1159), .Y(new_n22410_));
  OAI21X1  g19974(.A0(new_n22409_), .A1(pi0619), .B0(new_n22410_), .Y(new_n22411_));
  AND3X1   g19975(.A(new_n22411_), .B(new_n22327_), .C(new_n12517_), .Y(new_n22412_));
  AOI21X1  g19976(.A0(new_n22354_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n22413_));
  OAI21X1  g19977(.A0(new_n22409_), .A1(new_n12509_), .B0(new_n22413_), .Y(new_n22414_));
  AND3X1   g19978(.A(new_n22414_), .B(new_n22329_), .C(pi0648), .Y(new_n22415_));
  OR3X1    g19979(.A(new_n22415_), .B(new_n22412_), .C(new_n11766_), .Y(new_n22416_));
  AOI21X1  g19980(.A0(new_n22409_), .A1(new_n11766_), .B0(new_n13481_), .Y(new_n22417_));
  NAND2X1  g19981(.A(new_n22417_), .B(new_n22416_), .Y(new_n22418_));
  AOI21X1  g19982(.A0(new_n22297_), .A1(pi0626), .B0(new_n16218_), .Y(new_n22419_));
  OAI21X1  g19983(.A0(new_n22331_), .A1(pi0626), .B0(new_n22419_), .Y(new_n22420_));
  AOI21X1  g19984(.A0(new_n22297_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n22421_));
  OAI21X1  g19985(.A0(new_n22331_), .A1(new_n12542_), .B0(new_n22421_), .Y(new_n22422_));
  OR2X1    g19986(.A(new_n22356_), .B(new_n13439_), .Y(new_n22423_));
  NAND3X1  g19987(.A(new_n22423_), .B(new_n22422_), .C(new_n22420_), .Y(new_n22424_));
  AOI21X1  g19988(.A0(new_n22424_), .A1(pi0788), .B0(new_n14125_), .Y(new_n22425_));
  AOI22X1  g19989(.A0(new_n22425_), .A1(new_n22418_), .B0(new_n22367_), .B1(pi0792), .Y(new_n22426_));
  NAND2X1  g19990(.A(new_n22297_), .B(new_n12580_), .Y(new_n22427_));
  OAI21X1  g19991(.A0(new_n22332_), .A1(new_n12580_), .B0(new_n22427_), .Y(new_n22428_));
  OR2X1    g19992(.A(new_n22358_), .B(pi0792), .Y(new_n22429_));
  OAI21X1  g19993(.A0(new_n22365_), .A1(new_n22361_), .B0(pi0792), .Y(new_n22430_));
  AND2X1   g19994(.A(new_n22430_), .B(new_n22429_), .Y(new_n22431_));
  MX2X1    g19995(.A(new_n22431_), .B(new_n22298_), .S0(new_n12577_), .Y(new_n22432_));
  AND3X1   g19996(.A(new_n22430_), .B(new_n22429_), .C(new_n12577_), .Y(new_n22433_));
  AOI21X1  g19997(.A0(new_n22298_), .A1(pi0647), .B0(pi1157), .Y(new_n22434_));
  INVX1    g19998(.A(new_n22434_), .Y(new_n22435_));
  OR3X1    g19999(.A(new_n22435_), .B(new_n22433_), .C(new_n12592_), .Y(new_n22436_));
  OAI21X1  g20000(.A0(new_n22432_), .A1(new_n14242_), .B0(new_n22436_), .Y(new_n22437_));
  AOI21X1  g20001(.A0(new_n22428_), .A1(new_n14326_), .B0(new_n22437_), .Y(new_n22438_));
  OAI22X1  g20002(.A0(new_n22438_), .A1(new_n11763_), .B0(new_n22426_), .B1(new_n14121_), .Y(new_n22439_));
  AOI21X1  g20003(.A0(new_n22430_), .A1(new_n22429_), .B0(pi0787), .Y(new_n22440_));
  OAI22X1  g20004(.A0(new_n22435_), .A1(new_n22433_), .B0(new_n22432_), .B1(new_n12578_), .Y(new_n22441_));
  AOI21X1  g20005(.A0(new_n22441_), .A1(pi0787), .B0(new_n22440_), .Y(new_n22442_));
  AOI21X1  g20006(.A0(new_n22442_), .A1(pi0644), .B0(pi0715), .Y(new_n22443_));
  OAI21X1  g20007(.A0(new_n22439_), .A1(pi0644), .B0(new_n22443_), .Y(new_n22444_));
  MX2X1    g20008(.A(new_n22428_), .B(new_n22297_), .S0(new_n12604_), .Y(new_n22445_));
  AOI21X1  g20009(.A0(new_n22298_), .A1(pi0644), .B0(new_n12608_), .Y(new_n22446_));
  OAI21X1  g20010(.A0(new_n22445_), .A1(pi0644), .B0(new_n22446_), .Y(new_n22447_));
  AND2X1   g20011(.A(new_n22447_), .B(new_n11762_), .Y(new_n22448_));
  AOI21X1  g20012(.A0(new_n22442_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n22449_));
  OAI21X1  g20013(.A0(new_n22439_), .A1(new_n12612_), .B0(new_n22449_), .Y(new_n22450_));
  AOI21X1  g20014(.A0(new_n22298_), .A1(new_n12612_), .B0(pi0715), .Y(new_n22451_));
  OAI21X1  g20015(.A0(new_n22445_), .A1(new_n12612_), .B0(new_n22451_), .Y(new_n22452_));
  AND2X1   g20016(.A(new_n22452_), .B(pi1160), .Y(new_n22453_));
  AOI22X1  g20017(.A0(new_n22453_), .A1(new_n22450_), .B0(new_n22448_), .B1(new_n22444_), .Y(new_n22454_));
  MX2X1    g20018(.A(new_n22454_), .B(new_n22439_), .S0(new_n12766_), .Y(new_n22455_));
  MX2X1    g20019(.A(new_n22455_), .B(pi0200), .S0(po1038), .Y(po0357));
  INVX1    g20020(.A(pi0201), .Y(new_n22457_));
  NAND2X1  g20021(.A(pi0237), .B(pi0233), .Y(new_n22458_));
  AOI21X1  g20022(.A0(new_n4975_), .A1(pi0332), .B0(pi0059), .Y(new_n22459_));
  AOI21X1  g20023(.A0(pi0332), .A1(pi0074), .B0(pi0055), .Y(new_n22460_));
  INVX1    g20024(.A(new_n22460_), .Y(new_n22461_));
  MX2X1    g20025(.A(pi0587), .B(pi0947), .S0(pi0299), .Y(new_n22462_));
  MX2X1    g20026(.A(new_n22462_), .B(new_n5018_), .S0(pi0468), .Y(new_n22463_));
  AND3X1   g20027(.A(new_n22463_), .B(new_n8232_), .C(new_n2499_), .Y(new_n22464_));
  OAI21X1  g20028(.A0(new_n22464_), .A1(pi0332), .B0(new_n5839_), .Y(new_n22465_));
  OAI21X1  g20029(.A0(new_n5340_), .A1(new_n2986_), .B0(new_n2444_), .Y(new_n22466_));
  AOI22X1  g20030(.A0(new_n22466_), .A1(new_n11153_), .B0(new_n3086_), .B1(pi0332), .Y(new_n22467_));
  AOI21X1  g20031(.A0(new_n22467_), .A1(new_n22465_), .B0(pi0074), .Y(new_n22468_));
  OR4X1    g20032(.A(new_n5314_), .B(new_n3105_), .C(new_n2985_), .D(new_n2536_), .Y(new_n22469_));
  NAND3X1  g20033(.A(new_n22469_), .B(new_n2444_), .C(pi0055), .Y(new_n22470_));
  AND2X1   g20034(.A(new_n22470_), .B(new_n3123_), .Y(new_n22471_));
  OAI21X1  g20035(.A0(new_n22468_), .A1(new_n22461_), .B0(new_n22471_), .Y(new_n22472_));
  AOI21X1  g20036(.A0(new_n22469_), .A1(new_n2444_), .B0(new_n8381_), .Y(new_n22473_));
  AOI21X1  g20037(.A0(new_n8381_), .A1(pi0332), .B0(new_n3127_), .Y(new_n22474_));
  INVX1    g20038(.A(new_n22474_), .Y(new_n22475_));
  OAI21X1  g20039(.A0(new_n22475_), .A1(new_n22473_), .B0(new_n2436_), .Y(new_n22476_));
  AOI21X1  g20040(.A0(new_n22472_), .A1(new_n22459_), .B0(new_n22476_), .Y(new_n22477_));
  AOI21X1  g20041(.A0(pi0332), .A1(pi0057), .B0(new_n22477_), .Y(new_n22478_));
  NOR2X1   g20042(.A(new_n5018_), .B(pi0332), .Y(new_n22479_));
  NOR2X1   g20043(.A(new_n22479_), .B(pi0947), .Y(new_n22480_));
  INVX1    g20044(.A(new_n22480_), .Y(new_n22481_));
  AND3X1   g20045(.A(pi0332), .B(pi0210), .C(pi0096), .Y(new_n22482_));
  NOR2X1   g20046(.A(pi0841), .B(pi0070), .Y(new_n22483_));
  MX2X1    g20047(.A(new_n22483_), .B(pi0070), .S0(new_n2455_), .Y(new_n22484_));
  NOR2X1   g20048(.A(pi0096), .B(pi0032), .Y(new_n22485_));
  AOI21X1  g20049(.A0(new_n22485_), .A1(pi0070), .B0(pi0332), .Y(new_n22486_));
  INVX1    g20050(.A(new_n22486_), .Y(new_n22487_));
  AOI21X1  g20051(.A0(new_n22484_), .A1(new_n2777_), .B0(new_n22487_), .Y(new_n22488_));
  OR3X1    g20052(.A(new_n22488_), .B(new_n22482_), .C(new_n5023_), .Y(new_n22489_));
  AOI21X1  g20053(.A0(new_n22489_), .A1(new_n5018_), .B0(new_n22481_), .Y(new_n22490_));
  MX2X1    g20054(.A(new_n22488_), .B(new_n2444_), .S0(pi0468), .Y(new_n22491_));
  AND2X1   g20055(.A(new_n22491_), .B(new_n5348_), .Y(new_n22492_));
  INVX1    g20056(.A(new_n22492_), .Y(new_n22493_));
  NOR2X1   g20057(.A(new_n22488_), .B(new_n22482_), .Y(new_n22494_));
  INVX1    g20058(.A(new_n22494_), .Y(new_n22495_));
  AOI21X1  g20059(.A0(new_n22495_), .A1(new_n5018_), .B0(new_n5362_), .Y(new_n22496_));
  AOI21X1  g20060(.A0(new_n22496_), .A1(new_n22493_), .B0(new_n22490_), .Y(new_n22497_));
  INVX1    g20061(.A(new_n22497_), .Y(new_n22498_));
  INVX1    g20062(.A(new_n22482_), .Y(new_n22499_));
  NOR4X1   g20063(.A(new_n2691_), .B(new_n2689_), .C(pi0095), .D(pi0040), .Y(new_n22500_));
  OAI21X1  g20064(.A0(new_n22500_), .A1(pi0070), .B0(new_n22485_), .Y(new_n22501_));
  INVX1    g20065(.A(new_n22484_), .Y(new_n22502_));
  OAI21X1  g20066(.A0(pi0841), .A1(pi0070), .B0(pi0032), .Y(new_n22503_));
  NAND3X1  g20067(.A(new_n22503_), .B(new_n2746_), .C(new_n2523_), .Y(new_n22504_));
  OR3X1    g20068(.A(new_n22504_), .B(pi0051), .C(pi0035), .Y(new_n22505_));
  OAI21X1  g20069(.A0(new_n22505_), .A1(new_n2506_), .B0(new_n22502_), .Y(new_n22506_));
  AOI21X1  g20070(.A0(new_n22506_), .A1(new_n2777_), .B0(pi0332), .Y(new_n22507_));
  OAI21X1  g20071(.A0(new_n22501_), .A1(new_n2777_), .B0(new_n22507_), .Y(new_n22508_));
  AND2X1   g20072(.A(new_n22508_), .B(new_n22499_), .Y(new_n22509_));
  AOI21X1  g20073(.A0(new_n22509_), .A1(new_n5048_), .B0(new_n5348_), .Y(new_n22510_));
  MX2X1    g20074(.A(new_n22508_), .B(pi0332), .S0(pi0468), .Y(new_n22511_));
  NOR2X1   g20075(.A(new_n22511_), .B(new_n5018_), .Y(new_n22512_));
  OAI21X1  g20076(.A0(new_n22509_), .A1(new_n5348_), .B0(pi0947), .Y(new_n22513_));
  OAI22X1  g20077(.A0(new_n22513_), .A1(new_n22512_), .B0(new_n22510_), .B1(new_n22481_), .Y(new_n22514_));
  MX2X1    g20078(.A(new_n22514_), .B(new_n22498_), .S0(new_n3105_), .Y(new_n22515_));
  OR2X1    g20079(.A(new_n22515_), .B(new_n8381_), .Y(new_n22516_));
  AOI21X1  g20080(.A0(new_n22497_), .A1(new_n8381_), .B0(new_n3127_), .Y(new_n22517_));
  INVX1    g20081(.A(new_n2456_), .Y(new_n22518_));
  NAND2X1  g20082(.A(new_n2517_), .B(new_n2499_), .Y(new_n22519_));
  NOR3X1   g20083(.A(new_n22519_), .B(new_n22518_), .C(pi0095), .Y(new_n22520_));
  OAI21X1  g20084(.A0(new_n22520_), .A1(pi0070), .B0(new_n22485_), .Y(new_n22521_));
  OAI21X1  g20085(.A0(new_n22519_), .A1(new_n22504_), .B0(new_n22502_), .Y(new_n22522_));
  AOI21X1  g20086(.A0(new_n22522_), .A1(new_n2777_), .B0(pi0332), .Y(new_n22523_));
  OAI21X1  g20087(.A0(new_n22521_), .A1(new_n2777_), .B0(new_n22523_), .Y(new_n22524_));
  AND3X1   g20088(.A(new_n22524_), .B(new_n22499_), .C(new_n5048_), .Y(new_n22525_));
  OAI21X1  g20089(.A0(new_n22525_), .A1(new_n5348_), .B0(new_n22480_), .Y(new_n22526_));
  MX2X1    g20090(.A(new_n22524_), .B(pi0332), .S0(pi0468), .Y(new_n22527_));
  NAND2X1  g20091(.A(new_n22524_), .B(new_n22499_), .Y(new_n22528_));
  AOI21X1  g20092(.A0(new_n22528_), .A1(new_n5018_), .B0(new_n5362_), .Y(new_n22529_));
  OAI21X1  g20093(.A0(new_n22527_), .A1(new_n5018_), .B0(new_n22529_), .Y(new_n22530_));
  AND3X1   g20094(.A(new_n22530_), .B(new_n22526_), .C(pi0299), .Y(new_n22531_));
  AOI21X1  g20095(.A0(new_n22522_), .A1(new_n2954_), .B0(pi0332), .Y(new_n22532_));
  OAI21X1  g20096(.A0(new_n22521_), .A1(new_n2954_), .B0(new_n22532_), .Y(new_n22533_));
  NAND3X1  g20097(.A(pi0332), .B(pi0198), .C(pi0096), .Y(new_n22534_));
  AND2X1   g20098(.A(new_n22534_), .B(new_n22533_), .Y(new_n22535_));
  AOI21X1  g20099(.A0(new_n22535_), .A1(new_n5048_), .B0(new_n5348_), .Y(new_n22536_));
  OR3X1    g20100(.A(new_n22536_), .B(new_n22479_), .C(pi0587), .Y(new_n22537_));
  AOI21X1  g20101(.A0(new_n22534_), .A1(new_n22533_), .B0(new_n5348_), .Y(new_n22538_));
  OAI21X1  g20102(.A0(new_n8621_), .A1(new_n2444_), .B0(new_n5348_), .Y(new_n22539_));
  AOI21X1  g20103(.A0(new_n22533_), .A1(new_n8621_), .B0(new_n22539_), .Y(new_n22540_));
  OR3X1    g20104(.A(new_n22540_), .B(new_n22538_), .C(new_n5354_), .Y(new_n22541_));
  AND3X1   g20105(.A(new_n22541_), .B(new_n22537_), .C(new_n2933_), .Y(new_n22542_));
  OAI21X1  g20106(.A0(new_n22542_), .A1(new_n22531_), .B0(new_n5839_), .Y(new_n22543_));
  AND2X1   g20107(.A(new_n22514_), .B(pi0299), .Y(new_n22544_));
  NOR2X1   g20108(.A(new_n22479_), .B(pi0587), .Y(new_n22545_));
  AOI21X1  g20109(.A0(new_n22506_), .A1(new_n2954_), .B0(pi0332), .Y(new_n22546_));
  OAI21X1  g20110(.A0(new_n22501_), .A1(new_n2954_), .B0(new_n22546_), .Y(new_n22547_));
  AND3X1   g20111(.A(new_n22547_), .B(new_n22534_), .C(new_n5048_), .Y(new_n22548_));
  OAI21X1  g20112(.A0(new_n22548_), .A1(new_n5348_), .B0(new_n22545_), .Y(new_n22549_));
  AOI21X1  g20113(.A0(new_n22547_), .A1(new_n22534_), .B0(new_n5348_), .Y(new_n22550_));
  AOI21X1  g20114(.A0(new_n22547_), .A1(new_n8621_), .B0(new_n22539_), .Y(new_n22551_));
  OR3X1    g20115(.A(new_n22551_), .B(new_n22550_), .C(new_n5354_), .Y(new_n22552_));
  AOI21X1  g20116(.A0(new_n22552_), .A1(new_n22549_), .B0(pi0299), .Y(new_n22553_));
  OR3X1    g20117(.A(new_n22553_), .B(new_n22544_), .C(new_n11154_), .Y(new_n22554_));
  AOI21X1  g20118(.A0(new_n22554_), .A1(new_n22543_), .B0(pi0074), .Y(new_n22555_));
  NOR2X1   g20119(.A(new_n22497_), .B(new_n2933_), .Y(new_n22556_));
  AND2X1   g20120(.A(pi0198), .B(pi0096), .Y(new_n22557_));
  AOI21X1  g20121(.A0(new_n22484_), .A1(new_n2954_), .B0(new_n22487_), .Y(new_n22558_));
  AOI21X1  g20122(.A0(new_n22557_), .A1(pi0332), .B0(new_n22558_), .Y(new_n22559_));
  NOR2X1   g20123(.A(new_n22559_), .B(new_n5348_), .Y(new_n22560_));
  OR3X1    g20124(.A(new_n22558_), .B(new_n5345_), .C(new_n5352_), .Y(new_n22561_));
  AND2X1   g20125(.A(new_n22561_), .B(new_n22479_), .Y(new_n22562_));
  OR4X1    g20126(.A(new_n22562_), .B(new_n22560_), .C(new_n5345_), .D(pi0299), .Y(new_n22563_));
  OAI21X1  g20127(.A0(new_n3086_), .A1(pi0074), .B0(new_n22563_), .Y(new_n22564_));
  OAI21X1  g20128(.A0(new_n22564_), .A1(new_n22556_), .B0(new_n3107_), .Y(new_n22565_));
  AOI21X1  g20129(.A0(new_n22515_), .A1(pi0055), .B0(new_n4975_), .Y(new_n22566_));
  OAI21X1  g20130(.A0(new_n22565_), .A1(new_n22555_), .B0(new_n22566_), .Y(new_n22567_));
  AOI21X1  g20131(.A0(new_n22497_), .A1(new_n4975_), .B0(pi0059), .Y(new_n22568_));
  AOI22X1  g20132(.A0(new_n22568_), .A1(new_n22567_), .B0(new_n22517_), .B1(new_n22516_), .Y(new_n22569_));
  MX2X1    g20133(.A(new_n22569_), .B(new_n22497_), .S0(pi0057), .Y(new_n22570_));
  MX2X1    g20134(.A(new_n22570_), .B(new_n22478_), .S0(new_n22458_), .Y(new_n22571_));
  INVX1    g20135(.A(new_n11660_), .Y(new_n22572_));
  AOI21X1  g20136(.A0(new_n22557_), .A1(new_n5319_), .B0(new_n22572_), .Y(new_n22573_));
  AOI21X1  g20137(.A0(pi0210), .A1(pi0096), .B0(new_n11660_), .Y(new_n22574_));
  NOR2X1   g20138(.A(new_n11660_), .B(new_n5310_), .Y(new_n22575_));
  NOR4X1   g20139(.A(new_n22575_), .B(new_n22574_), .C(new_n22573_), .D(new_n22458_), .Y(new_n22576_));
  MX2X1    g20140(.A(new_n22576_), .B(new_n22571_), .S0(new_n22457_), .Y(po0358));
  INVX1    g20141(.A(pi0202), .Y(new_n22578_));
  INVX1    g20142(.A(pi0237), .Y(new_n22579_));
  OR2X1    g20143(.A(new_n22579_), .B(pi0233), .Y(new_n22580_));
  MX2X1    g20144(.A(new_n22570_), .B(new_n22478_), .S0(new_n22580_), .Y(new_n22581_));
  NOR4X1   g20145(.A(new_n22580_), .B(new_n22575_), .C(new_n22574_), .D(new_n22573_), .Y(new_n22582_));
  MX2X1    g20146(.A(new_n22582_), .B(new_n22581_), .S0(new_n22578_), .Y(po0359));
  INVX1    g20147(.A(pi0203), .Y(new_n22584_));
  OR2X1    g20148(.A(pi0237), .B(pi0233), .Y(new_n22585_));
  MX2X1    g20149(.A(new_n22570_), .B(new_n22478_), .S0(new_n22585_), .Y(new_n22586_));
  NOR4X1   g20150(.A(new_n22585_), .B(new_n22575_), .C(new_n22574_), .D(new_n22573_), .Y(new_n22587_));
  MX2X1    g20151(.A(new_n22587_), .B(new_n22586_), .S0(new_n22584_), .Y(po0360));
  INVX1    g20152(.A(pi0204), .Y(new_n22589_));
  MX2X1    g20153(.A(new_n5020_), .B(pi0602), .S0(new_n8621_), .Y(new_n22590_));
  MX2X1    g20154(.A(new_n22590_), .B(new_n5105_), .S0(pi0299), .Y(new_n22591_));
  AOI21X1  g20155(.A0(new_n22591_), .A1(new_n2987_), .B0(pi0332), .Y(new_n22592_));
  NOR2X1   g20156(.A(pi0602), .B(pi0299), .Y(new_n22593_));
  OAI21X1  g20157(.A0(pi0907), .A1(new_n2933_), .B0(new_n8621_), .Y(new_n22594_));
  OAI22X1  g20158(.A0(new_n22594_), .A1(new_n22593_), .B0(new_n5262_), .B1(new_n8621_), .Y(new_n22595_));
  NAND3X1  g20159(.A(new_n22595_), .B(new_n8232_), .C(new_n2499_), .Y(new_n22596_));
  AND2X1   g20160(.A(new_n22596_), .B(new_n2444_), .Y(new_n22597_));
  OAI22X1  g20161(.A0(new_n22597_), .A1(new_n5840_), .B0(new_n22592_), .B1(new_n11154_), .Y(new_n22598_));
  OAI21X1  g20162(.A0(new_n3085_), .A1(new_n2444_), .B0(new_n22460_), .Y(new_n22599_));
  AOI21X1  g20163(.A0(new_n22598_), .A1(new_n4982_), .B0(new_n22599_), .Y(new_n22600_));
  NAND2X1  g20164(.A(new_n5105_), .B(new_n3104_), .Y(new_n22601_));
  OAI21X1  g20165(.A0(new_n22601_), .A1(new_n2986_), .B0(new_n2444_), .Y(new_n22602_));
  OAI21X1  g20166(.A0(new_n22602_), .A1(new_n3107_), .B0(new_n3123_), .Y(new_n22603_));
  OAI21X1  g20167(.A0(new_n22603_), .A1(new_n22600_), .B0(new_n22459_), .Y(new_n22604_));
  AOI21X1  g20168(.A0(new_n22602_), .A1(new_n5306_), .B0(new_n22475_), .Y(new_n22605_));
  NOR2X1   g20169(.A(new_n22605_), .B(pi0057), .Y(new_n22606_));
  AOI22X1  g20170(.A0(new_n22606_), .A1(new_n22604_), .B0(pi0332), .B1(pi0057), .Y(new_n22607_));
  AOI21X1  g20171(.A0(new_n5262_), .A1(new_n2444_), .B0(pi0907), .Y(new_n22608_));
  INVX1    g20172(.A(new_n22608_), .Y(new_n22609_));
  AOI21X1  g20173(.A0(new_n22489_), .A1(new_n5020_), .B0(new_n22609_), .Y(new_n22610_));
  AND2X1   g20174(.A(new_n22491_), .B(new_n5262_), .Y(new_n22611_));
  INVX1    g20175(.A(new_n22611_), .Y(new_n22612_));
  AOI21X1  g20176(.A0(new_n22495_), .A1(new_n5020_), .B0(new_n5277_), .Y(new_n22613_));
  AOI21X1  g20177(.A0(new_n22613_), .A1(new_n22612_), .B0(new_n22610_), .Y(new_n22614_));
  INVX1    g20178(.A(new_n22614_), .Y(new_n22615_));
  NOR2X1   g20179(.A(new_n22511_), .B(new_n5020_), .Y(new_n22616_));
  OAI21X1  g20180(.A0(new_n22509_), .A1(new_n5262_), .B0(pi0907), .Y(new_n22617_));
  OAI21X1  g20181(.A0(new_n11863_), .A1(new_n2444_), .B0(pi0680), .Y(new_n22618_));
  AOI21X1  g20182(.A0(new_n22509_), .A1(new_n5048_), .B0(new_n22618_), .Y(new_n22619_));
  OAI22X1  g20183(.A0(new_n22619_), .A1(new_n22609_), .B0(new_n22617_), .B1(new_n22616_), .Y(new_n22620_));
  MX2X1    g20184(.A(new_n22620_), .B(new_n22615_), .S0(new_n3105_), .Y(new_n22621_));
  OR2X1    g20185(.A(new_n22621_), .B(new_n8381_), .Y(new_n22622_));
  AOI21X1  g20186(.A0(new_n22614_), .A1(new_n8381_), .B0(new_n3127_), .Y(new_n22623_));
  AOI21X1  g20187(.A0(new_n22557_), .A1(new_n5020_), .B0(new_n2444_), .Y(new_n22624_));
  OR2X1    g20188(.A(new_n22624_), .B(pi0299), .Y(new_n22625_));
  AND3X1   g20189(.A(new_n22547_), .B(new_n22534_), .C(new_n5197_), .Y(new_n22626_));
  OAI22X1  g20190(.A0(new_n22626_), .A1(new_n22625_), .B0(new_n22620_), .B1(new_n2933_), .Y(new_n22627_));
  NAND2X1  g20191(.A(new_n22627_), .B(new_n11153_), .Y(new_n22628_));
  AOI21X1  g20192(.A0(new_n22535_), .A1(new_n5197_), .B0(new_n22625_), .Y(new_n22629_));
  OAI21X1  g20193(.A0(new_n22525_), .A1(new_n5262_), .B0(new_n22608_), .Y(new_n22630_));
  AOI21X1  g20194(.A0(new_n22528_), .A1(new_n5020_), .B0(new_n5277_), .Y(new_n22631_));
  OAI21X1  g20195(.A0(new_n22527_), .A1(new_n5020_), .B0(new_n22631_), .Y(new_n22632_));
  AND3X1   g20196(.A(new_n22632_), .B(new_n22630_), .C(pi0299), .Y(new_n22633_));
  OAI21X1  g20197(.A0(new_n22633_), .A1(new_n22629_), .B0(new_n5839_), .Y(new_n22634_));
  AOI21X1  g20198(.A0(new_n22634_), .A1(new_n22628_), .B0(pi0074), .Y(new_n22635_));
  NOR2X1   g20199(.A(new_n22614_), .B(new_n2933_), .Y(new_n22636_));
  AOI21X1  g20200(.A0(new_n22590_), .A1(new_n22559_), .B0(new_n22624_), .Y(new_n22637_));
  OAI22X1  g20201(.A0(new_n22637_), .A1(pi0299), .B0(new_n3086_), .B1(pi0074), .Y(new_n22638_));
  OAI21X1  g20202(.A0(new_n22638_), .A1(new_n22636_), .B0(new_n3107_), .Y(new_n22639_));
  AOI21X1  g20203(.A0(new_n22621_), .A1(pi0055), .B0(new_n4975_), .Y(new_n22640_));
  OAI21X1  g20204(.A0(new_n22639_), .A1(new_n22635_), .B0(new_n22640_), .Y(new_n22641_));
  AOI21X1  g20205(.A0(new_n22614_), .A1(new_n4975_), .B0(pi0059), .Y(new_n22642_));
  AOI22X1  g20206(.A0(new_n22642_), .A1(new_n22641_), .B0(new_n22623_), .B1(new_n22622_), .Y(new_n22643_));
  MX2X1    g20207(.A(new_n22643_), .B(new_n22614_), .S0(pi0057), .Y(new_n22644_));
  MX2X1    g20208(.A(new_n22644_), .B(new_n22607_), .S0(new_n22458_), .Y(new_n22645_));
  AOI21X1  g20209(.A0(new_n22557_), .A1(new_n5197_), .B0(new_n22572_), .Y(new_n22646_));
  NOR2X1   g20210(.A(new_n11660_), .B(new_n5105_), .Y(new_n22647_));
  NOR4X1   g20211(.A(new_n22647_), .B(new_n22646_), .C(new_n22574_), .D(new_n22458_), .Y(new_n22648_));
  MX2X1    g20212(.A(new_n22648_), .B(new_n22645_), .S0(new_n22589_), .Y(po0361));
  INVX1    g20213(.A(pi0205), .Y(new_n22650_));
  MX2X1    g20214(.A(new_n22644_), .B(new_n22607_), .S0(new_n22580_), .Y(new_n22651_));
  NOR4X1   g20215(.A(new_n22647_), .B(new_n22646_), .C(new_n22580_), .D(new_n22574_), .Y(new_n22652_));
  MX2X1    g20216(.A(new_n22652_), .B(new_n22651_), .S0(new_n22650_), .Y(po0362));
  INVX1    g20217(.A(pi0206), .Y(new_n22654_));
  INVX1    g20218(.A(pi0233), .Y(new_n22655_));
  OR2X1    g20219(.A(pi0237), .B(new_n22655_), .Y(new_n22656_));
  MX2X1    g20220(.A(new_n22644_), .B(new_n22607_), .S0(new_n22656_), .Y(new_n22657_));
  NOR4X1   g20221(.A(new_n22656_), .B(new_n22647_), .C(new_n22646_), .D(new_n22574_), .Y(new_n22658_));
  MX2X1    g20222(.A(new_n22658_), .B(new_n22657_), .S0(new_n22654_), .Y(po0363));
  INVX1    g20223(.A(pi0207), .Y(new_n22660_));
  INVX1    g20224(.A(pi0623), .Y(new_n22661_));
  AND2X1   g20225(.A(new_n12447_), .B(new_n3103_), .Y(new_n22662_));
  INVX1    g20226(.A(new_n22662_), .Y(new_n22663_));
  AND2X1   g20227(.A(new_n13568_), .B(new_n3103_), .Y(new_n22664_));
  MX2X1    g20228(.A(new_n22664_), .B(new_n22662_), .S0(new_n12473_), .Y(new_n22665_));
  AOI21X1  g20229(.A0(new_n13568_), .A1(new_n3103_), .B0(new_n12473_), .Y(new_n22666_));
  AOI22X1  g20230(.A0(new_n22666_), .A1(new_n12462_), .B0(new_n12481_), .B1(new_n22663_), .Y(new_n22667_));
  AOI22X1  g20231(.A0(new_n22666_), .A1(pi0609), .B0(new_n12472_), .B1(new_n22663_), .Y(new_n22668_));
  MX2X1    g20232(.A(new_n22668_), .B(new_n22667_), .S0(new_n12463_), .Y(new_n22669_));
  MX2X1    g20233(.A(new_n22669_), .B(new_n22665_), .S0(new_n11768_), .Y(new_n22670_));
  OR2X1    g20234(.A(new_n22670_), .B(pi0781), .Y(new_n22671_));
  OAI21X1  g20235(.A0(new_n22663_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n22672_));
  AOI21X1  g20236(.A0(new_n22670_), .A1(new_n12486_), .B0(new_n22672_), .Y(new_n22673_));
  OAI21X1  g20237(.A0(new_n22663_), .A1(pi0618), .B0(pi1154), .Y(new_n22674_));
  AOI21X1  g20238(.A0(new_n22670_), .A1(pi0618), .B0(new_n22674_), .Y(new_n22675_));
  OAI21X1  g20239(.A0(new_n22675_), .A1(new_n22673_), .B0(pi0781), .Y(new_n22676_));
  AND2X1   g20240(.A(new_n22676_), .B(new_n22671_), .Y(new_n22677_));
  INVX1    g20241(.A(new_n22677_), .Y(new_n22678_));
  AOI21X1  g20242(.A0(new_n22662_), .A1(pi0619), .B0(pi1159), .Y(new_n22679_));
  OAI21X1  g20243(.A0(new_n22678_), .A1(pi0619), .B0(new_n22679_), .Y(new_n22680_));
  AOI21X1  g20244(.A0(new_n22662_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n22681_));
  OAI21X1  g20245(.A0(new_n22678_), .A1(new_n12509_), .B0(new_n22681_), .Y(new_n22682_));
  AND2X1   g20246(.A(new_n22682_), .B(new_n22680_), .Y(new_n22683_));
  MX2X1    g20247(.A(new_n22683_), .B(new_n22677_), .S0(new_n11766_), .Y(new_n22684_));
  AND3X1   g20248(.A(new_n12708_), .B(new_n12447_), .C(new_n3103_), .Y(new_n22685_));
  AOI21X1  g20249(.A0(new_n22684_), .A1(new_n16140_), .B0(new_n22685_), .Y(new_n22686_));
  MX2X1    g20250(.A(new_n22686_), .B(new_n22663_), .S0(new_n12580_), .Y(new_n22687_));
  INVX1    g20251(.A(new_n22687_), .Y(new_n22688_));
  NAND2X1  g20252(.A(new_n16617_), .B(new_n3103_), .Y(new_n22689_));
  OR4X1    g20253(.A(new_n22689_), .B(new_n14039_), .C(new_n14034_), .D(new_n12473_), .Y(new_n22690_));
  NOR4X1   g20254(.A(new_n22690_), .B(new_n14036_), .C(new_n12708_), .D(new_n12580_), .Y(new_n22691_));
  OAI21X1  g20255(.A0(new_n22691_), .A1(new_n22660_), .B0(pi0623), .Y(new_n22692_));
  AOI21X1  g20256(.A0(new_n22688_), .A1(new_n22660_), .B0(new_n22692_), .Y(new_n22693_));
  AOI21X1  g20257(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0207), .Y(new_n22694_));
  AOI21X1  g20258(.A0(new_n22694_), .A1(new_n22661_), .B0(new_n22693_), .Y(new_n22695_));
  NAND2X1  g20259(.A(new_n22695_), .B(new_n14326_), .Y(new_n22696_));
  INVX1    g20260(.A(pi0710), .Y(new_n22697_));
  NOR4X1   g20261(.A(new_n16582_), .B(new_n13508_), .C(new_n13489_), .D(new_n13433_), .Y(new_n22698_));
  INVX1    g20262(.A(new_n12737_), .Y(new_n22699_));
  OAI21X1  g20263(.A0(new_n16583_), .A1(new_n11770_), .B0(new_n11769_), .Y(new_n22700_));
  OAI21X1  g20264(.A0(new_n12832_), .A1(new_n11770_), .B0(new_n12363_), .Y(new_n22701_));
  OAI21X1  g20265(.A0(new_n16583_), .A1(new_n11770_), .B0(pi0625), .Y(new_n22702_));
  AOI21X1  g20266(.A0(new_n22702_), .A1(new_n22701_), .B0(new_n12364_), .Y(new_n22703_));
  OAI21X1  g20267(.A0(new_n12832_), .A1(new_n11770_), .B0(pi0625), .Y(new_n22704_));
  OAI21X1  g20268(.A0(new_n16583_), .A1(new_n11770_), .B0(new_n12363_), .Y(new_n22705_));
  AOI21X1  g20269(.A0(new_n22705_), .A1(new_n22704_), .B0(pi1153), .Y(new_n22706_));
  OAI21X1  g20270(.A0(new_n22706_), .A1(new_n22703_), .B0(pi0778), .Y(new_n22707_));
  NAND2X1  g20271(.A(new_n22707_), .B(new_n22700_), .Y(new_n22708_));
  MX2X1    g20272(.A(new_n22708_), .B(new_n22663_), .S0(new_n12490_), .Y(new_n22709_));
  MX2X1    g20273(.A(new_n22709_), .B(new_n22663_), .S0(new_n12513_), .Y(new_n22710_));
  INVX1    g20274(.A(new_n22710_), .Y(new_n22711_));
  MX2X1    g20275(.A(new_n22711_), .B(new_n22662_), .S0(new_n12531_), .Y(new_n22712_));
  AND3X1   g20276(.A(new_n12563_), .B(new_n12447_), .C(new_n3103_), .Y(new_n22713_));
  AOI21X1  g20277(.A0(new_n22712_), .A1(new_n13356_), .B0(new_n22713_), .Y(new_n22714_));
  OAI22X1  g20278(.A0(new_n22714_), .A1(new_n13508_), .B0(new_n22699_), .B1(new_n22663_), .Y(new_n22715_));
  INVX1    g20279(.A(new_n22715_), .Y(new_n22716_));
  MX2X1    g20280(.A(new_n22716_), .B(new_n22698_), .S0(pi0207), .Y(new_n22717_));
  MX2X1    g20281(.A(new_n22717_), .B(new_n22694_), .S0(new_n22697_), .Y(new_n22718_));
  INVX1    g20282(.A(new_n22718_), .Y(new_n22719_));
  AOI21X1  g20283(.A0(new_n22694_), .A1(pi0647), .B0(pi1157), .Y(new_n22720_));
  OAI21X1  g20284(.A0(new_n22719_), .A1(pi0647), .B0(new_n22720_), .Y(new_n22721_));
  AOI21X1  g20285(.A0(new_n22694_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n22722_));
  OAI21X1  g20286(.A0(new_n22719_), .A1(new_n12577_), .B0(new_n22722_), .Y(new_n22723_));
  MX2X1    g20287(.A(new_n22723_), .B(new_n22721_), .S0(pi0630), .Y(new_n22724_));
  AOI21X1  g20288(.A0(new_n22724_), .A1(new_n22696_), .B0(new_n11763_), .Y(new_n22725_));
  AOI21X1  g20289(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0628), .Y(new_n22726_));
  AOI21X1  g20290(.A0(new_n22714_), .A1(pi0628), .B0(new_n22726_), .Y(new_n22727_));
  OR2X1    g20291(.A(new_n22727_), .B(pi0629), .Y(new_n22728_));
  INVX1    g20292(.A(new_n22728_), .Y(new_n22729_));
  OAI21X1  g20293(.A0(new_n22729_), .A1(new_n22726_), .B0(pi1156), .Y(new_n22730_));
  AOI21X1  g20294(.A0(new_n12447_), .A1(new_n3103_), .B0(new_n12554_), .Y(new_n22731_));
  AOI21X1  g20295(.A0(new_n22714_), .A1(new_n12554_), .B0(new_n22731_), .Y(new_n22732_));
  INVX1    g20296(.A(new_n22732_), .Y(new_n22733_));
  AOI22X1  g20297(.A0(new_n22733_), .A1(new_n16374_), .B0(new_n22731_), .B1(new_n12555_), .Y(new_n22734_));
  AND2X1   g20298(.A(new_n22734_), .B(new_n22730_), .Y(new_n22735_));
  INVX1    g20299(.A(new_n22709_), .Y(new_n22736_));
  OAI21X1  g20300(.A0(new_n13543_), .A1(new_n11770_), .B0(new_n11769_), .Y(new_n22737_));
  NOR2X1   g20301(.A(new_n13543_), .B(new_n11770_), .Y(new_n22738_));
  MX2X1    g20302(.A(new_n22738_), .B(new_n22662_), .S0(pi0625), .Y(new_n22739_));
  NOR2X1   g20303(.A(new_n22703_), .B(pi0608), .Y(new_n22740_));
  OAI21X1  g20304(.A0(new_n22739_), .A1(pi1153), .B0(new_n22740_), .Y(new_n22741_));
  MX2X1    g20305(.A(new_n22738_), .B(new_n22662_), .S0(new_n12363_), .Y(new_n22742_));
  NOR2X1   g20306(.A(new_n22706_), .B(new_n12368_), .Y(new_n22743_));
  OAI21X1  g20307(.A0(new_n22742_), .A1(new_n12364_), .B0(new_n22743_), .Y(new_n22744_));
  NAND3X1  g20308(.A(new_n22744_), .B(new_n22741_), .C(pi0778), .Y(new_n22745_));
  AND2X1   g20309(.A(new_n22745_), .B(new_n22737_), .Y(new_n22746_));
  NAND2X1  g20310(.A(new_n22708_), .B(pi0609), .Y(new_n22747_));
  OAI21X1  g20311(.A0(new_n22746_), .A1(pi0609), .B0(new_n22747_), .Y(new_n22748_));
  OAI21X1  g20312(.A0(new_n22662_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n22749_));
  AOI21X1  g20313(.A0(new_n22748_), .A1(new_n12463_), .B0(new_n22749_), .Y(new_n22750_));
  NAND2X1  g20314(.A(new_n22708_), .B(new_n12462_), .Y(new_n22751_));
  OAI21X1  g20315(.A0(new_n22746_), .A1(new_n12462_), .B0(new_n22751_), .Y(new_n22752_));
  OAI21X1  g20316(.A0(new_n22662_), .A1(pi1155), .B0(pi0660), .Y(new_n22753_));
  AOI21X1  g20317(.A0(new_n22752_), .A1(pi1155), .B0(new_n22753_), .Y(new_n22754_));
  OR2X1    g20318(.A(new_n22754_), .B(new_n22750_), .Y(new_n22755_));
  MX2X1    g20319(.A(new_n22755_), .B(new_n22746_), .S0(new_n11768_), .Y(new_n22756_));
  MX2X1    g20320(.A(new_n22756_), .B(new_n22736_), .S0(pi0618), .Y(new_n22757_));
  AOI21X1  g20321(.A0(new_n22663_), .A1(pi1154), .B0(pi0627), .Y(new_n22758_));
  OAI21X1  g20322(.A0(new_n22757_), .A1(pi1154), .B0(new_n22758_), .Y(new_n22759_));
  MX2X1    g20323(.A(new_n22756_), .B(new_n22736_), .S0(new_n12486_), .Y(new_n22760_));
  AOI21X1  g20324(.A0(new_n22663_), .A1(new_n12487_), .B0(new_n12494_), .Y(new_n22761_));
  OAI21X1  g20325(.A0(new_n22760_), .A1(new_n12487_), .B0(new_n22761_), .Y(new_n22762_));
  AOI21X1  g20326(.A0(new_n22762_), .A1(new_n22759_), .B0(new_n11767_), .Y(new_n22763_));
  AND2X1   g20327(.A(new_n22756_), .B(new_n11767_), .Y(new_n22764_));
  NOR2X1   g20328(.A(new_n22764_), .B(new_n22763_), .Y(new_n22765_));
  AND2X1   g20329(.A(new_n22710_), .B(pi0619), .Y(new_n22766_));
  NOR3X1   g20330(.A(new_n22764_), .B(new_n22763_), .C(pi0619), .Y(new_n22767_));
  OAI21X1  g20331(.A0(new_n22767_), .A1(new_n22766_), .B0(new_n12510_), .Y(new_n22768_));
  AOI21X1  g20332(.A0(new_n22663_), .A1(pi1159), .B0(pi0648), .Y(new_n22769_));
  AND2X1   g20333(.A(new_n22710_), .B(new_n12509_), .Y(new_n22770_));
  NOR3X1   g20334(.A(new_n22764_), .B(new_n22763_), .C(new_n12509_), .Y(new_n22771_));
  OAI21X1  g20335(.A0(new_n22771_), .A1(new_n22770_), .B0(pi1159), .Y(new_n22772_));
  AOI21X1  g20336(.A0(new_n22663_), .A1(new_n12510_), .B0(new_n12517_), .Y(new_n22773_));
  AOI22X1  g20337(.A0(new_n22773_), .A1(new_n22772_), .B0(new_n22769_), .B1(new_n22768_), .Y(new_n22774_));
  MX2X1    g20338(.A(new_n22774_), .B(new_n22765_), .S0(new_n11766_), .Y(new_n22775_));
  AOI21X1  g20339(.A0(new_n22712_), .A1(pi0626), .B0(pi0641), .Y(new_n22776_));
  OAI21X1  g20340(.A0(new_n22775_), .A1(pi0626), .B0(new_n22776_), .Y(new_n22777_));
  AOI21X1  g20341(.A0(new_n22663_), .A1(pi0641), .B0(pi1158), .Y(new_n22778_));
  AOI21X1  g20342(.A0(new_n22712_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n22779_));
  OAI21X1  g20343(.A0(new_n22775_), .A1(new_n12542_), .B0(new_n22779_), .Y(new_n22780_));
  AOI21X1  g20344(.A0(new_n22663_), .A1(new_n12543_), .B0(new_n12548_), .Y(new_n22781_));
  AOI22X1  g20345(.A0(new_n22781_), .A1(new_n22780_), .B0(new_n22778_), .B1(new_n22777_), .Y(new_n22782_));
  NOR2X1   g20346(.A(new_n22782_), .B(new_n11765_), .Y(new_n22783_));
  OAI21X1  g20347(.A0(new_n22775_), .A1(pi0788), .B0(new_n14126_), .Y(new_n22784_));
  OAI22X1  g20348(.A0(new_n22784_), .A1(new_n22783_), .B0(new_n22735_), .B1(new_n11764_), .Y(new_n22785_));
  AND3X1   g20349(.A(new_n16664_), .B(new_n3103_), .C(new_n12363_), .Y(new_n22786_));
  OR4X1    g20350(.A(new_n16581_), .B(new_n12440_), .C(new_n11770_), .D(new_n12363_), .Y(new_n22787_));
  AOI21X1  g20351(.A0(new_n22787_), .A1(pi1153), .B0(pi0608), .Y(new_n22788_));
  OAI21X1  g20352(.A0(new_n22786_), .A1(pi1153), .B0(new_n22788_), .Y(new_n22789_));
  OAI21X1  g20353(.A0(new_n22150_), .A1(new_n12363_), .B0(pi1153), .Y(new_n22790_));
  OR4X1    g20354(.A(new_n16581_), .B(new_n12440_), .C(new_n11770_), .D(pi0625), .Y(new_n22791_));
  AOI21X1  g20355(.A0(new_n22791_), .A1(new_n12364_), .B0(new_n12368_), .Y(new_n22792_));
  AOI21X1  g20356(.A0(new_n22792_), .A1(new_n22790_), .B0(new_n11769_), .Y(new_n22793_));
  AOI22X1  g20357(.A0(new_n22793_), .A1(new_n22789_), .B0(new_n22150_), .B1(new_n11769_), .Y(new_n22794_));
  NOR2X1   g20358(.A(new_n22794_), .B(pi0609), .Y(new_n22795_));
  NOR4X1   g20359(.A(new_n16581_), .B(new_n13433_), .C(new_n12440_), .D(new_n11770_), .Y(new_n22796_));
  OAI21X1  g20360(.A0(new_n22796_), .A1(new_n12462_), .B0(new_n12489_), .Y(new_n22797_));
  NOR2X1   g20361(.A(new_n22794_), .B(new_n12462_), .Y(new_n22798_));
  OAI21X1  g20362(.A0(new_n22796_), .A1(pi0609), .B0(new_n12488_), .Y(new_n22799_));
  OAI22X1  g20363(.A0(new_n22799_), .A1(new_n22798_), .B0(new_n22797_), .B1(new_n22795_), .Y(new_n22800_));
  MX2X1    g20364(.A(new_n22800_), .B(new_n22794_), .S0(new_n11768_), .Y(new_n22801_));
  AOI21X1  g20365(.A0(new_n22796_), .A1(new_n13910_), .B0(new_n12486_), .Y(new_n22802_));
  NOR3X1   g20366(.A(new_n22802_), .B(pi1154), .C(pi0627), .Y(new_n22803_));
  OAI21X1  g20367(.A0(new_n22801_), .A1(pi0618), .B0(new_n22803_), .Y(new_n22804_));
  AOI21X1  g20368(.A0(new_n22796_), .A1(new_n13910_), .B0(pi0618), .Y(new_n22805_));
  NOR3X1   g20369(.A(new_n22805_), .B(new_n12487_), .C(new_n12494_), .Y(new_n22806_));
  OAI21X1  g20370(.A0(new_n22801_), .A1(new_n12486_), .B0(new_n22806_), .Y(new_n22807_));
  AND3X1   g20371(.A(new_n22807_), .B(new_n22804_), .C(pi0781), .Y(new_n22808_));
  OAI22X1  g20372(.A0(new_n22801_), .A1(pi0781), .B0(new_n16117_), .B1(new_n11766_), .Y(new_n22809_));
  NAND3X1  g20373(.A(new_n22796_), .B(new_n14053_), .C(new_n13910_), .Y(new_n22810_));
  NAND2X1  g20374(.A(new_n14036_), .B(new_n12530_), .Y(new_n22811_));
  OAI22X1  g20375(.A0(new_n22811_), .A1(new_n22810_), .B0(new_n22809_), .B1(new_n22808_), .Y(new_n22812_));
  NAND4X1  g20376(.A(new_n22796_), .B(new_n14051_), .C(new_n14053_), .D(new_n13910_), .Y(new_n22813_));
  AOI21X1  g20377(.A0(new_n22813_), .A1(pi0626), .B0(pi0641), .Y(new_n22814_));
  AND2X1   g20378(.A(new_n22814_), .B(new_n12548_), .Y(new_n22815_));
  OAI21X1  g20379(.A0(new_n22812_), .A1(pi0626), .B0(new_n22815_), .Y(new_n22816_));
  AOI21X1  g20380(.A0(new_n22813_), .A1(new_n12542_), .B0(new_n12543_), .Y(new_n22817_));
  AND2X1   g20381(.A(new_n22817_), .B(pi1158), .Y(new_n22818_));
  OAI21X1  g20382(.A0(new_n22812_), .A1(new_n12542_), .B0(new_n22818_), .Y(new_n22819_));
  AND3X1   g20383(.A(new_n22819_), .B(new_n22816_), .C(pi0788), .Y(new_n22820_));
  OAI21X1  g20384(.A0(new_n22812_), .A1(pi0788), .B0(new_n14126_), .Y(new_n22821_));
  OR2X1    g20385(.A(new_n22821_), .B(new_n22820_), .Y(new_n22822_));
  NOR3X1   g20386(.A(new_n16582_), .B(new_n13489_), .C(new_n13433_), .Y(new_n22823_));
  NAND4X1  g20387(.A(new_n22823_), .B(new_n12736_), .C(new_n12734_), .D(new_n12580_), .Y(new_n22824_));
  AND2X1   g20388(.A(new_n22824_), .B(new_n22822_), .Y(new_n22825_));
  OAI21X1  g20389(.A0(new_n22825_), .A1(new_n22660_), .B0(new_n22661_), .Y(new_n22826_));
  AOI21X1  g20390(.A0(new_n22785_), .A1(new_n22660_), .B0(new_n22826_), .Y(new_n22827_));
  OR4X1    g20391(.A(new_n13558_), .B(new_n13557_), .C(new_n13555_), .D(new_n11770_), .Y(new_n22828_));
  OAI21X1  g20392(.A0(new_n22828_), .A1(new_n12363_), .B0(pi1153), .Y(new_n22829_));
  AOI21X1  g20393(.A0(new_n22664_), .A1(new_n12363_), .B0(new_n22829_), .Y(new_n22830_));
  OR3X1    g20394(.A(new_n22830_), .B(new_n22706_), .C(new_n12368_), .Y(new_n22831_));
  OAI21X1  g20395(.A0(new_n22828_), .A1(pi0625), .B0(new_n12364_), .Y(new_n22832_));
  AOI21X1  g20396(.A0(new_n22664_), .A1(pi0625), .B0(new_n22832_), .Y(new_n22833_));
  OR3X1    g20397(.A(new_n22833_), .B(new_n22703_), .C(pi0608), .Y(new_n22834_));
  AND3X1   g20398(.A(new_n22834_), .B(new_n22831_), .C(pi0778), .Y(new_n22835_));
  AOI21X1  g20399(.A0(new_n22828_), .A1(new_n11769_), .B0(new_n22835_), .Y(new_n22836_));
  OAI21X1  g20400(.A0(new_n22836_), .A1(pi0609), .B0(new_n22747_), .Y(new_n22837_));
  OAI21X1  g20401(.A0(new_n22668_), .A1(new_n12463_), .B0(new_n12468_), .Y(new_n22838_));
  AOI21X1  g20402(.A0(new_n22837_), .A1(new_n12463_), .B0(new_n22838_), .Y(new_n22839_));
  OAI21X1  g20403(.A0(new_n22836_), .A1(new_n12462_), .B0(new_n22751_), .Y(new_n22840_));
  OAI21X1  g20404(.A0(new_n22667_), .A1(pi1155), .B0(pi0660), .Y(new_n22841_));
  AOI21X1  g20405(.A0(new_n22840_), .A1(pi1155), .B0(new_n22841_), .Y(new_n22842_));
  OR2X1    g20406(.A(new_n22842_), .B(new_n22839_), .Y(new_n22843_));
  MX2X1    g20407(.A(new_n22843_), .B(new_n22836_), .S0(new_n11768_), .Y(new_n22844_));
  MX2X1    g20408(.A(new_n22844_), .B(new_n22736_), .S0(pi0618), .Y(new_n22845_));
  NOR2X1   g20409(.A(new_n22675_), .B(pi0627), .Y(new_n22846_));
  OAI21X1  g20410(.A0(new_n22845_), .A1(pi1154), .B0(new_n22846_), .Y(new_n22847_));
  MX2X1    g20411(.A(new_n22844_), .B(new_n22736_), .S0(new_n12486_), .Y(new_n22848_));
  NOR2X1   g20412(.A(new_n22673_), .B(new_n12494_), .Y(new_n22849_));
  OAI21X1  g20413(.A0(new_n22848_), .A1(new_n12487_), .B0(new_n22849_), .Y(new_n22850_));
  AOI21X1  g20414(.A0(new_n22850_), .A1(new_n22847_), .B0(new_n11767_), .Y(new_n22851_));
  AND2X1   g20415(.A(new_n22844_), .B(new_n11767_), .Y(new_n22852_));
  NOR3X1   g20416(.A(new_n22852_), .B(new_n22851_), .C(pi0619), .Y(new_n22853_));
  OAI21X1  g20417(.A0(new_n22853_), .A1(new_n22766_), .B0(new_n12510_), .Y(new_n22854_));
  AND3X1   g20418(.A(new_n22854_), .B(new_n22682_), .C(new_n12517_), .Y(new_n22855_));
  INVX1    g20419(.A(new_n22770_), .Y(new_n22856_));
  OR3X1    g20420(.A(new_n22852_), .B(new_n22851_), .C(new_n12509_), .Y(new_n22857_));
  AOI21X1  g20421(.A0(new_n22857_), .A1(new_n22856_), .B0(new_n12510_), .Y(new_n22858_));
  AND2X1   g20422(.A(new_n22680_), .B(pi0648), .Y(new_n22859_));
  INVX1    g20423(.A(new_n22859_), .Y(new_n22860_));
  OAI21X1  g20424(.A0(new_n22860_), .A1(new_n22858_), .B0(pi0789), .Y(new_n22861_));
  NOR3X1   g20425(.A(new_n22852_), .B(new_n22851_), .C(pi0789), .Y(new_n22862_));
  NOR2X1   g20426(.A(new_n22862_), .B(new_n13481_), .Y(new_n22863_));
  OAI21X1  g20427(.A0(new_n22861_), .A1(new_n22855_), .B0(new_n22863_), .Y(new_n22864_));
  AND2X1   g20428(.A(new_n12636_), .B(new_n12639_), .Y(new_n22865_));
  NAND2X1  g20429(.A(new_n22865_), .B(new_n22684_), .Y(new_n22866_));
  AOI21X1  g20430(.A0(new_n22663_), .A1(new_n12543_), .B0(new_n14050_), .Y(new_n22867_));
  OAI21X1  g20431(.A0(new_n22712_), .A1(new_n12543_), .B0(new_n22867_), .Y(new_n22868_));
  AOI21X1  g20432(.A0(new_n22663_), .A1(pi0641), .B0(new_n14062_), .Y(new_n22869_));
  OAI21X1  g20433(.A0(new_n22712_), .A1(pi0641), .B0(new_n22869_), .Y(new_n22870_));
  AND3X1   g20434(.A(new_n22870_), .B(new_n22868_), .C(new_n22866_), .Y(new_n22871_));
  OAI21X1  g20435(.A0(new_n22871_), .A1(new_n11765_), .B0(new_n14126_), .Y(new_n22872_));
  INVX1    g20436(.A(new_n22872_), .Y(new_n22873_));
  NAND2X1  g20437(.A(new_n22686_), .B(new_n14249_), .Y(new_n22874_));
  AOI22X1  g20438(.A0(new_n22733_), .A1(new_n16374_), .B0(new_n22729_), .B1(pi1156), .Y(new_n22875_));
  AOI21X1  g20439(.A0(new_n22875_), .A1(new_n22874_), .B0(new_n11764_), .Y(new_n22876_));
  AOI21X1  g20440(.A0(new_n22873_), .A1(new_n22864_), .B0(new_n22876_), .Y(new_n22877_));
  OR3X1    g20441(.A(new_n22690_), .B(new_n14036_), .C(new_n12708_), .Y(new_n22878_));
  OAI21X1  g20442(.A0(new_n22823_), .A1(pi1156), .B0(new_n14247_), .Y(new_n22879_));
  AOI21X1  g20443(.A0(new_n22878_), .A1(pi1156), .B0(new_n22879_), .Y(new_n22880_));
  OAI21X1  g20444(.A0(new_n22823_), .A1(new_n12555_), .B0(new_n14248_), .Y(new_n22881_));
  AOI21X1  g20445(.A0(new_n22878_), .A1(new_n12555_), .B0(new_n22881_), .Y(new_n22882_));
  OAI21X1  g20446(.A0(new_n22882_), .A1(new_n22880_), .B0(pi0792), .Y(new_n22883_));
  AND2X1   g20447(.A(new_n22690_), .B(new_n12510_), .Y(new_n22884_));
  AND2X1   g20448(.A(new_n22810_), .B(pi1159), .Y(new_n22885_));
  NOR4X1   g20449(.A(new_n22885_), .B(new_n22884_), .C(new_n12517_), .D(pi0619), .Y(new_n22886_));
  AND2X1   g20450(.A(new_n22690_), .B(pi1159), .Y(new_n22887_));
  AND2X1   g20451(.A(new_n22810_), .B(new_n12510_), .Y(new_n22888_));
  NOR4X1   g20452(.A(new_n22888_), .B(new_n22887_), .C(pi0648), .D(new_n12509_), .Y(new_n22889_));
  OAI21X1  g20453(.A0(new_n22889_), .A1(new_n22886_), .B0(pi0789), .Y(new_n22890_));
  OR2X1    g20454(.A(new_n22802_), .B(pi1154), .Y(new_n22891_));
  NOR3X1   g20455(.A(new_n22689_), .B(new_n14034_), .C(new_n12473_), .Y(new_n22892_));
  AOI21X1  g20456(.A0(new_n22892_), .A1(new_n14038_), .B0(pi0627), .Y(new_n22893_));
  AOI21X1  g20457(.A0(new_n13554_), .A1(new_n3103_), .B0(pi0778), .Y(new_n22894_));
  AND3X1   g20458(.A(new_n13554_), .B(new_n3103_), .C(new_n12363_), .Y(new_n22895_));
  OAI21X1  g20459(.A0(new_n22689_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n22896_));
  OAI21X1  g20460(.A0(new_n22896_), .A1(new_n22895_), .B0(new_n22788_), .Y(new_n22897_));
  AND3X1   g20461(.A(new_n13554_), .B(new_n3103_), .C(pi0625), .Y(new_n22898_));
  OAI21X1  g20462(.A0(new_n22689_), .A1(pi0625), .B0(pi1153), .Y(new_n22899_));
  OAI21X1  g20463(.A0(new_n22899_), .A1(new_n22898_), .B0(new_n22792_), .Y(new_n22900_));
  AND3X1   g20464(.A(new_n22900_), .B(new_n22897_), .C(pi0778), .Y(new_n22901_));
  NOR2X1   g20465(.A(new_n22901_), .B(new_n22894_), .Y(new_n22902_));
  INVX1    g20466(.A(new_n22796_), .Y(new_n22903_));
  AOI21X1  g20467(.A0(new_n22903_), .A1(pi0609), .B0(pi1155), .Y(new_n22904_));
  OAI21X1  g20468(.A0(new_n22902_), .A1(pi0609), .B0(new_n22904_), .Y(new_n22905_));
  NAND4X1  g20469(.A(new_n16617_), .B(new_n14033_), .C(new_n12474_), .D(new_n3103_), .Y(new_n22906_));
  AND2X1   g20470(.A(new_n22906_), .B(new_n12468_), .Y(new_n22907_));
  AOI21X1  g20471(.A0(new_n22903_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n22908_));
  OAI21X1  g20472(.A0(new_n22902_), .A1(new_n12462_), .B0(new_n22908_), .Y(new_n22909_));
  NAND4X1  g20473(.A(new_n16617_), .B(new_n14032_), .C(new_n12474_), .D(new_n3103_), .Y(new_n22910_));
  AND2X1   g20474(.A(new_n22910_), .B(pi0660), .Y(new_n22911_));
  AOI22X1  g20475(.A0(new_n22911_), .A1(new_n22909_), .B0(new_n22907_), .B1(new_n22905_), .Y(new_n22912_));
  MX2X1    g20476(.A(new_n22912_), .B(new_n22902_), .S0(new_n11768_), .Y(new_n22913_));
  NOR2X1   g20477(.A(new_n22805_), .B(new_n12487_), .Y(new_n22914_));
  OAI21X1  g20478(.A0(new_n22913_), .A1(new_n12486_), .B0(new_n22914_), .Y(new_n22915_));
  AOI21X1  g20479(.A0(new_n22892_), .A1(new_n14037_), .B0(new_n12494_), .Y(new_n22916_));
  AOI22X1  g20480(.A0(new_n22916_), .A1(new_n22915_), .B0(new_n22893_), .B1(new_n22891_), .Y(new_n22917_));
  NOR2X1   g20481(.A(new_n22917_), .B(new_n11767_), .Y(new_n22918_));
  AOI21X1  g20482(.A0(new_n12494_), .A1(new_n12486_), .B0(new_n11767_), .Y(new_n22919_));
  OR4X1    g20483(.A(new_n22889_), .B(new_n22886_), .C(new_n16117_), .D(new_n11766_), .Y(new_n22920_));
  OAI21X1  g20484(.A0(new_n22919_), .A1(new_n22913_), .B0(new_n22920_), .Y(new_n22921_));
  OAI21X1  g20485(.A0(new_n22921_), .A1(new_n22918_), .B0(new_n22890_), .Y(new_n22922_));
  OAI21X1  g20486(.A0(new_n22922_), .A1(pi0626), .B0(new_n22814_), .Y(new_n22923_));
  OR4X1    g20487(.A(new_n22690_), .B(new_n14036_), .C(new_n12543_), .D(pi0626), .Y(new_n22924_));
  AND2X1   g20488(.A(new_n22924_), .B(new_n12548_), .Y(new_n22925_));
  OAI21X1  g20489(.A0(new_n22922_), .A1(new_n12542_), .B0(new_n22817_), .Y(new_n22926_));
  OR4X1    g20490(.A(new_n22690_), .B(new_n14036_), .C(pi0641), .D(new_n12542_), .Y(new_n22927_));
  AND2X1   g20491(.A(new_n22927_), .B(pi1158), .Y(new_n22928_));
  AOI22X1  g20492(.A0(new_n22928_), .A1(new_n22926_), .B0(new_n22925_), .B1(new_n22923_), .Y(new_n22929_));
  OR2X1    g20493(.A(new_n22922_), .B(pi0788), .Y(new_n22930_));
  AND2X1   g20494(.A(new_n22930_), .B(new_n14126_), .Y(new_n22931_));
  OAI21X1  g20495(.A0(new_n22929_), .A1(new_n11765_), .B0(new_n22931_), .Y(new_n22932_));
  AND2X1   g20496(.A(new_n22932_), .B(new_n22883_), .Y(new_n22933_));
  INVX1    g20497(.A(new_n22933_), .Y(new_n22934_));
  AOI21X1  g20498(.A0(new_n22934_), .A1(pi0207), .B0(new_n22661_), .Y(new_n22935_));
  OAI21X1  g20499(.A0(new_n22877_), .A1(pi0207), .B0(new_n22935_), .Y(new_n22936_));
  NAND2X1  g20500(.A(new_n22936_), .B(pi0710), .Y(new_n22937_));
  OR2X1    g20501(.A(new_n22937_), .B(new_n22827_), .Y(new_n22938_));
  INVX1    g20502(.A(new_n22695_), .Y(new_n22939_));
  AOI21X1  g20503(.A0(new_n22939_), .A1(new_n22697_), .B0(new_n14121_), .Y(new_n22940_));
  AOI21X1  g20504(.A0(new_n22940_), .A1(new_n22938_), .B0(new_n22725_), .Y(new_n22941_));
  NAND2X1  g20505(.A(new_n22723_), .B(new_n22721_), .Y(new_n22942_));
  MX2X1    g20506(.A(new_n22942_), .B(new_n22719_), .S0(new_n11763_), .Y(new_n22943_));
  OAI21X1  g20507(.A0(new_n22943_), .A1(pi0644), .B0(pi0715), .Y(new_n22944_));
  AOI21X1  g20508(.A0(new_n22941_), .A1(pi0644), .B0(new_n22944_), .Y(new_n22945_));
  MX2X1    g20509(.A(new_n22939_), .B(new_n22694_), .S0(new_n12604_), .Y(new_n22946_));
  INVX1    g20510(.A(new_n22694_), .Y(new_n22947_));
  OAI21X1  g20511(.A0(new_n22947_), .A1(pi0644), .B0(new_n12608_), .Y(new_n22948_));
  AOI21X1  g20512(.A0(new_n22946_), .A1(pi0644), .B0(new_n22948_), .Y(new_n22949_));
  OR2X1    g20513(.A(new_n22949_), .B(new_n11762_), .Y(new_n22950_));
  OAI21X1  g20514(.A0(new_n22943_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n22951_));
  AOI21X1  g20515(.A0(new_n22941_), .A1(new_n12612_), .B0(new_n22951_), .Y(new_n22952_));
  OAI21X1  g20516(.A0(new_n22947_), .A1(new_n12612_), .B0(pi0715), .Y(new_n22953_));
  AOI21X1  g20517(.A0(new_n22946_), .A1(new_n12612_), .B0(new_n22953_), .Y(new_n22954_));
  OR2X1    g20518(.A(new_n22954_), .B(pi1160), .Y(new_n22955_));
  OAI22X1  g20519(.A0(new_n22955_), .A1(new_n22952_), .B0(new_n22950_), .B1(new_n22945_), .Y(new_n22956_));
  MX2X1    g20520(.A(new_n22956_), .B(new_n22941_), .S0(new_n12766_), .Y(new_n22957_));
  MX2X1    g20521(.A(new_n22957_), .B(new_n22660_), .S0(po1038), .Y(po0364));
  INVX1    g20522(.A(pi0208), .Y(new_n22959_));
  INVX1    g20523(.A(pi0607), .Y(new_n22960_));
  OAI21X1  g20524(.A0(new_n22691_), .A1(new_n22959_), .B0(pi0607), .Y(new_n22961_));
  AOI21X1  g20525(.A0(new_n22688_), .A1(new_n22959_), .B0(new_n22961_), .Y(new_n22962_));
  AOI21X1  g20526(.A0(new_n12447_), .A1(new_n3103_), .B0(pi0208), .Y(new_n22963_));
  AOI21X1  g20527(.A0(new_n22963_), .A1(new_n22960_), .B0(new_n22962_), .Y(new_n22964_));
  NAND2X1  g20528(.A(new_n22964_), .B(new_n14326_), .Y(new_n22965_));
  INVX1    g20529(.A(pi0638), .Y(new_n22966_));
  MX2X1    g20530(.A(new_n22716_), .B(new_n22698_), .S0(pi0208), .Y(new_n22967_));
  MX2X1    g20531(.A(new_n22967_), .B(new_n22963_), .S0(new_n22966_), .Y(new_n22968_));
  INVX1    g20532(.A(new_n22968_), .Y(new_n22969_));
  AOI21X1  g20533(.A0(new_n22963_), .A1(pi0647), .B0(pi1157), .Y(new_n22970_));
  OAI21X1  g20534(.A0(new_n22969_), .A1(pi0647), .B0(new_n22970_), .Y(new_n22971_));
  AOI21X1  g20535(.A0(new_n22963_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n22972_));
  OAI21X1  g20536(.A0(new_n22969_), .A1(new_n12577_), .B0(new_n22972_), .Y(new_n22973_));
  MX2X1    g20537(.A(new_n22973_), .B(new_n22971_), .S0(pi0630), .Y(new_n22974_));
  AOI21X1  g20538(.A0(new_n22974_), .A1(new_n22965_), .B0(new_n11763_), .Y(new_n22975_));
  OAI21X1  g20539(.A0(new_n22825_), .A1(new_n22959_), .B0(new_n22960_), .Y(new_n22976_));
  AOI21X1  g20540(.A0(new_n22785_), .A1(new_n22959_), .B0(new_n22976_), .Y(new_n22977_));
  AOI21X1  g20541(.A0(new_n22934_), .A1(pi0208), .B0(new_n22960_), .Y(new_n22978_));
  OAI21X1  g20542(.A0(new_n22877_), .A1(pi0208), .B0(new_n22978_), .Y(new_n22979_));
  NAND2X1  g20543(.A(new_n22979_), .B(pi0638), .Y(new_n22980_));
  OR2X1    g20544(.A(new_n22980_), .B(new_n22977_), .Y(new_n22981_));
  INVX1    g20545(.A(new_n22964_), .Y(new_n22982_));
  AOI21X1  g20546(.A0(new_n22982_), .A1(new_n22966_), .B0(new_n14121_), .Y(new_n22983_));
  AOI21X1  g20547(.A0(new_n22983_), .A1(new_n22981_), .B0(new_n22975_), .Y(new_n22984_));
  NAND2X1  g20548(.A(new_n22973_), .B(new_n22971_), .Y(new_n22985_));
  MX2X1    g20549(.A(new_n22985_), .B(new_n22969_), .S0(new_n11763_), .Y(new_n22986_));
  OAI21X1  g20550(.A0(new_n22986_), .A1(pi0644), .B0(pi0715), .Y(new_n22987_));
  AOI21X1  g20551(.A0(new_n22984_), .A1(pi0644), .B0(new_n22987_), .Y(new_n22988_));
  MX2X1    g20552(.A(new_n22982_), .B(new_n22963_), .S0(new_n12604_), .Y(new_n22989_));
  INVX1    g20553(.A(new_n22963_), .Y(new_n22990_));
  OAI21X1  g20554(.A0(new_n22990_), .A1(pi0644), .B0(new_n12608_), .Y(new_n22991_));
  AOI21X1  g20555(.A0(new_n22989_), .A1(pi0644), .B0(new_n22991_), .Y(new_n22992_));
  OR2X1    g20556(.A(new_n22992_), .B(new_n11762_), .Y(new_n22993_));
  OAI21X1  g20557(.A0(new_n22986_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n22994_));
  AOI21X1  g20558(.A0(new_n22984_), .A1(new_n12612_), .B0(new_n22994_), .Y(new_n22995_));
  OAI21X1  g20559(.A0(new_n22990_), .A1(new_n12612_), .B0(pi0715), .Y(new_n22996_));
  AOI21X1  g20560(.A0(new_n22989_), .A1(new_n12612_), .B0(new_n22996_), .Y(new_n22997_));
  OR2X1    g20561(.A(new_n22997_), .B(pi1160), .Y(new_n22998_));
  OAI22X1  g20562(.A0(new_n22998_), .A1(new_n22995_), .B0(new_n22993_), .B1(new_n22988_), .Y(new_n22999_));
  MX2X1    g20563(.A(new_n22999_), .B(new_n22984_), .S0(new_n12766_), .Y(new_n23000_));
  MX2X1    g20564(.A(new_n23000_), .B(new_n22959_), .S0(po1038), .Y(po0365));
  INVX1    g20565(.A(pi0639), .Y(new_n23002_));
  MX2X1    g20566(.A(new_n22715_), .B(new_n22662_), .S0(new_n12577_), .Y(new_n23003_));
  OAI22X1  g20567(.A0(new_n23003_), .A1(pi0630), .B0(new_n22662_), .B1(pi0647), .Y(new_n23004_));
  NAND2X1  g20568(.A(new_n23004_), .B(pi1157), .Y(new_n23005_));
  AOI21X1  g20569(.A0(new_n12447_), .A1(new_n3103_), .B0(new_n12577_), .Y(new_n23006_));
  MX2X1    g20570(.A(new_n22715_), .B(new_n22662_), .S0(pi0647), .Y(new_n23007_));
  INVX1    g20571(.A(new_n23007_), .Y(new_n23008_));
  AOI22X1  g20572(.A0(new_n23008_), .A1(new_n14243_), .B0(new_n23006_), .B1(new_n12578_), .Y(new_n23009_));
  AOI21X1  g20573(.A0(new_n23009_), .A1(new_n23005_), .B0(new_n11763_), .Y(new_n23010_));
  AOI21X1  g20574(.A0(new_n22785_), .A1(new_n14122_), .B0(new_n23010_), .Y(new_n23011_));
  MX2X1    g20575(.A(new_n22715_), .B(new_n22662_), .S0(new_n13520_), .Y(new_n23012_));
  INVX1    g20576(.A(new_n23012_), .Y(new_n23013_));
  AOI21X1  g20577(.A0(new_n23013_), .A1(pi0644), .B0(pi0715), .Y(new_n23014_));
  OAI21X1  g20578(.A0(new_n23011_), .A1(pi0644), .B0(new_n23014_), .Y(new_n23015_));
  AOI21X1  g20579(.A0(new_n22662_), .A1(pi0715), .B0(pi1160), .Y(new_n23016_));
  AOI21X1  g20580(.A0(new_n23013_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n23017_));
  OAI21X1  g20581(.A0(new_n23011_), .A1(new_n12612_), .B0(new_n23017_), .Y(new_n23018_));
  AOI21X1  g20582(.A0(new_n22662_), .A1(new_n12608_), .B0(new_n11762_), .Y(new_n23019_));
  AOI22X1  g20583(.A0(new_n23019_), .A1(new_n23018_), .B0(new_n23016_), .B1(new_n23015_), .Y(new_n23020_));
  NOR2X1   g20584(.A(new_n23020_), .B(new_n12766_), .Y(new_n23021_));
  OAI21X1  g20585(.A0(new_n23011_), .A1(pi0790), .B0(new_n6489_), .Y(new_n23022_));
  OR3X1    g20586(.A(new_n23022_), .B(new_n23021_), .C(new_n23002_), .Y(new_n23023_));
  AND2X1   g20587(.A(new_n12447_), .B(new_n7625_), .Y(new_n23024_));
  AOI21X1  g20588(.A0(new_n23024_), .A1(new_n23002_), .B0(pi0622), .Y(new_n23025_));
  INVX1    g20589(.A(new_n23014_), .Y(new_n23026_));
  NOR3X1   g20590(.A(new_n23003_), .B(new_n12578_), .C(pi0630), .Y(new_n23027_));
  AOI21X1  g20591(.A0(new_n23008_), .A1(new_n14243_), .B0(new_n23027_), .Y(new_n23028_));
  OAI21X1  g20592(.A0(new_n22688_), .A1(new_n14239_), .B0(new_n23028_), .Y(new_n23029_));
  NAND2X1  g20593(.A(new_n23029_), .B(pi0787), .Y(new_n23030_));
  OAI21X1  g20594(.A0(new_n22877_), .A1(new_n14121_), .B0(new_n23030_), .Y(new_n23031_));
  AOI21X1  g20595(.A0(new_n23031_), .A1(new_n12612_), .B0(new_n23026_), .Y(new_n23032_));
  MX2X1    g20596(.A(new_n22688_), .B(new_n22662_), .S0(new_n12604_), .Y(new_n23033_));
  MX2X1    g20597(.A(new_n23033_), .B(new_n22662_), .S0(pi0644), .Y(new_n23034_));
  AOI21X1  g20598(.A0(new_n23034_), .A1(pi0715), .B0(pi1160), .Y(new_n23035_));
  INVX1    g20599(.A(new_n23035_), .Y(new_n23036_));
  INVX1    g20600(.A(new_n23017_), .Y(new_n23037_));
  AOI21X1  g20601(.A0(new_n23031_), .A1(pi0644), .B0(new_n23037_), .Y(new_n23038_));
  MX2X1    g20602(.A(new_n23033_), .B(new_n22662_), .S0(new_n12612_), .Y(new_n23039_));
  AOI21X1  g20603(.A0(new_n23039_), .A1(new_n12608_), .B0(new_n11762_), .Y(new_n23040_));
  INVX1    g20604(.A(new_n23040_), .Y(new_n23041_));
  OAI22X1  g20605(.A0(new_n23041_), .A1(new_n23038_), .B0(new_n23036_), .B1(new_n23032_), .Y(new_n23042_));
  AOI21X1  g20606(.A0(new_n23031_), .A1(new_n12766_), .B0(po1038), .Y(new_n23043_));
  INVX1    g20607(.A(new_n23043_), .Y(new_n23044_));
  AOI21X1  g20608(.A0(new_n23042_), .A1(pi0790), .B0(new_n23044_), .Y(new_n23045_));
  NAND2X1  g20609(.A(new_n23045_), .B(pi0639), .Y(new_n23046_));
  INVX1    g20610(.A(pi0622), .Y(new_n23047_));
  AND2X1   g20611(.A(new_n23039_), .B(pi1160), .Y(new_n23048_));
  INVX1    g20612(.A(new_n23048_), .Y(new_n23049_));
  AOI21X1  g20613(.A0(new_n23034_), .A1(new_n11762_), .B0(new_n12766_), .Y(new_n23050_));
  OAI21X1  g20614(.A0(new_n23033_), .A1(pi0790), .B0(new_n6489_), .Y(new_n23051_));
  AOI21X1  g20615(.A0(new_n23050_), .A1(new_n23049_), .B0(new_n23051_), .Y(new_n23052_));
  AOI21X1  g20616(.A0(new_n23052_), .A1(new_n23002_), .B0(new_n23047_), .Y(new_n23053_));
  AOI22X1  g20617(.A0(new_n23053_), .A1(new_n23046_), .B0(new_n23025_), .B1(new_n23023_), .Y(new_n23054_));
  AND2X1   g20618(.A(new_n22698_), .B(new_n14140_), .Y(new_n23055_));
  OAI21X1  g20619(.A0(new_n23055_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n23056_));
  AOI21X1  g20620(.A0(new_n22691_), .A1(pi0647), .B0(pi1157), .Y(new_n23057_));
  OAI21X1  g20621(.A0(new_n22933_), .A1(pi0647), .B0(new_n23057_), .Y(new_n23058_));
  AOI21X1  g20622(.A0(new_n22698_), .A1(pi0647), .B0(new_n12578_), .Y(new_n23059_));
  OR2X1    g20623(.A(new_n23059_), .B(pi0630), .Y(new_n23060_));
  INVX1    g20624(.A(new_n23060_), .Y(new_n23061_));
  AOI21X1  g20625(.A0(new_n22691_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n23062_));
  OAI21X1  g20626(.A0(new_n22933_), .A1(new_n12577_), .B0(new_n23062_), .Y(new_n23063_));
  AOI21X1  g20627(.A0(new_n22698_), .A1(new_n12577_), .B0(pi1157), .Y(new_n23064_));
  OR2X1    g20628(.A(new_n23064_), .B(new_n12592_), .Y(new_n23065_));
  INVX1    g20629(.A(new_n23065_), .Y(new_n23066_));
  AOI22X1  g20630(.A0(new_n23066_), .A1(new_n23063_), .B0(new_n23061_), .B1(new_n23058_), .Y(new_n23067_));
  MX2X1    g20631(.A(new_n23067_), .B(new_n22933_), .S0(new_n11763_), .Y(new_n23068_));
  AOI21X1  g20632(.A0(new_n23068_), .A1(new_n12612_), .B0(new_n23056_), .Y(new_n23069_));
  OR4X1    g20633(.A(new_n22690_), .B(new_n16164_), .C(new_n14036_), .D(new_n12708_), .Y(new_n23070_));
  OR2X1    g20634(.A(new_n12608_), .B(pi0644), .Y(new_n23071_));
  OAI21X1  g20635(.A0(new_n23071_), .A1(new_n23070_), .B0(new_n11762_), .Y(new_n23072_));
  OAI21X1  g20636(.A0(new_n23055_), .A1(pi0644), .B0(pi0715), .Y(new_n23073_));
  AOI21X1  g20637(.A0(new_n23068_), .A1(pi0644), .B0(new_n23073_), .Y(new_n23074_));
  OR2X1    g20638(.A(pi0715), .B(new_n12612_), .Y(new_n23075_));
  OAI21X1  g20639(.A0(new_n23075_), .A1(new_n23070_), .B0(pi1160), .Y(new_n23076_));
  OAI22X1  g20640(.A0(new_n23076_), .A1(new_n23074_), .B0(new_n23072_), .B1(new_n23069_), .Y(new_n23077_));
  AND2X1   g20641(.A(new_n23068_), .B(new_n12766_), .Y(new_n23078_));
  OR2X1    g20642(.A(new_n23078_), .B(po1038), .Y(new_n23079_));
  AOI21X1  g20643(.A0(new_n23077_), .A1(pi0790), .B0(new_n23079_), .Y(new_n23080_));
  NAND2X1  g20644(.A(pi0639), .B(pi0622), .Y(new_n23081_));
  AOI21X1  g20645(.A0(new_n22824_), .A1(new_n22822_), .B0(new_n14121_), .Y(new_n23082_));
  AND2X1   g20646(.A(new_n13519_), .B(new_n12604_), .Y(new_n23083_));
  AOI21X1  g20647(.A0(new_n23083_), .A1(new_n22698_), .B0(new_n23082_), .Y(new_n23084_));
  OR2X1    g20648(.A(new_n23073_), .B(new_n11762_), .Y(new_n23085_));
  AOI21X1  g20649(.A0(new_n23084_), .A1(pi0644), .B0(new_n23085_), .Y(new_n23086_));
  OR2X1    g20650(.A(new_n23056_), .B(pi1160), .Y(new_n23087_));
  AOI21X1  g20651(.A0(new_n23084_), .A1(new_n12612_), .B0(new_n23087_), .Y(new_n23088_));
  OR3X1    g20652(.A(new_n23088_), .B(new_n23086_), .C(new_n12766_), .Y(new_n23089_));
  AOI21X1  g20653(.A0(new_n23084_), .A1(new_n12766_), .B0(po1038), .Y(new_n23090_));
  AOI21X1  g20654(.A0(new_n23090_), .A1(new_n23089_), .B0(pi0622), .Y(new_n23091_));
  XOR2X1   g20655(.A(pi1160), .B(pi0644), .Y(new_n23092_));
  AND2X1   g20656(.A(new_n23092_), .B(pi0790), .Y(new_n23093_));
  NOR4X1   g20657(.A(new_n23093_), .B(new_n23070_), .C(po1038), .D(new_n23047_), .Y(new_n23094_));
  OAI21X1  g20658(.A0(new_n23094_), .A1(pi0639), .B0(pi0209), .Y(new_n23095_));
  NOR2X1   g20659(.A(new_n23095_), .B(new_n23091_), .Y(new_n23096_));
  OAI21X1  g20660(.A0(new_n23081_), .A1(new_n23080_), .B0(new_n23096_), .Y(new_n23097_));
  OAI21X1  g20661(.A0(new_n23054_), .A1(pi0209), .B0(new_n23097_), .Y(po0366));
  AOI22X1  g20662(.A0(new_n14453_), .A1(pi0634), .B0(pi0947), .B1(pi0633), .Y(new_n23099_));
  OAI21X1  g20663(.A0(new_n23099_), .A1(new_n12771_), .B0(pi0038), .Y(new_n23100_));
  AOI21X1  g20664(.A0(new_n12771_), .A1(pi0210), .B0(new_n23100_), .Y(new_n23101_));
  AND2X1   g20665(.A(new_n11825_), .B(pi0210), .Y(new_n23102_));
  NOR2X1   g20666(.A(new_n5021_), .B(new_n2777_), .Y(new_n23103_));
  AOI22X1  g20667(.A0(new_n23103_), .A1(new_n11917_), .B0(new_n23102_), .B1(new_n5021_), .Y(new_n23104_));
  NAND2X1  g20668(.A(new_n23104_), .B(new_n5277_), .Y(new_n23105_));
  MX2X1    g20669(.A(new_n21904_), .B(new_n2777_), .S0(new_n11825_), .Y(new_n23106_));
  OR2X1    g20670(.A(new_n23106_), .B(new_n6255_), .Y(new_n23107_));
  AND2X1   g20671(.A(new_n23107_), .B(pi0907), .Y(new_n23108_));
  MX2X1    g20672(.A(new_n2777_), .B(new_n21904_), .S0(new_n11899_), .Y(new_n23109_));
  OAI21X1  g20673(.A0(new_n23109_), .A1(new_n6256_), .B0(new_n23108_), .Y(new_n23110_));
  NAND3X1  g20674(.A(new_n23110_), .B(new_n23105_), .C(new_n5362_), .Y(new_n23111_));
  MX2X1    g20675(.A(new_n21784_), .B(new_n2777_), .S0(new_n11825_), .Y(new_n23112_));
  AOI21X1  g20676(.A0(new_n23112_), .A1(new_n5021_), .B0(new_n5362_), .Y(new_n23113_));
  INVX1    g20677(.A(new_n23112_), .Y(new_n23114_));
  OAI21X1  g20678(.A0(new_n23114_), .A1(new_n5021_), .B0(new_n6256_), .Y(new_n23115_));
  MX2X1    g20679(.A(new_n2777_), .B(new_n21784_), .S0(new_n11899_), .Y(new_n23116_));
  OAI21X1  g20680(.A0(new_n23116_), .A1(new_n5023_), .B0(new_n23115_), .Y(new_n23117_));
  AOI21X1  g20681(.A0(new_n23117_), .A1(new_n23113_), .B0(new_n5042_), .Y(new_n23118_));
  AOI21X1  g20682(.A0(new_n23106_), .A1(new_n5043_), .B0(new_n5277_), .Y(new_n23119_));
  INVX1    g20683(.A(new_n23119_), .Y(new_n23120_));
  AOI21X1  g20684(.A0(new_n23109_), .A1(new_n5044_), .B0(new_n23120_), .Y(new_n23121_));
  NOR3X1   g20685(.A(new_n11976_), .B(pi0907), .C(new_n2777_), .Y(new_n23122_));
  OAI21X1  g20686(.A0(new_n23122_), .A1(new_n23121_), .B0(new_n5362_), .Y(new_n23123_));
  OAI21X1  g20687(.A0(new_n23114_), .A1(new_n5044_), .B0(pi0947), .Y(new_n23124_));
  AOI21X1  g20688(.A0(new_n23116_), .A1(new_n5044_), .B0(new_n23124_), .Y(new_n23125_));
  NOR2X1   g20689(.A(new_n23125_), .B(new_n5041_), .Y(new_n23126_));
  AOI22X1  g20690(.A0(new_n23126_), .A1(new_n23123_), .B0(new_n23118_), .B1(new_n23111_), .Y(new_n23127_));
  MX2X1    g20691(.A(new_n23099_), .B(new_n2777_), .S0(new_n11825_), .Y(new_n23128_));
  AOI21X1  g20692(.A0(new_n23128_), .A1(new_n2951_), .B0(pi0223), .Y(new_n23129_));
  OAI21X1  g20693(.A0(new_n23127_), .A1(new_n2951_), .B0(new_n23129_), .Y(new_n23130_));
  MX2X1    g20694(.A(pi0634), .B(pi0210), .S0(new_n11835_), .Y(new_n23131_));
  OAI21X1  g20695(.A0(new_n23131_), .A1(new_n5043_), .B0(new_n23119_), .Y(new_n23132_));
  NOR3X1   g20696(.A(new_n11824_), .B(new_n5044_), .C(new_n2725_), .Y(new_n23133_));
  OR4X1    g20697(.A(new_n23133_), .B(new_n11834_), .C(new_n11831_), .D(new_n2777_), .Y(new_n23134_));
  AOI21X1  g20698(.A0(new_n23134_), .A1(new_n23132_), .B0(pi0947), .Y(new_n23135_));
  MX2X1    g20699(.A(new_n21784_), .B(new_n2777_), .S0(new_n11835_), .Y(new_n23136_));
  AOI21X1  g20700(.A0(new_n23136_), .A1(new_n5044_), .B0(new_n23124_), .Y(new_n23137_));
  OR3X1    g20701(.A(new_n23137_), .B(new_n23135_), .C(new_n5041_), .Y(new_n23138_));
  INVX1    g20702(.A(new_n12008_), .Y(new_n23139_));
  AOI22X1  g20703(.A0(new_n23103_), .A1(new_n23139_), .B0(new_n23102_), .B1(new_n5021_), .Y(new_n23140_));
  NAND2X1  g20704(.A(new_n23140_), .B(new_n5277_), .Y(new_n23141_));
  NAND2X1  g20705(.A(new_n23131_), .B(new_n6255_), .Y(new_n23142_));
  AOI21X1  g20706(.A0(new_n23142_), .A1(new_n23108_), .B0(pi0947), .Y(new_n23143_));
  NAND2X1  g20707(.A(new_n23143_), .B(new_n23141_), .Y(new_n23144_));
  OAI21X1  g20708(.A0(new_n23136_), .A1(new_n5023_), .B0(new_n23115_), .Y(new_n23145_));
  AOI21X1  g20709(.A0(new_n23145_), .A1(new_n23113_), .B0(new_n5042_), .Y(new_n23146_));
  AOI21X1  g20710(.A0(new_n23146_), .A1(new_n23144_), .B0(new_n2940_), .Y(new_n23147_));
  AOI21X1  g20711(.A0(new_n23147_), .A1(new_n23138_), .B0(pi0299), .Y(new_n23148_));
  AND2X1   g20712(.A(new_n23148_), .B(new_n23130_), .Y(new_n23149_));
  OAI21X1  g20713(.A0(new_n11976_), .A1(new_n2777_), .B0(new_n11952_), .Y(new_n23150_));
  AOI21X1  g20714(.A0(new_n23104_), .A1(new_n5057_), .B0(pi0907), .Y(new_n23151_));
  AOI21X1  g20715(.A0(new_n23151_), .A1(new_n23150_), .B0(new_n23121_), .Y(new_n23152_));
  NOR2X1   g20716(.A(new_n23125_), .B(new_n10044_), .Y(new_n23153_));
  OAI21X1  g20717(.A0(new_n23152_), .A1(pi0947), .B0(new_n23153_), .Y(new_n23154_));
  AOI21X1  g20718(.A0(new_n23128_), .A1(new_n10044_), .B0(pi0215), .Y(new_n23155_));
  AND2X1   g20719(.A(new_n23140_), .B(new_n5057_), .Y(new_n23156_));
  AND2X1   g20720(.A(new_n23134_), .B(new_n11952_), .Y(new_n23157_));
  OR2X1    g20721(.A(new_n23157_), .B(pi0907), .Y(new_n23158_));
  OAI21X1  g20722(.A0(new_n23158_), .A1(new_n23156_), .B0(new_n23132_), .Y(new_n23159_));
  AOI21X1  g20723(.A0(new_n23159_), .A1(new_n5362_), .B0(new_n23137_), .Y(new_n23160_));
  OAI21X1  g20724(.A0(new_n23160_), .A1(new_n2934_), .B0(pi0299), .Y(new_n23161_));
  AOI21X1  g20725(.A0(new_n23155_), .A1(new_n23154_), .B0(new_n23161_), .Y(new_n23162_));
  OR3X1    g20726(.A(new_n23162_), .B(new_n23149_), .C(new_n2939_), .Y(new_n23163_));
  INVX1    g20727(.A(new_n23099_), .Y(new_n23164_));
  AOI21X1  g20728(.A0(new_n23164_), .A1(new_n11820_), .B0(pi0299), .Y(new_n23165_));
  OAI21X1  g20729(.A0(new_n11820_), .A1(new_n2777_), .B0(new_n23165_), .Y(new_n23166_));
  AOI21X1  g20730(.A0(new_n23164_), .A1(new_n11960_), .B0(new_n2933_), .Y(new_n23167_));
  OAI21X1  g20731(.A0(new_n11818_), .A1(new_n2777_), .B0(new_n23167_), .Y(new_n23168_));
  AND2X1   g20732(.A(new_n23168_), .B(new_n2939_), .Y(new_n23169_));
  AOI21X1  g20733(.A0(new_n23169_), .A1(new_n23166_), .B0(pi0038), .Y(new_n23170_));
  AOI21X1  g20734(.A0(new_n23170_), .A1(new_n23163_), .B0(new_n23101_), .Y(new_n23171_));
  MX2X1    g20735(.A(new_n23171_), .B(pi0210), .S0(new_n9483_), .Y(po0367));
  INVX1    g20736(.A(pi0211), .Y(new_n23173_));
  OR2X1    g20737(.A(new_n14941_), .B(new_n11770_), .Y(new_n23174_));
  AND2X1   g20738(.A(new_n14939_), .B(new_n3103_), .Y(new_n23175_));
  AOI21X1  g20739(.A0(new_n23175_), .A1(pi0606), .B0(new_n22368_), .Y(new_n23176_));
  OAI21X1  g20740(.A0(new_n23174_), .A1(pi0606), .B0(new_n23176_), .Y(new_n23177_));
  OAI21X1  g20741(.A0(new_n14519_), .A1(new_n14518_), .B0(new_n3103_), .Y(new_n23178_));
  AOI21X1  g20742(.A0(new_n22662_), .A1(new_n22299_), .B0(pi0643), .Y(new_n23179_));
  OAI21X1  g20743(.A0(new_n23178_), .A1(new_n22299_), .B0(new_n23179_), .Y(new_n23180_));
  AND3X1   g20744(.A(new_n23180_), .B(new_n23177_), .C(new_n6489_), .Y(new_n23181_));
  NAND2X1  g20745(.A(new_n14932_), .B(new_n3103_), .Y(new_n23182_));
  AND2X1   g20746(.A(new_n14930_), .B(new_n3103_), .Y(new_n23183_));
  OAI21X1  g20747(.A0(new_n23183_), .A1(new_n22299_), .B0(pi0643), .Y(new_n23184_));
  AOI21X1  g20748(.A0(new_n23182_), .A1(new_n22299_), .B0(new_n23184_), .Y(new_n23185_));
  AND3X1   g20749(.A(new_n14536_), .B(new_n14523_), .C(new_n3103_), .Y(new_n23186_));
  AND3X1   g20750(.A(new_n23186_), .B(new_n22368_), .C(pi0606), .Y(new_n23187_));
  AND3X1   g20751(.A(new_n5102_), .B(new_n23173_), .C(new_n2436_), .Y(new_n23188_));
  OAI21X1  g20752(.A0(new_n23187_), .A1(new_n23185_), .B0(new_n23188_), .Y(new_n23189_));
  OAI21X1  g20753(.A0(new_n23181_), .A1(new_n23173_), .B0(new_n23189_), .Y(po0368));
  AOI21X1  g20754(.A0(new_n23175_), .A1(pi0607), .B0(new_n22966_), .Y(new_n23191_));
  OAI21X1  g20755(.A0(new_n23174_), .A1(pi0607), .B0(new_n23191_), .Y(new_n23192_));
  AOI21X1  g20756(.A0(new_n22662_), .A1(new_n22960_), .B0(pi0638), .Y(new_n23193_));
  OAI21X1  g20757(.A0(new_n23178_), .A1(new_n22960_), .B0(new_n23193_), .Y(new_n23194_));
  AND3X1   g20758(.A(new_n23194_), .B(new_n23192_), .C(new_n6489_), .Y(new_n23195_));
  OR2X1    g20759(.A(new_n23183_), .B(new_n22960_), .Y(new_n23196_));
  AOI21X1  g20760(.A0(new_n23182_), .A1(new_n22960_), .B0(new_n22966_), .Y(new_n23197_));
  AND2X1   g20761(.A(new_n22966_), .B(pi0607), .Y(new_n23198_));
  AOI22X1  g20762(.A0(new_n23198_), .A1(new_n23186_), .B0(new_n23197_), .B1(new_n23196_), .Y(new_n23199_));
  NAND3X1  g20763(.A(new_n5102_), .B(pi0212), .C(new_n2436_), .Y(new_n23200_));
  OAI22X1  g20764(.A0(new_n23200_), .A1(new_n23199_), .B0(new_n23195_), .B1(pi0212), .Y(po0369));
  AND3X1   g20765(.A(new_n5102_), .B(pi0213), .C(new_n2436_), .Y(new_n23202_));
  INVX1    g20766(.A(new_n23202_), .Y(new_n23203_));
  OR2X1    g20767(.A(new_n23183_), .B(new_n23047_), .Y(new_n23204_));
  AOI21X1  g20768(.A0(new_n23182_), .A1(new_n23047_), .B0(new_n23002_), .Y(new_n23205_));
  AND2X1   g20769(.A(new_n23002_), .B(pi0622), .Y(new_n23206_));
  AOI22X1  g20770(.A0(new_n23206_), .A1(new_n23186_), .B0(new_n23205_), .B1(new_n23204_), .Y(new_n23207_));
  AOI21X1  g20771(.A0(new_n23175_), .A1(pi0639), .B0(new_n23047_), .Y(new_n23208_));
  OAI21X1  g20772(.A0(new_n23178_), .A1(pi0639), .B0(new_n23208_), .Y(new_n23209_));
  AOI21X1  g20773(.A0(new_n22662_), .A1(new_n23002_), .B0(pi0622), .Y(new_n23210_));
  OAI21X1  g20774(.A0(new_n23174_), .A1(new_n23002_), .B0(new_n23210_), .Y(new_n23211_));
  AND3X1   g20775(.A(new_n23211_), .B(new_n23209_), .C(new_n6489_), .Y(new_n23212_));
  OAI22X1  g20776(.A0(new_n23212_), .A1(pi0213), .B0(new_n23207_), .B1(new_n23203_), .Y(po0370));
  AOI21X1  g20777(.A0(new_n23175_), .A1(pi0623), .B0(new_n22697_), .Y(new_n23214_));
  OAI21X1  g20778(.A0(new_n23174_), .A1(pi0623), .B0(new_n23214_), .Y(new_n23215_));
  AOI21X1  g20779(.A0(new_n22662_), .A1(new_n22661_), .B0(pi0710), .Y(new_n23216_));
  OAI21X1  g20780(.A0(new_n23178_), .A1(new_n22661_), .B0(new_n23216_), .Y(new_n23217_));
  AND3X1   g20781(.A(new_n23217_), .B(new_n23215_), .C(new_n6489_), .Y(new_n23218_));
  OR2X1    g20782(.A(new_n23183_), .B(new_n22661_), .Y(new_n23219_));
  AOI21X1  g20783(.A0(new_n23182_), .A1(new_n22661_), .B0(new_n22697_), .Y(new_n23220_));
  AND2X1   g20784(.A(new_n22697_), .B(pi0623), .Y(new_n23221_));
  AOI22X1  g20785(.A0(new_n23221_), .A1(new_n23186_), .B0(new_n23220_), .B1(new_n23219_), .Y(new_n23222_));
  NAND3X1  g20786(.A(new_n5102_), .B(pi0214), .C(new_n2436_), .Y(new_n23223_));
  OAI22X1  g20787(.A0(new_n23223_), .A1(new_n23222_), .B0(new_n23218_), .B1(pi0214), .Y(po0371));
  NOR3X1   g20788(.A(new_n14513_), .B(new_n11955_), .C(pi0947), .Y(new_n23225_));
  INVX1    g20789(.A(new_n23225_), .Y(new_n23226_));
  AND2X1   g20790(.A(pi0907), .B(pi0681), .Y(new_n23227_));
  AND2X1   g20791(.A(new_n23227_), .B(new_n5362_), .Y(new_n23228_));
  INVX1    g20792(.A(new_n11846_), .Y(new_n23229_));
  NOR2X1   g20793(.A(pi0681), .B(pi0661), .Y(new_n23230_));
  AOI21X1  g20794(.A0(new_n23230_), .A1(new_n11856_), .B0(pi0642), .Y(new_n23231_));
  OAI21X1  g20795(.A0(new_n23229_), .A1(new_n5020_), .B0(new_n23231_), .Y(new_n23232_));
  AOI21X1  g20796(.A0(new_n23232_), .A1(pi0947), .B0(new_n23228_), .Y(new_n23233_));
  AOI21X1  g20797(.A0(new_n23233_), .A1(new_n23226_), .B0(new_n2933_), .Y(new_n23234_));
  INVX1    g20798(.A(new_n23227_), .Y(new_n23235_));
  AND3X1   g20799(.A(new_n23235_), .B(new_n11933_), .C(new_n5362_), .Y(new_n23236_));
  AOI21X1  g20800(.A0(new_n11976_), .A1(new_n5016_), .B0(new_n5041_), .Y(new_n23237_));
  OAI21X1  g20801(.A0(new_n11917_), .A1(pi0642), .B0(new_n5020_), .Y(new_n23238_));
  NOR3X1   g20802(.A(new_n11824_), .B(new_n5017_), .C(new_n2725_), .Y(new_n23239_));
  AOI21X1  g20803(.A0(new_n23239_), .A1(new_n5016_), .B0(new_n5020_), .Y(new_n23240_));
  OAI21X1  g20804(.A0(new_n12001_), .A1(new_n11938_), .B0(new_n23240_), .Y(new_n23241_));
  AOI21X1  g20805(.A0(new_n23241_), .A1(new_n23238_), .B0(new_n5042_), .Y(new_n23242_));
  NOR3X1   g20806(.A(new_n23242_), .B(new_n23237_), .C(new_n5362_), .Y(new_n23243_));
  OR2X1    g20807(.A(new_n23243_), .B(new_n2951_), .Y(new_n23244_));
  AND2X1   g20808(.A(new_n11825_), .B(new_n2951_), .Y(new_n23245_));
  MX2X1    g20809(.A(new_n23235_), .B(new_n5016_), .S0(pi0947), .Y(new_n23246_));
  NOR2X1   g20810(.A(new_n23246_), .B(new_n2952_), .Y(new_n23247_));
  NOR3X1   g20811(.A(new_n23247_), .B(new_n23245_), .C(pi0223), .Y(new_n23248_));
  OAI21X1  g20812(.A0(new_n23244_), .A1(new_n23236_), .B0(new_n23248_), .Y(new_n23249_));
  INVX1    g20813(.A(new_n11878_), .Y(new_n23250_));
  OAI21X1  g20814(.A0(new_n12008_), .A1(new_n5262_), .B0(new_n5016_), .Y(new_n23251_));
  AOI21X1  g20815(.A0(new_n11854_), .A1(new_n5262_), .B0(new_n23251_), .Y(new_n23252_));
  AOI21X1  g20816(.A0(new_n23232_), .A1(new_n5042_), .B0(new_n5362_), .Y(new_n23253_));
  OAI21X1  g20817(.A0(new_n23252_), .A1(new_n5042_), .B0(new_n23253_), .Y(new_n23254_));
  OAI21X1  g20818(.A0(new_n23250_), .A1(pi0947), .B0(new_n23254_), .Y(new_n23255_));
  AOI21X1  g20819(.A0(new_n23227_), .A1(new_n5362_), .B0(new_n2940_), .Y(new_n23256_));
  AOI21X1  g20820(.A0(new_n23256_), .A1(new_n23255_), .B0(pi0299), .Y(new_n23257_));
  AOI21X1  g20821(.A0(new_n23257_), .A1(new_n23249_), .B0(new_n23234_), .Y(new_n23258_));
  NOR2X1   g20822(.A(new_n11863_), .B(new_n5016_), .Y(new_n23259_));
  NOR2X1   g20823(.A(new_n11900_), .B(new_n5019_), .Y(new_n23260_));
  NOR4X1   g20824(.A(new_n23260_), .B(new_n11872_), .C(new_n11867_), .D(new_n5016_), .Y(new_n23261_));
  AOI21X1  g20825(.A0(new_n23259_), .A1(new_n11880_), .B0(new_n23261_), .Y(new_n23262_));
  OAI21X1  g20826(.A0(new_n23262_), .A1(new_n5362_), .B0(new_n5041_), .Y(new_n23263_));
  AOI21X1  g20827(.A0(new_n23228_), .A1(new_n11941_), .B0(new_n23263_), .Y(new_n23264_));
  AOI21X1  g20828(.A0(new_n23227_), .A1(new_n11926_), .B0(pi0947), .Y(new_n23265_));
  MX2X1    g20829(.A(new_n11925_), .B(new_n11899_), .S0(new_n5020_), .Y(new_n23266_));
  NAND3X1  g20830(.A(new_n23266_), .B(new_n11863_), .C(pi0642), .Y(new_n23267_));
  AOI21X1  g20831(.A0(new_n23259_), .A1(new_n11925_), .B0(new_n5362_), .Y(new_n23268_));
  AOI21X1  g20832(.A0(new_n23268_), .A1(new_n23267_), .B0(new_n23265_), .Y(new_n23269_));
  OAI21X1  g20833(.A0(new_n23269_), .A1(new_n5041_), .B0(new_n2952_), .Y(new_n23270_));
  AOI21X1  g20834(.A0(new_n23247_), .A1(new_n11880_), .B0(pi0223), .Y(new_n23271_));
  OAI21X1  g20835(.A0(new_n23270_), .A1(new_n23264_), .B0(new_n23271_), .Y(new_n23272_));
  AOI21X1  g20836(.A0(new_n11854_), .A1(new_n5041_), .B0(new_n23235_), .Y(new_n23273_));
  NOR2X1   g20837(.A(new_n23273_), .B(pi0947), .Y(new_n23274_));
  OAI21X1  g20838(.A0(new_n11836_), .A1(new_n5362_), .B0(new_n11846_), .Y(new_n23275_));
  NOR4X1   g20839(.A(new_n11872_), .B(new_n11868_), .C(new_n11867_), .D(new_n5016_), .Y(new_n23276_));
  INVX1    g20840(.A(new_n23259_), .Y(new_n23277_));
  OAI21X1  g20841(.A0(new_n23277_), .A1(new_n11825_), .B0(pi0947), .Y(new_n23278_));
  OAI22X1  g20842(.A0(new_n23278_), .A1(new_n23276_), .B0(new_n23275_), .B1(new_n5041_), .Y(new_n23279_));
  OAI21X1  g20843(.A0(new_n23279_), .A1(new_n23274_), .B0(pi0223), .Y(new_n23280_));
  AOI21X1  g20844(.A0(new_n23280_), .A1(new_n23272_), .B0(pi0299), .Y(new_n23281_));
  OAI21X1  g20845(.A0(new_n23246_), .A1(new_n11948_), .B0(pi0299), .Y(new_n23282_));
  AOI21X1  g20846(.A0(new_n23269_), .A1(new_n10045_), .B0(new_n23282_), .Y(new_n23283_));
  OR3X1    g20847(.A(new_n23283_), .B(new_n23281_), .C(pi0215), .Y(new_n23284_));
  OAI21X1  g20848(.A0(new_n23258_), .A1(new_n2934_), .B0(new_n23284_), .Y(new_n23285_));
  OAI21X1  g20849(.A0(new_n23246_), .A1(new_n11961_), .B0(pi0299), .Y(new_n23286_));
  AOI21X1  g20850(.A0(new_n11961_), .A1(pi0215), .B0(new_n23286_), .Y(new_n23287_));
  NOR2X1   g20851(.A(new_n23246_), .B(new_n12306_), .Y(new_n23288_));
  OAI21X1  g20852(.A0(new_n11820_), .A1(new_n2934_), .B0(new_n2933_), .Y(new_n23289_));
  OAI21X1  g20853(.A0(new_n23289_), .A1(new_n23288_), .B0(new_n2939_), .Y(new_n23290_));
  OAI21X1  g20854(.A0(new_n23290_), .A1(new_n23287_), .B0(new_n2979_), .Y(new_n23291_));
  AOI21X1  g20855(.A0(new_n23285_), .A1(pi0039), .B0(new_n23291_), .Y(new_n23292_));
  NOR4X1   g20856(.A(new_n23246_), .B(new_n2986_), .C(new_n2725_), .D(pi0039), .Y(new_n23293_));
  OAI21X1  g20857(.A0(new_n12077_), .A1(new_n2934_), .B0(pi0038), .Y(new_n23294_));
  OAI21X1  g20858(.A0(new_n23294_), .A1(new_n23293_), .B0(new_n7625_), .Y(new_n23295_));
  OAI22X1  g20859(.A0(new_n23295_), .A1(new_n23292_), .B0(new_n7625_), .B1(new_n2934_), .Y(po0372));
  NAND2X1  g20860(.A(pi0907), .B(pi0662), .Y(new_n23297_));
  MX2X1    g20861(.A(new_n23297_), .B(new_n11838_), .S0(pi0947), .Y(new_n23298_));
  AOI21X1  g20862(.A0(new_n12771_), .A1(pi0216), .B0(new_n2979_), .Y(new_n23299_));
  OAI21X1  g20863(.A0(new_n23298_), .A1(new_n12771_), .B0(new_n23299_), .Y(new_n23300_));
  NAND2X1  g20864(.A(new_n14510_), .B(new_n5362_), .Y(new_n23301_));
  NOR2X1   g20865(.A(new_n23297_), .B(pi0947), .Y(new_n23302_));
  AOI21X1  g20866(.A0(new_n11976_), .A1(new_n11838_), .B0(new_n5362_), .Y(new_n23303_));
  NOR2X1   g20867(.A(new_n23303_), .B(new_n23302_), .Y(new_n23304_));
  AOI21X1  g20868(.A0(new_n23304_), .A1(new_n23301_), .B0(new_n2438_), .Y(new_n23305_));
  AND2X1   g20869(.A(pi0947), .B(pi0614), .Y(new_n23306_));
  AOI22X1  g20870(.A0(new_n23306_), .A1(new_n23266_), .B0(new_n23302_), .B1(new_n11926_), .Y(new_n23307_));
  OAI22X1  g20871(.A0(new_n23307_), .A1(new_n11419_), .B0(new_n23298_), .B1(new_n11948_), .Y(new_n23308_));
  OAI21X1  g20872(.A0(new_n23308_), .A1(new_n23305_), .B0(new_n2934_), .Y(new_n23309_));
  AOI22X1  g20873(.A0(new_n12195_), .A1(new_n5018_), .B0(new_n11871_), .B1(pi0614), .Y(new_n23310_));
  OAI21X1  g20874(.A0(new_n11836_), .A1(new_n5018_), .B0(new_n23310_), .Y(new_n23311_));
  NOR2X1   g20875(.A(new_n11835_), .B(pi0614), .Y(new_n23312_));
  AOI22X1  g20876(.A0(new_n23312_), .A1(new_n5020_), .B0(new_n23311_), .B1(new_n11905_), .Y(new_n23313_));
  AND2X1   g20877(.A(new_n23313_), .B(pi0947), .Y(new_n23314_));
  OR3X1    g20878(.A(new_n23314_), .B(new_n23302_), .C(new_n2438_), .Y(new_n23315_));
  OAI21X1  g20879(.A0(new_n23297_), .A1(new_n11846_), .B0(new_n5362_), .Y(new_n23316_));
  NOR2X1   g20880(.A(new_n11921_), .B(new_n5362_), .Y(new_n23317_));
  OAI21X1  g20881(.A0(new_n11919_), .A1(new_n11868_), .B0(new_n23317_), .Y(new_n23318_));
  NAND2X1  g20882(.A(new_n11836_), .B(pi0947), .Y(new_n23319_));
  NAND3X1  g20883(.A(new_n23319_), .B(new_n23318_), .C(new_n23316_), .Y(new_n23320_));
  AOI21X1  g20884(.A0(new_n23320_), .A1(new_n2438_), .B0(new_n2934_), .Y(new_n23321_));
  OAI21X1  g20885(.A0(new_n23315_), .A1(new_n23225_), .B0(new_n23321_), .Y(new_n23322_));
  AND3X1   g20886(.A(new_n23322_), .B(new_n23309_), .C(pi0299), .Y(new_n23323_));
  OR2X1    g20887(.A(new_n11908_), .B(new_n11907_), .Y(new_n23324_));
  AND2X1   g20888(.A(new_n11924_), .B(new_n5362_), .Y(new_n23325_));
  AOI22X1  g20889(.A0(new_n23325_), .A1(new_n23297_), .B0(new_n23324_), .B1(pi0947), .Y(new_n23326_));
  OAI21X1  g20890(.A0(new_n11931_), .A1(new_n11927_), .B0(new_n5362_), .Y(new_n23327_));
  NOR3X1   g20891(.A(new_n23303_), .B(new_n23302_), .C(new_n5041_), .Y(new_n23328_));
  AOI21X1  g20892(.A0(new_n23328_), .A1(new_n23327_), .B0(new_n2951_), .Y(new_n23329_));
  OAI21X1  g20893(.A0(new_n23326_), .A1(new_n5042_), .B0(new_n23329_), .Y(new_n23330_));
  OAI21X1  g20894(.A0(new_n23298_), .A1(new_n2952_), .B0(new_n2940_), .Y(new_n23331_));
  AOI21X1  g20895(.A0(new_n11825_), .A1(new_n2951_), .B0(new_n23331_), .Y(new_n23332_));
  OR3X1    g20896(.A(new_n11844_), .B(new_n11841_), .C(pi0616), .Y(new_n23333_));
  AND3X1   g20897(.A(new_n23333_), .B(new_n11874_), .C(new_n5262_), .Y(new_n23334_));
  OAI21X1  g20898(.A0(new_n12008_), .A1(new_n5262_), .B0(new_n11838_), .Y(new_n23335_));
  OAI21X1  g20899(.A0(new_n23335_), .A1(new_n23334_), .B0(new_n5041_), .Y(new_n23336_));
  AOI21X1  g20900(.A0(new_n23313_), .A1(new_n5042_), .B0(new_n5362_), .Y(new_n23337_));
  AOI22X1  g20901(.A0(new_n23337_), .A1(new_n23336_), .B0(new_n11878_), .B1(new_n5362_), .Y(new_n23338_));
  OAI21X1  g20902(.A0(new_n23297_), .A1(pi0947), .B0(pi0223), .Y(new_n23339_));
  OAI21X1  g20903(.A0(new_n23339_), .A1(new_n23338_), .B0(pi0216), .Y(new_n23340_));
  AOI21X1  g20904(.A0(new_n23332_), .A1(new_n23330_), .B0(new_n23340_), .Y(new_n23341_));
  INVX1    g20905(.A(new_n23302_), .Y(new_n23342_));
  AOI21X1  g20906(.A0(new_n11922_), .A1(pi0947), .B0(new_n5042_), .Y(new_n23343_));
  OAI21X1  g20907(.A0(new_n23342_), .A1(new_n11904_), .B0(new_n23343_), .Y(new_n23344_));
  AOI21X1  g20908(.A0(new_n23307_), .A1(new_n5042_), .B0(new_n2951_), .Y(new_n23345_));
  OR2X1    g20909(.A(new_n23298_), .B(new_n2952_), .Y(new_n23346_));
  OAI21X1  g20910(.A0(new_n23346_), .A1(new_n11825_), .B0(new_n2940_), .Y(new_n23347_));
  AOI21X1  g20911(.A0(new_n23345_), .A1(new_n23344_), .B0(new_n23347_), .Y(new_n23348_));
  OR2X1    g20912(.A(new_n23275_), .B(new_n5041_), .Y(new_n23349_));
  AND2X1   g20913(.A(new_n11854_), .B(new_n5041_), .Y(new_n23350_));
  OAI21X1  g20914(.A0(new_n23297_), .A1(new_n23350_), .B0(new_n5362_), .Y(new_n23351_));
  AND3X1   g20915(.A(new_n23351_), .B(new_n23318_), .C(new_n23349_), .Y(new_n23352_));
  OAI21X1  g20916(.A0(new_n23352_), .A1(new_n2940_), .B0(new_n2438_), .Y(new_n23353_));
  OAI21X1  g20917(.A0(new_n23353_), .A1(new_n23348_), .B0(new_n2933_), .Y(new_n23354_));
  OAI21X1  g20918(.A0(new_n23354_), .A1(new_n23341_), .B0(pi0039), .Y(new_n23355_));
  AND2X1   g20919(.A(new_n11961_), .B(pi0216), .Y(new_n23356_));
  OAI21X1  g20920(.A0(new_n23298_), .A1(new_n11961_), .B0(pi0299), .Y(new_n23357_));
  OR2X1    g20921(.A(new_n23357_), .B(new_n23356_), .Y(new_n23358_));
  OR2X1    g20922(.A(new_n23298_), .B(new_n12306_), .Y(new_n23359_));
  AOI21X1  g20923(.A0(new_n12306_), .A1(pi0216), .B0(pi0299), .Y(new_n23360_));
  AOI21X1  g20924(.A0(new_n23360_), .A1(new_n23359_), .B0(pi0039), .Y(new_n23361_));
  AOI21X1  g20925(.A0(new_n23361_), .A1(new_n23358_), .B0(pi0038), .Y(new_n23362_));
  OAI21X1  g20926(.A0(new_n23355_), .A1(new_n23323_), .B0(new_n23362_), .Y(new_n23363_));
  AND2X1   g20927(.A(new_n23363_), .B(new_n23300_), .Y(new_n23364_));
  MX2X1    g20928(.A(new_n23364_), .B(pi0216), .S0(new_n9483_), .Y(po0373));
  INVX1    g20929(.A(pi0695), .Y(new_n23366_));
  OR2X1    g20930(.A(new_n23022_), .B(new_n23021_), .Y(new_n23367_));
  OAI21X1  g20931(.A0(new_n23024_), .A1(new_n23366_), .B0(new_n9353_), .Y(new_n23368_));
  AOI21X1  g20932(.A0(new_n23367_), .A1(new_n23366_), .B0(new_n23368_), .Y(new_n23369_));
  INVX1    g20933(.A(pi0612), .Y(new_n23370_));
  AND3X1   g20934(.A(new_n23090_), .B(new_n23089_), .C(new_n23366_), .Y(new_n23371_));
  OAI21X1  g20935(.A0(new_n23371_), .A1(new_n9353_), .B0(new_n23370_), .Y(new_n23372_));
  NOR2X1   g20936(.A(new_n23045_), .B(pi0695), .Y(new_n23373_));
  OAI21X1  g20937(.A0(new_n23052_), .A1(new_n23366_), .B0(new_n9353_), .Y(new_n23374_));
  NOR2X1   g20938(.A(new_n23374_), .B(new_n23373_), .Y(new_n23375_));
  NOR4X1   g20939(.A(new_n23093_), .B(new_n23070_), .C(po1038), .D(new_n23366_), .Y(new_n23376_));
  OR2X1    g20940(.A(new_n23376_), .B(new_n9353_), .Y(new_n23377_));
  AOI21X1  g20941(.A0(new_n23080_), .A1(new_n23366_), .B0(new_n23377_), .Y(new_n23378_));
  OR3X1    g20942(.A(new_n23378_), .B(new_n23375_), .C(new_n23370_), .Y(new_n23379_));
  OAI21X1  g20943(.A0(new_n23372_), .A1(new_n23369_), .B0(new_n23379_), .Y(po0374));
  INVX1    g20944(.A(pi0218), .Y(new_n23381_));
  MX2X1    g20945(.A(new_n22644_), .B(new_n22607_), .S0(new_n22585_), .Y(new_n23382_));
  NOR4X1   g20946(.A(new_n22647_), .B(new_n22646_), .C(new_n22585_), .D(new_n22574_), .Y(new_n23383_));
  MX2X1    g20947(.A(new_n23383_), .B(new_n23382_), .S0(new_n23381_), .Y(po0375));
  NAND3X1  g20948(.A(new_n5102_), .B(new_n8422_), .C(new_n2436_), .Y(new_n23385_));
  OR2X1    g20949(.A(new_n23183_), .B(new_n22151_), .Y(new_n23386_));
  AOI21X1  g20950(.A0(new_n23182_), .A1(new_n22151_), .B0(new_n22139_), .Y(new_n23387_));
  AND2X1   g20951(.A(new_n22139_), .B(pi0617), .Y(new_n23388_));
  AOI22X1  g20952(.A0(new_n23388_), .A1(new_n23186_), .B0(new_n23387_), .B1(new_n23386_), .Y(new_n23389_));
  AOI21X1  g20953(.A0(new_n23175_), .A1(pi0617), .B0(new_n22139_), .Y(new_n23390_));
  OAI21X1  g20954(.A0(new_n23174_), .A1(pi0617), .B0(new_n23390_), .Y(new_n23391_));
  AOI21X1  g20955(.A0(new_n22662_), .A1(new_n22151_), .B0(pi0637), .Y(new_n23392_));
  OAI21X1  g20956(.A0(new_n23178_), .A1(new_n22151_), .B0(new_n23392_), .Y(new_n23393_));
  AND3X1   g20957(.A(new_n23393_), .B(new_n23391_), .C(new_n6489_), .Y(new_n23394_));
  OAI22X1  g20958(.A0(new_n23394_), .A1(new_n8422_), .B0(new_n23389_), .B1(new_n23385_), .Y(po0376));
  INVX1    g20959(.A(pi0220), .Y(new_n23396_));
  MX2X1    g20960(.A(new_n22570_), .B(new_n22478_), .S0(new_n22656_), .Y(new_n23397_));
  NOR4X1   g20961(.A(new_n22656_), .B(new_n22575_), .C(new_n22574_), .D(new_n22573_), .Y(new_n23398_));
  MX2X1    g20962(.A(new_n23398_), .B(new_n23397_), .S0(new_n23396_), .Y(po0377));
  AND2X1   g20963(.A(pi0907), .B(pi0661), .Y(new_n23400_));
  AND2X1   g20964(.A(pi0947), .B(pi0616), .Y(new_n23401_));
  AOI21X1  g20965(.A0(new_n23400_), .A1(new_n5362_), .B0(new_n23401_), .Y(new_n23402_));
  AOI21X1  g20966(.A0(new_n12771_), .A1(pi0221), .B0(new_n2979_), .Y(new_n23403_));
  OAI21X1  g20967(.A0(new_n23402_), .A1(new_n12771_), .B0(new_n23403_), .Y(new_n23404_));
  OR2X1    g20968(.A(new_n11903_), .B(new_n11864_), .Y(new_n23405_));
  NOR4X1   g20969(.A(pi0681), .B(pi0662), .C(pi0661), .D(pi0616), .Y(new_n23406_));
  OAI21X1  g20970(.A0(new_n11920_), .A1(new_n23324_), .B0(new_n23406_), .Y(new_n23407_));
  AOI21X1  g20971(.A0(new_n23407_), .A1(new_n23405_), .B0(new_n5362_), .Y(new_n23408_));
  OR3X1    g20972(.A(new_n23408_), .B(new_n23325_), .C(new_n5042_), .Y(new_n23409_));
  AND2X1   g20973(.A(new_n23400_), .B(new_n5362_), .Y(new_n23410_));
  MX2X1    g20974(.A(new_n11903_), .B(new_n11916_), .S0(new_n5023_), .Y(new_n23411_));
  OAI21X1  g20975(.A0(new_n13165_), .A1(pi0642), .B0(new_n23267_), .Y(new_n23412_));
  AOI21X1  g20976(.A0(new_n23412_), .A1(new_n23406_), .B0(new_n5362_), .Y(new_n23413_));
  OAI21X1  g20977(.A0(new_n23411_), .A1(new_n11864_), .B0(new_n23413_), .Y(new_n23414_));
  AOI21X1  g20978(.A0(new_n23414_), .A1(new_n23327_), .B0(new_n5041_), .Y(new_n23415_));
  NOR2X1   g20979(.A(new_n23415_), .B(new_n23410_), .Y(new_n23416_));
  AOI21X1  g20980(.A0(new_n23416_), .A1(new_n23409_), .B0(new_n2951_), .Y(new_n23417_));
  OR3X1    g20981(.A(new_n23402_), .B(new_n11824_), .C(new_n2725_), .Y(new_n23418_));
  OAI21X1  g20982(.A0(new_n23418_), .A1(new_n2952_), .B0(new_n2940_), .Y(new_n23419_));
  OR3X1    g20983(.A(new_n23419_), .B(new_n23417_), .C(new_n23245_), .Y(new_n23420_));
  AND2X1   g20984(.A(new_n11845_), .B(new_n11837_), .Y(new_n23421_));
  AOI21X1  g20985(.A0(new_n23230_), .A1(new_n11856_), .B0(pi0616), .Y(new_n23422_));
  OAI21X1  g20986(.A0(new_n23421_), .A1(new_n5020_), .B0(new_n23422_), .Y(new_n23423_));
  AND2X1   g20987(.A(new_n23423_), .B(pi0947), .Y(new_n23424_));
  AOI21X1  g20988(.A0(new_n11953_), .A1(new_n5362_), .B0(new_n23424_), .Y(new_n23425_));
  NAND2X1  g20989(.A(new_n11877_), .B(new_n5362_), .Y(new_n23426_));
  OAI21X1  g20990(.A0(new_n11870_), .A1(new_n11865_), .B0(pi0947), .Y(new_n23427_));
  AND2X1   g20991(.A(new_n23427_), .B(new_n5041_), .Y(new_n23428_));
  OR2X1    g20992(.A(new_n23410_), .B(new_n2940_), .Y(new_n23429_));
  AOI21X1  g20993(.A0(new_n23428_), .A1(new_n23426_), .B0(new_n23429_), .Y(new_n23430_));
  OAI21X1  g20994(.A0(new_n23425_), .A1(new_n5041_), .B0(new_n23430_), .Y(new_n23431_));
  AND2X1   g20995(.A(new_n23431_), .B(pi0221), .Y(new_n23432_));
  INVX1    g20996(.A(new_n23410_), .Y(new_n23433_));
  OAI22X1  g20997(.A0(new_n23260_), .A1(new_n11873_), .B0(new_n11874_), .B1(new_n11863_), .Y(new_n23434_));
  AOI21X1  g20998(.A0(new_n23434_), .A1(pi0947), .B0(new_n5042_), .Y(new_n23435_));
  OAI21X1  g20999(.A0(new_n23433_), .A1(new_n11904_), .B0(new_n23435_), .Y(new_n23436_));
  AOI22X1  g21000(.A0(new_n23401_), .A1(new_n23266_), .B0(new_n23410_), .B1(new_n11926_), .Y(new_n23437_));
  AOI21X1  g21001(.A0(new_n23437_), .A1(new_n5042_), .B0(new_n2951_), .Y(new_n23438_));
  AOI21X1  g21002(.A0(new_n23438_), .A1(new_n23436_), .B0(new_n23419_), .Y(new_n23439_));
  NAND2X1  g21003(.A(new_n11875_), .B(pi0947), .Y(new_n23440_));
  MX2X1    g21004(.A(new_n23400_), .B(new_n11875_), .S0(pi0947), .Y(new_n23441_));
  OAI21X1  g21005(.A0(new_n23275_), .A1(new_n5041_), .B0(new_n23441_), .Y(new_n23442_));
  AOI21X1  g21006(.A0(new_n23440_), .A1(new_n23350_), .B0(new_n23442_), .Y(new_n23443_));
  OAI21X1  g21007(.A0(new_n23443_), .A1(new_n2940_), .B0(new_n2437_), .Y(new_n23444_));
  OAI21X1  g21008(.A0(new_n23444_), .A1(new_n23439_), .B0(new_n2933_), .Y(new_n23445_));
  AOI21X1  g21009(.A0(new_n23432_), .A1(new_n23420_), .B0(new_n23445_), .Y(new_n23446_));
  OAI21X1  g21010(.A0(new_n23400_), .A1(new_n14510_), .B0(new_n5362_), .Y(new_n23447_));
  AND2X1   g21011(.A(new_n23414_), .B(pi0221), .Y(new_n23448_));
  NOR2X1   g21012(.A(new_n23437_), .B(new_n2438_), .Y(new_n23449_));
  OAI21X1  g21013(.A0(new_n23418_), .A1(pi0216), .B0(new_n2437_), .Y(new_n23450_));
  OAI21X1  g21014(.A0(new_n23450_), .A1(new_n23449_), .B0(new_n2934_), .Y(new_n23451_));
  AOI21X1  g21015(.A0(new_n23448_), .A1(new_n23447_), .B0(new_n23451_), .Y(new_n23452_));
  NOR4X1   g21016(.A(new_n23424_), .B(new_n23410_), .C(new_n23225_), .D(new_n2437_), .Y(new_n23453_));
  AOI21X1  g21017(.A0(new_n23441_), .A1(new_n23275_), .B0(pi0221), .Y(new_n23454_));
  OR2X1    g21018(.A(new_n23454_), .B(new_n2934_), .Y(new_n23455_));
  OAI21X1  g21019(.A0(new_n23455_), .A1(new_n23453_), .B0(pi0299), .Y(new_n23456_));
  OAI21X1  g21020(.A0(new_n23456_), .A1(new_n23452_), .B0(pi0039), .Y(new_n23457_));
  AND2X1   g21021(.A(new_n11961_), .B(pi0221), .Y(new_n23458_));
  OAI21X1  g21022(.A0(new_n23402_), .A1(new_n11961_), .B0(pi0299), .Y(new_n23459_));
  OR2X1    g21023(.A(new_n23459_), .B(new_n23458_), .Y(new_n23460_));
  OR2X1    g21024(.A(new_n23402_), .B(new_n12306_), .Y(new_n23461_));
  AOI21X1  g21025(.A0(new_n12306_), .A1(pi0221), .B0(pi0299), .Y(new_n23462_));
  AOI21X1  g21026(.A0(new_n23462_), .A1(new_n23461_), .B0(pi0039), .Y(new_n23463_));
  AOI21X1  g21027(.A0(new_n23463_), .A1(new_n23460_), .B0(pi0038), .Y(new_n23464_));
  OAI21X1  g21028(.A0(new_n23457_), .A1(new_n23446_), .B0(new_n23464_), .Y(new_n23465_));
  AND2X1   g21029(.A(new_n23465_), .B(new_n23404_), .Y(new_n23466_));
  MX2X1    g21030(.A(new_n23466_), .B(pi0221), .S0(new_n9483_), .Y(po0378));
  MX2X1    g21031(.A(new_n14779_), .B(new_n23250_), .S0(pi0223), .Y(new_n23468_));
  AOI21X1  g21032(.A0(new_n23468_), .A1(new_n2933_), .B0(new_n2939_), .Y(new_n23469_));
  OR2X1    g21033(.A(new_n12779_), .B(pi0038), .Y(new_n23470_));
  AOI21X1  g21034(.A0(new_n23469_), .A1(new_n11957_), .B0(new_n23470_), .Y(new_n23471_));
  NOR2X1   g21035(.A(new_n23471_), .B(new_n21749_), .Y(new_n23472_));
  NOR2X1   g21036(.A(new_n23472_), .B(new_n2941_), .Y(new_n23473_));
  OR2X1    g21037(.A(new_n3103_), .B(new_n2941_), .Y(new_n23474_));
  INVX1    g21038(.A(new_n23230_), .Y(new_n23475_));
  MX2X1    g21039(.A(new_n23411_), .B(new_n12156_), .S0(pi0616), .Y(new_n23476_));
  NOR3X1   g21040(.A(new_n11979_), .B(new_n11871_), .C(new_n11881_), .Y(new_n23477_));
  OAI21X1  g21041(.A0(new_n23477_), .A1(new_n11987_), .B0(new_n11986_), .Y(new_n23478_));
  AOI21X1  g21042(.A0(new_n23478_), .A1(new_n11850_), .B0(new_n23475_), .Y(new_n23479_));
  OAI21X1  g21043(.A0(new_n23476_), .A1(new_n11850_), .B0(new_n23479_), .Y(new_n23480_));
  INVX1    g21044(.A(new_n23480_), .Y(new_n23481_));
  AOI21X1  g21045(.A0(new_n23476_), .A1(new_n23475_), .B0(new_n23481_), .Y(new_n23482_));
  NAND2X1  g21046(.A(new_n23482_), .B(new_n5059_), .Y(new_n23483_));
  MX2X1    g21047(.A(new_n11992_), .B(new_n11940_), .S0(new_n11871_), .Y(new_n23484_));
  INVX1    g21048(.A(new_n23484_), .Y(new_n23485_));
  NOR3X1   g21049(.A(new_n23477_), .B(new_n5019_), .C(pi0662), .Y(new_n23486_));
  AOI21X1  g21050(.A0(new_n23486_), .A1(new_n11900_), .B0(new_n23475_), .Y(new_n23487_));
  OAI21X1  g21051(.A0(new_n23485_), .A1(new_n11850_), .B0(new_n23487_), .Y(new_n23488_));
  OAI21X1  g21052(.A0(new_n23484_), .A1(new_n23230_), .B0(new_n23488_), .Y(new_n23489_));
  OR2X1    g21053(.A(new_n23489_), .B(new_n5059_), .Y(new_n23490_));
  AND2X1   g21054(.A(new_n23490_), .B(pi0222), .Y(new_n23491_));
  AND2X1   g21055(.A(new_n23491_), .B(new_n23483_), .Y(new_n23492_));
  MX2X1    g21056(.A(new_n12050_), .B(new_n12047_), .S0(new_n5020_), .Y(new_n23493_));
  NOR2X1   g21057(.A(new_n23493_), .B(new_n11871_), .Y(new_n23494_));
  NOR2X1   g21058(.A(new_n23494_), .B(new_n5059_), .Y(new_n23495_));
  INVX1    g21059(.A(new_n23495_), .Y(new_n23496_));
  AND2X1   g21060(.A(new_n23477_), .B(new_n11925_), .Y(new_n23497_));
  INVX1    g21061(.A(new_n23497_), .Y(new_n23498_));
  INVX1    g21062(.A(new_n12134_), .Y(new_n23499_));
  AND3X1   g21063(.A(pi0680), .B(new_n11849_), .C(pi0616), .Y(new_n23500_));
  AOI21X1  g21064(.A0(new_n23500_), .A1(new_n23499_), .B0(new_n23475_), .Y(new_n23501_));
  OAI21X1  g21065(.A0(new_n23498_), .A1(new_n11850_), .B0(new_n23501_), .Y(new_n23502_));
  INVX1    g21066(.A(new_n23502_), .Y(new_n23503_));
  AOI21X1  g21067(.A0(new_n23498_), .A1(new_n23475_), .B0(new_n23503_), .Y(new_n23504_));
  OR2X1    g21068(.A(new_n23504_), .B(new_n5058_), .Y(new_n23505_));
  AND3X1   g21069(.A(new_n23505_), .B(new_n23496_), .C(new_n2941_), .Y(new_n23506_));
  NOR3X1   g21070(.A(new_n23506_), .B(new_n23492_), .C(new_n10044_), .Y(new_n23507_));
  NOR4X1   g21071(.A(new_n12048_), .B(new_n11824_), .C(new_n2725_), .D(new_n11871_), .Y(new_n23508_));
  INVX1    g21072(.A(new_n23508_), .Y(new_n23509_));
  AOI21X1  g21073(.A0(new_n11825_), .A1(pi0222), .B0(new_n10045_), .Y(new_n23510_));
  AOI21X1  g21074(.A0(new_n23510_), .A1(new_n23509_), .B0(pi0215), .Y(new_n23511_));
  INVX1    g21075(.A(new_n23511_), .Y(new_n23512_));
  OAI21X1  g21076(.A0(new_n11842_), .A1(new_n5262_), .B0(new_n12049_), .Y(new_n23513_));
  OR2X1    g21077(.A(new_n23513_), .B(new_n11871_), .Y(new_n23514_));
  NOR3X1   g21078(.A(new_n23514_), .B(new_n12389_), .C(pi0222), .Y(new_n23515_));
  AOI21X1  g21079(.A0(new_n12019_), .A1(pi0616), .B0(new_n11846_), .Y(new_n23516_));
  INVX1    g21080(.A(new_n23516_), .Y(new_n23517_));
  AOI21X1  g21081(.A0(new_n12019_), .A1(pi0616), .B0(new_n11856_), .Y(new_n23518_));
  OAI21X1  g21082(.A0(new_n23229_), .A1(new_n11850_), .B0(new_n23518_), .Y(new_n23519_));
  AND2X1   g21083(.A(new_n23519_), .B(new_n23230_), .Y(new_n23520_));
  AOI21X1  g21084(.A0(new_n23517_), .A1(new_n23475_), .B0(new_n23520_), .Y(new_n23521_));
  AND2X1   g21085(.A(new_n23521_), .B(new_n5059_), .Y(new_n23522_));
  INVX1    g21086(.A(new_n23522_), .Y(new_n23523_));
  AOI21X1  g21087(.A0(new_n11993_), .A1(pi0616), .B0(new_n11866_), .Y(new_n23524_));
  INVX1    g21088(.A(new_n23524_), .Y(new_n23525_));
  AOI21X1  g21089(.A0(new_n23486_), .A1(new_n12008_), .B0(new_n23475_), .Y(new_n23526_));
  OAI21X1  g21090(.A0(new_n23525_), .A1(new_n11850_), .B0(new_n23526_), .Y(new_n23527_));
  INVX1    g21091(.A(new_n23527_), .Y(new_n23528_));
  AOI21X1  g21092(.A0(new_n23525_), .A1(new_n23475_), .B0(new_n23528_), .Y(new_n23529_));
  AOI21X1  g21093(.A0(new_n23529_), .A1(new_n5058_), .B0(new_n2941_), .Y(new_n23530_));
  AOI21X1  g21094(.A0(new_n23530_), .A1(new_n23523_), .B0(new_n23515_), .Y(new_n23531_));
  OAI21X1  g21095(.A0(new_n23531_), .A1(new_n2934_), .B0(pi0299), .Y(new_n23532_));
  INVX1    g21096(.A(new_n23532_), .Y(new_n23533_));
  OAI21X1  g21097(.A0(new_n23512_), .A1(new_n23507_), .B0(new_n23533_), .Y(new_n23534_));
  OAI21X1  g21098(.A0(new_n23489_), .A1(new_n5042_), .B0(pi0222), .Y(new_n23535_));
  AOI21X1  g21099(.A0(new_n23482_), .A1(new_n5042_), .B0(new_n23535_), .Y(new_n23536_));
  OR3X1    g21100(.A(new_n23493_), .B(new_n5042_), .C(new_n11871_), .Y(new_n23537_));
  AOI21X1  g21101(.A0(new_n23504_), .A1(new_n5042_), .B0(new_n2942_), .Y(new_n23538_));
  AOI21X1  g21102(.A0(new_n23509_), .A1(new_n2942_), .B0(pi0222), .Y(new_n23539_));
  INVX1    g21103(.A(new_n23539_), .Y(new_n23540_));
  AOI21X1  g21104(.A0(new_n23538_), .A1(new_n23537_), .B0(new_n23540_), .Y(new_n23541_));
  NOR3X1   g21105(.A(new_n23541_), .B(new_n23536_), .C(pi0223), .Y(new_n23542_));
  NAND2X1  g21106(.A(new_n23521_), .B(new_n5042_), .Y(new_n23543_));
  AOI21X1  g21107(.A0(new_n23529_), .A1(new_n5041_), .B0(new_n2941_), .Y(new_n23544_));
  NOR3X1   g21108(.A(new_n23514_), .B(new_n12380_), .C(pi0222), .Y(new_n23545_));
  NOR2X1   g21109(.A(new_n23545_), .B(new_n2940_), .Y(new_n23546_));
  INVX1    g21110(.A(new_n23546_), .Y(new_n23547_));
  AOI21X1  g21111(.A0(new_n23544_), .A1(new_n23543_), .B0(new_n23547_), .Y(new_n23548_));
  OR2X1    g21112(.A(new_n23548_), .B(new_n23542_), .Y(new_n23549_));
  AOI21X1  g21113(.A0(new_n23549_), .A1(new_n2933_), .B0(new_n2939_), .Y(new_n23550_));
  NOR3X1   g21114(.A(new_n11974_), .B(new_n11967_), .C(new_n2941_), .Y(new_n23551_));
  AOI21X1  g21115(.A0(new_n16614_), .A1(new_n2941_), .B0(pi0039), .Y(new_n23552_));
  OAI21X1  g21116(.A0(new_n16614_), .A1(pi0616), .B0(new_n23552_), .Y(new_n23553_));
  OAI21X1  g21117(.A0(new_n23553_), .A1(new_n23551_), .B0(new_n2979_), .Y(new_n23554_));
  AOI21X1  g21118(.A0(new_n23550_), .A1(new_n23534_), .B0(new_n23554_), .Y(new_n23555_));
  AOI21X1  g21119(.A0(new_n12771_), .A1(pi0222), .B0(new_n2979_), .Y(new_n23556_));
  AND2X1   g21120(.A(new_n12079_), .B(pi0616), .Y(new_n23557_));
  INVX1    g21121(.A(new_n23557_), .Y(new_n23558_));
  AOI21X1  g21122(.A0(new_n23558_), .A1(new_n23556_), .B0(new_n11770_), .Y(new_n23559_));
  INVX1    g21123(.A(new_n23559_), .Y(new_n23560_));
  OAI21X1  g21124(.A0(new_n23560_), .A1(new_n23555_), .B0(new_n23474_), .Y(new_n23561_));
  MX2X1    g21125(.A(new_n23561_), .B(new_n23473_), .S0(new_n12473_), .Y(new_n23562_));
  INVX1    g21126(.A(new_n23473_), .Y(new_n23563_));
  AOI21X1  g21127(.A0(new_n23563_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n23564_));
  OAI21X1  g21128(.A0(new_n23562_), .A1(new_n12462_), .B0(new_n23564_), .Y(new_n23565_));
  AOI21X1  g21129(.A0(new_n23563_), .A1(pi0609), .B0(pi1155), .Y(new_n23566_));
  OAI21X1  g21130(.A0(new_n23562_), .A1(pi0609), .B0(new_n23566_), .Y(new_n23567_));
  NAND2X1  g21131(.A(new_n23567_), .B(new_n23565_), .Y(new_n23568_));
  MX2X1    g21132(.A(new_n23568_), .B(new_n23562_), .S0(new_n11768_), .Y(new_n23569_));
  AND2X1   g21133(.A(new_n23569_), .B(new_n11767_), .Y(new_n23570_));
  AOI21X1  g21134(.A0(new_n23563_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n23571_));
  OAI21X1  g21135(.A0(new_n23569_), .A1(new_n12486_), .B0(new_n23571_), .Y(new_n23572_));
  AOI21X1  g21136(.A0(new_n23563_), .A1(pi0618), .B0(pi1154), .Y(new_n23573_));
  OAI21X1  g21137(.A0(new_n23569_), .A1(pi0618), .B0(new_n23573_), .Y(new_n23574_));
  AOI21X1  g21138(.A0(new_n23574_), .A1(new_n23572_), .B0(new_n11767_), .Y(new_n23575_));
  OAI21X1  g21139(.A0(new_n23575_), .A1(new_n23570_), .B0(new_n11766_), .Y(new_n23576_));
  NOR3X1   g21140(.A(new_n23575_), .B(new_n23570_), .C(new_n12509_), .Y(new_n23577_));
  OAI21X1  g21141(.A0(new_n23473_), .A1(pi0619), .B0(pi1159), .Y(new_n23578_));
  NOR2X1   g21142(.A(new_n23578_), .B(new_n23577_), .Y(new_n23579_));
  NOR3X1   g21143(.A(new_n23575_), .B(new_n23570_), .C(pi0619), .Y(new_n23580_));
  OAI21X1  g21144(.A0(new_n23473_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n23581_));
  NOR2X1   g21145(.A(new_n23581_), .B(new_n23580_), .Y(new_n23582_));
  OAI21X1  g21146(.A0(new_n23582_), .A1(new_n23579_), .B0(pi0789), .Y(new_n23583_));
  AND2X1   g21147(.A(new_n23583_), .B(new_n23576_), .Y(new_n23584_));
  INVX1    g21148(.A(new_n23584_), .Y(new_n23585_));
  MX2X1    g21149(.A(new_n23585_), .B(new_n23473_), .S0(new_n12708_), .Y(new_n23586_));
  NAND2X1  g21150(.A(new_n23586_), .B(new_n14249_), .Y(new_n23587_));
  AND2X1   g21151(.A(pi0680), .B(pi0661), .Y(new_n23588_));
  INVX1    g21152(.A(new_n23588_), .Y(new_n23589_));
  AND3X1   g21153(.A(new_n23589_), .B(new_n12322_), .C(new_n12318_), .Y(new_n23590_));
  AOI21X1  g21154(.A0(new_n12322_), .A1(new_n12318_), .B0(pi0222), .Y(new_n23591_));
  OAI21X1  g21155(.A0(new_n12310_), .A1(new_n2941_), .B0(new_n2933_), .Y(new_n23592_));
  OR3X1    g21156(.A(new_n23592_), .B(new_n23591_), .C(new_n23590_), .Y(new_n23593_));
  AND3X1   g21157(.A(new_n23589_), .B(new_n12327_), .C(new_n12326_), .Y(new_n23594_));
  AOI21X1  g21158(.A0(new_n12327_), .A1(new_n12326_), .B0(pi0222), .Y(new_n23595_));
  OAI21X1  g21159(.A0(new_n12312_), .A1(new_n2941_), .B0(pi0299), .Y(new_n23596_));
  OR3X1    g21160(.A(new_n23596_), .B(new_n23595_), .C(new_n23594_), .Y(new_n23597_));
  AND3X1   g21161(.A(new_n23597_), .B(new_n23593_), .C(new_n2939_), .Y(new_n23598_));
  AOI22X1  g21162(.A0(new_n23260_), .A1(new_n11849_), .B0(new_n11904_), .B1(new_n11851_), .Y(new_n23599_));
  NAND2X1  g21163(.A(new_n11904_), .B(pi0681), .Y(new_n23600_));
  MX2X1    g21164(.A(new_n12814_), .B(new_n23600_), .S0(new_n11848_), .Y(new_n23601_));
  OAI21X1  g21165(.A0(new_n23599_), .A1(new_n23475_), .B0(new_n23601_), .Y(new_n23602_));
  OR2X1    g21166(.A(new_n23602_), .B(new_n5042_), .Y(new_n23603_));
  MX2X1    g21167(.A(new_n12263_), .B(new_n11926_), .S0(new_n5019_), .Y(new_n23604_));
  MX2X1    g21168(.A(new_n23604_), .B(new_n11932_), .S0(new_n11848_), .Y(new_n23605_));
  AOI21X1  g21169(.A0(new_n23605_), .A1(new_n5042_), .B0(new_n2941_), .Y(new_n23606_));
  OR3X1    g21170(.A(new_n23589_), .B(new_n12370_), .C(new_n5042_), .Y(new_n23607_));
  OR4X1    g21171(.A(new_n12275_), .B(new_n12132_), .C(new_n5041_), .D(new_n11848_), .Y(new_n23608_));
  AND3X1   g21172(.A(new_n23608_), .B(new_n23607_), .C(pi0224), .Y(new_n23609_));
  NOR4X1   g21173(.A(new_n12275_), .B(new_n11824_), .C(new_n2725_), .D(new_n11848_), .Y(new_n23610_));
  OAI21X1  g21174(.A0(new_n23610_), .A1(pi0224), .B0(new_n2941_), .Y(new_n23611_));
  OAI21X1  g21175(.A0(new_n23611_), .A1(new_n23609_), .B0(new_n2940_), .Y(new_n23612_));
  AOI21X1  g21176(.A0(new_n23606_), .A1(new_n23603_), .B0(new_n23612_), .Y(new_n23613_));
  AOI22X1  g21177(.A0(new_n12396_), .A1(new_n12280_), .B0(new_n11854_), .B1(new_n5019_), .Y(new_n23614_));
  MX2X1    g21178(.A(new_n23614_), .B(new_n11877_), .S0(new_n11848_), .Y(new_n23615_));
  NAND2X1  g21179(.A(new_n23615_), .B(new_n5041_), .Y(new_n23616_));
  NOR2X1   g21180(.A(new_n23475_), .B(new_n11858_), .Y(new_n23617_));
  OR2X1    g21181(.A(new_n12418_), .B(new_n12107_), .Y(new_n23618_));
  MX2X1    g21182(.A(new_n23618_), .B(new_n11847_), .S0(new_n11848_), .Y(new_n23619_));
  OR3X1    g21183(.A(new_n23619_), .B(new_n23617_), .C(new_n5041_), .Y(new_n23620_));
  AND3X1   g21184(.A(new_n23620_), .B(new_n23616_), .C(pi0222), .Y(new_n23621_));
  OR2X1    g21185(.A(new_n11848_), .B(pi0222), .Y(new_n23622_));
  OAI21X1  g21186(.A0(new_n23622_), .A1(new_n12382_), .B0(pi0223), .Y(new_n23623_));
  NOR2X1   g21187(.A(new_n23623_), .B(new_n23621_), .Y(new_n23624_));
  OAI21X1  g21188(.A0(new_n23624_), .A1(new_n23613_), .B0(new_n2933_), .Y(new_n23625_));
  AOI21X1  g21189(.A0(new_n23605_), .A1(new_n5059_), .B0(new_n2941_), .Y(new_n23626_));
  OAI21X1  g21190(.A0(new_n23602_), .A1(new_n5059_), .B0(new_n23626_), .Y(new_n23627_));
  AOI21X1  g21191(.A0(new_n12375_), .A1(pi0661), .B0(new_n5058_), .Y(new_n23628_));
  INVX1    g21192(.A(new_n12370_), .Y(new_n23629_));
  AOI21X1  g21193(.A0(new_n23588_), .A1(new_n23629_), .B0(new_n5059_), .Y(new_n23630_));
  OR3X1    g21194(.A(new_n23630_), .B(new_n23628_), .C(pi0222), .Y(new_n23631_));
  AND3X1   g21195(.A(new_n23631_), .B(new_n23627_), .C(new_n10045_), .Y(new_n23632_));
  INVX1    g21196(.A(new_n23510_), .Y(new_n23633_));
  OAI21X1  g21197(.A0(new_n23610_), .A1(new_n23633_), .B0(new_n2934_), .Y(new_n23634_));
  AND2X1   g21198(.A(new_n23615_), .B(new_n5058_), .Y(new_n23635_));
  NOR3X1   g21199(.A(new_n23619_), .B(new_n23617_), .C(new_n5058_), .Y(new_n23636_));
  OR3X1    g21200(.A(new_n23636_), .B(new_n23635_), .C(new_n2941_), .Y(new_n23637_));
  OAI21X1  g21201(.A0(new_n23622_), .A1(new_n12391_), .B0(new_n23637_), .Y(new_n23638_));
  AOI21X1  g21202(.A0(new_n23638_), .A1(pi0215), .B0(new_n2933_), .Y(new_n23639_));
  OAI21X1  g21203(.A0(new_n23634_), .A1(new_n23632_), .B0(new_n23639_), .Y(new_n23640_));
  AOI21X1  g21204(.A0(new_n23640_), .A1(new_n23625_), .B0(new_n2939_), .Y(new_n23641_));
  OAI21X1  g21205(.A0(new_n23641_), .A1(new_n23598_), .B0(new_n2979_), .Y(new_n23642_));
  NAND3X1  g21206(.A(new_n12439_), .B(new_n5782_), .C(pi0661), .Y(new_n23643_));
  AOI21X1  g21207(.A0(new_n23643_), .A1(new_n23556_), .B0(new_n11770_), .Y(new_n23644_));
  AOI22X1  g21208(.A0(new_n23644_), .A1(new_n23642_), .B0(new_n11770_), .B1(pi0222), .Y(new_n23645_));
  OR2X1    g21209(.A(new_n23645_), .B(pi0778), .Y(new_n23646_));
  OAI21X1  g21210(.A0(new_n23473_), .A1(pi0625), .B0(pi1153), .Y(new_n23647_));
  AOI21X1  g21211(.A0(new_n23645_), .A1(pi0625), .B0(new_n23647_), .Y(new_n23648_));
  OAI21X1  g21212(.A0(new_n23473_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n23649_));
  AOI21X1  g21213(.A0(new_n23645_), .A1(new_n12363_), .B0(new_n23649_), .Y(new_n23650_));
  OAI21X1  g21214(.A0(new_n23650_), .A1(new_n23648_), .B0(pi0778), .Y(new_n23651_));
  AND2X1   g21215(.A(new_n23651_), .B(new_n23646_), .Y(new_n23652_));
  MX2X1    g21216(.A(new_n23652_), .B(new_n23563_), .S0(new_n12490_), .Y(new_n23653_));
  MX2X1    g21217(.A(new_n23653_), .B(new_n23563_), .S0(new_n12513_), .Y(new_n23654_));
  AND2X1   g21218(.A(new_n23654_), .B(new_n14051_), .Y(new_n23655_));
  AOI22X1  g21219(.A0(new_n23655_), .A1(new_n13356_), .B0(new_n23563_), .B1(new_n21878_), .Y(new_n23656_));
  INVX1    g21220(.A(new_n16374_), .Y(new_n23657_));
  AOI21X1  g21221(.A0(new_n23563_), .A1(pi0628), .B0(new_n23657_), .Y(new_n23658_));
  OAI21X1  g21222(.A0(new_n23656_), .A1(pi0628), .B0(new_n23658_), .Y(new_n23659_));
  AOI21X1  g21223(.A0(new_n23563_), .A1(new_n12554_), .B0(new_n21973_), .Y(new_n23660_));
  OAI21X1  g21224(.A0(new_n23656_), .A1(new_n12554_), .B0(new_n23660_), .Y(new_n23661_));
  NAND3X1  g21225(.A(new_n23661_), .B(new_n23659_), .C(new_n23587_), .Y(new_n23662_));
  OR2X1    g21226(.A(new_n23578_), .B(new_n23577_), .Y(new_n23663_));
  NOR2X1   g21227(.A(new_n23476_), .B(pi0680), .Y(new_n23664_));
  AOI22X1  g21228(.A0(new_n12123_), .A1(new_n5023_), .B0(new_n12084_), .B1(new_n11977_), .Y(new_n23665_));
  INVX1    g21229(.A(new_n23665_), .Y(new_n23666_));
  AOI22X1  g21230(.A0(new_n12126_), .A1(new_n11979_), .B0(new_n11916_), .B1(pi0603), .Y(new_n23667_));
  OAI21X1  g21231(.A0(new_n23666_), .A1(pi0603), .B0(new_n23667_), .Y(new_n23668_));
  AOI21X1  g21232(.A0(new_n11991_), .A1(new_n11925_), .B0(new_n23666_), .Y(new_n23669_));
  INVX1    g21233(.A(new_n23669_), .Y(new_n23670_));
  AOI21X1  g21234(.A0(new_n23670_), .A1(pi0642), .B0(new_n21816_), .Y(new_n23671_));
  OAI21X1  g21235(.A0(new_n23668_), .A1(pi0642), .B0(new_n23671_), .Y(new_n23672_));
  INVX1    g21236(.A(new_n23672_), .Y(new_n23673_));
  INVX1    g21237(.A(new_n12224_), .Y(new_n23674_));
  NOR2X1   g21238(.A(new_n23665_), .B(new_n23674_), .Y(new_n23675_));
  INVX1    g21239(.A(new_n23675_), .Y(new_n23676_));
  AOI21X1  g21240(.A0(new_n23676_), .A1(pi0616), .B0(new_n5019_), .Y(new_n23677_));
  OAI21X1  g21241(.A0(new_n23670_), .A1(new_n12189_), .B0(new_n23677_), .Y(new_n23678_));
  OAI21X1  g21242(.A0(new_n23678_), .A1(new_n23673_), .B0(pi0661), .Y(new_n23679_));
  NOR2X1   g21243(.A(new_n23679_), .B(new_n23664_), .Y(new_n23680_));
  AND2X1   g21244(.A(pi0681), .B(new_n11848_), .Y(new_n23681_));
  AND2X1   g21245(.A(new_n23681_), .B(new_n23476_), .Y(new_n23682_));
  NOR3X1   g21246(.A(new_n23682_), .B(new_n23680_), .C(new_n23481_), .Y(new_n23683_));
  INVX1    g21247(.A(new_n23488_), .Y(new_n23684_));
  INVX1    g21248(.A(new_n12085_), .Y(new_n23685_));
  AOI21X1  g21249(.A0(new_n23685_), .A1(new_n11901_), .B0(pi0642), .Y(new_n23686_));
  OAI21X1  g21250(.A0(new_n23686_), .A1(new_n12090_), .B0(new_n11838_), .Y(new_n23687_));
  AOI21X1  g21251(.A0(new_n23687_), .A1(new_n12089_), .B0(pi0616), .Y(new_n23688_));
  OAI21X1  g21252(.A0(new_n12268_), .A1(new_n11871_), .B0(pi0680), .Y(new_n23689_));
  OAI21X1  g21253(.A0(new_n23689_), .A1(new_n23688_), .B0(pi0661), .Y(new_n23690_));
  AOI21X1  g21254(.A0(new_n23484_), .A1(new_n5019_), .B0(new_n23690_), .Y(new_n23691_));
  INVX1    g21255(.A(new_n23681_), .Y(new_n23692_));
  NOR2X1   g21256(.A(new_n23692_), .B(new_n23484_), .Y(new_n23693_));
  NOR3X1   g21257(.A(new_n23693_), .B(new_n23691_), .C(new_n23684_), .Y(new_n23694_));
  OR2X1    g21258(.A(new_n23694_), .B(new_n5059_), .Y(new_n23695_));
  AND2X1   g21259(.A(new_n23695_), .B(pi0222), .Y(new_n23696_));
  OAI21X1  g21260(.A0(new_n23683_), .A1(new_n5058_), .B0(new_n23696_), .Y(new_n23697_));
  AND2X1   g21261(.A(new_n13155_), .B(new_n13154_), .Y(new_n23698_));
  AND2X1   g21262(.A(new_n12219_), .B(pi0616), .Y(new_n23699_));
  OR2X1    g21263(.A(new_n23699_), .B(new_n5019_), .Y(new_n23700_));
  AOI21X1  g21264(.A0(new_n23497_), .A1(new_n5019_), .B0(new_n11848_), .Y(new_n23701_));
  OAI21X1  g21265(.A0(new_n23700_), .A1(new_n23698_), .B0(new_n23701_), .Y(new_n23702_));
  INVX1    g21266(.A(new_n23477_), .Y(new_n23703_));
  OAI21X1  g21267(.A0(new_n23703_), .A1(new_n11978_), .B0(new_n23681_), .Y(new_n23704_));
  AND3X1   g21268(.A(new_n23704_), .B(new_n23702_), .C(new_n23502_), .Y(new_n23705_));
  INVX1    g21269(.A(new_n23705_), .Y(new_n23706_));
  AND2X1   g21270(.A(new_n12182_), .B(pi0680), .Y(new_n23707_));
  OAI21X1  g21271(.A0(new_n12225_), .A1(new_n11871_), .B0(new_n23707_), .Y(new_n23708_));
  AOI21X1  g21272(.A0(new_n23508_), .A1(new_n5019_), .B0(new_n11848_), .Y(new_n23709_));
  AND3X1   g21273(.A(new_n23500_), .B(new_n11991_), .C(new_n11900_), .Y(new_n23710_));
  AND2X1   g21274(.A(new_n23508_), .B(new_n11851_), .Y(new_n23711_));
  NOR3X1   g21275(.A(new_n23711_), .B(new_n23710_), .C(new_n23475_), .Y(new_n23712_));
  AOI21X1  g21276(.A0(new_n23681_), .A1(new_n23509_), .B0(new_n23712_), .Y(new_n23713_));
  INVX1    g21277(.A(new_n23713_), .Y(new_n23714_));
  AOI21X1  g21278(.A0(new_n23709_), .A1(new_n23708_), .B0(new_n23714_), .Y(new_n23715_));
  AOI21X1  g21279(.A0(new_n23715_), .A1(new_n5058_), .B0(pi0222), .Y(new_n23716_));
  OAI21X1  g21280(.A0(new_n23706_), .A1(new_n5058_), .B0(new_n23716_), .Y(new_n23717_));
  AOI21X1  g21281(.A0(new_n23717_), .A1(new_n23697_), .B0(new_n10044_), .Y(new_n23718_));
  OR2X1    g21282(.A(new_n23588_), .B(new_n23477_), .Y(new_n23719_));
  MX2X1    g21283(.A(new_n12225_), .B(new_n12174_), .S0(new_n11871_), .Y(new_n23720_));
  AND2X1   g21284(.A(new_n23720_), .B(new_n23719_), .Y(new_n23721_));
  OAI21X1  g21285(.A0(new_n23721_), .A1(new_n23633_), .B0(new_n2934_), .Y(new_n23722_));
  AOI21X1  g21286(.A0(new_n23524_), .A1(new_n5019_), .B0(new_n11848_), .Y(new_n23723_));
  OAI21X1  g21287(.A0(new_n23689_), .A1(new_n12102_), .B0(new_n23723_), .Y(new_n23724_));
  OR2X1    g21288(.A(new_n23692_), .B(new_n23524_), .Y(new_n23725_));
  AND3X1   g21289(.A(new_n23725_), .B(new_n23724_), .C(new_n23527_), .Y(new_n23726_));
  OAI21X1  g21290(.A0(new_n23674_), .A1(new_n12110_), .B0(pi0616), .Y(new_n23727_));
  AND2X1   g21291(.A(new_n23727_), .B(pi0680), .Y(new_n23728_));
  AOI21X1  g21292(.A0(new_n23728_), .A1(new_n12112_), .B0(new_n11848_), .Y(new_n23729_));
  OAI21X1  g21293(.A0(new_n23517_), .A1(pi0680), .B0(new_n23729_), .Y(new_n23730_));
  AOI22X1  g21294(.A0(new_n23681_), .A1(new_n23517_), .B0(new_n23519_), .B1(new_n23230_), .Y(new_n23731_));
  AND2X1   g21295(.A(new_n23731_), .B(new_n23730_), .Y(new_n23732_));
  INVX1    g21296(.A(new_n23732_), .Y(new_n23733_));
  AOI21X1  g21297(.A0(new_n23733_), .A1(new_n5059_), .B0(new_n2941_), .Y(new_n23734_));
  OAI21X1  g21298(.A0(new_n23726_), .A1(new_n5059_), .B0(new_n23734_), .Y(new_n23735_));
  AOI21X1  g21299(.A0(new_n12177_), .A1(new_n12050_), .B0(new_n11836_), .Y(new_n23736_));
  OR2X1    g21300(.A(new_n23736_), .B(new_n11871_), .Y(new_n23737_));
  NAND4X1  g21301(.A(new_n23737_), .B(new_n12193_), .C(new_n12190_), .D(pi0680), .Y(new_n23738_));
  NOR3X1   g21302(.A(new_n12050_), .B(new_n11836_), .C(new_n11871_), .Y(new_n23739_));
  AOI21X1  g21303(.A0(new_n23739_), .A1(new_n5019_), .B0(new_n11848_), .Y(new_n23740_));
  OAI21X1  g21304(.A0(new_n23509_), .A1(new_n11835_), .B0(new_n5020_), .Y(new_n23741_));
  OAI21X1  g21305(.A0(new_n23739_), .A1(pi0661), .B0(new_n23741_), .Y(new_n23742_));
  AOI21X1  g21306(.A0(new_n23740_), .A1(new_n23738_), .B0(new_n23742_), .Y(new_n23743_));
  OR3X1    g21307(.A(new_n23589_), .B(new_n12084_), .C(new_n12015_), .Y(new_n23744_));
  AND2X1   g21308(.A(new_n23744_), .B(new_n23514_), .Y(new_n23745_));
  OAI21X1  g21309(.A0(new_n23745_), .A1(new_n5059_), .B0(new_n2941_), .Y(new_n23746_));
  AOI21X1  g21310(.A0(new_n23743_), .A1(new_n5059_), .B0(new_n23746_), .Y(new_n23747_));
  NOR2X1   g21311(.A(new_n23747_), .B(new_n2934_), .Y(new_n23748_));
  AOI21X1  g21312(.A0(new_n23748_), .A1(new_n23735_), .B0(new_n2933_), .Y(new_n23749_));
  OAI21X1  g21313(.A0(new_n23722_), .A1(new_n23718_), .B0(new_n23749_), .Y(new_n23750_));
  OR2X1    g21314(.A(new_n23720_), .B(new_n23589_), .Y(new_n23751_));
  AOI21X1  g21315(.A0(new_n23589_), .A1(new_n23509_), .B0(pi0222), .Y(new_n23752_));
  AOI21X1  g21316(.A0(new_n23752_), .A1(new_n23751_), .B0(new_n3138_), .Y(new_n23753_));
  NAND4X1  g21317(.A(new_n23704_), .B(new_n23702_), .C(new_n23502_), .D(new_n5042_), .Y(new_n23754_));
  AOI21X1  g21318(.A0(new_n23715_), .A1(new_n5041_), .B0(new_n2942_), .Y(new_n23755_));
  AOI21X1  g21319(.A0(new_n23755_), .A1(new_n23754_), .B0(new_n23753_), .Y(new_n23756_));
  NOR4X1   g21320(.A(new_n23682_), .B(new_n23680_), .C(new_n23481_), .D(new_n5041_), .Y(new_n23757_));
  NOR4X1   g21321(.A(new_n23693_), .B(new_n23691_), .C(new_n23684_), .D(new_n5042_), .Y(new_n23758_));
  NOR3X1   g21322(.A(new_n23758_), .B(new_n23757_), .C(new_n2941_), .Y(new_n23759_));
  OAI21X1  g21323(.A0(new_n23759_), .A1(new_n23756_), .B0(new_n2940_), .Y(new_n23760_));
  AOI21X1  g21324(.A0(new_n23733_), .A1(new_n5042_), .B0(new_n2941_), .Y(new_n23761_));
  OAI21X1  g21325(.A0(new_n23726_), .A1(new_n5042_), .B0(new_n23761_), .Y(new_n23762_));
  OAI21X1  g21326(.A0(new_n23745_), .A1(new_n5042_), .B0(new_n2941_), .Y(new_n23763_));
  AOI21X1  g21327(.A0(new_n23743_), .A1(new_n5042_), .B0(new_n23763_), .Y(new_n23764_));
  NOR2X1   g21328(.A(new_n23764_), .B(new_n2940_), .Y(new_n23765_));
  AOI21X1  g21329(.A0(new_n23765_), .A1(new_n23762_), .B0(pi0299), .Y(new_n23766_));
  AOI21X1  g21330(.A0(new_n23766_), .A1(new_n23760_), .B0(new_n2939_), .Y(new_n23767_));
  AND2X1   g21331(.A(new_n23767_), .B(new_n23750_), .Y(new_n23768_));
  OR2X1    g21332(.A(new_n12325_), .B(new_n11848_), .Y(new_n23769_));
  AOI21X1  g21333(.A0(new_n12041_), .A1(pi0616), .B0(pi0222), .Y(new_n23770_));
  OR3X1    g21334(.A(new_n12324_), .B(new_n12323_), .C(new_n12316_), .Y(new_n23771_));
  AND2X1   g21335(.A(new_n12310_), .B(new_n11881_), .Y(new_n23772_));
  NOR3X1   g21336(.A(new_n23772_), .B(new_n12324_), .C(new_n12126_), .Y(new_n23773_));
  AOI21X1  g21337(.A0(new_n12041_), .A1(new_n11871_), .B0(new_n23773_), .Y(new_n23774_));
  OAI21X1  g21338(.A0(new_n23588_), .A1(new_n23771_), .B0(new_n23774_), .Y(new_n23775_));
  AOI22X1  g21339(.A0(new_n23775_), .A1(pi0222), .B0(new_n23770_), .B1(new_n23769_), .Y(new_n23776_));
  OR3X1    g21340(.A(new_n23588_), .B(new_n12330_), .C(new_n12328_), .Y(new_n23777_));
  AND2X1   g21341(.A(new_n11965_), .B(pi0603), .Y(new_n23778_));
  AND2X1   g21342(.A(new_n12312_), .B(new_n11881_), .Y(new_n23779_));
  NOR3X1   g21343(.A(new_n23779_), .B(new_n12126_), .C(new_n23778_), .Y(new_n23780_));
  AOI21X1  g21344(.A0(new_n12044_), .A1(new_n11871_), .B0(new_n23780_), .Y(new_n23781_));
  AND2X1   g21345(.A(new_n23781_), .B(new_n23777_), .Y(new_n23782_));
  AOI21X1  g21346(.A0(new_n12044_), .A1(pi0616), .B0(pi0222), .Y(new_n23783_));
  OAI21X1  g21347(.A0(new_n12331_), .A1(new_n11848_), .B0(new_n23783_), .Y(new_n23784_));
  OAI21X1  g21348(.A0(new_n23782_), .A1(new_n2941_), .B0(new_n23784_), .Y(new_n23785_));
  AOI21X1  g21349(.A0(new_n23785_), .A1(pi0299), .B0(pi0039), .Y(new_n23786_));
  OAI21X1  g21350(.A0(new_n23776_), .A1(pi0299), .B0(new_n23786_), .Y(new_n23787_));
  AND2X1   g21351(.A(new_n23787_), .B(new_n2979_), .Y(new_n23788_));
  INVX1    g21352(.A(new_n23788_), .Y(new_n23789_));
  NOR4X1   g21353(.A(new_n23674_), .B(new_n2985_), .C(new_n2725_), .D(new_n2536_), .Y(new_n23790_));
  INVX1    g21354(.A(new_n23790_), .Y(new_n23791_));
  AND3X1   g21355(.A(new_n23588_), .B(pi0616), .C(new_n2939_), .Y(new_n23792_));
  AOI21X1  g21356(.A0(new_n11871_), .A1(new_n2941_), .B0(new_n23792_), .Y(new_n23793_));
  AOI22X1  g21357(.A0(new_n23589_), .A1(new_n23703_), .B0(new_n12352_), .B1(new_n11871_), .Y(new_n23794_));
  MX2X1    g21358(.A(pi0222), .B(new_n23794_), .S0(new_n12077_), .Y(new_n23795_));
  OAI21X1  g21359(.A0(new_n23793_), .A1(new_n23791_), .B0(new_n23795_), .Y(new_n23796_));
  AOI21X1  g21360(.A0(new_n23796_), .A1(pi0038), .B0(new_n11770_), .Y(new_n23797_));
  OAI21X1  g21361(.A0(new_n23789_), .A1(new_n23768_), .B0(new_n23797_), .Y(new_n23798_));
  AND2X1   g21362(.A(new_n23798_), .B(new_n23474_), .Y(new_n23799_));
  INVX1    g21363(.A(new_n23799_), .Y(new_n23800_));
  INVX1    g21364(.A(new_n23561_), .Y(new_n23801_));
  AOI21X1  g21365(.A0(new_n23801_), .A1(pi0625), .B0(pi1153), .Y(new_n23802_));
  OAI21X1  g21366(.A0(new_n23800_), .A1(pi0625), .B0(new_n23802_), .Y(new_n23803_));
  NOR2X1   g21367(.A(new_n23648_), .B(pi0608), .Y(new_n23804_));
  AOI21X1  g21368(.A0(new_n23801_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n23805_));
  OAI21X1  g21369(.A0(new_n23800_), .A1(new_n12363_), .B0(new_n23805_), .Y(new_n23806_));
  NOR2X1   g21370(.A(new_n23650_), .B(new_n12368_), .Y(new_n23807_));
  AOI22X1  g21371(.A0(new_n23807_), .A1(new_n23806_), .B0(new_n23804_), .B1(new_n23803_), .Y(new_n23808_));
  MX2X1    g21372(.A(new_n23808_), .B(new_n23800_), .S0(new_n11769_), .Y(new_n23809_));
  AOI21X1  g21373(.A0(new_n23652_), .A1(pi0609), .B0(pi1155), .Y(new_n23810_));
  OAI21X1  g21374(.A0(new_n23809_), .A1(pi0609), .B0(new_n23810_), .Y(new_n23811_));
  AND2X1   g21375(.A(new_n23565_), .B(new_n12468_), .Y(new_n23812_));
  AOI21X1  g21376(.A0(new_n23652_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n23813_));
  OAI21X1  g21377(.A0(new_n23809_), .A1(new_n12462_), .B0(new_n23813_), .Y(new_n23814_));
  AND2X1   g21378(.A(new_n23567_), .B(pi0660), .Y(new_n23815_));
  AOI22X1  g21379(.A0(new_n23815_), .A1(new_n23814_), .B0(new_n23812_), .B1(new_n23811_), .Y(new_n23816_));
  MX2X1    g21380(.A(new_n23816_), .B(new_n23809_), .S0(new_n11768_), .Y(new_n23817_));
  AOI21X1  g21381(.A0(new_n23653_), .A1(pi0618), .B0(pi1154), .Y(new_n23818_));
  OAI21X1  g21382(.A0(new_n23817_), .A1(pi0618), .B0(new_n23818_), .Y(new_n23819_));
  AND2X1   g21383(.A(new_n23572_), .B(new_n12494_), .Y(new_n23820_));
  AOI21X1  g21384(.A0(new_n23653_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n23821_));
  OAI21X1  g21385(.A0(new_n23817_), .A1(new_n12486_), .B0(new_n23821_), .Y(new_n23822_));
  AND2X1   g21386(.A(new_n23574_), .B(pi0627), .Y(new_n23823_));
  AOI22X1  g21387(.A0(new_n23823_), .A1(new_n23822_), .B0(new_n23820_), .B1(new_n23819_), .Y(new_n23824_));
  MX2X1    g21388(.A(new_n23824_), .B(new_n23817_), .S0(new_n11767_), .Y(new_n23825_));
  AOI21X1  g21389(.A0(new_n23654_), .A1(pi0619), .B0(pi1159), .Y(new_n23826_));
  OAI21X1  g21390(.A0(new_n23825_), .A1(pi0619), .B0(new_n23826_), .Y(new_n23827_));
  AND3X1   g21391(.A(new_n23827_), .B(new_n23663_), .C(new_n12517_), .Y(new_n23828_));
  OR2X1    g21392(.A(new_n23825_), .B(new_n12509_), .Y(new_n23829_));
  AOI21X1  g21393(.A0(new_n23654_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n23830_));
  OAI21X1  g21394(.A0(new_n23581_), .A1(new_n23580_), .B0(pi0648), .Y(new_n23831_));
  AOI21X1  g21395(.A0(new_n23830_), .A1(new_n23829_), .B0(new_n23831_), .Y(new_n23832_));
  NOR3X1   g21396(.A(new_n23832_), .B(new_n23828_), .C(new_n11766_), .Y(new_n23833_));
  NAND2X1  g21397(.A(new_n23825_), .B(new_n11766_), .Y(new_n23834_));
  AOI21X1  g21398(.A0(new_n23563_), .A1(pi0626), .B0(new_n16218_), .Y(new_n23835_));
  OAI21X1  g21399(.A0(new_n23585_), .A1(pi0626), .B0(new_n23835_), .Y(new_n23836_));
  AOI21X1  g21400(.A0(new_n23563_), .A1(new_n12542_), .B0(new_n16222_), .Y(new_n23837_));
  OAI21X1  g21401(.A0(new_n23585_), .A1(new_n12542_), .B0(new_n23837_), .Y(new_n23838_));
  OAI21X1  g21402(.A0(new_n23473_), .A1(new_n14051_), .B0(new_n12637_), .Y(new_n23839_));
  OR2X1    g21403(.A(new_n23839_), .B(new_n23655_), .Y(new_n23840_));
  AND3X1   g21404(.A(new_n23840_), .B(new_n23838_), .C(new_n23836_), .Y(new_n23841_));
  OAI21X1  g21405(.A0(new_n23841_), .A1(new_n11765_), .B0(new_n23834_), .Y(new_n23842_));
  OR2X1    g21406(.A(new_n23842_), .B(new_n23833_), .Y(new_n23843_));
  AOI21X1  g21407(.A0(new_n23841_), .A1(new_n13481_), .B0(new_n14125_), .Y(new_n23844_));
  AOI22X1  g21408(.A0(new_n23844_), .A1(new_n23843_), .B0(new_n23662_), .B1(pi0792), .Y(new_n23845_));
  MX2X1    g21409(.A(new_n23586_), .B(new_n23473_), .S0(new_n12580_), .Y(new_n23846_));
  OAI22X1  g21410(.A0(new_n23656_), .A1(new_n13508_), .B0(new_n23473_), .B1(new_n22699_), .Y(new_n23847_));
  OAI21X1  g21411(.A0(new_n23473_), .A1(pi0647), .B0(pi1157), .Y(new_n23848_));
  AOI21X1  g21412(.A0(new_n23847_), .A1(pi0647), .B0(new_n23848_), .Y(new_n23849_));
  OAI21X1  g21413(.A0(new_n23473_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n23850_));
  AOI21X1  g21414(.A0(new_n23847_), .A1(new_n12577_), .B0(new_n23850_), .Y(new_n23851_));
  MX2X1    g21415(.A(new_n23851_), .B(new_n23849_), .S0(new_n12592_), .Y(new_n23852_));
  AOI21X1  g21416(.A0(new_n23846_), .A1(new_n14326_), .B0(new_n23852_), .Y(new_n23853_));
  OAI22X1  g21417(.A0(new_n23853_), .A1(new_n11763_), .B0(new_n23845_), .B1(new_n14121_), .Y(new_n23854_));
  NOR2X1   g21418(.A(new_n23851_), .B(new_n23849_), .Y(new_n23855_));
  MX2X1    g21419(.A(new_n23855_), .B(new_n23847_), .S0(new_n11763_), .Y(new_n23856_));
  AOI21X1  g21420(.A0(new_n23856_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n23857_));
  OAI21X1  g21421(.A0(new_n23854_), .A1(new_n12612_), .B0(new_n23857_), .Y(new_n23858_));
  MX2X1    g21422(.A(new_n23846_), .B(new_n23473_), .S0(new_n12604_), .Y(new_n23859_));
  AOI21X1  g21423(.A0(new_n23563_), .A1(new_n12612_), .B0(pi0715), .Y(new_n23860_));
  OAI21X1  g21424(.A0(new_n23859_), .A1(new_n12612_), .B0(new_n23860_), .Y(new_n23861_));
  AND2X1   g21425(.A(new_n23861_), .B(pi1160), .Y(new_n23862_));
  AOI21X1  g21426(.A0(new_n23856_), .A1(pi0644), .B0(pi0715), .Y(new_n23863_));
  OAI21X1  g21427(.A0(new_n23854_), .A1(pi0644), .B0(new_n23863_), .Y(new_n23864_));
  AOI21X1  g21428(.A0(new_n23563_), .A1(pi0644), .B0(new_n12608_), .Y(new_n23865_));
  OAI21X1  g21429(.A0(new_n23859_), .A1(pi0644), .B0(new_n23865_), .Y(new_n23866_));
  AND2X1   g21430(.A(new_n23866_), .B(new_n11762_), .Y(new_n23867_));
  AOI22X1  g21431(.A0(new_n23867_), .A1(new_n23864_), .B0(new_n23862_), .B1(new_n23858_), .Y(new_n23868_));
  MX2X1    g21432(.A(new_n23868_), .B(new_n23854_), .S0(new_n12766_), .Y(new_n23869_));
  MX2X1    g21433(.A(new_n23869_), .B(pi0222), .S0(po1038), .Y(po0379));
  AOI21X1  g21434(.A0(new_n23250_), .A1(new_n2933_), .B0(new_n2939_), .Y(new_n23871_));
  AND2X1   g21435(.A(new_n23871_), .B(new_n11957_), .Y(new_n23872_));
  NOR3X1   g21436(.A(new_n23872_), .B(new_n12779_), .C(new_n10655_), .Y(new_n23873_));
  OAI21X1  g21437(.A0(new_n23873_), .A1(new_n21749_), .B0(pi0223), .Y(new_n23874_));
  INVX1    g21438(.A(new_n23874_), .Y(new_n23875_));
  NOR3X1   g21439(.A(new_n11979_), .B(new_n5016_), .C(new_n11881_), .Y(new_n23876_));
  NOR4X1   g21440(.A(new_n23876_), .B(new_n11824_), .C(new_n5017_), .D(new_n2725_), .Y(new_n23877_));
  INVX1    g21441(.A(new_n23877_), .Y(new_n23878_));
  NOR2X1   g21442(.A(new_n11992_), .B(new_n5016_), .Y(new_n23879_));
  NOR2X1   g21443(.A(new_n23879_), .B(new_n21816_), .Y(new_n23880_));
  OAI21X1  g21444(.A0(new_n11901_), .A1(pi0642), .B0(new_n23880_), .Y(new_n23881_));
  AND3X1   g21445(.A(new_n23881_), .B(new_n23878_), .C(pi0681), .Y(new_n23882_));
  AOI21X1  g21446(.A0(new_n23881_), .A1(new_n23878_), .B0(new_n11928_), .Y(new_n23883_));
  OAI21X1  g21447(.A0(new_n11997_), .A1(new_n5016_), .B0(new_n11900_), .Y(new_n23884_));
  OAI21X1  g21448(.A0(new_n23884_), .A1(new_n11929_), .B0(new_n11859_), .Y(new_n23885_));
  OAI21X1  g21449(.A0(new_n23885_), .A1(new_n23883_), .B0(new_n5058_), .Y(new_n23886_));
  NOR2X1   g21450(.A(new_n23886_), .B(new_n23882_), .Y(new_n23887_));
  MX2X1    g21451(.A(new_n11985_), .B(new_n11926_), .S0(new_n5016_), .Y(new_n23888_));
  NOR2X1   g21452(.A(new_n23888_), .B(new_n11859_), .Y(new_n23889_));
  AND2X1   g21453(.A(new_n23888_), .B(new_n11929_), .Y(new_n23890_));
  NOR3X1   g21454(.A(new_n23876_), .B(new_n11916_), .C(new_n11929_), .Y(new_n23891_));
  NOR3X1   g21455(.A(new_n23891_), .B(new_n23890_), .C(pi0681), .Y(new_n23892_));
  NOR3X1   g21456(.A(new_n23892_), .B(new_n23889_), .C(new_n5058_), .Y(new_n23893_));
  OR3X1    g21457(.A(new_n23893_), .B(new_n23887_), .C(new_n2940_), .Y(new_n23894_));
  NOR4X1   g21458(.A(new_n12048_), .B(new_n11824_), .C(new_n2725_), .D(new_n5016_), .Y(new_n23895_));
  INVX1    g21459(.A(new_n23895_), .Y(new_n23896_));
  AOI21X1  g21460(.A0(new_n23895_), .A1(new_n11929_), .B0(pi0681), .Y(new_n23897_));
  INVX1    g21461(.A(new_n23897_), .Y(new_n23898_));
  NOR4X1   g21462(.A(new_n5019_), .B(pi0662), .C(pi0661), .D(new_n5016_), .Y(new_n23899_));
  AND3X1   g21463(.A(new_n23899_), .B(new_n11991_), .C(new_n11900_), .Y(new_n23900_));
  OR2X1    g21464(.A(new_n23900_), .B(new_n23898_), .Y(new_n23901_));
  INVX1    g21465(.A(new_n23901_), .Y(new_n23902_));
  AOI21X1  g21466(.A0(new_n23896_), .A1(pi0681), .B0(new_n23902_), .Y(new_n23903_));
  NAND2X1  g21467(.A(new_n23903_), .B(new_n14456_), .Y(new_n23904_));
  AND2X1   g21468(.A(new_n23876_), .B(new_n11925_), .Y(new_n23905_));
  INVX1    g21469(.A(new_n23905_), .Y(new_n23906_));
  AOI21X1  g21470(.A0(new_n23899_), .A1(new_n23499_), .B0(pi0681), .Y(new_n23907_));
  OAI21X1  g21471(.A0(new_n23906_), .A1(new_n11928_), .B0(new_n23907_), .Y(new_n23908_));
  INVX1    g21472(.A(new_n23908_), .Y(new_n23909_));
  AOI21X1  g21473(.A0(new_n23906_), .A1(pi0681), .B0(new_n23909_), .Y(new_n23910_));
  AOI21X1  g21474(.A0(new_n23910_), .A1(new_n14458_), .B0(pi0947), .Y(new_n23911_));
  NAND2X1  g21475(.A(new_n23911_), .B(new_n23904_), .Y(new_n23912_));
  OR2X1    g21476(.A(new_n23910_), .B(new_n5362_), .Y(new_n23913_));
  AND2X1   g21477(.A(new_n23913_), .B(new_n2940_), .Y(new_n23914_));
  AOI21X1  g21478(.A0(new_n23914_), .A1(new_n23912_), .B0(new_n10044_), .Y(new_n23915_));
  AOI21X1  g21479(.A0(new_n11825_), .A1(pi0223), .B0(new_n10045_), .Y(new_n23916_));
  AOI21X1  g21480(.A0(new_n23916_), .A1(new_n23896_), .B0(pi0215), .Y(new_n23917_));
  INVX1    g21481(.A(new_n23917_), .Y(new_n23918_));
  AOI21X1  g21482(.A0(new_n23915_), .A1(new_n23894_), .B0(new_n23918_), .Y(new_n23919_));
  AOI21X1  g21483(.A0(new_n23899_), .A1(new_n12060_), .B0(new_n23898_), .Y(new_n23920_));
  AOI21X1  g21484(.A0(new_n12019_), .A1(pi0642), .B0(new_n11929_), .Y(new_n23921_));
  AOI21X1  g21485(.A0(new_n23921_), .A1(new_n12195_), .B0(pi0681), .Y(new_n23922_));
  AOI21X1  g21486(.A0(new_n23922_), .A1(new_n11836_), .B0(new_n23920_), .Y(new_n23923_));
  OR2X1    g21487(.A(new_n12050_), .B(new_n11836_), .Y(new_n23924_));
  OAI21X1  g21488(.A0(new_n23924_), .A1(new_n5016_), .B0(pi0681), .Y(new_n23925_));
  AND2X1   g21489(.A(new_n23925_), .B(new_n23923_), .Y(new_n23926_));
  INVX1    g21490(.A(new_n23926_), .Y(new_n23927_));
  NOR2X1   g21491(.A(new_n23920_), .B(new_n5059_), .Y(new_n23928_));
  AOI21X1  g21492(.A0(new_n23928_), .A1(new_n23895_), .B0(pi0947), .Y(new_n23929_));
  OAI21X1  g21493(.A0(new_n23927_), .A1(new_n14456_), .B0(new_n23929_), .Y(new_n23930_));
  AOI21X1  g21494(.A0(new_n23927_), .A1(pi0947), .B0(pi0223), .Y(new_n23931_));
  OAI21X1  g21495(.A0(new_n23879_), .A1(new_n23525_), .B0(new_n23878_), .Y(new_n23932_));
  INVX1    g21496(.A(new_n23932_), .Y(new_n23933_));
  NAND2X1  g21497(.A(new_n23932_), .B(new_n11929_), .Y(new_n23934_));
  NOR4X1   g21498(.A(new_n23876_), .B(new_n2985_), .C(new_n2725_), .D(new_n2536_), .Y(new_n23935_));
  AND2X1   g21499(.A(new_n23935_), .B(new_n11928_), .Y(new_n23936_));
  AOI21X1  g21500(.A0(new_n23936_), .A1(new_n12008_), .B0(pi0681), .Y(new_n23937_));
  AOI22X1  g21501(.A0(new_n23937_), .A1(new_n23934_), .B0(new_n23933_), .B1(pi0681), .Y(new_n23938_));
  AND2X1   g21502(.A(new_n23938_), .B(new_n5058_), .Y(new_n23939_));
  INVX1    g21503(.A(new_n23939_), .Y(new_n23940_));
  MX2X1    g21504(.A(new_n12020_), .B(new_n23229_), .S0(new_n5016_), .Y(new_n23941_));
  INVX1    g21505(.A(new_n23941_), .Y(new_n23942_));
  OAI21X1  g21506(.A0(new_n23942_), .A1(new_n11928_), .B0(new_n23922_), .Y(new_n23943_));
  INVX1    g21507(.A(new_n23943_), .Y(new_n23944_));
  AOI21X1  g21508(.A0(new_n23942_), .A1(pi0681), .B0(new_n23944_), .Y(new_n23945_));
  AOI21X1  g21509(.A0(new_n23945_), .A1(new_n5059_), .B0(new_n2940_), .Y(new_n23946_));
  AOI22X1  g21510(.A0(new_n23946_), .A1(new_n23940_), .B0(new_n23931_), .B1(new_n23930_), .Y(new_n23947_));
  OAI21X1  g21511(.A0(new_n23947_), .A1(new_n2934_), .B0(pi0299), .Y(new_n23948_));
  AND2X1   g21512(.A(new_n23903_), .B(new_n5041_), .Y(new_n23949_));
  INVX1    g21513(.A(new_n23949_), .Y(new_n23950_));
  AOI21X1  g21514(.A0(new_n23910_), .A1(new_n5042_), .B0(new_n2951_), .Y(new_n23951_));
  AOI21X1  g21515(.A0(new_n23896_), .A1(new_n2951_), .B0(pi0223), .Y(new_n23952_));
  INVX1    g21516(.A(new_n23952_), .Y(new_n23953_));
  AOI21X1  g21517(.A0(new_n23951_), .A1(new_n23950_), .B0(new_n23953_), .Y(new_n23954_));
  AOI21X1  g21518(.A0(new_n23945_), .A1(new_n5042_), .B0(new_n2940_), .Y(new_n23955_));
  INVX1    g21519(.A(new_n23955_), .Y(new_n23956_));
  AOI21X1  g21520(.A0(new_n23938_), .A1(new_n5041_), .B0(new_n23956_), .Y(new_n23957_));
  NOR3X1   g21521(.A(new_n23957_), .B(new_n23954_), .C(pi0299), .Y(new_n23958_));
  NOR2X1   g21522(.A(new_n23958_), .B(new_n2939_), .Y(new_n23959_));
  OAI21X1  g21523(.A0(new_n23948_), .A1(new_n23919_), .B0(new_n23959_), .Y(new_n23960_));
  AND2X1   g21524(.A(pi0642), .B(new_n2940_), .Y(new_n23961_));
  AOI21X1  g21525(.A0(new_n23961_), .A1(new_n12041_), .B0(pi0299), .Y(new_n23962_));
  INVX1    g21526(.A(new_n23962_), .Y(new_n23963_));
  AOI21X1  g21527(.A0(new_n12041_), .A1(new_n5016_), .B0(new_n2940_), .Y(new_n23964_));
  AND3X1   g21528(.A(new_n23964_), .B(new_n11973_), .C(new_n11968_), .Y(new_n23965_));
  AOI21X1  g21529(.A0(new_n23961_), .A1(new_n12044_), .B0(new_n2933_), .Y(new_n23966_));
  NOR3X1   g21530(.A(new_n12043_), .B(new_n12042_), .C(new_n11840_), .Y(new_n23967_));
  NOR3X1   g21531(.A(new_n23967_), .B(new_n11966_), .C(new_n2940_), .Y(new_n23968_));
  INVX1    g21532(.A(new_n23968_), .Y(new_n23969_));
  AOI21X1  g21533(.A0(new_n23969_), .A1(new_n23966_), .B0(pi0039), .Y(new_n23970_));
  OAI21X1  g21534(.A0(new_n23965_), .A1(new_n23963_), .B0(new_n23970_), .Y(new_n23971_));
  NAND3X1  g21535(.A(new_n23971_), .B(new_n23960_), .C(new_n2979_), .Y(new_n23972_));
  INVX1    g21536(.A(new_n23935_), .Y(new_n23973_));
  AOI21X1  g21537(.A0(pi0223), .A1(pi0039), .B0(new_n2979_), .Y(new_n23974_));
  INVX1    g21538(.A(new_n23974_), .Y(new_n23975_));
  AOI21X1  g21539(.A0(new_n13175_), .A1(new_n2940_), .B0(pi0039), .Y(new_n23976_));
  AOI21X1  g21540(.A0(new_n23976_), .A1(new_n23973_), .B0(new_n23975_), .Y(new_n23977_));
  OR2X1    g21541(.A(new_n23977_), .B(new_n11770_), .Y(new_n23978_));
  INVX1    g21542(.A(new_n23978_), .Y(new_n23979_));
  AOI22X1  g21543(.A0(new_n23979_), .A1(new_n23972_), .B0(new_n11770_), .B1(pi0223), .Y(new_n23980_));
  MX2X1    g21544(.A(new_n23980_), .B(new_n23874_), .S0(new_n12473_), .Y(new_n23981_));
  INVX1    g21545(.A(new_n23981_), .Y(new_n23982_));
  AOI21X1  g21546(.A0(new_n23874_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n23983_));
  OAI21X1  g21547(.A0(new_n23982_), .A1(new_n12462_), .B0(new_n23983_), .Y(new_n23984_));
  AOI21X1  g21548(.A0(new_n23874_), .A1(pi0609), .B0(pi1155), .Y(new_n23985_));
  OAI21X1  g21549(.A0(new_n23982_), .A1(pi0609), .B0(new_n23985_), .Y(new_n23986_));
  NAND2X1  g21550(.A(new_n23986_), .B(new_n23984_), .Y(new_n23987_));
  MX2X1    g21551(.A(new_n23987_), .B(new_n23982_), .S0(new_n11768_), .Y(new_n23988_));
  AOI21X1  g21552(.A0(new_n23874_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n23989_));
  OAI21X1  g21553(.A0(new_n23988_), .A1(new_n12486_), .B0(new_n23989_), .Y(new_n23990_));
  AOI21X1  g21554(.A0(new_n23874_), .A1(pi0618), .B0(pi1154), .Y(new_n23991_));
  OAI21X1  g21555(.A0(new_n23988_), .A1(pi0618), .B0(new_n23991_), .Y(new_n23992_));
  AOI21X1  g21556(.A0(new_n23992_), .A1(new_n23990_), .B0(new_n11767_), .Y(new_n23993_));
  AOI21X1  g21557(.A0(new_n23988_), .A1(new_n11767_), .B0(new_n23993_), .Y(new_n23994_));
  OAI21X1  g21558(.A0(new_n23875_), .A1(pi0619), .B0(pi1159), .Y(new_n23995_));
  AOI21X1  g21559(.A0(new_n23994_), .A1(pi0619), .B0(new_n23995_), .Y(new_n23996_));
  OAI21X1  g21560(.A0(new_n23875_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n23997_));
  AOI21X1  g21561(.A0(new_n23994_), .A1(new_n12509_), .B0(new_n23997_), .Y(new_n23998_));
  OAI21X1  g21562(.A0(new_n23998_), .A1(new_n23996_), .B0(pi0789), .Y(new_n23999_));
  OAI21X1  g21563(.A0(new_n23994_), .A1(pi0789), .B0(new_n23999_), .Y(new_n24000_));
  MX2X1    g21564(.A(new_n24000_), .B(new_n23875_), .S0(new_n12708_), .Y(new_n24001_));
  MX2X1    g21565(.A(new_n24001_), .B(new_n23875_), .S0(new_n12580_), .Y(new_n24002_));
  AND2X1   g21566(.A(pi0681), .B(pi0680), .Y(new_n24003_));
  INVX1    g21567(.A(new_n24003_), .Y(new_n24004_));
  AND3X1   g21568(.A(new_n24004_), .B(new_n12322_), .C(new_n12318_), .Y(new_n24005_));
  AOI21X1  g21569(.A0(new_n12322_), .A1(new_n12318_), .B0(pi0223), .Y(new_n24006_));
  OAI21X1  g21570(.A0(new_n12310_), .A1(new_n2940_), .B0(new_n2933_), .Y(new_n24007_));
  NOR3X1   g21571(.A(new_n24007_), .B(new_n24006_), .C(new_n24005_), .Y(new_n24008_));
  AND3X1   g21572(.A(new_n24004_), .B(new_n12327_), .C(new_n12326_), .Y(new_n24009_));
  AOI21X1  g21573(.A0(new_n12327_), .A1(new_n12326_), .B0(pi0223), .Y(new_n24010_));
  OAI21X1  g21574(.A0(new_n12312_), .A1(new_n2940_), .B0(pi0299), .Y(new_n24011_));
  NOR3X1   g21575(.A(new_n24011_), .B(new_n24010_), .C(new_n24009_), .Y(new_n24012_));
  NOR3X1   g21576(.A(new_n24012_), .B(new_n24008_), .C(pi0039), .Y(new_n24013_));
  OR4X1    g21577(.A(new_n12275_), .B(new_n11824_), .C(new_n2725_), .D(new_n11859_), .Y(new_n24014_));
  AND2X1   g21578(.A(new_n24014_), .B(new_n23916_), .Y(new_n24015_));
  AND2X1   g21579(.A(new_n11942_), .B(new_n5058_), .Y(new_n24016_));
  OAI21X1  g21580(.A0(new_n12814_), .A1(new_n11859_), .B0(new_n24016_), .Y(new_n24017_));
  NOR2X1   g21581(.A(new_n23604_), .B(new_n11859_), .Y(new_n24018_));
  NOR3X1   g21582(.A(new_n24018_), .B(new_n11931_), .C(new_n5058_), .Y(new_n24019_));
  NOR2X1   g21583(.A(new_n24019_), .B(new_n2940_), .Y(new_n24020_));
  OR3X1    g21584(.A(new_n12275_), .B(new_n12132_), .C(new_n11859_), .Y(new_n24021_));
  AND2X1   g21585(.A(new_n24021_), .B(new_n5059_), .Y(new_n24022_));
  NOR2X1   g21586(.A(new_n24004_), .B(new_n12370_), .Y(new_n24023_));
  OAI21X1  g21587(.A0(new_n24023_), .A1(new_n5059_), .B0(new_n2940_), .Y(new_n24024_));
  OAI21X1  g21588(.A0(new_n24024_), .A1(new_n24022_), .B0(new_n10045_), .Y(new_n24025_));
  AOI21X1  g21589(.A0(new_n24020_), .A1(new_n24017_), .B0(new_n24025_), .Y(new_n24026_));
  OAI21X1  g21590(.A0(new_n24026_), .A1(new_n24015_), .B0(new_n2934_), .Y(new_n24027_));
  AND2X1   g21591(.A(new_n23618_), .B(pi0681), .Y(new_n24028_));
  OR3X1    g21592(.A(new_n24028_), .B(new_n11861_), .C(new_n5058_), .Y(new_n24029_));
  NOR2X1   g21593(.A(new_n23614_), .B(new_n11859_), .Y(new_n24030_));
  NOR2X1   g21594(.A(new_n24030_), .B(new_n11876_), .Y(new_n24031_));
  AOI21X1  g21595(.A0(new_n24031_), .A1(new_n5058_), .B0(new_n2940_), .Y(new_n24032_));
  AND2X1   g21596(.A(pi0681), .B(new_n2940_), .Y(new_n24033_));
  AOI21X1  g21597(.A0(new_n24033_), .A1(new_n12390_), .B0(new_n2934_), .Y(new_n24034_));
  INVX1    g21598(.A(new_n24034_), .Y(new_n24035_));
  AOI21X1  g21599(.A0(new_n24032_), .A1(new_n24029_), .B0(new_n24035_), .Y(new_n24036_));
  NOR2X1   g21600(.A(new_n24036_), .B(new_n2933_), .Y(new_n24037_));
  NAND2X1  g21601(.A(new_n24037_), .B(new_n24027_), .Y(new_n24038_));
  NOR4X1   g21602(.A(new_n12275_), .B(new_n11824_), .C(new_n2725_), .D(new_n11859_), .Y(new_n24039_));
  NOR3X1   g21603(.A(new_n24004_), .B(new_n12370_), .C(new_n5042_), .Y(new_n24040_));
  OAI21X1  g21604(.A0(new_n24021_), .A1(new_n5041_), .B0(new_n2952_), .Y(new_n24041_));
  OAI22X1  g21605(.A0(new_n24041_), .A1(new_n24040_), .B0(new_n24039_), .B1(new_n2952_), .Y(new_n24042_));
  AND2X1   g21606(.A(new_n24042_), .B(new_n2940_), .Y(new_n24043_));
  INVX1    g21607(.A(new_n24043_), .Y(new_n24044_));
  OAI21X1  g21608(.A0(new_n24028_), .A1(new_n11861_), .B0(new_n5042_), .Y(new_n24045_));
  OAI21X1  g21609(.A0(new_n24031_), .A1(new_n5042_), .B0(pi0223), .Y(new_n24046_));
  INVX1    g21610(.A(new_n24046_), .Y(new_n24047_));
  AOI21X1  g21611(.A0(new_n24047_), .A1(new_n24045_), .B0(pi0299), .Y(new_n24048_));
  AOI21X1  g21612(.A0(new_n24048_), .A1(new_n24044_), .B0(new_n2939_), .Y(new_n24049_));
  AND2X1   g21613(.A(new_n24049_), .B(new_n24038_), .Y(new_n24050_));
  OAI21X1  g21614(.A0(new_n24050_), .A1(new_n24013_), .B0(new_n2979_), .Y(new_n24051_));
  AND3X1   g21615(.A(new_n12439_), .B(new_n5782_), .C(pi0681), .Y(new_n24052_));
  INVX1    g21616(.A(new_n24052_), .Y(new_n24053_));
  AOI21X1  g21617(.A0(new_n12771_), .A1(pi0223), .B0(new_n2979_), .Y(new_n24054_));
  AOI21X1  g21618(.A0(new_n24054_), .A1(new_n24053_), .B0(new_n11770_), .Y(new_n24055_));
  AOI22X1  g21619(.A0(new_n24055_), .A1(new_n24051_), .B0(new_n11770_), .B1(pi0223), .Y(new_n24056_));
  INVX1    g21620(.A(new_n24056_), .Y(new_n24057_));
  AOI21X1  g21621(.A0(new_n23874_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n24058_));
  OAI21X1  g21622(.A0(new_n24057_), .A1(new_n12363_), .B0(new_n24058_), .Y(new_n24059_));
  AOI21X1  g21623(.A0(new_n23874_), .A1(pi0625), .B0(pi1153), .Y(new_n24060_));
  OAI21X1  g21624(.A0(new_n24057_), .A1(pi0625), .B0(new_n24060_), .Y(new_n24061_));
  AND2X1   g21625(.A(new_n24061_), .B(new_n24059_), .Y(new_n24062_));
  MX2X1    g21626(.A(new_n24062_), .B(new_n24056_), .S0(new_n11769_), .Y(new_n24063_));
  MX2X1    g21627(.A(new_n24063_), .B(new_n23874_), .S0(new_n12490_), .Y(new_n24064_));
  MX2X1    g21628(.A(new_n24064_), .B(new_n23874_), .S0(new_n12513_), .Y(new_n24065_));
  AND2X1   g21629(.A(new_n24065_), .B(new_n14051_), .Y(new_n24066_));
  AOI22X1  g21630(.A0(new_n24066_), .A1(new_n13356_), .B0(new_n23874_), .B1(new_n21878_), .Y(new_n24067_));
  OAI22X1  g21631(.A0(new_n24067_), .A1(new_n13508_), .B0(new_n23875_), .B1(new_n22699_), .Y(new_n24068_));
  OAI21X1  g21632(.A0(new_n23875_), .A1(pi0647), .B0(pi1157), .Y(new_n24069_));
  AOI21X1  g21633(.A0(new_n24068_), .A1(pi0647), .B0(new_n24069_), .Y(new_n24070_));
  OAI21X1  g21634(.A0(new_n23875_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n24071_));
  AOI21X1  g21635(.A0(new_n24068_), .A1(new_n12577_), .B0(new_n24071_), .Y(new_n24072_));
  MX2X1    g21636(.A(new_n24072_), .B(new_n24070_), .S0(new_n12592_), .Y(new_n24073_));
  AOI21X1  g21637(.A0(new_n24002_), .A1(new_n14326_), .B0(new_n24073_), .Y(new_n24074_));
  NAND2X1  g21638(.A(new_n24001_), .B(new_n14249_), .Y(new_n24075_));
  AOI21X1  g21639(.A0(new_n23874_), .A1(pi0628), .B0(new_n23657_), .Y(new_n24076_));
  OAI21X1  g21640(.A0(new_n24067_), .A1(pi0628), .B0(new_n24076_), .Y(new_n24077_));
  AOI21X1  g21641(.A0(new_n23874_), .A1(new_n12554_), .B0(new_n21973_), .Y(new_n24078_));
  OAI21X1  g21642(.A0(new_n24067_), .A1(new_n12554_), .B0(new_n24078_), .Y(new_n24079_));
  NAND3X1  g21643(.A(new_n24079_), .B(new_n24077_), .C(new_n24075_), .Y(new_n24080_));
  OAI21X1  g21644(.A0(new_n23874_), .A1(pi0626), .B0(new_n16221_), .Y(new_n24081_));
  AOI21X1  g21645(.A0(new_n24000_), .A1(pi0626), .B0(new_n24081_), .Y(new_n24082_));
  AND2X1   g21646(.A(new_n24000_), .B(new_n12542_), .Y(new_n24083_));
  OAI21X1  g21647(.A0(new_n23874_), .A1(new_n12542_), .B0(new_n16217_), .Y(new_n24084_));
  AOI21X1  g21648(.A0(new_n23874_), .A1(new_n12531_), .B0(new_n24066_), .Y(new_n24085_));
  OAI22X1  g21649(.A0(new_n24085_), .A1(new_n13439_), .B0(new_n24084_), .B1(new_n24083_), .Y(new_n24086_));
  OAI21X1  g21650(.A0(new_n24086_), .A1(new_n24082_), .B0(pi0788), .Y(new_n24087_));
  INVX1    g21651(.A(new_n23239_), .Y(new_n24088_));
  OR2X1    g21652(.A(new_n12268_), .B(new_n5016_), .Y(new_n24089_));
  AOI21X1  g21653(.A0(new_n24089_), .A1(new_n23685_), .B0(new_n24088_), .Y(new_n24090_));
  NOR2X1   g21654(.A(new_n24090_), .B(new_n5019_), .Y(new_n24091_));
  INVX1    g21655(.A(new_n24091_), .Y(new_n24092_));
  OAI21X1  g21656(.A0(new_n12225_), .A1(new_n5016_), .B0(new_n5017_), .Y(new_n24093_));
  AOI21X1  g21657(.A0(new_n12180_), .A1(new_n5016_), .B0(new_n24093_), .Y(new_n24094_));
  OAI22X1  g21658(.A0(new_n24094_), .A1(new_n24092_), .B0(new_n23895_), .B1(pi0680), .Y(new_n24095_));
  AOI21X1  g21659(.A0(new_n24095_), .A1(pi0681), .B0(new_n23902_), .Y(new_n24096_));
  OAI21X1  g21660(.A0(new_n23906_), .A1(pi0680), .B0(pi0681), .Y(new_n24097_));
  NOR2X1   g21661(.A(new_n5017_), .B(pi0642), .Y(new_n24098_));
  AOI21X1  g21662(.A0(new_n12219_), .A1(pi0642), .B0(new_n5019_), .Y(new_n24099_));
  OAI21X1  g21663(.A0(new_n13153_), .A1(new_n12001_), .B0(new_n24099_), .Y(new_n24100_));
  AOI21X1  g21664(.A0(new_n24098_), .A1(new_n12161_), .B0(new_n24100_), .Y(new_n24101_));
  OAI21X1  g21665(.A0(new_n24101_), .A1(new_n24097_), .B0(new_n23908_), .Y(new_n24102_));
  AOI21X1  g21666(.A0(new_n24102_), .A1(new_n5059_), .B0(pi0223), .Y(new_n24103_));
  OAI21X1  g21667(.A0(new_n24096_), .A1(new_n5059_), .B0(new_n24103_), .Y(new_n24104_));
  OR2X1    g21668(.A(new_n23885_), .B(new_n23883_), .Y(new_n24105_));
  MX2X1    g21669(.A(new_n23674_), .B(new_n12085_), .S0(new_n5016_), .Y(new_n24106_));
  NOR4X1   g21670(.A(new_n24106_), .B(new_n2985_), .C(new_n2725_), .D(new_n2536_), .Y(new_n24107_));
  AND2X1   g21671(.A(new_n24107_), .B(new_n12274_), .Y(new_n24108_));
  OAI21X1  g21672(.A0(new_n24108_), .A1(new_n5017_), .B0(pi0680), .Y(new_n24109_));
  AOI21X1  g21673(.A0(new_n24089_), .A1(new_n12119_), .B0(new_n21816_), .Y(new_n24110_));
  OAI22X1  g21674(.A0(new_n24110_), .A1(new_n24109_), .B0(new_n24003_), .B1(new_n23882_), .Y(new_n24111_));
  NAND3X1  g21675(.A(new_n24111_), .B(new_n24105_), .C(new_n5058_), .Y(new_n24112_));
  NOR2X1   g21676(.A(new_n23892_), .B(new_n5058_), .Y(new_n24113_));
  NAND2X1  g21677(.A(new_n23668_), .B(new_n11999_), .Y(new_n24114_));
  OAI21X1  g21678(.A0(new_n23675_), .A1(new_n5016_), .B0(pi0680), .Y(new_n24115_));
  AOI21X1  g21679(.A0(new_n24098_), .A1(new_n23669_), .B0(new_n24115_), .Y(new_n24116_));
  NAND2X1  g21680(.A(new_n24116_), .B(new_n24114_), .Y(new_n24117_));
  OAI21X1  g21681(.A0(new_n24003_), .A1(new_n23889_), .B0(new_n24117_), .Y(new_n24118_));
  AOI21X1  g21682(.A0(new_n24118_), .A1(new_n24113_), .B0(new_n2940_), .Y(new_n24119_));
  AOI21X1  g21683(.A0(new_n24119_), .A1(new_n24112_), .B0(new_n10044_), .Y(new_n24120_));
  AOI21X1  g21684(.A0(new_n23685_), .A1(new_n5016_), .B0(new_n24004_), .Y(new_n24121_));
  AOI22X1  g21685(.A0(new_n24121_), .A1(new_n23791_), .B0(new_n24004_), .B1(new_n23876_), .Y(new_n24122_));
  NOR3X1   g21686(.A(new_n24122_), .B(new_n11825_), .C(pi0223), .Y(new_n24123_));
  AOI21X1  g21687(.A0(new_n24107_), .A1(new_n24003_), .B0(new_n2940_), .Y(new_n24124_));
  OAI21X1  g21688(.A0(new_n24003_), .A1(new_n23973_), .B0(new_n24124_), .Y(new_n24125_));
  NAND2X1  g21689(.A(new_n24125_), .B(new_n23916_), .Y(new_n24126_));
  OAI21X1  g21690(.A0(new_n24126_), .A1(new_n24123_), .B0(new_n2934_), .Y(new_n24127_));
  AOI21X1  g21691(.A0(new_n24120_), .A1(new_n24104_), .B0(new_n24127_), .Y(new_n24128_));
  OAI21X1  g21692(.A0(new_n23933_), .A1(new_n11928_), .B0(new_n23937_), .Y(new_n24129_));
  OAI21X1  g21693(.A0(new_n23933_), .A1(pi0680), .B0(pi0681), .Y(new_n24130_));
  NOR2X1   g21694(.A(new_n12268_), .B(new_n5016_), .Y(new_n24131_));
  AOI21X1  g21695(.A0(new_n12100_), .A1(new_n11838_), .B0(new_n24131_), .Y(new_n24132_));
  NOR2X1   g21696(.A(new_n24132_), .B(pi0616), .Y(new_n24133_));
  NOR2X1   g21697(.A(new_n24133_), .B(new_n24109_), .Y(new_n24134_));
  OAI21X1  g21698(.A0(new_n24134_), .A1(new_n24130_), .B0(new_n24129_), .Y(new_n24135_));
  NOR2X1   g21699(.A(new_n12111_), .B(new_n5017_), .Y(new_n24136_));
  NOR2X1   g21700(.A(new_n23674_), .B(new_n12110_), .Y(new_n24137_));
  NOR2X1   g21701(.A(new_n24137_), .B(new_n5016_), .Y(new_n24138_));
  OAI21X1  g21702(.A0(new_n12097_), .A1(new_n12001_), .B0(pi0680), .Y(new_n24139_));
  NOR3X1   g21703(.A(new_n24139_), .B(new_n24138_), .C(new_n24136_), .Y(new_n24140_));
  OR2X1    g21704(.A(new_n24140_), .B(new_n11859_), .Y(new_n24141_));
  AOI21X1  g21705(.A0(new_n23941_), .A1(new_n5019_), .B0(new_n24141_), .Y(new_n24142_));
  NOR2X1   g21706(.A(new_n24142_), .B(new_n23944_), .Y(new_n24143_));
  OAI21X1  g21707(.A0(new_n24143_), .A1(new_n5058_), .B0(pi0223), .Y(new_n24144_));
  AOI21X1  g21708(.A0(new_n24135_), .A1(new_n5058_), .B0(new_n24144_), .Y(new_n24145_));
  INVX1    g21709(.A(new_n23928_), .Y(new_n24146_));
  OAI21X1  g21710(.A0(new_n24093_), .A1(new_n12192_), .B0(new_n24091_), .Y(new_n24147_));
  OAI21X1  g21711(.A0(new_n23895_), .A1(pi0680), .B0(new_n24147_), .Y(new_n24148_));
  AOI21X1  g21712(.A0(new_n24148_), .A1(pi0681), .B0(new_n24146_), .Y(new_n24149_));
  AND3X1   g21713(.A(new_n12245_), .B(new_n12179_), .C(new_n12011_), .Y(new_n24150_));
  OR2X1    g21714(.A(new_n24150_), .B(new_n12001_), .Y(new_n24151_));
  OAI21X1  g21715(.A0(new_n23736_), .A1(new_n5016_), .B0(pi0680), .Y(new_n24152_));
  AOI21X1  g21716(.A0(new_n24098_), .A1(new_n12191_), .B0(new_n24152_), .Y(new_n24153_));
  AOI22X1  g21717(.A0(new_n24153_), .A1(new_n24151_), .B0(new_n24004_), .B1(new_n23925_), .Y(new_n24154_));
  NAND2X1  g21718(.A(new_n23923_), .B(new_n5059_), .Y(new_n24155_));
  OAI21X1  g21719(.A0(new_n24155_), .A1(new_n24154_), .B0(new_n2940_), .Y(new_n24156_));
  OAI21X1  g21720(.A0(new_n24156_), .A1(new_n24149_), .B0(pi0215), .Y(new_n24157_));
  OAI21X1  g21721(.A0(new_n24157_), .A1(new_n24145_), .B0(pi0299), .Y(new_n24158_));
  NOR2X1   g21722(.A(new_n24102_), .B(new_n5041_), .Y(new_n24159_));
  AND2X1   g21723(.A(new_n24096_), .B(new_n5041_), .Y(new_n24160_));
  OR2X1    g21724(.A(new_n24160_), .B(new_n2951_), .Y(new_n24161_));
  OAI21X1  g21725(.A0(new_n24122_), .A1(new_n11825_), .B0(new_n2951_), .Y(new_n24162_));
  AND2X1   g21726(.A(new_n24162_), .B(new_n2940_), .Y(new_n24163_));
  OAI21X1  g21727(.A0(new_n24161_), .A1(new_n24159_), .B0(new_n24163_), .Y(new_n24164_));
  OR2X1    g21728(.A(new_n24135_), .B(new_n5042_), .Y(new_n24165_));
  AOI21X1  g21729(.A0(new_n24143_), .A1(new_n5042_), .B0(new_n2940_), .Y(new_n24166_));
  AOI21X1  g21730(.A0(new_n24166_), .A1(new_n24165_), .B0(pi0299), .Y(new_n24167_));
  AOI21X1  g21731(.A0(new_n24167_), .A1(new_n24164_), .B0(new_n2939_), .Y(new_n24168_));
  OAI21X1  g21732(.A0(new_n24158_), .A1(new_n24128_), .B0(new_n24168_), .Y(new_n24169_));
  INVX1    g21733(.A(new_n23773_), .Y(new_n24170_));
  OR4X1    g21734(.A(new_n24003_), .B(new_n12324_), .C(new_n12323_), .D(new_n12316_), .Y(new_n24171_));
  NAND3X1  g21735(.A(new_n24171_), .B(new_n23964_), .C(new_n24170_), .Y(new_n24172_));
  AOI21X1  g21736(.A0(new_n24033_), .A1(new_n12793_), .B0(new_n23963_), .Y(new_n24173_));
  AND2X1   g21737(.A(new_n24173_), .B(new_n24172_), .Y(new_n24174_));
  NAND2X1  g21738(.A(new_n24033_), .B(new_n12794_), .Y(new_n24175_));
  NOR3X1   g21739(.A(new_n24003_), .B(new_n12330_), .C(new_n12328_), .Y(new_n24176_));
  OR4X1    g21740(.A(new_n24176_), .B(new_n23967_), .C(new_n23780_), .D(new_n2940_), .Y(new_n24177_));
  AND3X1   g21741(.A(new_n24177_), .B(new_n24175_), .C(new_n23966_), .Y(new_n24178_));
  OR3X1    g21742(.A(new_n24178_), .B(new_n24174_), .C(pi0039), .Y(new_n24179_));
  AND3X1   g21743(.A(new_n24179_), .B(new_n24169_), .C(new_n2979_), .Y(new_n24180_));
  NAND2X1  g21744(.A(new_n24125_), .B(new_n24122_), .Y(new_n24181_));
  AOI21X1  g21745(.A0(new_n24181_), .A1(new_n23976_), .B0(new_n23975_), .Y(new_n24182_));
  OR2X1    g21746(.A(new_n24182_), .B(new_n11770_), .Y(new_n24183_));
  OAI22X1  g21747(.A0(new_n24183_), .A1(new_n24180_), .B0(new_n3103_), .B1(new_n2940_), .Y(new_n24184_));
  OR2X1    g21748(.A(new_n24184_), .B(pi0625), .Y(new_n24185_));
  AOI21X1  g21749(.A0(new_n23980_), .A1(pi0625), .B0(pi1153), .Y(new_n24186_));
  AOI21X1  g21750(.A0(new_n24186_), .A1(new_n24185_), .B0(pi0608), .Y(new_n24187_));
  OR2X1    g21751(.A(new_n24184_), .B(new_n12363_), .Y(new_n24188_));
  AOI21X1  g21752(.A0(new_n23980_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n24189_));
  AOI21X1  g21753(.A0(new_n24189_), .A1(new_n24188_), .B0(new_n12368_), .Y(new_n24190_));
  AOI22X1  g21754(.A0(new_n24190_), .A1(new_n24061_), .B0(new_n24187_), .B1(new_n24059_), .Y(new_n24191_));
  MX2X1    g21755(.A(new_n24191_), .B(new_n24184_), .S0(new_n11769_), .Y(new_n24192_));
  AOI21X1  g21756(.A0(new_n24063_), .A1(pi0609), .B0(pi1155), .Y(new_n24193_));
  OAI21X1  g21757(.A0(new_n24192_), .A1(pi0609), .B0(new_n24193_), .Y(new_n24194_));
  AND3X1   g21758(.A(new_n24194_), .B(new_n23984_), .C(new_n12468_), .Y(new_n24195_));
  AOI21X1  g21759(.A0(new_n24063_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n24196_));
  OAI21X1  g21760(.A0(new_n24192_), .A1(new_n12462_), .B0(new_n24196_), .Y(new_n24197_));
  AND3X1   g21761(.A(new_n24197_), .B(new_n23986_), .C(pi0660), .Y(new_n24198_));
  OAI21X1  g21762(.A0(new_n24198_), .A1(new_n24195_), .B0(pi0785), .Y(new_n24199_));
  OAI21X1  g21763(.A0(new_n24192_), .A1(pi0785), .B0(new_n24199_), .Y(new_n24200_));
  INVX1    g21764(.A(new_n24064_), .Y(new_n24201_));
  OAI21X1  g21765(.A0(new_n24201_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n24202_));
  AOI21X1  g21766(.A0(new_n24200_), .A1(new_n12486_), .B0(new_n24202_), .Y(new_n24203_));
  NAND2X1  g21767(.A(new_n23990_), .B(new_n12494_), .Y(new_n24204_));
  OAI21X1  g21768(.A0(new_n24201_), .A1(pi0618), .B0(pi1154), .Y(new_n24205_));
  AOI21X1  g21769(.A0(new_n24200_), .A1(pi0618), .B0(new_n24205_), .Y(new_n24206_));
  NAND2X1  g21770(.A(new_n23992_), .B(pi0627), .Y(new_n24207_));
  OAI22X1  g21771(.A0(new_n24207_), .A1(new_n24206_), .B0(new_n24204_), .B1(new_n24203_), .Y(new_n24208_));
  MX2X1    g21772(.A(new_n24208_), .B(new_n24200_), .S0(new_n11767_), .Y(new_n24209_));
  NAND2X1  g21773(.A(new_n24209_), .B(new_n12509_), .Y(new_n24210_));
  AOI21X1  g21774(.A0(new_n24065_), .A1(pi0619), .B0(pi1159), .Y(new_n24211_));
  OR2X1    g21775(.A(new_n23996_), .B(pi0648), .Y(new_n24212_));
  AOI21X1  g21776(.A0(new_n24211_), .A1(new_n24210_), .B0(new_n24212_), .Y(new_n24213_));
  AND2X1   g21777(.A(new_n24065_), .B(new_n12509_), .Y(new_n24214_));
  OR2X1    g21778(.A(new_n24214_), .B(new_n12510_), .Y(new_n24215_));
  AOI21X1  g21779(.A0(new_n24209_), .A1(pi0619), .B0(new_n24215_), .Y(new_n24216_));
  OR2X1    g21780(.A(new_n23998_), .B(new_n12517_), .Y(new_n24217_));
  OAI21X1  g21781(.A0(new_n24217_), .A1(new_n24216_), .B0(pi0789), .Y(new_n24218_));
  OR2X1    g21782(.A(new_n24209_), .B(pi0789), .Y(new_n24219_));
  AND2X1   g21783(.A(new_n24219_), .B(new_n12709_), .Y(new_n24220_));
  OAI21X1  g21784(.A0(new_n24218_), .A1(new_n24213_), .B0(new_n24220_), .Y(new_n24221_));
  AOI22X1  g21785(.A0(new_n24221_), .A1(new_n24087_), .B0(new_n24080_), .B1(pi0792), .Y(new_n24222_));
  OAI21X1  g21786(.A0(new_n24080_), .A1(new_n14126_), .B0(new_n14122_), .Y(new_n24223_));
  OAI22X1  g21787(.A0(new_n24223_), .A1(new_n24222_), .B0(new_n24074_), .B1(new_n11763_), .Y(new_n24224_));
  NOR2X1   g21788(.A(new_n24072_), .B(new_n24070_), .Y(new_n24225_));
  MX2X1    g21789(.A(new_n24225_), .B(new_n24068_), .S0(new_n11763_), .Y(new_n24226_));
  AOI21X1  g21790(.A0(new_n24226_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n24227_));
  OAI21X1  g21791(.A0(new_n24224_), .A1(new_n12612_), .B0(new_n24227_), .Y(new_n24228_));
  MX2X1    g21792(.A(new_n24002_), .B(new_n23875_), .S0(new_n12604_), .Y(new_n24229_));
  AOI21X1  g21793(.A0(new_n23874_), .A1(new_n12612_), .B0(pi0715), .Y(new_n24230_));
  OAI21X1  g21794(.A0(new_n24229_), .A1(new_n12612_), .B0(new_n24230_), .Y(new_n24231_));
  AND2X1   g21795(.A(new_n24231_), .B(pi1160), .Y(new_n24232_));
  AOI21X1  g21796(.A0(new_n24226_), .A1(pi0644), .B0(pi0715), .Y(new_n24233_));
  OAI21X1  g21797(.A0(new_n24224_), .A1(pi0644), .B0(new_n24233_), .Y(new_n24234_));
  AOI21X1  g21798(.A0(new_n23874_), .A1(pi0644), .B0(new_n12608_), .Y(new_n24235_));
  OAI21X1  g21799(.A0(new_n24229_), .A1(pi0644), .B0(new_n24235_), .Y(new_n24236_));
  AND2X1   g21800(.A(new_n24236_), .B(new_n11762_), .Y(new_n24237_));
  AOI22X1  g21801(.A0(new_n24237_), .A1(new_n24234_), .B0(new_n24232_), .B1(new_n24228_), .Y(new_n24238_));
  MX2X1    g21802(.A(new_n24238_), .B(new_n24224_), .S0(new_n12766_), .Y(new_n24239_));
  MX2X1    g21803(.A(new_n24239_), .B(pi0223), .S0(po1038), .Y(po0380));
  NOR2X1   g21804(.A(new_n23472_), .B(new_n2942_), .Y(new_n24241_));
  NOR3X1   g21805(.A(new_n11979_), .B(new_n11838_), .C(new_n11881_), .Y(new_n24242_));
  OR3X1    g21806(.A(new_n24242_), .B(new_n11824_), .C(new_n2725_), .Y(new_n24243_));
  AND2X1   g21807(.A(new_n24243_), .B(new_n5348_), .Y(new_n24244_));
  AOI21X1  g21808(.A0(new_n11903_), .A1(new_n11871_), .B0(new_n24244_), .Y(new_n24245_));
  NOR2X1   g21809(.A(new_n24245_), .B(new_n11863_), .Y(new_n24246_));
  OAI21X1  g21810(.A0(new_n24242_), .A1(new_n11917_), .B0(pi0680), .Y(new_n24247_));
  OAI21X1  g21811(.A0(new_n24245_), .A1(pi0680), .B0(new_n24247_), .Y(new_n24248_));
  AOI21X1  g21812(.A0(new_n24248_), .A1(new_n11863_), .B0(new_n24246_), .Y(new_n24249_));
  NAND2X1  g21813(.A(new_n24249_), .B(new_n5058_), .Y(new_n24250_));
  AOI21X1  g21814(.A0(new_n11899_), .A1(new_n5023_), .B0(new_n21816_), .Y(new_n24251_));
  OAI21X1  g21815(.A0(new_n11902_), .A1(new_n5023_), .B0(new_n24251_), .Y(new_n24252_));
  AND2X1   g21816(.A(pi0616), .B(new_n11838_), .Y(new_n24253_));
  AOI22X1  g21817(.A0(new_n24253_), .A1(new_n11978_), .B0(new_n12156_), .B1(pi0614), .Y(new_n24254_));
  AOI21X1  g21818(.A0(new_n24254_), .A1(new_n24252_), .B0(new_n11863_), .Y(new_n24255_));
  AND2X1   g21819(.A(new_n24254_), .B(new_n24252_), .Y(new_n24256_));
  AOI21X1  g21820(.A0(new_n23499_), .A1(pi0614), .B0(new_n5019_), .Y(new_n24257_));
  AOI22X1  g21821(.A0(new_n24257_), .A1(new_n11916_), .B0(new_n24242_), .B1(pi0680), .Y(new_n24258_));
  OAI21X1  g21822(.A0(new_n24256_), .A1(pi0680), .B0(new_n24258_), .Y(new_n24259_));
  AOI21X1  g21823(.A0(new_n24259_), .A1(new_n11863_), .B0(new_n24255_), .Y(new_n24260_));
  AOI21X1  g21824(.A0(new_n24260_), .A1(new_n5059_), .B0(new_n2942_), .Y(new_n24261_));
  AND2X1   g21825(.A(new_n24242_), .B(new_n11925_), .Y(new_n24262_));
  AOI21X1  g21826(.A0(new_n24242_), .A1(new_n11925_), .B0(pi0680), .Y(new_n24263_));
  OAI21X1  g21827(.A0(new_n24263_), .A1(new_n24257_), .B0(new_n11863_), .Y(new_n24264_));
  OAI21X1  g21828(.A0(new_n24262_), .A1(new_n11863_), .B0(new_n24264_), .Y(new_n24265_));
  NOR2X1   g21829(.A(new_n23493_), .B(new_n11838_), .Y(new_n24266_));
  OAI21X1  g21830(.A0(new_n24266_), .A1(new_n5059_), .B0(new_n2942_), .Y(new_n24267_));
  AOI21X1  g21831(.A0(new_n24265_), .A1(new_n5059_), .B0(new_n24267_), .Y(new_n24268_));
  OR2X1    g21832(.A(new_n24268_), .B(new_n10044_), .Y(new_n24269_));
  AOI21X1  g21833(.A0(new_n24261_), .A1(new_n24250_), .B0(new_n24269_), .Y(new_n24270_));
  AOI21X1  g21834(.A0(new_n11825_), .A1(pi0224), .B0(new_n10045_), .Y(new_n24271_));
  INVX1    g21835(.A(new_n24271_), .Y(new_n24272_));
  NOR4X1   g21836(.A(new_n12048_), .B(new_n11824_), .C(new_n2725_), .D(new_n11838_), .Y(new_n24273_));
  OAI21X1  g21837(.A0(new_n24273_), .A1(new_n24272_), .B0(new_n2934_), .Y(new_n24274_));
  OR3X1    g21838(.A(new_n23513_), .B(new_n11838_), .C(pi0224), .Y(new_n24275_));
  NOR2X1   g21839(.A(new_n24244_), .B(new_n11866_), .Y(new_n24276_));
  INVX1    g21840(.A(new_n24276_), .Y(new_n24277_));
  OAI21X1  g21841(.A0(new_n24244_), .A1(new_n11866_), .B0(new_n5019_), .Y(new_n24278_));
  AOI21X1  g21842(.A0(new_n24242_), .A1(pi0680), .B0(new_n11868_), .Y(new_n24279_));
  AOI21X1  g21843(.A0(new_n24279_), .A1(new_n24278_), .B0(new_n11867_), .Y(new_n24280_));
  AOI21X1  g21844(.A0(new_n24277_), .A1(new_n11867_), .B0(new_n24280_), .Y(new_n24281_));
  AND2X1   g21845(.A(new_n24281_), .B(new_n5058_), .Y(new_n24282_));
  OAI21X1  g21846(.A0(new_n12020_), .A1(new_n11838_), .B0(new_n23311_), .Y(new_n24283_));
  NAND2X1  g21847(.A(new_n24283_), .B(new_n5019_), .Y(new_n24284_));
  NAND2X1  g21848(.A(new_n12022_), .B(pi0680), .Y(new_n24285_));
  OAI21X1  g21849(.A0(new_n24285_), .A1(new_n23312_), .B0(new_n24284_), .Y(new_n24286_));
  MX2X1    g21850(.A(new_n24286_), .B(new_n24283_), .S0(new_n11867_), .Y(new_n24287_));
  OAI21X1  g21851(.A0(new_n24287_), .A1(new_n5058_), .B0(pi0224), .Y(new_n24288_));
  OAI22X1  g21852(.A0(new_n24288_), .A1(new_n24282_), .B0(new_n24275_), .B1(new_n12389_), .Y(new_n24289_));
  AOI21X1  g21853(.A0(new_n24289_), .A1(pi0215), .B0(new_n2933_), .Y(new_n24290_));
  OAI21X1  g21854(.A0(new_n24274_), .A1(new_n24270_), .B0(new_n24290_), .Y(new_n24291_));
  OAI21X1  g21855(.A0(new_n24287_), .A1(new_n5041_), .B0(pi0224), .Y(new_n24292_));
  AOI21X1  g21856(.A0(new_n24281_), .A1(new_n5041_), .B0(new_n24292_), .Y(new_n24293_));
  OAI21X1  g21857(.A0(new_n24275_), .A1(new_n12380_), .B0(pi0223), .Y(new_n24294_));
  NAND2X1  g21858(.A(new_n24249_), .B(new_n5041_), .Y(new_n24295_));
  AOI21X1  g21859(.A0(new_n24260_), .A1(new_n5042_), .B0(new_n2942_), .Y(new_n24296_));
  AND2X1   g21860(.A(new_n24296_), .B(new_n24295_), .Y(new_n24297_));
  AND2X1   g21861(.A(new_n24265_), .B(new_n5042_), .Y(new_n24298_));
  AND2X1   g21862(.A(new_n2942_), .B(pi0222), .Y(new_n24299_));
  OAI21X1  g21863(.A0(new_n24266_), .A1(new_n5042_), .B0(new_n24299_), .Y(new_n24300_));
  AOI21X1  g21864(.A0(new_n12066_), .A1(pi0614), .B0(pi0223), .Y(new_n24301_));
  OAI21X1  g21865(.A0(new_n24300_), .A1(new_n24298_), .B0(new_n24301_), .Y(new_n24302_));
  OAI22X1  g21866(.A0(new_n24302_), .A1(new_n24297_), .B0(new_n24294_), .B1(new_n24293_), .Y(new_n24303_));
  AOI21X1  g21867(.A0(new_n24303_), .A1(new_n2933_), .B0(new_n2939_), .Y(new_n24304_));
  AOI21X1  g21868(.A0(new_n12041_), .A1(new_n11838_), .B0(new_n2942_), .Y(new_n24305_));
  NAND3X1  g21869(.A(new_n24305_), .B(new_n11973_), .C(new_n11968_), .Y(new_n24306_));
  NAND3X1  g21870(.A(new_n12041_), .B(pi0614), .C(new_n2942_), .Y(new_n24307_));
  AND3X1   g21871(.A(new_n24307_), .B(new_n24306_), .C(new_n2933_), .Y(new_n24308_));
  NOR4X1   g21872(.A(new_n12043_), .B(new_n12042_), .C(new_n11838_), .D(new_n11881_), .Y(new_n24309_));
  OAI21X1  g21873(.A0(new_n11965_), .A1(new_n2942_), .B0(new_n24309_), .Y(new_n24310_));
  OAI21X1  g21874(.A0(new_n11819_), .A1(new_n2942_), .B0(new_n24310_), .Y(new_n24311_));
  OAI21X1  g21875(.A0(new_n24311_), .A1(new_n2933_), .B0(new_n2939_), .Y(new_n24312_));
  OAI21X1  g21876(.A0(new_n24312_), .A1(new_n24308_), .B0(new_n2979_), .Y(new_n24313_));
  AOI21X1  g21877(.A0(new_n24304_), .A1(new_n24291_), .B0(new_n24313_), .Y(new_n24314_));
  AOI21X1  g21878(.A0(new_n12771_), .A1(pi0224), .B0(new_n2979_), .Y(new_n24315_));
  INVX1    g21879(.A(new_n24315_), .Y(new_n24316_));
  AOI21X1  g21880(.A0(new_n12079_), .A1(pi0614), .B0(new_n24316_), .Y(new_n24317_));
  OR2X1    g21881(.A(new_n24317_), .B(new_n11770_), .Y(new_n24318_));
  OAI22X1  g21882(.A0(new_n24318_), .A1(new_n24314_), .B0(new_n3103_), .B1(new_n2942_), .Y(new_n24319_));
  MX2X1    g21883(.A(new_n24319_), .B(new_n24241_), .S0(new_n12473_), .Y(new_n24320_));
  INVX1    g21884(.A(new_n24320_), .Y(new_n24321_));
  INVX1    g21885(.A(new_n24241_), .Y(new_n24322_));
  AOI21X1  g21886(.A0(new_n24322_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n24323_));
  OAI21X1  g21887(.A0(new_n24320_), .A1(new_n12462_), .B0(new_n24323_), .Y(new_n24324_));
  AOI21X1  g21888(.A0(new_n24322_), .A1(pi0609), .B0(pi1155), .Y(new_n24325_));
  OAI21X1  g21889(.A0(new_n24320_), .A1(pi0609), .B0(new_n24325_), .Y(new_n24326_));
  AND2X1   g21890(.A(new_n24326_), .B(new_n24324_), .Y(new_n24327_));
  MX2X1    g21891(.A(new_n24327_), .B(new_n24321_), .S0(new_n11768_), .Y(new_n24328_));
  NOR2X1   g21892(.A(new_n24328_), .B(pi0781), .Y(new_n24329_));
  INVX1    g21893(.A(new_n24328_), .Y(new_n24330_));
  AOI21X1  g21894(.A0(new_n24322_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n24331_));
  OAI21X1  g21895(.A0(new_n24330_), .A1(new_n12486_), .B0(new_n24331_), .Y(new_n24332_));
  AOI21X1  g21896(.A0(new_n24322_), .A1(pi0618), .B0(pi1154), .Y(new_n24333_));
  OAI21X1  g21897(.A0(new_n24330_), .A1(pi0618), .B0(new_n24333_), .Y(new_n24334_));
  AOI21X1  g21898(.A0(new_n24334_), .A1(new_n24332_), .B0(new_n11767_), .Y(new_n24335_));
  OAI21X1  g21899(.A0(new_n24335_), .A1(new_n24329_), .B0(new_n11766_), .Y(new_n24336_));
  NOR3X1   g21900(.A(new_n24335_), .B(new_n24329_), .C(new_n12509_), .Y(new_n24337_));
  OAI21X1  g21901(.A0(new_n24241_), .A1(pi0619), .B0(pi1159), .Y(new_n24338_));
  NOR2X1   g21902(.A(new_n24338_), .B(new_n24337_), .Y(new_n24339_));
  NOR3X1   g21903(.A(new_n24335_), .B(new_n24329_), .C(pi0619), .Y(new_n24340_));
  OAI21X1  g21904(.A0(new_n24241_), .A1(new_n12509_), .B0(new_n12510_), .Y(new_n24341_));
  NOR2X1   g21905(.A(new_n24341_), .B(new_n24340_), .Y(new_n24342_));
  OAI21X1  g21906(.A0(new_n24342_), .A1(new_n24339_), .B0(pi0789), .Y(new_n24343_));
  AND2X1   g21907(.A(new_n24343_), .B(new_n24336_), .Y(new_n24344_));
  INVX1    g21908(.A(new_n24344_), .Y(new_n24345_));
  MX2X1    g21909(.A(new_n24345_), .B(new_n24241_), .S0(new_n12708_), .Y(new_n24346_));
  NAND2X1  g21910(.A(new_n24346_), .B(new_n14249_), .Y(new_n24347_));
  AND2X1   g21911(.A(pi0680), .B(pi0662), .Y(new_n24348_));
  INVX1    g21912(.A(new_n24348_), .Y(new_n24349_));
  AND3X1   g21913(.A(new_n24349_), .B(new_n12322_), .C(new_n12318_), .Y(new_n24350_));
  AOI21X1  g21914(.A0(new_n12322_), .A1(new_n12318_), .B0(pi0224), .Y(new_n24351_));
  OAI21X1  g21915(.A0(new_n12310_), .A1(new_n2942_), .B0(new_n2933_), .Y(new_n24352_));
  NOR3X1   g21916(.A(new_n24352_), .B(new_n24351_), .C(new_n24350_), .Y(new_n24353_));
  AND3X1   g21917(.A(new_n24349_), .B(new_n12327_), .C(new_n12326_), .Y(new_n24354_));
  AOI21X1  g21918(.A0(new_n12327_), .A1(new_n12326_), .B0(pi0224), .Y(new_n24355_));
  NOR2X1   g21919(.A(new_n12312_), .B(new_n2942_), .Y(new_n24356_));
  NOR4X1   g21920(.A(new_n24356_), .B(new_n24355_), .C(new_n24354_), .D(new_n2933_), .Y(new_n24357_));
  OR3X1    g21921(.A(new_n24357_), .B(new_n24353_), .C(pi0039), .Y(new_n24358_));
  OAI21X1  g21922(.A0(new_n24349_), .A1(new_n12177_), .B0(new_n24271_), .Y(new_n24359_));
  MX2X1    g21923(.A(new_n12814_), .B(new_n11924_), .S0(new_n11849_), .Y(new_n24360_));
  OAI21X1  g21924(.A0(new_n23604_), .A1(new_n11850_), .B0(new_n11932_), .Y(new_n24361_));
  OAI21X1  g21925(.A0(new_n24361_), .A1(new_n5058_), .B0(pi0224), .Y(new_n24362_));
  AOI21X1  g21926(.A0(new_n24360_), .A1(new_n5058_), .B0(new_n24362_), .Y(new_n24363_));
  AND3X1   g21927(.A(new_n12205_), .B(new_n11926_), .C(pi0662), .Y(new_n24364_));
  NOR2X1   g21928(.A(new_n24364_), .B(new_n5058_), .Y(new_n24365_));
  NOR2X1   g21929(.A(new_n24349_), .B(new_n12370_), .Y(new_n24366_));
  OAI21X1  g21930(.A0(new_n24366_), .A1(new_n5059_), .B0(new_n2942_), .Y(new_n24367_));
  OAI21X1  g21931(.A0(new_n24367_), .A1(new_n24365_), .B0(new_n10045_), .Y(new_n24368_));
  OAI21X1  g21932(.A0(new_n24368_), .A1(new_n24363_), .B0(new_n24359_), .Y(new_n24369_));
  AND2X1   g21933(.A(new_n24369_), .B(new_n2934_), .Y(new_n24370_));
  MX2X1    g21934(.A(new_n23618_), .B(new_n11953_), .S0(new_n11849_), .Y(new_n24371_));
  MX2X1    g21935(.A(new_n23614_), .B(new_n11877_), .S0(new_n11849_), .Y(new_n24372_));
  AOI21X1  g21936(.A0(new_n24372_), .A1(new_n5058_), .B0(new_n2942_), .Y(new_n24373_));
  OAI21X1  g21937(.A0(new_n24371_), .A1(new_n5058_), .B0(new_n24373_), .Y(new_n24374_));
  AND2X1   g21938(.A(pi0662), .B(new_n2942_), .Y(new_n24375_));
  AOI21X1  g21939(.A0(new_n24375_), .A1(new_n12390_), .B0(new_n2934_), .Y(new_n24376_));
  AOI21X1  g21940(.A0(new_n24376_), .A1(new_n24374_), .B0(new_n2933_), .Y(new_n24377_));
  INVX1    g21941(.A(new_n24377_), .Y(new_n24378_));
  OAI21X1  g21942(.A0(new_n24361_), .A1(new_n5041_), .B0(pi0224), .Y(new_n24379_));
  AOI21X1  g21943(.A0(new_n24360_), .A1(new_n5041_), .B0(new_n24379_), .Y(new_n24380_));
  OR2X1    g21944(.A(new_n24364_), .B(new_n5041_), .Y(new_n24381_));
  OAI21X1  g21945(.A0(new_n24349_), .A1(new_n12370_), .B0(new_n5041_), .Y(new_n24382_));
  AND3X1   g21946(.A(new_n24382_), .B(new_n24381_), .C(new_n24299_), .Y(new_n24383_));
  AND2X1   g21947(.A(new_n12369_), .B(pi0662), .Y(new_n24384_));
  NOR4X1   g21948(.A(new_n24384_), .B(new_n24383_), .C(new_n24380_), .D(pi0223), .Y(new_n24385_));
  INVX1    g21949(.A(new_n24385_), .Y(new_n24386_));
  AOI21X1  g21950(.A0(new_n24372_), .A1(new_n5041_), .B0(new_n2942_), .Y(new_n24387_));
  OAI21X1  g21951(.A0(new_n24371_), .A1(new_n5041_), .B0(new_n24387_), .Y(new_n24388_));
  AOI21X1  g21952(.A0(new_n24375_), .A1(new_n12381_), .B0(new_n2940_), .Y(new_n24389_));
  AOI21X1  g21953(.A0(new_n24389_), .A1(new_n24388_), .B0(pi0299), .Y(new_n24390_));
  AOI21X1  g21954(.A0(new_n24390_), .A1(new_n24386_), .B0(new_n2939_), .Y(new_n24391_));
  OAI21X1  g21955(.A0(new_n24378_), .A1(new_n24370_), .B0(new_n24391_), .Y(new_n24392_));
  AOI21X1  g21956(.A0(new_n24392_), .A1(new_n24358_), .B0(pi0038), .Y(new_n24393_));
  AND3X1   g21957(.A(new_n12439_), .B(new_n5782_), .C(pi0662), .Y(new_n24394_));
  OAI21X1  g21958(.A0(new_n24394_), .A1(new_n24316_), .B0(new_n3103_), .Y(new_n24395_));
  OAI22X1  g21959(.A0(new_n24395_), .A1(new_n24393_), .B0(new_n3103_), .B1(new_n2942_), .Y(new_n24396_));
  INVX1    g21960(.A(new_n24396_), .Y(new_n24397_));
  OR2X1    g21961(.A(new_n24396_), .B(new_n12363_), .Y(new_n24398_));
  AOI21X1  g21962(.A0(new_n24322_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n24399_));
  OR2X1    g21963(.A(new_n24396_), .B(pi0625), .Y(new_n24400_));
  AOI21X1  g21964(.A0(new_n24322_), .A1(pi0625), .B0(pi1153), .Y(new_n24401_));
  AOI22X1  g21965(.A0(new_n24401_), .A1(new_n24400_), .B0(new_n24399_), .B1(new_n24398_), .Y(new_n24402_));
  MX2X1    g21966(.A(new_n24402_), .B(new_n24397_), .S0(new_n11769_), .Y(new_n24403_));
  MX2X1    g21967(.A(new_n24403_), .B(new_n24322_), .S0(new_n12490_), .Y(new_n24404_));
  MX2X1    g21968(.A(new_n24404_), .B(new_n24322_), .S0(new_n12513_), .Y(new_n24405_));
  AND3X1   g21969(.A(new_n24405_), .B(new_n13356_), .C(new_n14051_), .Y(new_n24406_));
  AOI21X1  g21970(.A0(new_n24322_), .A1(new_n21878_), .B0(new_n24406_), .Y(new_n24407_));
  AOI21X1  g21971(.A0(new_n24322_), .A1(pi0628), .B0(new_n23657_), .Y(new_n24408_));
  OAI21X1  g21972(.A0(new_n24407_), .A1(pi0628), .B0(new_n24408_), .Y(new_n24409_));
  AOI21X1  g21973(.A0(new_n24322_), .A1(new_n12554_), .B0(new_n21973_), .Y(new_n24410_));
  OAI21X1  g21974(.A0(new_n24407_), .A1(new_n12554_), .B0(new_n24410_), .Y(new_n24411_));
  NAND3X1  g21975(.A(new_n24411_), .B(new_n24409_), .C(new_n24347_), .Y(new_n24412_));
  MX2X1    g21976(.A(new_n23790_), .B(new_n16396_), .S0(new_n11838_), .Y(new_n24413_));
  AOI21X1  g21977(.A0(new_n24413_), .A1(new_n12274_), .B0(new_n11871_), .Y(new_n24414_));
  OR2X1    g21978(.A(new_n12268_), .B(new_n11838_), .Y(new_n24415_));
  AOI21X1  g21979(.A0(new_n24415_), .A1(new_n23687_), .B0(pi0616), .Y(new_n24416_));
  NOR2X1   g21980(.A(new_n24416_), .B(new_n24414_), .Y(new_n24417_));
  MX2X1    g21981(.A(new_n24417_), .B(new_n24245_), .S0(new_n5019_), .Y(new_n24418_));
  NOR2X1   g21982(.A(new_n23230_), .B(pi0662), .Y(new_n24419_));
  INVX1    g21983(.A(new_n24419_), .Y(new_n24420_));
  NOR2X1   g21984(.A(new_n24420_), .B(new_n24245_), .Y(new_n24421_));
  AOI21X1  g21985(.A0(new_n24248_), .A1(new_n11863_), .B0(new_n24421_), .Y(new_n24422_));
  OAI21X1  g21986(.A0(new_n24418_), .A1(new_n11849_), .B0(new_n24422_), .Y(new_n24423_));
  INVX1    g21987(.A(new_n24266_), .Y(new_n24424_));
  NOR2X1   g21988(.A(new_n12225_), .B(new_n11871_), .Y(new_n24425_));
  NOR3X1   g21989(.A(new_n12174_), .B(new_n11871_), .C(pi0614), .Y(new_n24426_));
  OAI21X1  g21990(.A0(new_n24426_), .A1(new_n24425_), .B0(pi0680), .Y(new_n24427_));
  OAI21X1  g21991(.A0(new_n24273_), .A1(new_n23707_), .B0(new_n24427_), .Y(new_n24428_));
  MX2X1    g21992(.A(new_n24428_), .B(new_n24424_), .S0(new_n11849_), .Y(new_n24429_));
  AOI21X1  g21993(.A0(new_n24429_), .A1(new_n2942_), .B0(new_n5059_), .Y(new_n24430_));
  OAI21X1  g21994(.A0(new_n24423_), .A1(new_n2942_), .B0(new_n24430_), .Y(new_n24431_));
  OAI21X1  g21995(.A0(new_n12219_), .A1(new_n11838_), .B0(pi0680), .Y(new_n24432_));
  AOI21X1  g21996(.A0(new_n13156_), .A1(new_n11838_), .B0(new_n24432_), .Y(new_n24433_));
  OR2X1    g21997(.A(new_n24433_), .B(new_n24263_), .Y(new_n24434_));
  OAI21X1  g21998(.A0(new_n24420_), .A1(new_n24262_), .B0(new_n24264_), .Y(new_n24435_));
  AOI21X1  g21999(.A0(new_n24434_), .A1(pi0662), .B0(new_n24435_), .Y(new_n24436_));
  AOI21X1  g22000(.A0(new_n24254_), .A1(new_n24252_), .B0(pi0680), .Y(new_n24437_));
  AOI22X1  g22001(.A0(new_n24253_), .A1(new_n23669_), .B0(new_n23676_), .B1(pi0614), .Y(new_n24438_));
  AOI21X1  g22002(.A0(new_n24438_), .A1(new_n23672_), .B0(new_n5019_), .Y(new_n24439_));
  OAI21X1  g22003(.A0(new_n24439_), .A1(new_n24437_), .B0(pi0662), .Y(new_n24440_));
  AOI21X1  g22004(.A0(new_n24254_), .A1(new_n24252_), .B0(new_n24420_), .Y(new_n24441_));
  AOI21X1  g22005(.A0(new_n24259_), .A1(new_n11863_), .B0(new_n24441_), .Y(new_n24442_));
  AND2X1   g22006(.A(new_n24442_), .B(new_n24440_), .Y(new_n24443_));
  AOI21X1  g22007(.A0(new_n24443_), .A1(pi0224), .B0(new_n5058_), .Y(new_n24444_));
  OAI21X1  g22008(.A0(new_n24436_), .A1(pi0224), .B0(new_n24444_), .Y(new_n24445_));
  NAND3X1  g22009(.A(new_n24445_), .B(new_n24431_), .C(new_n10045_), .Y(new_n24446_));
  AOI21X1  g22010(.A0(new_n24348_), .A1(new_n12174_), .B0(new_n24273_), .Y(new_n24447_));
  OR2X1    g22011(.A(new_n24447_), .B(pi0224), .Y(new_n24448_));
  OR2X1    g22012(.A(new_n24348_), .B(new_n24242_), .Y(new_n24449_));
  OAI21X1  g22013(.A0(new_n24449_), .A1(new_n13175_), .B0(pi0224), .Y(new_n24450_));
  AOI21X1  g22014(.A0(new_n24413_), .A1(new_n24348_), .B0(new_n24450_), .Y(new_n24451_));
  NOR2X1   g22015(.A(new_n24451_), .B(new_n24272_), .Y(new_n24452_));
  AOI21X1  g22016(.A0(new_n24452_), .A1(new_n24448_), .B0(pi0215), .Y(new_n24453_));
  AOI21X1  g22017(.A0(new_n24415_), .A1(new_n12101_), .B0(pi0616), .Y(new_n24454_));
  OAI21X1  g22018(.A0(new_n24454_), .A1(new_n24414_), .B0(pi0680), .Y(new_n24455_));
  AND2X1   g22019(.A(new_n24455_), .B(new_n24278_), .Y(new_n24456_));
  AOI21X1  g22020(.A0(new_n24419_), .A1(new_n24277_), .B0(new_n24280_), .Y(new_n24457_));
  OAI21X1  g22021(.A0(new_n24456_), .A1(new_n11849_), .B0(new_n24457_), .Y(new_n24458_));
  OAI21X1  g22022(.A0(new_n24137_), .A1(new_n11838_), .B0(new_n12112_), .Y(new_n24459_));
  MX2X1    g22023(.A(new_n24459_), .B(new_n24283_), .S0(new_n5019_), .Y(new_n24460_));
  NAND2X1  g22024(.A(new_n24460_), .B(pi0662), .Y(new_n24461_));
  AOI22X1  g22025(.A0(new_n24419_), .A1(new_n24283_), .B0(new_n24286_), .B1(new_n11863_), .Y(new_n24462_));
  AOI21X1  g22026(.A0(new_n24462_), .A1(new_n24461_), .B0(new_n5058_), .Y(new_n24463_));
  OR2X1    g22027(.A(new_n24463_), .B(new_n2942_), .Y(new_n24464_));
  AOI21X1  g22028(.A0(new_n24458_), .A1(new_n5058_), .B0(new_n24464_), .Y(new_n24465_));
  OR2X1    g22029(.A(new_n23513_), .B(new_n11838_), .Y(new_n24466_));
  AND2X1   g22030(.A(new_n12198_), .B(pi0680), .Y(new_n24467_));
  OAI21X1  g22031(.A0(new_n24467_), .A1(new_n24273_), .B0(new_n24427_), .Y(new_n24468_));
  MX2X1    g22032(.A(new_n24468_), .B(new_n24466_), .S0(new_n11849_), .Y(new_n24469_));
  NOR2X1   g22033(.A(new_n24469_), .B(new_n5059_), .Y(new_n24470_));
  OAI21X1  g22034(.A0(new_n24466_), .A1(new_n11836_), .B0(new_n11849_), .Y(new_n24471_));
  NOR3X1   g22035(.A(new_n12187_), .B(new_n11871_), .C(pi0614), .Y(new_n24472_));
  OAI21X1  g22036(.A0(new_n23736_), .A1(new_n11838_), .B0(pi0680), .Y(new_n24473_));
  NOR2X1   g22037(.A(new_n24473_), .B(new_n24472_), .Y(new_n24474_));
  AND2X1   g22038(.A(new_n24474_), .B(new_n12193_), .Y(new_n24475_));
  OR2X1    g22039(.A(pi0680), .B(new_n11838_), .Y(new_n24476_));
  OAI21X1  g22040(.A0(new_n24476_), .A1(new_n23924_), .B0(pi0662), .Y(new_n24477_));
  OAI21X1  g22041(.A0(new_n24477_), .A1(new_n24475_), .B0(new_n24471_), .Y(new_n24478_));
  OAI21X1  g22042(.A0(new_n24478_), .A1(new_n5058_), .B0(new_n2942_), .Y(new_n24479_));
  OAI21X1  g22043(.A0(new_n24479_), .A1(new_n24470_), .B0(pi0215), .Y(new_n24480_));
  OAI21X1  g22044(.A0(new_n24480_), .A1(new_n24465_), .B0(pi0299), .Y(new_n24481_));
  AOI21X1  g22045(.A0(new_n24453_), .A1(new_n24446_), .B0(new_n24481_), .Y(new_n24482_));
  AOI21X1  g22046(.A0(new_n24443_), .A1(new_n5042_), .B0(new_n2942_), .Y(new_n24483_));
  OAI21X1  g22047(.A0(new_n24423_), .A1(new_n5042_), .B0(new_n24483_), .Y(new_n24484_));
  OR2X1    g22048(.A(new_n24436_), .B(new_n5041_), .Y(new_n24485_));
  INVX1    g22049(.A(new_n24299_), .Y(new_n24486_));
  AOI21X1  g22050(.A0(new_n24429_), .A1(new_n5041_), .B0(new_n24486_), .Y(new_n24487_));
  OAI21X1  g22051(.A0(new_n24448_), .A1(pi0222), .B0(new_n2940_), .Y(new_n24488_));
  AOI21X1  g22052(.A0(new_n24487_), .A1(new_n24485_), .B0(new_n24488_), .Y(new_n24489_));
  AOI21X1  g22053(.A0(new_n24469_), .A1(new_n2942_), .B0(new_n5042_), .Y(new_n24490_));
  OAI21X1  g22054(.A0(new_n24458_), .A1(new_n2942_), .B0(new_n24490_), .Y(new_n24491_));
  NAND3X1  g22055(.A(new_n24462_), .B(new_n24461_), .C(pi0224), .Y(new_n24492_));
  AOI21X1  g22056(.A0(new_n24478_), .A1(new_n2942_), .B0(new_n5041_), .Y(new_n24493_));
  AOI21X1  g22057(.A0(new_n24493_), .A1(new_n24492_), .B0(new_n2940_), .Y(new_n24494_));
  AOI22X1  g22058(.A0(new_n24494_), .A1(new_n24491_), .B0(new_n24489_), .B1(new_n24484_), .Y(new_n24495_));
  OAI21X1  g22059(.A0(new_n24495_), .A1(pi0299), .B0(pi0039), .Y(new_n24496_));
  OAI22X1  g22060(.A0(new_n24349_), .A1(new_n23771_), .B0(new_n16612_), .B1(new_n11838_), .Y(new_n24497_));
  OR4X1    g22061(.A(new_n24348_), .B(new_n12324_), .C(new_n12323_), .D(new_n12316_), .Y(new_n24498_));
  AND3X1   g22062(.A(new_n24498_), .B(new_n24305_), .C(new_n24170_), .Y(new_n24499_));
  AOI21X1  g22063(.A0(new_n24497_), .A1(new_n2942_), .B0(new_n24499_), .Y(new_n24500_));
  NOR4X1   g22064(.A(new_n12043_), .B(new_n12042_), .C(pi0614), .D(new_n11881_), .Y(new_n24501_));
  OAI21X1  g22065(.A0(new_n24501_), .A1(new_n23780_), .B0(pi0224), .Y(new_n24502_));
  OAI21X1  g22066(.A0(new_n12330_), .A1(new_n12328_), .B0(new_n2942_), .Y(new_n24503_));
  OAI21X1  g22067(.A0(new_n24503_), .A1(new_n24309_), .B0(new_n24502_), .Y(new_n24504_));
  AND2X1   g22068(.A(new_n24504_), .B(new_n24348_), .Y(new_n24505_));
  OAI21X1  g22069(.A0(new_n24348_), .A1(new_n24311_), .B0(pi0299), .Y(new_n24506_));
  OAI22X1  g22070(.A0(new_n24506_), .A1(new_n24505_), .B0(new_n24500_), .B1(pi0299), .Y(new_n24507_));
  AOI21X1  g22071(.A0(new_n24507_), .A1(new_n2939_), .B0(pi0038), .Y(new_n24508_));
  OAI21X1  g22072(.A0(new_n24496_), .A1(new_n24482_), .B0(new_n24508_), .Y(new_n24509_));
  NAND3X1  g22073(.A(new_n12141_), .B(new_n12077_), .C(pi0662), .Y(new_n24510_));
  AOI21X1  g22074(.A0(new_n24510_), .A1(new_n24317_), .B0(new_n11770_), .Y(new_n24511_));
  AOI22X1  g22075(.A0(new_n24511_), .A1(new_n24509_), .B0(new_n11770_), .B1(pi0224), .Y(new_n24512_));
  AND2X1   g22076(.A(new_n24512_), .B(new_n12363_), .Y(new_n24513_));
  OAI21X1  g22077(.A0(new_n24319_), .A1(new_n12363_), .B0(new_n12364_), .Y(new_n24514_));
  AOI21X1  g22078(.A0(new_n24399_), .A1(new_n24398_), .B0(pi0608), .Y(new_n24515_));
  OAI21X1  g22079(.A0(new_n24514_), .A1(new_n24513_), .B0(new_n24515_), .Y(new_n24516_));
  AND2X1   g22080(.A(new_n24512_), .B(pi0625), .Y(new_n24517_));
  OAI21X1  g22081(.A0(new_n24319_), .A1(pi0625), .B0(pi1153), .Y(new_n24518_));
  AOI21X1  g22082(.A0(new_n24401_), .A1(new_n24400_), .B0(new_n12368_), .Y(new_n24519_));
  OAI21X1  g22083(.A0(new_n24518_), .A1(new_n24517_), .B0(new_n24519_), .Y(new_n24520_));
  AOI21X1  g22084(.A0(new_n24520_), .A1(new_n24516_), .B0(new_n11769_), .Y(new_n24521_));
  AOI21X1  g22085(.A0(new_n24512_), .A1(new_n11769_), .B0(new_n24521_), .Y(new_n24522_));
  AOI21X1  g22086(.A0(new_n24403_), .A1(pi0609), .B0(pi1155), .Y(new_n24523_));
  OAI21X1  g22087(.A0(new_n24522_), .A1(pi0609), .B0(new_n24523_), .Y(new_n24524_));
  AND3X1   g22088(.A(new_n24524_), .B(new_n24324_), .C(new_n12468_), .Y(new_n24525_));
  AOI21X1  g22089(.A0(new_n24403_), .A1(new_n12462_), .B0(new_n12463_), .Y(new_n24526_));
  OAI21X1  g22090(.A0(new_n24522_), .A1(new_n12462_), .B0(new_n24526_), .Y(new_n24527_));
  AND3X1   g22091(.A(new_n24527_), .B(new_n24326_), .C(pi0660), .Y(new_n24528_));
  OAI21X1  g22092(.A0(new_n24528_), .A1(new_n24525_), .B0(pi0785), .Y(new_n24529_));
  OAI21X1  g22093(.A0(new_n24522_), .A1(pi0785), .B0(new_n24529_), .Y(new_n24530_));
  INVX1    g22094(.A(new_n24404_), .Y(new_n24531_));
  OAI21X1  g22095(.A0(new_n24531_), .A1(new_n12486_), .B0(new_n12487_), .Y(new_n24532_));
  AOI21X1  g22096(.A0(new_n24530_), .A1(new_n12486_), .B0(new_n24532_), .Y(new_n24533_));
  NAND2X1  g22097(.A(new_n24332_), .B(new_n12494_), .Y(new_n24534_));
  OAI21X1  g22098(.A0(new_n24531_), .A1(pi0618), .B0(pi1154), .Y(new_n24535_));
  AOI21X1  g22099(.A0(new_n24530_), .A1(pi0618), .B0(new_n24535_), .Y(new_n24536_));
  NAND2X1  g22100(.A(new_n24334_), .B(pi0627), .Y(new_n24537_));
  OAI22X1  g22101(.A0(new_n24537_), .A1(new_n24536_), .B0(new_n24534_), .B1(new_n24533_), .Y(new_n24538_));
  MX2X1    g22102(.A(new_n24538_), .B(new_n24530_), .S0(new_n11767_), .Y(new_n24539_));
  NAND2X1  g22103(.A(new_n24539_), .B(new_n12509_), .Y(new_n24540_));
  AOI21X1  g22104(.A0(new_n24405_), .A1(pi0619), .B0(pi1159), .Y(new_n24541_));
  OAI21X1  g22105(.A0(new_n24338_), .A1(new_n24337_), .B0(new_n12517_), .Y(new_n24542_));
  AOI21X1  g22106(.A0(new_n24541_), .A1(new_n24540_), .B0(new_n24542_), .Y(new_n24543_));
  AND2X1   g22107(.A(new_n24405_), .B(new_n12509_), .Y(new_n24544_));
  OR2X1    g22108(.A(new_n24544_), .B(new_n12510_), .Y(new_n24545_));
  AOI21X1  g22109(.A0(new_n24539_), .A1(pi0619), .B0(new_n24545_), .Y(new_n24546_));
  OAI21X1  g22110(.A0(new_n24341_), .A1(new_n24340_), .B0(pi0648), .Y(new_n24547_));
  OAI21X1  g22111(.A0(new_n24547_), .A1(new_n24546_), .B0(pi0789), .Y(new_n24548_));
  OR2X1    g22112(.A(new_n24539_), .B(pi0789), .Y(new_n24549_));
  AND2X1   g22113(.A(new_n24549_), .B(new_n12709_), .Y(new_n24550_));
  OAI21X1  g22114(.A0(new_n24548_), .A1(new_n24543_), .B0(new_n24550_), .Y(new_n24551_));
  OAI21X1  g22115(.A0(new_n24322_), .A1(pi0626), .B0(new_n16221_), .Y(new_n24552_));
  AOI21X1  g22116(.A0(new_n24345_), .A1(pi0626), .B0(new_n24552_), .Y(new_n24553_));
  OAI21X1  g22117(.A0(new_n24322_), .A1(new_n12542_), .B0(new_n16217_), .Y(new_n24554_));
  AOI21X1  g22118(.A0(new_n24345_), .A1(new_n12542_), .B0(new_n24554_), .Y(new_n24555_));
  MX2X1    g22119(.A(new_n24405_), .B(new_n24322_), .S0(new_n12531_), .Y(new_n24556_));
  AND2X1   g22120(.A(new_n24556_), .B(new_n12637_), .Y(new_n24557_));
  OR3X1    g22121(.A(new_n24557_), .B(new_n24555_), .C(new_n24553_), .Y(new_n24558_));
  AOI21X1  g22122(.A0(new_n24558_), .A1(pi0788), .B0(new_n14125_), .Y(new_n24559_));
  AOI22X1  g22123(.A0(new_n24559_), .A1(new_n24551_), .B0(new_n24412_), .B1(pi0792), .Y(new_n24560_));
  MX2X1    g22124(.A(new_n24346_), .B(new_n24241_), .S0(new_n12580_), .Y(new_n24561_));
  OAI22X1  g22125(.A0(new_n24407_), .A1(new_n13508_), .B0(new_n24241_), .B1(new_n22699_), .Y(new_n24562_));
  OAI21X1  g22126(.A0(new_n24241_), .A1(pi0647), .B0(pi1157), .Y(new_n24563_));
  AOI21X1  g22127(.A0(new_n24562_), .A1(pi0647), .B0(new_n24563_), .Y(new_n24564_));
  OAI21X1  g22128(.A0(new_n24241_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n24565_));
  AOI21X1  g22129(.A0(new_n24562_), .A1(new_n12577_), .B0(new_n24565_), .Y(new_n24566_));
  MX2X1    g22130(.A(new_n24566_), .B(new_n24564_), .S0(new_n12592_), .Y(new_n24567_));
  AOI21X1  g22131(.A0(new_n24561_), .A1(new_n14326_), .B0(new_n24567_), .Y(new_n24568_));
  OAI22X1  g22132(.A0(new_n24568_), .A1(new_n11763_), .B0(new_n24560_), .B1(new_n14121_), .Y(new_n24569_));
  NOR2X1   g22133(.A(new_n24566_), .B(new_n24564_), .Y(new_n24570_));
  MX2X1    g22134(.A(new_n24570_), .B(new_n24562_), .S0(new_n11763_), .Y(new_n24571_));
  AOI21X1  g22135(.A0(new_n24571_), .A1(new_n12612_), .B0(new_n12608_), .Y(new_n24572_));
  OAI21X1  g22136(.A0(new_n24569_), .A1(new_n12612_), .B0(new_n24572_), .Y(new_n24573_));
  MX2X1    g22137(.A(new_n24561_), .B(new_n24241_), .S0(new_n12604_), .Y(new_n24574_));
  AOI21X1  g22138(.A0(new_n24322_), .A1(new_n12612_), .B0(pi0715), .Y(new_n24575_));
  OAI21X1  g22139(.A0(new_n24574_), .A1(new_n12612_), .B0(new_n24575_), .Y(new_n24576_));
  AND2X1   g22140(.A(new_n24576_), .B(pi1160), .Y(new_n24577_));
  AOI21X1  g22141(.A0(new_n24571_), .A1(pi0644), .B0(pi0715), .Y(new_n24578_));
  OAI21X1  g22142(.A0(new_n24569_), .A1(pi0644), .B0(new_n24578_), .Y(new_n24579_));
  AOI21X1  g22143(.A0(new_n24322_), .A1(pi0644), .B0(new_n12608_), .Y(new_n24580_));
  OAI21X1  g22144(.A0(new_n24574_), .A1(pi0644), .B0(new_n24580_), .Y(new_n24581_));
  AND2X1   g22145(.A(new_n24581_), .B(new_n11762_), .Y(new_n24582_));
  AOI22X1  g22146(.A0(new_n24582_), .A1(new_n24579_), .B0(new_n24577_), .B1(new_n24573_), .Y(new_n24583_));
  MX2X1    g22147(.A(new_n24583_), .B(new_n24569_), .S0(new_n12766_), .Y(new_n24584_));
  MX2X1    g22148(.A(new_n24584_), .B(pi0224), .S0(po1038), .Y(po0381));
  OR2X1    g22149(.A(new_n5814_), .B(pi0056), .Y(new_n24586_));
  AOI21X1  g22150(.A0(new_n5071_), .A1(new_n7564_), .B0(pi0137), .Y(new_n24587_));
  NOR4X1   g22151(.A(new_n24587_), .B(new_n5075_), .C(new_n2986_), .D(pi0039), .Y(new_n24588_));
  NAND2X1  g22152(.A(new_n8450_), .B(new_n2852_), .Y(new_n24589_));
  OAI21X1  g22153(.A0(new_n24589_), .A1(new_n2687_), .B0(new_n2533_), .Y(new_n24590_));
  AOI21X1  g22154(.A0(new_n24590_), .A1(new_n2528_), .B0(new_n2710_), .Y(new_n24591_));
  OAI21X1  g22155(.A0(new_n24591_), .A1(pi0095), .B0(new_n2794_), .Y(new_n24592_));
  INVX1    g22156(.A(new_n8538_), .Y(new_n24593_));
  OAI21X1  g22157(.A0(new_n8450_), .A1(new_n22518_), .B0(new_n2782_), .Y(new_n24594_));
  AND3X1   g22158(.A(new_n24594_), .B(new_n2714_), .C(new_n2523_), .Y(new_n24595_));
  NOR3X1   g22159(.A(new_n2762_), .B(new_n2710_), .C(pi0095), .Y(new_n24596_));
  OR2X1    g22160(.A(new_n5905_), .B(new_n22518_), .Y(new_n24597_));
  NOR4X1   g22161(.A(new_n24597_), .B(new_n2689_), .C(new_n2535_), .D(pi0051), .Y(new_n24598_));
  AOI22X1  g22162(.A0(new_n24598_), .A1(new_n24596_), .B0(new_n24595_), .B1(new_n2762_), .Y(new_n24599_));
  INVX1    g22163(.A(new_n24599_), .Y(new_n24600_));
  INVX1    g22164(.A(new_n24595_), .Y(new_n24601_));
  OAI21X1  g22165(.A0(new_n24597_), .A1(new_n2512_), .B0(new_n2455_), .Y(new_n24602_));
  AOI21X1  g22166(.A0(new_n24602_), .A1(new_n24596_), .B0(pi1093), .Y(new_n24603_));
  AOI22X1  g22167(.A0(new_n24599_), .A1(new_n24603_), .B0(new_n24601_), .B1(pi1093), .Y(new_n24604_));
  OR3X1    g22168(.A(new_n2761_), .B(new_n2756_), .C(new_n2782_), .Y(new_n24605_));
  AND2X1   g22169(.A(new_n24605_), .B(new_n24603_), .Y(new_n24606_));
  OAI21X1  g22170(.A0(new_n24597_), .A1(new_n2736_), .B0(new_n2455_), .Y(new_n24607_));
  NAND2X1  g22171(.A(new_n24605_), .B(pi1093), .Y(new_n24608_));
  AOI21X1  g22172(.A0(new_n24607_), .A1(new_n24596_), .B0(new_n24608_), .Y(new_n24609_));
  OAI21X1  g22173(.A0(new_n24609_), .A1(new_n24606_), .B0(new_n8515_), .Y(new_n24610_));
  OAI22X1  g22174(.A0(new_n24610_), .A1(new_n24600_), .B0(new_n24604_), .B1(new_n24593_), .Y(new_n24611_));
  AOI21X1  g22175(.A0(new_n24592_), .A1(pi0137), .B0(new_n24611_), .Y(new_n24612_));
  AOI21X1  g22176(.A0(new_n2711_), .A1(new_n2794_), .B0(new_n2452_), .Y(new_n24613_));
  NOR2X1   g22177(.A(new_n2783_), .B(new_n5032_), .Y(new_n24614_));
  OAI21X1  g22178(.A0(new_n24614_), .A1(new_n24606_), .B0(new_n8538_), .Y(new_n24615_));
  NAND2X1  g22179(.A(new_n24615_), .B(new_n24610_), .Y(new_n24616_));
  NOR2X1   g22180(.A(new_n24616_), .B(new_n24613_), .Y(new_n24617_));
  MX2X1    g22181(.A(new_n24617_), .B(new_n24612_), .S0(pi0332), .Y(new_n24618_));
  NAND2X1  g22182(.A(new_n24618_), .B(new_n3038_), .Y(new_n24619_));
  MX2X1    g22183(.A(new_n24601_), .B(new_n24592_), .S0(pi0137), .Y(new_n24620_));
  NAND2X1  g22184(.A(new_n24620_), .B(pi0332), .Y(new_n24621_));
  OAI21X1  g22185(.A0(new_n24613_), .A1(new_n2784_), .B0(new_n2444_), .Y(new_n24622_));
  NAND3X1  g22186(.A(new_n24622_), .B(new_n24621_), .C(new_n2815_), .Y(new_n24623_));
  AND2X1   g22187(.A(new_n24623_), .B(new_n2777_), .Y(new_n24624_));
  AOI21X1  g22188(.A0(new_n2794_), .A1(new_n2694_), .B0(new_n2452_), .Y(new_n24625_));
  OR2X1    g22189(.A(new_n24625_), .B(new_n2750_), .Y(new_n24626_));
  AOI21X1  g22190(.A0(new_n24590_), .A1(new_n2528_), .B0(new_n2481_), .Y(new_n24627_));
  OAI21X1  g22191(.A0(new_n24627_), .A1(pi0095), .B0(new_n2825_), .Y(new_n24628_));
  NOR3X1   g22192(.A(new_n2481_), .B(pi0137), .C(pi0095), .Y(new_n24629_));
  AOI21X1  g22193(.A0(new_n24629_), .A1(new_n24594_), .B0(new_n2444_), .Y(new_n24630_));
  AOI22X1  g22194(.A0(new_n24630_), .A1(new_n24628_), .B0(new_n24626_), .B1(new_n2444_), .Y(new_n24631_));
  OAI21X1  g22195(.A0(new_n24631_), .A1(new_n2777_), .B0(pi0299), .Y(new_n24632_));
  AOI21X1  g22196(.A0(new_n24624_), .A1(new_n24619_), .B0(new_n24632_), .Y(new_n24633_));
  NAND3X1  g22197(.A(new_n24622_), .B(new_n24621_), .C(new_n5069_), .Y(new_n24634_));
  AOI21X1  g22198(.A0(new_n24618_), .A1(new_n5070_), .B0(pi0198), .Y(new_n24635_));
  OAI21X1  g22199(.A0(new_n24631_), .A1(new_n2954_), .B0(new_n2933_), .Y(new_n24636_));
  AOI21X1  g22200(.A0(new_n24635_), .A1(new_n24634_), .B0(new_n24636_), .Y(new_n24637_));
  OAI21X1  g22201(.A0(new_n24637_), .A1(new_n24633_), .B0(new_n2939_), .Y(new_n24638_));
  AOI21X1  g22202(.A0(new_n2998_), .A1(pi0039), .B0(pi0038), .Y(new_n24639_));
  OAI21X1  g22203(.A0(pi0137), .A1(new_n2979_), .B0(new_n4988_), .Y(new_n24640_));
  AOI21X1  g22204(.A0(new_n24639_), .A1(new_n24638_), .B0(new_n24640_), .Y(new_n24641_));
  OAI21X1  g22205(.A0(new_n24641_), .A1(new_n24588_), .B0(new_n3131_), .Y(new_n24642_));
  NOR4X1   g22206(.A(new_n3132_), .B(new_n2985_), .C(new_n2536_), .D(new_n2452_), .Y(new_n24643_));
  AOI21X1  g22207(.A0(new_n24643_), .A1(pi0087), .B0(pi0075), .Y(new_n24644_));
  NOR4X1   g22208(.A(new_n24587_), .B(new_n5778_), .C(new_n2986_), .D(pi0039), .Y(new_n24645_));
  OAI21X1  g22209(.A0(new_n24645_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n24646_));
  AOI21X1  g22210(.A0(new_n24644_), .A1(new_n24642_), .B0(new_n24646_), .Y(new_n24647_));
  AND3X1   g22211(.A(new_n24643_), .B(new_n3077_), .C(pi0092), .Y(new_n24648_));
  OR2X1    g22212(.A(new_n24648_), .B(pi0054), .Y(new_n24649_));
  NAND3X1  g22213(.A(new_n24643_), .B(new_n3077_), .C(new_n3079_), .Y(new_n24650_));
  AOI21X1  g22214(.A0(new_n24650_), .A1(pi0054), .B0(pi0074), .Y(new_n24651_));
  OAI21X1  g22215(.A0(new_n24649_), .A1(new_n24647_), .B0(new_n24651_), .Y(new_n24652_));
  AND2X1   g22216(.A(new_n4983_), .B(pi0074), .Y(new_n24653_));
  AOI21X1  g22217(.A0(new_n24653_), .A1(new_n24643_), .B0(pi0055), .Y(new_n24654_));
  AOI21X1  g22218(.A0(new_n24654_), .A1(new_n24652_), .B0(new_n24586_), .Y(new_n24655_));
  AND3X1   g22219(.A(new_n24643_), .B(new_n3113_), .C(pi0056), .Y(new_n24656_));
  OAI21X1  g22220(.A0(new_n24656_), .A1(new_n24655_), .B0(new_n3222_), .Y(new_n24657_));
  NAND3X1  g22221(.A(new_n24643_), .B(new_n5096_), .C(pi0062), .Y(new_n24658_));
  AND2X1   g22222(.A(new_n24658_), .B(new_n3223_), .Y(new_n24659_));
  AND3X1   g22223(.A(new_n24643_), .B(new_n5096_), .C(new_n3222_), .Y(new_n24660_));
  OAI21X1  g22224(.A0(new_n24660_), .A1(new_n3223_), .B0(new_n4974_), .Y(new_n24661_));
  AOI21X1  g22225(.A0(new_n24659_), .A1(new_n24657_), .B0(new_n24661_), .Y(po0382));
  AND2X1   g22226(.A(pi0231), .B(pi0228), .Y(new_n24663_));
  INVX1    g22227(.A(pi0231), .Y(new_n24664_));
  AOI21X1  g22228(.A0(new_n2846_), .A1(new_n2509_), .B0(pi0070), .Y(new_n24665_));
  OAI21X1  g22229(.A0(new_n24665_), .A1(pi0051), .B0(new_n2537_), .Y(new_n24666_));
  AOI21X1  g22230(.A0(new_n24666_), .A1(new_n2852_), .B0(new_n4990_), .Y(new_n24667_));
  OAI21X1  g22231(.A0(new_n24667_), .A1(new_n2795_), .B0(new_n5013_), .Y(new_n24668_));
  AOI21X1  g22232(.A0(new_n24668_), .A1(new_n2523_), .B0(new_n3237_), .Y(new_n24669_));
  AOI21X1  g22233(.A0(new_n2986_), .A1(pi0039), .B0(pi0038), .Y(new_n24670_));
  OAI21X1  g22234(.A0(new_n24669_), .A1(pi0039), .B0(new_n24670_), .Y(new_n24671_));
  MX2X1    g22235(.A(new_n24671_), .B(new_n24664_), .S0(pi0228), .Y(new_n24672_));
  INVX1    g22236(.A(new_n24663_), .Y(new_n24673_));
  OAI21X1  g22237(.A0(new_n3604_), .A1(new_n3060_), .B0(new_n24673_), .Y(new_n24674_));
  AOI21X1  g22238(.A0(new_n24674_), .A1(pi0100), .B0(pi0087), .Y(new_n24675_));
  OAI21X1  g22239(.A0(new_n24672_), .A1(pi0100), .B0(new_n24675_), .Y(new_n24676_));
  OR3X1    g22240(.A(new_n24663_), .B(new_n5819_), .C(new_n3131_), .Y(new_n24677_));
  AND3X1   g22241(.A(new_n24677_), .B(new_n24676_), .C(new_n3073_), .Y(new_n24678_));
  AOI21X1  g22242(.A0(new_n6777_), .A1(new_n5827_), .B0(new_n24663_), .Y(new_n24679_));
  OAI21X1  g22243(.A0(new_n24679_), .A1(new_n3073_), .B0(new_n3079_), .Y(new_n24680_));
  OR2X1    g22244(.A(new_n24663_), .B(new_n3079_), .Y(new_n24681_));
  OAI22X1  g22245(.A0(new_n24681_), .A1(new_n5834_), .B0(new_n24680_), .B1(new_n24678_), .Y(new_n24682_));
  OAI21X1  g22246(.A0(new_n24663_), .A1(new_n3091_), .B0(new_n4982_), .Y(new_n24683_));
  AOI21X1  g22247(.A0(new_n24682_), .A1(new_n3091_), .B0(new_n24683_), .Y(new_n24684_));
  OAI21X1  g22248(.A0(new_n24663_), .A1(new_n5841_), .B0(pi0074), .Y(new_n24685_));
  NAND2X1  g22249(.A(new_n24685_), .B(new_n3107_), .Y(new_n24686_));
  AOI21X1  g22250(.A0(new_n24673_), .A1(pi0055), .B0(pi0056), .Y(new_n24687_));
  OAI21X1  g22251(.A0(new_n24686_), .A1(new_n24684_), .B0(new_n24687_), .Y(new_n24688_));
  OAI21X1  g22252(.A0(new_n24663_), .A1(new_n5845_), .B0(pi0056), .Y(new_n24689_));
  AND2X1   g22253(.A(new_n24689_), .B(new_n3222_), .Y(new_n24690_));
  NOR3X1   g22254(.A(new_n24663_), .B(new_n5820_), .C(new_n3222_), .Y(new_n24691_));
  AOI21X1  g22255(.A0(new_n24690_), .A1(new_n24688_), .B0(new_n24691_), .Y(new_n24692_));
  MX2X1    g22256(.A(new_n24692_), .B(new_n24663_), .S0(new_n3374_), .Y(po0383));
  AND2X1   g22257(.A(new_n5150_), .B(new_n2479_), .Y(new_n24694_));
  OR4X1    g22258(.A(new_n8190_), .B(new_n8183_), .C(new_n5225_), .D(new_n2514_), .Y(new_n24695_));
  NOR2X1   g22259(.A(new_n11891_), .B(new_n2514_), .Y(new_n24696_));
  OAI21X1  g22260(.A0(new_n7671_), .A1(new_n2503_), .B0(new_n2515_), .Y(new_n24697_));
  AOI21X1  g22261(.A0(new_n24696_), .A1(new_n8198_), .B0(new_n24697_), .Y(new_n24698_));
  NAND2X1  g22262(.A(new_n24698_), .B(new_n24695_), .Y(new_n24699_));
  AOI21X1  g22263(.A0(new_n24699_), .A1(new_n24694_), .B0(pi0072), .Y(new_n24700_));
  OR2X1    g22264(.A(new_n24700_), .B(new_n5170_), .Y(new_n24701_));
  AOI21X1  g22265(.A0(new_n2704_), .A1(pi1093), .B0(new_n5237_), .Y(new_n24702_));
  INVX1    g22266(.A(new_n5239_), .Y(new_n24703_));
  NAND4X1  g22267(.A(new_n9485_), .B(new_n5927_), .C(new_n5169_), .D(new_n2479_), .Y(new_n24704_));
  AOI21X1  g22268(.A0(new_n24704_), .A1(new_n24703_), .B0(new_n5032_), .Y(new_n24705_));
  AOI21X1  g22269(.A0(new_n24697_), .A1(new_n24694_), .B0(pi0072), .Y(new_n24706_));
  NOR3X1   g22270(.A(new_n8190_), .B(new_n8183_), .C(new_n2514_), .Y(new_n24707_));
  AND3X1   g22271(.A(new_n24707_), .B(new_n5150_), .C(new_n2479_), .Y(new_n24708_));
  AOI22X1  g22272(.A0(new_n24708_), .A1(new_n5928_), .B0(new_n5032_), .B1(pi0829), .Y(new_n24709_));
  AOI21X1  g22273(.A0(new_n24709_), .A1(new_n24706_), .B0(new_n5170_), .Y(new_n24710_));
  INVX1    g22274(.A(new_n24708_), .Y(new_n24711_));
  AOI21X1  g22275(.A0(new_n24711_), .A1(new_n24706_), .B0(new_n5170_), .Y(new_n24712_));
  OAI22X1  g22276(.A0(new_n24712_), .A1(new_n9462_), .B0(new_n24710_), .B1(new_n24705_), .Y(new_n24713_));
  AOI21X1  g22277(.A0(new_n24702_), .A1(new_n24701_), .B0(new_n24713_), .Y(new_n24714_));
  OAI21X1  g22278(.A0(new_n24714_), .A1(pi0039), .B0(new_n8487_), .Y(po0384));
  OR2X1    g22279(.A(new_n8456_), .B(new_n8453_), .Y(new_n24716_));
  AND2X1   g22280(.A(new_n24716_), .B(pi0039), .Y(new_n24717_));
  NOR2X1   g22281(.A(new_n6740_), .B(new_n2759_), .Y(new_n24718_));
  OR3X1    g22282(.A(pi0095), .B(pi0039), .C(pi0032), .Y(new_n24719_));
  NOR4X1   g22283(.A(new_n24719_), .B(new_n24718_), .C(new_n8500_), .D(new_n2520_), .Y(new_n24720_));
  AOI21X1  g22284(.A0(new_n24717_), .A1(new_n5235_), .B0(new_n24720_), .Y(new_n24721_));
  OAI22X1  g22285(.A0(new_n24721_), .A1(new_n7629_), .B0(new_n2793_), .B1(pi0039), .Y(po0385));
  OAI21X1  g22286(.A0(new_n4986_), .A1(new_n2979_), .B0(new_n7625_), .Y(new_n24723_));
  INVX1    g22287(.A(new_n11824_), .Y(new_n24724_));
  NOR3X1   g22288(.A(new_n5031_), .B(new_n5922_), .C(new_n5032_), .Y(new_n24725_));
  AND2X1   g22289(.A(new_n24725_), .B(new_n11884_), .Y(new_n24726_));
  OAI21X1  g22290(.A0(new_n24725_), .A1(new_n11823_), .B0(pi1091), .Y(new_n24727_));
  OR2X1    g22291(.A(new_n24727_), .B(new_n24726_), .Y(new_n24728_));
  AOI21X1  g22292(.A0(new_n11826_), .A1(new_n5231_), .B0(pi1091), .Y(new_n24729_));
  OAI21X1  g22293(.A0(new_n11892_), .A1(new_n5231_), .B0(new_n24729_), .Y(new_n24730_));
  AND2X1   g22294(.A(new_n24730_), .B(new_n24728_), .Y(new_n24731_));
  MX2X1    g22295(.A(new_n24731_), .B(new_n2987_), .S0(pi0120), .Y(new_n24732_));
  MX2X1    g22296(.A(new_n24732_), .B(new_n24724_), .S0(new_n5043_), .Y(new_n24733_));
  NOR2X1   g22297(.A(new_n11824_), .B(new_n6255_), .Y(new_n24734_));
  AOI21X1  g22298(.A0(new_n24732_), .A1(new_n6255_), .B0(new_n24734_), .Y(new_n24735_));
  AOI21X1  g22299(.A0(new_n24735_), .A1(new_n5041_), .B0(new_n2951_), .Y(new_n24736_));
  OAI21X1  g22300(.A0(new_n24733_), .A1(new_n5041_), .B0(new_n24736_), .Y(new_n24737_));
  AOI21X1  g22301(.A0(new_n24724_), .A1(new_n2951_), .B0(pi0223), .Y(new_n24738_));
  NOR2X1   g22302(.A(new_n11824_), .B(new_n5044_), .Y(new_n24739_));
  INVX1    g22303(.A(new_n24739_), .Y(new_n24740_));
  AND2X1   g22304(.A(new_n5035_), .B(pi0120), .Y(new_n24741_));
  NOR2X1   g22305(.A(new_n24741_), .B(new_n11824_), .Y(new_n24742_));
  INVX1    g22306(.A(new_n24742_), .Y(new_n24743_));
  AOI21X1  g22307(.A0(new_n24743_), .A1(new_n24740_), .B0(new_n5041_), .Y(new_n24744_));
  NOR2X1   g22308(.A(new_n24742_), .B(new_n24734_), .Y(new_n24745_));
  OAI21X1  g22309(.A0(new_n24745_), .A1(new_n5042_), .B0(pi0223), .Y(new_n24746_));
  OAI21X1  g22310(.A0(new_n24746_), .A1(new_n24744_), .B0(new_n2933_), .Y(new_n24747_));
  AOI21X1  g22311(.A0(new_n24738_), .A1(new_n24737_), .B0(new_n24747_), .Y(new_n24748_));
  AOI21X1  g22312(.A0(new_n24735_), .A1(new_n5058_), .B0(new_n10044_), .Y(new_n24749_));
  OAI21X1  g22313(.A0(new_n24733_), .A1(new_n5058_), .B0(new_n24749_), .Y(new_n24750_));
  NOR2X1   g22314(.A(new_n12425_), .B(pi0215), .Y(new_n24751_));
  AOI21X1  g22315(.A0(new_n24743_), .A1(new_n24740_), .B0(new_n5058_), .Y(new_n24752_));
  OAI21X1  g22316(.A0(new_n24745_), .A1(new_n5059_), .B0(pi0215), .Y(new_n24753_));
  OAI21X1  g22317(.A0(new_n24753_), .A1(new_n24752_), .B0(pi0299), .Y(new_n24754_));
  AOI21X1  g22318(.A0(new_n24751_), .A1(new_n24750_), .B0(new_n24754_), .Y(new_n24755_));
  OAI21X1  g22319(.A0(new_n24755_), .A1(new_n24748_), .B0(pi0039), .Y(new_n24756_));
  AND2X1   g22320(.A(pi1091), .B(pi0829), .Y(new_n24757_));
  AOI21X1  g22321(.A0(new_n24757_), .A1(new_n11814_), .B0(pi0824), .Y(new_n24758_));
  INVX1    g22322(.A(new_n24758_), .Y(new_n24759_));
  OR2X1    g22323(.A(new_n11811_), .B(new_n11809_), .Y(new_n24760_));
  AOI21X1  g22324(.A0(new_n24760_), .A1(pi0824), .B0(new_n5232_), .Y(new_n24761_));
  AOI21X1  g22325(.A0(new_n24761_), .A1(new_n24759_), .B0(new_n11803_), .Y(new_n24762_));
  AOI22X1  g22326(.A0(new_n24758_), .A1(new_n24757_), .B0(new_n24760_), .B1(pi0824), .Y(new_n24763_));
  OR2X1    g22327(.A(new_n5232_), .B(new_n5230_), .Y(new_n24764_));
  OAI22X1  g22328(.A0(new_n24764_), .A1(new_n24763_), .B0(new_n5232_), .B1(new_n5009_), .Y(new_n24765_));
  NOR2X1   g22329(.A(new_n5232_), .B(new_n5009_), .Y(new_n24766_));
  NOR3X1   g22330(.A(new_n11788_), .B(new_n5927_), .C(new_n7250_), .Y(new_n24767_));
  OAI21X1  g22331(.A0(new_n24767_), .A1(new_n11801_), .B0(new_n24766_), .Y(new_n24768_));
  AND2X1   g22332(.A(new_n24768_), .B(pi1093), .Y(new_n24769_));
  OAI21X1  g22333(.A0(new_n24765_), .A1(new_n24762_), .B0(new_n24769_), .Y(new_n24770_));
  OR3X1    g22334(.A(new_n11788_), .B(new_n5882_), .C(new_n7250_), .Y(new_n24771_));
  NOR4X1   g22335(.A(new_n6954_), .B(new_n2553_), .C(new_n2728_), .D(pi0091), .Y(new_n24772_));
  AOI21X1  g22336(.A0(new_n24772_), .A1(new_n11782_), .B0(pi0040), .Y(new_n24773_));
  OAI21X1  g22337(.A0(new_n24773_), .A1(new_n7683_), .B0(pi0252), .Y(new_n24774_));
  AND2X1   g22338(.A(new_n11778_), .B(new_n5882_), .Y(new_n24775_));
  AOI21X1  g22339(.A0(new_n24775_), .A1(new_n24774_), .B0(pi1093), .Y(new_n24776_));
  AOI21X1  g22340(.A0(new_n24776_), .A1(new_n24771_), .B0(pi0039), .Y(new_n24777_));
  AOI21X1  g22341(.A0(new_n24777_), .A1(new_n24770_), .B0(pi0038), .Y(new_n24778_));
  AOI21X1  g22342(.A0(new_n24778_), .A1(new_n24756_), .B0(new_n24723_), .Y(po0387));
  INVX1    g22343(.A(new_n5785_), .Y(new_n24780_));
  OAI21X1  g22344(.A0(new_n2660_), .A1(pi0081), .B0(new_n5140_), .Y(new_n24781_));
  AOI21X1  g22345(.A0(new_n24781_), .A1(new_n5139_), .B0(new_n2666_), .Y(new_n24782_));
  OAI21X1  g22346(.A0(new_n24782_), .A1(new_n5154_), .B0(new_n2670_), .Y(new_n24783_));
  AOI21X1  g22347(.A0(new_n24783_), .A1(new_n2488_), .B0(new_n2575_), .Y(new_n24784_));
  OAI21X1  g22348(.A0(new_n24784_), .A1(pi0086), .B0(new_n2574_), .Y(new_n24785_));
  AOI21X1  g22349(.A0(new_n24785_), .A1(new_n2571_), .B0(new_n2565_), .Y(new_n24786_));
  OAI21X1  g22350(.A0(new_n24786_), .A1(pi0108), .B0(new_n2563_), .Y(new_n24787_));
  AOI21X1  g22351(.A0(new_n24787_), .A1(new_n2678_), .B0(new_n2557_), .Y(new_n24788_));
  OAI21X1  g22352(.A0(new_n24788_), .A1(new_n2556_), .B0(new_n2554_), .Y(new_n24789_));
  AOI21X1  g22353(.A0(new_n24789_), .A1(new_n2545_), .B0(new_n2836_), .Y(new_n24790_));
  OAI21X1  g22354(.A0(new_n24790_), .A1(new_n2525_), .B0(new_n11110_), .Y(new_n24791_));
  AOI21X1  g22355(.A0(new_n24791_), .A1(new_n2535_), .B0(new_n2848_), .Y(new_n24792_));
  OAI21X1  g22356(.A0(new_n24792_), .A1(pi0051), .B0(new_n2537_), .Y(new_n24793_));
  AOI21X1  g22357(.A0(new_n24793_), .A1(new_n2852_), .B0(new_n4990_), .Y(new_n24794_));
  OAI21X1  g22358(.A0(new_n7584_), .A1(pi1082), .B0(new_n2455_), .Y(new_n24795_));
  OAI21X1  g22359(.A0(new_n24795_), .A1(new_n24794_), .B0(new_n3176_), .Y(new_n24796_));
  AOI21X1  g22360(.A0(new_n24796_), .A1(new_n2523_), .B0(new_n2696_), .Y(new_n24797_));
  MX2X1    g22361(.A(new_n5062_), .B(new_n5049_), .S0(new_n2933_), .Y(new_n24798_));
  OR3X1    g22362(.A(new_n5034_), .B(new_n5031_), .C(new_n5230_), .Y(po0950));
  NOR3X1   g22363(.A(po0950), .B(new_n24798_), .C(new_n5223_), .Y(new_n24800_));
  NOR4X1   g22364(.A(new_n24800_), .B(new_n8420_), .C(new_n7634_), .D(pi0287), .Y(new_n24801_));
  AOI21X1  g22365(.A0(new_n2986_), .A1(pi0039), .B0(new_n24801_), .Y(new_n24802_));
  OAI21X1  g22366(.A0(new_n24797_), .A1(pi0039), .B0(new_n24802_), .Y(new_n24803_));
  AOI21X1  g22367(.A0(new_n24803_), .A1(new_n2979_), .B0(new_n4989_), .Y(new_n24804_));
  NOR2X1   g22368(.A(new_n5076_), .B(pi0087), .Y(new_n24805_));
  INVX1    g22369(.A(new_n24805_), .Y(new_n24806_));
  OAI21X1  g22370(.A0(new_n24806_), .A1(new_n24804_), .B0(new_n5090_), .Y(new_n24807_));
  AOI21X1  g22371(.A0(new_n24807_), .A1(new_n3084_), .B0(new_n24780_), .Y(new_n24808_));
  MX2X1    g22372(.A(new_n24808_), .B(new_n5809_), .S0(pi0054), .Y(new_n24809_));
  OAI21X1  g22373(.A0(new_n24809_), .A1(new_n7552_), .B0(new_n11168_), .Y(new_n24810_));
  AOI21X1  g22374(.A0(new_n24810_), .A1(new_n3118_), .B0(new_n4980_), .Y(new_n24811_));
  OAI21X1  g22375(.A0(new_n24811_), .A1(pi0062), .B0(new_n11167_), .Y(new_n24812_));
  AOI21X1  g22376(.A0(new_n24812_), .A1(new_n3223_), .B0(new_n4977_), .Y(po0389));
  INVX1    g22377(.A(pi0230), .Y(new_n24814_));
  INVX1    g22378(.A(pi0213), .Y(new_n24815_));
  NOR2X1   g22379(.A(pi0214), .B(pi0212), .Y(new_n24816_));
  NOR2X1   g22380(.A(new_n24816_), .B(pi0211), .Y(new_n24817_));
  NOR2X1   g22381(.A(new_n24817_), .B(new_n8422_), .Y(new_n24818_));
  NOR2X1   g22382(.A(new_n24818_), .B(new_n6489_), .Y(new_n24819_));
  INVX1    g22383(.A(pi1142), .Y(new_n24820_));
  INVX1    g22384(.A(pi1143), .Y(new_n24821_));
  MX2X1    g22385(.A(new_n2439_), .B(new_n24821_), .S0(pi0211), .Y(new_n24822_));
  INVX1    g22386(.A(pi0212), .Y(new_n24823_));
  XOR2X1   g22387(.A(pi0214), .B(new_n24823_), .Y(new_n24824_));
  NOR2X1   g22388(.A(new_n24824_), .B(new_n24822_), .Y(new_n24825_));
  AND2X1   g22389(.A(pi1143), .B(new_n23173_), .Y(new_n24826_));
  AOI21X1  g22390(.A0(new_n24826_), .A1(new_n7996_), .B0(new_n24825_), .Y(new_n24827_));
  OAI22X1  g22391(.A0(new_n24827_), .A1(pi0219), .B0(new_n7963_), .B1(new_n24820_), .Y(new_n24828_));
  AND2X1   g22392(.A(new_n24828_), .B(new_n24819_), .Y(new_n24829_));
  INVX1    g22393(.A(new_n24829_), .Y(new_n24830_));
  NOR2X1   g22394(.A(new_n24822_), .B(new_n2933_), .Y(new_n24831_));
  AOI21X1  g22395(.A0(pi1142), .A1(pi0199), .B0(pi0200), .Y(new_n24832_));
  OAI21X1  g22396(.A0(new_n2439_), .A1(pi0199), .B0(new_n24832_), .Y(new_n24833_));
  AOI21X1  g22397(.A0(pi1143), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n24834_));
  INVX1    g22398(.A(new_n24834_), .Y(new_n24835_));
  AOI21X1  g22399(.A0(new_n24835_), .A1(new_n24833_), .B0(pi0299), .Y(new_n24836_));
  OR2X1    g22400(.A(new_n24821_), .B(pi0199), .Y(new_n24837_));
  AND2X1   g22401(.A(new_n24837_), .B(new_n24832_), .Y(new_n24838_));
  AND2X1   g22402(.A(new_n2933_), .B(pi0207), .Y(new_n24839_));
  INVX1    g22403(.A(new_n24839_), .Y(new_n24840_));
  AOI21X1  g22404(.A0(pi1142), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n24841_));
  OR3X1    g22405(.A(new_n24841_), .B(new_n24840_), .C(new_n24838_), .Y(new_n24842_));
  OAI21X1  g22406(.A0(new_n24836_), .A1(pi0207), .B0(new_n24842_), .Y(new_n24843_));
  AND2X1   g22407(.A(new_n22959_), .B(pi0207), .Y(new_n24844_));
  AND3X1   g22408(.A(new_n24844_), .B(new_n24835_), .C(new_n24833_), .Y(new_n24845_));
  AOI21X1  g22409(.A0(new_n24843_), .A1(pi0208), .B0(new_n24845_), .Y(new_n24846_));
  NOR2X1   g22410(.A(new_n24846_), .B(pi0299), .Y(new_n24847_));
  NOR3X1   g22411(.A(new_n24847_), .B(new_n24831_), .C(pi0214), .Y(new_n24848_));
  INVX1    g22412(.A(pi0214), .Y(new_n24849_));
  MX2X1    g22413(.A(pi1143), .B(pi1142), .S0(pi0211), .Y(new_n24850_));
  AND2X1   g22414(.A(new_n24850_), .B(pi0299), .Y(new_n24851_));
  OR2X1    g22415(.A(new_n24851_), .B(new_n24849_), .Y(new_n24852_));
  OAI21X1  g22416(.A0(new_n24852_), .A1(new_n24847_), .B0(pi0212), .Y(new_n24853_));
  NOR2X1   g22417(.A(new_n24853_), .B(new_n24848_), .Y(new_n24854_));
  NOR2X1   g22418(.A(new_n24847_), .B(pi0214), .Y(new_n24855_));
  OAI21X1  g22419(.A0(new_n24847_), .A1(new_n24831_), .B0(new_n24823_), .Y(new_n24856_));
  OAI21X1  g22420(.A0(new_n24856_), .A1(new_n24855_), .B0(new_n8422_), .Y(new_n24857_));
  OR3X1    g22421(.A(new_n24846_), .B(new_n24817_), .C(pi0299), .Y(new_n24858_));
  NAND2X1  g22422(.A(new_n24846_), .B(new_n2933_), .Y(new_n24859_));
  AND2X1   g22423(.A(new_n24820_), .B(pi0299), .Y(new_n24860_));
  NOR3X1   g22424(.A(new_n24860_), .B(new_n24816_), .C(pi0211), .Y(new_n24861_));
  AOI21X1  g22425(.A0(new_n24861_), .A1(new_n24859_), .B0(new_n8422_), .Y(new_n24862_));
  AOI21X1  g22426(.A0(new_n24862_), .A1(new_n24858_), .B0(po1038), .Y(new_n24863_));
  OAI21X1  g22427(.A0(new_n24857_), .A1(new_n24854_), .B0(new_n24863_), .Y(new_n24864_));
  NAND2X1  g22428(.A(new_n24864_), .B(new_n24830_), .Y(new_n24865_));
  INVX1    g22429(.A(pi0209), .Y(new_n24866_));
  MX2X1    g22430(.A(pi1157), .B(pi1156), .S0(pi0211), .Y(new_n24867_));
  AOI21X1  g22431(.A0(new_n24867_), .A1(pi0214), .B0(pi0212), .Y(new_n24868_));
  MX2X1    g22432(.A(new_n12555_), .B(new_n12463_), .S0(pi0211), .Y(new_n24869_));
  MX2X1    g22433(.A(new_n12463_), .B(new_n12487_), .S0(pi0211), .Y(new_n24870_));
  MX2X1    g22434(.A(new_n24870_), .B(new_n24869_), .S0(new_n24849_), .Y(new_n24871_));
  AOI21X1  g22435(.A0(new_n24871_), .A1(pi0212), .B0(new_n24868_), .Y(new_n24872_));
  NOR2X1   g22436(.A(new_n24872_), .B(pi0219), .Y(new_n24873_));
  AND2X1   g22437(.A(pi0214), .B(new_n23173_), .Y(new_n24874_));
  AOI21X1  g22438(.A0(new_n24874_), .A1(pi1155), .B0(pi0212), .Y(new_n24875_));
  AOI21X1  g22439(.A0(pi1154), .A1(new_n23173_), .B0(pi0214), .Y(new_n24876_));
  INVX1    g22440(.A(new_n7996_), .Y(new_n24877_));
  AND2X1   g22441(.A(pi1153), .B(new_n23173_), .Y(new_n24878_));
  NOR2X1   g22442(.A(new_n24878_), .B(new_n24877_), .Y(new_n24879_));
  NOR3X1   g22443(.A(new_n24879_), .B(new_n24876_), .C(new_n24875_), .Y(new_n24880_));
  OAI21X1  g22444(.A0(new_n24880_), .A1(new_n8422_), .B0(po1038), .Y(new_n24881_));
  OAI21X1  g22445(.A0(new_n24881_), .A1(new_n24873_), .B0(new_n24815_), .Y(new_n24882_));
  INVX1    g22446(.A(new_n24882_), .Y(new_n24883_));
  AND2X1   g22447(.A(pi0299), .B(new_n8422_), .Y(new_n24884_));
  NAND2X1  g22448(.A(new_n24884_), .B(new_n24872_), .Y(new_n24885_));
  AND2X1   g22449(.A(pi0214), .B(new_n24823_), .Y(new_n24886_));
  AND2X1   g22450(.A(pi1155), .B(pi0299), .Y(new_n24887_));
  OAI21X1  g22451(.A0(new_n12364_), .A1(new_n2933_), .B0(pi0214), .Y(new_n24888_));
  AND2X1   g22452(.A(pi1154), .B(pi0299), .Y(new_n24889_));
  INVX1    g22453(.A(new_n24889_), .Y(new_n24890_));
  AOI21X1  g22454(.A0(new_n24890_), .A1(new_n24849_), .B0(new_n24823_), .Y(new_n24891_));
  AOI22X1  g22455(.A0(new_n24891_), .A1(new_n24888_), .B0(new_n24887_), .B1(new_n24886_), .Y(new_n24892_));
  AND2X1   g22456(.A(pi0219), .B(new_n23173_), .Y(new_n24893_));
  INVX1    g22457(.A(new_n24893_), .Y(new_n24894_));
  OAI21X1  g22458(.A0(new_n24894_), .A1(new_n24892_), .B0(new_n24885_), .Y(new_n24895_));
  OAI21X1  g22459(.A0(new_n24895_), .A1(new_n24847_), .B0(new_n6489_), .Y(new_n24896_));
  AOI21X1  g22460(.A0(new_n24896_), .A1(new_n24883_), .B0(new_n24866_), .Y(new_n24897_));
  OAI21X1  g22461(.A0(new_n24865_), .A1(new_n24815_), .B0(new_n24897_), .Y(new_n24898_));
  AND3X1   g22462(.A(pi1155), .B(new_n7937_), .C(pi0199), .Y(new_n24899_));
  AOI21X1  g22463(.A0(new_n24899_), .A1(new_n2933_), .B0(pi1156), .Y(new_n24900_));
  INVX1    g22464(.A(new_n24900_), .Y(new_n24901_));
  OR2X1    g22465(.A(pi1155), .B(pi0200), .Y(new_n24902_));
  XOR2X1   g22466(.A(pi0200), .B(pi0199), .Y(new_n24903_));
  AND2X1   g22467(.A(new_n24903_), .B(new_n2933_), .Y(new_n24904_));
  NAND4X1  g22468(.A(new_n24904_), .B(new_n24902_), .C(new_n24901_), .D(pi0207), .Y(new_n24905_));
  AND2X1   g22469(.A(new_n24905_), .B(new_n22959_), .Y(new_n24906_));
  AOI21X1  g22470(.A0(pi0200), .A1(pi0199), .B0(pi0299), .Y(new_n24907_));
  OR2X1    g22471(.A(new_n24907_), .B(new_n12364_), .Y(new_n24908_));
  AND2X1   g22472(.A(new_n24908_), .B(pi1154), .Y(new_n24909_));
  AND3X1   g22473(.A(new_n8423_), .B(pi1155), .C(new_n7937_), .Y(new_n24910_));
  INVX1    g22474(.A(new_n24903_), .Y(new_n24911_));
  NOR2X1   g22475(.A(new_n8423_), .B(pi1153), .Y(new_n24912_));
  NOR3X1   g22476(.A(new_n24912_), .B(new_n24911_), .C(new_n12487_), .Y(new_n24913_));
  NOR2X1   g22477(.A(new_n24913_), .B(new_n24910_), .Y(new_n24914_));
  INVX1    g22478(.A(new_n24914_), .Y(new_n24915_));
  NOR2X1   g22479(.A(pi0299), .B(pi0200), .Y(new_n24916_));
  INVX1    g22480(.A(new_n24916_), .Y(new_n24917_));
  AND2X1   g22481(.A(new_n12364_), .B(pi0199), .Y(new_n24918_));
  OAI21X1  g22482(.A0(pi1155), .A1(pi0199), .B0(new_n12487_), .Y(new_n24919_));
  NOR3X1   g22483(.A(new_n24919_), .B(new_n24918_), .C(new_n24917_), .Y(new_n24920_));
  AOI21X1  g22484(.A0(new_n24915_), .A1(new_n24909_), .B0(new_n24920_), .Y(new_n24921_));
  NOR4X1   g22485(.A(new_n12463_), .B(pi0299), .C(new_n7937_), .D(pi0199), .Y(new_n24922_));
  NOR2X1   g22486(.A(new_n24922_), .B(pi1154), .Y(new_n24923_));
  INVX1    g22487(.A(new_n24923_), .Y(new_n24924_));
  OAI21X1  g22488(.A0(new_n12463_), .A1(pi0199), .B0(pi0200), .Y(new_n24925_));
  AND2X1   g22489(.A(new_n24925_), .B(new_n9445_), .Y(new_n24926_));
  OAI21X1  g22490(.A0(pi1155), .A1(new_n7937_), .B0(new_n8423_), .Y(new_n24927_));
  NOR2X1   g22491(.A(new_n24927_), .B(new_n12555_), .Y(new_n24928_));
  AOI21X1  g22492(.A0(new_n24926_), .A1(new_n24924_), .B0(new_n24928_), .Y(new_n24929_));
  MX2X1    g22493(.A(new_n24929_), .B(new_n24921_), .S0(pi0207), .Y(new_n24930_));
  AOI21X1  g22494(.A0(new_n24930_), .A1(pi0208), .B0(new_n24906_), .Y(new_n24931_));
  OR2X1    g22495(.A(new_n24931_), .B(pi1157), .Y(new_n24932_));
  INVX1    g22496(.A(new_n24907_), .Y(new_n24933_));
  AND2X1   g22497(.A(new_n12463_), .B(pi0199), .Y(new_n24934_));
  NOR3X1   g22498(.A(new_n24934_), .B(new_n24933_), .C(new_n12555_), .Y(new_n24935_));
  NOR3X1   g22499(.A(new_n24934_), .B(new_n24917_), .C(pi1156), .Y(new_n24936_));
  NOR2X1   g22500(.A(new_n24936_), .B(new_n24935_), .Y(new_n24937_));
  NOR2X1   g22501(.A(new_n24937_), .B(new_n22660_), .Y(new_n24938_));
  NOR2X1   g22502(.A(new_n24938_), .B(pi0208), .Y(new_n24939_));
  AOI21X1  g22503(.A0(new_n24930_), .A1(pi0208), .B0(new_n24939_), .Y(new_n24940_));
  OAI21X1  g22504(.A0(new_n24940_), .A1(new_n12578_), .B0(new_n24932_), .Y(new_n24941_));
  AND2X1   g22505(.A(new_n24941_), .B(pi0211), .Y(new_n24942_));
  AOI21X1  g22506(.A0(new_n24941_), .A1(new_n24849_), .B0(pi0212), .Y(new_n24943_));
  INVX1    g22507(.A(new_n24874_), .Y(new_n24944_));
  NOR3X1   g22508(.A(new_n24902_), .B(pi0299), .C(new_n7871_), .Y(new_n24945_));
  AND2X1   g22509(.A(new_n2933_), .B(pi0200), .Y(new_n24946_));
  MX2X1    g22510(.A(new_n24946_), .B(new_n9445_), .S0(new_n12364_), .Y(new_n24947_));
  INVX1    g22511(.A(new_n24947_), .Y(new_n24948_));
  AOI22X1  g22512(.A0(new_n24948_), .A1(pi1155), .B0(new_n24945_), .B1(pi1153), .Y(new_n24949_));
  AND2X1   g22513(.A(new_n2933_), .B(pi0199), .Y(new_n24950_));
  INVX1    g22514(.A(new_n24950_), .Y(new_n24951_));
  NOR3X1   g22515(.A(new_n24918_), .B(new_n24911_), .C(pi0299), .Y(new_n24952_));
  AOI21X1  g22516(.A0(new_n24951_), .A1(pi1155), .B0(new_n24952_), .Y(new_n24953_));
  MX2X1    g22517(.A(new_n24953_), .B(new_n24949_), .S0(new_n12487_), .Y(new_n24954_));
  INVX1    g22518(.A(new_n24887_), .Y(new_n24955_));
  AND3X1   g22519(.A(new_n24929_), .B(new_n24955_), .C(new_n22660_), .Y(new_n24956_));
  OR2X1    g22520(.A(new_n24956_), .B(new_n22959_), .Y(new_n24957_));
  AOI21X1  g22521(.A0(new_n24954_), .A1(pi0207), .B0(new_n24957_), .Y(new_n24958_));
  AOI21X1  g22522(.A0(new_n2933_), .A1(pi0200), .B0(new_n12463_), .Y(new_n24959_));
  OAI21X1  g22523(.A0(new_n24959_), .A1(new_n8423_), .B0(pi1156), .Y(new_n24960_));
  AOI21X1  g22524(.A0(new_n7937_), .A1(pi0199), .B0(pi0299), .Y(new_n24961_));
  AOI21X1  g22525(.A0(new_n2933_), .A1(pi0200), .B0(pi1156), .Y(new_n24962_));
  OAI21X1  g22526(.A0(new_n24961_), .A1(pi1155), .B0(new_n24962_), .Y(new_n24963_));
  AND2X1   g22527(.A(new_n24963_), .B(new_n24960_), .Y(new_n24964_));
  AOI21X1  g22528(.A0(new_n24955_), .A1(new_n22660_), .B0(pi0208), .Y(new_n24965_));
  NAND2X1  g22529(.A(new_n24965_), .B(pi1157), .Y(new_n24966_));
  AOI21X1  g22530(.A0(new_n24964_), .A1(pi0207), .B0(new_n24966_), .Y(new_n24967_));
  INVX1    g22531(.A(new_n24965_), .Y(new_n24968_));
  NOR3X1   g22532(.A(new_n24899_), .B(pi1156), .C(pi0299), .Y(new_n24969_));
  NOR2X1   g22533(.A(new_n24903_), .B(pi0299), .Y(new_n24970_));
  NOR2X1   g22534(.A(new_n8423_), .B(pi1155), .Y(new_n24971_));
  NOR4X1   g22535(.A(new_n24971_), .B(new_n24970_), .C(new_n24969_), .D(new_n24968_), .Y(new_n24972_));
  OR4X1    g22536(.A(new_n24972_), .B(new_n24967_), .C(new_n24958_), .D(new_n24944_), .Y(new_n24973_));
  NOR2X1   g22537(.A(pi0214), .B(pi0211), .Y(new_n24974_));
  MX2X1    g22538(.A(new_n24970_), .B(new_n24961_), .S0(new_n12463_), .Y(new_n24975_));
  OAI21X1  g22539(.A0(new_n24975_), .A1(new_n12487_), .B0(new_n24929_), .Y(new_n24976_));
  AOI21X1  g22540(.A0(new_n24953_), .A1(new_n2933_), .B0(new_n12487_), .Y(new_n24977_));
  OR2X1    g22541(.A(new_n24977_), .B(new_n24920_), .Y(new_n24978_));
  MX2X1    g22542(.A(new_n24978_), .B(new_n24976_), .S0(new_n22660_), .Y(new_n24979_));
  NAND2X1  g22543(.A(new_n24979_), .B(pi0208), .Y(new_n24980_));
  MX2X1    g22544(.A(new_n24946_), .B(new_n9445_), .S0(new_n12463_), .Y(new_n24981_));
  AOI21X1  g22545(.A0(pi1155), .A1(new_n7937_), .B0(new_n24951_), .Y(new_n24982_));
  MX2X1    g22546(.A(new_n24982_), .B(new_n24981_), .S0(new_n12555_), .Y(new_n24983_));
  NOR2X1   g22547(.A(pi0299), .B(pi0207), .Y(new_n24984_));
  NOR2X1   g22548(.A(new_n24984_), .B(pi0208), .Y(new_n24985_));
  INVX1    g22549(.A(new_n24985_), .Y(new_n24986_));
  AOI21X1  g22550(.A0(new_n24983_), .A1(pi0207), .B0(new_n24986_), .Y(new_n24987_));
  AOI21X1  g22551(.A0(new_n12487_), .A1(pi0299), .B0(new_n12578_), .Y(new_n24988_));
  AOI21X1  g22552(.A0(new_n24905_), .A1(new_n24890_), .B0(pi0208), .Y(new_n24989_));
  AOI22X1  g22553(.A0(new_n24989_), .A1(new_n12578_), .B0(new_n24988_), .B1(new_n24987_), .Y(new_n24990_));
  NAND3X1  g22554(.A(new_n24990_), .B(new_n24980_), .C(new_n24974_), .Y(new_n24991_));
  INVX1    g22555(.A(new_n24961_), .Y(new_n24992_));
  AOI21X1  g22556(.A0(new_n24992_), .A1(pi1153), .B0(new_n24915_), .Y(new_n24993_));
  NOR2X1   g22557(.A(new_n24993_), .B(new_n22660_), .Y(new_n24994_));
  OR2X1    g22558(.A(new_n24975_), .B(new_n12487_), .Y(new_n24995_));
  MX2X1    g22559(.A(new_n24950_), .B(new_n9445_), .S0(new_n12463_), .Y(new_n24996_));
  OR2X1    g22560(.A(new_n24996_), .B(new_n12555_), .Y(new_n24997_));
  AOI21X1  g22561(.A0(pi0200), .A1(new_n7871_), .B0(pi0299), .Y(new_n24998_));
  MX2X1    g22562(.A(new_n24998_), .B(new_n2933_), .S0(new_n12463_), .Y(new_n24999_));
  AND3X1   g22563(.A(new_n24999_), .B(new_n24997_), .C(new_n24995_), .Y(new_n25000_));
  AND2X1   g22564(.A(new_n12364_), .B(pi0299), .Y(new_n25001_));
  NOR3X1   g22565(.A(new_n25001_), .B(new_n25000_), .C(pi0207), .Y(new_n25002_));
  OAI21X1  g22566(.A0(new_n25002_), .A1(new_n24994_), .B0(pi0208), .Y(new_n25003_));
  AND2X1   g22567(.A(pi0200), .B(new_n7871_), .Y(new_n25004_));
  OR4X1    g22568(.A(new_n24899_), .B(new_n25004_), .C(new_n12555_), .D(pi0299), .Y(new_n25005_));
  AND3X1   g22569(.A(new_n25005_), .B(new_n24901_), .C(pi0207), .Y(new_n25006_));
  OAI21X1  g22570(.A0(new_n25006_), .A1(pi0299), .B0(new_n22959_), .Y(new_n25007_));
  NAND2X1  g22571(.A(new_n25007_), .B(new_n12578_), .Y(new_n25008_));
  NOR2X1   g22572(.A(new_n24987_), .B(new_n12578_), .Y(new_n25009_));
  NOR2X1   g22573(.A(new_n25009_), .B(new_n25001_), .Y(new_n25010_));
  AOI21X1  g22574(.A0(new_n25010_), .A1(new_n25008_), .B0(new_n24944_), .Y(new_n25011_));
  AOI21X1  g22575(.A0(new_n25011_), .A1(new_n25003_), .B0(new_n24823_), .Y(new_n25012_));
  AOI22X1  g22576(.A0(new_n25012_), .A1(new_n24991_), .B0(new_n24973_), .B1(new_n24943_), .Y(new_n25013_));
  OAI21X1  g22577(.A0(new_n25013_), .A1(new_n24942_), .B0(pi0219), .Y(new_n25014_));
  AND2X1   g22578(.A(new_n25000_), .B(new_n22660_), .Y(new_n25015_));
  AND2X1   g22579(.A(new_n24993_), .B(new_n24839_), .Y(new_n25016_));
  OR3X1    g22580(.A(new_n25016_), .B(new_n25015_), .C(new_n22959_), .Y(new_n25017_));
  AOI21X1  g22581(.A0(new_n25017_), .A1(new_n25009_), .B0(pi0211), .Y(new_n25018_));
  AND2X1   g22582(.A(new_n25018_), .B(new_n24932_), .Y(new_n25019_));
  OAI21X1  g22583(.A0(new_n24922_), .A1(pi1154), .B0(new_n24926_), .Y(new_n25020_));
  AND2X1   g22584(.A(new_n24997_), .B(new_n25020_), .Y(new_n25021_));
  AND2X1   g22585(.A(pi1156), .B(pi0299), .Y(new_n25022_));
  INVX1    g22586(.A(new_n25022_), .Y(new_n25023_));
  MX2X1    g22587(.A(new_n25023_), .B(new_n25021_), .S0(new_n22660_), .Y(new_n25024_));
  OAI21X1  g22588(.A0(new_n24921_), .A1(new_n22660_), .B0(new_n25024_), .Y(new_n25025_));
  AND2X1   g22589(.A(pi1157), .B(new_n22959_), .Y(new_n25026_));
  OAI21X1  g22590(.A0(new_n25022_), .A1(new_n24938_), .B0(new_n25026_), .Y(new_n25027_));
  OAI21X1  g22591(.A0(new_n25007_), .A1(new_n24900_), .B0(new_n25027_), .Y(new_n25028_));
  AOI21X1  g22592(.A0(new_n25025_), .A1(pi0208), .B0(new_n25028_), .Y(new_n25029_));
  OAI21X1  g22593(.A0(new_n25029_), .A1(new_n23173_), .B0(pi0214), .Y(new_n25030_));
  OAI21X1  g22594(.A0(new_n25030_), .A1(new_n25019_), .B0(new_n24943_), .Y(new_n25031_));
  AND2X1   g22595(.A(pi0214), .B(pi0211), .Y(new_n25032_));
  INVX1    g22596(.A(new_n25032_), .Y(new_n25033_));
  AOI21X1  g22597(.A0(new_n24990_), .A1(new_n24980_), .B0(new_n25033_), .Y(new_n25034_));
  OR3X1    g22598(.A(new_n24972_), .B(new_n24967_), .C(new_n24958_), .Y(new_n25035_));
  XOR2X1   g22599(.A(pi0214), .B(pi0211), .Y(new_n25036_));
  AND2X1   g22600(.A(new_n25036_), .B(new_n25035_), .Y(new_n25037_));
  INVX1    g22601(.A(new_n24974_), .Y(new_n25038_));
  NOR2X1   g22602(.A(new_n25029_), .B(new_n25038_), .Y(new_n25039_));
  OR3X1    g22603(.A(new_n25039_), .B(new_n25037_), .C(new_n25034_), .Y(new_n25040_));
  AOI21X1  g22604(.A0(new_n25040_), .A1(pi0212), .B0(pi0219), .Y(new_n25041_));
  AOI21X1  g22605(.A0(new_n25041_), .A1(new_n25031_), .B0(po1038), .Y(new_n25042_));
  AOI21X1  g22606(.A0(new_n25042_), .A1(new_n25014_), .B0(new_n24882_), .Y(new_n25043_));
  AND2X1   g22607(.A(new_n7996_), .B(new_n23173_), .Y(new_n25044_));
  NAND2X1  g22608(.A(new_n24921_), .B(pi0207), .Y(new_n25045_));
  AND2X1   g22609(.A(pi1143), .B(pi0299), .Y(new_n25046_));
  OAI21X1  g22610(.A0(new_n24903_), .A1(pi0299), .B0(pi1155), .Y(new_n25047_));
  AND2X1   g22611(.A(new_n24821_), .B(pi0299), .Y(new_n25048_));
  AND2X1   g22612(.A(new_n25046_), .B(new_n12463_), .Y(new_n25049_));
  NOR3X1   g22613(.A(new_n25049_), .B(new_n24945_), .C(new_n12487_), .Y(new_n25050_));
  OAI21X1  g22614(.A0(new_n25048_), .A1(new_n25047_), .B0(new_n25050_), .Y(new_n25051_));
  INVX1    g22615(.A(new_n25046_), .Y(new_n25052_));
  AOI21X1  g22616(.A0(new_n25052_), .A1(new_n24923_), .B0(pi1156), .Y(new_n25053_));
  OAI21X1  g22617(.A0(new_n25048_), .A1(new_n24996_), .B0(new_n12487_), .Y(new_n25054_));
  AOI21X1  g22618(.A0(new_n24925_), .A1(new_n2933_), .B0(new_n12487_), .Y(new_n25055_));
  AOI21X1  g22619(.A0(new_n25055_), .A1(new_n25052_), .B0(new_n12555_), .Y(new_n25056_));
  AOI22X1  g22620(.A0(new_n25056_), .A1(new_n25054_), .B0(new_n25053_), .B1(new_n25051_), .Y(new_n25057_));
  AOI21X1  g22621(.A0(new_n25057_), .A1(new_n22660_), .B0(new_n22959_), .Y(new_n25058_));
  OAI21X1  g22622(.A0(new_n25046_), .A1(new_n25045_), .B0(new_n25058_), .Y(new_n25059_));
  NOR3X1   g22623(.A(new_n25048_), .B(new_n25007_), .C(pi1157), .Y(new_n25060_));
  NOR2X1   g22624(.A(new_n9445_), .B(pi1155), .Y(new_n25061_));
  NOR3X1   g22625(.A(new_n25061_), .B(new_n24959_), .C(new_n24935_), .Y(new_n25062_));
  OAI21X1  g22626(.A0(pi1143), .A1(new_n2933_), .B0(pi0207), .Y(new_n25063_));
  OAI21X1  g22627(.A0(new_n25063_), .A1(new_n25062_), .B0(new_n25052_), .Y(new_n25064_));
  AOI21X1  g22628(.A0(new_n25064_), .A1(new_n25026_), .B0(new_n25060_), .Y(new_n25065_));
  AND3X1   g22629(.A(new_n25065_), .B(new_n25059_), .C(new_n25044_), .Y(new_n25066_));
  AOI21X1  g22630(.A0(new_n25065_), .A1(new_n25059_), .B0(new_n23173_), .Y(new_n25067_));
  AND2X1   g22631(.A(pi1144), .B(pi0299), .Y(new_n25068_));
  AND2X1   g22632(.A(new_n2439_), .B(pi0299), .Y(new_n25069_));
  AND2X1   g22633(.A(new_n25068_), .B(new_n12463_), .Y(new_n25070_));
  NOR3X1   g22634(.A(new_n25070_), .B(new_n24945_), .C(new_n12487_), .Y(new_n25071_));
  OAI21X1  g22635(.A0(new_n25069_), .A1(new_n25047_), .B0(new_n25071_), .Y(new_n25072_));
  INVX1    g22636(.A(new_n25068_), .Y(new_n25073_));
  AOI21X1  g22637(.A0(new_n25073_), .A1(new_n24923_), .B0(pi1156), .Y(new_n25074_));
  OAI21X1  g22638(.A0(new_n25069_), .A1(new_n24996_), .B0(new_n12487_), .Y(new_n25075_));
  AOI21X1  g22639(.A0(new_n25073_), .A1(new_n25055_), .B0(new_n12555_), .Y(new_n25076_));
  AOI22X1  g22640(.A0(new_n25076_), .A1(new_n25075_), .B0(new_n25074_), .B1(new_n25072_), .Y(new_n25077_));
  AOI21X1  g22641(.A0(new_n25077_), .A1(new_n22660_), .B0(new_n22959_), .Y(new_n25078_));
  OAI21X1  g22642(.A0(new_n25068_), .A1(new_n25045_), .B0(new_n25078_), .Y(new_n25079_));
  NOR3X1   g22643(.A(new_n25069_), .B(new_n25007_), .C(pi1157), .Y(new_n25080_));
  OAI21X1  g22644(.A0(pi1144), .A1(new_n2933_), .B0(pi0207), .Y(new_n25081_));
  OAI21X1  g22645(.A0(new_n25081_), .A1(new_n25062_), .B0(new_n25073_), .Y(new_n25082_));
  AOI21X1  g22646(.A0(new_n25082_), .A1(new_n25026_), .B0(new_n25080_), .Y(new_n25083_));
  AOI21X1  g22647(.A0(new_n25083_), .A1(new_n25079_), .B0(pi0211), .Y(new_n25084_));
  XOR2X1   g22648(.A(pi0214), .B(pi0212), .Y(new_n25085_));
  INVX1    g22649(.A(new_n25085_), .Y(new_n25086_));
  NOR3X1   g22650(.A(new_n25086_), .B(new_n25084_), .C(new_n25067_), .Y(new_n25087_));
  OAI21X1  g22651(.A0(new_n25087_), .A1(new_n25066_), .B0(new_n8422_), .Y(new_n25088_));
  OAI22X1  g22652(.A0(new_n8422_), .A1(new_n23173_), .B0(pi0214), .B1(pi0212), .Y(new_n25089_));
  NAND2X1  g22653(.A(new_n25089_), .B(new_n24941_), .Y(new_n25090_));
  OAI22X1  g22654(.A0(new_n24987_), .A1(new_n12578_), .B0(pi1142), .B1(new_n2933_), .Y(new_n25091_));
  AOI21X1  g22655(.A0(new_n25007_), .A1(new_n12578_), .B0(new_n25091_), .Y(new_n25092_));
  AOI21X1  g22656(.A0(pi1142), .A1(pi0299), .B0(new_n22660_), .Y(new_n25093_));
  OAI21X1  g22657(.A0(new_n24954_), .A1(pi0299), .B0(new_n25093_), .Y(new_n25094_));
  AND2X1   g22658(.A(new_n24997_), .B(new_n24995_), .Y(new_n25095_));
  INVX1    g22659(.A(new_n24922_), .Y(new_n25096_));
  OAI21X1  g22660(.A0(new_n24820_), .A1(new_n2933_), .B0(new_n25096_), .Y(new_n25097_));
  NOR2X1   g22661(.A(pi1156), .B(pi1154), .Y(new_n25098_));
  AOI21X1  g22662(.A0(new_n25098_), .A1(new_n25097_), .B0(pi0207), .Y(new_n25099_));
  OAI21X1  g22663(.A0(new_n25095_), .A1(new_n24860_), .B0(new_n25099_), .Y(new_n25100_));
  AND3X1   g22664(.A(new_n25100_), .B(new_n25094_), .C(pi0208), .Y(new_n25101_));
  NOR4X1   g22665(.A(new_n25101_), .B(new_n25092_), .C(new_n25089_), .D(new_n7963_), .Y(new_n25102_));
  NOR2X1   g22666(.A(new_n25102_), .B(po1038), .Y(new_n25103_));
  AND3X1   g22667(.A(new_n25103_), .B(new_n25090_), .C(new_n25088_), .Y(new_n25104_));
  OR2X1    g22668(.A(new_n24829_), .B(new_n24815_), .Y(new_n25105_));
  OAI21X1  g22669(.A0(new_n25105_), .A1(new_n25104_), .B0(new_n24866_), .Y(new_n25106_));
  OAI21X1  g22670(.A0(new_n25106_), .A1(new_n25043_), .B0(new_n24898_), .Y(new_n25107_));
  MX2X1    g22671(.A(new_n25107_), .B(new_n22655_), .S0(new_n24814_), .Y(po0390));
  NOR2X1   g22672(.A(new_n24816_), .B(pi0219), .Y(new_n25109_));
  INVX1    g22673(.A(new_n25109_), .Y(new_n25110_));
  MX2X1    g22674(.A(new_n12487_), .B(new_n12364_), .S0(pi0211), .Y(new_n25111_));
  AND2X1   g22675(.A(new_n25111_), .B(new_n24877_), .Y(new_n25112_));
  NOR3X1   g22676(.A(new_n25112_), .B(new_n25110_), .C(new_n24879_), .Y(new_n25113_));
  AOI21X1  g22677(.A0(new_n25113_), .A1(po1038), .B0(pi1152), .Y(new_n25114_));
  XOR2X1   g22678(.A(pi0208), .B(pi0207), .Y(new_n25115_));
  INVX1    g22679(.A(new_n25115_), .Y(new_n25116_));
  INVX1    g22680(.A(new_n24910_), .Y(new_n25117_));
  OAI21X1  g22681(.A0(new_n24902_), .A1(pi0199), .B0(new_n24907_), .Y(new_n25118_));
  AOI21X1  g22682(.A0(new_n25117_), .A1(new_n12487_), .B0(new_n25118_), .Y(new_n25119_));
  AND2X1   g22683(.A(new_n25119_), .B(pi0207), .Y(new_n25120_));
  INVX1    g22684(.A(new_n25120_), .Y(new_n25121_));
  AOI22X1  g22685(.A0(new_n25121_), .A1(new_n25116_), .B0(new_n24929_), .B1(new_n7827_), .Y(new_n25122_));
  INVX1    g22686(.A(new_n25122_), .Y(new_n25123_));
  AOI21X1  g22687(.A0(new_n25123_), .A1(new_n24849_), .B0(pi0212), .Y(new_n25124_));
  INVX1    g22688(.A(new_n25124_), .Y(new_n25125_));
  AND2X1   g22689(.A(new_n24889_), .B(new_n22660_), .Y(new_n25126_));
  AOI21X1  g22690(.A0(new_n24995_), .A1(new_n24929_), .B0(new_n22660_), .Y(new_n25127_));
  OR2X1    g22691(.A(new_n25127_), .B(new_n25126_), .Y(new_n25128_));
  AND2X1   g22692(.A(new_n25128_), .B(new_n22959_), .Y(new_n25129_));
  AND2X1   g22693(.A(pi0200), .B(pi0199), .Y(new_n25130_));
  AOI21X1  g22694(.A0(new_n8055_), .A1(new_n12463_), .B0(new_n25130_), .Y(new_n25131_));
  NOR2X1   g22695(.A(new_n25131_), .B(pi0299), .Y(new_n25132_));
  AOI21X1  g22696(.A0(new_n25117_), .A1(new_n12487_), .B0(new_n25132_), .Y(new_n25133_));
  MX2X1    g22697(.A(new_n25133_), .B(new_n24976_), .S0(new_n22660_), .Y(new_n25134_));
  AOI21X1  g22698(.A0(new_n25134_), .A1(pi0208), .B0(new_n25129_), .Y(new_n25135_));
  INVX1    g22699(.A(new_n25015_), .Y(new_n25136_));
  AND3X1   g22700(.A(new_n24999_), .B(new_n25095_), .C(pi0207), .Y(new_n25137_));
  INVX1    g22701(.A(new_n25137_), .Y(new_n25138_));
  OR2X1    g22702(.A(new_n25133_), .B(new_n24840_), .Y(new_n25139_));
  AND2X1   g22703(.A(new_n25139_), .B(pi0208), .Y(new_n25140_));
  AOI22X1  g22704(.A0(new_n25140_), .A1(new_n25136_), .B0(new_n25138_), .B1(new_n24985_), .Y(new_n25141_));
  OR2X1    g22705(.A(new_n25141_), .B(new_n25001_), .Y(new_n25142_));
  MX2X1    g22706(.A(new_n25142_), .B(new_n25135_), .S0(new_n23173_), .Y(new_n25143_));
  AOI21X1  g22707(.A0(new_n25143_), .A1(pi0214), .B0(new_n25125_), .Y(new_n25144_));
  OR2X1    g22708(.A(new_n25144_), .B(pi0219), .Y(new_n25145_));
  OAI21X1  g22709(.A0(new_n25141_), .A1(new_n25001_), .B0(new_n23173_), .Y(new_n25146_));
  NAND2X1  g22710(.A(new_n25146_), .B(pi0214), .Y(new_n25147_));
  NOR2X1   g22711(.A(new_n25122_), .B(new_n23173_), .Y(new_n25148_));
  OAI22X1  g22712(.A0(new_n25148_), .A1(new_n25147_), .B0(new_n25143_), .B1(pi0214), .Y(new_n25149_));
  AOI21X1  g22713(.A0(new_n25149_), .A1(pi0212), .B0(new_n25145_), .Y(new_n25150_));
  OAI21X1  g22714(.A0(new_n25122_), .A1(new_n8422_), .B0(new_n6489_), .Y(new_n25151_));
  OAI21X1  g22715(.A0(new_n25151_), .A1(new_n25150_), .B0(new_n25114_), .Y(new_n25152_));
  INVX1    g22716(.A(pi1152), .Y(new_n25153_));
  NOR2X1   g22717(.A(new_n24876_), .B(new_n24874_), .Y(new_n25154_));
  AOI21X1  g22718(.A0(new_n25038_), .A1(pi1153), .B0(new_n25154_), .Y(new_n25155_));
  INVX1    g22719(.A(new_n25111_), .Y(new_n25156_));
  AOI21X1  g22720(.A0(new_n25156_), .A1(new_n24886_), .B0(pi0219), .Y(new_n25157_));
  OAI21X1  g22721(.A0(new_n25155_), .A1(new_n24823_), .B0(new_n25157_), .Y(new_n25158_));
  AOI21X1  g22722(.A0(new_n25158_), .A1(new_n24819_), .B0(new_n25153_), .Y(new_n25159_));
  OAI22X1  g22723(.A0(new_n25147_), .A1(new_n25141_), .B0(new_n25143_), .B1(pi0214), .Y(new_n25160_));
  AND2X1   g22724(.A(new_n25160_), .B(pi0212), .Y(new_n25161_));
  INVX1    g22725(.A(new_n24817_), .Y(new_n25162_));
  AOI21X1  g22726(.A0(new_n25122_), .A1(new_n25162_), .B0(new_n8422_), .Y(new_n25163_));
  OAI21X1  g22727(.A0(new_n25141_), .A1(new_n25162_), .B0(new_n25163_), .Y(new_n25164_));
  AND2X1   g22728(.A(new_n25164_), .B(new_n6489_), .Y(new_n25165_));
  OAI21X1  g22729(.A0(new_n25161_), .A1(new_n25145_), .B0(new_n25165_), .Y(new_n25166_));
  AOI21X1  g22730(.A0(new_n25166_), .A1(new_n25159_), .B0(pi0213), .Y(new_n25167_));
  OR2X1    g22731(.A(new_n25021_), .B(new_n22660_), .Y(new_n25168_));
  AOI21X1  g22732(.A0(new_n25168_), .A1(new_n25023_), .B0(pi0208), .Y(new_n25169_));
  AOI21X1  g22733(.A0(new_n25121_), .A1(new_n25024_), .B0(new_n22959_), .Y(new_n25170_));
  OR2X1    g22734(.A(new_n25170_), .B(new_n25169_), .Y(new_n25171_));
  AND2X1   g22735(.A(new_n24929_), .B(new_n24955_), .Y(new_n25172_));
  OR2X1    g22736(.A(new_n24887_), .B(new_n22660_), .Y(new_n25173_));
  OAI21X1  g22737(.A0(new_n25173_), .A1(new_n25119_), .B0(pi0208), .Y(new_n25174_));
  OAI22X1  g22738(.A0(new_n25174_), .A1(new_n24956_), .B0(new_n25172_), .B1(new_n24968_), .Y(new_n25175_));
  MX2X1    g22739(.A(new_n25175_), .B(new_n25171_), .S0(new_n23173_), .Y(new_n25176_));
  OAI21X1  g22740(.A0(new_n25176_), .A1(new_n24849_), .B0(new_n25124_), .Y(new_n25177_));
  OR2X1    g22741(.A(new_n25176_), .B(pi0214), .Y(new_n25178_));
  AOI21X1  g22742(.A0(new_n25175_), .A1(new_n23173_), .B0(new_n24849_), .Y(new_n25179_));
  OAI21X1  g22743(.A0(new_n25135_), .A1(new_n23173_), .B0(new_n25179_), .Y(new_n25180_));
  NAND3X1  g22744(.A(new_n25180_), .B(new_n25178_), .C(pi0212), .Y(new_n25181_));
  AND3X1   g22745(.A(new_n25181_), .B(new_n25177_), .C(new_n8422_), .Y(new_n25182_));
  INVX1    g22746(.A(new_n25163_), .Y(new_n25183_));
  NOR3X1   g22747(.A(new_n25135_), .B(new_n24816_), .C(pi0211), .Y(new_n25184_));
  OAI21X1  g22748(.A0(new_n25184_), .A1(new_n25183_), .B0(new_n23202_), .Y(new_n25185_));
  OAI21X1  g22749(.A0(new_n25185_), .A1(new_n25182_), .B0(pi0209), .Y(new_n25186_));
  AOI21X1  g22750(.A0(new_n25167_), .A1(new_n25152_), .B0(new_n25186_), .Y(new_n25187_));
  INVX1    g22751(.A(new_n24816_), .Y(new_n25188_));
  NOR4X1   g22752(.A(new_n12364_), .B(pi0299), .C(new_n7937_), .D(pi0199), .Y(new_n25189_));
  NOR2X1   g22753(.A(new_n25189_), .B(pi1154), .Y(new_n25190_));
  OR3X1    g22754(.A(new_n12487_), .B(pi0299), .C(new_n7937_), .Y(new_n25191_));
  AOI21X1  g22755(.A0(pi1153), .A1(new_n7871_), .B0(new_n25191_), .Y(new_n25192_));
  OAI21X1  g22756(.A0(new_n25192_), .A1(new_n25190_), .B0(new_n24961_), .Y(new_n25193_));
  OR2X1    g22757(.A(new_n25193_), .B(pi0207), .Y(new_n25194_));
  AND2X1   g22758(.A(new_n7937_), .B(pi0199), .Y(new_n25195_));
  INVX1    g22759(.A(new_n25195_), .Y(new_n25196_));
  NOR2X1   g22760(.A(pi1153), .B(pi0200), .Y(new_n25197_));
  OR2X1    g22761(.A(new_n25197_), .B(pi0199), .Y(new_n25198_));
  AND2X1   g22762(.A(new_n25198_), .B(new_n2933_), .Y(new_n25199_));
  AND3X1   g22763(.A(new_n25199_), .B(new_n25196_), .C(pi0207), .Y(new_n25200_));
  NOR2X1   g22764(.A(new_n25200_), .B(new_n22959_), .Y(new_n25201_));
  AOI22X1  g22765(.A0(new_n25201_), .A1(new_n25194_), .B0(new_n25193_), .B1(new_n24985_), .Y(new_n25202_));
  INVX1    g22766(.A(new_n25202_), .Y(new_n25203_));
  NOR3X1   g22767(.A(pi0299), .B(pi0200), .C(pi0199), .Y(new_n25204_));
  OR2X1    g22768(.A(new_n25204_), .B(pi1153), .Y(new_n25205_));
  AND3X1   g22769(.A(new_n25205_), .B(new_n24908_), .C(pi1154), .Y(new_n25206_));
  NOR2X1   g22770(.A(pi1153), .B(pi0199), .Y(new_n25207_));
  NOR4X1   g22771(.A(new_n25207_), .B(new_n25130_), .C(new_n8055_), .D(pi0299), .Y(new_n25208_));
  NOR2X1   g22772(.A(new_n25208_), .B(new_n25206_), .Y(new_n25209_));
  INVX1    g22773(.A(new_n25209_), .Y(new_n25210_));
  NOR2X1   g22774(.A(pi0208), .B(pi0207), .Y(new_n25211_));
  OR3X1    g22775(.A(pi1153), .B(pi0200), .C(pi0199), .Y(new_n25212_));
  AND2X1   g22776(.A(new_n25212_), .B(new_n24907_), .Y(new_n25213_));
  INVX1    g22777(.A(new_n25213_), .Y(new_n25214_));
  AOI21X1  g22778(.A0(new_n25214_), .A1(new_n7826_), .B0(new_n25211_), .Y(new_n25215_));
  OAI21X1  g22779(.A0(new_n25210_), .A1(new_n7826_), .B0(new_n25215_), .Y(new_n25216_));
  INVX1    g22780(.A(new_n25216_), .Y(new_n25217_));
  MX2X1    g22781(.A(new_n25217_), .B(new_n25203_), .S0(new_n23173_), .Y(new_n25218_));
  OAI21X1  g22782(.A0(new_n25216_), .A1(new_n25188_), .B0(pi0219), .Y(new_n25219_));
  AOI21X1  g22783(.A0(new_n25218_), .A1(new_n25188_), .B0(new_n25219_), .Y(new_n25220_));
  NOR2X1   g22784(.A(new_n25220_), .B(po1038), .Y(new_n25221_));
  OAI21X1  g22785(.A0(new_n25208_), .A1(new_n25206_), .B0(pi0207), .Y(new_n25222_));
  NAND2X1  g22786(.A(new_n25222_), .B(new_n24890_), .Y(new_n25223_));
  AND2X1   g22787(.A(new_n12487_), .B(pi0299), .Y(new_n25224_));
  INVX1    g22788(.A(new_n25224_), .Y(new_n25225_));
  AOI21X1  g22789(.A0(new_n25199_), .A1(new_n25196_), .B0(new_n22660_), .Y(new_n25226_));
  NAND2X1  g22790(.A(new_n25226_), .B(new_n25225_), .Y(new_n25227_));
  NOR2X1   g22791(.A(new_n9445_), .B(new_n12487_), .Y(new_n25228_));
  NOR3X1   g22792(.A(new_n25228_), .B(new_n25208_), .C(new_n25206_), .Y(new_n25229_));
  OAI21X1  g22793(.A0(new_n25229_), .A1(pi0207), .B0(new_n25227_), .Y(new_n25230_));
  MX2X1    g22794(.A(new_n25230_), .B(new_n25223_), .S0(new_n22959_), .Y(new_n25231_));
  AND2X1   g22795(.A(new_n25231_), .B(new_n23173_), .Y(new_n25232_));
  AND3X1   g22796(.A(pi1153), .B(pi0299), .C(new_n22660_), .Y(new_n25233_));
  OAI22X1  g22797(.A0(new_n24916_), .A1(pi1153), .B0(new_n24903_), .B1(pi0299), .Y(new_n25234_));
  NOR2X1   g22798(.A(new_n24916_), .B(pi1153), .Y(new_n25235_));
  OAI21X1  g22799(.A0(pi0299), .A1(new_n7871_), .B0(pi1154), .Y(new_n25236_));
  OR2X1    g22800(.A(new_n25236_), .B(new_n25235_), .Y(new_n25237_));
  AND2X1   g22801(.A(new_n25237_), .B(new_n25234_), .Y(new_n25238_));
  INVX1    g22802(.A(new_n25238_), .Y(new_n25239_));
  AOI21X1  g22803(.A0(new_n25239_), .A1(pi0207), .B0(new_n25233_), .Y(new_n25240_));
  NOR2X1   g22804(.A(new_n9445_), .B(pi1153), .Y(new_n25241_));
  INVX1    g22805(.A(new_n25241_), .Y(new_n25242_));
  AOI21X1  g22806(.A0(new_n25130_), .A1(new_n2933_), .B0(new_n22660_), .Y(new_n25243_));
  AOI22X1  g22807(.A0(new_n25243_), .A1(new_n25242_), .B0(new_n25239_), .B1(new_n22660_), .Y(new_n25244_));
  MX2X1    g22808(.A(new_n25244_), .B(new_n25240_), .S0(new_n22959_), .Y(new_n25245_));
  NOR2X1   g22809(.A(new_n25245_), .B(new_n23173_), .Y(new_n25246_));
  NOR2X1   g22810(.A(new_n25246_), .B(new_n25232_), .Y(new_n25247_));
  NOR2X1   g22811(.A(new_n25245_), .B(pi0211), .Y(new_n25248_));
  OAI21X1  g22812(.A0(new_n25202_), .A1(new_n23173_), .B0(pi0214), .Y(new_n25249_));
  OAI21X1  g22813(.A0(new_n25249_), .A1(new_n25248_), .B0(pi0212), .Y(new_n25250_));
  AOI21X1  g22814(.A0(new_n25247_), .A1(new_n24849_), .B0(new_n25250_), .Y(new_n25251_));
  AOI21X1  g22815(.A0(new_n25216_), .A1(new_n24849_), .B0(pi0212), .Y(new_n25252_));
  INVX1    g22816(.A(new_n25252_), .Y(new_n25253_));
  AOI21X1  g22817(.A0(new_n25247_), .A1(pi0214), .B0(new_n25253_), .Y(new_n25254_));
  OR3X1    g22818(.A(new_n25254_), .B(new_n25251_), .C(pi0219), .Y(new_n25255_));
  NAND2X1  g22819(.A(new_n25255_), .B(new_n25221_), .Y(new_n25256_));
  OR2X1    g22820(.A(pi1154), .B(new_n12364_), .Y(new_n25257_));
  OAI22X1  g22821(.A0(new_n25257_), .A1(new_n24998_), .B0(new_n25236_), .B1(new_n25235_), .Y(new_n25258_));
  AOI21X1  g22822(.A0(new_n25258_), .A1(pi0207), .B0(new_n25233_), .Y(new_n25259_));
  NOR2X1   g22823(.A(new_n9445_), .B(new_n22660_), .Y(new_n25260_));
  AOI22X1  g22824(.A0(new_n25260_), .A1(pi1153), .B0(new_n25258_), .B1(new_n22660_), .Y(new_n25261_));
  MX2X1    g22825(.A(new_n25261_), .B(new_n25259_), .S0(new_n22959_), .Y(new_n25262_));
  INVX1    g22826(.A(new_n25189_), .Y(new_n25263_));
  AOI21X1  g22827(.A0(new_n2933_), .A1(pi0199), .B0(new_n12364_), .Y(new_n25264_));
  OAI21X1  g22828(.A0(new_n25264_), .A1(new_n25241_), .B0(pi1154), .Y(new_n25265_));
  AOI21X1  g22829(.A0(new_n25265_), .A1(new_n25263_), .B0(new_n22660_), .Y(new_n25266_));
  OR2X1    g22830(.A(new_n25266_), .B(new_n25126_), .Y(new_n25267_));
  NAND3X1  g22831(.A(new_n25265_), .B(new_n25263_), .C(new_n22660_), .Y(new_n25268_));
  OAI21X1  g22832(.A0(new_n8058_), .A1(new_n12364_), .B0(new_n2933_), .Y(new_n25269_));
  AOI21X1  g22833(.A0(new_n25269_), .A1(new_n25225_), .B0(new_n22660_), .Y(new_n25270_));
  NOR2X1   g22834(.A(new_n25270_), .B(new_n22959_), .Y(new_n25271_));
  AOI22X1  g22835(.A0(new_n25271_), .A1(new_n25268_), .B0(new_n25267_), .B1(new_n22959_), .Y(new_n25272_));
  MX2X1    g22836(.A(new_n25272_), .B(new_n25262_), .S0(pi0211), .Y(new_n25273_));
  AOI22X1  g22837(.A0(new_n25273_), .A1(new_n25085_), .B0(new_n25262_), .B1(new_n25044_), .Y(new_n25274_));
  INVX1    g22838(.A(new_n8423_), .Y(new_n25275_));
  AOI21X1  g22839(.A0(new_n12364_), .A1(pi0200), .B0(new_n25275_), .Y(new_n25276_));
  MX2X1    g22840(.A(new_n25276_), .B(new_n25189_), .S0(new_n12487_), .Y(new_n25277_));
  AND3X1   g22841(.A(new_n2933_), .B(pi0208), .C(pi0207), .Y(new_n25278_));
  NOR2X1   g22842(.A(new_n9445_), .B(new_n12364_), .Y(new_n25279_));
  AOI22X1  g22843(.A0(new_n25279_), .A1(new_n25278_), .B0(new_n25277_), .B1(new_n25115_), .Y(new_n25280_));
  INVX1    g22844(.A(new_n25280_), .Y(new_n25281_));
  OAI21X1  g22845(.A0(new_n25281_), .A1(new_n8422_), .B0(new_n6489_), .Y(new_n25282_));
  AOI21X1  g22846(.A0(pi0214), .A1(new_n23173_), .B0(new_n25085_), .Y(new_n25283_));
  AOI21X1  g22847(.A0(new_n25283_), .A1(new_n25280_), .B0(new_n25282_), .Y(new_n25284_));
  OAI21X1  g22848(.A0(new_n25274_), .A1(pi0219), .B0(new_n25284_), .Y(new_n25285_));
  AOI22X1  g22849(.A0(new_n25285_), .A1(new_n25114_), .B0(new_n25256_), .B1(new_n25159_), .Y(new_n25286_));
  AND3X1   g22850(.A(new_n5102_), .B(new_n25153_), .C(new_n2436_), .Y(new_n25287_));
  AND2X1   g22851(.A(new_n12463_), .B(pi0299), .Y(new_n25288_));
  AND3X1   g22852(.A(pi1153), .B(pi0200), .C(new_n7871_), .Y(new_n25289_));
  OAI21X1  g22853(.A0(new_n25289_), .A1(pi0299), .B0(new_n12487_), .Y(new_n25290_));
  OR2X1    g22854(.A(new_n25290_), .B(new_n25288_), .Y(new_n25291_));
  OR2X1    g22855(.A(new_n25265_), .B(new_n24971_), .Y(new_n25292_));
  AND3X1   g22856(.A(new_n25292_), .B(new_n25291_), .C(pi0207), .Y(new_n25293_));
  NOR2X1   g22857(.A(new_n25293_), .B(new_n24968_), .Y(new_n25294_));
  AND3X1   g22858(.A(new_n25292_), .B(new_n25291_), .C(new_n22660_), .Y(new_n25295_));
  INVX1    g22859(.A(new_n25288_), .Y(new_n25296_));
  AOI21X1  g22860(.A0(new_n25269_), .A1(new_n25296_), .B0(new_n22660_), .Y(new_n25297_));
  NOR3X1   g22861(.A(new_n25297_), .B(new_n25295_), .C(new_n22959_), .Y(new_n25298_));
  OR3X1    g22862(.A(new_n25298_), .B(new_n25294_), .C(pi0211), .Y(new_n25299_));
  AOI21X1  g22863(.A0(new_n25272_), .A1(pi0211), .B0(new_n24877_), .Y(new_n25300_));
  OR3X1    g22864(.A(new_n25298_), .B(new_n25294_), .C(new_n23173_), .Y(new_n25301_));
  AOI21X1  g22865(.A0(pi1156), .A1(pi0299), .B0(pi0211), .Y(new_n25302_));
  AOI21X1  g22866(.A0(new_n25302_), .A1(new_n25280_), .B0(new_n24824_), .Y(new_n25303_));
  AOI22X1  g22867(.A0(new_n25303_), .A1(new_n25301_), .B0(new_n25300_), .B1(new_n25299_), .Y(new_n25304_));
  NAND2X1  g22868(.A(new_n25272_), .B(new_n23173_), .Y(new_n25305_));
  OAI21X1  g22869(.A0(pi0214), .A1(pi0212), .B0(pi0219), .Y(new_n25306_));
  AOI21X1  g22870(.A0(new_n25280_), .A1(pi0211), .B0(new_n25306_), .Y(new_n25307_));
  AOI22X1  g22871(.A0(new_n25307_), .A1(new_n25305_), .B0(new_n25281_), .B1(new_n24816_), .Y(new_n25308_));
  OAI21X1  g22872(.A0(new_n25304_), .A1(pi0219), .B0(new_n25308_), .Y(new_n25309_));
  AOI22X1  g22873(.A0(new_n25232_), .A1(new_n25188_), .B0(new_n25217_), .B1(new_n25162_), .Y(new_n25310_));
  AND2X1   g22874(.A(new_n25231_), .B(pi0211), .Y(new_n25311_));
  AOI22X1  g22875(.A0(new_n25201_), .A1(new_n25194_), .B0(new_n25193_), .B1(new_n24965_), .Y(new_n25312_));
  NOR2X1   g22876(.A(pi1154), .B(pi0199), .Y(new_n25313_));
  AND3X1   g22877(.A(new_n25313_), .B(new_n24984_), .C(new_n7937_), .Y(new_n25314_));
  NOR4X1   g22878(.A(new_n25314_), .B(new_n25312_), .C(new_n25288_), .D(pi0211), .Y(new_n25315_));
  OR2X1    g22879(.A(new_n25315_), .B(new_n24877_), .Y(new_n25316_));
  OR4X1    g22880(.A(new_n25314_), .B(new_n25312_), .C(new_n25288_), .D(new_n23173_), .Y(new_n25317_));
  OAI21X1  g22881(.A0(new_n25210_), .A1(new_n25022_), .B0(new_n22660_), .Y(new_n25318_));
  OAI21X1  g22882(.A0(pi1156), .A1(new_n2933_), .B0(new_n25226_), .Y(new_n25319_));
  NAND3X1  g22883(.A(new_n25319_), .B(new_n25318_), .C(pi0208), .Y(new_n25320_));
  AOI21X1  g22884(.A0(pi1156), .A1(pi0299), .B0(pi0208), .Y(new_n25321_));
  AOI21X1  g22885(.A0(new_n25321_), .A1(new_n25222_), .B0(pi0211), .Y(new_n25322_));
  AOI21X1  g22886(.A0(new_n25322_), .A1(new_n25320_), .B0(new_n24824_), .Y(new_n25323_));
  AND3X1   g22887(.A(new_n25216_), .B(new_n24849_), .C(new_n24823_), .Y(new_n25324_));
  OR2X1    g22888(.A(new_n25324_), .B(pi0219), .Y(new_n25325_));
  AOI21X1  g22889(.A0(new_n25323_), .A1(new_n25317_), .B0(new_n25325_), .Y(new_n25326_));
  OAI21X1  g22890(.A0(new_n25316_), .A1(new_n25311_), .B0(new_n25326_), .Y(new_n25327_));
  OAI21X1  g22891(.A0(new_n25310_), .A1(new_n8422_), .B0(new_n25327_), .Y(new_n25328_));
  AND3X1   g22892(.A(new_n5102_), .B(pi1152), .C(new_n2436_), .Y(new_n25329_));
  AOI22X1  g22893(.A0(new_n25329_), .A1(new_n25328_), .B0(new_n25309_), .B1(new_n25287_), .Y(new_n25330_));
  OAI21X1  g22894(.A0(new_n25330_), .A1(new_n24815_), .B0(new_n24866_), .Y(new_n25331_));
  AOI21X1  g22895(.A0(new_n25286_), .A1(new_n24815_), .B0(new_n25331_), .Y(new_n25332_));
  NOR2X1   g22896(.A(new_n24871_), .B(new_n24823_), .Y(new_n25333_));
  NOR3X1   g22897(.A(new_n24869_), .B(new_n24849_), .C(pi0212), .Y(new_n25334_));
  OR2X1    g22898(.A(new_n25334_), .B(pi0219), .Y(new_n25335_));
  NOR2X1   g22899(.A(new_n25335_), .B(new_n25333_), .Y(new_n25336_));
  AOI21X1  g22900(.A0(pi1154), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n25337_));
  OR4X1    g22901(.A(new_n25337_), .B(new_n24818_), .C(new_n6489_), .D(new_n24815_), .Y(new_n25338_));
  OAI22X1  g22902(.A0(new_n25338_), .A1(new_n25336_), .B0(new_n25332_), .B1(new_n25187_), .Y(new_n25339_));
  MX2X1    g22903(.A(new_n25339_), .B(pi0234), .S0(new_n24814_), .Y(po0391));
  NOR2X1   g22904(.A(new_n24998_), .B(new_n12463_), .Y(new_n25341_));
  OAI21X1  g22905(.A0(new_n25341_), .A1(new_n24928_), .B0(pi0207), .Y(new_n25342_));
  NOR4X1   g22906(.A(new_n24971_), .B(new_n24970_), .C(new_n24969_), .D(pi0207), .Y(new_n25343_));
  INVX1    g22907(.A(new_n25343_), .Y(new_n25344_));
  AOI21X1  g22908(.A0(new_n25344_), .A1(new_n25342_), .B0(new_n22959_), .Y(new_n25345_));
  OAI21X1  g22909(.A0(new_n25345_), .A1(new_n24972_), .B0(new_n12578_), .Y(new_n25346_));
  AND2X1   g22910(.A(pi1157), .B(pi0208), .Y(new_n25347_));
  OAI21X1  g22911(.A0(new_n24964_), .A1(pi0207), .B0(new_n25342_), .Y(new_n25348_));
  AOI21X1  g22912(.A0(new_n25348_), .A1(new_n25347_), .B0(new_n24967_), .Y(new_n25349_));
  AOI21X1  g22913(.A0(new_n25349_), .A1(new_n25346_), .B0(new_n23173_), .Y(new_n25350_));
  AND2X1   g22914(.A(new_n25005_), .B(new_n24901_), .Y(new_n25351_));
  MX2X1    g22915(.A(new_n24996_), .B(new_n25096_), .S0(new_n12555_), .Y(new_n25352_));
  NOR2X1   g22916(.A(new_n25352_), .B(new_n22660_), .Y(new_n25353_));
  AOI21X1  g22917(.A0(new_n25351_), .A1(new_n22660_), .B0(new_n25353_), .Y(new_n25354_));
  OAI22X1  g22918(.A0(new_n25354_), .A1(new_n22959_), .B0(new_n25007_), .B1(new_n24900_), .Y(new_n25355_));
  NOR2X1   g22919(.A(new_n24982_), .B(new_n12555_), .Y(new_n25356_));
  OAI21X1  g22920(.A0(new_n25356_), .A1(new_n24936_), .B0(new_n22660_), .Y(new_n25357_));
  OAI21X1  g22921(.A0(new_n25352_), .A1(new_n22660_), .B0(new_n25357_), .Y(new_n25358_));
  NAND2X1  g22922(.A(new_n25358_), .B(new_n25347_), .Y(new_n25359_));
  NAND2X1  g22923(.A(new_n25359_), .B(new_n25027_), .Y(new_n25360_));
  AOI21X1  g22924(.A0(new_n25355_), .A1(new_n12578_), .B0(new_n25360_), .Y(new_n25361_));
  OAI21X1  g22925(.A0(new_n25361_), .A1(pi0211), .B0(new_n7996_), .Y(new_n25362_));
  NOR2X1   g22926(.A(new_n25362_), .B(new_n25350_), .Y(new_n25363_));
  AND2X1   g22927(.A(new_n24922_), .B(new_n12555_), .Y(new_n25364_));
  NOR3X1   g22928(.A(new_n25364_), .B(new_n24928_), .C(new_n7827_), .Y(new_n25365_));
  AND3X1   g22929(.A(new_n24903_), .B(new_n24902_), .C(new_n2933_), .Y(new_n25366_));
  AOI21X1  g22930(.A0(new_n25366_), .A1(new_n24901_), .B0(pi0207), .Y(new_n25367_));
  NOR3X1   g22931(.A(new_n25367_), .B(new_n25365_), .C(new_n24906_), .Y(new_n25368_));
  NOR3X1   g22932(.A(new_n24936_), .B(new_n24935_), .C(pi0207), .Y(new_n25369_));
  NOR3X1   g22933(.A(new_n25369_), .B(new_n25365_), .C(new_n24939_), .Y(new_n25370_));
  MX2X1    g22934(.A(new_n25370_), .B(new_n25368_), .S0(new_n12578_), .Y(new_n25371_));
  AOI21X1  g22935(.A0(new_n24983_), .A1(new_n22660_), .B0(new_n22959_), .Y(new_n25372_));
  NAND3X1  g22936(.A(new_n24999_), .B(new_n24997_), .C(pi0207), .Y(new_n25373_));
  AOI21X1  g22937(.A0(new_n25373_), .A1(new_n25372_), .B0(new_n24987_), .Y(new_n25374_));
  NAND2X1  g22938(.A(new_n25374_), .B(pi1157), .Y(new_n25375_));
  NOR2X1   g22939(.A(new_n25368_), .B(pi1157), .Y(new_n25376_));
  NOR2X1   g22940(.A(new_n25376_), .B(pi0211), .Y(new_n25377_));
  AOI21X1  g22941(.A0(new_n25377_), .A1(new_n25375_), .B0(new_n25086_), .Y(new_n25378_));
  OAI21X1  g22942(.A0(new_n25361_), .A1(new_n23173_), .B0(new_n25378_), .Y(new_n25379_));
  OAI21X1  g22943(.A0(new_n25371_), .A1(new_n25188_), .B0(new_n25379_), .Y(new_n25380_));
  OAI21X1  g22944(.A0(new_n25380_), .A1(new_n25363_), .B0(new_n8422_), .Y(new_n25381_));
  AND3X1   g22945(.A(new_n25349_), .B(new_n25346_), .C(new_n23173_), .Y(new_n25382_));
  INVX1    g22946(.A(new_n24824_), .Y(new_n25383_));
  OAI21X1  g22947(.A0(new_n25371_), .A1(new_n23173_), .B0(new_n25383_), .Y(new_n25384_));
  AOI21X1  g22948(.A0(new_n25371_), .A1(new_n24824_), .B0(new_n8422_), .Y(new_n25385_));
  OAI21X1  g22949(.A0(new_n25384_), .A1(new_n25382_), .B0(new_n25385_), .Y(new_n25386_));
  AND3X1   g22950(.A(new_n25386_), .B(new_n25381_), .C(pi0209), .Y(new_n25387_));
  AOI21X1  g22951(.A0(new_n24993_), .A1(new_n24839_), .B0(new_n24986_), .Y(new_n25388_));
  AND3X1   g22952(.A(new_n25290_), .B(new_n25265_), .C(pi0207), .Y(new_n25389_));
  OR2X1    g22953(.A(new_n25389_), .B(new_n22959_), .Y(new_n25390_));
  AOI21X1  g22954(.A0(new_n24993_), .A1(new_n24984_), .B0(new_n25390_), .Y(new_n25391_));
  OAI21X1  g22955(.A0(new_n25391_), .A1(new_n25388_), .B0(pi1157), .Y(new_n25392_));
  OAI21X1  g22956(.A0(new_n25211_), .A1(new_n24921_), .B0(new_n7827_), .Y(new_n25393_));
  OAI21X1  g22957(.A0(new_n25277_), .A1(new_n7827_), .B0(new_n25393_), .Y(new_n25394_));
  INVX1    g22958(.A(new_n25394_), .Y(new_n25395_));
  AOI21X1  g22959(.A0(new_n25395_), .A1(new_n12578_), .B0(pi0211), .Y(new_n25396_));
  AND3X1   g22960(.A(new_n25394_), .B(new_n25023_), .C(pi0211), .Y(new_n25397_));
  AOI21X1  g22961(.A0(new_n25396_), .A1(new_n25392_), .B0(new_n25397_), .Y(new_n25398_));
  AND2X1   g22962(.A(new_n24954_), .B(new_n22660_), .Y(new_n25399_));
  OR2X1    g22963(.A(new_n25293_), .B(new_n22959_), .Y(new_n25400_));
  OAI22X1  g22964(.A0(new_n25400_), .A1(new_n25399_), .B0(new_n24968_), .B1(new_n24954_), .Y(new_n25401_));
  NAND2X1  g22965(.A(new_n25401_), .B(pi0211), .Y(new_n25402_));
  AOI21X1  g22966(.A0(new_n25394_), .A1(new_n25023_), .B0(pi0211), .Y(new_n25403_));
  NOR2X1   g22967(.A(new_n25403_), .B(new_n24877_), .Y(new_n25404_));
  AOI22X1  g22968(.A0(new_n25404_), .A1(new_n25402_), .B0(new_n25394_), .B1(new_n24816_), .Y(new_n25405_));
  OAI21X1  g22969(.A0(new_n25398_), .A1(new_n25086_), .B0(new_n25405_), .Y(new_n25406_));
  AOI21X1  g22970(.A0(new_n25394_), .A1(pi0211), .B0(new_n24824_), .Y(new_n25407_));
  OAI21X1  g22971(.A0(new_n25401_), .A1(pi0211), .B0(new_n25407_), .Y(new_n25408_));
  AOI21X1  g22972(.A0(new_n25395_), .A1(new_n24824_), .B0(new_n8422_), .Y(new_n25409_));
  AND2X1   g22973(.A(new_n25409_), .B(new_n25408_), .Y(new_n25410_));
  OR2X1    g22974(.A(new_n25410_), .B(pi0209), .Y(new_n25411_));
  AOI21X1  g22975(.A0(new_n25406_), .A1(new_n8422_), .B0(new_n25411_), .Y(new_n25412_));
  OAI21X1  g22976(.A0(new_n25412_), .A1(new_n25387_), .B0(new_n6489_), .Y(new_n25413_));
  NAND3X1  g22977(.A(new_n24867_), .B(pi0214), .C(new_n24823_), .Y(new_n25414_));
  NAND2X1  g22978(.A(new_n24867_), .B(new_n24849_), .Y(new_n25415_));
  OAI21X1  g22979(.A0(new_n24869_), .A1(new_n24849_), .B0(new_n25415_), .Y(new_n25416_));
  AOI21X1  g22980(.A0(new_n25416_), .A1(pi0212), .B0(pi0219), .Y(new_n25417_));
  NAND2X1  g22981(.A(new_n25417_), .B(new_n25414_), .Y(new_n25418_));
  AOI21X1  g22982(.A0(pi1155), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n25419_));
  NOR2X1   g22983(.A(new_n25085_), .B(new_n8422_), .Y(new_n25420_));
  NOR3X1   g22984(.A(new_n25420_), .B(new_n25419_), .C(new_n6489_), .Y(new_n25421_));
  AOI21X1  g22985(.A0(new_n25421_), .A1(new_n25418_), .B0(new_n24815_), .Y(new_n25422_));
  INVX1    g22986(.A(new_n25384_), .Y(new_n25423_));
  NOR2X1   g22987(.A(new_n25374_), .B(new_n12578_), .Y(new_n25424_));
  INVX1    g22988(.A(new_n25424_), .Y(new_n25425_));
  OAI21X1  g22989(.A0(new_n25355_), .A1(pi0299), .B0(new_n12578_), .Y(new_n25426_));
  AOI21X1  g22990(.A0(new_n25426_), .A1(new_n25425_), .B0(new_n25001_), .Y(new_n25427_));
  OAI21X1  g22991(.A0(new_n25427_), .A1(pi0211), .B0(new_n25423_), .Y(new_n25428_));
  AND2X1   g22992(.A(new_n25428_), .B(new_n25385_), .Y(new_n25429_));
  NAND2X1  g22993(.A(new_n25427_), .B(pi0211), .Y(new_n25430_));
  INVX1    g22994(.A(new_n24988_), .Y(new_n25431_));
  NOR2X1   g22995(.A(new_n24999_), .B(new_n24923_), .Y(new_n25432_));
  OAI21X1  g22996(.A0(new_n25432_), .A1(new_n24928_), .B0(pi0207), .Y(new_n25433_));
  AOI21X1  g22997(.A0(new_n25005_), .A1(pi1154), .B0(new_n25366_), .Y(new_n25434_));
  OR3X1    g22998(.A(new_n25434_), .B(new_n24969_), .C(pi0207), .Y(new_n25435_));
  AOI21X1  g22999(.A0(new_n25435_), .A1(new_n25433_), .B0(new_n22959_), .Y(new_n25436_));
  OAI21X1  g23000(.A0(new_n25436_), .A1(new_n24989_), .B0(new_n12578_), .Y(new_n25437_));
  OAI21X1  g23001(.A0(new_n25374_), .A1(new_n25431_), .B0(new_n25437_), .Y(new_n25438_));
  AOI21X1  g23002(.A0(new_n25438_), .A1(new_n23173_), .B0(new_n24877_), .Y(new_n25439_));
  NAND2X1  g23003(.A(new_n25439_), .B(new_n25430_), .Y(new_n25440_));
  NOR2X1   g23004(.A(new_n25371_), .B(new_n25188_), .Y(new_n25441_));
  NOR2X1   g23005(.A(new_n25438_), .B(new_n23173_), .Y(new_n25442_));
  OR2X1    g23006(.A(new_n25442_), .B(new_n25382_), .Y(new_n25443_));
  AOI21X1  g23007(.A0(new_n25443_), .A1(new_n25085_), .B0(new_n25441_), .Y(new_n25444_));
  AOI21X1  g23008(.A0(new_n25444_), .A1(new_n25440_), .B0(pi0219), .Y(new_n25445_));
  OAI21X1  g23009(.A0(new_n25445_), .A1(new_n25429_), .B0(pi0209), .Y(new_n25446_));
  INVX1    g23010(.A(new_n25407_), .Y(new_n25447_));
  OAI21X1  g23011(.A0(new_n25233_), .A1(new_n24994_), .B0(new_n22959_), .Y(new_n25448_));
  NAND2X1  g23012(.A(new_n25258_), .B(pi0207), .Y(new_n25449_));
  OAI21X1  g23013(.A0(new_n24993_), .A1(pi0207), .B0(new_n25449_), .Y(new_n25450_));
  NAND2X1  g23014(.A(new_n25450_), .B(pi0208), .Y(new_n25451_));
  AND3X1   g23015(.A(new_n25451_), .B(new_n25448_), .C(new_n23173_), .Y(new_n25452_));
  OAI21X1  g23016(.A0(new_n25452_), .A1(new_n25447_), .B0(new_n25409_), .Y(new_n25453_));
  AOI21X1  g23017(.A0(new_n24978_), .A1(pi0207), .B0(new_n25126_), .Y(new_n25454_));
  OR2X1    g23018(.A(new_n25454_), .B(pi0208), .Y(new_n25455_));
  AOI21X1  g23019(.A0(new_n24978_), .A1(new_n22660_), .B0(new_n25266_), .Y(new_n25456_));
  OR2X1    g23020(.A(new_n25456_), .B(new_n22959_), .Y(new_n25457_));
  NAND3X1  g23021(.A(new_n25457_), .B(new_n25455_), .C(pi0211), .Y(new_n25458_));
  OAI21X1  g23022(.A0(new_n25401_), .A1(pi0211), .B0(new_n25458_), .Y(new_n25459_));
  AOI21X1  g23023(.A0(new_n25457_), .A1(new_n25455_), .B0(pi0211), .Y(new_n25460_));
  AOI21X1  g23024(.A0(new_n25451_), .A1(new_n25448_), .B0(new_n23173_), .Y(new_n25461_));
  OR3X1    g23025(.A(new_n25461_), .B(new_n25460_), .C(new_n24877_), .Y(new_n25462_));
  OAI21X1  g23026(.A0(new_n25395_), .A1(new_n25188_), .B0(new_n25462_), .Y(new_n25463_));
  AOI21X1  g23027(.A0(new_n25459_), .A1(new_n25383_), .B0(new_n25463_), .Y(new_n25464_));
  OAI21X1  g23028(.A0(new_n25464_), .A1(pi0219), .B0(new_n25453_), .Y(new_n25465_));
  AOI21X1  g23029(.A0(new_n25465_), .A1(new_n24866_), .B0(po1038), .Y(new_n25466_));
  AOI21X1  g23030(.A0(pi1153), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n25467_));
  OR2X1    g23031(.A(new_n25467_), .B(new_n6489_), .Y(new_n25468_));
  AOI21X1  g23032(.A0(new_n25156_), .A1(new_n7996_), .B0(pi0219), .Y(new_n25469_));
  OAI21X1  g23033(.A0(new_n25086_), .A1(new_n24870_), .B0(new_n25469_), .Y(new_n25470_));
  OAI21X1  g23034(.A0(new_n25085_), .A1(new_n8422_), .B0(new_n25470_), .Y(new_n25471_));
  OAI21X1  g23035(.A0(new_n25471_), .A1(new_n25468_), .B0(new_n24815_), .Y(new_n25472_));
  AOI21X1  g23036(.A0(new_n25466_), .A1(new_n25446_), .B0(new_n25472_), .Y(new_n25473_));
  AOI21X1  g23037(.A0(new_n25422_), .A1(new_n25413_), .B0(new_n25473_), .Y(new_n25474_));
  MX2X1    g23038(.A(new_n25474_), .B(pi0235), .S0(new_n24814_), .Y(po0392));
  OAI21X1  g23039(.A0(new_n24671_), .A1(pi0100), .B0(new_n24805_), .Y(new_n25476_));
  AOI21X1  g23040(.A0(new_n25476_), .A1(new_n5090_), .B0(pi0075), .Y(new_n25477_));
  OAI21X1  g23041(.A0(new_n25477_), .A1(new_n5780_), .B0(new_n3079_), .Y(new_n25478_));
  AOI21X1  g23042(.A0(new_n25478_), .A1(new_n11150_), .B0(pi0074), .Y(new_n25479_));
  OAI21X1  g23043(.A0(new_n25479_), .A1(new_n4985_), .B0(new_n3118_), .Y(new_n25480_));
  AOI21X1  g23044(.A0(new_n25480_), .A1(new_n4981_), .B0(pi0062), .Y(new_n25481_));
  NOR2X1   g23045(.A(new_n25481_), .B(new_n9834_), .Y(po0393));
  MX2X1    g23046(.A(pi1158), .B(pi1157), .S0(pi0211), .Y(new_n25483_));
  NAND3X1  g23047(.A(new_n25483_), .B(pi0214), .C(new_n24823_), .Y(new_n25484_));
  AND2X1   g23048(.A(new_n25484_), .B(new_n25417_), .Y(new_n25485_));
  OR4X1    g23049(.A(new_n12555_), .B(new_n24849_), .C(pi0212), .D(pi0211), .Y(new_n25486_));
  AOI21X1  g23050(.A0(new_n25486_), .A1(pi0219), .B0(new_n6489_), .Y(new_n25487_));
  AND2X1   g23051(.A(pi1154), .B(new_n23173_), .Y(new_n25488_));
  AOI22X1  g23052(.A0(new_n24974_), .A1(pi1155), .B0(new_n25488_), .B1(pi0214), .Y(new_n25489_));
  NOR3X1   g23053(.A(new_n25489_), .B(new_n6489_), .C(new_n24823_), .Y(new_n25490_));
  NOR2X1   g23054(.A(new_n25490_), .B(new_n25487_), .Y(new_n25491_));
  OAI21X1  g23055(.A0(new_n25491_), .A1(new_n25485_), .B0(new_n24815_), .Y(new_n25492_));
  NOR3X1   g23056(.A(new_n25485_), .B(new_n2933_), .C(pi0219), .Y(new_n25493_));
  AOI21X1  g23057(.A0(pi1143), .A1(pi0199), .B0(pi0200), .Y(new_n25494_));
  OAI21X1  g23058(.A0(new_n2439_), .A1(pi0199), .B0(new_n25494_), .Y(new_n25495_));
  AND3X1   g23059(.A(new_n25495_), .B(new_n25278_), .C(new_n24835_), .Y(new_n25496_));
  OAI21X1  g23060(.A0(new_n3309_), .A1(pi0199), .B0(new_n25494_), .Y(new_n25497_));
  OAI21X1  g23061(.A0(new_n2439_), .A1(pi0199), .B0(pi0200), .Y(new_n25498_));
  AND3X1   g23062(.A(new_n25498_), .B(new_n25497_), .C(new_n25115_), .Y(new_n25499_));
  OAI21X1  g23063(.A0(new_n25499_), .A1(new_n25496_), .B0(new_n2933_), .Y(new_n25500_));
  INVX1    g23064(.A(new_n25500_), .Y(new_n25501_));
  NAND3X1  g23065(.A(new_n25022_), .B(pi0214), .C(new_n24823_), .Y(new_n25502_));
  AOI21X1  g23066(.A0(new_n24955_), .A1(new_n24849_), .B0(new_n24823_), .Y(new_n25503_));
  OAI21X1  g23067(.A0(new_n24889_), .A1(new_n24849_), .B0(new_n25503_), .Y(new_n25504_));
  AOI21X1  g23068(.A0(new_n25504_), .A1(new_n25502_), .B0(new_n24894_), .Y(new_n25505_));
  OR3X1    g23069(.A(new_n25505_), .B(new_n25501_), .C(new_n25493_), .Y(new_n25506_));
  AOI21X1  g23070(.A0(new_n25506_), .A1(new_n6489_), .B0(new_n25492_), .Y(new_n25507_));
  MX2X1    g23071(.A(pi1145), .B(pi1144), .S0(pi0211), .Y(new_n25508_));
  OAI21X1  g23072(.A0(new_n25508_), .A1(new_n7996_), .B0(new_n25188_), .Y(new_n25509_));
  AOI21X1  g23073(.A0(new_n24822_), .A1(new_n7996_), .B0(new_n25509_), .Y(new_n25510_));
  OAI21X1  g23074(.A0(new_n24821_), .A1(pi0211), .B0(pi0219), .Y(new_n25511_));
  AND2X1   g23075(.A(new_n25511_), .B(new_n24819_), .Y(new_n25512_));
  OAI21X1  g23076(.A0(new_n25510_), .A1(pi0219), .B0(new_n25512_), .Y(new_n25513_));
  NOR4X1   g23077(.A(new_n25306_), .B(new_n24821_), .C(new_n2933_), .D(pi0211), .Y(new_n25514_));
  AOI21X1  g23078(.A0(new_n25510_), .A1(new_n24884_), .B0(new_n25514_), .Y(new_n25515_));
  AND2X1   g23079(.A(new_n25515_), .B(new_n25500_), .Y(new_n25516_));
  OAI21X1  g23080(.A0(new_n25516_), .A1(po1038), .B0(new_n25513_), .Y(new_n25517_));
  OAI21X1  g23081(.A0(new_n25517_), .A1(new_n24815_), .B0(pi0209), .Y(new_n25518_));
  OR2X1    g23082(.A(pi1158), .B(pi0199), .Y(new_n25519_));
  AOI22X1  g23083(.A0(new_n25519_), .A1(pi1156), .B0(new_n25204_), .B1(pi1158), .Y(new_n25520_));
  NOR4X1   g23084(.A(new_n25520_), .B(new_n24917_), .C(pi0208), .D(new_n22660_), .Y(new_n25521_));
  AND2X1   g23085(.A(new_n24929_), .B(pi0207), .Y(new_n25522_));
  NOR3X1   g23086(.A(new_n25522_), .B(new_n25367_), .C(new_n22959_), .Y(new_n25523_));
  OAI21X1  g23087(.A0(new_n25523_), .A1(new_n25521_), .B0(new_n12578_), .Y(new_n25524_));
  AOI21X1  g23088(.A0(new_n12548_), .A1(new_n7937_), .B0(pi0199), .Y(new_n25525_));
  AOI21X1  g23089(.A0(new_n25195_), .A1(pi1156), .B0(new_n25525_), .Y(new_n25526_));
  OR2X1    g23090(.A(new_n25526_), .B(new_n24840_), .Y(new_n25527_));
  NOR2X1   g23091(.A(new_n25369_), .B(new_n22959_), .Y(new_n25528_));
  INVX1    g23092(.A(new_n25528_), .Y(new_n25529_));
  OAI22X1  g23093(.A0(new_n25529_), .A1(new_n25522_), .B0(new_n25527_), .B1(pi0208), .Y(new_n25530_));
  NAND2X1  g23094(.A(new_n25530_), .B(pi1157), .Y(new_n25531_));
  AND3X1   g23095(.A(new_n25531_), .B(new_n25524_), .C(new_n25162_), .Y(new_n25532_));
  INVX1    g23096(.A(new_n24886_), .Y(new_n25533_));
  INVX1    g23097(.A(new_n25347_), .Y(new_n25534_));
  AOI21X1  g23098(.A0(new_n25357_), .A1(new_n25168_), .B0(new_n25534_), .Y(new_n25535_));
  AOI21X1  g23099(.A0(new_n25351_), .A1(new_n22660_), .B0(new_n22959_), .Y(new_n25536_));
  INVX1    g23100(.A(new_n25321_), .Y(new_n25537_));
  NOR3X1   g23101(.A(new_n25520_), .B(new_n22660_), .C(pi0200), .Y(new_n25538_));
  OAI21X1  g23102(.A0(new_n25538_), .A1(new_n25537_), .B0(new_n12578_), .Y(new_n25539_));
  AOI21X1  g23103(.A0(new_n25536_), .A1(new_n25168_), .B0(new_n25539_), .Y(new_n25540_));
  INVX1    g23104(.A(new_n25026_), .Y(new_n25541_));
  AOI21X1  g23105(.A0(new_n25527_), .A1(new_n25023_), .B0(new_n25541_), .Y(new_n25542_));
  OR4X1    g23106(.A(new_n25542_), .B(new_n25540_), .C(new_n25535_), .D(new_n25533_), .Y(new_n25543_));
  OAI21X1  g23107(.A0(new_n25172_), .A1(new_n22660_), .B0(new_n25344_), .Y(new_n25544_));
  AND2X1   g23108(.A(new_n25544_), .B(pi0208), .Y(new_n25545_));
  AND2X1   g23109(.A(new_n24887_), .B(new_n22959_), .Y(new_n25546_));
  OR3X1    g23110(.A(new_n25546_), .B(new_n25545_), .C(new_n25521_), .Y(new_n25547_));
  MX2X1    g23111(.A(new_n25172_), .B(new_n24964_), .S0(new_n22660_), .Y(new_n25548_));
  AND2X1   g23112(.A(new_n25130_), .B(new_n2933_), .Y(new_n25549_));
  AOI21X1  g23113(.A0(new_n24903_), .A1(new_n2933_), .B0(pi1158), .Y(new_n25550_));
  NOR3X1   g23114(.A(new_n25550_), .B(new_n25549_), .C(new_n12555_), .Y(new_n25551_));
  OAI21X1  g23115(.A0(new_n25551_), .A1(new_n25525_), .B0(new_n24839_), .Y(new_n25552_));
  AND2X1   g23116(.A(new_n25552_), .B(new_n24955_), .Y(new_n25553_));
  OAI22X1  g23117(.A0(new_n25553_), .A1(new_n25541_), .B0(new_n25548_), .B1(new_n25534_), .Y(new_n25554_));
  AOI21X1  g23118(.A0(new_n25547_), .A1(new_n12578_), .B0(new_n25554_), .Y(new_n25555_));
  OR3X1    g23119(.A(new_n25224_), .B(new_n24983_), .C(pi0207), .Y(new_n25556_));
  NOR2X1   g23120(.A(new_n25521_), .B(pi1157), .Y(new_n25557_));
  AOI22X1  g23121(.A0(new_n25557_), .A1(new_n25435_), .B0(new_n25556_), .B1(pi1157), .Y(new_n25558_));
  OR3X1    g23122(.A(new_n25558_), .B(new_n25127_), .C(new_n22959_), .Y(new_n25559_));
  AOI21X1  g23123(.A0(pi1154), .A1(pi0299), .B0(pi0208), .Y(new_n25560_));
  OAI21X1  g23124(.A0(new_n25557_), .A1(new_n25552_), .B0(new_n25560_), .Y(new_n25561_));
  AND2X1   g23125(.A(new_n25561_), .B(pi0214), .Y(new_n25562_));
  AOI21X1  g23126(.A0(new_n25562_), .A1(new_n25559_), .B0(new_n24823_), .Y(new_n25563_));
  OAI21X1  g23127(.A0(new_n25555_), .A1(pi0214), .B0(new_n25563_), .Y(new_n25564_));
  AOI21X1  g23128(.A0(new_n25564_), .A1(new_n25543_), .B0(pi0211), .Y(new_n25565_));
  OAI21X1  g23129(.A0(new_n25565_), .A1(new_n25532_), .B0(pi0219), .Y(new_n25566_));
  NAND3X1  g23130(.A(new_n25531_), .B(new_n25524_), .C(new_n24849_), .Y(new_n25567_));
  AND2X1   g23131(.A(new_n25567_), .B(new_n24823_), .Y(new_n25568_));
  AOI21X1  g23132(.A0(new_n25526_), .A1(new_n2933_), .B0(new_n24986_), .Y(new_n25569_));
  AOI21X1  g23133(.A0(new_n25372_), .A1(new_n25138_), .B0(new_n25569_), .Y(new_n25570_));
  OAI21X1  g23134(.A0(new_n25570_), .A1(new_n12578_), .B0(new_n25524_), .Y(new_n25571_));
  NOR2X1   g23135(.A(new_n25571_), .B(new_n23173_), .Y(new_n25572_));
  NAND4X1  g23136(.A(new_n24999_), .B(new_n24997_), .C(new_n24995_), .D(pi1158), .Y(new_n25573_));
  AOI21X1  g23137(.A0(new_n24929_), .A1(new_n12548_), .B0(new_n22660_), .Y(new_n25574_));
  AND2X1   g23138(.A(new_n25574_), .B(new_n25573_), .Y(new_n25575_));
  AOI21X1  g23139(.A0(new_n25005_), .A1(new_n24901_), .B0(pi0299), .Y(new_n25576_));
  OAI21X1  g23140(.A0(pi1158), .A1(new_n2933_), .B0(new_n22660_), .Y(new_n25577_));
  OAI21X1  g23141(.A0(new_n25577_), .A1(new_n25576_), .B0(pi0208), .Y(new_n25578_));
  OAI21X1  g23142(.A0(new_n25260_), .A1(pi0299), .B0(pi1158), .Y(new_n25579_));
  NAND3X1  g23143(.A(new_n25195_), .B(new_n24839_), .C(pi1156), .Y(new_n25580_));
  AND3X1   g23144(.A(new_n25580_), .B(new_n25579_), .C(new_n22959_), .Y(new_n25581_));
  NOR2X1   g23145(.A(new_n25581_), .B(pi1157), .Y(new_n25582_));
  OAI21X1  g23146(.A0(new_n25578_), .A1(new_n25575_), .B0(new_n25582_), .Y(new_n25583_));
  AND2X1   g23147(.A(new_n12548_), .B(pi0299), .Y(new_n25584_));
  NOR3X1   g23148(.A(new_n25584_), .B(new_n24983_), .C(pi0207), .Y(new_n25585_));
  OR2X1    g23149(.A(new_n25585_), .B(new_n25575_), .Y(new_n25586_));
  INVX1    g23150(.A(new_n25579_), .Y(new_n25587_));
  NOR3X1   g23151(.A(new_n24962_), .B(new_n24911_), .C(pi0299), .Y(new_n25588_));
  INVX1    g23152(.A(new_n25588_), .Y(new_n25589_));
  AOI21X1  g23153(.A0(new_n25204_), .A1(pi1158), .B0(new_n12578_), .Y(new_n25590_));
  AOI21X1  g23154(.A0(new_n25590_), .A1(new_n25589_), .B0(new_n22660_), .Y(new_n25591_));
  NOR2X1   g23155(.A(new_n25591_), .B(new_n25587_), .Y(new_n25592_));
  OAI21X1  g23156(.A0(new_n25592_), .A1(new_n25541_), .B0(new_n23173_), .Y(new_n25593_));
  AOI21X1  g23157(.A0(new_n25586_), .A1(new_n25347_), .B0(new_n25593_), .Y(new_n25594_));
  AOI21X1  g23158(.A0(new_n25594_), .A1(new_n25583_), .B0(new_n25572_), .Y(new_n25595_));
  OAI21X1  g23159(.A0(new_n25595_), .A1(new_n24849_), .B0(new_n25568_), .Y(new_n25596_));
  OR3X1    g23160(.A(new_n25542_), .B(new_n25540_), .C(new_n25535_), .Y(new_n25597_));
  AOI22X1  g23161(.A0(new_n25571_), .A1(new_n24974_), .B0(new_n25597_), .B1(new_n25036_), .Y(new_n25598_));
  OAI21X1  g23162(.A0(new_n25555_), .A1(new_n25033_), .B0(new_n25598_), .Y(new_n25599_));
  AOI21X1  g23163(.A0(new_n25599_), .A1(pi0212), .B0(pi0219), .Y(new_n25600_));
  AOI21X1  g23164(.A0(new_n25600_), .A1(new_n25596_), .B0(po1038), .Y(new_n25601_));
  AOI21X1  g23165(.A0(new_n25601_), .A1(new_n25566_), .B0(new_n25492_), .Y(new_n25602_));
  AND2X1   g23166(.A(new_n3309_), .B(pi0299), .Y(new_n25603_));
  OAI21X1  g23167(.A0(new_n25603_), .A1(new_n24975_), .B0(pi1154), .Y(new_n25604_));
  AND2X1   g23168(.A(pi1145), .B(pi0299), .Y(new_n25605_));
  INVX1    g23169(.A(new_n25605_), .Y(new_n25606_));
  AOI21X1  g23170(.A0(new_n25606_), .A1(new_n24923_), .B0(pi1156), .Y(new_n25607_));
  OAI21X1  g23171(.A0(new_n25603_), .A1(new_n24996_), .B0(new_n12487_), .Y(new_n25608_));
  AOI21X1  g23172(.A0(new_n25606_), .A1(new_n25055_), .B0(new_n12555_), .Y(new_n25609_));
  AOI22X1  g23173(.A0(new_n25609_), .A1(new_n25608_), .B0(new_n25607_), .B1(new_n25604_), .Y(new_n25610_));
  OR2X1    g23174(.A(new_n25610_), .B(new_n22660_), .Y(new_n25611_));
  AND2X1   g23175(.A(pi1157), .B(new_n7937_), .Y(new_n25612_));
  INVX1    g23176(.A(new_n25612_), .Y(new_n25613_));
  OAI21X1  g23177(.A0(new_n25613_), .A1(pi0199), .B0(new_n25576_), .Y(new_n25614_));
  AOI21X1  g23178(.A0(new_n3309_), .A1(pi0299), .B0(pi0207), .Y(new_n25615_));
  AOI21X1  g23179(.A0(new_n25615_), .A1(new_n25614_), .B0(new_n22959_), .Y(new_n25616_));
  OR4X1    g23180(.A(new_n12555_), .B(pi0299), .C(pi0200), .D(new_n7871_), .Y(new_n25617_));
  AOI21X1  g23181(.A0(new_n25204_), .A1(pi1158), .B0(pi1157), .Y(new_n25618_));
  NAND2X1  g23182(.A(new_n25618_), .B(new_n25617_), .Y(new_n25619_));
  OR2X1    g23183(.A(new_n25605_), .B(pi0208), .Y(new_n25620_));
  AOI21X1  g23184(.A0(new_n25619_), .A1(new_n25591_), .B0(new_n25620_), .Y(new_n25621_));
  AOI21X1  g23185(.A0(new_n25616_), .A1(new_n25611_), .B0(new_n25621_), .Y(new_n25622_));
  OAI21X1  g23186(.A0(new_n25538_), .A1(pi1157), .B0(new_n22959_), .Y(new_n25623_));
  OR2X1    g23187(.A(new_n25623_), .B(new_n25552_), .Y(new_n25624_));
  AND3X1   g23188(.A(new_n25624_), .B(new_n25073_), .C(new_n22959_), .Y(new_n25625_));
  NOR2X1   g23189(.A(new_n25077_), .B(new_n22660_), .Y(new_n25626_));
  INVX1    g23190(.A(new_n25626_), .Y(new_n25627_));
  AOI21X1  g23191(.A0(new_n2439_), .A1(pi0299), .B0(pi0207), .Y(new_n25628_));
  AOI21X1  g23192(.A0(new_n25628_), .A1(new_n25614_), .B0(new_n22959_), .Y(new_n25629_));
  AOI21X1  g23193(.A0(new_n25629_), .A1(new_n25627_), .B0(new_n25625_), .Y(new_n25630_));
  MX2X1    g23194(.A(new_n25630_), .B(new_n25622_), .S0(new_n23173_), .Y(new_n25631_));
  OAI21X1  g23195(.A0(new_n25631_), .A1(new_n24849_), .B0(new_n25568_), .Y(new_n25632_));
  OR2X1    g23196(.A(new_n25631_), .B(pi0214), .Y(new_n25633_));
  NAND2X1  g23197(.A(new_n25630_), .B(new_n23173_), .Y(new_n25634_));
  AND3X1   g23198(.A(new_n25624_), .B(new_n25052_), .C(new_n22959_), .Y(new_n25635_));
  OR2X1    g23199(.A(new_n25057_), .B(new_n22660_), .Y(new_n25636_));
  AOI21X1  g23200(.A0(new_n24821_), .A1(pi0299), .B0(pi0207), .Y(new_n25637_));
  AOI21X1  g23201(.A0(new_n25637_), .A1(new_n25614_), .B0(new_n22959_), .Y(new_n25638_));
  AOI21X1  g23202(.A0(new_n25638_), .A1(new_n25636_), .B0(new_n25635_), .Y(new_n25639_));
  AOI21X1  g23203(.A0(new_n25639_), .A1(pi0211), .B0(new_n24849_), .Y(new_n25640_));
  AOI21X1  g23204(.A0(new_n25640_), .A1(new_n25634_), .B0(new_n24823_), .Y(new_n25641_));
  AOI21X1  g23205(.A0(new_n25641_), .A1(new_n25633_), .B0(pi0219), .Y(new_n25642_));
  NOR2X1   g23206(.A(new_n25639_), .B(new_n25162_), .Y(new_n25643_));
  OAI21X1  g23207(.A0(new_n25643_), .A1(new_n25532_), .B0(pi0219), .Y(new_n25644_));
  NAND2X1  g23208(.A(new_n25644_), .B(new_n6489_), .Y(new_n25645_));
  AOI21X1  g23209(.A0(new_n25642_), .A1(new_n25632_), .B0(new_n25645_), .Y(new_n25646_));
  NAND2X1  g23210(.A(new_n25513_), .B(pi0213), .Y(new_n25647_));
  OAI21X1  g23211(.A0(new_n25647_), .A1(new_n25646_), .B0(new_n24866_), .Y(new_n25648_));
  OAI22X1  g23212(.A0(new_n25648_), .A1(new_n25602_), .B0(new_n25518_), .B1(new_n25507_), .Y(new_n25649_));
  MX2X1    g23213(.A(new_n25649_), .B(new_n22579_), .S0(new_n24814_), .Y(po0394));
  INVX1    g23214(.A(new_n24819_), .Y(new_n25651_));
  NOR2X1   g23215(.A(pi1153), .B(pi0211), .Y(new_n25652_));
  AOI21X1  g23216(.A0(new_n25652_), .A1(pi0219), .B0(new_n25651_), .Y(new_n25653_));
  NOR4X1   g23217(.A(new_n25211_), .B(new_n7826_), .C(pi0299), .D(pi0200), .Y(new_n25654_));
  AOI21X1  g23218(.A0(new_n25278_), .A1(new_n24903_), .B0(new_n25654_), .Y(new_n25655_));
  AOI21X1  g23219(.A0(new_n8055_), .A1(new_n12364_), .B0(new_n25655_), .Y(new_n25656_));
  INVX1    g23220(.A(new_n25656_), .Y(new_n25657_));
  AOI21X1  g23221(.A0(new_n25657_), .A1(new_n24849_), .B0(pi0212), .Y(new_n25658_));
  MX2X1    g23222(.A(new_n24961_), .B(new_n24946_), .S0(pi1153), .Y(new_n25659_));
  OAI22X1  g23223(.A0(new_n25659_), .A1(new_n12463_), .B0(new_n25207_), .B1(new_n24917_), .Y(new_n25660_));
  NOR3X1   g23224(.A(new_n24903_), .B(pi0299), .C(new_n22660_), .Y(new_n25661_));
  OAI21X1  g23225(.A0(new_n25661_), .A1(new_n22959_), .B0(new_n24968_), .Y(new_n25662_));
  AOI22X1  g23226(.A0(new_n25662_), .A1(new_n25660_), .B0(new_n25278_), .B1(new_n24903_), .Y(new_n25663_));
  OR2X1    g23227(.A(new_n24870_), .B(new_n2933_), .Y(new_n25664_));
  AND2X1   g23228(.A(new_n25664_), .B(pi0214), .Y(new_n25665_));
  OAI21X1  g23229(.A0(new_n25663_), .A1(pi0299), .B0(new_n25665_), .Y(new_n25666_));
  AND2X1   g23230(.A(new_n25666_), .B(new_n25658_), .Y(new_n25667_));
  AOI21X1  g23231(.A0(pi0207), .A1(new_n7937_), .B0(pi0299), .Y(new_n25668_));
  AND2X1   g23232(.A(new_n24984_), .B(pi0200), .Y(new_n25669_));
  NOR3X1   g23233(.A(new_n25669_), .B(new_n25661_), .C(new_n22959_), .Y(new_n25670_));
  INVX1    g23234(.A(new_n25670_), .Y(new_n25671_));
  OAI21X1  g23235(.A0(new_n25668_), .A1(pi0208), .B0(new_n25671_), .Y(new_n25672_));
  AOI21X1  g23236(.A0(new_n25672_), .A1(new_n25242_), .B0(new_n25033_), .Y(new_n25673_));
  INVX1    g23237(.A(new_n25036_), .Y(new_n25674_));
  NOR3X1   g23238(.A(new_n25656_), .B(new_n25674_), .C(new_n24889_), .Y(new_n25675_));
  OR3X1    g23239(.A(new_n25675_), .B(new_n25673_), .C(new_n24823_), .Y(new_n25676_));
  AOI21X1  g23240(.A0(new_n25663_), .A1(new_n24974_), .B0(new_n25676_), .Y(new_n25677_));
  OR3X1    g23241(.A(new_n25677_), .B(new_n25667_), .C(pi0219), .Y(new_n25678_));
  AND3X1   g23242(.A(new_n5102_), .B(pi1151), .C(new_n2436_), .Y(new_n25679_));
  INVX1    g23243(.A(new_n25672_), .Y(new_n25680_));
  MX2X1    g23244(.A(new_n25680_), .B(new_n25655_), .S0(pi0211), .Y(new_n25681_));
  NOR2X1   g23245(.A(new_n25656_), .B(new_n25188_), .Y(new_n25682_));
  NOR3X1   g23246(.A(new_n25682_), .B(new_n25681_), .C(new_n25241_), .Y(new_n25683_));
  OR2X1    g23247(.A(new_n25683_), .B(new_n8422_), .Y(new_n25684_));
  AND3X1   g23248(.A(new_n25684_), .B(new_n25679_), .C(new_n25678_), .Y(new_n25685_));
  AND3X1   g23249(.A(new_n25204_), .B(new_n25115_), .C(pi1153), .Y(new_n25686_));
  OAI21X1  g23250(.A0(new_n25686_), .A1(new_n24889_), .B0(new_n23173_), .Y(new_n25687_));
  AOI21X1  g23251(.A0(new_n25115_), .A1(new_n8055_), .B0(pi0299), .Y(new_n25688_));
  OR3X1    g23252(.A(new_n25688_), .B(new_n12364_), .C(new_n23173_), .Y(new_n25689_));
  NAND3X1  g23253(.A(new_n25689_), .B(new_n25687_), .C(new_n7996_), .Y(new_n25690_));
  INVX1    g23254(.A(new_n25686_), .Y(new_n25691_));
  NAND3X1  g23255(.A(new_n25691_), .B(new_n25664_), .C(new_n25383_), .Y(new_n25692_));
  AOI21X1  g23256(.A0(new_n25692_), .A1(new_n25690_), .B0(pi0219), .Y(new_n25693_));
  INVX1    g23257(.A(pi1151), .Y(new_n25694_));
  AND3X1   g23258(.A(new_n5102_), .B(new_n25694_), .C(new_n2436_), .Y(new_n25695_));
  AOI21X1  g23259(.A0(new_n25204_), .A1(new_n25115_), .B0(pi0214), .Y(new_n25696_));
  AND2X1   g23260(.A(new_n25696_), .B(new_n24823_), .Y(new_n25697_));
  NOR4X1   g23261(.A(new_n25697_), .B(new_n25688_), .C(new_n9446_), .D(new_n12364_), .Y(new_n25698_));
  OAI21X1  g23262(.A0(new_n25698_), .A1(new_n25109_), .B0(new_n25695_), .Y(new_n25699_));
  OAI21X1  g23263(.A0(new_n25699_), .A1(new_n25693_), .B0(new_n25153_), .Y(new_n25700_));
  NOR2X1   g23264(.A(new_n25700_), .B(new_n25685_), .Y(new_n25701_));
  INVX1    g23265(.A(new_n25233_), .Y(new_n25702_));
  OAI21X1  g23266(.A0(new_n25264_), .A1(new_n8467_), .B0(pi0207), .Y(new_n25703_));
  AND2X1   g23267(.A(new_n25703_), .B(new_n25702_), .Y(new_n25704_));
  AOI21X1  g23268(.A0(pi0207), .A1(pi0200), .B0(pi0199), .Y(new_n25705_));
  OAI21X1  g23269(.A0(new_n25705_), .A1(pi0299), .B0(pi0208), .Y(new_n25706_));
  NOR3X1   g23270(.A(pi0207), .B(pi0200), .C(pi0199), .Y(new_n25707_));
  OAI21X1  g23271(.A0(new_n25707_), .A1(pi0299), .B0(new_n12364_), .Y(new_n25708_));
  INVX1    g23272(.A(new_n25708_), .Y(new_n25709_));
  OAI22X1  g23273(.A0(new_n25709_), .A1(new_n25706_), .B0(new_n25704_), .B1(pi0208), .Y(new_n25710_));
  AND2X1   g23274(.A(new_n25710_), .B(pi0211), .Y(new_n25711_));
  MX2X1    g23275(.A(new_n25199_), .B(new_n9445_), .S0(pi0207), .Y(new_n25712_));
  OAI22X1  g23276(.A0(new_n25712_), .A1(new_n22959_), .B0(new_n25199_), .B1(new_n24986_), .Y(new_n25713_));
  AND3X1   g23277(.A(new_n25713_), .B(new_n25225_), .C(new_n23173_), .Y(new_n25714_));
  OR2X1    g23278(.A(new_n25714_), .B(new_n25711_), .Y(new_n25715_));
  NAND2X1  g23279(.A(new_n24870_), .B(pi0299), .Y(new_n25716_));
  AND2X1   g23280(.A(new_n25713_), .B(new_n25383_), .Y(new_n25717_));
  AOI22X1  g23281(.A0(new_n25717_), .A1(new_n25716_), .B0(new_n25715_), .B1(new_n7996_), .Y(new_n25718_));
  AOI21X1  g23282(.A0(pi0207), .A1(new_n7937_), .B0(new_n25115_), .Y(new_n25719_));
  NOR2X1   g23283(.A(new_n25719_), .B(new_n25275_), .Y(new_n25720_));
  INVX1    g23284(.A(new_n25720_), .Y(new_n25721_));
  AOI21X1  g23285(.A0(new_n25197_), .A1(new_n7827_), .B0(new_n25721_), .Y(new_n25722_));
  AND3X1   g23286(.A(pi1153), .B(pi0299), .C(new_n23173_), .Y(new_n25723_));
  AOI21X1  g23287(.A0(new_n25723_), .A1(new_n25188_), .B0(new_n25722_), .Y(new_n25724_));
  OAI22X1  g23288(.A0(new_n25724_), .A1(new_n25109_), .B0(new_n25718_), .B1(pi0219), .Y(new_n25725_));
  INVX1    g23289(.A(new_n25199_), .Y(new_n25726_));
  NOR3X1   g23290(.A(new_n25243_), .B(new_n25726_), .C(new_n25195_), .Y(new_n25727_));
  OAI22X1  g23291(.A0(new_n25727_), .A1(new_n22959_), .B0(new_n25200_), .B1(new_n24986_), .Y(new_n25728_));
  AND3X1   g23292(.A(new_n25728_), .B(new_n25296_), .C(new_n23173_), .Y(new_n25729_));
  AND3X1   g23293(.A(new_n25728_), .B(new_n25225_), .C(pi0211), .Y(new_n25730_));
  OAI21X1  g23294(.A0(new_n25730_), .A1(new_n25729_), .B0(new_n25383_), .Y(new_n25731_));
  AND3X1   g23295(.A(new_n24903_), .B(new_n2933_), .C(pi0207), .Y(new_n25732_));
  NOR4X1   g23296(.A(new_n25707_), .B(new_n25130_), .C(pi0299), .D(new_n22959_), .Y(new_n25733_));
  NOR2X1   g23297(.A(new_n25733_), .B(new_n25732_), .Y(new_n25734_));
  NAND2X1  g23298(.A(new_n25734_), .B(new_n25689_), .Y(new_n25735_));
  OAI21X1  g23299(.A0(new_n25735_), .A1(new_n25714_), .B0(new_n7996_), .Y(new_n25736_));
  NOR3X1   g23300(.A(new_n25733_), .B(new_n25732_), .C(pi0214), .Y(new_n25737_));
  AOI21X1  g23301(.A0(new_n25737_), .A1(new_n25691_), .B0(pi0212), .Y(new_n25738_));
  AOI21X1  g23302(.A0(new_n25738_), .A1(new_n24849_), .B0(pi0219), .Y(new_n25739_));
  AND3X1   g23303(.A(new_n25739_), .B(new_n25736_), .C(new_n25731_), .Y(new_n25740_));
  OR3X1    g23304(.A(new_n25733_), .B(new_n25732_), .C(new_n8422_), .Y(new_n25741_));
  OAI21X1  g23305(.A0(new_n25741_), .A1(new_n25698_), .B0(new_n25679_), .Y(new_n25742_));
  OAI21X1  g23306(.A0(new_n25742_), .A1(new_n25740_), .B0(pi1152), .Y(new_n25743_));
  AOI21X1  g23307(.A0(new_n25725_), .A1(new_n25695_), .B0(new_n25743_), .Y(new_n25744_));
  OAI21X1  g23308(.A0(new_n25744_), .A1(new_n25701_), .B0(new_n24866_), .Y(new_n25745_));
  AND3X1   g23309(.A(new_n24904_), .B(new_n12487_), .C(pi1153), .Y(new_n25746_));
  OR3X1    g23310(.A(new_n25746_), .B(new_n25228_), .C(new_n25206_), .Y(new_n25747_));
  AND2X1   g23311(.A(new_n25747_), .B(pi0207), .Y(new_n25748_));
  AOI21X1  g23312(.A0(new_n24978_), .A1(new_n22660_), .B0(new_n25748_), .Y(new_n25749_));
  MX2X1    g23313(.A(new_n25749_), .B(new_n25454_), .S0(new_n22959_), .Y(new_n25750_));
  NOR2X1   g23314(.A(new_n25228_), .B(new_n25206_), .Y(new_n25751_));
  AOI21X1  g23315(.A0(new_n12364_), .A1(new_n2933_), .B0(pi1154), .Y(new_n25752_));
  OAI21X1  g23316(.A0(new_n24903_), .A1(pi0299), .B0(new_n25752_), .Y(new_n25753_));
  AND2X1   g23317(.A(new_n25753_), .B(pi0207), .Y(new_n25754_));
  AOI21X1  g23318(.A0(new_n25754_), .A1(new_n25751_), .B0(new_n22959_), .Y(new_n25755_));
  INVX1    g23319(.A(new_n25755_), .Y(new_n25756_));
  AOI21X1  g23320(.A0(new_n25297_), .A1(new_n24933_), .B0(new_n25756_), .Y(new_n25757_));
  INVX1    g23321(.A(new_n25757_), .Y(new_n25758_));
  OAI22X1  g23322(.A0(new_n25758_), .A1(new_n25399_), .B0(new_n24968_), .B1(new_n24954_), .Y(new_n25759_));
  AOI21X1  g23323(.A0(new_n25759_), .A1(new_n23173_), .B0(new_n25533_), .Y(new_n25760_));
  OAI21X1  g23324(.A0(new_n25750_), .A1(new_n23173_), .B0(new_n25760_), .Y(new_n25761_));
  OR2X1    g23325(.A(new_n25750_), .B(new_n25674_), .Y(new_n25762_));
  NAND2X1  g23326(.A(new_n25759_), .B(new_n24974_), .Y(new_n25763_));
  NOR2X1   g23327(.A(new_n24970_), .B(new_n12364_), .Y(new_n25764_));
  NOR2X1   g23328(.A(new_n25764_), .B(new_n25206_), .Y(new_n25765_));
  MX2X1    g23329(.A(new_n25765_), .B(new_n24993_), .S0(new_n22660_), .Y(new_n25766_));
  OAI21X1  g23330(.A0(new_n25766_), .A1(new_n22959_), .B0(new_n25448_), .Y(new_n25767_));
  AOI21X1  g23331(.A0(new_n25767_), .A1(new_n25032_), .B0(new_n24823_), .Y(new_n25768_));
  NAND3X1  g23332(.A(new_n25768_), .B(new_n25763_), .C(new_n25762_), .Y(new_n25769_));
  AOI21X1  g23333(.A0(new_n25769_), .A1(new_n25761_), .B0(pi0219), .Y(new_n25770_));
  INVX1    g23334(.A(new_n25393_), .Y(new_n25771_));
  NOR3X1   g23335(.A(new_n25746_), .B(new_n25206_), .C(new_n7827_), .Y(new_n25772_));
  NOR2X1   g23336(.A(new_n25772_), .B(new_n25771_), .Y(new_n25773_));
  MX2X1    g23337(.A(new_n25773_), .B(new_n25767_), .S0(new_n23173_), .Y(new_n25774_));
  NOR3X1   g23338(.A(new_n25773_), .B(pi0214), .C(pi0212), .Y(new_n25775_));
  NOR2X1   g23339(.A(new_n25775_), .B(po1038), .Y(new_n25776_));
  OAI21X1  g23340(.A0(new_n25774_), .A1(new_n25306_), .B0(new_n25776_), .Y(new_n25777_));
  OAI21X1  g23341(.A0(new_n25777_), .A1(new_n25770_), .B0(pi0209), .Y(new_n25778_));
  AOI22X1  g23342(.A0(new_n25778_), .A1(new_n25745_), .B0(new_n25653_), .B1(new_n25470_), .Y(new_n25779_));
  AND3X1   g23343(.A(new_n25085_), .B(pi1153), .C(new_n23173_), .Y(new_n25780_));
  NOR3X1   g23344(.A(new_n25780_), .B(new_n7962_), .C(pi0219), .Y(new_n25781_));
  OAI21X1  g23345(.A0(new_n25781_), .A1(new_n25651_), .B0(pi1151), .Y(new_n25782_));
  INVX1    g23346(.A(new_n25773_), .Y(new_n25783_));
  AOI21X1  g23347(.A0(new_n24993_), .A1(new_n24984_), .B0(new_n25756_), .Y(new_n25784_));
  NOR2X1   g23348(.A(new_n25784_), .B(new_n25388_), .Y(new_n25785_));
  MX2X1    g23349(.A(new_n25785_), .B(new_n25783_), .S0(pi0211), .Y(new_n25786_));
  AOI21X1  g23350(.A0(new_n25786_), .A1(new_n25188_), .B0(new_n25775_), .Y(new_n25787_));
  OAI21X1  g23351(.A0(new_n25787_), .A1(new_n8422_), .B0(new_n6489_), .Y(new_n25788_));
  MX2X1    g23352(.A(new_n25774_), .B(new_n25773_), .S0(new_n24849_), .Y(new_n25789_));
  AND2X1   g23353(.A(new_n25774_), .B(new_n24849_), .Y(new_n25790_));
  NOR2X1   g23354(.A(new_n25785_), .B(new_n23173_), .Y(new_n25791_));
  AOI21X1  g23355(.A0(new_n25773_), .A1(new_n23173_), .B0(new_n25791_), .Y(new_n25792_));
  OAI21X1  g23356(.A0(new_n25792_), .A1(new_n24849_), .B0(pi0212), .Y(new_n25793_));
  OAI22X1  g23357(.A0(new_n25793_), .A1(new_n25790_), .B0(new_n25789_), .B1(pi0212), .Y(new_n25794_));
  AOI21X1  g23358(.A0(new_n25794_), .A1(new_n8422_), .B0(new_n25788_), .Y(new_n25795_));
  AOI21X1  g23359(.A0(new_n5102_), .A1(new_n2436_), .B0(pi0219), .Y(new_n25796_));
  AOI21X1  g23360(.A0(new_n25780_), .A1(new_n25796_), .B0(pi1151), .Y(new_n25797_));
  AND2X1   g23361(.A(new_n25085_), .B(new_n8422_), .Y(new_n25798_));
  INVX1    g23362(.A(new_n25798_), .Y(new_n25799_));
  AOI21X1  g23363(.A0(new_n25799_), .A1(new_n25783_), .B0(po1038), .Y(new_n25800_));
  OAI21X1  g23364(.A0(new_n25799_), .A1(new_n25774_), .B0(new_n25800_), .Y(new_n25801_));
  AOI21X1  g23365(.A0(new_n25801_), .A1(new_n25797_), .B0(pi1152), .Y(new_n25802_));
  OAI21X1  g23366(.A0(new_n25795_), .A1(new_n25782_), .B0(new_n25802_), .Y(new_n25803_));
  NOR4X1   g23367(.A(new_n24816_), .B(new_n7962_), .C(new_n6489_), .D(pi0219), .Y(new_n25804_));
  MX2X1    g23368(.A(new_n25652_), .B(pi0211), .S0(new_n7996_), .Y(new_n25805_));
  INVX1    g23369(.A(new_n25805_), .Y(new_n25806_));
  AOI21X1  g23370(.A0(new_n25806_), .A1(new_n25804_), .B0(pi1151), .Y(new_n25807_));
  INVX1    g23371(.A(new_n25807_), .Y(new_n25808_));
  AOI21X1  g23372(.A0(new_n25767_), .A1(new_n23173_), .B0(new_n25791_), .Y(new_n25809_));
  NAND2X1  g23373(.A(new_n25809_), .B(pi0214), .Y(new_n25810_));
  AOI21X1  g23374(.A0(new_n25783_), .A1(new_n24849_), .B0(pi0212), .Y(new_n25811_));
  AOI21X1  g23375(.A0(new_n25811_), .A1(new_n25810_), .B0(pi0219), .Y(new_n25812_));
  MX2X1    g23376(.A(new_n25809_), .B(new_n25786_), .S0(pi0214), .Y(new_n25813_));
  OAI21X1  g23377(.A0(new_n25813_), .A1(new_n24823_), .B0(new_n25812_), .Y(new_n25814_));
  AOI21X1  g23378(.A0(new_n25783_), .A1(pi0219), .B0(po1038), .Y(new_n25815_));
  AOI21X1  g23379(.A0(new_n25815_), .A1(new_n25814_), .B0(new_n25808_), .Y(new_n25816_));
  INVX1    g23380(.A(new_n25788_), .Y(new_n25817_));
  INVX1    g23381(.A(new_n25804_), .Y(new_n25818_));
  NOR3X1   g23382(.A(new_n24818_), .B(new_n7963_), .C(new_n6489_), .Y(new_n25819_));
  NOR2X1   g23383(.A(new_n25819_), .B(new_n25694_), .Y(new_n25820_));
  OAI21X1  g23384(.A0(new_n25805_), .A1(new_n25818_), .B0(new_n25820_), .Y(new_n25821_));
  MX2X1    g23385(.A(new_n25809_), .B(new_n25785_), .S0(pi0214), .Y(new_n25822_));
  OAI21X1  g23386(.A0(new_n25822_), .A1(new_n24823_), .B0(new_n25812_), .Y(new_n25823_));
  AOI21X1  g23387(.A0(new_n25823_), .A1(new_n25817_), .B0(new_n25821_), .Y(new_n25824_));
  OR3X1    g23388(.A(new_n25824_), .B(new_n25816_), .C(new_n25153_), .Y(new_n25825_));
  AND3X1   g23389(.A(new_n25825_), .B(new_n25803_), .C(pi0209), .Y(new_n25826_));
  NOR3X1   g23390(.A(new_n25681_), .B(new_n25241_), .C(pi0214), .Y(new_n25827_));
  OR2X1    g23391(.A(new_n25686_), .B(new_n9446_), .Y(new_n25828_));
  OAI21X1  g23392(.A0(new_n25828_), .A1(new_n25656_), .B0(pi0214), .Y(new_n25829_));
  AND2X1   g23393(.A(new_n25829_), .B(pi0212), .Y(new_n25830_));
  INVX1    g23394(.A(new_n25830_), .Y(new_n25831_));
  OAI22X1  g23395(.A0(new_n25831_), .A1(new_n25827_), .B0(new_n25683_), .B1(pi0212), .Y(new_n25832_));
  AND2X1   g23396(.A(pi0299), .B(new_n23173_), .Y(new_n25833_));
  NOR3X1   g23397(.A(new_n25833_), .B(new_n25686_), .C(new_n25656_), .Y(new_n25834_));
  NOR2X1   g23398(.A(new_n25834_), .B(new_n25682_), .Y(new_n25835_));
  INVX1    g23399(.A(new_n25835_), .Y(new_n25836_));
  AOI21X1  g23400(.A0(new_n25836_), .A1(pi0219), .B0(po1038), .Y(new_n25837_));
  INVX1    g23401(.A(new_n25837_), .Y(new_n25838_));
  AOI21X1  g23402(.A0(new_n25832_), .A1(new_n8422_), .B0(new_n25838_), .Y(new_n25839_));
  NAND2X1  g23403(.A(new_n25698_), .B(new_n25696_), .Y(new_n25840_));
  NOR2X1   g23404(.A(new_n25696_), .B(new_n24823_), .Y(new_n25841_));
  AOI21X1  g23405(.A0(new_n25841_), .A1(new_n25828_), .B0(pi0219), .Y(new_n25842_));
  AND2X1   g23406(.A(new_n25204_), .B(new_n25115_), .Y(new_n25843_));
  AOI21X1  g23407(.A0(new_n25723_), .A1(new_n24886_), .B0(new_n25843_), .Y(new_n25844_));
  NAND3X1  g23408(.A(new_n25844_), .B(new_n25842_), .C(new_n25840_), .Y(new_n25845_));
  INVX1    g23409(.A(new_n25843_), .Y(new_n25846_));
  AOI21X1  g23410(.A0(new_n25846_), .A1(pi0219), .B0(po1038), .Y(new_n25847_));
  NAND3X1  g23411(.A(new_n25847_), .B(new_n25845_), .C(new_n25698_), .Y(new_n25848_));
  AOI21X1  g23412(.A0(new_n25848_), .A1(new_n25797_), .B0(pi1152), .Y(new_n25849_));
  OAI21X1  g23413(.A0(new_n25839_), .A1(new_n25782_), .B0(new_n25849_), .Y(new_n25850_));
  OR3X1    g23414(.A(new_n25733_), .B(new_n25732_), .C(new_n25686_), .Y(new_n25851_));
  AOI21X1  g23415(.A0(new_n25728_), .A1(new_n23173_), .B0(new_n25851_), .Y(new_n25852_));
  AOI22X1  g23416(.A0(new_n25852_), .A1(pi0214), .B0(new_n25737_), .B1(new_n25691_), .Y(new_n25853_));
  NOR2X1   g23417(.A(new_n25853_), .B(pi0212), .Y(new_n25854_));
  OAI21X1  g23418(.A0(new_n25854_), .A1(new_n25852_), .B0(pi0219), .Y(new_n25855_));
  AND2X1   g23419(.A(new_n25855_), .B(new_n6489_), .Y(new_n25856_));
  NAND2X1  g23420(.A(new_n25728_), .B(pi0211), .Y(new_n25857_));
  OAI21X1  g23421(.A0(new_n25688_), .A1(new_n12364_), .B0(new_n25857_), .Y(new_n25858_));
  OR3X1    g23422(.A(new_n25733_), .B(new_n25732_), .C(new_n24849_), .Y(new_n25859_));
  OAI21X1  g23423(.A0(new_n25859_), .A1(new_n25858_), .B0(new_n25738_), .Y(new_n25860_));
  INVX1    g23424(.A(new_n25737_), .Y(new_n25861_));
  NOR2X1   g23425(.A(new_n25728_), .B(new_n24849_), .Y(new_n25862_));
  NOR2X1   g23426(.A(new_n25862_), .B(new_n24823_), .Y(new_n25863_));
  OAI21X1  g23427(.A0(new_n25858_), .A1(new_n25861_), .B0(new_n25863_), .Y(new_n25864_));
  NAND3X1  g23428(.A(new_n25864_), .B(new_n25860_), .C(new_n8422_), .Y(new_n25865_));
  AOI21X1  g23429(.A0(new_n25865_), .A1(new_n25856_), .B0(new_n25821_), .Y(new_n25866_));
  INVX1    g23430(.A(new_n25722_), .Y(new_n25867_));
  AOI21X1  g23431(.A0(new_n25867_), .A1(pi0219), .B0(po1038), .Y(new_n25868_));
  OAI21X1  g23432(.A0(new_n25710_), .A1(pi0211), .B0(new_n25717_), .Y(new_n25869_));
  AND3X1   g23433(.A(new_n7996_), .B(pi0299), .C(new_n23173_), .Y(new_n25870_));
  OR2X1    g23434(.A(new_n25870_), .B(pi0219), .Y(new_n25871_));
  AOI21X1  g23435(.A0(new_n25722_), .A1(new_n25086_), .B0(new_n25871_), .Y(new_n25872_));
  NAND2X1  g23436(.A(new_n25872_), .B(new_n25869_), .Y(new_n25873_));
  AOI21X1  g23437(.A0(new_n25873_), .A1(new_n25868_), .B0(new_n25808_), .Y(new_n25874_));
  OR2X1    g23438(.A(new_n25874_), .B(new_n25153_), .Y(new_n25875_));
  OAI21X1  g23439(.A0(new_n25875_), .A1(new_n25866_), .B0(new_n25850_), .Y(new_n25876_));
  OAI21X1  g23440(.A0(new_n25876_), .A1(pi0209), .B0(new_n24815_), .Y(new_n25877_));
  OAI22X1  g23441(.A0(new_n25877_), .A1(new_n25826_), .B0(new_n25779_), .B1(new_n24815_), .Y(new_n25878_));
  MX2X1    g23442(.A(new_n25878_), .B(pi0238), .S0(new_n24814_), .Y(po0395));
  INVX1    g23443(.A(new_n24844_), .Y(new_n25880_));
  NOR2X1   g23444(.A(new_n24929_), .B(new_n25880_), .Y(new_n25881_));
  AOI21X1  g23445(.A0(new_n25881_), .A1(new_n24849_), .B0(pi0212), .Y(new_n25882_));
  AND2X1   g23446(.A(new_n25882_), .B(new_n8422_), .Y(new_n25883_));
  NAND2X1  g23447(.A(pi1158), .B(pi0299), .Y(new_n25884_));
  NAND3X1  g23448(.A(new_n25574_), .B(new_n25573_), .C(new_n22959_), .Y(new_n25885_));
  OAI21X1  g23449(.A0(new_n25884_), .A1(new_n24844_), .B0(new_n25885_), .Y(new_n25886_));
  AOI21X1  g23450(.A0(pi0299), .A1(pi0208), .B0(new_n12578_), .Y(new_n25887_));
  OAI21X1  g23451(.A0(new_n25137_), .A1(new_n24986_), .B0(new_n25887_), .Y(new_n25888_));
  INVX1    g23452(.A(new_n25881_), .Y(new_n25889_));
  AOI21X1  g23453(.A0(new_n25889_), .A1(new_n12578_), .B0(new_n23173_), .Y(new_n25890_));
  AOI22X1  g23454(.A0(new_n25890_), .A1(new_n25888_), .B0(new_n25886_), .B1(new_n23173_), .Y(new_n25891_));
  OAI21X1  g23455(.A0(new_n25891_), .A1(new_n24849_), .B0(new_n25883_), .Y(new_n25892_));
  NAND2X1  g23456(.A(new_n25882_), .B(pi0219), .Y(new_n25893_));
  AOI21X1  g23457(.A0(new_n25889_), .A1(pi0211), .B0(new_n24849_), .Y(new_n25894_));
  NOR3X1   g23458(.A(new_n25169_), .B(new_n25022_), .C(pi0211), .Y(new_n25895_));
  INVX1    g23459(.A(new_n25895_), .Y(new_n25896_));
  AOI21X1  g23460(.A0(new_n25896_), .A1(new_n25894_), .B0(new_n25893_), .Y(new_n25897_));
  AOI21X1  g23461(.A0(new_n25889_), .A1(pi0212), .B0(po1038), .Y(new_n25898_));
  NAND2X1  g23462(.A(new_n25898_), .B(new_n24866_), .Y(new_n25899_));
  NOR2X1   g23463(.A(new_n25899_), .B(new_n25897_), .Y(new_n25900_));
  NOR3X1   g23464(.A(new_n25557_), .B(new_n25527_), .C(pi0208), .Y(new_n25901_));
  INVX1    g23465(.A(new_n25901_), .Y(new_n25902_));
  OAI21X1  g23466(.A0(new_n25902_), .A1(pi0214), .B0(new_n24823_), .Y(new_n25903_));
  OR2X1    g23467(.A(new_n25903_), .B(pi0219), .Y(new_n25904_));
  MX2X1    g23468(.A(new_n25884_), .B(pi1157), .S0(new_n22959_), .Y(new_n25905_));
  NOR2X1   g23469(.A(new_n25905_), .B(new_n25581_), .Y(new_n25906_));
  OR2X1    g23470(.A(new_n25906_), .B(new_n25593_), .Y(new_n25907_));
  INVX1    g23471(.A(new_n25887_), .Y(new_n25908_));
  OAI22X1  g23472(.A0(new_n25908_), .A1(new_n25569_), .B0(new_n25521_), .B1(pi1157), .Y(new_n25909_));
  AOI21X1  g23473(.A0(new_n25909_), .A1(pi0211), .B0(new_n24849_), .Y(new_n25910_));
  AOI21X1  g23474(.A0(new_n25910_), .A1(new_n25907_), .B0(new_n25904_), .Y(new_n25911_));
  OR2X1    g23475(.A(new_n25903_), .B(new_n8422_), .Y(new_n25912_));
  OR2X1    g23476(.A(new_n25901_), .B(new_n23173_), .Y(new_n25913_));
  AOI21X1  g23477(.A0(new_n25902_), .A1(new_n25302_), .B0(new_n24849_), .Y(new_n25914_));
  AOI21X1  g23478(.A0(new_n25914_), .A1(new_n25913_), .B0(new_n25912_), .Y(new_n25915_));
  OAI21X1  g23479(.A0(new_n25901_), .A1(new_n24823_), .B0(new_n6489_), .Y(new_n25916_));
  OR4X1    g23480(.A(new_n25916_), .B(new_n25915_), .C(new_n25911_), .D(new_n24866_), .Y(new_n25917_));
  NAND2X1  g23481(.A(new_n25484_), .B(new_n8422_), .Y(new_n25918_));
  AOI21X1  g23482(.A0(new_n25918_), .A1(new_n25487_), .B0(new_n24815_), .Y(new_n25919_));
  NAND2X1  g23483(.A(new_n25919_), .B(new_n25917_), .Y(new_n25920_));
  AOI21X1  g23484(.A0(new_n25900_), .A1(new_n25892_), .B0(new_n25920_), .Y(new_n25921_));
  NOR2X1   g23485(.A(new_n24887_), .B(new_n23173_), .Y(new_n25922_));
  OAI21X1  g23486(.A0(new_n25623_), .A1(new_n25552_), .B0(new_n25922_), .Y(new_n25923_));
  AOI21X1  g23487(.A0(new_n25923_), .A1(new_n25914_), .B0(new_n25904_), .Y(new_n25924_));
  NAND3X1  g23488(.A(new_n25624_), .B(new_n24890_), .C(new_n23173_), .Y(new_n25925_));
  AND3X1   g23489(.A(new_n25925_), .B(new_n25913_), .C(pi0214), .Y(new_n25926_));
  NOR3X1   g23490(.A(new_n25926_), .B(new_n25903_), .C(new_n8422_), .Y(new_n25927_));
  OR3X1    g23491(.A(new_n25927_), .B(new_n25924_), .C(new_n25916_), .Y(new_n25928_));
  OAI21X1  g23492(.A0(new_n25129_), .A1(new_n24889_), .B0(new_n25894_), .Y(new_n25929_));
  NAND3X1  g23493(.A(new_n25929_), .B(new_n25882_), .C(pi0219), .Y(new_n25930_));
  OAI21X1  g23494(.A0(new_n25172_), .A1(new_n24968_), .B0(new_n25922_), .Y(new_n25931_));
  NAND2X1  g23495(.A(new_n25931_), .B(pi0214), .Y(new_n25932_));
  OAI21X1  g23496(.A0(new_n25932_), .A1(new_n25895_), .B0(new_n25883_), .Y(new_n25933_));
  NAND3X1  g23497(.A(new_n25933_), .B(new_n25930_), .C(new_n25898_), .Y(new_n25934_));
  MX2X1    g23498(.A(new_n25934_), .B(new_n25928_), .S0(pi0209), .Y(new_n25935_));
  NOR2X1   g23499(.A(new_n25337_), .B(new_n6489_), .Y(new_n25936_));
  NAND3X1  g23500(.A(new_n25936_), .B(new_n25335_), .C(new_n24886_), .Y(new_n25937_));
  AND2X1   g23501(.A(new_n25937_), .B(new_n24815_), .Y(new_n25938_));
  AOI21X1  g23502(.A0(new_n25938_), .A1(new_n25935_), .B0(new_n25921_), .Y(new_n25939_));
  MX2X1    g23503(.A(new_n25939_), .B(pi0239), .S0(new_n24814_), .Y(po0396));
  AOI21X1  g23504(.A0(new_n25720_), .A1(new_n6489_), .B0(new_n25847_), .Y(new_n25941_));
  NAND3X1  g23505(.A(new_n8423_), .B(new_n22959_), .C(pi0207), .Y(new_n25942_));
  AND3X1   g23506(.A(new_n25942_), .B(new_n25706_), .C(new_n2933_), .Y(new_n25943_));
  INVX1    g23507(.A(new_n25943_), .Y(new_n25944_));
  OAI21X1  g23508(.A0(new_n25719_), .A1(new_n25275_), .B0(new_n24849_), .Y(new_n25945_));
  NAND2X1  g23509(.A(new_n25945_), .B(new_n24823_), .Y(new_n25946_));
  AND2X1   g23510(.A(new_n25943_), .B(pi0214), .Y(new_n25947_));
  OAI21X1  g23511(.A0(new_n25947_), .A1(new_n25946_), .B0(new_n8422_), .Y(new_n25948_));
  NOR2X1   g23512(.A(new_n25943_), .B(pi0211), .Y(new_n25949_));
  NOR3X1   g23513(.A(new_n25719_), .B(new_n25275_), .C(new_n23173_), .Y(new_n25950_));
  NOR3X1   g23514(.A(new_n25950_), .B(new_n25949_), .C(new_n24849_), .Y(new_n25951_));
  NOR2X1   g23515(.A(new_n25951_), .B(new_n24823_), .Y(new_n25952_));
  AOI21X1  g23516(.A0(new_n25952_), .A1(new_n25944_), .B0(new_n25948_), .Y(new_n25953_));
  OAI21X1  g23517(.A0(new_n25953_), .A1(new_n25941_), .B0(new_n25818_), .Y(new_n25954_));
  INVX1    g23518(.A(pi1149), .Y(new_n25955_));
  AOI21X1  g23519(.A0(new_n5102_), .A1(new_n2436_), .B0(pi0211), .Y(new_n25956_));
  NOR2X1   g23520(.A(new_n25956_), .B(new_n25796_), .Y(new_n25957_));
  NOR2X1   g23521(.A(new_n25957_), .B(new_n24816_), .Y(new_n25958_));
  NOR2X1   g23522(.A(new_n24816_), .B(new_n2933_), .Y(new_n25959_));
  INVX1    g23523(.A(new_n25959_), .Y(new_n25960_));
  NOR3X1   g23524(.A(new_n25960_), .B(new_n24818_), .C(po1038), .Y(new_n25961_));
  NOR3X1   g23525(.A(new_n25211_), .B(new_n25130_), .C(pi0299), .Y(new_n25962_));
  AND2X1   g23526(.A(new_n25962_), .B(new_n6489_), .Y(new_n25963_));
  NOR3X1   g23527(.A(new_n25963_), .B(new_n25961_), .C(new_n25958_), .Y(new_n25964_));
  AOI21X1  g23528(.A0(new_n25964_), .A1(pi1147), .B0(new_n25955_), .Y(new_n25965_));
  OAI21X1  g23529(.A0(new_n25954_), .A1(pi1147), .B0(new_n25965_), .Y(new_n25966_));
  AOI22X1  g23530(.A0(new_n25036_), .A1(pi0212), .B0(new_n24886_), .B1(pi0211), .Y(new_n25967_));
  NOR3X1   g23531(.A(new_n25967_), .B(new_n6489_), .C(pi0219), .Y(new_n25968_));
  NAND2X1  g23532(.A(new_n24998_), .B(new_n7827_), .Y(new_n25969_));
  OAI21X1  g23533(.A0(new_n25260_), .A1(new_n25115_), .B0(new_n25969_), .Y(new_n25970_));
  NOR3X1   g23534(.A(new_n25970_), .B(new_n25707_), .C(pi0299), .Y(new_n25971_));
  AND3X1   g23535(.A(pi0299), .B(pi0214), .C(pi0211), .Y(new_n25972_));
  OAI21X1  g23536(.A0(new_n25972_), .A1(new_n25971_), .B0(new_n24823_), .Y(new_n25973_));
  NAND2X1  g23537(.A(new_n25973_), .B(new_n8422_), .Y(new_n25974_));
  AOI21X1  g23538(.A0(new_n25970_), .A1(new_n2933_), .B0(new_n24849_), .Y(new_n25975_));
  AOI21X1  g23539(.A0(new_n25971_), .A1(new_n24849_), .B0(pi0212), .Y(new_n25976_));
  INVX1    g23540(.A(new_n25976_), .Y(new_n25977_));
  AND2X1   g23541(.A(new_n25970_), .B(new_n2933_), .Y(new_n25978_));
  INVX1    g23542(.A(new_n25978_), .Y(new_n25979_));
  AOI21X1  g23543(.A0(new_n25979_), .A1(new_n23173_), .B0(new_n25971_), .Y(new_n25980_));
  OAI21X1  g23544(.A0(new_n25980_), .A1(new_n24849_), .B0(pi0212), .Y(new_n25981_));
  AOI21X1  g23545(.A0(new_n25970_), .A1(new_n2933_), .B0(pi0214), .Y(new_n25982_));
  OAI22X1  g23546(.A0(new_n25982_), .A1(new_n25981_), .B0(new_n25977_), .B1(new_n25975_), .Y(new_n25983_));
  INVX1    g23547(.A(new_n25983_), .Y(new_n25984_));
  OR3X1    g23548(.A(new_n25975_), .B(new_n25971_), .C(new_n9446_), .Y(new_n25985_));
  AND2X1   g23549(.A(new_n25985_), .B(pi0212), .Y(new_n25986_));
  AOI21X1  g23550(.A0(new_n25986_), .A1(new_n25984_), .B0(new_n25974_), .Y(new_n25987_));
  OR2X1    g23551(.A(new_n25971_), .B(new_n8422_), .Y(new_n25988_));
  AND2X1   g23552(.A(new_n25988_), .B(new_n6489_), .Y(new_n25989_));
  INVX1    g23553(.A(new_n25989_), .Y(new_n25990_));
  NOR2X1   g23554(.A(new_n25990_), .B(new_n25987_), .Y(new_n25991_));
  NOR3X1   g23555(.A(new_n25991_), .B(new_n25968_), .C(pi1147), .Y(new_n25992_));
  INVX1    g23556(.A(pi1147), .Y(new_n25993_));
  OR3X1    g23557(.A(new_n24849_), .B(pi0212), .C(new_n23173_), .Y(new_n25994_));
  OAI21X1  g23558(.A0(pi0214), .A1(pi0211), .B0(pi0212), .Y(new_n25995_));
  AND3X1   g23559(.A(new_n25995_), .B(new_n25994_), .C(new_n8422_), .Y(new_n25996_));
  OR4X1    g23560(.A(new_n25996_), .B(new_n25960_), .C(new_n24818_), .D(po1038), .Y(new_n25997_));
  NOR2X1   g23561(.A(new_n25734_), .B(po1038), .Y(new_n25998_));
  INVX1    g23562(.A(new_n25998_), .Y(new_n25999_));
  NOR3X1   g23563(.A(new_n25996_), .B(new_n24818_), .C(new_n6489_), .Y(new_n26000_));
  INVX1    g23564(.A(new_n26000_), .Y(new_n26001_));
  AND3X1   g23565(.A(new_n26001_), .B(new_n25999_), .C(new_n25997_), .Y(new_n26002_));
  INVX1    g23566(.A(new_n26002_), .Y(new_n26003_));
  OAI21X1  g23567(.A0(new_n26003_), .A1(new_n25993_), .B0(new_n25955_), .Y(new_n26004_));
  OAI21X1  g23568(.A0(new_n26004_), .A1(new_n25992_), .B0(new_n25966_), .Y(new_n26005_));
  AND2X1   g23569(.A(new_n25085_), .B(new_n23173_), .Y(new_n26006_));
  NOR3X1   g23570(.A(new_n26006_), .B(new_n7962_), .C(pi0219), .Y(new_n26007_));
  NOR3X1   g23571(.A(new_n26007_), .B(new_n24818_), .C(new_n6489_), .Y(new_n26008_));
  INVX1    g23572(.A(new_n26008_), .Y(new_n26009_));
  OR2X1    g23573(.A(new_n25655_), .B(pi0211), .Y(new_n26010_));
  AOI21X1  g23574(.A0(new_n25672_), .A1(pi0211), .B0(new_n24849_), .Y(new_n26011_));
  AOI21X1  g23575(.A0(new_n26011_), .A1(new_n26010_), .B0(new_n24877_), .Y(new_n26012_));
  AOI21X1  g23576(.A0(new_n25655_), .A1(new_n24849_), .B0(pi0212), .Y(new_n26013_));
  INVX1    g23577(.A(new_n26013_), .Y(new_n26014_));
  AOI21X1  g23578(.A0(new_n25681_), .A1(pi0214), .B0(new_n26014_), .Y(new_n26015_));
  INVX1    g23579(.A(new_n25681_), .Y(new_n26016_));
  AOI21X1  g23580(.A0(new_n26011_), .A1(new_n26010_), .B0(new_n24823_), .Y(new_n26017_));
  AND2X1   g23581(.A(new_n26017_), .B(new_n26016_), .Y(new_n26018_));
  NOR4X1   g23582(.A(new_n26018_), .B(new_n26015_), .C(new_n26012_), .D(pi0219), .Y(new_n26019_));
  INVX1    g23583(.A(new_n26015_), .Y(new_n26020_));
  AOI21X1  g23584(.A0(new_n26016_), .A1(pi0212), .B0(new_n8422_), .Y(new_n26021_));
  AOI21X1  g23585(.A0(new_n26021_), .A1(new_n26020_), .B0(po1038), .Y(new_n26022_));
  INVX1    g23586(.A(new_n26022_), .Y(new_n26023_));
  OR2X1    g23587(.A(new_n26023_), .B(new_n26019_), .Y(new_n26024_));
  AND3X1   g23588(.A(new_n26024_), .B(new_n26009_), .C(pi1147), .Y(new_n26025_));
  AND3X1   g23589(.A(new_n25115_), .B(new_n11660_), .C(new_n8055_), .Y(new_n26026_));
  NOR2X1   g23590(.A(new_n11660_), .B(pi0219), .Y(new_n26027_));
  AOI21X1  g23591(.A0(new_n26027_), .A1(new_n26006_), .B0(new_n26026_), .Y(new_n26028_));
  INVX1    g23592(.A(new_n26028_), .Y(new_n26029_));
  OAI21X1  g23593(.A0(new_n26029_), .A1(pi1147), .B0(pi1149), .Y(new_n26030_));
  AND2X1   g23594(.A(pi0207), .B(pi0200), .Y(new_n26031_));
  OAI21X1  g23595(.A0(new_n26031_), .A1(new_n24992_), .B0(pi0208), .Y(new_n26032_));
  AOI21X1  g23596(.A0(new_n26032_), .A1(new_n7871_), .B0(new_n25734_), .Y(new_n26033_));
  NOR2X1   g23597(.A(new_n26033_), .B(pi0299), .Y(new_n26034_));
  INVX1    g23598(.A(new_n26034_), .Y(new_n26035_));
  INVX1    g23599(.A(new_n25734_), .Y(new_n26036_));
  OR2X1    g23600(.A(new_n25972_), .B(pi0212), .Y(new_n26037_));
  NOR3X1   g23601(.A(new_n25833_), .B(new_n25733_), .C(new_n25732_), .Y(new_n26038_));
  NOR2X1   g23602(.A(new_n26038_), .B(new_n25737_), .Y(new_n26039_));
  INVX1    g23603(.A(new_n9446_), .Y(new_n26040_));
  OAI21X1  g23604(.A0(new_n26040_), .A1(pi0214), .B0(pi0212), .Y(new_n26041_));
  OAI22X1  g23605(.A0(new_n26041_), .A1(new_n26039_), .B0(new_n26037_), .B1(new_n26036_), .Y(new_n26042_));
  OAI21X1  g23606(.A0(new_n26034_), .A1(new_n26042_), .B0(new_n8422_), .Y(new_n26043_));
  OR2X1    g23607(.A(new_n26043_), .B(pi0211), .Y(new_n26044_));
  NOR4X1   g23608(.A(new_n25733_), .B(new_n25732_), .C(new_n9446_), .D(new_n24849_), .Y(new_n26045_));
  NOR4X1   g23609(.A(new_n25833_), .B(new_n25733_), .C(new_n25732_), .D(pi0214), .Y(new_n26046_));
  OR3X1    g23610(.A(new_n26046_), .B(new_n26045_), .C(new_n24823_), .Y(new_n26047_));
  NOR3X1   g23611(.A(new_n26038_), .B(new_n25737_), .C(pi0212), .Y(new_n26048_));
  NOR2X1   g23612(.A(new_n26048_), .B(pi0219), .Y(new_n26049_));
  AND2X1   g23613(.A(new_n26049_), .B(new_n26047_), .Y(new_n26050_));
  INVX1    g23614(.A(new_n25833_), .Y(new_n26051_));
  NOR2X1   g23615(.A(new_n24818_), .B(po1038), .Y(new_n26052_));
  INVX1    g23616(.A(new_n26052_), .Y(new_n26053_));
  AOI21X1  g23617(.A0(new_n26051_), .A1(pi0219), .B0(new_n26053_), .Y(new_n26054_));
  INVX1    g23618(.A(new_n26054_), .Y(new_n26055_));
  AOI21X1  g23619(.A0(new_n26055_), .A1(new_n25999_), .B0(new_n26050_), .Y(new_n26056_));
  AND3X1   g23620(.A(new_n26056_), .B(new_n26044_), .C(new_n26035_), .Y(new_n26057_));
  OR2X1    g23621(.A(new_n26057_), .B(new_n25819_), .Y(new_n26058_));
  NAND3X1  g23622(.A(new_n26058_), .B(new_n25955_), .C(pi1147), .Y(new_n26059_));
  OAI21X1  g23623(.A0(new_n26030_), .A1(new_n26025_), .B0(new_n26059_), .Y(new_n26060_));
  MX2X1    g23624(.A(new_n26060_), .B(new_n26005_), .S0(pi1148), .Y(new_n26061_));
  AND2X1   g23625(.A(pi1146), .B(pi0211), .Y(new_n26062_));
  MX2X1    g23626(.A(new_n3140_), .B(new_n3309_), .S0(pi0211), .Y(new_n26063_));
  INVX1    g23627(.A(new_n26063_), .Y(new_n26064_));
  MX2X1    g23628(.A(new_n26062_), .B(new_n26064_), .S0(pi0214), .Y(new_n26065_));
  AOI22X1  g23629(.A0(new_n26065_), .A1(pi0212), .B0(new_n26062_), .B1(new_n24886_), .Y(new_n26066_));
  AND2X1   g23630(.A(pi1145), .B(new_n23173_), .Y(new_n26067_));
  OAI22X1  g23631(.A0(new_n26067_), .A1(new_n8422_), .B0(new_n5103_), .B1(pi0057), .Y(new_n26068_));
  AOI21X1  g23632(.A0(new_n26066_), .A1(new_n25306_), .B0(new_n26068_), .Y(new_n26069_));
  NOR4X1   g23633(.A(new_n24816_), .B(new_n7996_), .C(pi0219), .D(pi0211), .Y(new_n26070_));
  AND2X1   g23634(.A(new_n26070_), .B(po1038), .Y(new_n26071_));
  NOR3X1   g23635(.A(new_n26071_), .B(new_n26069_), .C(new_n25993_), .Y(new_n26072_));
  INVX1    g23636(.A(new_n26072_), .Y(new_n26073_));
  AOI21X1  g23637(.A0(new_n25605_), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n26074_));
  OR3X1    g23638(.A(new_n26074_), .B(new_n24818_), .C(po1038), .Y(new_n26075_));
  NOR2X1   g23639(.A(new_n26063_), .B(new_n2933_), .Y(new_n26076_));
  OAI21X1  g23640(.A0(new_n26076_), .A1(new_n26036_), .B0(new_n7996_), .Y(new_n26077_));
  AND3X1   g23641(.A(pi1146), .B(pi0299), .C(pi0211), .Y(new_n26078_));
  NOR4X1   g23642(.A(new_n26078_), .B(new_n25833_), .C(new_n25733_), .D(new_n25732_), .Y(new_n26079_));
  OR2X1    g23643(.A(new_n26079_), .B(new_n25086_), .Y(new_n26080_));
  AOI21X1  g23644(.A0(new_n26036_), .A1(new_n24816_), .B0(pi0219), .Y(new_n26081_));
  AND3X1   g23645(.A(new_n26081_), .B(new_n26080_), .C(new_n26077_), .Y(new_n26082_));
  AOI21X1  g23646(.A0(new_n26075_), .A1(new_n25999_), .B0(new_n26082_), .Y(new_n26083_));
  INVX1    g23647(.A(pi1148), .Y(new_n26084_));
  NOR4X1   g23648(.A(new_n25970_), .B(new_n25707_), .C(po1038), .D(pi0299), .Y(new_n26085_));
  INVX1    g23649(.A(new_n26085_), .Y(new_n26086_));
  OR3X1    g23650(.A(new_n26066_), .B(new_n23385_), .C(new_n2933_), .Y(new_n26087_));
  OAI21X1  g23651(.A0(new_n26075_), .A1(new_n8422_), .B0(new_n26087_), .Y(new_n26088_));
  NOR3X1   g23652(.A(new_n26088_), .B(new_n26069_), .C(pi1147), .Y(new_n26089_));
  AOI21X1  g23653(.A0(new_n26089_), .A1(new_n26086_), .B0(new_n26084_), .Y(new_n26090_));
  OAI21X1  g23654(.A0(new_n26083_), .A1(new_n26073_), .B0(new_n26090_), .Y(new_n26091_));
  INVX1    g23655(.A(new_n26077_), .Y(new_n26092_));
  AOI21X1  g23656(.A0(new_n9446_), .A1(new_n3140_), .B0(new_n25086_), .Y(new_n26093_));
  NOR2X1   g23657(.A(new_n26034_), .B(pi0219), .Y(new_n26094_));
  OAI21X1  g23658(.A0(new_n26093_), .A1(new_n26092_), .B0(new_n26094_), .Y(new_n26095_));
  NOR4X1   g23659(.A(new_n25306_), .B(new_n3309_), .C(new_n2933_), .D(pi0211), .Y(new_n26096_));
  AOI21X1  g23660(.A0(new_n26033_), .A1(new_n25110_), .B0(new_n26096_), .Y(new_n26097_));
  AOI21X1  g23661(.A0(new_n26097_), .A1(new_n26095_), .B0(po1038), .Y(new_n26098_));
  NOR2X1   g23662(.A(new_n26089_), .B(pi1148), .Y(new_n26099_));
  OAI21X1  g23663(.A0(new_n26098_), .A1(new_n26073_), .B0(new_n26099_), .Y(new_n26100_));
  AOI21X1  g23664(.A0(new_n26100_), .A1(new_n26091_), .B0(pi1149), .Y(new_n26101_));
  AOI21X1  g23665(.A0(new_n25655_), .A1(pi0219), .B0(po1038), .Y(new_n26102_));
  INVX1    g23666(.A(new_n26102_), .Y(new_n26103_));
  NAND2X1  g23667(.A(new_n26103_), .B(new_n26075_), .Y(new_n26104_));
  NAND2X1  g23668(.A(new_n25672_), .B(new_n23173_), .Y(new_n26105_));
  AND2X1   g23669(.A(pi1146), .B(pi0299), .Y(new_n26106_));
  OAI22X1  g23670(.A0(new_n25671_), .A1(pi0299), .B0(new_n24917_), .B1(new_n25880_), .Y(new_n26107_));
  OAI21X1  g23671(.A0(new_n26107_), .A1(new_n26106_), .B0(pi0211), .Y(new_n26108_));
  AND3X1   g23672(.A(new_n26108_), .B(new_n26105_), .C(pi0214), .Y(new_n26109_));
  NOR2X1   g23673(.A(new_n26109_), .B(new_n26014_), .Y(new_n26110_));
  AND3X1   g23674(.A(new_n26108_), .B(new_n26105_), .C(new_n24849_), .Y(new_n26111_));
  OAI21X1  g23675(.A0(new_n26063_), .A1(new_n2933_), .B0(pi0214), .Y(new_n26112_));
  OAI21X1  g23676(.A0(new_n26112_), .A1(new_n26107_), .B0(pi0212), .Y(new_n26113_));
  OAI21X1  g23677(.A0(new_n26113_), .A1(new_n26111_), .B0(new_n8422_), .Y(new_n26114_));
  OAI21X1  g23678(.A0(new_n26114_), .A1(new_n26110_), .B0(new_n26104_), .Y(new_n26115_));
  NOR4X1   g23679(.A(new_n26088_), .B(new_n26069_), .C(new_n26026_), .D(pi1147), .Y(new_n26116_));
  OR2X1    g23680(.A(new_n26116_), .B(pi1148), .Y(new_n26117_));
  AOI21X1  g23681(.A0(new_n26115_), .A1(new_n26072_), .B0(new_n26117_), .Y(new_n26118_));
  NOR2X1   g23682(.A(new_n26069_), .B(pi1147), .Y(new_n26119_));
  INVX1    g23683(.A(new_n26119_), .Y(new_n26120_));
  OR3X1    g23684(.A(new_n25943_), .B(new_n24816_), .C(pi0211), .Y(new_n26121_));
  AOI21X1  g23685(.A0(new_n25720_), .A1(new_n25162_), .B0(new_n8422_), .Y(new_n26122_));
  AOI21X1  g23686(.A0(new_n26122_), .A1(new_n26121_), .B0(po1038), .Y(new_n26123_));
  NAND2X1  g23687(.A(new_n26123_), .B(new_n8423_), .Y(new_n26124_));
  NAND2X1  g23688(.A(new_n26124_), .B(new_n26075_), .Y(new_n26125_));
  NOR2X1   g23689(.A(new_n26078_), .B(new_n25720_), .Y(new_n26126_));
  NOR2X1   g23690(.A(new_n26126_), .B(new_n25946_), .Y(new_n26127_));
  OR2X1    g23691(.A(new_n25943_), .B(new_n24823_), .Y(new_n26128_));
  NOR2X1   g23692(.A(new_n26065_), .B(new_n25720_), .Y(new_n26129_));
  OAI21X1  g23693(.A0(new_n26129_), .A1(new_n26128_), .B0(new_n8422_), .Y(new_n26130_));
  OR2X1    g23694(.A(new_n26130_), .B(new_n26127_), .Y(new_n26131_));
  AOI21X1  g23695(.A0(new_n26131_), .A1(new_n26125_), .B0(new_n26120_), .Y(new_n26132_));
  INVX1    g23696(.A(new_n25962_), .Y(new_n26133_));
  AOI21X1  g23697(.A0(new_n26133_), .A1(pi0219), .B0(po1038), .Y(new_n26134_));
  INVX1    g23698(.A(new_n26134_), .Y(new_n26135_));
  OR2X1    g23699(.A(new_n25962_), .B(new_n23173_), .Y(new_n26136_));
  AND2X1   g23700(.A(pi0299), .B(pi0214), .Y(new_n26137_));
  NOR2X1   g23701(.A(new_n26137_), .B(new_n25962_), .Y(new_n26138_));
  NOR2X1   g23702(.A(new_n26138_), .B(pi0212), .Y(new_n26139_));
  NAND2X1  g23703(.A(new_n26139_), .B(new_n26136_), .Y(new_n26140_));
  AOI21X1  g23704(.A0(new_n26133_), .A1(new_n2933_), .B0(new_n24823_), .Y(new_n26141_));
  NOR2X1   g23705(.A(new_n25995_), .B(new_n2933_), .Y(new_n26142_));
  INVX1    g23706(.A(new_n26142_), .Y(new_n26143_));
  AOI21X1  g23707(.A0(new_n26143_), .A1(new_n26141_), .B0(pi0219), .Y(new_n26144_));
  AOI21X1  g23708(.A0(new_n26144_), .A1(new_n26140_), .B0(new_n26135_), .Y(new_n26145_));
  NOR3X1   g23709(.A(new_n26145_), .B(new_n26088_), .C(new_n26073_), .Y(new_n26146_));
  NOR3X1   g23710(.A(new_n26146_), .B(new_n26132_), .C(new_n26084_), .Y(new_n26147_));
  OR2X1    g23711(.A(new_n26147_), .B(new_n26118_), .Y(new_n26148_));
  AOI21X1  g23712(.A0(new_n26148_), .A1(pi1149), .B0(new_n26101_), .Y(new_n26149_));
  OAI21X1  g23713(.A0(new_n26149_), .A1(pi0213), .B0(pi0209), .Y(new_n26150_));
  AOI21X1  g23714(.A0(new_n26061_), .A1(pi0213), .B0(new_n26150_), .Y(new_n26151_));
  AOI21X1  g23715(.A0(pi1146), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n26152_));
  AND3X1   g23716(.A(new_n3309_), .B(new_n7937_), .C(pi0199), .Y(new_n26153_));
  NOR3X1   g23717(.A(new_n26153_), .B(new_n26152_), .C(pi0299), .Y(new_n26154_));
  INVX1    g23718(.A(new_n26154_), .Y(new_n26155_));
  NOR4X1   g23719(.A(new_n26153_), .B(new_n26152_), .C(pi0299), .D(pi0207), .Y(new_n26156_));
  AOI21X1  g23720(.A0(pi1145), .A1(pi0199), .B0(pi0200), .Y(new_n26157_));
  OAI21X1  g23721(.A0(new_n3140_), .A1(pi0199), .B0(new_n26157_), .Y(new_n26158_));
  OAI21X1  g23722(.A0(new_n3309_), .A1(pi0199), .B0(pi0200), .Y(new_n26159_));
  AND3X1   g23723(.A(new_n26159_), .B(new_n26158_), .C(new_n24839_), .Y(new_n26160_));
  NOR3X1   g23724(.A(new_n26160_), .B(new_n26156_), .C(new_n26106_), .Y(new_n26161_));
  OAI22X1  g23725(.A0(new_n26161_), .A1(new_n22959_), .B0(new_n26155_), .B1(new_n25880_), .Y(new_n26162_));
  OR2X1    g23726(.A(new_n26162_), .B(pi0299), .Y(new_n26163_));
  AND2X1   g23727(.A(new_n26163_), .B(pi0211), .Y(new_n26164_));
  INVX1    g23728(.A(new_n26164_), .Y(new_n26165_));
  AND2X1   g23729(.A(new_n26157_), .B(new_n26156_), .Y(new_n26166_));
  OR3X1    g23730(.A(new_n26166_), .B(new_n26161_), .C(new_n22959_), .Y(new_n26167_));
  NOR3X1   g23731(.A(new_n26157_), .B(new_n26152_), .C(pi0299), .Y(new_n26168_));
  INVX1    g23732(.A(new_n26168_), .Y(new_n26169_));
  OAI21X1  g23733(.A0(new_n26169_), .A1(new_n25880_), .B0(new_n26167_), .Y(new_n26170_));
  OAI21X1  g23734(.A0(new_n26170_), .A1(pi0299), .B0(pi0214), .Y(new_n26171_));
  AOI21X1  g23735(.A0(new_n26171_), .A1(new_n26165_), .B0(new_n24823_), .Y(new_n26172_));
  AND2X1   g23736(.A(new_n26163_), .B(new_n25032_), .Y(new_n26173_));
  INVX1    g23737(.A(new_n26160_), .Y(new_n26174_));
  AOI22X1  g23738(.A0(new_n26174_), .A1(new_n25116_), .B0(new_n26155_), .B1(new_n7827_), .Y(new_n26175_));
  OR4X1    g23739(.A(new_n26175_), .B(new_n26173_), .C(new_n26172_), .D(pi0219), .Y(new_n26176_));
  AOI22X1  g23740(.A0(new_n26169_), .A1(new_n7827_), .B0(new_n26174_), .B1(new_n25116_), .Y(new_n26177_));
  AOI21X1  g23741(.A0(new_n26177_), .A1(new_n24816_), .B0(new_n26176_), .Y(new_n26178_));
  NOR2X1   g23742(.A(new_n26170_), .B(pi0299), .Y(new_n26179_));
  AOI21X1  g23743(.A0(new_n26163_), .A1(new_n23173_), .B0(new_n26175_), .Y(new_n26180_));
  AND2X1   g23744(.A(new_n26180_), .B(pi0214), .Y(new_n26181_));
  OR2X1    g23745(.A(new_n26181_), .B(new_n26179_), .Y(new_n26182_));
  AOI21X1  g23746(.A0(new_n26177_), .A1(new_n24849_), .B0(pi0212), .Y(new_n26183_));
  AOI22X1  g23747(.A0(new_n26183_), .A1(new_n26171_), .B0(new_n26182_), .B1(pi0212), .Y(new_n26184_));
  INVX1    g23748(.A(new_n26177_), .Y(new_n26185_));
  AOI21X1  g23749(.A0(new_n26185_), .A1(pi0219), .B0(po1038), .Y(new_n26186_));
  OAI21X1  g23750(.A0(new_n26184_), .A1(pi0219), .B0(new_n26186_), .Y(new_n26187_));
  OR2X1    g23751(.A(new_n26187_), .B(new_n26178_), .Y(new_n26188_));
  NOR2X1   g23752(.A(new_n25968_), .B(pi1147), .Y(new_n26189_));
  AOI21X1  g23753(.A0(new_n26175_), .A1(new_n25162_), .B0(new_n8422_), .Y(new_n26190_));
  NAND3X1  g23754(.A(new_n26163_), .B(new_n25188_), .C(new_n23173_), .Y(new_n26191_));
  AOI21X1  g23755(.A0(new_n26191_), .A1(new_n26190_), .B0(po1038), .Y(new_n26192_));
  AND2X1   g23756(.A(new_n26192_), .B(new_n26176_), .Y(new_n26193_));
  OR2X1    g23757(.A(new_n26000_), .B(new_n25993_), .Y(new_n26194_));
  OAI21X1  g23758(.A0(new_n26194_), .A1(new_n26193_), .B0(new_n25955_), .Y(new_n26195_));
  AOI21X1  g23759(.A0(new_n26189_), .A1(new_n26188_), .B0(new_n26195_), .Y(new_n26196_));
  NOR2X1   g23760(.A(new_n25804_), .B(pi1147), .Y(new_n26197_));
  OR3X1    g23761(.A(new_n26175_), .B(new_n25959_), .C(pi0219), .Y(new_n26198_));
  OAI21X1  g23762(.A0(new_n25957_), .A1(new_n24816_), .B0(pi1147), .Y(new_n26199_));
  AOI21X1  g23763(.A0(new_n26198_), .A1(new_n26192_), .B0(new_n26199_), .Y(new_n26200_));
  OR2X1    g23764(.A(new_n26200_), .B(new_n25955_), .Y(new_n26201_));
  AOI21X1  g23765(.A0(new_n26197_), .A1(new_n26187_), .B0(new_n26201_), .Y(new_n26202_));
  OR3X1    g23766(.A(new_n26202_), .B(new_n26196_), .C(new_n26084_), .Y(new_n26203_));
  AND3X1   g23767(.A(new_n5102_), .B(new_n25993_), .C(new_n2436_), .Y(new_n26204_));
  NOR3X1   g23768(.A(new_n26175_), .B(new_n26164_), .C(new_n24849_), .Y(new_n26205_));
  AND2X1   g23769(.A(new_n26163_), .B(new_n23173_), .Y(new_n26206_));
  NOR3X1   g23770(.A(new_n26206_), .B(new_n26175_), .C(pi0214), .Y(new_n26207_));
  OR3X1    g23771(.A(new_n26207_), .B(new_n26205_), .C(new_n24823_), .Y(new_n26208_));
  OAI21X1  g23772(.A0(new_n26175_), .A1(pi0214), .B0(new_n24823_), .Y(new_n26209_));
  OR2X1    g23773(.A(new_n26209_), .B(new_n26180_), .Y(new_n26210_));
  AND3X1   g23774(.A(new_n26210_), .B(new_n26208_), .C(new_n8422_), .Y(new_n26211_));
  INVX1    g23775(.A(new_n26211_), .Y(new_n26212_));
  AND2X1   g23776(.A(new_n26212_), .B(new_n26193_), .Y(new_n26213_));
  OR2X1    g23777(.A(new_n26213_), .B(new_n25819_), .Y(new_n26214_));
  AOI22X1  g23778(.A0(new_n26214_), .A1(pi1147), .B0(new_n26204_), .B1(new_n26177_), .Y(new_n26215_));
  AOI21X1  g23779(.A0(new_n26212_), .A1(new_n26192_), .B0(new_n26008_), .Y(new_n26216_));
  INVX1    g23780(.A(new_n26070_), .Y(new_n26217_));
  INVX1    g23781(.A(new_n26204_), .Y(new_n26218_));
  OAI22X1  g23782(.A0(new_n26218_), .A1(new_n26185_), .B0(new_n26217_), .B1(pi1147), .Y(new_n26219_));
  NAND2X1  g23783(.A(new_n26070_), .B(new_n11660_), .Y(new_n26220_));
  OAI21X1  g23784(.A0(new_n26220_), .A1(new_n26170_), .B0(new_n26219_), .Y(new_n26221_));
  OAI21X1  g23785(.A0(new_n26216_), .A1(new_n25993_), .B0(new_n26221_), .Y(new_n26222_));
  AOI21X1  g23786(.A0(new_n26222_), .A1(pi1149), .B0(pi1148), .Y(new_n26223_));
  OAI21X1  g23787(.A0(new_n26215_), .A1(pi1149), .B0(new_n26223_), .Y(new_n26224_));
  NAND3X1  g23788(.A(new_n26224_), .B(new_n26203_), .C(pi0213), .Y(new_n26225_));
  AOI21X1  g23789(.A0(new_n26177_), .A1(new_n24816_), .B0(new_n8422_), .Y(new_n26226_));
  AOI21X1  g23790(.A0(new_n26177_), .A1(new_n25188_), .B0(new_n24817_), .Y(new_n26227_));
  OR2X1    g23791(.A(new_n25605_), .B(pi0211), .Y(new_n26228_));
  AOI21X1  g23792(.A0(new_n26170_), .A1(new_n2933_), .B0(new_n26228_), .Y(new_n26229_));
  OAI21X1  g23793(.A0(new_n26229_), .A1(new_n26227_), .B0(new_n26226_), .Y(new_n26230_));
  OR2X1    g23794(.A(new_n26177_), .B(new_n26078_), .Y(new_n26231_));
  AOI21X1  g23795(.A0(new_n26185_), .A1(new_n24849_), .B0(pi0212), .Y(new_n26232_));
  AOI21X1  g23796(.A0(new_n26232_), .A1(new_n26231_), .B0(pi0219), .Y(new_n26233_));
  AOI21X1  g23797(.A0(new_n26170_), .A1(new_n2933_), .B0(new_n26112_), .Y(new_n26234_));
  OAI21X1  g23798(.A0(new_n26231_), .A1(pi0214), .B0(pi0212), .Y(new_n26235_));
  OAI21X1  g23799(.A0(new_n26235_), .A1(new_n26234_), .B0(new_n26233_), .Y(new_n26236_));
  NAND3X1  g23800(.A(new_n26236_), .B(new_n26230_), .C(new_n6489_), .Y(new_n26237_));
  NOR2X1   g23801(.A(new_n26162_), .B(new_n26112_), .Y(new_n26238_));
  OAI22X1  g23802(.A0(new_n26238_), .A1(new_n26173_), .B0(new_n26165_), .B1(new_n25603_), .Y(new_n26239_));
  OR4X1    g23803(.A(new_n26162_), .B(new_n26078_), .C(new_n25833_), .D(pi0214), .Y(new_n26240_));
  AND3X1   g23804(.A(new_n26240_), .B(new_n26239_), .C(pi0212), .Y(new_n26241_));
  NAND2X1  g23805(.A(new_n26233_), .B(new_n26210_), .Y(new_n26242_));
  INVX1    g23806(.A(new_n25603_), .Y(new_n26243_));
  NAND4X1  g23807(.A(new_n26163_), .B(new_n26243_), .C(new_n25188_), .D(new_n23173_), .Y(new_n26244_));
  AOI21X1  g23808(.A0(new_n26244_), .A1(new_n26190_), .B0(po1038), .Y(new_n26245_));
  OAI21X1  g23809(.A0(new_n26242_), .A1(new_n26241_), .B0(new_n26245_), .Y(new_n26246_));
  AOI22X1  g23810(.A0(new_n26246_), .A1(new_n26072_), .B0(new_n26237_), .B1(new_n26119_), .Y(new_n26247_));
  AOI21X1  g23811(.A0(new_n26247_), .A1(new_n24815_), .B0(pi0209), .Y(new_n26248_));
  AOI21X1  g23812(.A0(new_n26248_), .A1(new_n26225_), .B0(new_n26151_), .Y(new_n26249_));
  MX2X1    g23813(.A(new_n26249_), .B(pi0240), .S0(new_n24814_), .Y(po0397));
  OR2X1    g23814(.A(new_n26070_), .B(new_n6489_), .Y(new_n26251_));
  AND2X1   g23815(.A(new_n26251_), .B(pi1151), .Y(new_n26252_));
  AOI21X1  g23816(.A0(new_n26070_), .A1(new_n25728_), .B0(new_n25851_), .Y(new_n26253_));
  OAI21X1  g23817(.A0(new_n26253_), .A1(new_n25153_), .B0(new_n6489_), .Y(new_n26254_));
  AND2X1   g23818(.A(new_n26006_), .B(new_n24884_), .Y(new_n26255_));
  OR2X1    g23819(.A(new_n26255_), .B(new_n25656_), .Y(new_n26256_));
  AOI22X1  g23820(.A0(new_n26256_), .A1(new_n26252_), .B0(new_n25695_), .B1(new_n25686_), .Y(new_n26257_));
  NAND3X1  g23821(.A(new_n25722_), .B(new_n25695_), .C(pi1152), .Y(new_n26258_));
  OAI21X1  g23822(.A0(new_n26257_), .A1(pi1152), .B0(new_n26258_), .Y(new_n26259_));
  AOI21X1  g23823(.A0(new_n26254_), .A1(new_n26252_), .B0(new_n26259_), .Y(new_n26260_));
  OR2X1    g23824(.A(new_n26260_), .B(pi1150), .Y(new_n26261_));
  NOR2X1   g23825(.A(new_n25804_), .B(new_n25694_), .Y(new_n26262_));
  INVX1    g23826(.A(new_n26262_), .Y(new_n26263_));
  AOI21X1  g23827(.A0(new_n25691_), .A1(pi0219), .B0(po1038), .Y(new_n26264_));
  INVX1    g23828(.A(new_n26264_), .Y(new_n26265_));
  OAI21X1  g23829(.A0(new_n25728_), .A1(new_n24849_), .B0(new_n25738_), .Y(new_n26266_));
  AND2X1   g23830(.A(new_n26266_), .B(new_n8422_), .Y(new_n26267_));
  INVX1    g23831(.A(new_n26267_), .Y(new_n26268_));
  OAI21X1  g23832(.A0(new_n25728_), .A1(pi0214), .B0(pi0212), .Y(new_n26269_));
  AOI21X1  g23833(.A0(new_n25852_), .A1(pi0214), .B0(new_n26269_), .Y(new_n26270_));
  OAI21X1  g23834(.A0(new_n26270_), .A1(new_n26268_), .B0(pi1152), .Y(new_n26271_));
  INVX1    g23835(.A(new_n25658_), .Y(new_n26272_));
  AOI21X1  g23836(.A0(new_n25672_), .A1(new_n25242_), .B0(pi0299), .Y(new_n26273_));
  AOI21X1  g23837(.A0(new_n25680_), .A1(new_n24849_), .B0(new_n24823_), .Y(new_n26274_));
  OAI21X1  g23838(.A0(new_n26016_), .A1(new_n24849_), .B0(new_n26274_), .Y(new_n26275_));
  AOI21X1  g23839(.A0(new_n26275_), .A1(new_n26272_), .B0(new_n26273_), .Y(new_n26276_));
  AOI21X1  g23840(.A0(new_n25655_), .A1(pi0219), .B0(pi1152), .Y(new_n26277_));
  OAI21X1  g23841(.A0(new_n26276_), .A1(pi0219), .B0(new_n26277_), .Y(new_n26278_));
  AOI22X1  g23842(.A0(new_n26278_), .A1(new_n26271_), .B0(new_n26265_), .B1(new_n25999_), .Y(new_n26279_));
  INVX1    g23843(.A(pi1150), .Y(new_n26280_));
  NOR2X1   g23844(.A(new_n25968_), .B(pi1151), .Y(new_n26281_));
  NOR3X1   g23845(.A(new_n25696_), .B(new_n25688_), .C(pi0212), .Y(new_n26282_));
  AOI21X1  g23846(.A0(new_n26282_), .A1(new_n26051_), .B0(pi0219), .Y(new_n26283_));
  INVX1    g23847(.A(new_n26283_), .Y(new_n26284_));
  OAI21X1  g23848(.A0(new_n25688_), .A1(new_n9446_), .B0(pi0214), .Y(new_n26285_));
  AND2X1   g23849(.A(new_n25696_), .B(new_n23173_), .Y(new_n26286_));
  NOR3X1   g23850(.A(new_n26286_), .B(new_n25688_), .C(new_n24823_), .Y(new_n26287_));
  AOI21X1  g23851(.A0(new_n26287_), .A1(new_n26285_), .B0(new_n26284_), .Y(new_n26288_));
  AND2X1   g23852(.A(new_n25842_), .B(new_n25691_), .Y(new_n26289_));
  AOI21X1  g23853(.A0(new_n26289_), .A1(new_n2933_), .B0(new_n26288_), .Y(new_n26290_));
  NAND2X1  g23854(.A(new_n26290_), .B(new_n26264_), .Y(new_n26291_));
  OAI21X1  g23855(.A0(new_n26290_), .A1(new_n25722_), .B0(new_n25868_), .Y(new_n26292_));
  MX2X1    g23856(.A(new_n26292_), .B(new_n26291_), .S0(new_n25153_), .Y(new_n26293_));
  AOI21X1  g23857(.A0(new_n26293_), .A1(new_n26281_), .B0(new_n26280_), .Y(new_n26294_));
  OAI21X1  g23858(.A0(new_n26279_), .A1(new_n26263_), .B0(new_n26294_), .Y(new_n26295_));
  AOI21X1  g23859(.A0(new_n26295_), .A1(new_n26261_), .B0(pi1149), .Y(new_n26296_));
  OR4X1    g23860(.A(new_n25733_), .B(new_n25732_), .C(new_n25686_), .D(new_n24823_), .Y(new_n26297_));
  AOI21X1  g23861(.A0(new_n25728_), .A1(new_n25674_), .B0(new_n26297_), .Y(new_n26298_));
  OAI21X1  g23862(.A0(new_n26298_), .A1(new_n25854_), .B0(new_n8422_), .Y(new_n26299_));
  AND3X1   g23863(.A(new_n26299_), .B(new_n25856_), .C(pi1152), .Y(new_n26300_));
  NOR2X1   g23864(.A(new_n26008_), .B(new_n25694_), .Y(new_n26301_));
  OAI21X1  g23865(.A0(new_n25834_), .A1(pi0214), .B0(new_n25830_), .Y(new_n26302_));
  OAI21X1  g23866(.A0(new_n25834_), .A1(new_n25682_), .B0(new_n24823_), .Y(new_n26303_));
  AOI21X1  g23867(.A0(new_n26303_), .A1(new_n26302_), .B0(pi0219), .Y(new_n26304_));
  NAND2X1  g23868(.A(new_n25837_), .B(new_n25153_), .Y(new_n26305_));
  OAI21X1  g23869(.A0(new_n26305_), .A1(new_n26304_), .B0(new_n26301_), .Y(new_n26306_));
  AOI21X1  g23870(.A0(new_n26265_), .A1(new_n26055_), .B0(new_n26289_), .Y(new_n26307_));
  NAND2X1  g23871(.A(new_n26307_), .B(new_n25153_), .Y(new_n26308_));
  OR3X1    g23872(.A(new_n26264_), .B(new_n26054_), .C(new_n25868_), .Y(new_n26309_));
  AOI21X1  g23873(.A0(new_n25842_), .A1(new_n25867_), .B0(new_n25153_), .Y(new_n26310_));
  NOR2X1   g23874(.A(new_n25819_), .B(pi1151), .Y(new_n26311_));
  INVX1    g23875(.A(new_n26311_), .Y(new_n26312_));
  AOI21X1  g23876(.A0(new_n26310_), .A1(new_n26309_), .B0(new_n26312_), .Y(new_n26313_));
  AOI21X1  g23877(.A0(new_n26313_), .A1(new_n26308_), .B0(pi1150), .Y(new_n26314_));
  OAI21X1  g23878(.A0(new_n26306_), .A1(new_n26300_), .B0(new_n26314_), .Y(new_n26315_));
  NAND2X1  g23879(.A(new_n25728_), .B(pi0212), .Y(new_n26316_));
  AOI21X1  g23880(.A0(new_n26316_), .A1(new_n26267_), .B0(new_n25153_), .Y(new_n26317_));
  NOR2X1   g23881(.A(new_n25958_), .B(new_n25694_), .Y(new_n26318_));
  NOR2X1   g23882(.A(new_n26273_), .B(new_n25682_), .Y(new_n26319_));
  NOR2X1   g23883(.A(new_n26319_), .B(pi0219), .Y(new_n26320_));
  OAI21X1  g23884(.A0(new_n26320_), .A1(new_n26305_), .B0(new_n26318_), .Y(new_n26321_));
  AOI21X1  g23885(.A0(new_n26317_), .A1(new_n25856_), .B0(new_n26321_), .Y(new_n26322_));
  NOR2X1   g23886(.A(new_n26000_), .B(pi1151), .Y(new_n26323_));
  INVX1    g23887(.A(new_n26323_), .Y(new_n26324_));
  AOI21X1  g23888(.A0(new_n26290_), .A1(new_n26264_), .B0(pi1152), .Y(new_n26325_));
  INVX1    g23889(.A(new_n26307_), .Y(new_n26326_));
  NOR2X1   g23890(.A(new_n25713_), .B(new_n24877_), .Y(new_n26327_));
  NOR2X1   g23891(.A(new_n25686_), .B(new_n9446_), .Y(new_n26328_));
  OR2X1    g23892(.A(new_n26328_), .B(new_n25697_), .Y(new_n26329_));
  NOR2X1   g23893(.A(new_n25722_), .B(new_n7996_), .Y(new_n26330_));
  AOI21X1  g23894(.A0(new_n26330_), .A1(new_n26329_), .B0(new_n26327_), .Y(new_n26331_));
  OAI21X1  g23895(.A0(new_n26331_), .A1(pi0219), .B0(new_n26309_), .Y(new_n26332_));
  AOI22X1  g23896(.A0(new_n26332_), .A1(pi1152), .B0(new_n26326_), .B1(new_n26325_), .Y(new_n26333_));
  OAI21X1  g23897(.A0(new_n26333_), .A1(new_n26324_), .B0(pi1150), .Y(new_n26334_));
  OR2X1    g23898(.A(new_n26334_), .B(new_n26322_), .Y(new_n26335_));
  AOI21X1  g23899(.A0(new_n26335_), .A1(new_n26315_), .B0(new_n25955_), .Y(new_n26336_));
  OAI21X1  g23900(.A0(new_n26336_), .A1(new_n26296_), .B0(new_n24815_), .Y(new_n26337_));
  AOI21X1  g23901(.A0(new_n25876_), .A1(pi0213), .B0(new_n24866_), .Y(new_n26338_));
  OAI21X1  g23902(.A0(new_n25990_), .A1(new_n25987_), .B0(new_n26281_), .Y(new_n26339_));
  OAI21X1  g23903(.A0(new_n25953_), .A1(new_n25941_), .B0(new_n26262_), .Y(new_n26340_));
  AND3X1   g23904(.A(new_n26340_), .B(new_n26339_), .C(pi1150), .Y(new_n26341_));
  NOR3X1   g23905(.A(new_n26028_), .B(new_n25694_), .C(pi1150), .Y(new_n26342_));
  OR3X1    g23906(.A(new_n26342_), .B(new_n26341_), .C(pi1149), .Y(new_n26343_));
  AND2X1   g23907(.A(new_n26301_), .B(new_n26024_), .Y(new_n26344_));
  OAI21X1  g23908(.A0(new_n26312_), .A1(new_n26057_), .B0(new_n26280_), .Y(new_n26345_));
  NOR4X1   g23909(.A(new_n25963_), .B(new_n25961_), .C(new_n25958_), .D(new_n25694_), .Y(new_n26346_));
  INVX1    g23910(.A(new_n26346_), .Y(new_n26347_));
  AOI21X1  g23911(.A0(new_n26002_), .A1(new_n25694_), .B0(new_n26280_), .Y(new_n26348_));
  AOI21X1  g23912(.A0(new_n26348_), .A1(new_n26347_), .B0(new_n25955_), .Y(new_n26349_));
  OAI21X1  g23913(.A0(new_n26345_), .A1(new_n26344_), .B0(new_n26349_), .Y(new_n26350_));
  NAND3X1  g23914(.A(new_n26350_), .B(new_n26343_), .C(new_n24815_), .Y(new_n26351_));
  INVX1    g23915(.A(new_n25001_), .Y(new_n26352_));
  NAND3X1  g23916(.A(new_n25672_), .B(new_n26352_), .C(new_n23173_), .Y(new_n26353_));
  OAI21X1  g23917(.A0(new_n25655_), .A1(new_n23173_), .B0(new_n26353_), .Y(new_n26354_));
  OAI22X1  g23918(.A0(new_n26354_), .A1(new_n26012_), .B0(new_n26017_), .B1(new_n26013_), .Y(new_n26355_));
  AOI21X1  g23919(.A0(new_n26355_), .A1(new_n8422_), .B0(new_n26023_), .Y(new_n26356_));
  AND2X1   g23920(.A(new_n25652_), .B(pi0299), .Y(new_n26357_));
  OAI21X1  g23921(.A0(new_n26255_), .A1(new_n26033_), .B0(new_n6489_), .Y(new_n26358_));
  OAI21X1  g23922(.A0(new_n26358_), .A1(new_n26357_), .B0(new_n25797_), .Y(new_n26359_));
  AND2X1   g23923(.A(new_n26359_), .B(new_n25153_), .Y(new_n26360_));
  OAI21X1  g23924(.A0(new_n26356_), .A1(new_n25782_), .B0(new_n26360_), .Y(new_n26361_));
  INVX1    g23925(.A(new_n25821_), .Y(new_n26362_));
  AOI22X1  g23926(.A0(new_n26011_), .A1(new_n26010_), .B0(new_n25655_), .B1(new_n24849_), .Y(new_n26363_));
  NOR4X1   g23927(.A(new_n26363_), .B(new_n26142_), .C(new_n25683_), .D(pi0219), .Y(new_n26364_));
  OAI21X1  g23928(.A0(new_n26364_), .A1(new_n26023_), .B0(new_n26362_), .Y(new_n26365_));
  INVX1    g23929(.A(new_n24904_), .Y(new_n26366_));
  INVX1    g23930(.A(new_n26033_), .Y(new_n26367_));
  AOI22X1  g23931(.A0(new_n26367_), .A1(new_n25960_), .B0(new_n25805_), .B1(new_n26366_), .Y(new_n26368_));
  AOI21X1  g23932(.A0(new_n26367_), .A1(pi0219), .B0(po1038), .Y(new_n26369_));
  OAI21X1  g23933(.A0(new_n26368_), .A1(pi0219), .B0(new_n26369_), .Y(new_n26370_));
  AOI21X1  g23934(.A0(new_n26370_), .A1(new_n25807_), .B0(new_n25153_), .Y(new_n26371_));
  AOI21X1  g23935(.A0(new_n26371_), .A1(new_n26365_), .B0(pi1150), .Y(new_n26372_));
  NOR4X1   g23936(.A(new_n26142_), .B(new_n25962_), .C(pi1153), .D(pi0219), .Y(new_n26373_));
  AOI21X1  g23937(.A0(new_n7962_), .A1(pi0299), .B0(pi0219), .Y(new_n26374_));
  INVX1    g23938(.A(new_n26374_), .Y(new_n26375_));
  AOI21X1  g23939(.A0(new_n26375_), .A1(new_n26054_), .B0(new_n26145_), .Y(new_n26376_));
  NOR2X1   g23940(.A(new_n26376_), .B(new_n26373_), .Y(new_n26377_));
  AND3X1   g23941(.A(new_n26006_), .B(new_n24884_), .C(pi1153), .Y(new_n26378_));
  INVX1    g23942(.A(new_n26378_), .Y(new_n26379_));
  AOI21X1  g23943(.A0(new_n26379_), .A1(new_n25797_), .B0(pi1152), .Y(new_n26380_));
  NOR2X1   g23944(.A(new_n25998_), .B(pi1151), .Y(new_n26381_));
  NOR2X1   g23945(.A(new_n26381_), .B(pi1152), .Y(new_n26382_));
  OAI22X1  g23946(.A0(new_n26382_), .A1(new_n26380_), .B0(new_n26377_), .B1(new_n25782_), .Y(new_n26383_));
  OR2X1    g23947(.A(new_n25963_), .B(new_n25961_), .Y(new_n26384_));
  OR4X1    g23948(.A(new_n26142_), .B(new_n25962_), .C(pi0219), .D(pi0211), .Y(new_n26385_));
  AND2X1   g23949(.A(new_n26385_), .B(new_n26384_), .Y(new_n26386_));
  NOR3X1   g23950(.A(new_n26386_), .B(new_n26377_), .C(new_n25821_), .Y(new_n26387_));
  AND2X1   g23951(.A(new_n25741_), .B(new_n6489_), .Y(new_n26388_));
  OR2X1    g23952(.A(new_n26038_), .B(new_n24877_), .Y(new_n26389_));
  NOR3X1   g23953(.A(new_n25733_), .B(new_n25732_), .C(pi0299), .Y(new_n26390_));
  OR3X1    g23954(.A(new_n26390_), .B(new_n26357_), .C(new_n24824_), .Y(new_n26391_));
  NAND3X1  g23955(.A(new_n26391_), .B(new_n26389_), .C(new_n26081_), .Y(new_n26392_));
  AOI21X1  g23956(.A0(new_n26392_), .A1(new_n26388_), .B0(new_n25808_), .Y(new_n26393_));
  OR3X1    g23957(.A(new_n26393_), .B(new_n26387_), .C(new_n25153_), .Y(new_n26394_));
  AND3X1   g23958(.A(new_n26394_), .B(new_n26383_), .C(pi1150), .Y(new_n26395_));
  OR2X1    g23959(.A(new_n26395_), .B(new_n25955_), .Y(new_n26396_));
  AOI21X1  g23960(.A0(new_n26372_), .A1(new_n26361_), .B0(new_n26396_), .Y(new_n26397_));
  NOR3X1   g23961(.A(new_n26357_), .B(new_n25978_), .C(new_n24849_), .Y(new_n26398_));
  NOR3X1   g23962(.A(new_n26357_), .B(new_n25978_), .C(pi0214), .Y(new_n26399_));
  OAI22X1  g23963(.A0(new_n26399_), .A1(new_n25981_), .B0(new_n26398_), .B1(new_n25977_), .Y(new_n26400_));
  AOI21X1  g23964(.A0(new_n26400_), .A1(new_n8422_), .B0(new_n25990_), .Y(new_n26401_));
  INVX1    g23965(.A(new_n26123_), .Y(new_n26402_));
  NOR2X1   g23966(.A(new_n25943_), .B(new_n23173_), .Y(new_n26403_));
  OAI21X1  g23967(.A0(new_n24986_), .A1(new_n24950_), .B0(new_n25706_), .Y(new_n26404_));
  AND3X1   g23968(.A(new_n26404_), .B(new_n26352_), .C(new_n23173_), .Y(new_n26405_));
  NOR2X1   g23969(.A(new_n26405_), .B(new_n26403_), .Y(new_n26406_));
  AOI21X1  g23970(.A0(new_n26406_), .A1(pi0214), .B0(new_n25946_), .Y(new_n26407_));
  AOI21X1  g23971(.A0(new_n26406_), .A1(new_n24849_), .B0(new_n26128_), .Y(new_n26408_));
  NOR3X1   g23972(.A(new_n26408_), .B(new_n26407_), .C(pi0219), .Y(new_n26409_));
  OAI21X1  g23973(.A0(new_n26409_), .A1(new_n26402_), .B0(new_n26362_), .Y(new_n26410_));
  AND2X1   g23974(.A(new_n26410_), .B(pi1152), .Y(new_n26411_));
  OAI21X1  g23975(.A0(new_n26401_), .A1(new_n25808_), .B0(new_n26411_), .Y(new_n26412_));
  OAI21X1  g23976(.A0(new_n25978_), .A1(new_n25001_), .B0(new_n23173_), .Y(new_n26413_));
  NOR2X1   g23977(.A(new_n25980_), .B(new_n25799_), .Y(new_n26414_));
  AOI22X1  g23978(.A0(new_n26414_), .A1(new_n26413_), .B0(new_n25971_), .B1(new_n25799_), .Y(new_n26415_));
  OAI21X1  g23979(.A0(new_n26415_), .A1(po1038), .B0(new_n25797_), .Y(new_n26416_));
  INVX1    g23980(.A(new_n25782_), .Y(new_n26417_));
  NOR3X1   g23981(.A(new_n26403_), .B(new_n25720_), .C(new_n24849_), .Y(new_n26418_));
  OAI21X1  g23982(.A0(new_n25949_), .A1(new_n25945_), .B0(pi0212), .Y(new_n26419_));
  NOR3X1   g23983(.A(new_n26419_), .B(new_n26418_), .C(new_n26406_), .Y(new_n26420_));
  NOR2X1   g23984(.A(new_n26405_), .B(new_n25950_), .Y(new_n26421_));
  OAI21X1  g23985(.A0(new_n26421_), .A1(new_n25946_), .B0(new_n8422_), .Y(new_n26422_));
  OAI21X1  g23986(.A0(new_n26422_), .A1(new_n26420_), .B0(new_n26123_), .Y(new_n26423_));
  AOI21X1  g23987(.A0(new_n26423_), .A1(new_n26417_), .B0(pi1152), .Y(new_n26424_));
  AOI21X1  g23988(.A0(new_n26424_), .A1(new_n26416_), .B0(new_n26280_), .Y(new_n26425_));
  NOR3X1   g23989(.A(new_n25697_), .B(new_n25688_), .C(new_n9446_), .Y(new_n26426_));
  OR2X1    g23990(.A(new_n26426_), .B(new_n8422_), .Y(new_n26427_));
  AND2X1   g23991(.A(new_n26427_), .B(new_n6489_), .Y(new_n26428_));
  NAND2X1  g23992(.A(new_n26428_), .B(new_n25845_), .Y(new_n26429_));
  OAI21X1  g23993(.A0(new_n26287_), .A1(new_n26284_), .B0(new_n26428_), .Y(new_n26430_));
  NAND3X1  g23994(.A(new_n26430_), .B(new_n26429_), .C(new_n26362_), .Y(new_n26431_));
  NOR3X1   g23995(.A(new_n24816_), .B(new_n7962_), .C(pi0219), .Y(new_n26432_));
  INVX1    g23996(.A(new_n26432_), .Y(new_n26433_));
  OR3X1    g23997(.A(new_n25805_), .B(new_n26433_), .C(new_n2933_), .Y(new_n26434_));
  AOI21X1  g23998(.A0(new_n26434_), .A1(new_n25807_), .B0(new_n25153_), .Y(new_n26435_));
  INVX1    g23999(.A(new_n26380_), .Y(new_n26436_));
  AOI21X1  g24000(.A0(new_n26428_), .A1(new_n25845_), .B0(new_n25782_), .Y(new_n26437_));
  OAI21X1  g24001(.A0(new_n26437_), .A1(new_n26436_), .B0(new_n26280_), .Y(new_n26438_));
  AOI21X1  g24002(.A0(new_n26435_), .A1(new_n26431_), .B0(new_n26438_), .Y(new_n26439_));
  OR2X1    g24003(.A(new_n26439_), .B(pi1149), .Y(new_n26440_));
  AOI21X1  g24004(.A0(new_n26425_), .A1(new_n26412_), .B0(new_n26440_), .Y(new_n26441_));
  OAI21X1  g24005(.A0(new_n26441_), .A1(new_n26397_), .B0(pi0213), .Y(new_n26442_));
  AND3X1   g24006(.A(new_n26442_), .B(new_n26351_), .C(new_n24866_), .Y(new_n26443_));
  AOI21X1  g24007(.A0(new_n26338_), .A1(new_n26337_), .B0(new_n26443_), .Y(new_n26444_));
  MX2X1    g24008(.A(new_n26444_), .B(pi0241), .S0(new_n24814_), .Y(po0398));
  MX2X1    g24009(.A(new_n26064_), .B(new_n25508_), .S0(pi0214), .Y(new_n26446_));
  NOR3X1   g24010(.A(new_n26063_), .B(new_n24849_), .C(pi0212), .Y(new_n26447_));
  OR2X1    g24011(.A(new_n26447_), .B(pi0219), .Y(new_n26448_));
  AOI21X1  g24012(.A0(new_n26446_), .A1(pi0212), .B0(new_n26448_), .Y(new_n26449_));
  AOI21X1  g24013(.A0(pi1144), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n26450_));
  NOR3X1   g24014(.A(new_n26450_), .B(new_n26449_), .C(new_n25651_), .Y(new_n26451_));
  INVX1    g24015(.A(new_n26451_), .Y(new_n26452_));
  AOI21X1  g24016(.A0(pi1144), .A1(pi0199), .B0(pi0200), .Y(new_n26453_));
  OAI21X1  g24017(.A0(new_n3140_), .A1(pi0199), .B0(new_n26453_), .Y(new_n26454_));
  AND3X1   g24018(.A(new_n26454_), .B(new_n26159_), .C(new_n2933_), .Y(new_n26455_));
  OAI21X1  g24019(.A0(new_n3309_), .A1(pi0199), .B0(new_n26453_), .Y(new_n26456_));
  NAND3X1  g24020(.A(new_n26456_), .B(new_n25498_), .C(new_n2933_), .Y(new_n26457_));
  AOI21X1  g24021(.A0(new_n26457_), .A1(pi0207), .B0(new_n22959_), .Y(new_n26458_));
  OAI21X1  g24022(.A0(new_n26455_), .A1(pi0207), .B0(new_n26458_), .Y(new_n26459_));
  NAND4X1  g24023(.A(new_n26454_), .B(new_n26159_), .C(new_n24844_), .D(new_n2933_), .Y(new_n26460_));
  AND3X1   g24024(.A(new_n26460_), .B(new_n26459_), .C(new_n25606_), .Y(new_n26461_));
  NOR2X1   g24025(.A(new_n26461_), .B(pi0211), .Y(new_n26462_));
  AND3X1   g24026(.A(new_n26460_), .B(new_n26459_), .C(new_n25073_), .Y(new_n26463_));
  OAI21X1  g24027(.A0(new_n26463_), .A1(new_n23173_), .B0(pi0214), .Y(new_n26464_));
  INVX1    g24028(.A(new_n26106_), .Y(new_n26465_));
  AND3X1   g24029(.A(new_n26460_), .B(new_n26459_), .C(new_n26465_), .Y(new_n26466_));
  MX2X1    g24030(.A(new_n26466_), .B(new_n26461_), .S0(pi0211), .Y(new_n26467_));
  AOI21X1  g24031(.A0(new_n26467_), .A1(new_n24849_), .B0(new_n24823_), .Y(new_n26468_));
  OAI21X1  g24032(.A0(new_n26464_), .A1(new_n26462_), .B0(new_n26468_), .Y(new_n26469_));
  NAND4X1  g24033(.A(new_n26454_), .B(new_n26159_), .C(new_n25115_), .D(new_n2933_), .Y(new_n26470_));
  AND3X1   g24034(.A(new_n26470_), .B(new_n26459_), .C(new_n24849_), .Y(new_n26471_));
  NOR2X1   g24035(.A(new_n26471_), .B(pi0212), .Y(new_n26472_));
  NAND2X1  g24036(.A(new_n26467_), .B(pi0214), .Y(new_n26473_));
  AOI21X1  g24037(.A0(new_n26473_), .A1(new_n26472_), .B0(pi0219), .Y(new_n26474_));
  AND2X1   g24038(.A(new_n26474_), .B(new_n26469_), .Y(new_n26475_));
  AND2X1   g24039(.A(new_n26470_), .B(new_n26459_), .Y(new_n26476_));
  INVX1    g24040(.A(new_n26476_), .Y(new_n26477_));
  AOI21X1  g24041(.A0(new_n26477_), .A1(new_n25162_), .B0(new_n8422_), .Y(new_n26478_));
  OAI21X1  g24042(.A0(new_n26463_), .A1(new_n25162_), .B0(new_n26478_), .Y(new_n26479_));
  NAND2X1  g24043(.A(new_n26479_), .B(new_n6489_), .Y(new_n26480_));
  OAI21X1  g24044(.A0(new_n26480_), .A1(new_n26475_), .B0(new_n26452_), .Y(new_n26481_));
  AOI21X1  g24045(.A0(pi1142), .A1(pi0299), .B0(new_n25162_), .Y(new_n26482_));
  AOI22X1  g24046(.A0(new_n26482_), .A1(new_n26460_), .B0(new_n26470_), .B1(pi0211), .Y(new_n26483_));
  OAI22X1  g24047(.A0(new_n25086_), .A1(new_n24831_), .B0(new_n24851_), .B1(new_n24877_), .Y(new_n26484_));
  AND2X1   g24048(.A(new_n26460_), .B(new_n8422_), .Y(new_n26485_));
  AOI22X1  g24049(.A0(new_n26485_), .A1(new_n26484_), .B0(new_n26470_), .B1(new_n24816_), .Y(new_n26486_));
  OAI21X1  g24050(.A0(new_n26483_), .A1(new_n8422_), .B0(new_n26486_), .Y(new_n26487_));
  AOI21X1  g24051(.A0(new_n26487_), .A1(new_n26459_), .B0(po1038), .Y(new_n26488_));
  OR2X1    g24052(.A(new_n24829_), .B(pi0213), .Y(new_n26489_));
  OAI22X1  g24053(.A0(new_n26489_), .A1(new_n26488_), .B0(new_n26481_), .B1(new_n24815_), .Y(new_n26490_));
  AND2X1   g24054(.A(new_n24816_), .B(pi0219), .Y(new_n26491_));
  OR3X1    g24055(.A(new_n26491_), .B(new_n26450_), .C(new_n26449_), .Y(new_n26492_));
  AOI21X1  g24056(.A0(new_n26492_), .A1(pi0299), .B0(po1038), .Y(new_n26493_));
  AOI21X1  g24057(.A0(new_n26493_), .A1(new_n24859_), .B0(new_n26451_), .Y(new_n26494_));
  OAI21X1  g24058(.A0(new_n26494_), .A1(new_n24815_), .B0(new_n24866_), .Y(new_n26495_));
  AOI21X1  g24059(.A0(new_n24865_), .A1(new_n24815_), .B0(new_n26495_), .Y(new_n26496_));
  AOI21X1  g24060(.A0(new_n26490_), .A1(pi0209), .B0(new_n26496_), .Y(new_n26497_));
  MX2X1    g24061(.A(new_n26497_), .B(pi0242), .S0(new_n24814_), .Y(po0399));
  INVX1    g24062(.A(pi0243), .Y(new_n26499_));
  INVX1    g24063(.A(pi0271), .Y(new_n26500_));
  AOI21X1  g24064(.A0(new_n5124_), .A1(new_n2594_), .B0(new_n5117_), .Y(new_n26501_));
  AND3X1   g24065(.A(new_n26501_), .B(pi0802), .C(pi0276), .Y(new_n26502_));
  NOR2X1   g24066(.A(new_n26502_), .B(pi1091), .Y(new_n26503_));
  NOR2X1   g24067(.A(new_n26503_), .B(new_n26500_), .Y(new_n26504_));
  AOI21X1  g24068(.A0(new_n26504_), .A1(pi0273), .B0(pi1091), .Y(new_n26505_));
  OR2X1    g24069(.A(new_n26505_), .B(pi0200), .Y(new_n26506_));
  OR2X1    g24070(.A(new_n26505_), .B(new_n7871_), .Y(new_n26507_));
  OR3X1    g24071(.A(pi0085), .B(pi0083), .C(pi0081), .Y(new_n26508_));
  NAND4X1  g24072(.A(new_n26508_), .B(pi0802), .C(pi0314), .D(pi0276), .Y(new_n26509_));
  NOR2X1   g24073(.A(new_n26509_), .B(pi1091), .Y(new_n26510_));
  INVX1    g24074(.A(new_n26510_), .Y(new_n26511_));
  OAI21X1  g24075(.A0(new_n26504_), .A1(pi1091), .B0(pi0273), .Y(new_n26512_));
  INVX1    g24076(.A(pi0273), .Y(new_n26513_));
  NOR4X1   g24077(.A(new_n26509_), .B(pi1091), .C(new_n26513_), .D(new_n26500_), .Y(new_n26514_));
  INVX1    g24078(.A(new_n26514_), .Y(new_n26515_));
  AND2X1   g24079(.A(new_n26515_), .B(new_n26512_), .Y(new_n26516_));
  AOI21X1  g24080(.A0(new_n26516_), .A1(new_n2702_), .B0(pi0199), .Y(new_n26517_));
  INVX1    g24081(.A(new_n26517_), .Y(new_n26518_));
  AOI21X1  g24082(.A0(new_n26518_), .A1(new_n26507_), .B0(new_n26511_), .Y(new_n26519_));
  NOR2X1   g24083(.A(new_n26519_), .B(pi0299), .Y(new_n26520_));
  AND3X1   g24084(.A(new_n26520_), .B(new_n26507_), .C(new_n26506_), .Y(new_n26521_));
  NOR2X1   g24085(.A(new_n26514_), .B(new_n2933_), .Y(new_n26522_));
  OAI22X1  g24086(.A0(new_n26522_), .A1(new_n26521_), .B0(pi1091), .B1(new_n26499_), .Y(new_n26523_));
  NOR2X1   g24087(.A(new_n26510_), .B(pi0200), .Y(new_n26524_));
  AOI21X1  g24088(.A0(new_n26518_), .A1(new_n26507_), .B0(new_n26524_), .Y(new_n26525_));
  NOR2X1   g24089(.A(new_n26525_), .B(pi0299), .Y(new_n26526_));
  AND2X1   g24090(.A(new_n26526_), .B(new_n26507_), .Y(new_n26527_));
  AND3X1   g24091(.A(new_n26502_), .B(new_n2702_), .C(pi0271), .Y(new_n26528_));
  AOI21X1  g24092(.A0(new_n26528_), .A1(pi0273), .B0(new_n2933_), .Y(new_n26529_));
  AND3X1   g24093(.A(new_n26520_), .B(new_n26518_), .C(new_n26506_), .Y(new_n26530_));
  NOR3X1   g24094(.A(new_n26530_), .B(new_n26529_), .C(new_n26527_), .Y(new_n26531_));
  INVX1    g24095(.A(new_n26531_), .Y(new_n26532_));
  AND2X1   g24096(.A(new_n26520_), .B(new_n26506_), .Y(new_n26533_));
  INVX1    g24097(.A(new_n26533_), .Y(new_n26534_));
  AND2X1   g24098(.A(new_n26505_), .B(pi0299), .Y(new_n26535_));
  INVX1    g24099(.A(new_n26535_), .Y(new_n26536_));
  AOI21X1  g24100(.A0(new_n26536_), .A1(new_n26534_), .B0(new_n26499_), .Y(new_n26537_));
  AOI21X1  g24101(.A0(new_n26537_), .A1(new_n26532_), .B0(new_n12463_), .Y(new_n26538_));
  AND3X1   g24102(.A(new_n26515_), .B(new_n26505_), .C(pi0299), .Y(new_n26539_));
  NOR3X1   g24103(.A(new_n26539_), .B(new_n26530_), .C(new_n12463_), .Y(new_n26540_));
  MX2X1    g24104(.A(new_n26525_), .B(new_n26514_), .S0(pi0299), .Y(new_n26541_));
  NAND2X1  g24105(.A(new_n26541_), .B(new_n26499_), .Y(new_n26542_));
  OAI22X1  g24106(.A0(new_n26542_), .A1(new_n26521_), .B0(new_n26540_), .B1(new_n26538_), .Y(new_n26543_));
  NOR3X1   g24107(.A(new_n26525_), .B(new_n26517_), .C(pi0299), .Y(new_n26544_));
  OR3X1    g24108(.A(new_n26544_), .B(new_n26539_), .C(new_n26521_), .Y(new_n26545_));
  NOR4X1   g24109(.A(new_n26530_), .B(new_n26527_), .C(new_n26522_), .D(new_n26499_), .Y(new_n26546_));
  AOI21X1  g24110(.A0(new_n26545_), .A1(new_n26499_), .B0(new_n26546_), .Y(new_n26547_));
  OR2X1    g24111(.A(new_n26547_), .B(pi1155), .Y(new_n26548_));
  NAND3X1  g24112(.A(new_n26548_), .B(new_n26543_), .C(new_n26523_), .Y(new_n26549_));
  AND2X1   g24113(.A(new_n26549_), .B(pi1156), .Y(new_n26550_));
  NOR2X1   g24114(.A(new_n26544_), .B(new_n26535_), .Y(new_n26551_));
  NOR2X1   g24115(.A(new_n26551_), .B(pi0243), .Y(new_n26552_));
  INVX1    g24116(.A(new_n26522_), .Y(new_n26553_));
  OAI21X1  g24117(.A0(new_n26519_), .A1(pi0299), .B0(new_n26553_), .Y(new_n26554_));
  AOI21X1  g24118(.A0(new_n26554_), .A1(new_n26552_), .B0(pi1155), .Y(new_n26555_));
  AND2X1   g24119(.A(new_n26520_), .B(new_n26507_), .Y(new_n26556_));
  NOR4X1   g24120(.A(new_n26533_), .B(new_n26522_), .C(new_n26556_), .D(new_n26499_), .Y(new_n26557_));
  INVX1    g24121(.A(new_n26557_), .Y(new_n26558_));
  AOI21X1  g24122(.A0(new_n26558_), .A1(new_n26555_), .B0(pi1156), .Y(new_n26559_));
  INVX1    g24123(.A(new_n26559_), .Y(new_n26560_));
  AOI21X1  g24124(.A0(new_n26520_), .A1(new_n26506_), .B0(new_n26522_), .Y(new_n26561_));
  NOR2X1   g24125(.A(new_n26539_), .B(new_n26526_), .Y(new_n26562_));
  OAI21X1  g24126(.A0(new_n26562_), .A1(pi0243), .B0(pi1155), .Y(new_n26563_));
  AOI21X1  g24127(.A0(new_n26561_), .A1(pi0243), .B0(new_n26563_), .Y(new_n26564_));
  OAI21X1  g24128(.A0(new_n26564_), .A1(new_n26560_), .B0(pi1157), .Y(new_n26565_));
  NOR2X1   g24129(.A(new_n26554_), .B(pi1155), .Y(new_n26566_));
  NOR2X1   g24130(.A(pi1091), .B(pi0243), .Y(new_n26567_));
  AND2X1   g24131(.A(new_n26528_), .B(pi0273), .Y(new_n26568_));
  MX2X1    g24132(.A(new_n26568_), .B(new_n26519_), .S0(new_n2933_), .Y(new_n26569_));
  INVX1    g24133(.A(new_n26569_), .Y(new_n26570_));
  AOI21X1  g24134(.A0(new_n26570_), .A1(new_n26567_), .B0(pi1155), .Y(new_n26571_));
  OAI22X1  g24135(.A0(new_n26571_), .A1(new_n26566_), .B0(new_n26554_), .B1(new_n26499_), .Y(new_n26572_));
  AND2X1   g24136(.A(new_n26572_), .B(new_n12555_), .Y(new_n26573_));
  AND2X1   g24137(.A(new_n2702_), .B(pi0243), .Y(new_n26574_));
  NOR4X1   g24138(.A(new_n26505_), .B(new_n26574_), .C(new_n12463_), .D(new_n7871_), .Y(new_n26575_));
  NOR2X1   g24139(.A(new_n26575_), .B(new_n26564_), .Y(new_n26576_));
  NAND2X1  g24140(.A(new_n26576_), .B(new_n26573_), .Y(new_n26577_));
  AND3X1   g24141(.A(new_n26561_), .B(new_n26511_), .C(new_n12463_), .Y(new_n26578_));
  NOR3X1   g24142(.A(new_n26519_), .B(new_n26517_), .C(pi0299), .Y(new_n26579_));
  NOR2X1   g24143(.A(new_n26579_), .B(new_n26539_), .Y(new_n26580_));
  INVX1    g24144(.A(new_n26580_), .Y(new_n26581_));
  AOI21X1  g24145(.A0(new_n26520_), .A1(new_n26507_), .B0(new_n26522_), .Y(new_n26582_));
  MX2X1    g24146(.A(new_n26582_), .B(new_n26581_), .S0(pi0243), .Y(new_n26583_));
  NOR3X1   g24147(.A(new_n26583_), .B(new_n26578_), .C(new_n12555_), .Y(new_n26584_));
  NOR2X1   g24148(.A(new_n26584_), .B(pi1157), .Y(new_n26585_));
  AOI21X1  g24149(.A0(new_n26585_), .A1(new_n26577_), .B0(new_n23173_), .Y(new_n26586_));
  OAI21X1  g24150(.A0(new_n26565_), .A1(new_n26550_), .B0(new_n26586_), .Y(new_n26587_));
  AOI21X1  g24151(.A0(new_n26548_), .A1(new_n26543_), .B0(new_n12555_), .Y(new_n26588_));
  AOI21X1  g24152(.A0(new_n26520_), .A1(new_n26506_), .B0(new_n26539_), .Y(new_n26589_));
  OAI21X1  g24153(.A0(new_n26589_), .A1(new_n26499_), .B0(new_n26542_), .Y(new_n26590_));
  OAI21X1  g24154(.A0(new_n26590_), .A1(new_n26560_), .B0(pi1157), .Y(new_n26591_));
  NOR4X1   g24155(.A(new_n26541_), .B(new_n26539_), .C(new_n26533_), .D(pi1155), .Y(new_n26592_));
  OR4X1    g24156(.A(new_n26592_), .B(new_n26583_), .C(new_n26578_), .D(new_n12555_), .Y(new_n26593_));
  OAI21X1  g24157(.A0(new_n26590_), .A1(new_n26583_), .B0(pi1155), .Y(new_n26594_));
  AOI21X1  g24158(.A0(new_n26594_), .A1(new_n26573_), .B0(pi1157), .Y(new_n26595_));
  AOI21X1  g24159(.A0(new_n26595_), .A1(new_n26593_), .B0(pi0211), .Y(new_n26596_));
  OAI21X1  g24160(.A0(new_n26591_), .A1(new_n26588_), .B0(new_n26596_), .Y(new_n26597_));
  AND2X1   g24161(.A(new_n26597_), .B(new_n8422_), .Y(new_n26598_));
  INVX1    g24162(.A(pi0263), .Y(new_n26599_));
  AND3X1   g24163(.A(pi0267), .B(pi0254), .C(pi0253), .Y(new_n26600_));
  AND2X1   g24164(.A(new_n26600_), .B(new_n26599_), .Y(new_n26601_));
  MX2X1    g24165(.A(new_n26568_), .B(new_n26525_), .S0(new_n2933_), .Y(new_n26602_));
  INVX1    g24166(.A(new_n26602_), .Y(new_n26603_));
  OR4X1    g24167(.A(new_n26603_), .B(new_n26535_), .C(new_n26521_), .D(pi0243), .Y(new_n26604_));
  NAND2X1  g24168(.A(new_n26604_), .B(new_n26538_), .Y(new_n26605_));
  NOR2X1   g24169(.A(new_n26535_), .B(new_n26521_), .Y(new_n26606_));
  INVX1    g24170(.A(new_n26606_), .Y(new_n26607_));
  MX2X1    g24171(.A(new_n26607_), .B(new_n26531_), .S0(pi0243), .Y(new_n26608_));
  OAI21X1  g24172(.A0(new_n26551_), .A1(pi0243), .B0(new_n26523_), .Y(new_n26609_));
  OAI21X1  g24173(.A0(new_n26609_), .A1(new_n26608_), .B0(new_n12463_), .Y(new_n26610_));
  AOI21X1  g24174(.A0(new_n26610_), .A1(new_n26605_), .B0(new_n12555_), .Y(new_n26611_));
  OR2X1    g24175(.A(new_n26544_), .B(new_n26529_), .Y(new_n26612_));
  OAI21X1  g24176(.A0(new_n26556_), .A1(new_n26499_), .B0(new_n12463_), .Y(new_n26613_));
  AOI21X1  g24177(.A0(new_n26612_), .A1(new_n26499_), .B0(new_n26613_), .Y(new_n26614_));
  AND3X1   g24178(.A(new_n26602_), .B(pi1155), .C(new_n26499_), .Y(new_n26615_));
  NOR4X1   g24179(.A(new_n26615_), .B(new_n26614_), .C(new_n26537_), .D(pi1156), .Y(new_n26616_));
  OR4X1    g24180(.A(new_n26616_), .B(new_n26611_), .C(new_n12578_), .D(pi0211), .Y(new_n26617_));
  INVX1    g24181(.A(new_n26608_), .Y(new_n26618_));
  NOR3X1   g24182(.A(new_n26530_), .B(new_n26529_), .C(new_n26499_), .Y(new_n26619_));
  OAI22X1  g24183(.A0(new_n26619_), .A1(new_n26563_), .B0(new_n26552_), .B1(pi1155), .Y(new_n26620_));
  AOI21X1  g24184(.A0(new_n26620_), .A1(new_n26618_), .B0(new_n12555_), .Y(new_n26621_));
  NOR2X1   g24185(.A(new_n26562_), .B(pi0243), .Y(new_n26622_));
  AOI21X1  g24186(.A0(new_n26520_), .A1(new_n26506_), .B0(new_n26529_), .Y(new_n26623_));
  AND2X1   g24187(.A(new_n26623_), .B(pi0243), .Y(new_n26624_));
  OAI21X1  g24188(.A0(new_n26624_), .A1(new_n26622_), .B0(pi1155), .Y(new_n26625_));
  NOR3X1   g24189(.A(new_n26533_), .B(new_n26529_), .C(new_n26556_), .Y(new_n26626_));
  AOI21X1  g24190(.A0(new_n26626_), .A1(pi0243), .B0(new_n26552_), .Y(new_n26627_));
  AOI21X1  g24191(.A0(new_n26627_), .A1(new_n26625_), .B0(pi1156), .Y(new_n26628_));
  OR4X1    g24192(.A(new_n26628_), .B(new_n26621_), .C(new_n12578_), .D(new_n23173_), .Y(new_n26629_));
  NOR3X1   g24193(.A(new_n26579_), .B(new_n26529_), .C(new_n12463_), .Y(new_n26630_));
  NOR3X1   g24194(.A(new_n26579_), .B(new_n26529_), .C(new_n26526_), .Y(new_n26631_));
  OAI21X1  g24195(.A0(new_n26631_), .A1(new_n26630_), .B0(pi0243), .Y(new_n26632_));
  AOI21X1  g24196(.A0(new_n26520_), .A1(new_n26507_), .B0(new_n26535_), .Y(new_n26633_));
  OR3X1    g24197(.A(new_n26633_), .B(new_n26578_), .C(pi0243), .Y(new_n26634_));
  AOI21X1  g24198(.A0(new_n26634_), .A1(new_n26632_), .B0(new_n12555_), .Y(new_n26635_));
  OR4X1    g24199(.A(new_n26579_), .B(new_n26533_), .C(new_n26529_), .D(new_n26499_), .Y(new_n26636_));
  OR2X1    g24200(.A(new_n26535_), .B(new_n26527_), .Y(new_n26637_));
  AOI21X1  g24201(.A0(new_n26637_), .A1(new_n26499_), .B0(new_n12463_), .Y(new_n26638_));
  OAI21X1  g24202(.A0(new_n26570_), .A1(new_n26499_), .B0(new_n26571_), .Y(new_n26639_));
  NAND2X1  g24203(.A(new_n26639_), .B(new_n12555_), .Y(new_n26640_));
  AOI21X1  g24204(.A0(new_n26638_), .A1(new_n26636_), .B0(new_n26640_), .Y(new_n26641_));
  OR3X1    g24205(.A(new_n26641_), .B(new_n26635_), .C(pi1157), .Y(new_n26642_));
  AND3X1   g24206(.A(new_n26642_), .B(new_n26629_), .C(new_n26617_), .Y(new_n26643_));
  OAI21X1  g24207(.A0(new_n26643_), .A1(new_n8422_), .B0(new_n26601_), .Y(new_n26644_));
  AOI21X1  g24208(.A0(new_n26598_), .A1(new_n26587_), .B0(new_n26644_), .Y(new_n26645_));
  AOI21X1  g24209(.A0(new_n25130_), .A1(new_n2933_), .B0(new_n12555_), .Y(new_n26646_));
  AND2X1   g24210(.A(pi1091), .B(new_n2933_), .Y(new_n26647_));
  AOI21X1  g24211(.A0(new_n26647_), .A1(new_n25131_), .B0(new_n26567_), .Y(new_n26648_));
  NOR2X1   g24212(.A(new_n26648_), .B(new_n12555_), .Y(new_n26649_));
  NOR2X1   g24213(.A(new_n25204_), .B(new_n2702_), .Y(new_n26650_));
  AOI21X1  g24214(.A0(new_n26650_), .A1(new_n26646_), .B0(new_n26649_), .Y(new_n26651_));
  AND3X1   g24215(.A(new_n2933_), .B(new_n7937_), .C(pi0199), .Y(new_n26652_));
  MX2X1    g24216(.A(new_n26652_), .B(new_n26499_), .S0(new_n2702_), .Y(new_n26653_));
  MX2X1    g24217(.A(pi1155), .B(new_n26499_), .S0(new_n2702_), .Y(new_n26654_));
  AND2X1   g24218(.A(new_n26654_), .B(new_n24916_), .Y(new_n26655_));
  OAI21X1  g24219(.A0(new_n26655_), .A1(new_n26653_), .B0(new_n12555_), .Y(new_n26656_));
  AOI21X1  g24220(.A0(new_n26656_), .A1(new_n26651_), .B0(new_n12578_), .Y(new_n26657_));
  OAI21X1  g24221(.A0(new_n25204_), .A1(new_n2702_), .B0(new_n26654_), .Y(new_n26658_));
  NAND2X1  g24222(.A(new_n26658_), .B(new_n12555_), .Y(new_n26659_));
  AND2X1   g24223(.A(pi1091), .B(pi0199), .Y(new_n26660_));
  AND2X1   g24224(.A(new_n26660_), .B(new_n2933_), .Y(new_n26661_));
  NOR3X1   g24225(.A(new_n26661_), .B(new_n26574_), .C(new_n12463_), .Y(new_n26662_));
  NOR2X1   g24226(.A(new_n26662_), .B(new_n12555_), .Y(new_n26663_));
  AOI21X1  g24227(.A0(new_n2702_), .A1(pi0243), .B0(pi1155), .Y(new_n26664_));
  OR3X1    g24228(.A(new_n25004_), .B(new_n2702_), .C(pi0299), .Y(new_n26665_));
  NAND2X1  g24229(.A(new_n26665_), .B(new_n26664_), .Y(new_n26666_));
  AOI21X1  g24230(.A0(new_n26666_), .A1(new_n26663_), .B0(pi1157), .Y(new_n26667_));
  AOI21X1  g24231(.A0(new_n26667_), .A1(new_n26659_), .B0(new_n26657_), .Y(new_n26668_));
  NAND2X1  g24232(.A(new_n26653_), .B(new_n12463_), .Y(new_n26669_));
  AND2X1   g24233(.A(pi1091), .B(pi0200), .Y(new_n26670_));
  AND2X1   g24234(.A(new_n26670_), .B(new_n2933_), .Y(new_n26671_));
  OR3X1    g24235(.A(new_n26671_), .B(new_n26574_), .C(new_n12463_), .Y(new_n26672_));
  AND2X1   g24236(.A(new_n26672_), .B(new_n12555_), .Y(new_n26673_));
  AOI22X1  g24237(.A0(new_n26673_), .A1(new_n26669_), .B0(new_n26663_), .B1(new_n26648_), .Y(new_n26674_));
  NOR2X1   g24238(.A(new_n26674_), .B(new_n12578_), .Y(new_n26675_));
  OR2X1    g24239(.A(new_n8467_), .B(new_n2702_), .Y(new_n26676_));
  AOI21X1  g24240(.A0(new_n26676_), .A1(new_n26664_), .B0(new_n26662_), .Y(new_n26677_));
  NOR4X1   g24241(.A(pi1156), .B(new_n2702_), .C(pi0299), .D(new_n7937_), .Y(new_n26678_));
  NOR2X1   g24242(.A(new_n26678_), .B(new_n26677_), .Y(new_n26679_));
  OAI21X1  g24243(.A0(new_n26679_), .A1(pi1157), .B0(new_n23173_), .Y(new_n26680_));
  OAI22X1  g24244(.A0(new_n26680_), .A1(new_n26675_), .B0(new_n26668_), .B1(new_n23173_), .Y(new_n26681_));
  NOR3X1   g24245(.A(new_n26649_), .B(new_n12578_), .C(new_n23173_), .Y(new_n26682_));
  AOI21X1  g24246(.A0(new_n26682_), .A1(new_n26656_), .B0(new_n8422_), .Y(new_n26683_));
  AND2X1   g24247(.A(pi1091), .B(pi0299), .Y(new_n26684_));
  INVX1    g24248(.A(new_n26684_), .Y(new_n26685_));
  AOI21X1  g24249(.A0(new_n26685_), .A1(new_n26679_), .B0(pi1157), .Y(new_n26686_));
  OAI21X1  g24250(.A0(new_n24992_), .A1(new_n2702_), .B0(new_n26664_), .Y(new_n26687_));
  AOI21X1  g24251(.A0(new_n26687_), .A1(new_n26672_), .B0(pi1156), .Y(new_n26688_));
  NOR3X1   g24252(.A(new_n26688_), .B(new_n12578_), .C(pi0211), .Y(new_n26689_));
  AOI21X1  g24253(.A0(new_n26689_), .A1(new_n26651_), .B0(new_n26686_), .Y(new_n26690_));
  AOI22X1  g24254(.A0(new_n26690_), .A1(new_n26683_), .B0(new_n26681_), .B1(new_n8422_), .Y(new_n26691_));
  OAI21X1  g24255(.A0(new_n26691_), .A1(new_n26601_), .B0(new_n6489_), .Y(new_n26692_));
  INVX1    g24256(.A(new_n26601_), .Y(new_n26693_));
  INVX1    g24257(.A(new_n26505_), .Y(new_n26694_));
  AND2X1   g24258(.A(new_n26502_), .B(new_n2702_), .Y(new_n26695_));
  NOR4X1   g24259(.A(new_n26695_), .B(new_n26574_), .C(new_n12578_), .D(pi0211), .Y(new_n26696_));
  AOI21X1  g24260(.A0(new_n26568_), .A1(pi0243), .B0(new_n26696_), .Y(new_n26697_));
  OAI21X1  g24261(.A0(new_n26694_), .A1(pi0243), .B0(new_n26697_), .Y(new_n26698_));
  NAND3X1  g24262(.A(new_n26515_), .B(new_n26512_), .C(new_n26574_), .Y(new_n26699_));
  MX2X1    g24263(.A(new_n12555_), .B(new_n12463_), .S0(new_n23173_), .Y(new_n26700_));
  INVX1    g24264(.A(new_n26700_), .Y(new_n26701_));
  OAI21X1  g24265(.A0(new_n26701_), .A1(new_n2702_), .B0(new_n8422_), .Y(new_n26702_));
  AOI21X1  g24266(.A0(new_n26514_), .A1(new_n26499_), .B0(new_n26702_), .Y(new_n26703_));
  AOI22X1  g24267(.A0(new_n26703_), .A1(new_n26699_), .B0(new_n26698_), .B1(pi0219), .Y(new_n26704_));
  AOI22X1  g24268(.A0(new_n26701_), .A1(new_n8422_), .B0(new_n24893_), .B1(pi1157), .Y(new_n26705_));
  MX2X1    g24269(.A(new_n26705_), .B(pi0243), .S0(new_n2702_), .Y(new_n26706_));
  OR2X1    g24270(.A(new_n26706_), .B(new_n26601_), .Y(new_n26707_));
  AND2X1   g24271(.A(new_n26707_), .B(po1038), .Y(new_n26708_));
  OAI21X1  g24272(.A0(new_n26704_), .A1(new_n26693_), .B0(new_n26708_), .Y(new_n26709_));
  AND3X1   g24273(.A(pi0283), .B(pi0275), .C(pi0272), .Y(new_n26710_));
  AND2X1   g24274(.A(new_n26710_), .B(pi0268), .Y(new_n26711_));
  AND2X1   g24275(.A(new_n26711_), .B(new_n26709_), .Y(new_n26712_));
  OAI21X1  g24276(.A0(new_n26692_), .A1(new_n26645_), .B0(new_n26712_), .Y(new_n26713_));
  NAND2X1  g24277(.A(new_n26691_), .B(new_n6489_), .Y(new_n26714_));
  AOI21X1  g24278(.A0(new_n26706_), .A1(po1038), .B0(new_n26711_), .Y(new_n26715_));
  AOI21X1  g24279(.A0(new_n26715_), .A1(new_n26714_), .B0(pi0230), .Y(new_n26716_));
  OR2X1    g24280(.A(new_n26705_), .B(new_n11660_), .Y(new_n26717_));
  OAI22X1  g24281(.A0(new_n8058_), .A1(pi1155), .B0(pi1156), .B1(new_n7937_), .Y(new_n26718_));
  AOI21X1  g24282(.A0(new_n25613_), .A1(pi0199), .B0(new_n26718_), .Y(new_n26719_));
  AOI21X1  g24283(.A0(new_n26719_), .A1(new_n11660_), .B0(new_n24814_), .Y(new_n26720_));
  AOI22X1  g24284(.A0(new_n26720_), .A1(new_n26717_), .B0(new_n26716_), .B1(new_n26713_), .Y(po0400));
  INVX1    g24285(.A(new_n25069_), .Y(new_n26722_));
  AOI22X1  g24286(.A0(new_n26206_), .A1(new_n26243_), .B0(new_n26164_), .B1(new_n26722_), .Y(new_n26723_));
  OAI21X1  g24287(.A0(new_n26723_), .A1(new_n26179_), .B0(pi0214), .Y(new_n26724_));
  AND2X1   g24288(.A(new_n26724_), .B(new_n26232_), .Y(new_n26725_));
  AOI21X1  g24289(.A0(new_n26137_), .A1(new_n24822_), .B0(new_n24823_), .Y(new_n26726_));
  INVX1    g24290(.A(new_n26726_), .Y(new_n26727_));
  AOI21X1  g24291(.A0(new_n26723_), .A1(new_n24849_), .B0(new_n26727_), .Y(new_n26728_));
  OAI21X1  g24292(.A0(new_n26170_), .A1(pi0299), .B0(new_n26728_), .Y(new_n26729_));
  NAND2X1  g24293(.A(new_n26729_), .B(new_n8422_), .Y(new_n26730_));
  OR2X1    g24294(.A(new_n25046_), .B(pi0211), .Y(new_n26731_));
  AOI21X1  g24295(.A0(new_n26170_), .A1(new_n2933_), .B0(new_n26731_), .Y(new_n26732_));
  OAI21X1  g24296(.A0(new_n26732_), .A1(new_n26227_), .B0(new_n26226_), .Y(new_n26733_));
  AND2X1   g24297(.A(new_n26733_), .B(new_n26204_), .Y(new_n26734_));
  OAI21X1  g24298(.A0(new_n26730_), .A1(new_n26725_), .B0(new_n26734_), .Y(new_n26735_));
  AND2X1   g24299(.A(new_n26728_), .B(new_n26163_), .Y(new_n26736_));
  AOI21X1  g24300(.A0(new_n26723_), .A1(pi0214), .B0(new_n26209_), .Y(new_n26737_));
  OR2X1    g24301(.A(new_n26737_), .B(pi0219), .Y(new_n26738_));
  OR2X1    g24302(.A(new_n25511_), .B(new_n2933_), .Y(new_n26739_));
  AND3X1   g24303(.A(new_n26739_), .B(new_n26192_), .C(pi1147), .Y(new_n26740_));
  OAI21X1  g24304(.A0(new_n26738_), .A1(new_n26736_), .B0(new_n26740_), .Y(new_n26741_));
  NAND4X1  g24305(.A(new_n26741_), .B(new_n26735_), .C(new_n25513_), .D(new_n24815_), .Y(new_n26742_));
  OAI21X1  g24306(.A0(new_n26247_), .A1(new_n24815_), .B0(new_n26742_), .Y(new_n26743_));
  AOI21X1  g24307(.A0(new_n26087_), .A1(new_n26119_), .B0(new_n26072_), .Y(new_n26744_));
  NOR2X1   g24308(.A(new_n26066_), .B(new_n2933_), .Y(new_n26745_));
  OAI21X1  g24309(.A0(pi1146), .A1(new_n23173_), .B0(pi0299), .Y(new_n26746_));
  OAI21X1  g24310(.A0(new_n26076_), .A1(new_n24877_), .B0(new_n25109_), .Y(new_n26747_));
  AOI21X1  g24311(.A0(new_n26746_), .A1(new_n24877_), .B0(new_n26747_), .Y(new_n26748_));
  OAI21X1  g24312(.A0(new_n26745_), .A1(new_n26120_), .B0(new_n26748_), .Y(new_n26749_));
  NOR2X1   g24313(.A(new_n26096_), .B(new_n25501_), .Y(new_n26750_));
  AOI21X1  g24314(.A0(new_n26750_), .A1(new_n26749_), .B0(po1038), .Y(new_n26751_));
  OAI21X1  g24315(.A0(new_n26751_), .A1(new_n26744_), .B0(pi0213), .Y(new_n26752_));
  AOI21X1  g24316(.A0(new_n25517_), .A1(new_n24815_), .B0(pi0209), .Y(new_n26753_));
  AOI22X1  g24317(.A0(new_n26753_), .A1(new_n26752_), .B0(new_n26743_), .B1(pi0209), .Y(new_n26754_));
  MX2X1    g24318(.A(new_n26754_), .B(pi0244), .S0(new_n24814_), .Y(po0401));
  NOR4X1   g24319(.A(new_n24818_), .B(new_n7963_), .C(new_n6489_), .D(new_n3140_), .Y(new_n26756_));
  NOR2X1   g24320(.A(new_n26756_), .B(pi1147), .Y(new_n26757_));
  OAI21X1  g24321(.A0(new_n26007_), .A1(new_n25818_), .B0(new_n26757_), .Y(new_n26758_));
  OR3X1    g24322(.A(new_n26466_), .B(new_n24816_), .C(pi0211), .Y(new_n26759_));
  AOI21X1  g24323(.A0(new_n26759_), .A1(new_n26478_), .B0(po1038), .Y(new_n26760_));
  NOR2X1   g24324(.A(new_n26078_), .B(new_n24849_), .Y(new_n26761_));
  OAI21X1  g24325(.A0(new_n26467_), .A1(pi0299), .B0(new_n26761_), .Y(new_n26762_));
  NAND2X1  g24326(.A(new_n26762_), .B(pi0212), .Y(new_n26763_));
  AND2X1   g24327(.A(new_n26461_), .B(new_n2933_), .Y(new_n26764_));
  OAI21X1  g24328(.A0(new_n26764_), .A1(pi0211), .B0(new_n26476_), .Y(new_n26765_));
  NOR2X1   g24329(.A(new_n26765_), .B(pi0214), .Y(new_n26766_));
  AOI21X1  g24330(.A0(new_n26765_), .A1(new_n26472_), .B0(pi0219), .Y(new_n26767_));
  OAI21X1  g24331(.A0(new_n26766_), .A1(new_n26763_), .B0(new_n26767_), .Y(new_n26768_));
  AOI21X1  g24332(.A0(new_n26768_), .A1(new_n26760_), .B0(new_n26758_), .Y(new_n26769_));
  NOR3X1   g24333(.A(new_n26756_), .B(new_n25804_), .C(new_n25993_), .Y(new_n26770_));
  INVX1    g24334(.A(new_n26770_), .Y(new_n26771_));
  MX2X1    g24335(.A(new_n26764_), .B(new_n26466_), .S0(pi0211), .Y(new_n26772_));
  MX2X1    g24336(.A(new_n26772_), .B(new_n26764_), .S0(new_n24849_), .Y(new_n26773_));
  OR3X1    g24337(.A(new_n26764_), .B(new_n26471_), .C(pi0212), .Y(new_n26774_));
  AND2X1   g24338(.A(new_n26774_), .B(new_n8422_), .Y(new_n26775_));
  OAI21X1  g24339(.A0(new_n26773_), .A1(new_n24823_), .B0(new_n26775_), .Y(new_n26776_));
  AOI21X1  g24340(.A0(new_n26776_), .A1(new_n26760_), .B0(new_n26771_), .Y(new_n26777_));
  NOR3X1   g24341(.A(new_n26777_), .B(new_n26769_), .C(new_n26084_), .Y(new_n26778_));
  AOI21X1  g24342(.A0(new_n26001_), .A1(pi1147), .B0(new_n26770_), .Y(new_n26779_));
  AND3X1   g24343(.A(new_n26470_), .B(new_n26459_), .C(new_n26040_), .Y(new_n26780_));
  MX2X1    g24344(.A(new_n26780_), .B(new_n26772_), .S0(pi0214), .Y(new_n26781_));
  OR3X1    g24345(.A(new_n26780_), .B(new_n26471_), .C(pi0212), .Y(new_n26782_));
  AND2X1   g24346(.A(new_n26782_), .B(new_n8422_), .Y(new_n26783_));
  OAI21X1  g24347(.A0(new_n26781_), .A1(new_n24823_), .B0(new_n26783_), .Y(new_n26784_));
  AOI21X1  g24348(.A0(new_n26784_), .A1(new_n26760_), .B0(new_n26779_), .Y(new_n26785_));
  INVX1    g24349(.A(new_n26757_), .Y(new_n26786_));
  AOI21X1  g24350(.A0(new_n26477_), .A1(new_n24823_), .B0(pi0219), .Y(new_n26787_));
  OAI21X1  g24351(.A0(new_n26763_), .A1(new_n26471_), .B0(new_n26787_), .Y(new_n26788_));
  AOI21X1  g24352(.A0(new_n26788_), .A1(new_n26760_), .B0(new_n26786_), .Y(new_n26789_));
  NOR3X1   g24353(.A(new_n26789_), .B(new_n26785_), .C(pi1148), .Y(new_n26790_));
  OAI21X1  g24354(.A0(new_n26790_), .A1(new_n26778_), .B0(pi0213), .Y(new_n26791_));
  AOI21X1  g24355(.A0(new_n26481_), .A1(new_n24815_), .B0(pi0209), .Y(new_n26792_));
  AOI21X1  g24356(.A0(pi1146), .A1(pi0199), .B0(pi0200), .Y(new_n26793_));
  OR4X1    g24357(.A(new_n26793_), .B(new_n26152_), .C(pi0299), .D(new_n22660_), .Y(new_n26794_));
  OAI21X1  g24358(.A0(new_n24961_), .A1(new_n3140_), .B0(new_n26794_), .Y(new_n26795_));
  AND2X1   g24359(.A(new_n26795_), .B(pi0208), .Y(new_n26796_));
  AND3X1   g24360(.A(new_n3140_), .B(new_n7937_), .C(pi0199), .Y(new_n26797_));
  NOR4X1   g24361(.A(new_n26797_), .B(new_n26152_), .C(pi0299), .D(new_n22959_), .Y(new_n26798_));
  NOR2X1   g24362(.A(new_n26798_), .B(pi0207), .Y(new_n26799_));
  NOR4X1   g24363(.A(new_n26799_), .B(new_n26797_), .C(new_n24917_), .D(new_n7826_), .Y(new_n26800_));
  AND2X1   g24364(.A(new_n26106_), .B(new_n22959_), .Y(new_n26801_));
  NOR3X1   g24365(.A(new_n26801_), .B(new_n26800_), .C(new_n26796_), .Y(new_n26802_));
  NOR2X1   g24366(.A(new_n26802_), .B(pi0299), .Y(new_n26803_));
  INVX1    g24367(.A(new_n26803_), .Y(new_n26804_));
  AOI21X1  g24368(.A0(new_n26804_), .A1(new_n24849_), .B0(pi0212), .Y(new_n26805_));
  NOR3X1   g24369(.A(new_n26793_), .B(new_n26152_), .C(pi0299), .Y(new_n26806_));
  OAI21X1  g24370(.A0(new_n25654_), .A1(new_n7826_), .B0(new_n26806_), .Y(new_n26807_));
  NOR2X1   g24371(.A(new_n26806_), .B(pi0299), .Y(new_n26808_));
  NOR2X1   g24372(.A(new_n26808_), .B(new_n26802_), .Y(new_n26809_));
  NOR3X1   g24373(.A(new_n26809_), .B(pi0299), .C(pi0211), .Y(new_n26810_));
  AOI21X1  g24374(.A0(new_n26807_), .A1(pi0211), .B0(new_n26810_), .Y(new_n26811_));
  OR2X1    g24375(.A(new_n26811_), .B(new_n26803_), .Y(new_n26812_));
  AOI21X1  g24376(.A0(new_n26812_), .A1(new_n26805_), .B0(pi0219), .Y(new_n26813_));
  NOR3X1   g24377(.A(new_n26803_), .B(new_n26078_), .C(new_n24849_), .Y(new_n26814_));
  OAI21X1  g24378(.A0(new_n26812_), .A1(pi0214), .B0(pi0212), .Y(new_n26815_));
  OAI21X1  g24379(.A0(new_n26815_), .A1(new_n26814_), .B0(new_n26813_), .Y(new_n26816_));
  AOI21X1  g24380(.A0(new_n26803_), .A1(new_n25162_), .B0(new_n8422_), .Y(new_n26817_));
  OR2X1    g24381(.A(new_n26802_), .B(new_n25162_), .Y(new_n26818_));
  AOI21X1  g24382(.A0(new_n26818_), .A1(new_n26817_), .B0(po1038), .Y(new_n26819_));
  AOI21X1  g24383(.A0(new_n26819_), .A1(new_n26816_), .B0(new_n26758_), .Y(new_n26820_));
  NOR2X1   g24384(.A(new_n26797_), .B(new_n24933_), .Y(new_n26821_));
  NOR2X1   g24385(.A(new_n26821_), .B(new_n7826_), .Y(new_n26822_));
  NOR4X1   g24386(.A(new_n26797_), .B(new_n26152_), .C(pi0299), .D(new_n22660_), .Y(new_n26823_));
  INVX1    g24387(.A(new_n26823_), .Y(new_n26824_));
  AOI21X1  g24388(.A0(new_n26824_), .A1(new_n25116_), .B0(new_n26822_), .Y(new_n26825_));
  OR2X1    g24389(.A(new_n26825_), .B(pi0214), .Y(new_n26826_));
  AND2X1   g24390(.A(new_n26826_), .B(new_n24823_), .Y(new_n26827_));
  NOR3X1   g24391(.A(new_n26793_), .B(new_n25130_), .C(pi0299), .Y(new_n26828_));
  AOI21X1  g24392(.A0(new_n26828_), .A1(new_n22660_), .B0(new_n26106_), .Y(new_n26829_));
  AOI21X1  g24393(.A0(new_n26829_), .A1(new_n26824_), .B0(new_n22959_), .Y(new_n26830_));
  AOI21X1  g24394(.A0(new_n26821_), .A1(new_n24844_), .B0(new_n26798_), .Y(new_n26831_));
  INVX1    g24395(.A(new_n26831_), .Y(new_n26832_));
  NOR3X1   g24396(.A(new_n26832_), .B(new_n26830_), .C(pi0299), .Y(new_n26833_));
  INVX1    g24397(.A(new_n26833_), .Y(new_n26834_));
  AOI21X1  g24398(.A0(new_n26834_), .A1(new_n26827_), .B0(pi0219), .Y(new_n26835_));
  OR2X1    g24399(.A(new_n26833_), .B(new_n24823_), .Y(new_n26836_));
  AOI21X1  g24400(.A0(new_n26830_), .A1(new_n2933_), .B0(new_n26832_), .Y(new_n26837_));
  AND3X1   g24401(.A(new_n26837_), .B(new_n26465_), .C(new_n25032_), .Y(new_n26838_));
  OR2X1    g24402(.A(new_n26838_), .B(new_n26836_), .Y(new_n26839_));
  AOI21X1  g24403(.A0(new_n26825_), .A1(new_n25162_), .B0(new_n8422_), .Y(new_n26840_));
  INVX1    g24404(.A(new_n26840_), .Y(new_n26841_));
  AOI21X1  g24405(.A0(new_n26837_), .A1(new_n26465_), .B0(new_n25162_), .Y(new_n26842_));
  OAI21X1  g24406(.A0(new_n26842_), .A1(new_n26841_), .B0(new_n6489_), .Y(new_n26843_));
  AOI21X1  g24407(.A0(new_n26839_), .A1(new_n26835_), .B0(new_n26843_), .Y(new_n26844_));
  OAI21X1  g24408(.A0(new_n26844_), .A1(new_n26771_), .B0(pi1148), .Y(new_n26845_));
  INVX1    g24409(.A(new_n26828_), .Y(new_n26846_));
  AOI22X1  g24410(.A0(new_n26846_), .A1(new_n7827_), .B0(new_n26824_), .B1(new_n25116_), .Y(new_n26847_));
  NOR2X1   g24411(.A(new_n26847_), .B(new_n9446_), .Y(new_n26848_));
  AOI21X1  g24412(.A0(new_n26847_), .A1(new_n24849_), .B0(pi0212), .Y(new_n26849_));
  OAI21X1  g24413(.A0(new_n26848_), .A1(new_n24849_), .B0(new_n26849_), .Y(new_n26850_));
  OAI22X1  g24414(.A0(new_n26846_), .A1(new_n25880_), .B0(new_n26465_), .B1(pi0208), .Y(new_n26851_));
  NOR3X1   g24415(.A(new_n26851_), .B(new_n26830_), .C(pi0299), .Y(new_n26852_));
  NOR2X1   g24416(.A(new_n26852_), .B(new_n24849_), .Y(new_n26853_));
  NOR2X1   g24417(.A(new_n26833_), .B(pi0211), .Y(new_n26854_));
  NOR2X1   g24418(.A(new_n26854_), .B(new_n26825_), .Y(new_n26855_));
  INVX1    g24419(.A(new_n26855_), .Y(new_n26856_));
  AOI21X1  g24420(.A0(new_n26856_), .A1(new_n26853_), .B0(new_n24823_), .Y(new_n26857_));
  OAI21X1  g24421(.A0(new_n26848_), .A1(pi0214), .B0(new_n26857_), .Y(new_n26858_));
  AOI21X1  g24422(.A0(new_n26858_), .A1(new_n26850_), .B0(pi0219), .Y(new_n26859_));
  OAI21X1  g24423(.A0(new_n25036_), .A1(pi1146), .B0(new_n26142_), .Y(new_n26860_));
  NOR2X1   g24424(.A(new_n26851_), .B(new_n26830_), .Y(new_n26861_));
  AOI21X1  g24425(.A0(new_n26847_), .A1(new_n25188_), .B0(new_n24817_), .Y(new_n26862_));
  AND3X1   g24426(.A(new_n26847_), .B(new_n24849_), .C(new_n24823_), .Y(new_n26863_));
  NOR2X1   g24427(.A(new_n26863_), .B(new_n8422_), .Y(new_n26864_));
  OAI21X1  g24428(.A0(new_n26862_), .A1(new_n26861_), .B0(new_n26864_), .Y(new_n26865_));
  NAND2X1  g24429(.A(new_n26865_), .B(new_n6489_), .Y(new_n26866_));
  AOI21X1  g24430(.A0(new_n26860_), .A1(new_n26859_), .B0(new_n26866_), .Y(new_n26867_));
  AND2X1   g24431(.A(new_n7962_), .B(pi0299), .Y(new_n26868_));
  OAI21X1  g24432(.A0(new_n26803_), .A1(new_n26868_), .B0(new_n26795_), .Y(new_n26869_));
  AND2X1   g24433(.A(new_n26869_), .B(new_n8422_), .Y(new_n26870_));
  NAND2X1  g24434(.A(new_n26807_), .B(pi0219), .Y(new_n26871_));
  AOI21X1  g24435(.A0(new_n26807_), .A1(pi0211), .B0(new_n24816_), .Y(new_n26872_));
  AOI22X1  g24436(.A0(new_n26872_), .A1(new_n26809_), .B0(new_n26871_), .B1(new_n25306_), .Y(new_n26873_));
  OR3X1    g24437(.A(new_n26873_), .B(new_n26870_), .C(po1038), .Y(new_n26874_));
  AOI21X1  g24438(.A0(new_n26874_), .A1(new_n26757_), .B0(pi1148), .Y(new_n26875_));
  OAI21X1  g24439(.A0(new_n26867_), .A1(new_n26779_), .B0(new_n26875_), .Y(new_n26876_));
  OAI21X1  g24440(.A0(new_n26845_), .A1(new_n26820_), .B0(new_n26876_), .Y(new_n26877_));
  NAND2X1  g24441(.A(new_n26877_), .B(pi0213), .Y(new_n26878_));
  MX2X1    g24442(.A(new_n26802_), .B(new_n26063_), .S0(pi0299), .Y(new_n26879_));
  OAI21X1  g24443(.A0(new_n26809_), .A1(pi0299), .B0(pi0214), .Y(new_n26880_));
  OAI22X1  g24444(.A0(new_n26880_), .A1(new_n26879_), .B0(new_n26807_), .B1(pi0214), .Y(new_n26881_));
  AND2X1   g24445(.A(new_n26446_), .B(pi0299), .Y(new_n26882_));
  OAI21X1  g24446(.A0(new_n26882_), .A1(new_n26803_), .B0(pi0212), .Y(new_n26883_));
  OAI21X1  g24447(.A0(new_n26883_), .A1(new_n26808_), .B0(new_n8422_), .Y(new_n26884_));
  AOI21X1  g24448(.A0(new_n26881_), .A1(new_n24823_), .B0(new_n26884_), .Y(new_n26885_));
  MX2X1    g24449(.A(new_n26809_), .B(pi1144), .S0(pi0299), .Y(new_n26886_));
  OR2X1    g24450(.A(new_n26886_), .B(pi0211), .Y(new_n26887_));
  AOI22X1  g24451(.A0(new_n26887_), .A1(new_n26872_), .B0(new_n26871_), .B1(new_n25306_), .Y(new_n26888_));
  NOR3X1   g24452(.A(new_n26888_), .B(new_n26885_), .C(new_n26218_), .Y(new_n26889_));
  INVX1    g24453(.A(new_n26853_), .Y(new_n26890_));
  INVX1    g24454(.A(new_n26837_), .Y(new_n26891_));
  NOR2X1   g24455(.A(new_n26891_), .B(new_n26076_), .Y(new_n26892_));
  NOR2X1   g24456(.A(new_n26892_), .B(new_n26890_), .Y(new_n26893_));
  AOI21X1  g24457(.A0(new_n26847_), .A1(new_n24849_), .B0(new_n26893_), .Y(new_n26894_));
  INVX1    g24458(.A(new_n26852_), .Y(new_n26895_));
  INVX1    g24459(.A(new_n26882_), .Y(new_n26896_));
  AOI21X1  g24460(.A0(new_n26896_), .A1(new_n26837_), .B0(new_n24823_), .Y(new_n26897_));
  AOI21X1  g24461(.A0(new_n26897_), .A1(new_n26895_), .B0(pi0219), .Y(new_n26898_));
  OAI21X1  g24462(.A0(new_n26894_), .A1(pi0212), .B0(new_n26898_), .Y(new_n26899_));
  INVX1    g24463(.A(new_n26862_), .Y(new_n26900_));
  AOI21X1  g24464(.A0(new_n26837_), .A1(new_n25073_), .B0(new_n26852_), .Y(new_n26901_));
  OAI21X1  g24465(.A0(new_n26901_), .A1(pi0211), .B0(new_n26900_), .Y(new_n26902_));
  NAND3X1  g24466(.A(new_n5102_), .B(pi1147), .C(new_n2436_), .Y(new_n26903_));
  AOI21X1  g24467(.A0(new_n26902_), .A1(new_n26864_), .B0(new_n26903_), .Y(new_n26904_));
  AND2X1   g24468(.A(new_n26904_), .B(new_n26899_), .Y(new_n26905_));
  OR4X1    g24469(.A(new_n26905_), .B(new_n26889_), .C(new_n26451_), .D(pi1148), .Y(new_n26906_));
  OAI21X1  g24470(.A0(new_n26803_), .A1(new_n26076_), .B0(new_n26805_), .Y(new_n26907_));
  AND3X1   g24471(.A(new_n26907_), .B(new_n26883_), .C(new_n8422_), .Y(new_n26908_));
  INVX1    g24472(.A(new_n26817_), .Y(new_n26909_));
  NOR4X1   g24473(.A(new_n26801_), .B(new_n26800_), .C(new_n26796_), .D(pi0299), .Y(new_n26910_));
  NOR2X1   g24474(.A(new_n26910_), .B(new_n25162_), .Y(new_n26911_));
  AOI21X1  g24475(.A0(new_n26911_), .A1(new_n26722_), .B0(new_n26909_), .Y(new_n26912_));
  OR3X1    g24476(.A(new_n26912_), .B(new_n26908_), .C(new_n26218_), .Y(new_n26913_));
  OR3X1    g24477(.A(new_n26891_), .B(new_n26076_), .C(new_n24849_), .Y(new_n26914_));
  AND2X1   g24478(.A(new_n26914_), .B(new_n26827_), .Y(new_n26915_));
  OR3X1    g24479(.A(new_n26915_), .B(new_n26897_), .C(pi0219), .Y(new_n26916_));
  OAI21X1  g24480(.A0(new_n26891_), .A1(new_n25068_), .B0(new_n24817_), .Y(new_n26917_));
  AOI21X1  g24481(.A0(new_n26917_), .A1(new_n26840_), .B0(new_n26903_), .Y(new_n26918_));
  OR2X1    g24482(.A(new_n26451_), .B(new_n26084_), .Y(new_n26919_));
  AOI21X1  g24483(.A0(new_n26918_), .A1(new_n26916_), .B0(new_n26919_), .Y(new_n26920_));
  AOI21X1  g24484(.A0(new_n26920_), .A1(new_n26913_), .B0(pi0213), .Y(new_n26921_));
  AOI21X1  g24485(.A0(new_n26921_), .A1(new_n26906_), .B0(new_n24866_), .Y(new_n26922_));
  AOI22X1  g24486(.A0(new_n26922_), .A1(new_n26878_), .B0(new_n26792_), .B1(new_n26791_), .Y(new_n26923_));
  MX2X1    g24487(.A(new_n26923_), .B(pi0245), .S0(new_n24814_), .Y(po0402));
  AOI21X1  g24488(.A0(new_n25964_), .A1(pi1150), .B0(new_n25955_), .Y(new_n26925_));
  OAI21X1  g24489(.A0(new_n26003_), .A1(pi1150), .B0(new_n26925_), .Y(new_n26926_));
  AND3X1   g24490(.A(new_n26024_), .B(new_n26009_), .C(pi1150), .Y(new_n26927_));
  OAI21X1  g24491(.A0(new_n26058_), .A1(pi1150), .B0(new_n25955_), .Y(new_n26928_));
  OAI21X1  g24492(.A0(new_n26928_), .A1(new_n26927_), .B0(new_n26926_), .Y(new_n26929_));
  NOR3X1   g24493(.A(new_n25991_), .B(new_n25968_), .C(pi1150), .Y(new_n26930_));
  OAI21X1  g24494(.A0(new_n25954_), .A1(new_n26280_), .B0(pi1149), .Y(new_n26931_));
  OR2X1    g24495(.A(new_n26280_), .B(pi1149), .Y(new_n26932_));
  OAI22X1  g24496(.A0(new_n26932_), .A1(new_n26028_), .B0(new_n26931_), .B1(new_n26930_), .Y(new_n26933_));
  MX2X1    g24497(.A(new_n26933_), .B(new_n26929_), .S0(pi1148), .Y(new_n26934_));
  NAND2X1  g24498(.A(new_n26934_), .B(pi0213), .Y(new_n26935_));
  AND2X1   g24499(.A(new_n26771_), .B(new_n26758_), .Y(new_n26936_));
  AOI21X1  g24500(.A0(new_n26465_), .A1(pi0219), .B0(new_n26053_), .Y(new_n26937_));
  AND2X1   g24501(.A(new_n26032_), .B(new_n7871_), .Y(new_n26938_));
  NOR2X1   g24502(.A(new_n26938_), .B(new_n25999_), .Y(new_n26939_));
  NOR2X1   g24503(.A(new_n26939_), .B(new_n26937_), .Y(new_n26940_));
  AOI21X1  g24504(.A0(new_n9446_), .A1(new_n3140_), .B0(new_n26034_), .Y(new_n26941_));
  OAI22X1  g24505(.A0(new_n26941_), .A1(new_n25383_), .B0(new_n26033_), .B1(new_n25959_), .Y(new_n26942_));
  AOI21X1  g24506(.A0(new_n26942_), .A1(new_n8422_), .B0(new_n26940_), .Y(new_n26943_));
  INVX1    g24507(.A(new_n26758_), .Y(new_n26944_));
  NOR3X1   g24508(.A(new_n26033_), .B(pi0299), .C(pi0219), .Y(new_n26945_));
  OR2X1    g24509(.A(new_n26050_), .B(new_n26945_), .Y(new_n26946_));
  AOI21X1  g24510(.A0(new_n26946_), .A1(new_n26944_), .B0(pi1150), .Y(new_n26947_));
  OAI21X1  g24511(.A0(new_n26943_), .A1(new_n26936_), .B0(new_n26947_), .Y(new_n26948_));
  OR2X1    g24512(.A(new_n26937_), .B(new_n26102_), .Y(new_n26949_));
  INVX1    g24513(.A(new_n26274_), .Y(new_n26950_));
  OAI21X1  g24514(.A0(new_n25655_), .A1(pi0212), .B0(new_n8422_), .Y(new_n26951_));
  NOR2X1   g24515(.A(new_n26951_), .B(new_n26282_), .Y(new_n26952_));
  OAI21X1  g24516(.A0(new_n26950_), .A1(new_n26109_), .B0(new_n26952_), .Y(new_n26953_));
  AOI21X1  g24517(.A0(new_n26953_), .A1(new_n26949_), .B0(new_n26771_), .Y(new_n26954_));
  NOR2X1   g24518(.A(new_n26015_), .B(pi0219), .Y(new_n26955_));
  AND3X1   g24519(.A(new_n26108_), .B(new_n26010_), .C(pi0214), .Y(new_n26956_));
  OAI21X1  g24520(.A0(new_n26016_), .A1(pi0214), .B0(pi0212), .Y(new_n26957_));
  OAI21X1  g24521(.A0(new_n26957_), .A1(new_n26956_), .B0(new_n26955_), .Y(new_n26958_));
  AOI21X1  g24522(.A0(new_n26958_), .A1(new_n26949_), .B0(new_n26758_), .Y(new_n26959_));
  OR3X1    g24523(.A(new_n26959_), .B(new_n26954_), .C(new_n26280_), .Y(new_n26960_));
  AOI21X1  g24524(.A0(new_n26960_), .A1(new_n26948_), .B0(new_n26084_), .Y(new_n26961_));
  OR2X1    g24525(.A(new_n26062_), .B(pi0219), .Y(new_n26962_));
  AND3X1   g24526(.A(new_n26962_), .B(new_n26937_), .C(new_n26375_), .Y(new_n26963_));
  OAI22X1  g24527(.A0(new_n26963_), .A1(new_n26786_), .B0(new_n26937_), .B1(new_n26779_), .Y(new_n26964_));
  NAND4X1  g24528(.A(new_n25115_), .B(new_n11660_), .C(new_n8055_), .D(pi1150), .Y(new_n26965_));
  NAND3X1  g24529(.A(new_n25204_), .B(new_n25115_), .C(pi1150), .Y(new_n26966_));
  OR4X1    g24530(.A(new_n2933_), .B(new_n24849_), .C(pi0212), .D(new_n23173_), .Y(new_n26967_));
  NAND4X1  g24531(.A(new_n26967_), .B(new_n26966_), .C(new_n26860_), .D(new_n8422_), .Y(new_n26968_));
  OAI21X1  g24532(.A0(new_n26968_), .A1(new_n26779_), .B0(new_n26084_), .Y(new_n26969_));
  AOI21X1  g24533(.A0(new_n26965_), .A1(new_n26964_), .B0(new_n26969_), .Y(new_n26970_));
  OAI21X1  g24534(.A0(new_n26970_), .A1(new_n26961_), .B0(new_n25955_), .Y(new_n26971_));
  AOI21X1  g24535(.A0(new_n26137_), .A1(new_n26062_), .B0(new_n25971_), .Y(new_n26972_));
  AOI22X1  g24536(.A0(new_n25988_), .A1(new_n6489_), .B0(new_n25979_), .B1(new_n26052_), .Y(new_n26973_));
  INVX1    g24537(.A(new_n26973_), .Y(new_n26974_));
  OAI21X1  g24538(.A0(new_n25988_), .A1(pi1146), .B0(new_n26974_), .Y(new_n26975_));
  AOI21X1  g24539(.A0(new_n26972_), .A1(new_n25987_), .B0(new_n26975_), .Y(new_n26976_));
  OAI22X1  g24540(.A0(new_n25972_), .A1(new_n25971_), .B0(new_n25688_), .B1(pi0212), .Y(new_n26977_));
  AOI21X1  g24541(.A0(new_n26977_), .A1(new_n8422_), .B0(new_n26973_), .Y(new_n26978_));
  OAI21X1  g24542(.A0(new_n25971_), .A1(pi1146), .B0(new_n26978_), .Y(new_n26979_));
  AOI21X1  g24543(.A0(new_n26979_), .A1(new_n26757_), .B0(pi1150), .Y(new_n26980_));
  OAI21X1  g24544(.A0(new_n26976_), .A1(new_n26779_), .B0(new_n26980_), .Y(new_n26981_));
  OR4X1    g24545(.A(new_n25719_), .B(new_n25275_), .C(new_n5103_), .D(pi0057), .Y(new_n26982_));
  OR3X1    g24546(.A(new_n26403_), .B(new_n25720_), .C(pi0214), .Y(new_n26983_));
  AOI21X1  g24547(.A0(new_n26983_), .A1(new_n25952_), .B0(pi0219), .Y(new_n26984_));
  OAI21X1  g24548(.A0(new_n26403_), .A1(new_n25720_), .B0(new_n25945_), .Y(new_n26985_));
  OAI21X1  g24549(.A0(new_n26985_), .A1(pi0212), .B0(new_n26984_), .Y(new_n26986_));
  NAND3X1  g24550(.A(new_n25705_), .B(new_n2933_), .C(pi0208), .Y(new_n26987_));
  NAND3X1  g24551(.A(new_n26987_), .B(new_n26465_), .C(new_n25942_), .Y(new_n26988_));
  AOI21X1  g24552(.A0(new_n26123_), .A1(new_n8423_), .B0(new_n26937_), .Y(new_n26989_));
  AOI21X1  g24553(.A0(new_n26985_), .A1(new_n26984_), .B0(new_n26989_), .Y(new_n26990_));
  OAI21X1  g24554(.A0(new_n26988_), .A1(new_n26986_), .B0(new_n26990_), .Y(new_n26991_));
  NOR2X1   g24555(.A(new_n26419_), .B(new_n26418_), .Y(new_n26992_));
  OAI21X1  g24556(.A0(new_n25951_), .A1(new_n25946_), .B0(new_n8422_), .Y(new_n26993_));
  OAI21X1  g24557(.A0(new_n26993_), .A1(new_n26992_), .B0(new_n26123_), .Y(new_n26994_));
  AOI21X1  g24558(.A0(new_n26991_), .A1(new_n26982_), .B0(new_n26994_), .Y(new_n26995_));
  INVX1    g24559(.A(new_n26779_), .Y(new_n26996_));
  AOI21X1  g24560(.A0(new_n26991_), .A1(new_n26996_), .B0(new_n26280_), .Y(new_n26997_));
  OAI21X1  g24561(.A0(new_n26995_), .A1(new_n26786_), .B0(new_n26997_), .Y(new_n26998_));
  AND3X1   g24562(.A(new_n26998_), .B(new_n26981_), .C(new_n26084_), .Y(new_n26999_));
  INVX1    g24563(.A(new_n26936_), .Y(new_n27000_));
  NOR4X1   g24564(.A(new_n26046_), .B(new_n26045_), .C(new_n26038_), .D(new_n24823_), .Y(new_n27001_));
  INVX1    g24565(.A(new_n27001_), .Y(new_n27002_));
  AOI21X1  g24566(.A0(new_n27002_), .A1(new_n26042_), .B0(new_n26944_), .Y(new_n27003_));
  NOR4X1   g24567(.A(new_n26078_), .B(new_n25733_), .C(new_n25732_), .D(new_n24849_), .Y(new_n27004_));
  NOR3X1   g24568(.A(new_n27004_), .B(new_n26046_), .C(new_n24823_), .Y(new_n27005_));
  OR3X1    g24569(.A(new_n27005_), .B(new_n26048_), .C(pi0219), .Y(new_n27006_));
  OAI22X1  g24570(.A0(new_n27006_), .A1(new_n27003_), .B0(new_n26937_), .B1(new_n25998_), .Y(new_n27007_));
  AOI21X1  g24571(.A0(new_n27007_), .A1(new_n27000_), .B0(pi1150), .Y(new_n27008_));
  NOR3X1   g24572(.A(new_n26963_), .B(new_n26758_), .C(new_n26145_), .Y(new_n27009_));
  OAI21X1  g24573(.A0(new_n26136_), .A1(new_n24849_), .B0(new_n26141_), .Y(new_n27010_));
  NOR2X1   g24574(.A(new_n26139_), .B(pi0219), .Y(new_n27011_));
  AOI21X1  g24575(.A0(new_n27011_), .A1(new_n27010_), .B0(new_n26135_), .Y(new_n27012_));
  NOR4X1   g24576(.A(new_n25960_), .B(new_n24818_), .C(po1038), .D(new_n3140_), .Y(new_n27013_));
  OR4X1    g24577(.A(new_n27013_), .B(new_n26756_), .C(new_n25804_), .D(new_n25993_), .Y(new_n27014_));
  OAI21X1  g24578(.A0(new_n27014_), .A1(new_n27012_), .B0(pi1150), .Y(new_n27015_));
  OAI21X1  g24579(.A0(new_n27015_), .A1(new_n27009_), .B0(pi1148), .Y(new_n27016_));
  OAI21X1  g24580(.A0(new_n27016_), .A1(new_n27008_), .B0(pi1149), .Y(new_n27017_));
  OAI21X1  g24581(.A0(new_n27017_), .A1(new_n26999_), .B0(new_n26971_), .Y(new_n27018_));
  AOI21X1  g24582(.A0(new_n27018_), .A1(new_n24815_), .B0(new_n24866_), .Y(new_n27019_));
  INVX1    g24583(.A(new_n26807_), .Y(new_n27020_));
  AOI21X1  g24584(.A0(new_n27020_), .A1(new_n24849_), .B0(pi0212), .Y(new_n27021_));
  AND2X1   g24585(.A(new_n26807_), .B(new_n26040_), .Y(new_n27022_));
  OAI21X1  g24586(.A0(new_n27022_), .A1(new_n24849_), .B0(new_n27021_), .Y(new_n27023_));
  AOI21X1  g24587(.A0(new_n26811_), .A1(pi0214), .B0(new_n24823_), .Y(new_n27024_));
  OAI21X1  g24588(.A0(new_n27022_), .A1(pi0214), .B0(new_n27024_), .Y(new_n27025_));
  AOI21X1  g24589(.A0(new_n27025_), .A1(new_n27023_), .B0(pi0219), .Y(new_n27026_));
  NAND2X1  g24590(.A(new_n26871_), .B(new_n26204_), .Y(new_n27027_));
  NOR2X1   g24591(.A(new_n27027_), .B(new_n27026_), .Y(new_n27028_));
  NOR2X1   g24592(.A(new_n26847_), .B(new_n8422_), .Y(new_n27029_));
  NOR3X1   g24593(.A(new_n27029_), .B(new_n26903_), .C(new_n26859_), .Y(new_n27030_));
  OR4X1    g24594(.A(new_n27030_), .B(new_n27028_), .C(new_n25968_), .D(pi1150), .Y(new_n27031_));
  OAI21X1  g24595(.A0(new_n26809_), .A1(pi0299), .B0(new_n24849_), .Y(new_n27032_));
  AOI22X1  g24596(.A0(new_n27032_), .A1(new_n27024_), .B0(new_n27021_), .B1(new_n26880_), .Y(new_n27033_));
  OAI21X1  g24597(.A0(new_n27033_), .A1(pi0219), .B0(new_n26871_), .Y(new_n27034_));
  OR2X1    g24598(.A(new_n26852_), .B(pi0214), .Y(new_n27035_));
  AOI22X1  g24599(.A0(new_n27035_), .A1(new_n26857_), .B0(new_n26890_), .B1(new_n26849_), .Y(new_n27036_));
  MX2X1    g24600(.A(new_n27036_), .B(new_n26847_), .S0(pi0219), .Y(new_n27037_));
  OAI21X1  g24601(.A0(new_n27037_), .A1(new_n25993_), .B0(new_n6489_), .Y(new_n27038_));
  AOI21X1  g24602(.A0(new_n27034_), .A1(new_n25993_), .B0(new_n27038_), .Y(new_n27039_));
  OR2X1    g24603(.A(new_n25804_), .B(new_n26280_), .Y(new_n27040_));
  OAI21X1  g24604(.A0(new_n27040_), .A1(new_n27039_), .B0(new_n27031_), .Y(new_n27041_));
  AND2X1   g24605(.A(new_n26070_), .B(pi1150), .Y(new_n27042_));
  NOR3X1   g24606(.A(new_n26808_), .B(new_n26802_), .C(pi1147), .Y(new_n27043_));
  OR2X1    g24607(.A(new_n27043_), .B(new_n22572_), .Y(new_n27044_));
  NOR2X1   g24608(.A(new_n26847_), .B(new_n25993_), .Y(new_n27045_));
  OAI21X1  g24609(.A0(new_n27042_), .A1(new_n26807_), .B0(new_n25993_), .Y(new_n27046_));
  NAND2X1  g24610(.A(new_n27046_), .B(new_n6489_), .Y(new_n27047_));
  OAI21X1  g24611(.A0(new_n27047_), .A1(new_n27045_), .B0(new_n25955_), .Y(new_n27048_));
  AOI21X1  g24612(.A0(new_n27044_), .A1(new_n27042_), .B0(new_n27048_), .Y(new_n27049_));
  AOI21X1  g24613(.A0(new_n27041_), .A1(pi1149), .B0(new_n27049_), .Y(new_n27050_));
  OAI21X1  g24614(.A0(new_n26911_), .A1(new_n26909_), .B0(new_n26204_), .Y(new_n27051_));
  INVX1    g24615(.A(new_n27051_), .Y(new_n27052_));
  NOR4X1   g24616(.A(new_n27020_), .B(new_n26803_), .C(new_n9446_), .D(new_n24849_), .Y(new_n27053_));
  OAI21X1  g24617(.A0(new_n27053_), .A1(new_n26815_), .B0(new_n26813_), .Y(new_n27054_));
  AND2X1   g24618(.A(new_n27054_), .B(new_n27052_), .Y(new_n27055_));
  AOI21X1  g24619(.A0(new_n26854_), .A1(new_n25188_), .B0(new_n26841_), .Y(new_n27056_));
  OR2X1    g24620(.A(new_n27056_), .B(new_n26903_), .Y(new_n27057_));
  NOR2X1   g24621(.A(new_n9446_), .B(new_n24849_), .Y(new_n27058_));
  AOI21X1  g24622(.A0(new_n27058_), .A1(new_n26837_), .B0(new_n24823_), .Y(new_n27059_));
  OAI21X1  g24623(.A0(new_n26856_), .A1(pi0214), .B0(new_n27059_), .Y(new_n27060_));
  AOI21X1  g24624(.A0(new_n26856_), .A1(new_n26827_), .B0(pi0219), .Y(new_n27061_));
  AOI21X1  g24625(.A0(new_n27061_), .A1(new_n27060_), .B0(new_n27057_), .Y(new_n27062_));
  OR3X1    g24626(.A(new_n27062_), .B(new_n26008_), .C(new_n26280_), .Y(new_n27063_));
  AND2X1   g24627(.A(new_n26825_), .B(new_n24823_), .Y(new_n27064_));
  OR2X1    g24628(.A(new_n27064_), .B(pi0219), .Y(new_n27065_));
  AOI21X1  g24629(.A0(new_n27059_), .A1(new_n26826_), .B0(new_n27065_), .Y(new_n27066_));
  OR3X1    g24630(.A(new_n27066_), .B(new_n27056_), .C(new_n26903_), .Y(new_n27067_));
  OR3X1    g24631(.A(new_n26803_), .B(new_n26868_), .C(pi0219), .Y(new_n27068_));
  OR2X1    g24632(.A(new_n25819_), .B(pi1150), .Y(new_n27069_));
  AOI21X1  g24633(.A0(new_n27068_), .A1(new_n27052_), .B0(new_n27069_), .Y(new_n27070_));
  AOI21X1  g24634(.A0(new_n27070_), .A1(new_n27067_), .B0(pi1149), .Y(new_n27071_));
  OAI21X1  g24635(.A0(new_n27063_), .A1(new_n27055_), .B0(new_n27071_), .Y(new_n27072_));
  AOI21X1  g24636(.A0(new_n26836_), .A1(new_n26835_), .B0(new_n27056_), .Y(new_n27073_));
  NOR2X1   g24637(.A(new_n25089_), .B(new_n5102_), .Y(new_n27074_));
  OR3X1    g24638(.A(new_n27074_), .B(new_n25993_), .C(pi0057), .Y(new_n27075_));
  AOI21X1  g24639(.A0(new_n27073_), .A1(new_n5102_), .B0(new_n27075_), .Y(new_n27076_));
  NAND2X1  g24640(.A(new_n25089_), .B(pi0057), .Y(new_n27077_));
  NOR4X1   g24641(.A(new_n26804_), .B(new_n25109_), .C(new_n24817_), .D(new_n5103_), .Y(new_n27078_));
  NOR3X1   g24642(.A(new_n27074_), .B(pi1147), .C(pi0057), .Y(new_n27079_));
  OAI21X1  g24643(.A0(new_n26910_), .A1(new_n25089_), .B0(new_n27079_), .Y(new_n27080_));
  OAI21X1  g24644(.A0(new_n27080_), .A1(new_n27078_), .B0(new_n27077_), .Y(new_n27081_));
  OAI21X1  g24645(.A0(new_n27081_), .A1(new_n27076_), .B0(pi1150), .Y(new_n27082_));
  NOR3X1   g24646(.A(new_n27020_), .B(new_n26803_), .C(new_n9446_), .Y(new_n27083_));
  AOI21X1  g24647(.A0(new_n27083_), .A1(new_n26880_), .B0(new_n24823_), .Y(new_n27084_));
  INVX1    g24648(.A(new_n26805_), .Y(new_n27085_));
  OAI21X1  g24649(.A0(new_n27053_), .A1(new_n27085_), .B0(new_n8422_), .Y(new_n27086_));
  OAI21X1  g24650(.A0(new_n27086_), .A1(new_n27084_), .B0(new_n27052_), .Y(new_n27087_));
  AND3X1   g24651(.A(new_n26385_), .B(new_n6489_), .C(pi1147), .Y(new_n27088_));
  OR2X1    g24652(.A(new_n26000_), .B(pi1150), .Y(new_n27089_));
  AOI21X1  g24653(.A0(new_n27088_), .A1(new_n27073_), .B0(new_n27089_), .Y(new_n27090_));
  AOI21X1  g24654(.A0(new_n27090_), .A1(new_n27087_), .B0(new_n25955_), .Y(new_n27091_));
  AOI21X1  g24655(.A0(new_n27091_), .A1(new_n27082_), .B0(new_n26084_), .Y(new_n27092_));
  AOI21X1  g24656(.A0(new_n27092_), .A1(new_n27072_), .B0(new_n24815_), .Y(new_n27093_));
  OAI21X1  g24657(.A0(new_n27050_), .A1(pi1148), .B0(new_n27093_), .Y(new_n27094_));
  AOI21X1  g24658(.A0(new_n26877_), .A1(new_n24815_), .B0(pi0209), .Y(new_n27095_));
  AOI22X1  g24659(.A0(new_n27095_), .A1(new_n27094_), .B0(new_n27019_), .B1(new_n26935_), .Y(new_n27096_));
  MX2X1    g24660(.A(new_n27096_), .B(pi0246), .S0(new_n24814_), .Y(po0403));
  NAND2X1  g24661(.A(new_n26339_), .B(new_n25993_), .Y(new_n27098_));
  INVX1    g24662(.A(new_n25941_), .Y(new_n27099_));
  NOR2X1   g24663(.A(new_n25968_), .B(new_n25694_), .Y(new_n27100_));
  INVX1    g24664(.A(new_n27100_), .Y(new_n27101_));
  AOI21X1  g24665(.A0(new_n26986_), .A1(new_n27099_), .B0(new_n27101_), .Y(new_n27102_));
  OR2X1    g24666(.A(new_n26000_), .B(new_n25694_), .Y(new_n27103_));
  AOI21X1  g24667(.A0(new_n26985_), .A1(new_n26984_), .B0(new_n26402_), .Y(new_n27104_));
  NOR2X1   g24668(.A(new_n27104_), .B(new_n27103_), .Y(new_n27105_));
  INVX1    g24669(.A(new_n27105_), .Y(new_n27106_));
  OAI21X1  g24670(.A0(new_n25986_), .A1(new_n25974_), .B0(new_n26974_), .Y(new_n27107_));
  NAND3X1  g24671(.A(new_n27107_), .B(new_n26001_), .C(new_n25694_), .Y(new_n27108_));
  NAND3X1  g24672(.A(new_n27108_), .B(new_n27106_), .C(pi1147), .Y(new_n27109_));
  AND2X1   g24673(.A(new_n27109_), .B(new_n25955_), .Y(new_n27110_));
  OAI21X1  g24674(.A0(new_n27102_), .A1(new_n27098_), .B0(new_n27110_), .Y(new_n27111_));
  OR3X1    g24675(.A(new_n27001_), .B(new_n26048_), .C(pi0219), .Y(new_n27112_));
  AND2X1   g24676(.A(new_n27112_), .B(new_n26388_), .Y(new_n27113_));
  NAND2X1  g24677(.A(new_n26042_), .B(new_n8422_), .Y(new_n27114_));
  AND2X1   g24678(.A(new_n26388_), .B(new_n27114_), .Y(new_n27115_));
  NOR4X1   g24679(.A(new_n27115_), .B(new_n27113_), .C(new_n25804_), .D(pi1151), .Y(new_n27116_));
  OAI21X1  g24680(.A0(new_n27012_), .A1(new_n26263_), .B0(new_n25993_), .Y(new_n27117_));
  NOR2X1   g24681(.A(new_n26346_), .B(new_n25993_), .Y(new_n27118_));
  OR4X1    g24682(.A(new_n25998_), .B(new_n25961_), .C(new_n25958_), .D(pi1151), .Y(new_n27119_));
  AOI21X1  g24683(.A0(new_n27119_), .A1(new_n27118_), .B0(new_n25955_), .Y(new_n27120_));
  OAI21X1  g24684(.A0(new_n27117_), .A1(new_n27116_), .B0(new_n27120_), .Y(new_n27121_));
  NAND3X1  g24685(.A(new_n27121_), .B(new_n27111_), .C(pi1150), .Y(new_n27122_));
  OAI21X1  g24686(.A0(new_n25680_), .A1(new_n24823_), .B0(new_n26952_), .Y(new_n27123_));
  NAND2X1  g24687(.A(new_n27123_), .B(new_n26022_), .Y(new_n27124_));
  AOI21X1  g24688(.A0(new_n27124_), .A1(new_n26318_), .B0(new_n25993_), .Y(new_n27125_));
  AND2X1   g24689(.A(new_n26056_), .B(new_n26035_), .Y(new_n27126_));
  OAI21X1  g24690(.A0(new_n26038_), .A1(new_n25737_), .B0(new_n24824_), .Y(new_n27127_));
  AND3X1   g24691(.A(new_n27127_), .B(new_n26369_), .C(new_n26035_), .Y(new_n27128_));
  NOR4X1   g24692(.A(new_n27128_), .B(new_n27126_), .C(new_n25958_), .D(pi1151), .Y(new_n27129_));
  INVX1    g24693(.A(new_n27129_), .Y(new_n27130_));
  AOI21X1  g24694(.A0(new_n26952_), .A1(new_n26275_), .B0(new_n26103_), .Y(new_n27131_));
  NOR3X1   g24695(.A(new_n27131_), .B(new_n25804_), .C(new_n25694_), .Y(new_n27132_));
  NOR3X1   g24696(.A(new_n27128_), .B(new_n25804_), .C(pi1151), .Y(new_n27133_));
  OR2X1    g24697(.A(new_n27133_), .B(pi1147), .Y(new_n27134_));
  OAI21X1  g24698(.A0(new_n27134_), .A1(new_n27132_), .B0(pi1149), .Y(new_n27135_));
  AOI21X1  g24699(.A0(new_n27130_), .A1(new_n27125_), .B0(new_n27135_), .Y(new_n27136_));
  NOR3X1   g24700(.A(new_n25967_), .B(new_n11660_), .C(pi0219), .Y(new_n27137_));
  OR2X1    g24701(.A(new_n27137_), .B(pi1151), .Y(new_n27138_));
  AND2X1   g24702(.A(new_n27138_), .B(new_n25993_), .Y(new_n27139_));
  INVX1    g24703(.A(new_n25847_), .Y(new_n27140_));
  NOR2X1   g24704(.A(new_n26288_), .B(new_n27140_), .Y(new_n27141_));
  OAI21X1  g24705(.A0(new_n27141_), .A1(new_n27101_), .B0(new_n27139_), .Y(new_n27142_));
  AND3X1   g24706(.A(new_n26430_), .B(new_n26001_), .C(pi1151), .Y(new_n27143_));
  AND2X1   g24707(.A(new_n26323_), .B(new_n25997_), .Y(new_n27144_));
  OR3X1    g24708(.A(new_n27144_), .B(new_n27143_), .C(new_n25993_), .Y(new_n27145_));
  AND3X1   g24709(.A(new_n27145_), .B(new_n27142_), .C(new_n25955_), .Y(new_n27146_));
  OR3X1    g24710(.A(new_n27146_), .B(new_n27136_), .C(pi1150), .Y(new_n27147_));
  AOI21X1  g24711(.A0(new_n27147_), .A1(new_n27122_), .B0(new_n26084_), .Y(new_n27148_));
  AOI21X1  g24712(.A0(new_n26301_), .A1(new_n26024_), .B0(new_n25993_), .Y(new_n27149_));
  NOR2X1   g24713(.A(new_n26008_), .B(pi1151), .Y(new_n27150_));
  INVX1    g24714(.A(new_n27150_), .Y(new_n27151_));
  OAI21X1  g24715(.A0(new_n27151_), .A1(new_n27126_), .B0(new_n27149_), .Y(new_n27152_));
  INVX1    g24716(.A(new_n26071_), .Y(new_n27153_));
  NOR3X1   g24717(.A(new_n26018_), .B(new_n26015_), .C(pi0219), .Y(new_n27154_));
  OR2X1    g24718(.A(new_n26103_), .B(new_n27154_), .Y(new_n27155_));
  AND3X1   g24719(.A(new_n27155_), .B(new_n27153_), .C(pi1151), .Y(new_n27156_));
  AOI21X1  g24720(.A0(new_n26070_), .A1(po1038), .B0(pi1151), .Y(new_n27157_));
  AND2X1   g24721(.A(new_n27157_), .B(new_n26358_), .Y(new_n27158_));
  OR3X1    g24722(.A(new_n27158_), .B(new_n27156_), .C(pi1147), .Y(new_n27159_));
  AND3X1   g24723(.A(new_n27159_), .B(new_n27152_), .C(new_n26280_), .Y(new_n27160_));
  AOI21X1  g24724(.A0(new_n26376_), .A1(new_n26301_), .B0(new_n25993_), .Y(new_n27161_));
  OR3X1    g24725(.A(new_n26056_), .B(new_n26008_), .C(pi1151), .Y(new_n27162_));
  NOR3X1   g24726(.A(new_n27113_), .B(new_n26071_), .C(pi1151), .Y(new_n27163_));
  NOR3X1   g24727(.A(new_n26145_), .B(new_n26071_), .C(new_n25694_), .Y(new_n27164_));
  OR3X1    g24728(.A(new_n27164_), .B(new_n27163_), .C(pi1147), .Y(new_n27165_));
  NAND2X1  g24729(.A(new_n27165_), .B(pi1150), .Y(new_n27166_));
  AOI21X1  g24730(.A0(new_n27162_), .A1(new_n27161_), .B0(new_n27166_), .Y(new_n27167_));
  OAI21X1  g24731(.A0(new_n27167_), .A1(new_n27160_), .B0(pi1149), .Y(new_n27168_));
  INVX1    g24732(.A(new_n25820_), .Y(new_n27169_));
  OR2X1    g24733(.A(new_n26993_), .B(new_n26992_), .Y(new_n27170_));
  AOI21X1  g24734(.A0(new_n27104_), .A1(new_n27170_), .B0(new_n27169_), .Y(new_n27171_));
  NOR3X1   g24735(.A(new_n26978_), .B(new_n25819_), .C(pi1151), .Y(new_n27172_));
  NOR3X1   g24736(.A(new_n27172_), .B(new_n27171_), .C(new_n25993_), .Y(new_n27173_));
  OAI21X1  g24737(.A0(new_n26085_), .A1(pi1151), .B0(new_n25993_), .Y(new_n27174_));
  AND2X1   g24738(.A(new_n26982_), .B(pi1151), .Y(new_n27175_));
  OAI21X1  g24739(.A0(new_n27175_), .A1(new_n27174_), .B0(pi1150), .Y(new_n27176_));
  OAI21X1  g24740(.A0(new_n26375_), .A1(new_n25843_), .B0(new_n26428_), .Y(new_n27177_));
  AOI21X1  g24741(.A0(new_n26375_), .A1(new_n26054_), .B0(new_n26312_), .Y(new_n27178_));
  OR2X1    g24742(.A(new_n27178_), .B(new_n25993_), .Y(new_n27179_));
  AOI21X1  g24743(.A0(new_n27177_), .A1(new_n25820_), .B0(new_n27179_), .Y(new_n27180_));
  INVX1    g24744(.A(new_n26026_), .Y(new_n27181_));
  OR2X1    g24745(.A(new_n25694_), .B(pi1147), .Y(new_n27182_));
  OAI21X1  g24746(.A0(new_n27182_), .A1(new_n27181_), .B0(new_n26280_), .Y(new_n27183_));
  OAI22X1  g24747(.A0(new_n27183_), .A1(new_n27180_), .B0(new_n27176_), .B1(new_n27173_), .Y(new_n27184_));
  AOI21X1  g24748(.A0(new_n27184_), .A1(new_n25955_), .B0(pi1148), .Y(new_n27185_));
  AOI21X1  g24749(.A0(new_n27185_), .A1(new_n27168_), .B0(new_n27148_), .Y(new_n27186_));
  NAND3X1  g24750(.A(new_n26350_), .B(new_n26343_), .C(pi0213), .Y(new_n27187_));
  AND2X1   g24751(.A(new_n27187_), .B(pi0209), .Y(new_n27188_));
  OAI21X1  g24752(.A0(new_n27186_), .A1(pi0213), .B0(new_n27188_), .Y(new_n27189_));
  NOR3X1   g24753(.A(new_n27113_), .B(new_n26071_), .C(new_n25694_), .Y(new_n27190_));
  NOR3X1   g24754(.A(new_n27190_), .B(new_n26381_), .C(new_n25993_), .Y(new_n27191_));
  AOI21X1  g24755(.A0(new_n25971_), .A1(new_n25799_), .B0(po1038), .Y(new_n27192_));
  OAI21X1  g24756(.A0(new_n25980_), .A1(new_n25799_), .B0(new_n27192_), .Y(new_n27193_));
  AND2X1   g24757(.A(new_n27193_), .B(new_n26251_), .Y(new_n27194_));
  INVX1    g24758(.A(new_n27194_), .Y(new_n27195_));
  OAI21X1  g24759(.A0(new_n27195_), .A1(new_n27174_), .B0(new_n26280_), .Y(new_n27196_));
  AOI21X1  g24760(.A0(new_n25989_), .A1(new_n25984_), .B0(new_n26263_), .Y(new_n27197_));
  INVX1    g24761(.A(new_n27197_), .Y(new_n27198_));
  AND3X1   g24762(.A(new_n27198_), .B(new_n26339_), .C(new_n25993_), .Y(new_n27199_));
  NOR3X1   g24763(.A(new_n27115_), .B(new_n27113_), .C(new_n26263_), .Y(new_n27200_));
  INVX1    g24764(.A(new_n26281_), .Y(new_n27201_));
  OAI21X1  g24765(.A0(new_n27115_), .A1(new_n27201_), .B0(pi1147), .Y(new_n27202_));
  OAI21X1  g24766(.A0(new_n27202_), .A1(new_n27200_), .B0(pi1150), .Y(new_n27203_));
  OAI22X1  g24767(.A0(new_n27203_), .A1(new_n27199_), .B0(new_n27196_), .B1(new_n27191_), .Y(new_n27204_));
  AOI21X1  g24768(.A0(new_n27104_), .A1(new_n27170_), .B0(new_n26312_), .Y(new_n27205_));
  AND3X1   g24769(.A(new_n26994_), .B(new_n26009_), .C(pi1151), .Y(new_n27206_));
  OR2X1    g24770(.A(new_n27206_), .B(pi1147), .Y(new_n27207_));
  OAI21X1  g24771(.A0(new_n26133_), .A1(po1038), .B0(new_n27178_), .Y(new_n27208_));
  AOI21X1  g24772(.A0(new_n27208_), .A1(new_n27161_), .B0(pi1150), .Y(new_n27209_));
  OAI21X1  g24773(.A0(new_n27207_), .A1(new_n27205_), .B0(new_n27209_), .Y(new_n27210_));
  AOI21X1  g24774(.A0(new_n25944_), .A1(pi0212), .B0(new_n25948_), .Y(new_n27211_));
  OAI21X1  g24775(.A0(new_n27211_), .A1(new_n26402_), .B0(new_n26318_), .Y(new_n27212_));
  AND2X1   g24776(.A(new_n27212_), .B(new_n25993_), .Y(new_n27213_));
  OAI21X1  g24777(.A0(new_n27104_), .A1(new_n26324_), .B0(new_n27213_), .Y(new_n27214_));
  AOI21X1  g24778(.A0(new_n26385_), .A1(new_n26384_), .B0(new_n26000_), .Y(new_n27215_));
  NAND2X1  g24779(.A(new_n27215_), .B(new_n25694_), .Y(new_n27216_));
  AOI21X1  g24780(.A0(new_n27216_), .A1(new_n27118_), .B0(new_n26280_), .Y(new_n27217_));
  NAND2X1  g24781(.A(new_n27217_), .B(new_n27214_), .Y(new_n27218_));
  AOI21X1  g24782(.A0(new_n27218_), .A1(new_n27210_), .B0(new_n25955_), .Y(new_n27219_));
  OR2X1    g24783(.A(new_n27219_), .B(new_n26084_), .Y(new_n27220_));
  AOI21X1  g24784(.A0(new_n27204_), .A1(new_n25955_), .B0(new_n27220_), .Y(new_n27221_));
  OR2X1    g24785(.A(new_n26287_), .B(pi0219), .Y(new_n27222_));
  OAI21X1  g24786(.A0(new_n27222_), .A1(new_n26363_), .B0(new_n26022_), .Y(new_n27223_));
  OAI21X1  g24787(.A0(new_n27223_), .A1(new_n26019_), .B0(new_n26311_), .Y(new_n27224_));
  NAND2X1  g24788(.A(new_n25847_), .B(new_n26426_), .Y(new_n27225_));
  OAI21X1  g24789(.A0(new_n27225_), .A1(new_n7996_), .B0(new_n27177_), .Y(new_n27226_));
  NOR3X1   g24790(.A(new_n27226_), .B(new_n26008_), .C(new_n25694_), .Y(new_n27227_));
  AND2X1   g24791(.A(new_n27177_), .B(new_n26311_), .Y(new_n27228_));
  OR2X1    g24792(.A(new_n27228_), .B(pi1147), .Y(new_n27229_));
  OAI21X1  g24793(.A0(new_n27229_), .A1(new_n27227_), .B0(new_n26280_), .Y(new_n27230_));
  AOI21X1  g24794(.A0(new_n27224_), .A1(new_n27149_), .B0(new_n27230_), .Y(new_n27231_));
  NAND3X1  g24795(.A(new_n27223_), .B(new_n26001_), .C(new_n25694_), .Y(new_n27232_));
  AND3X1   g24796(.A(new_n27225_), .B(new_n26430_), .C(new_n26318_), .Y(new_n27233_));
  AND2X1   g24797(.A(new_n26430_), .B(new_n26323_), .Y(new_n27234_));
  NOR3X1   g24798(.A(new_n27234_), .B(new_n27233_), .C(pi1147), .Y(new_n27235_));
  OR2X1    g24799(.A(new_n27235_), .B(new_n26280_), .Y(new_n27236_));
  AOI21X1  g24800(.A0(new_n27232_), .A1(new_n27125_), .B0(new_n27236_), .Y(new_n27237_));
  OAI21X1  g24801(.A0(new_n27237_), .A1(new_n27231_), .B0(pi1149), .Y(new_n27238_));
  AOI21X1  g24802(.A0(new_n26369_), .A1(new_n26043_), .B0(new_n25968_), .Y(new_n27239_));
  OAI21X1  g24803(.A0(new_n27128_), .A1(new_n26263_), .B0(pi1147), .Y(new_n27240_));
  AOI21X1  g24804(.A0(new_n27239_), .A1(new_n25694_), .B0(new_n27240_), .Y(new_n27241_));
  INVX1    g24805(.A(new_n27139_), .Y(new_n27242_));
  AOI21X1  g24806(.A0(new_n26432_), .A1(new_n22572_), .B0(new_n25694_), .Y(new_n27243_));
  OAI21X1  g24807(.A0(new_n27243_), .A1(new_n27242_), .B0(pi1150), .Y(new_n27244_));
  OAI21X1  g24808(.A0(new_n26939_), .A1(pi1151), .B0(pi1147), .Y(new_n27245_));
  AOI21X1  g24809(.A0(new_n26358_), .A1(new_n27153_), .B0(new_n27245_), .Y(new_n27246_));
  OR4X1    g24810(.A(new_n25086_), .B(new_n11660_), .C(pi0219), .D(pi0211), .Y(new_n27247_));
  OAI21X1  g24811(.A0(new_n27182_), .A1(new_n27247_), .B0(new_n26280_), .Y(new_n27248_));
  OAI22X1  g24812(.A0(new_n27248_), .A1(new_n27246_), .B0(new_n27244_), .B1(new_n27241_), .Y(new_n27249_));
  AOI21X1  g24813(.A0(new_n27249_), .A1(new_n25955_), .B0(pi1148), .Y(new_n27250_));
  AOI21X1  g24814(.A0(new_n27250_), .A1(new_n27238_), .B0(new_n27221_), .Y(new_n27251_));
  AOI21X1  g24815(.A0(new_n26061_), .A1(new_n24815_), .B0(pi0209), .Y(new_n27252_));
  OAI21X1  g24816(.A0(new_n27251_), .A1(new_n24815_), .B0(new_n27252_), .Y(new_n27253_));
  AND2X1   g24817(.A(new_n27253_), .B(new_n27189_), .Y(new_n27254_));
  MX2X1    g24818(.A(new_n27254_), .B(pi0247), .S0(new_n24814_), .Y(po0404));
  OR3X1    g24819(.A(new_n27234_), .B(new_n27105_), .C(new_n25153_), .Y(new_n27256_));
  NAND3X1  g24820(.A(new_n27107_), .B(new_n26001_), .C(pi1151), .Y(new_n27257_));
  AOI21X1  g24821(.A0(new_n26323_), .A1(new_n25997_), .B0(pi1152), .Y(new_n27258_));
  AOI21X1  g24822(.A0(new_n27258_), .A1(new_n27257_), .B0(pi1150), .Y(new_n27259_));
  AND2X1   g24823(.A(new_n27259_), .B(new_n27256_), .Y(new_n27260_));
  NOR2X1   g24824(.A(new_n25958_), .B(pi1151), .Y(new_n27261_));
  OR2X1    g24825(.A(new_n26346_), .B(new_n25153_), .Y(new_n27262_));
  AOI21X1  g24826(.A0(new_n27261_), .A1(new_n27124_), .B0(new_n27262_), .Y(new_n27263_));
  NOR4X1   g24827(.A(new_n25998_), .B(new_n25961_), .C(new_n25958_), .D(new_n25694_), .Y(new_n27264_));
  OR2X1    g24828(.A(new_n27264_), .B(pi1152), .Y(new_n27265_));
  OAI21X1  g24829(.A0(new_n27265_), .A1(new_n27129_), .B0(pi1150), .Y(new_n27266_));
  OAI21X1  g24830(.A0(new_n27266_), .A1(new_n27263_), .B0(pi1148), .Y(new_n27267_));
  INVX1    g24831(.A(new_n27137_), .Y(new_n27268_));
  OAI21X1  g24832(.A0(new_n27101_), .A1(new_n25991_), .B0(new_n25153_), .Y(new_n27269_));
  AOI21X1  g24833(.A0(new_n27268_), .A1(new_n25694_), .B0(new_n27269_), .Y(new_n27270_));
  OAI21X1  g24834(.A0(new_n27141_), .A1(new_n27201_), .B0(pi1152), .Y(new_n27271_));
  OAI21X1  g24835(.A0(new_n27271_), .A1(new_n27102_), .B0(new_n26280_), .Y(new_n27272_));
  NOR2X1   g24836(.A(new_n27272_), .B(new_n27270_), .Y(new_n27273_));
  NOR3X1   g24837(.A(new_n27131_), .B(new_n25804_), .C(pi1151), .Y(new_n27274_));
  OAI21X1  g24838(.A0(new_n27012_), .A1(new_n26263_), .B0(pi1152), .Y(new_n27275_));
  NOR2X1   g24839(.A(new_n27275_), .B(new_n27274_), .Y(new_n27276_));
  NOR3X1   g24840(.A(new_n27200_), .B(new_n27133_), .C(pi1152), .Y(new_n27277_));
  OR2X1    g24841(.A(new_n27277_), .B(new_n26280_), .Y(new_n27278_));
  OAI21X1  g24842(.A0(new_n27278_), .A1(new_n27276_), .B0(new_n26084_), .Y(new_n27279_));
  OAI22X1  g24843(.A0(new_n27279_), .A1(new_n27273_), .B0(new_n27267_), .B1(new_n27260_), .Y(new_n27280_));
  NAND2X1  g24844(.A(new_n26376_), .B(new_n26301_), .Y(new_n27281_));
  OAI21X1  g24845(.A0(new_n26023_), .A1(new_n26019_), .B0(new_n27150_), .Y(new_n27282_));
  AND2X1   g24846(.A(new_n27282_), .B(pi1152), .Y(new_n27283_));
  AOI21X1  g24847(.A0(new_n26056_), .A1(new_n26035_), .B0(new_n27151_), .Y(new_n27284_));
  NOR3X1   g24848(.A(new_n26056_), .B(new_n26008_), .C(new_n25694_), .Y(new_n27285_));
  NOR3X1   g24849(.A(new_n27285_), .B(new_n27284_), .C(pi1152), .Y(new_n27286_));
  AOI21X1  g24850(.A0(new_n27283_), .A1(new_n27281_), .B0(new_n27286_), .Y(new_n27287_));
  OAI21X1  g24851(.A0(new_n27228_), .A1(new_n27171_), .B0(pi1152), .Y(new_n27288_));
  NOR3X1   g24852(.A(new_n26978_), .B(new_n25819_), .C(new_n25694_), .Y(new_n27289_));
  OAI21X1  g24853(.A0(new_n27289_), .A1(new_n27178_), .B0(new_n25153_), .Y(new_n27290_));
  NAND3X1  g24854(.A(new_n27290_), .B(new_n27288_), .C(new_n26280_), .Y(new_n27291_));
  AND2X1   g24855(.A(new_n27291_), .B(pi1148), .Y(new_n27292_));
  OAI21X1  g24856(.A0(new_n27287_), .A1(new_n26280_), .B0(new_n27292_), .Y(new_n27293_));
  AND3X1   g24857(.A(new_n27155_), .B(new_n27153_), .C(new_n25694_), .Y(new_n27294_));
  NOR3X1   g24858(.A(new_n27294_), .B(new_n27164_), .C(new_n25153_), .Y(new_n27295_));
  NOR3X1   g24859(.A(new_n27190_), .B(new_n27158_), .C(pi1152), .Y(new_n27296_));
  OR2X1    g24860(.A(new_n27296_), .B(new_n26280_), .Y(new_n27297_));
  AND2X1   g24861(.A(new_n25153_), .B(pi1151), .Y(new_n27298_));
  INVX1    g24862(.A(new_n27298_), .Y(new_n27299_));
  OR2X1    g24863(.A(new_n26026_), .B(pi1151), .Y(new_n27300_));
  AOI21X1  g24864(.A0(new_n26982_), .A1(pi1151), .B0(new_n25153_), .Y(new_n27301_));
  AOI21X1  g24865(.A0(new_n27301_), .A1(new_n27300_), .B0(pi1150), .Y(new_n27302_));
  OAI21X1  g24866(.A0(new_n27299_), .A1(new_n26086_), .B0(new_n27302_), .Y(new_n27303_));
  OAI21X1  g24867(.A0(new_n27297_), .A1(new_n27295_), .B0(new_n27303_), .Y(new_n27304_));
  AOI21X1  g24868(.A0(new_n27304_), .A1(new_n26084_), .B0(pi1149), .Y(new_n27305_));
  AOI22X1  g24869(.A0(new_n27305_), .A1(new_n27293_), .B0(new_n27280_), .B1(pi1149), .Y(new_n27306_));
  OR2X1    g24870(.A(new_n27306_), .B(pi0213), .Y(new_n27307_));
  OAI21X1  g24871(.A0(new_n25991_), .A1(new_n25968_), .B0(new_n27298_), .Y(new_n27308_));
  AND2X1   g24872(.A(new_n27247_), .B(new_n25694_), .Y(new_n27309_));
  AOI21X1  g24873(.A0(new_n27309_), .A1(new_n27181_), .B0(new_n25153_), .Y(new_n27310_));
  AOI21X1  g24874(.A0(new_n27310_), .A1(new_n26340_), .B0(pi1150), .Y(new_n27311_));
  NAND3X1  g24875(.A(new_n27282_), .B(new_n26347_), .C(pi1152), .Y(new_n27312_));
  AOI21X1  g24876(.A0(new_n26002_), .A1(pi1151), .B0(pi1152), .Y(new_n27313_));
  OAI21X1  g24877(.A0(new_n26312_), .A1(new_n26057_), .B0(new_n27313_), .Y(new_n27314_));
  AND2X1   g24878(.A(new_n27314_), .B(pi1150), .Y(new_n27315_));
  AOI22X1  g24879(.A0(new_n27315_), .A1(new_n27312_), .B0(new_n27311_), .B1(new_n27308_), .Y(new_n27316_));
  AOI21X1  g24880(.A0(new_n27316_), .A1(pi0213), .B0(new_n24866_), .Y(new_n27317_));
  NOR2X1   g24881(.A(new_n26085_), .B(pi1151), .Y(new_n27318_));
  AOI21X1  g24882(.A0(new_n27195_), .A1(new_n25694_), .B0(new_n25153_), .Y(new_n27319_));
  AOI21X1  g24883(.A0(new_n27319_), .A1(new_n27198_), .B0(pi1150), .Y(new_n27320_));
  OAI21X1  g24884(.A0(new_n27269_), .A1(new_n27318_), .B0(new_n27320_), .Y(new_n27321_));
  OR3X1    g24885(.A(new_n27205_), .B(new_n27105_), .C(pi1152), .Y(new_n27322_));
  NAND3X1  g24886(.A(new_n26994_), .B(new_n26009_), .C(new_n25694_), .Y(new_n27323_));
  AND2X1   g24887(.A(new_n27212_), .B(pi1152), .Y(new_n27324_));
  AOI21X1  g24888(.A0(new_n27324_), .A1(new_n27323_), .B0(new_n26280_), .Y(new_n27325_));
  AOI21X1  g24889(.A0(new_n27325_), .A1(new_n27322_), .B0(new_n25955_), .Y(new_n27326_));
  NOR2X1   g24890(.A(new_n27233_), .B(new_n25153_), .Y(new_n27327_));
  OAI21X1  g24891(.A0(new_n27226_), .A1(new_n27151_), .B0(new_n27327_), .Y(new_n27328_));
  OR3X1    g24892(.A(new_n27228_), .B(new_n27143_), .C(pi1152), .Y(new_n27329_));
  AND3X1   g24893(.A(new_n27329_), .B(new_n27328_), .C(pi1150), .Y(new_n27330_));
  NOR3X1   g24894(.A(new_n27309_), .B(new_n27243_), .C(new_n25153_), .Y(new_n27331_));
  OAI21X1  g24895(.A0(new_n27299_), .A1(new_n27268_), .B0(new_n26280_), .Y(new_n27332_));
  OAI21X1  g24896(.A0(new_n27332_), .A1(new_n27331_), .B0(new_n25955_), .Y(new_n27333_));
  OAI21X1  g24897(.A0(new_n27333_), .A1(new_n27330_), .B0(new_n26084_), .Y(new_n27334_));
  AOI21X1  g24898(.A0(new_n27326_), .A1(new_n27321_), .B0(new_n27334_), .Y(new_n27335_));
  NAND2X1  g24899(.A(new_n27124_), .B(new_n26318_), .Y(new_n27336_));
  AND3X1   g24900(.A(new_n27282_), .B(new_n27336_), .C(pi1152), .Y(new_n27337_));
  NAND3X1  g24901(.A(new_n27223_), .B(new_n26001_), .C(pi1151), .Y(new_n27338_));
  AND3X1   g24902(.A(new_n27338_), .B(new_n27224_), .C(new_n25153_), .Y(new_n27339_));
  OR3X1    g24903(.A(new_n27339_), .B(new_n27337_), .C(new_n26280_), .Y(new_n27340_));
  AND2X1   g24904(.A(new_n27239_), .B(pi1151), .Y(new_n27341_));
  OAI21X1  g24905(.A0(new_n26939_), .A1(pi1151), .B0(new_n25153_), .Y(new_n27342_));
  OR2X1    g24906(.A(new_n27342_), .B(new_n27341_), .Y(new_n27343_));
  AOI21X1  g24907(.A0(new_n27157_), .A1(new_n26358_), .B0(new_n25153_), .Y(new_n27344_));
  OAI21X1  g24908(.A0(new_n27128_), .A1(new_n26263_), .B0(new_n27344_), .Y(new_n27345_));
  AND2X1   g24909(.A(new_n27345_), .B(new_n26280_), .Y(new_n27346_));
  AOI21X1  g24910(.A0(new_n27346_), .A1(new_n27343_), .B0(pi1149), .Y(new_n27347_));
  NOR3X1   g24911(.A(new_n27200_), .B(new_n27163_), .C(new_n25153_), .Y(new_n27348_));
  INVX1    g24912(.A(new_n26382_), .Y(new_n27349_));
  AOI21X1  g24913(.A0(new_n26388_), .A1(new_n27114_), .B0(new_n27101_), .Y(new_n27350_));
  OAI21X1  g24914(.A0(new_n27350_), .A1(new_n27349_), .B0(new_n26280_), .Y(new_n27351_));
  NOR2X1   g24915(.A(new_n27351_), .B(new_n27348_), .Y(new_n27352_));
  AOI21X1  g24916(.A0(new_n27150_), .A1(new_n26376_), .B0(new_n27262_), .Y(new_n27353_));
  AND2X1   g24917(.A(new_n27215_), .B(pi1151), .Y(new_n27354_));
  NAND2X1  g24918(.A(new_n27208_), .B(new_n25153_), .Y(new_n27355_));
  OAI21X1  g24919(.A0(new_n27355_), .A1(new_n27354_), .B0(pi1150), .Y(new_n27356_));
  OAI21X1  g24920(.A0(new_n27356_), .A1(new_n27353_), .B0(pi1149), .Y(new_n27357_));
  OAI21X1  g24921(.A0(new_n27357_), .A1(new_n27352_), .B0(pi1148), .Y(new_n27358_));
  AOI21X1  g24922(.A0(new_n27347_), .A1(new_n27340_), .B0(new_n27358_), .Y(new_n27359_));
  OR3X1    g24923(.A(new_n27359_), .B(new_n27335_), .C(new_n24815_), .Y(new_n27360_));
  AOI21X1  g24924(.A0(new_n26934_), .A1(new_n24815_), .B0(pi0209), .Y(new_n27361_));
  AOI22X1  g24925(.A0(new_n27361_), .A1(new_n27360_), .B0(new_n27317_), .B1(new_n27307_), .Y(new_n27362_));
  MX2X1    g24926(.A(new_n27362_), .B(pi0248), .S0(new_n24814_), .Y(po0405));
  NAND2X1  g24927(.A(new_n27316_), .B(new_n24815_), .Y(new_n27364_));
  AND2X1   g24928(.A(new_n25111_), .B(pi0299), .Y(new_n27365_));
  NOR3X1   g24929(.A(new_n27365_), .B(new_n26034_), .C(new_n25737_), .Y(new_n27366_));
  NOR3X1   g24930(.A(new_n27365_), .B(new_n26034_), .C(pi0214), .Y(new_n27367_));
  NOR2X1   g24931(.A(new_n26033_), .B(new_n25833_), .Y(new_n27368_));
  OR2X1    g24932(.A(new_n26357_), .B(new_n24849_), .Y(new_n27369_));
  OAI21X1  g24933(.A0(new_n27369_), .A1(new_n27368_), .B0(pi0212), .Y(new_n27370_));
  OAI22X1  g24934(.A0(new_n27370_), .A1(new_n27367_), .B0(new_n27366_), .B1(pi0212), .Y(new_n27371_));
  OAI21X1  g24935(.A0(new_n26033_), .A1(new_n8422_), .B0(new_n5102_), .Y(new_n27372_));
  AOI21X1  g24936(.A0(new_n27371_), .A1(new_n8422_), .B0(new_n27372_), .Y(new_n27373_));
  NOR4X1   g24937(.A(new_n25112_), .B(new_n25110_), .C(new_n24879_), .D(new_n5102_), .Y(new_n27374_));
  OR4X1    g24938(.A(new_n27374_), .B(new_n27373_), .C(pi1151), .D(pi0057), .Y(new_n27375_));
  NOR2X1   g24939(.A(new_n25113_), .B(new_n2436_), .Y(new_n27376_));
  OR2X1    g24940(.A(new_n27365_), .B(new_n26390_), .Y(new_n27377_));
  OAI21X1  g24941(.A0(new_n25859_), .A1(new_n25723_), .B0(pi0212), .Y(new_n27378_));
  AOI21X1  g24942(.A0(new_n27377_), .A1(new_n24849_), .B0(new_n27378_), .Y(new_n27379_));
  OR2X1    g24943(.A(new_n25737_), .B(pi0212), .Y(new_n27380_));
  AOI21X1  g24944(.A0(new_n27377_), .A1(pi0214), .B0(new_n27380_), .Y(new_n27381_));
  OR3X1    g24945(.A(new_n27381_), .B(new_n27379_), .C(pi0219), .Y(new_n27382_));
  NAND3X1  g24946(.A(new_n27382_), .B(new_n25741_), .C(new_n5102_), .Y(new_n27383_));
  NOR3X1   g24947(.A(new_n27374_), .B(new_n25694_), .C(pi0057), .Y(new_n27384_));
  AOI21X1  g24948(.A0(new_n27384_), .A1(new_n27383_), .B0(new_n27376_), .Y(new_n27385_));
  AOI21X1  g24949(.A0(new_n27385_), .A1(new_n27375_), .B0(pi1152), .Y(new_n27386_));
  NAND2X1  g24950(.A(new_n26353_), .B(new_n26011_), .Y(new_n27387_));
  OAI21X1  g24951(.A0(new_n27365_), .A1(new_n25680_), .B0(new_n24849_), .Y(new_n27388_));
  AND3X1   g24952(.A(new_n27388_), .B(new_n27387_), .C(pi0212), .Y(new_n27389_));
  NOR4X1   g24953(.A(new_n27365_), .B(new_n25696_), .C(new_n25688_), .D(pi0212), .Y(new_n27390_));
  OR3X1    g24954(.A(new_n27390_), .B(new_n27389_), .C(new_n26951_), .Y(new_n27391_));
  AND3X1   g24955(.A(new_n27391_), .B(new_n26022_), .C(new_n25694_), .Y(new_n27392_));
  OR2X1    g24956(.A(new_n25962_), .B(pi0219), .Y(new_n27393_));
  OR3X1    g24957(.A(new_n25111_), .B(new_n7996_), .C(new_n2933_), .Y(new_n27394_));
  OAI21X1  g24958(.A0(new_n25155_), .A1(new_n24823_), .B0(new_n27394_), .Y(new_n27395_));
  AOI21X1  g24959(.A0(new_n27395_), .A1(new_n25959_), .B0(new_n27393_), .Y(new_n27396_));
  OAI21X1  g24960(.A0(new_n26134_), .A1(new_n26054_), .B0(pi1151), .Y(new_n27397_));
  OAI21X1  g24961(.A0(new_n27397_), .A1(new_n27396_), .B0(new_n25159_), .Y(new_n27398_));
  OAI21X1  g24962(.A0(new_n27398_), .A1(new_n27392_), .B0(pi1150), .Y(new_n27399_));
  OR3X1    g24963(.A(new_n25978_), .B(new_n25224_), .C(pi0211), .Y(new_n27400_));
  OR3X1    g24964(.A(new_n25978_), .B(new_n25001_), .C(new_n23173_), .Y(new_n27401_));
  AND3X1   g24965(.A(new_n27401_), .B(new_n27400_), .C(new_n25085_), .Y(new_n27402_));
  INVX1    g24966(.A(new_n25283_), .Y(new_n27403_));
  OAI22X1  g24967(.A0(new_n26413_), .A1(new_n24877_), .B0(new_n25971_), .B1(new_n27403_), .Y(new_n27404_));
  OAI21X1  g24968(.A0(new_n27404_), .A1(new_n27402_), .B0(new_n8422_), .Y(new_n27405_));
  AND3X1   g24969(.A(new_n25988_), .B(new_n6489_), .C(pi1151), .Y(new_n27406_));
  NOR2X1   g24970(.A(new_n25111_), .B(new_n2933_), .Y(new_n27407_));
  AOI21X1  g24971(.A0(new_n27407_), .A1(new_n24877_), .B0(new_n25723_), .Y(new_n27408_));
  OR4X1    g24972(.A(new_n25112_), .B(new_n25110_), .C(po1038), .D(pi1151), .Y(new_n27409_));
  OAI21X1  g24973(.A0(new_n27409_), .A1(new_n27408_), .B0(new_n25114_), .Y(new_n27410_));
  AOI21X1  g24974(.A0(new_n27406_), .A1(new_n27405_), .B0(new_n27410_), .Y(new_n27411_));
  OAI21X1  g24975(.A0(new_n27407_), .A1(new_n25945_), .B0(pi0212), .Y(new_n27412_));
  AOI21X1  g24976(.A0(new_n26406_), .A1(pi0214), .B0(new_n27412_), .Y(new_n27413_));
  OAI21X1  g24977(.A0(new_n25721_), .A1(pi0212), .B0(new_n8422_), .Y(new_n27414_));
  OR3X1    g24978(.A(new_n27414_), .B(new_n27413_), .C(new_n27390_), .Y(new_n27415_));
  INVX1    g24979(.A(new_n25679_), .Y(new_n27416_));
  AOI21X1  g24980(.A0(new_n26122_), .A1(new_n26121_), .B0(new_n27416_), .Y(new_n27417_));
  OR2X1    g24981(.A(new_n27409_), .B(new_n27408_), .Y(new_n27418_));
  AND2X1   g24982(.A(new_n27418_), .B(new_n25159_), .Y(new_n27419_));
  OAI21X1  g24983(.A0(new_n27177_), .A1(pi1151), .B0(new_n27419_), .Y(new_n27420_));
  AOI21X1  g24984(.A0(new_n27417_), .A1(new_n27415_), .B0(new_n27420_), .Y(new_n27421_));
  OR3X1    g24985(.A(new_n27421_), .B(new_n27411_), .C(pi1150), .Y(new_n27422_));
  OAI21X1  g24986(.A0(new_n27399_), .A1(new_n27386_), .B0(new_n27422_), .Y(new_n27423_));
  AOI21X1  g24987(.A0(new_n27423_), .A1(pi0213), .B0(pi0209), .Y(new_n27424_));
  AND3X1   g24988(.A(new_n25290_), .B(new_n25265_), .C(new_n22660_), .Y(new_n27425_));
  OR3X1    g24989(.A(new_n25279_), .B(new_n25001_), .C(new_n22660_), .Y(new_n27426_));
  AND2X1   g24990(.A(new_n27426_), .B(pi0208), .Y(new_n27427_));
  INVX1    g24991(.A(new_n27427_), .Y(new_n27428_));
  OAI22X1  g24992(.A0(new_n27428_), .A1(new_n27425_), .B0(new_n25389_), .B1(new_n24986_), .Y(new_n27429_));
  AND3X1   g24993(.A(new_n27429_), .B(pi0214), .C(pi0211), .Y(new_n27430_));
  AOI21X1  g24994(.A0(new_n25281_), .A1(new_n25033_), .B0(new_n27430_), .Y(new_n27431_));
  OAI21X1  g24995(.A0(new_n27431_), .A1(pi0212), .B0(new_n8422_), .Y(new_n27432_));
  INVX1    g24996(.A(new_n27432_), .Y(new_n27433_));
  MX2X1    g24997(.A(new_n27429_), .B(new_n25281_), .S0(pi0211), .Y(new_n27434_));
  INVX1    g24998(.A(new_n27429_), .Y(new_n27435_));
  AOI21X1  g24999(.A0(new_n25281_), .A1(new_n23173_), .B0(pi0214), .Y(new_n27436_));
  OAI21X1  g25000(.A0(new_n27435_), .A1(new_n23173_), .B0(new_n27436_), .Y(new_n27437_));
  AND2X1   g25001(.A(new_n27437_), .B(pi0212), .Y(new_n27438_));
  OAI21X1  g25002(.A0(new_n27434_), .A1(new_n24849_), .B0(new_n27438_), .Y(new_n27439_));
  AOI21X1  g25003(.A0(new_n27439_), .A1(new_n27433_), .B0(new_n25282_), .Y(new_n27440_));
  NOR3X1   g25004(.A(new_n25280_), .B(po1038), .C(pi1152), .Y(new_n27441_));
  OAI22X1  g25005(.A0(new_n27441_), .A1(new_n27298_), .B0(new_n27440_), .B1(new_n27101_), .Y(new_n27442_));
  NAND2X1  g25006(.A(new_n25202_), .B(pi0214), .Y(new_n27443_));
  AOI21X1  g25007(.A0(new_n27443_), .A1(new_n25252_), .B0(pi0219), .Y(new_n27444_));
  AOI21X1  g25008(.A0(new_n25202_), .A1(new_n24849_), .B0(new_n24823_), .Y(new_n27445_));
  OAI21X1  g25009(.A0(new_n25218_), .A1(new_n24849_), .B0(new_n27445_), .Y(new_n27446_));
  OAI21X1  g25010(.A0(new_n25217_), .A1(new_n8422_), .B0(new_n6489_), .Y(new_n27447_));
  AOI21X1  g25011(.A0(new_n27446_), .A1(new_n27444_), .B0(new_n27447_), .Y(new_n27448_));
  AOI21X1  g25012(.A0(new_n25799_), .A1(new_n25216_), .B0(po1038), .Y(new_n27449_));
  OAI21X1  g25013(.A0(new_n25799_), .A1(new_n25218_), .B0(new_n27449_), .Y(new_n27450_));
  AOI21X1  g25014(.A0(new_n27450_), .A1(new_n27157_), .B0(new_n25153_), .Y(new_n27451_));
  OAI21X1  g25015(.A0(new_n27448_), .A1(new_n26263_), .B0(new_n27451_), .Y(new_n27452_));
  AOI21X1  g25016(.A0(new_n27452_), .A1(new_n27442_), .B0(pi1150), .Y(new_n27453_));
  NAND2X1  g25017(.A(new_n27434_), .B(new_n25188_), .Y(new_n27454_));
  AOI21X1  g25018(.A0(new_n25281_), .A1(new_n24816_), .B0(new_n8422_), .Y(new_n27455_));
  AOI21X1  g25019(.A0(new_n27455_), .A1(new_n27454_), .B0(po1038), .Y(new_n27456_));
  OAI21X1  g25020(.A0(new_n27429_), .A1(new_n24849_), .B0(new_n27438_), .Y(new_n27457_));
  NAND2X1  g25021(.A(new_n27457_), .B(new_n27433_), .Y(new_n27458_));
  AOI21X1  g25022(.A0(new_n27458_), .A1(new_n27456_), .B0(new_n27103_), .Y(new_n27459_));
  AOI21X1  g25023(.A0(new_n25281_), .A1(new_n24823_), .B0(pi0219), .Y(new_n27460_));
  OAI21X1  g25024(.A0(new_n27431_), .A1(new_n24823_), .B0(new_n27460_), .Y(new_n27461_));
  AOI21X1  g25025(.A0(new_n27461_), .A1(new_n27456_), .B0(new_n26312_), .Y(new_n27462_));
  OR3X1    g25026(.A(new_n27462_), .B(new_n27459_), .C(pi1152), .Y(new_n27463_));
  INVX1    g25027(.A(new_n25221_), .Y(new_n27464_));
  MX2X1    g25028(.A(new_n25218_), .B(new_n25217_), .S0(new_n24849_), .Y(new_n27465_));
  MX2X1    g25029(.A(new_n25216_), .B(new_n25202_), .S0(pi0211), .Y(new_n27466_));
  AOI21X1  g25030(.A0(new_n25218_), .A1(new_n24849_), .B0(new_n24823_), .Y(new_n27467_));
  OAI21X1  g25031(.A0(new_n27466_), .A1(new_n24849_), .B0(new_n27467_), .Y(new_n27468_));
  OAI21X1  g25032(.A0(new_n27465_), .A1(pi0212), .B0(new_n27468_), .Y(new_n27469_));
  AOI21X1  g25033(.A0(new_n27469_), .A1(new_n8422_), .B0(new_n27464_), .Y(new_n27470_));
  OAI21X1  g25034(.A0(new_n25202_), .A1(new_n24823_), .B0(new_n27444_), .Y(new_n27471_));
  NAND2X1  g25035(.A(new_n27471_), .B(new_n25221_), .Y(new_n27472_));
  AOI21X1  g25036(.A0(new_n27472_), .A1(new_n26318_), .B0(new_n25153_), .Y(new_n27473_));
  OAI21X1  g25037(.A0(new_n27470_), .A1(new_n27151_), .B0(new_n27473_), .Y(new_n27474_));
  AOI21X1  g25038(.A0(new_n27474_), .A1(new_n27463_), .B0(new_n26280_), .Y(new_n27475_));
  OAI21X1  g25039(.A0(new_n27475_), .A1(new_n27453_), .B0(new_n24815_), .Y(new_n27476_));
  AOI21X1  g25040(.A0(new_n25286_), .A1(pi0213), .B0(new_n24866_), .Y(new_n27477_));
  AOI22X1  g25041(.A0(new_n27477_), .A1(new_n27476_), .B0(new_n27424_), .B1(new_n27364_), .Y(new_n27478_));
  MX2X1    g25042(.A(new_n27478_), .B(pi0249), .S0(new_n24814_), .Y(po0406));
  NOR4X1   g25043(.A(new_n7766_), .B(new_n3378_), .C(new_n5881_), .D(new_n7763_), .Y(new_n27480_));
  OAI21X1  g25044(.A0(new_n27480_), .A1(new_n5076_), .B0(new_n3073_), .Y(new_n27481_));
  NAND3X1  g25045(.A(new_n5804_), .B(new_n3007_), .C(pi0075), .Y(new_n27482_));
  NAND3X1  g25046(.A(new_n6722_), .B(new_n7779_), .C(new_n3131_), .Y(new_n27483_));
  AOI21X1  g25047(.A0(new_n27482_), .A1(new_n27481_), .B0(new_n27483_), .Y(po0407));
  INVX1    g25048(.A(pi0476), .Y(new_n27485_));
  AOI22X1  g25049(.A0(new_n25004_), .A1(new_n27485_), .B0(new_n8055_), .B1(pi0897), .Y(new_n27486_));
  INVX1    g25050(.A(pi1053), .Y(new_n27487_));
  OR2X1    g25051(.A(new_n27487_), .B(pi0200), .Y(new_n27488_));
  AOI21X1  g25052(.A0(pi1039), .A1(pi0200), .B0(pi0199), .Y(new_n27489_));
  AND2X1   g25053(.A(new_n27489_), .B(new_n27488_), .Y(new_n27490_));
  INVX1    g25054(.A(new_n27490_), .Y(new_n27491_));
  MX2X1    g25055(.A(new_n27491_), .B(pi0251), .S0(new_n27486_), .Y(po0408));
  OAI21X1  g25056(.A0(new_n5023_), .A1(new_n5021_), .B0(new_n8541_), .Y(new_n27493_));
  NOR3X1   g25057(.A(new_n2985_), .B(new_n2536_), .C(pi0287), .Y(new_n27494_));
  INVX1    g25058(.A(new_n27494_), .Y(new_n27495_));
  INVX1    g25059(.A(pi1001), .Y(new_n27496_));
  OR2X1    g25060(.A(pi0984), .B(pi0979), .Y(new_n27497_));
  OR2X1    g25061(.A(new_n27497_), .B(new_n27496_), .Y(new_n27498_));
  OR4X1    g25062(.A(new_n27498_), .B(new_n27495_), .C(new_n5031_), .D(new_n5029_), .Y(new_n27499_));
  OR2X1    g25063(.A(pi1093), .B(new_n5024_), .Y(new_n27500_));
  AOI21X1  g25064(.A0(new_n27499_), .A1(new_n3035_), .B0(new_n27500_), .Y(new_n27501_));
  MX2X1    g25065(.A(new_n5236_), .B(new_n5235_), .S0(new_n27501_), .Y(new_n27502_));
  OAI21X1  g25066(.A0(new_n27502_), .A1(new_n6256_), .B0(new_n27493_), .Y(new_n27503_));
  MX2X1    g25067(.A(new_n27502_), .B(new_n8542_), .S0(new_n5043_), .Y(new_n27504_));
  OAI21X1  g25068(.A0(new_n27504_), .A1(new_n5058_), .B0(pi0299), .Y(new_n27505_));
  AOI21X1  g25069(.A0(new_n27503_), .A1(new_n5058_), .B0(new_n27505_), .Y(new_n27506_));
  OAI21X1  g25070(.A0(new_n27504_), .A1(new_n5041_), .B0(new_n2933_), .Y(new_n27507_));
  AOI21X1  g25071(.A0(new_n27503_), .A1(new_n5041_), .B0(new_n27507_), .Y(new_n27508_));
  OR3X1    g25072(.A(new_n27508_), .B(new_n27506_), .C(new_n8170_), .Y(new_n27509_));
  AOI21X1  g25073(.A0(new_n8541_), .A1(new_n8170_), .B0(new_n6713_), .Y(new_n27510_));
  OR4X1    g25074(.A(new_n27498_), .B(new_n5029_), .C(new_n2939_), .D(pi0038), .Y(new_n27511_));
  OR4X1    g25075(.A(new_n27511_), .B(new_n14616_), .C(new_n5034_), .D(new_n5031_), .Y(new_n27512_));
  OR2X1    g25076(.A(new_n27512_), .B(new_n24798_), .Y(new_n27513_));
  OAI21X1  g25077(.A0(new_n27513_), .A1(new_n27495_), .B0(new_n3035_), .Y(new_n27514_));
  AND2X1   g25078(.A(pi1092), .B(new_n2436_), .Y(new_n27515_));
  OAI21X1  g25079(.A0(new_n8540_), .A1(new_n2436_), .B0(new_n6713_), .Y(new_n27516_));
  AOI21X1  g25080(.A0(new_n27515_), .A1(new_n27514_), .B0(new_n27516_), .Y(new_n27517_));
  AOI21X1  g25081(.A0(new_n27510_), .A1(new_n27509_), .B0(new_n27517_), .Y(po0409));
  OR3X1    g25082(.A(new_n24961_), .B(new_n24884_), .C(new_n9446_), .Y(new_n27519_));
  NOR2X1   g25083(.A(new_n27519_), .B(po1038), .Y(new_n27520_));
  AOI21X1  g25084(.A0(new_n25956_), .A1(pi0219), .B0(new_n27520_), .Y(new_n27521_));
  INVX1    g25085(.A(new_n27521_), .Y(new_n27522_));
  AOI21X1  g25086(.A0(new_n27522_), .A1(pi1153), .B0(pi1151), .Y(new_n27523_));
  INVX1    g25087(.A(new_n7997_), .Y(new_n27524_));
  NOR2X1   g25088(.A(new_n24918_), .B(new_n24917_), .Y(new_n27525_));
  OAI22X1  g25089(.A0(new_n24948_), .A1(new_n27524_), .B0(new_n27525_), .B1(new_n23173_), .Y(new_n27526_));
  INVX1    g25090(.A(new_n27526_), .Y(new_n27527_));
  OAI22X1  g25091(.A0(new_n8423_), .A1(pi1153), .B0(pi0299), .B1(new_n7937_), .Y(new_n27528_));
  AOI21X1  g25092(.A0(new_n27528_), .A1(new_n24893_), .B0(po1038), .Y(new_n27529_));
  AND2X1   g25093(.A(new_n8422_), .B(pi0211), .Y(new_n27530_));
  OAI21X1  g25094(.A0(new_n25468_), .A1(new_n27530_), .B0(pi1151), .Y(new_n27531_));
  AOI21X1  g25095(.A0(new_n27529_), .A1(new_n27527_), .B0(new_n27531_), .Y(new_n27532_));
  OAI21X1  g25096(.A0(new_n27532_), .A1(new_n27523_), .B0(new_n25153_), .Y(new_n27533_));
  NOR4X1   g25097(.A(new_n24970_), .B(new_n12364_), .C(new_n8422_), .D(pi0211), .Y(new_n27534_));
  NOR4X1   g25098(.A(new_n27534_), .B(new_n24952_), .C(new_n8468_), .D(pi1151), .Y(new_n27535_));
  MX2X1    g25099(.A(pi0200), .B(pi0211), .S0(pi0299), .Y(new_n27536_));
  NOR2X1   g25100(.A(new_n27536_), .B(new_n12364_), .Y(new_n27537_));
  MX2X1    g25101(.A(new_n8422_), .B(new_n7871_), .S0(new_n2933_), .Y(new_n27538_));
  NOR3X1   g25102(.A(new_n27538_), .B(new_n27537_), .C(new_n25694_), .Y(new_n27539_));
  OR2X1    g25103(.A(new_n27539_), .B(po1038), .Y(new_n27540_));
  AOI21X1  g25104(.A0(new_n7997_), .A1(new_n25694_), .B0(new_n25467_), .Y(new_n27541_));
  AOI21X1  g25105(.A0(new_n27541_), .A1(po1038), .B0(new_n25153_), .Y(new_n27542_));
  OAI21X1  g25106(.A0(new_n27540_), .A1(new_n27535_), .B0(new_n27542_), .Y(new_n27543_));
  AOI21X1  g25107(.A0(new_n27543_), .A1(new_n27533_), .B0(new_n24814_), .Y(new_n27544_));
  INVX1    g25108(.A(pi0253), .Y(new_n27545_));
  NOR4X1   g25109(.A(new_n26539_), .B(new_n26526_), .C(new_n26522_), .D(new_n26521_), .Y(new_n27546_));
  OR2X1    g25110(.A(new_n27546_), .B(new_n12364_), .Y(new_n27547_));
  OR2X1    g25111(.A(new_n26582_), .B(pi1153), .Y(new_n27548_));
  AND3X1   g25112(.A(new_n27548_), .B(new_n27547_), .C(new_n8422_), .Y(new_n27549_));
  AOI21X1  g25113(.A0(new_n26526_), .A1(new_n26507_), .B0(new_n26539_), .Y(new_n27550_));
  INVX1    g25114(.A(new_n27550_), .Y(new_n27551_));
  AOI21X1  g25115(.A0(new_n26522_), .A1(new_n23173_), .B0(new_n27551_), .Y(new_n27552_));
  NOR3X1   g25116(.A(new_n26544_), .B(new_n26535_), .C(new_n26521_), .Y(new_n27553_));
  AOI21X1  g25117(.A0(new_n27553_), .A1(new_n27552_), .B0(new_n12364_), .Y(new_n27554_));
  NOR2X1   g25118(.A(new_n26633_), .B(pi1153), .Y(new_n27555_));
  NOR3X1   g25119(.A(new_n27555_), .B(new_n27554_), .C(new_n8422_), .Y(new_n27556_));
  OR3X1    g25120(.A(new_n27556_), .B(new_n27549_), .C(new_n27545_), .Y(new_n27557_));
  NOR2X1   g25121(.A(new_n26579_), .B(new_n26529_), .Y(new_n27558_));
  INVX1    g25122(.A(new_n27558_), .Y(new_n27559_));
  NOR2X1   g25123(.A(new_n26530_), .B(new_n26529_), .Y(new_n27560_));
  NOR4X1   g25124(.A(new_n26535_), .B(new_n26533_), .C(new_n26556_), .D(pi0211), .Y(new_n27561_));
  OAI21X1  g25125(.A0(new_n27561_), .A1(new_n27560_), .B0(pi1153), .Y(new_n27562_));
  AND3X1   g25126(.A(new_n27562_), .B(new_n27559_), .C(pi0219), .Y(new_n27563_));
  OR3X1    g25127(.A(new_n26539_), .B(new_n26530_), .C(new_n12364_), .Y(new_n27564_));
  NOR3X1   g25128(.A(new_n26579_), .B(new_n26539_), .C(pi1153), .Y(new_n27565_));
  INVX1    g25129(.A(new_n27565_), .Y(new_n27566_));
  AND3X1   g25130(.A(new_n27566_), .B(new_n27564_), .C(new_n8422_), .Y(new_n27567_));
  OR3X1    g25131(.A(new_n27567_), .B(new_n27563_), .C(pi0253), .Y(new_n27568_));
  AOI21X1  g25132(.A0(new_n27568_), .A1(new_n27557_), .B0(po1038), .Y(new_n27569_));
  AOI21X1  g25133(.A0(new_n26516_), .A1(new_n2702_), .B0(pi0219), .Y(new_n27570_));
  INVX1    g25134(.A(new_n27570_), .Y(new_n27571_));
  AOI21X1  g25135(.A0(new_n26515_), .A1(new_n23173_), .B0(new_n27571_), .Y(new_n27572_));
  NOR4X1   g25136(.A(new_n27572_), .B(new_n26505_), .C(new_n6489_), .D(pi0219), .Y(new_n27573_));
  NAND2X1  g25137(.A(pi1091), .B(pi0219), .Y(new_n27574_));
  AOI21X1  g25138(.A0(pi1153), .A1(new_n23173_), .B0(new_n27574_), .Y(new_n27575_));
  OR3X1    g25139(.A(new_n27575_), .B(new_n27570_), .C(new_n26568_), .Y(new_n27576_));
  AOI21X1  g25140(.A0(new_n26568_), .A1(pi0211), .B0(new_n8422_), .Y(new_n27577_));
  OAI21X1  g25141(.A0(new_n26505_), .A1(pi0211), .B0(new_n27577_), .Y(new_n27578_));
  NOR2X1   g25142(.A(new_n26514_), .B(pi0219), .Y(new_n27579_));
  NOR2X1   g25143(.A(new_n27579_), .B(new_n27575_), .Y(new_n27580_));
  AOI21X1  g25144(.A0(new_n27580_), .A1(new_n27578_), .B0(pi0253), .Y(new_n27581_));
  OR2X1    g25145(.A(new_n27581_), .B(new_n6489_), .Y(new_n27582_));
  AOI21X1  g25146(.A0(new_n27576_), .A1(pi0253), .B0(new_n27582_), .Y(new_n27583_));
  NOR3X1   g25147(.A(new_n27583_), .B(new_n27573_), .C(new_n25694_), .Y(new_n27584_));
  INVX1    g25148(.A(new_n27584_), .Y(new_n27585_));
  INVX1    g25149(.A(new_n26530_), .Y(new_n27586_));
  OAI21X1  g25150(.A0(new_n26544_), .A1(new_n26539_), .B0(new_n12364_), .Y(new_n27587_));
  AND3X1   g25151(.A(new_n27587_), .B(new_n27552_), .C(new_n27586_), .Y(new_n27588_));
  NAND3X1  g25152(.A(new_n26526_), .B(new_n26507_), .C(pi0219), .Y(new_n27589_));
  OAI21X1  g25153(.A0(new_n27588_), .A1(pi0219), .B0(new_n27589_), .Y(new_n27590_));
  OAI21X1  g25154(.A0(new_n27590_), .A1(new_n27563_), .B0(new_n27545_), .Y(new_n27591_));
  NOR2X1   g25155(.A(new_n26544_), .B(new_n26521_), .Y(new_n27592_));
  INVX1    g25156(.A(new_n27592_), .Y(new_n27593_));
  NOR2X1   g25157(.A(new_n26522_), .B(new_n26521_), .Y(new_n27594_));
  INVX1    g25158(.A(new_n27594_), .Y(new_n27595_));
  INVX1    g25159(.A(new_n27561_), .Y(new_n27596_));
  AOI21X1  g25160(.A0(new_n27596_), .A1(new_n27595_), .B0(new_n27571_), .Y(new_n27597_));
  INVX1    g25161(.A(new_n27597_), .Y(new_n27598_));
  AOI21X1  g25162(.A0(new_n27587_), .A1(new_n27593_), .B0(new_n27598_), .Y(new_n27599_));
  OR3X1    g25163(.A(new_n26535_), .B(new_n26521_), .C(new_n8422_), .Y(new_n27600_));
  AOI21X1  g25164(.A0(new_n27554_), .A1(new_n26612_), .B0(new_n27600_), .Y(new_n27601_));
  OAI21X1  g25165(.A0(new_n27601_), .A1(new_n27599_), .B0(pi0253), .Y(new_n27602_));
  AND3X1   g25166(.A(new_n27602_), .B(new_n27591_), .C(new_n6489_), .Y(new_n27603_));
  OAI22X1  g25167(.A0(new_n27603_), .A1(pi1151), .B0(new_n27585_), .B1(new_n27569_), .Y(new_n27604_));
  OAI21X1  g25168(.A0(new_n26505_), .A1(pi0211), .B0(new_n27579_), .Y(new_n27605_));
  AND2X1   g25169(.A(new_n27605_), .B(new_n27570_), .Y(new_n27606_));
  NOR2X1   g25170(.A(new_n26505_), .B(new_n8422_), .Y(new_n27607_));
  NOR2X1   g25171(.A(new_n27607_), .B(new_n6489_), .Y(new_n27608_));
  INVX1    g25172(.A(new_n27608_), .Y(new_n27609_));
  NOR2X1   g25173(.A(new_n27609_), .B(new_n27606_), .Y(new_n27610_));
  AOI21X1  g25174(.A0(new_n27610_), .A1(new_n26694_), .B0(new_n27583_), .Y(new_n27611_));
  AOI21X1  g25175(.A0(new_n27611_), .A1(new_n27604_), .B0(new_n25153_), .Y(new_n27612_));
  AND2X1   g25176(.A(new_n27562_), .B(new_n27559_), .Y(new_n27613_));
  OAI22X1  g25177(.A0(new_n27598_), .A1(new_n27567_), .B0(new_n27613_), .B1(new_n8422_), .Y(new_n27614_));
  AOI21X1  g25178(.A0(new_n27614_), .A1(new_n26534_), .B0(pi0253), .Y(new_n27615_));
  AND2X1   g25179(.A(new_n27570_), .B(new_n27552_), .Y(new_n27616_));
  OAI21X1  g25180(.A0(new_n26562_), .A1(new_n12364_), .B0(new_n27616_), .Y(new_n27617_));
  AOI21X1  g25181(.A0(new_n27553_), .A1(new_n27552_), .B0(new_n26602_), .Y(new_n27618_));
  NAND2X1  g25182(.A(new_n27618_), .B(pi1153), .Y(new_n27619_));
  OAI21X1  g25183(.A0(new_n26535_), .A1(new_n26527_), .B0(new_n12364_), .Y(new_n27620_));
  NAND3X1  g25184(.A(new_n27620_), .B(new_n27619_), .C(pi0219), .Y(new_n27621_));
  AOI21X1  g25185(.A0(new_n27621_), .A1(new_n27617_), .B0(new_n27545_), .Y(new_n27622_));
  OR3X1    g25186(.A(new_n27622_), .B(new_n27615_), .C(po1038), .Y(new_n27623_));
  OR3X1    g25187(.A(new_n27613_), .B(new_n26556_), .C(new_n8422_), .Y(new_n27624_));
  INVX1    g25188(.A(new_n26582_), .Y(new_n27625_));
  AND2X1   g25189(.A(new_n26554_), .B(new_n12364_), .Y(new_n27626_));
  OR4X1    g25190(.A(new_n27626_), .B(new_n27625_), .C(new_n26533_), .D(pi0219), .Y(new_n27627_));
  AND2X1   g25191(.A(new_n27627_), .B(new_n27545_), .Y(new_n27628_));
  NOR2X1   g25192(.A(new_n26544_), .B(new_n26529_), .Y(new_n27629_));
  AND2X1   g25193(.A(new_n27553_), .B(new_n27552_), .Y(new_n27630_));
  AOI21X1  g25194(.A0(new_n27559_), .A1(new_n2702_), .B0(pi1153), .Y(new_n27631_));
  NOR3X1   g25195(.A(new_n26544_), .B(new_n26539_), .C(pi0219), .Y(new_n27632_));
  NOR4X1   g25196(.A(new_n27632_), .B(new_n27631_), .C(new_n27630_), .D(new_n27629_), .Y(new_n27633_));
  OAI21X1  g25197(.A0(new_n27633_), .A1(new_n27545_), .B0(new_n6489_), .Y(new_n27634_));
  AOI21X1  g25198(.A0(new_n27628_), .A1(new_n27624_), .B0(new_n27634_), .Y(new_n27635_));
  OR2X1    g25199(.A(new_n27583_), .B(pi1151), .Y(new_n27636_));
  OAI21X1  g25200(.A0(new_n27636_), .A1(new_n27635_), .B0(new_n25153_), .Y(new_n27637_));
  AOI21X1  g25201(.A0(new_n27623_), .A1(new_n27584_), .B0(new_n27637_), .Y(new_n27638_));
  OAI21X1  g25202(.A0(new_n27638_), .A1(new_n27612_), .B0(new_n26711_), .Y(new_n27639_));
  NOR2X1   g25203(.A(new_n26650_), .B(pi1153), .Y(new_n27640_));
  OAI21X1  g25204(.A0(new_n26671_), .A1(new_n12364_), .B0(new_n24893_), .Y(new_n27641_));
  OAI22X1  g25205(.A0(new_n27641_), .A1(new_n27640_), .B0(new_n27527_), .B1(new_n2702_), .Y(new_n27642_));
  NAND2X1  g25206(.A(new_n27642_), .B(pi0253), .Y(new_n27643_));
  OAI21X1  g25207(.A0(new_n27537_), .A1(new_n9448_), .B0(pi1091), .Y(new_n27644_));
  AOI21X1  g25208(.A0(new_n27644_), .A1(new_n27545_), .B0(po1038), .Y(new_n27645_));
  NOR2X1   g25209(.A(pi1091), .B(pi0253), .Y(new_n27646_));
  OR2X1    g25210(.A(new_n27646_), .B(new_n6489_), .Y(new_n27647_));
  AND2X1   g25211(.A(pi1091), .B(pi0211), .Y(new_n27648_));
  INVX1    g25212(.A(new_n27648_), .Y(new_n27649_));
  OR2X1    g25213(.A(pi1153), .B(new_n2702_), .Y(new_n27650_));
  OAI21X1  g25214(.A0(new_n27650_), .A1(new_n8422_), .B0(new_n27649_), .Y(new_n27651_));
  OAI21X1  g25215(.A0(new_n27651_), .A1(new_n27647_), .B0(pi1151), .Y(new_n27652_));
  AOI21X1  g25216(.A0(new_n27645_), .A1(new_n27643_), .B0(new_n27652_), .Y(new_n27653_));
  NOR4X1   g25217(.A(new_n27646_), .B(new_n27575_), .C(new_n6489_), .D(new_n8422_), .Y(new_n27654_));
  NOR4X1   g25218(.A(new_n27519_), .B(po1038), .C(new_n12364_), .D(new_n2702_), .Y(new_n27655_));
  AND2X1   g25219(.A(new_n2702_), .B(pi0253), .Y(new_n27656_));
  NOR4X1   g25220(.A(new_n27656_), .B(new_n27655_), .C(new_n27654_), .D(pi1151), .Y(new_n27657_));
  OAI21X1  g25221(.A0(new_n27657_), .A1(new_n27653_), .B0(new_n25153_), .Y(new_n27658_));
  OAI21X1  g25222(.A0(new_n8467_), .A1(new_n2702_), .B0(new_n12364_), .Y(new_n27659_));
  NOR3X1   g25223(.A(new_n24903_), .B(new_n2702_), .C(pi0299), .Y(new_n27660_));
  NOR2X1   g25224(.A(new_n27660_), .B(new_n12364_), .Y(new_n27661_));
  NOR2X1   g25225(.A(new_n27661_), .B(new_n24894_), .Y(new_n27662_));
  NAND2X1  g25226(.A(new_n27662_), .B(new_n27659_), .Y(new_n27663_));
  INVX1    g25227(.A(new_n27530_), .Y(new_n27664_));
  NOR4X1   g25228(.A(new_n24952_), .B(new_n27664_), .C(new_n2702_), .D(pi0299), .Y(new_n27665_));
  NOR2X1   g25229(.A(new_n27665_), .B(new_n27545_), .Y(new_n27666_));
  NOR3X1   g25230(.A(new_n24970_), .B(new_n12364_), .C(new_n2702_), .Y(new_n27667_));
  AND3X1   g25231(.A(new_n25207_), .B(new_n24946_), .C(pi1091), .Y(new_n27668_));
  OR3X1    g25232(.A(new_n27668_), .B(new_n27667_), .C(new_n24894_), .Y(new_n27669_));
  NOR4X1   g25233(.A(new_n24918_), .B(new_n24911_), .C(new_n2702_), .D(pi0299), .Y(new_n27670_));
  OR3X1    g25234(.A(new_n27670_), .B(new_n26684_), .C(new_n23173_), .Y(new_n27671_));
  AND3X1   g25235(.A(new_n27671_), .B(new_n27669_), .C(new_n27545_), .Y(new_n27672_));
  AOI21X1  g25236(.A0(new_n27666_), .A1(new_n27663_), .B0(new_n27672_), .Y(new_n27673_));
  XOR2X1   g25237(.A(pi0219), .B(new_n23173_), .Y(new_n27674_));
  INVX1    g25238(.A(new_n27674_), .Y(new_n27675_));
  NOR3X1   g25239(.A(new_n27675_), .B(new_n27670_), .C(new_n27656_), .Y(new_n27676_));
  OR4X1    g25240(.A(new_n27676_), .B(new_n27673_), .C(po1038), .D(pi1151), .Y(new_n27677_));
  OAI21X1  g25241(.A0(pi1091), .A1(new_n27545_), .B0(new_n27536_), .Y(new_n27678_));
  AOI21X1  g25242(.A0(new_n27678_), .A1(new_n27650_), .B0(new_n27538_), .Y(new_n27679_));
  OAI21X1  g25243(.A0(pi1091), .A1(pi0253), .B0(new_n6489_), .Y(new_n27680_));
  OAI22X1  g25244(.A0(new_n27680_), .A1(new_n27679_), .B0(new_n27647_), .B1(new_n27575_), .Y(new_n27681_));
  AND3X1   g25245(.A(pi1091), .B(new_n8422_), .C(new_n23173_), .Y(new_n27682_));
  NOR4X1   g25246(.A(new_n27682_), .B(new_n27646_), .C(new_n27575_), .D(new_n6489_), .Y(new_n27683_));
  OR2X1    g25247(.A(new_n27683_), .B(new_n25153_), .Y(new_n27684_));
  AOI21X1  g25248(.A0(new_n27681_), .A1(pi1151), .B0(new_n27684_), .Y(new_n27685_));
  AOI21X1  g25249(.A0(new_n27685_), .A1(new_n27677_), .B0(new_n26711_), .Y(new_n27686_));
  AOI21X1  g25250(.A0(new_n27686_), .A1(new_n27658_), .B0(pi0230), .Y(new_n27687_));
  AOI21X1  g25251(.A0(new_n27687_), .A1(new_n27639_), .B0(new_n27544_), .Y(po0410));
  INVX1    g25252(.A(new_n25190_), .Y(new_n27689_));
  OAI22X1  g25253(.A0(new_n25257_), .A1(new_n24998_), .B0(new_n25234_), .B1(new_n12487_), .Y(new_n27690_));
  OAI21X1  g25254(.A0(pi0219), .A1(new_n23173_), .B0(new_n25208_), .Y(new_n27691_));
  OAI21X1  g25255(.A0(new_n24894_), .A1(new_n2933_), .B0(new_n27691_), .Y(new_n27692_));
  AOI22X1  g25256(.A0(new_n27692_), .A1(new_n27689_), .B0(new_n27690_), .B1(new_n27530_), .Y(new_n27693_));
  AOI21X1  g25257(.A0(pi1153), .A1(pi0211), .B0(pi0219), .Y(new_n27694_));
  NOR2X1   g25258(.A(new_n27694_), .B(new_n25337_), .Y(new_n27695_));
  AOI21X1  g25259(.A0(new_n27695_), .A1(po1038), .B0(pi1152), .Y(new_n27696_));
  OAI21X1  g25260(.A0(new_n27693_), .A1(po1038), .B0(new_n27696_), .Y(new_n27697_));
  NAND2X1  g25261(.A(pi1154), .B(pi0211), .Y(new_n27698_));
  MX2X1    g25262(.A(new_n24916_), .B(new_n24907_), .S0(pi1153), .Y(new_n27699_));
  NOR2X1   g25263(.A(new_n27699_), .B(new_n27698_), .Y(new_n27700_));
  NOR2X1   g25264(.A(new_n25276_), .B(pi1154), .Y(new_n27701_));
  OR3X1    g25265(.A(new_n27701_), .B(new_n27700_), .C(new_n25192_), .Y(new_n27702_));
  OR2X1    g25266(.A(new_n12487_), .B(pi0200), .Y(new_n27703_));
  AOI22X1  g25267(.A0(new_n27703_), .A1(new_n24950_), .B0(new_n26051_), .B1(new_n25235_), .Y(new_n27704_));
  OAI21X1  g25268(.A0(new_n27704_), .A1(pi0219), .B0(new_n6489_), .Y(new_n27705_));
  AOI21X1  g25269(.A0(new_n27702_), .A1(pi0219), .B0(new_n27705_), .Y(new_n27706_));
  AND3X1   g25270(.A(new_n12364_), .B(new_n8422_), .C(pi0211), .Y(new_n27707_));
  NOR3X1   g25271(.A(new_n27707_), .B(new_n25337_), .C(new_n6489_), .Y(new_n27708_));
  OR2X1    g25272(.A(new_n27708_), .B(new_n25153_), .Y(new_n27709_));
  OAI21X1  g25273(.A0(new_n27709_), .A1(new_n27706_), .B0(new_n27697_), .Y(new_n27710_));
  INVX1    g25274(.A(new_n26711_), .Y(new_n27711_));
  AOI21X1  g25275(.A0(new_n27588_), .A1(new_n12364_), .B0(new_n26582_), .Y(new_n27712_));
  INVX1    g25276(.A(pi0254), .Y(new_n27713_));
  NOR3X1   g25277(.A(new_n26514_), .B(new_n2933_), .C(pi0211), .Y(new_n27714_));
  NOR4X1   g25278(.A(new_n27714_), .B(new_n27551_), .C(new_n26526_), .D(new_n12487_), .Y(new_n27715_));
  AOI21X1  g25279(.A0(new_n27715_), .A1(new_n27547_), .B0(new_n27713_), .Y(new_n27716_));
  OAI21X1  g25280(.A0(new_n27712_), .A1(pi1154), .B0(new_n27716_), .Y(new_n27717_));
  NOR4X1   g25281(.A(new_n26535_), .B(new_n26530_), .C(new_n26527_), .D(new_n12487_), .Y(new_n27718_));
  OAI21X1  g25282(.A0(new_n26553_), .A1(new_n23173_), .B0(new_n26534_), .Y(new_n27719_));
  AOI21X1  g25283(.A0(new_n27719_), .A1(new_n12364_), .B0(pi0254), .Y(new_n27720_));
  OAI21X1  g25284(.A0(new_n27718_), .A1(new_n26580_), .B0(new_n27720_), .Y(new_n27721_));
  AOI21X1  g25285(.A0(new_n27721_), .A1(new_n27717_), .B0(pi0219), .Y(new_n27722_));
  NOR3X1   g25286(.A(new_n27618_), .B(new_n27554_), .C(new_n12487_), .Y(new_n27723_));
  OR2X1    g25287(.A(new_n26633_), .B(new_n12364_), .Y(new_n27724_));
  AND3X1   g25288(.A(new_n27724_), .B(new_n27620_), .C(new_n12487_), .Y(new_n27725_));
  OR3X1    g25289(.A(new_n27725_), .B(new_n27723_), .C(new_n27713_), .Y(new_n27726_));
  INVX1    g25290(.A(new_n25488_), .Y(new_n27727_));
  INVX1    g25291(.A(new_n27555_), .Y(new_n27728_));
  NOR3X1   g25292(.A(new_n26535_), .B(new_n26530_), .C(new_n26527_), .Y(new_n27729_));
  AOI21X1  g25293(.A0(new_n27729_), .A1(new_n27728_), .B0(new_n27727_), .Y(new_n27730_));
  NAND2X1  g25294(.A(new_n27730_), .B(new_n26506_), .Y(new_n27731_));
  NOR2X1   g25295(.A(new_n26569_), .B(pi1153), .Y(new_n27732_));
  NOR4X1   g25296(.A(new_n27732_), .B(new_n26579_), .C(new_n26529_), .D(new_n26526_), .Y(new_n27733_));
  NOR2X1   g25297(.A(new_n27733_), .B(pi1154), .Y(new_n27734_));
  OAI21X1  g25298(.A0(new_n27559_), .A1(new_n26533_), .B0(new_n27734_), .Y(new_n27735_));
  NOR3X1   g25299(.A(new_n26530_), .B(new_n26529_), .C(new_n12364_), .Y(new_n27736_));
  OR3X1    g25300(.A(new_n27736_), .B(new_n26623_), .C(new_n27698_), .Y(new_n27737_));
  NAND4X1  g25301(.A(new_n27737_), .B(new_n27735_), .C(new_n27731_), .D(new_n27713_), .Y(new_n27738_));
  AOI21X1  g25302(.A0(new_n27738_), .A1(new_n27726_), .B0(new_n8422_), .Y(new_n27739_));
  OR3X1    g25303(.A(new_n27739_), .B(new_n27722_), .C(new_n27545_), .Y(new_n27740_));
  AOI21X1  g25304(.A0(new_n26660_), .A1(new_n2933_), .B0(new_n12364_), .Y(new_n27741_));
  OR2X1    g25305(.A(new_n27741_), .B(pi1154), .Y(new_n27742_));
  OAI22X1  g25306(.A0(new_n26650_), .A1(pi1153), .B0(new_n25242_), .B1(pi0211), .Y(new_n27743_));
  OR3X1    g25307(.A(new_n24916_), .B(new_n27698_), .C(new_n2702_), .Y(new_n27744_));
  OAI22X1  g25308(.A0(new_n27744_), .A1(new_n25264_), .B0(new_n27743_), .B1(new_n27742_), .Y(new_n27745_));
  AND2X1   g25309(.A(pi1091), .B(new_n23173_), .Y(new_n27746_));
  INVX1    g25310(.A(new_n27746_), .Y(new_n27747_));
  OAI21X1  g25311(.A0(new_n27747_), .A1(new_n12487_), .B0(new_n27574_), .Y(new_n27748_));
  AOI22X1  g25312(.A0(new_n27748_), .A1(new_n27702_), .B0(new_n27745_), .B1(new_n8422_), .Y(new_n27749_));
  NOR2X1   g25313(.A(new_n27536_), .B(new_n12487_), .Y(new_n27750_));
  OR3X1    g25314(.A(new_n27750_), .B(new_n25276_), .C(new_n8422_), .Y(new_n27751_));
  OAI21X1  g25315(.A0(new_n27704_), .A1(pi0219), .B0(new_n27751_), .Y(new_n27752_));
  OAI21X1  g25316(.A0(new_n27752_), .A1(new_n2702_), .B0(new_n27713_), .Y(new_n27753_));
  OAI21X1  g25317(.A0(new_n27749_), .A1(new_n27713_), .B0(new_n27753_), .Y(new_n27754_));
  AOI21X1  g25318(.A0(new_n27754_), .A1(new_n27545_), .B0(po1038), .Y(new_n27755_));
  OAI21X1  g25319(.A0(new_n26695_), .A1(pi0211), .B0(new_n27607_), .Y(new_n27756_));
  AND2X1   g25320(.A(new_n26514_), .B(new_n8422_), .Y(new_n27757_));
  INVX1    g25321(.A(new_n27757_), .Y(new_n27758_));
  AND2X1   g25322(.A(new_n25337_), .B(pi1091), .Y(new_n27759_));
  NOR4X1   g25323(.A(pi1153), .B(new_n2702_), .C(pi0219), .D(new_n23173_), .Y(new_n27760_));
  NOR3X1   g25324(.A(new_n27760_), .B(new_n27759_), .C(new_n27713_), .Y(new_n27761_));
  AND3X1   g25325(.A(new_n27761_), .B(new_n27758_), .C(new_n27756_), .Y(new_n27762_));
  INVX1    g25326(.A(new_n27578_), .Y(new_n27763_));
  AND2X1   g25327(.A(pi1153), .B(pi1091), .Y(new_n27764_));
  NOR2X1   g25328(.A(new_n27764_), .B(new_n27605_), .Y(new_n27765_));
  NOR4X1   g25329(.A(new_n27765_), .B(new_n27759_), .C(new_n27763_), .D(pi0254), .Y(new_n27766_));
  NOR3X1   g25330(.A(new_n27766_), .B(new_n27762_), .C(new_n27545_), .Y(new_n27767_));
  AOI22X1  g25331(.A0(new_n5102_), .A1(new_n2436_), .B0(new_n2702_), .B1(new_n27713_), .Y(new_n27768_));
  OAI21X1  g25332(.A0(new_n27695_), .A1(new_n2702_), .B0(new_n27768_), .Y(new_n27769_));
  OAI21X1  g25333(.A0(new_n5103_), .A1(pi0057), .B0(new_n27682_), .Y(new_n27770_));
  OR2X1    g25334(.A(new_n6489_), .B(new_n27545_), .Y(new_n27771_));
  AND3X1   g25335(.A(new_n27771_), .B(new_n27770_), .C(new_n27769_), .Y(new_n27772_));
  OAI21X1  g25336(.A0(new_n27772_), .A1(new_n27767_), .B0(pi1152), .Y(new_n27773_));
  AOI21X1  g25337(.A0(new_n27755_), .A1(new_n27740_), .B0(new_n27773_), .Y(new_n27774_));
  NOR4X1   g25338(.A(new_n26533_), .B(new_n26529_), .C(new_n26556_), .D(pi1154), .Y(new_n27775_));
  NOR3X1   g25339(.A(new_n26544_), .B(new_n26535_), .C(pi1153), .Y(new_n27776_));
  OR3X1    g25340(.A(new_n27776_), .B(new_n27775_), .C(new_n27553_), .Y(new_n27777_));
  AOI21X1  g25341(.A0(new_n26612_), .A1(new_n25488_), .B0(new_n8422_), .Y(new_n27778_));
  OR3X1    g25342(.A(new_n27776_), .B(new_n27561_), .C(new_n27594_), .Y(new_n27779_));
  OR4X1    g25343(.A(new_n26525_), .B(new_n26517_), .C(new_n12487_), .D(pi0299), .Y(new_n27780_));
  AND2X1   g25344(.A(new_n27780_), .B(new_n8422_), .Y(new_n27781_));
  AOI22X1  g25345(.A0(new_n27781_), .A1(new_n27779_), .B0(new_n27778_), .B1(new_n27777_), .Y(new_n27782_));
  AOI21X1  g25346(.A0(new_n27728_), .A1(new_n26531_), .B0(new_n27698_), .Y(new_n27783_));
  NOR4X1   g25347(.A(new_n27783_), .B(new_n27734_), .C(new_n27730_), .D(new_n8422_), .Y(new_n27784_));
  NOR4X1   g25348(.A(new_n27626_), .B(new_n26579_), .C(new_n26539_), .D(new_n26526_), .Y(new_n27785_));
  NOR2X1   g25349(.A(new_n27785_), .B(pi1154), .Y(new_n27786_));
  NOR3X1   g25350(.A(new_n26533_), .B(new_n26522_), .C(new_n26556_), .Y(new_n27787_));
  OR3X1    g25351(.A(new_n27787_), .B(new_n27785_), .C(new_n12487_), .Y(new_n27788_));
  AND3X1   g25352(.A(new_n26526_), .B(new_n26507_), .C(pi1154), .Y(new_n27789_));
  OAI21X1  g25353(.A0(new_n27789_), .A1(new_n26522_), .B0(new_n23173_), .Y(new_n27790_));
  NAND3X1  g25354(.A(new_n27790_), .B(new_n27788_), .C(new_n8422_), .Y(new_n27791_));
  OAI21X1  g25355(.A0(new_n27791_), .A1(new_n27786_), .B0(new_n27713_), .Y(new_n27792_));
  OAI22X1  g25356(.A0(new_n27792_), .A1(new_n27784_), .B0(new_n27782_), .B1(new_n27713_), .Y(new_n27793_));
  AND3X1   g25357(.A(new_n26652_), .B(new_n12364_), .C(pi1091), .Y(new_n27794_));
  OR2X1    g25358(.A(new_n27794_), .B(new_n27667_), .Y(new_n27795_));
  AND3X1   g25359(.A(new_n27795_), .B(new_n27742_), .C(pi0211), .Y(new_n27796_));
  AOI21X1  g25360(.A0(new_n25208_), .A1(pi1091), .B0(new_n12487_), .Y(new_n27797_));
  AOI21X1  g25361(.A0(new_n27764_), .A1(new_n8467_), .B0(pi1154), .Y(new_n27798_));
  NOR3X1   g25362(.A(new_n27798_), .B(new_n27797_), .C(pi0211), .Y(new_n27799_));
  OAI21X1  g25363(.A0(new_n27799_), .A1(new_n27796_), .B0(new_n8422_), .Y(new_n27800_));
  AND2X1   g25364(.A(new_n27797_), .B(pi0211), .Y(new_n27801_));
  NOR3X1   g25365(.A(new_n24961_), .B(pi1153), .C(new_n2702_), .Y(new_n27802_));
  NOR3X1   g25366(.A(new_n27802_), .B(new_n27667_), .C(new_n27727_), .Y(new_n27803_));
  NOR4X1   g25367(.A(new_n27803_), .B(new_n27801_), .C(new_n27798_), .D(new_n8422_), .Y(new_n27804_));
  INVX1    g25368(.A(new_n27804_), .Y(new_n27805_));
  AOI21X1  g25369(.A0(new_n27805_), .A1(new_n27800_), .B0(pi0254), .Y(new_n27806_));
  OAI21X1  g25370(.A0(pi0219), .A1(new_n23173_), .B0(pi1091), .Y(new_n27807_));
  OAI21X1  g25371(.A0(new_n27807_), .A1(new_n25189_), .B0(new_n12487_), .Y(new_n27808_));
  NOR2X1   g25372(.A(new_n26652_), .B(new_n2702_), .Y(new_n27809_));
  MX2X1    g25373(.A(new_n27660_), .B(new_n27809_), .S0(new_n12364_), .Y(new_n27810_));
  AOI21X1  g25374(.A0(new_n24903_), .A1(new_n2933_), .B0(new_n2702_), .Y(new_n27811_));
  OR2X1    g25375(.A(new_n27811_), .B(new_n27810_), .Y(new_n27812_));
  AND2X1   g25376(.A(new_n27812_), .B(new_n27674_), .Y(new_n27813_));
  NOR4X1   g25377(.A(new_n27661_), .B(new_n24992_), .C(new_n24894_), .D(new_n2702_), .Y(new_n27814_));
  NOR2X1   g25378(.A(new_n27814_), .B(new_n12487_), .Y(new_n27815_));
  INVX1    g25379(.A(new_n27815_), .Y(new_n27816_));
  OAI21X1  g25380(.A0(new_n27816_), .A1(new_n27813_), .B0(new_n27808_), .Y(new_n27817_));
  AND2X1   g25381(.A(new_n12487_), .B(pi1091), .Y(new_n27818_));
  AOI21X1  g25382(.A0(new_n27818_), .A1(new_n24998_), .B0(new_n27810_), .Y(new_n27819_));
  OAI21X1  g25383(.A0(new_n27819_), .A1(new_n27664_), .B0(pi0254), .Y(new_n27820_));
  INVX1    g25384(.A(new_n27820_), .Y(new_n27821_));
  AOI21X1  g25385(.A0(new_n27821_), .A1(new_n27817_), .B0(new_n27806_), .Y(new_n27822_));
  AND2X1   g25386(.A(new_n27822_), .B(new_n27545_), .Y(new_n27823_));
  OR2X1    g25387(.A(new_n27823_), .B(po1038), .Y(new_n27824_));
  AOI21X1  g25388(.A0(new_n27793_), .A1(pi0253), .B0(new_n27824_), .Y(new_n27825_));
  NAND2X1  g25389(.A(new_n27605_), .B(new_n27570_), .Y(new_n27826_));
  NAND2X1  g25390(.A(new_n27762_), .B(new_n27826_), .Y(new_n27827_));
  OR2X1    g25391(.A(new_n27572_), .B(pi0219), .Y(new_n27828_));
  AOI21X1  g25392(.A0(new_n27766_), .A1(new_n27828_), .B0(new_n27545_), .Y(new_n27829_));
  AOI22X1  g25393(.A0(new_n27829_), .A1(new_n27827_), .B0(new_n27771_), .B1(new_n27769_), .Y(new_n27830_));
  NOR3X1   g25394(.A(new_n27830_), .B(new_n27825_), .C(pi1152), .Y(new_n27831_));
  OR3X1    g25395(.A(new_n27831_), .B(new_n27774_), .C(new_n27711_), .Y(new_n27832_));
  AND2X1   g25396(.A(new_n27769_), .B(new_n25153_), .Y(new_n27833_));
  OAI21X1  g25397(.A0(new_n27822_), .A1(po1038), .B0(new_n27833_), .Y(new_n27834_));
  AND3X1   g25398(.A(new_n27770_), .B(new_n27769_), .C(pi1152), .Y(new_n27835_));
  OAI21X1  g25399(.A0(new_n27754_), .A1(po1038), .B0(new_n27835_), .Y(new_n27836_));
  NAND3X1  g25400(.A(new_n27836_), .B(new_n27834_), .C(new_n27711_), .Y(new_n27837_));
  AND2X1   g25401(.A(new_n27837_), .B(new_n24814_), .Y(new_n27838_));
  AOI22X1  g25402(.A0(new_n27838_), .A1(new_n27832_), .B0(new_n27710_), .B1(pi0230), .Y(po0411));
  MX2X1    g25403(.A(pi1049), .B(pi1036), .S0(pi0200), .Y(new_n27840_));
  MX2X1    g25404(.A(new_n27840_), .B(pi0255), .S0(new_n27486_), .Y(po0412));
  MX2X1    g25405(.A(pi1048), .B(pi1070), .S0(pi0200), .Y(new_n27842_));
  MX2X1    g25406(.A(new_n27842_), .B(pi0256), .S0(new_n27486_), .Y(po0413));
  MX2X1    g25407(.A(pi1084), .B(pi1065), .S0(pi0200), .Y(new_n27844_));
  MX2X1    g25408(.A(new_n27844_), .B(pi0257), .S0(new_n27486_), .Y(po0414));
  MX2X1    g25409(.A(pi1072), .B(pi1062), .S0(pi0200), .Y(new_n27846_));
  MX2X1    g25410(.A(new_n27846_), .B(pi0258), .S0(new_n27486_), .Y(po0415));
  MX2X1    g25411(.A(pi1059), .B(pi1069), .S0(pi0200), .Y(new_n27848_));
  MX2X1    g25412(.A(new_n27848_), .B(pi0259), .S0(new_n27486_), .Y(po0416));
  INVX1    g25413(.A(pi1044), .Y(new_n27850_));
  AOI21X1  g25414(.A0(pi1067), .A1(pi0200), .B0(pi0199), .Y(new_n27851_));
  OAI21X1  g25415(.A0(new_n27850_), .A1(pi0200), .B0(new_n27851_), .Y(new_n27852_));
  MX2X1    g25416(.A(new_n27852_), .B(pi0260), .S0(new_n27486_), .Y(po0417));
  INVX1    g25417(.A(pi1037), .Y(new_n27854_));
  AOI21X1  g25418(.A0(pi1040), .A1(pi0200), .B0(pi0199), .Y(new_n27855_));
  OAI21X1  g25419(.A0(new_n27854_), .A1(pi0200), .B0(new_n27855_), .Y(new_n27856_));
  MX2X1    g25420(.A(new_n27856_), .B(pi0261), .S0(new_n27486_), .Y(po0418));
  MX2X1    g25421(.A(new_n24820_), .B(pi0262), .S0(new_n5032_), .Y(new_n27858_));
  OR2X1    g25422(.A(new_n27858_), .B(pi0228), .Y(new_n27859_));
  AOI21X1  g25423(.A0(pi0262), .A1(pi0123), .B0(new_n2793_), .Y(new_n27860_));
  OAI21X1  g25424(.A0(pi1142), .A1(pi0123), .B0(new_n27860_), .Y(new_n27861_));
  AND2X1   g25425(.A(new_n27861_), .B(new_n27859_), .Y(new_n27862_));
  INVX1    g25426(.A(new_n27862_), .Y(new_n27863_));
  INVX1    g25427(.A(pi0123), .Y(new_n27864_));
  MX2X1    g25428(.A(pi1093), .B(new_n27864_), .S0(pi0228), .Y(new_n27865_));
  OAI22X1  g25429(.A0(new_n27865_), .A1(pi0262), .B0(new_n26433_), .B1(new_n2933_), .Y(new_n27866_));
  AOI21X1  g25430(.A0(new_n27865_), .A1(pi0199), .B0(new_n24840_), .Y(new_n27867_));
  OR2X1    g25431(.A(new_n27867_), .B(new_n27866_), .Y(new_n27868_));
  OR3X1    g25432(.A(new_n27865_), .B(pi0262), .C(pi0207), .Y(new_n27869_));
  AOI22X1  g25433(.A0(new_n27869_), .A1(new_n22959_), .B0(new_n26432_), .B1(pi0299), .Y(new_n27870_));
  AOI21X1  g25434(.A0(new_n27868_), .A1(new_n27863_), .B0(new_n27870_), .Y(new_n27871_));
  AND2X1   g25435(.A(new_n27866_), .B(pi0299), .Y(new_n27872_));
  OAI21X1  g25436(.A0(new_n26031_), .A1(pi0199), .B0(new_n27865_), .Y(new_n27873_));
  NAND2X1  g25437(.A(new_n27873_), .B(new_n2933_), .Y(new_n27874_));
  OAI21X1  g25438(.A0(new_n27874_), .A1(new_n27862_), .B0(pi0208), .Y(new_n27875_));
  OAI21X1  g25439(.A0(new_n27875_), .A1(new_n27872_), .B0(new_n6489_), .Y(new_n27876_));
  AND2X1   g25440(.A(new_n27865_), .B(new_n26433_), .Y(new_n27877_));
  OR3X1    g25441(.A(new_n27877_), .B(new_n27862_), .C(new_n6489_), .Y(new_n27878_));
  OAI21X1  g25442(.A0(new_n27876_), .A1(new_n27871_), .B0(new_n27878_), .Y(po0419));
  AND2X1   g25443(.A(new_n26561_), .B(new_n12463_), .Y(new_n27880_));
  OR3X1    g25444(.A(new_n27880_), .B(new_n26540_), .C(new_n12487_), .Y(new_n27881_));
  NOR3X1   g25445(.A(new_n26579_), .B(new_n26539_), .C(new_n26526_), .Y(new_n27882_));
  OAI21X1  g25446(.A0(new_n26554_), .A1(pi1155), .B0(new_n12487_), .Y(new_n27883_));
  AOI21X1  g25447(.A0(new_n27882_), .A1(pi1155), .B0(new_n27883_), .Y(new_n27884_));
  AND2X1   g25448(.A(new_n26589_), .B(new_n12463_), .Y(new_n27885_));
  NOR3X1   g25449(.A(new_n27885_), .B(new_n26540_), .C(new_n12487_), .Y(new_n27886_));
  INVX1    g25450(.A(new_n27886_), .Y(new_n27887_));
  AOI21X1  g25451(.A0(new_n27887_), .A1(new_n27780_), .B0(pi1156), .Y(new_n27888_));
  OR4X1    g25452(.A(new_n26533_), .B(new_n26522_), .C(new_n26556_), .D(new_n12555_), .Y(new_n27889_));
  OAI21X1  g25453(.A0(new_n27888_), .A1(new_n27884_), .B0(new_n27889_), .Y(new_n27890_));
  AOI21X1  g25454(.A0(new_n27890_), .A1(new_n27881_), .B0(new_n23173_), .Y(new_n27891_));
  AND2X1   g25455(.A(new_n27780_), .B(new_n12555_), .Y(new_n27892_));
  NOR4X1   g25456(.A(new_n26579_), .B(new_n26526_), .C(new_n26522_), .D(new_n12463_), .Y(new_n27893_));
  OR2X1    g25457(.A(new_n27893_), .B(new_n27883_), .Y(new_n27894_));
  AND3X1   g25458(.A(new_n27894_), .B(new_n27892_), .C(new_n27887_), .Y(new_n27895_));
  OAI21X1  g25459(.A0(new_n27894_), .A1(new_n27787_), .B0(pi1156), .Y(new_n27896_));
  OAI21X1  g25460(.A0(new_n27896_), .A1(new_n27886_), .B0(new_n23173_), .Y(new_n27897_));
  OAI21X1  g25461(.A0(new_n27897_), .A1(new_n27895_), .B0(new_n8422_), .Y(new_n27898_));
  AOI21X1  g25462(.A0(new_n26536_), .A1(new_n26534_), .B0(new_n26630_), .Y(new_n27899_));
  INVX1    g25463(.A(new_n27899_), .Y(new_n27900_));
  OAI21X1  g25464(.A0(new_n27789_), .A1(new_n26531_), .B0(new_n27900_), .Y(new_n27901_));
  OAI21X1  g25465(.A0(new_n27901_), .A1(new_n26579_), .B0(new_n12555_), .Y(new_n27902_));
  OR2X1    g25466(.A(new_n27729_), .B(new_n12463_), .Y(new_n27903_));
  INVX1    g25467(.A(new_n26633_), .Y(new_n27904_));
  OAI21X1  g25468(.A0(new_n27904_), .A1(new_n26533_), .B0(new_n12463_), .Y(new_n27905_));
  AND3X1   g25469(.A(new_n27905_), .B(new_n27903_), .C(new_n12487_), .Y(new_n27906_));
  AND2X1   g25470(.A(pi1156), .B(new_n23173_), .Y(new_n27907_));
  OAI21X1  g25471(.A0(new_n27899_), .A1(new_n12487_), .B0(new_n27907_), .Y(new_n27908_));
  OR2X1    g25472(.A(new_n27908_), .B(new_n27906_), .Y(new_n27909_));
  AND2X1   g25473(.A(pi1156), .B(pi0211), .Y(new_n27910_));
  AOI21X1  g25474(.A0(new_n27901_), .A1(new_n27910_), .B0(new_n8422_), .Y(new_n27911_));
  NAND3X1  g25475(.A(new_n27911_), .B(new_n27909_), .C(new_n27902_), .Y(new_n27912_));
  AND2X1   g25476(.A(new_n27912_), .B(pi0263), .Y(new_n27913_));
  OAI21X1  g25477(.A0(new_n27898_), .A1(new_n27891_), .B0(new_n27913_), .Y(new_n27914_));
  NOR4X1   g25478(.A(new_n27558_), .B(new_n26580_), .C(pi1155), .D(pi1091), .Y(new_n27915_));
  INVX1    g25479(.A(new_n27915_), .Y(new_n27916_));
  AOI21X1  g25480(.A0(new_n27595_), .A1(pi1155), .B0(pi1154), .Y(new_n27917_));
  AOI21X1  g25481(.A0(new_n27917_), .A1(new_n27916_), .B0(pi1156), .Y(new_n27918_));
  AOI21X1  g25482(.A0(new_n26526_), .A1(new_n26507_), .B0(new_n26522_), .Y(new_n27919_));
  NOR3X1   g25483(.A(new_n27558_), .B(pi1155), .C(pi1091), .Y(new_n27920_));
  INVX1    g25484(.A(new_n27920_), .Y(new_n27921_));
  AOI21X1  g25485(.A0(new_n27625_), .A1(pi1155), .B0(new_n12487_), .Y(new_n27922_));
  AOI21X1  g25486(.A0(new_n26607_), .A1(pi1155), .B0(pi1154), .Y(new_n27923_));
  AOI22X1  g25487(.A0(new_n27923_), .A1(new_n27921_), .B0(new_n27922_), .B1(new_n27919_), .Y(new_n27924_));
  AOI22X1  g25488(.A0(new_n26551_), .A1(new_n12463_), .B0(new_n27592_), .B1(new_n26553_), .Y(new_n27925_));
  OAI21X1  g25489(.A0(new_n27925_), .A1(pi1154), .B0(pi1156), .Y(new_n27926_));
  NAND2X1  g25490(.A(new_n27922_), .B(new_n27919_), .Y(new_n27927_));
  NAND2X1  g25491(.A(new_n27923_), .B(new_n26551_), .Y(new_n27928_));
  OAI21X1  g25492(.A0(new_n27927_), .A1(new_n26524_), .B0(new_n27928_), .Y(new_n27929_));
  OAI21X1  g25493(.A0(new_n27929_), .A1(new_n27926_), .B0(new_n23173_), .Y(new_n27930_));
  AOI21X1  g25494(.A0(new_n27924_), .A1(new_n27918_), .B0(new_n27930_), .Y(new_n27931_));
  AOI21X1  g25495(.A0(new_n27922_), .A1(new_n26562_), .B0(new_n27926_), .Y(new_n27932_));
  INVX1    g25496(.A(new_n27918_), .Y(new_n27933_));
  AND2X1   g25497(.A(new_n27922_), .B(new_n27550_), .Y(new_n27934_));
  OAI21X1  g25498(.A0(new_n27934_), .A1(new_n27933_), .B0(pi0211), .Y(new_n27935_));
  OAI21X1  g25499(.A0(new_n27935_), .A1(new_n27932_), .B0(new_n8422_), .Y(new_n27936_));
  AND2X1   g25500(.A(new_n26521_), .B(pi1155), .Y(new_n27937_));
  OR3X1    g25501(.A(new_n27937_), .B(new_n26637_), .C(new_n12487_), .Y(new_n27938_));
  OAI21X1  g25502(.A0(new_n27938_), .A1(new_n26526_), .B0(new_n27928_), .Y(new_n27939_));
  NAND2X1  g25503(.A(new_n27939_), .B(new_n27910_), .Y(new_n27940_));
  NAND2X1  g25504(.A(new_n27923_), .B(new_n27921_), .Y(new_n27941_));
  AOI21X1  g25505(.A0(new_n27938_), .A1(new_n27941_), .B0(pi1156), .Y(new_n27942_));
  INVX1    g25506(.A(new_n27907_), .Y(new_n27943_));
  OR3X1    g25507(.A(new_n26579_), .B(new_n26529_), .C(pi1154), .Y(new_n27944_));
  AND2X1   g25508(.A(new_n27944_), .B(new_n26603_), .Y(new_n27945_));
  NOR3X1   g25509(.A(new_n27945_), .B(new_n27937_), .C(new_n27943_), .Y(new_n27946_));
  NOR3X1   g25510(.A(new_n27946_), .B(new_n27942_), .C(new_n8422_), .Y(new_n27947_));
  AOI21X1  g25511(.A0(new_n27947_), .A1(new_n27940_), .B0(pi0263), .Y(new_n27948_));
  OAI21X1  g25512(.A0(new_n27936_), .A1(new_n27931_), .B0(new_n27948_), .Y(new_n27949_));
  AND3X1   g25513(.A(new_n27949_), .B(new_n27914_), .C(new_n26600_), .Y(new_n27950_));
  INVX1    g25514(.A(new_n26671_), .Y(new_n27951_));
  AOI21X1  g25515(.A0(new_n25130_), .A1(new_n2933_), .B0(new_n12463_), .Y(new_n27952_));
  NAND2X1  g25516(.A(new_n27811_), .B(new_n12487_), .Y(new_n27953_));
  OAI21X1  g25517(.A0(new_n27952_), .A1(new_n27951_), .B0(new_n27953_), .Y(new_n27954_));
  OR2X1    g25518(.A(new_n27954_), .B(new_n26684_), .Y(new_n27955_));
  AND2X1   g25519(.A(new_n27955_), .B(new_n27910_), .Y(new_n27956_));
  OR2X1    g25520(.A(new_n12463_), .B(pi0199), .Y(new_n27957_));
  AOI21X1  g25521(.A0(new_n27957_), .A1(new_n24946_), .B0(new_n12487_), .Y(new_n27958_));
  NOR3X1   g25522(.A(new_n27958_), .B(new_n27943_), .C(new_n2702_), .Y(new_n27959_));
  OAI21X1  g25523(.A0(new_n24975_), .A1(pi1154), .B0(new_n27959_), .Y(new_n27960_));
  NOR2X1   g25524(.A(new_n27818_), .B(new_n26650_), .Y(new_n27961_));
  NOR3X1   g25525(.A(new_n27961_), .B(new_n24922_), .C(pi1156), .Y(new_n27962_));
  NOR2X1   g25526(.A(new_n27962_), .B(new_n8422_), .Y(new_n27963_));
  AND2X1   g25527(.A(new_n27963_), .B(new_n27960_), .Y(new_n27964_));
  INVX1    g25528(.A(new_n27964_), .Y(new_n27965_));
  OAI21X1  g25529(.A0(new_n25313_), .A1(new_n24917_), .B0(new_n27648_), .Y(new_n27966_));
  NOR2X1   g25530(.A(new_n27966_), .B(new_n25341_), .Y(new_n27967_));
  AOI21X1  g25531(.A0(new_n27954_), .A1(new_n23173_), .B0(new_n27967_), .Y(new_n27968_));
  NOR2X1   g25532(.A(new_n27968_), .B(new_n12555_), .Y(new_n27969_));
  NOR3X1   g25533(.A(new_n27961_), .B(new_n25341_), .C(new_n23173_), .Y(new_n27970_));
  NOR2X1   g25534(.A(new_n25228_), .B(new_n24922_), .Y(new_n27971_));
  AOI21X1  g25535(.A0(new_n27971_), .A1(new_n27746_), .B0(new_n27970_), .Y(new_n27972_));
  OAI21X1  g25536(.A0(new_n27972_), .A1(pi1156), .B0(new_n8422_), .Y(new_n27973_));
  OAI22X1  g25537(.A0(new_n27973_), .A1(new_n27969_), .B0(new_n27965_), .B1(new_n27956_), .Y(new_n27974_));
  NOR3X1   g25538(.A(new_n25061_), .B(new_n24975_), .C(pi1154), .Y(new_n27975_));
  AOI21X1  g25539(.A0(new_n24951_), .A1(pi1155), .B0(new_n24916_), .Y(new_n27976_));
  OAI21X1  g25540(.A0(new_n27976_), .A1(new_n12487_), .B0(pi1156), .Y(new_n27977_));
  NOR3X1   g25541(.A(new_n27961_), .B(new_n25341_), .C(pi1156), .Y(new_n27978_));
  NOR2X1   g25542(.A(new_n27978_), .B(new_n23173_), .Y(new_n27979_));
  OAI21X1  g25543(.A0(new_n27977_), .A1(new_n27975_), .B0(new_n27979_), .Y(new_n27980_));
  AND2X1   g25544(.A(new_n12463_), .B(pi0200), .Y(new_n27981_));
  OAI22X1  g25545(.A0(new_n25589_), .A1(new_n27981_), .B0(new_n9445_), .B1(new_n12487_), .Y(new_n27982_));
  AOI21X1  g25546(.A0(new_n27982_), .A1(new_n23173_), .B0(pi0219), .Y(new_n27983_));
  AND2X1   g25547(.A(new_n27983_), .B(new_n27980_), .Y(new_n27984_));
  AOI21X1  g25548(.A0(new_n24925_), .A1(pi1154), .B0(new_n12555_), .Y(new_n27985_));
  NOR2X1   g25549(.A(new_n27985_), .B(pi0299), .Y(new_n27986_));
  AND3X1   g25550(.A(new_n24925_), .B(new_n9445_), .C(new_n12487_), .Y(new_n27987_));
  NOR3X1   g25551(.A(new_n27987_), .B(new_n27986_), .C(new_n25833_), .Y(new_n27988_));
  NOR2X1   g25552(.A(new_n27988_), .B(new_n12555_), .Y(new_n27989_));
  NOR3X1   g25553(.A(new_n27985_), .B(new_n27971_), .C(pi0299), .Y(new_n27990_));
  NOR3X1   g25554(.A(new_n27990_), .B(new_n27989_), .C(new_n8422_), .Y(new_n27991_));
  NOR4X1   g25555(.A(new_n27991_), .B(new_n27984_), .C(new_n2702_), .D(new_n26599_), .Y(new_n27992_));
  AOI21X1  g25556(.A0(new_n27974_), .A1(new_n26599_), .B0(new_n27992_), .Y(new_n27993_));
  OAI21X1  g25557(.A0(new_n27993_), .A1(new_n26600_), .B0(new_n6489_), .Y(new_n27994_));
  NAND2X1  g25558(.A(pi1155), .B(pi0211), .Y(new_n27995_));
  OAI21X1  g25559(.A0(new_n27818_), .A1(pi0211), .B0(new_n27995_), .Y(new_n27996_));
  AOI21X1  g25560(.A0(new_n26505_), .A1(pi0211), .B0(new_n27996_), .Y(new_n27997_));
  OAI21X1  g25561(.A0(new_n27997_), .A1(new_n26514_), .B0(new_n8422_), .Y(new_n27998_));
  AND3X1   g25562(.A(new_n27998_), .B(new_n27756_), .C(new_n26599_), .Y(new_n27999_));
  INVX1    g25563(.A(new_n27579_), .Y(new_n28000_));
  AOI22X1  g25564(.A0(new_n27746_), .A1(pi1154), .B0(pi1155), .B1(pi0211), .Y(new_n28001_));
  AOI21X1  g25565(.A0(new_n26505_), .A1(pi0211), .B0(new_n28001_), .Y(new_n28002_));
  OR2X1    g25566(.A(new_n28002_), .B(new_n28000_), .Y(new_n28003_));
  AND3X1   g25567(.A(new_n28003_), .B(new_n27578_), .C(pi0263), .Y(new_n28004_));
  INVX1    g25568(.A(new_n26600_), .Y(new_n28005_));
  AOI21X1  g25569(.A0(pi1156), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n28006_));
  AOI21X1  g25570(.A0(new_n28006_), .A1(pi1091), .B0(new_n28005_), .Y(new_n28007_));
  OAI21X1  g25571(.A0(new_n28004_), .A1(new_n27999_), .B0(new_n28007_), .Y(new_n28008_));
  AOI21X1  g25572(.A0(pi1155), .A1(pi0211), .B0(pi0219), .Y(new_n28009_));
  AOI21X1  g25573(.A0(new_n28009_), .A1(new_n27727_), .B0(new_n28006_), .Y(new_n28010_));
  MX2X1    g25574(.A(new_n28010_), .B(new_n26599_), .S0(new_n2702_), .Y(new_n28011_));
  AOI21X1  g25575(.A0(new_n28011_), .A1(new_n28005_), .B0(new_n6489_), .Y(new_n28012_));
  AOI21X1  g25576(.A0(new_n28012_), .A1(new_n28008_), .B0(new_n27711_), .Y(new_n28013_));
  OAI21X1  g25577(.A0(new_n27994_), .A1(new_n27950_), .B0(new_n28013_), .Y(new_n28014_));
  OAI21X1  g25578(.A0(new_n28011_), .A1(new_n6489_), .B0(new_n27711_), .Y(new_n28015_));
  AOI21X1  g25579(.A0(new_n27993_), .A1(new_n6489_), .B0(new_n28015_), .Y(new_n28016_));
  NOR2X1   g25580(.A(new_n28016_), .B(pi0230), .Y(new_n28017_));
  INVX1    g25581(.A(new_n27983_), .Y(new_n28018_));
  OR3X1    g25582(.A(pi1154), .B(pi0200), .C(pi0199), .Y(new_n28019_));
  OAI21X1  g25583(.A0(new_n24927_), .A1(new_n24923_), .B0(new_n12555_), .Y(new_n28020_));
  NAND4X1  g25584(.A(new_n28020_), .B(new_n28019_), .C(new_n24925_), .D(new_n2933_), .Y(new_n28021_));
  AOI21X1  g25585(.A0(new_n28021_), .A1(new_n24955_), .B0(new_n23173_), .Y(new_n28022_));
  AOI21X1  g25586(.A0(new_n25833_), .A1(pi1156), .B0(new_n8422_), .Y(new_n28023_));
  AOI21X1  g25587(.A0(new_n28023_), .A1(new_n28021_), .B0(po1038), .Y(new_n28024_));
  OAI21X1  g25588(.A0(new_n28022_), .A1(new_n28018_), .B0(new_n28024_), .Y(new_n28025_));
  AOI21X1  g25589(.A0(new_n28010_), .A1(po1038), .B0(new_n24814_), .Y(new_n28026_));
  AOI22X1  g25590(.A0(new_n28026_), .A1(new_n28025_), .B0(new_n28017_), .B1(new_n28014_), .Y(po0420));
  AND2X1   g25591(.A(new_n26508_), .B(pi0314), .Y(new_n28028_));
  INVX1    g25592(.A(new_n28028_), .Y(new_n28029_));
  AOI21X1  g25593(.A0(new_n28029_), .A1(pi0264), .B0(pi1091), .Y(new_n28030_));
  OAI21X1  g25594(.A0(new_n28029_), .A1(pi0796), .B0(new_n28030_), .Y(new_n28031_));
  NAND2X1  g25595(.A(pi1141), .B(pi1091), .Y(new_n28032_));
  AOI21X1  g25596(.A0(new_n28032_), .A1(new_n28031_), .B0(pi0200), .Y(new_n28033_));
  AND2X1   g25597(.A(pi1142), .B(pi1091), .Y(new_n28034_));
  INVX1    g25598(.A(new_n28034_), .Y(new_n28035_));
  AOI21X1  g25599(.A0(new_n28035_), .A1(new_n28031_), .B0(new_n7937_), .Y(new_n28036_));
  OR3X1    g25600(.A(new_n28036_), .B(new_n28033_), .C(pi0199), .Y(new_n28037_));
  INVX1    g25601(.A(new_n26501_), .Y(new_n28038_));
  AOI21X1  g25602(.A0(new_n28038_), .A1(pi0264), .B0(pi1091), .Y(new_n28039_));
  OAI21X1  g25603(.A0(new_n28038_), .A1(pi0796), .B0(new_n28039_), .Y(new_n28040_));
  AND2X1   g25604(.A(pi1143), .B(pi1091), .Y(new_n28041_));
  AOI21X1  g25605(.A0(new_n28041_), .A1(new_n7937_), .B0(new_n7871_), .Y(new_n28042_));
  AOI21X1  g25606(.A0(new_n28042_), .A1(new_n28040_), .B0(new_n22572_), .Y(new_n28043_));
  AOI21X1  g25607(.A0(new_n28032_), .A1(new_n28031_), .B0(pi0211), .Y(new_n28044_));
  AOI21X1  g25608(.A0(new_n28035_), .A1(new_n28031_), .B0(new_n23173_), .Y(new_n28045_));
  OR3X1    g25609(.A(new_n28045_), .B(new_n28044_), .C(pi0219), .Y(new_n28046_));
  AOI21X1  g25610(.A0(new_n27746_), .A1(new_n24826_), .B0(new_n8422_), .Y(new_n28047_));
  AOI21X1  g25611(.A0(new_n28047_), .A1(new_n28040_), .B0(new_n11660_), .Y(new_n28048_));
  AOI22X1  g25612(.A0(new_n28048_), .A1(new_n28046_), .B0(new_n28043_), .B1(new_n28037_), .Y(new_n28049_));
  AOI21X1  g25613(.A0(pi1142), .A1(pi0211), .B0(pi0219), .Y(new_n28050_));
  OAI21X1  g25614(.A0(new_n3759_), .A1(pi0211), .B0(new_n28050_), .Y(new_n28051_));
  AOI21X1  g25615(.A0(new_n28051_), .A1(new_n25511_), .B0(new_n11660_), .Y(new_n28052_));
  OR2X1    g25616(.A(new_n3759_), .B(pi0199), .Y(new_n28053_));
  AOI21X1  g25617(.A0(new_n28053_), .A1(new_n25494_), .B0(new_n24841_), .Y(new_n28054_));
  OAI21X1  g25618(.A0(new_n28054_), .A1(new_n22572_), .B0(pi0230), .Y(new_n28055_));
  OAI22X1  g25619(.A0(new_n28055_), .A1(new_n28052_), .B0(new_n28049_), .B1(pi0230), .Y(po0421));
  AOI21X1  g25620(.A0(new_n28029_), .A1(pi0265), .B0(pi1091), .Y(new_n28057_));
  OAI21X1  g25621(.A0(new_n28029_), .A1(pi0819), .B0(new_n28057_), .Y(new_n28058_));
  AOI21X1  g25622(.A0(new_n28058_), .A1(new_n28035_), .B0(pi0200), .Y(new_n28059_));
  INVX1    g25623(.A(new_n28041_), .Y(new_n28060_));
  AOI21X1  g25624(.A0(new_n28058_), .A1(new_n28060_), .B0(new_n7937_), .Y(new_n28061_));
  OR3X1    g25625(.A(new_n28061_), .B(new_n28059_), .C(pi0199), .Y(new_n28062_));
  AOI21X1  g25626(.A0(new_n28038_), .A1(pi0265), .B0(pi1091), .Y(new_n28063_));
  OAI21X1  g25627(.A0(new_n28038_), .A1(pi0819), .B0(new_n28063_), .Y(new_n28064_));
  AND2X1   g25628(.A(pi1144), .B(pi1091), .Y(new_n28065_));
  AOI21X1  g25629(.A0(new_n28065_), .A1(new_n7937_), .B0(new_n7871_), .Y(new_n28066_));
  AOI21X1  g25630(.A0(new_n28066_), .A1(new_n28064_), .B0(new_n22572_), .Y(new_n28067_));
  AOI21X1  g25631(.A0(new_n28058_), .A1(new_n28035_), .B0(pi0211), .Y(new_n28068_));
  AOI21X1  g25632(.A0(new_n28058_), .A1(new_n28060_), .B0(new_n23173_), .Y(new_n28069_));
  OR3X1    g25633(.A(new_n28069_), .B(new_n28068_), .C(pi0219), .Y(new_n28070_));
  AOI21X1  g25634(.A0(pi1091), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n28071_));
  OR2X1    g25635(.A(new_n28071_), .B(new_n26450_), .Y(new_n28072_));
  AOI21X1  g25636(.A0(new_n28072_), .A1(new_n28064_), .B0(new_n11660_), .Y(new_n28073_));
  AOI22X1  g25637(.A0(new_n28073_), .A1(new_n28070_), .B0(new_n28067_), .B1(new_n28062_), .Y(new_n28074_));
  INVX1    g25638(.A(new_n26450_), .Y(new_n28075_));
  AOI21X1  g25639(.A0(pi1143), .A1(pi0211), .B0(pi0219), .Y(new_n28076_));
  OAI21X1  g25640(.A0(new_n24820_), .A1(pi0211), .B0(new_n28076_), .Y(new_n28077_));
  AOI21X1  g25641(.A0(new_n28077_), .A1(new_n28075_), .B0(new_n11660_), .Y(new_n28078_));
  OR2X1    g25642(.A(new_n24820_), .B(pi0199), .Y(new_n28079_));
  AOI21X1  g25643(.A0(new_n26453_), .A1(new_n28079_), .B0(new_n24834_), .Y(new_n28080_));
  OAI21X1  g25644(.A0(new_n28080_), .A1(new_n22572_), .B0(pi0230), .Y(new_n28081_));
  OAI22X1  g25645(.A0(new_n28081_), .A1(new_n28078_), .B0(new_n28074_), .B1(pi0230), .Y(po0422));
  AOI21X1  g25646(.A0(pi1136), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n28083_));
  AND2X1   g25647(.A(new_n4622_), .B(pi0211), .Y(new_n28084_));
  OR3X1    g25648(.A(new_n28084_), .B(new_n28083_), .C(new_n7997_), .Y(new_n28085_));
  AOI21X1  g25649(.A0(pi1135), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n28086_));
  AOI21X1  g25650(.A0(pi1136), .A1(pi0199), .B0(pi0200), .Y(new_n28087_));
  OR2X1    g25651(.A(new_n28087_), .B(pi0299), .Y(new_n28088_));
  OAI22X1  g25652(.A0(new_n28088_), .A1(new_n28086_), .B0(new_n28085_), .B1(new_n2933_), .Y(new_n28089_));
  OAI21X1  g25653(.A0(new_n28085_), .A1(new_n6489_), .B0(pi0230), .Y(new_n28090_));
  AOI21X1  g25654(.A0(new_n28089_), .A1(new_n6489_), .B0(new_n28090_), .Y(new_n28091_));
  OAI21X1  g25655(.A0(new_n28029_), .A1(pi0948), .B0(new_n2702_), .Y(new_n28092_));
  AOI21X1  g25656(.A0(new_n28029_), .A1(new_n4470_), .B0(new_n28092_), .Y(new_n28093_));
  AND2X1   g25657(.A(pi1136), .B(pi1091), .Y(new_n28094_));
  NOR2X1   g25658(.A(new_n26501_), .B(pi0266), .Y(new_n28095_));
  OAI21X1  g25659(.A0(new_n28038_), .A1(pi0948), .B0(new_n2702_), .Y(new_n28096_));
  OAI21X1  g25660(.A0(new_n28096_), .A1(new_n28095_), .B0(pi0199), .Y(new_n28097_));
  OAI22X1  g25661(.A0(new_n28097_), .A1(new_n28094_), .B0(new_n28093_), .B1(pi0199), .Y(new_n28098_));
  NOR2X1   g25662(.A(new_n28098_), .B(pi0200), .Y(new_n28099_));
  AND2X1   g25663(.A(pi1135), .B(pi1091), .Y(new_n28100_));
  OR3X1    g25664(.A(new_n28100_), .B(new_n28093_), .C(pi0199), .Y(new_n28101_));
  AND3X1   g25665(.A(new_n28101_), .B(new_n28097_), .C(pi0200), .Y(new_n28102_));
  OAI21X1  g25666(.A0(new_n28102_), .A1(new_n28099_), .B0(new_n11660_), .Y(new_n28103_));
  OAI22X1  g25667(.A0(new_n28096_), .A1(new_n28095_), .B0(new_n28083_), .B1(new_n28071_), .Y(new_n28104_));
  AND2X1   g25668(.A(new_n28104_), .B(new_n22572_), .Y(new_n28105_));
  NOR2X1   g25669(.A(new_n28093_), .B(pi0219), .Y(new_n28106_));
  OAI21X1  g25670(.A0(new_n27649_), .A1(new_n4622_), .B0(new_n28106_), .Y(new_n28107_));
  AOI21X1  g25671(.A0(new_n28107_), .A1(new_n28105_), .B0(pi0230), .Y(new_n28108_));
  AOI21X1  g25672(.A0(new_n28108_), .A1(new_n28103_), .B0(new_n28091_), .Y(new_n28109_));
  AND3X1   g25673(.A(new_n4554_), .B(new_n7937_), .C(pi0199), .Y(new_n28110_));
  OR3X1    g25674(.A(new_n28110_), .B(new_n28086_), .C(new_n22572_), .Y(new_n28111_));
  OR3X1    g25675(.A(new_n28084_), .B(new_n28083_), .C(new_n11660_), .Y(new_n28112_));
  AND2X1   g25676(.A(new_n28112_), .B(pi0230), .Y(new_n28113_));
  OR2X1    g25677(.A(new_n2702_), .B(pi0199), .Y(new_n28114_));
  AOI21X1  g25678(.A0(new_n28114_), .A1(new_n28098_), .B0(pi0200), .Y(new_n28115_));
  OAI21X1  g25679(.A0(new_n28115_), .A1(new_n28102_), .B0(new_n11660_), .Y(new_n28116_));
  OAI21X1  g25680(.A0(new_n28084_), .A1(new_n2702_), .B0(new_n28106_), .Y(new_n28117_));
  AOI21X1  g25681(.A0(new_n28117_), .A1(new_n28105_), .B0(pi0230), .Y(new_n28118_));
  AOI22X1  g25682(.A0(new_n28118_), .A1(new_n28116_), .B0(new_n28113_), .B1(new_n28111_), .Y(new_n28119_));
  MX2X1    g25683(.A(new_n28119_), .B(new_n28109_), .S0(new_n4747_), .Y(po0423));
  AND2X1   g25684(.A(pi0254), .B(pi0253), .Y(new_n28121_));
  INVX1    g25685(.A(new_n28121_), .Y(new_n28122_));
  NOR4X1   g25686(.A(new_n27732_), .B(new_n26579_), .C(new_n26533_), .D(new_n26529_), .Y(new_n28123_));
  NOR3X1   g25687(.A(new_n28123_), .B(new_n26626_), .C(pi1154), .Y(new_n28124_));
  NOR4X1   g25688(.A(new_n27736_), .B(new_n26531_), .C(new_n12463_), .D(new_n12487_), .Y(new_n28125_));
  OAI21X1  g25689(.A0(new_n28125_), .A1(new_n28124_), .B0(pi0211), .Y(new_n28126_));
  INVX1    g25690(.A(pi0267), .Y(new_n28127_));
  NOR3X1   g25691(.A(new_n26535_), .B(new_n26533_), .C(new_n12364_), .Y(new_n28128_));
  AND2X1   g25692(.A(pi1155), .B(new_n23173_), .Y(new_n28129_));
  OAI21X1  g25693(.A0(new_n27904_), .A1(new_n26533_), .B0(new_n28129_), .Y(new_n28130_));
  OR3X1    g25694(.A(new_n28130_), .B(new_n28128_), .C(new_n27718_), .Y(new_n28131_));
  NOR4X1   g25695(.A(new_n26579_), .B(new_n26529_), .C(new_n26526_), .D(new_n12487_), .Y(new_n28132_));
  OR3X1    g25696(.A(new_n28132_), .B(new_n28123_), .C(pi1155), .Y(new_n28133_));
  AND3X1   g25697(.A(new_n28133_), .B(new_n28131_), .C(new_n28127_), .Y(new_n28134_));
  AOI21X1  g25698(.A0(new_n27566_), .A1(new_n27551_), .B0(new_n26607_), .Y(new_n28135_));
  NOR2X1   g25699(.A(new_n28135_), .B(new_n12487_), .Y(new_n28136_));
  OAI21X1  g25700(.A0(new_n26535_), .A1(new_n26527_), .B0(new_n12487_), .Y(new_n28137_));
  OAI21X1  g25701(.A0(new_n28137_), .A1(new_n27631_), .B0(new_n12463_), .Y(new_n28138_));
  OR2X1    g25702(.A(new_n28138_), .B(new_n28136_), .Y(new_n28139_));
  OR2X1    g25703(.A(new_n27630_), .B(new_n27629_), .Y(new_n28140_));
  OAI21X1  g25704(.A0(new_n26562_), .A1(new_n12364_), .B0(pi1155), .Y(new_n28141_));
  AOI21X1  g25705(.A0(new_n27944_), .A1(new_n26521_), .B0(new_n28141_), .Y(new_n28142_));
  AOI21X1  g25706(.A0(new_n28142_), .A1(new_n28140_), .B0(new_n28127_), .Y(new_n28143_));
  AOI22X1  g25707(.A0(new_n28143_), .A1(new_n28139_), .B0(new_n28134_), .B1(new_n28126_), .Y(new_n28144_));
  OR2X1    g25708(.A(new_n28144_), .B(new_n8422_), .Y(new_n28145_));
  INVX1    g25709(.A(new_n26561_), .Y(new_n28146_));
  NOR2X1   g25710(.A(new_n28135_), .B(new_n27595_), .Y(new_n28147_));
  OAI21X1  g25711(.A0(new_n28147_), .A1(new_n27903_), .B0(pi1154), .Y(new_n28148_));
  AOI21X1  g25712(.A0(new_n27548_), .A1(new_n12487_), .B0(new_n12463_), .Y(new_n28149_));
  OAI21X1  g25713(.A0(new_n28149_), .A1(new_n28146_), .B0(new_n28148_), .Y(new_n28150_));
  OR3X1    g25714(.A(new_n28123_), .B(new_n27882_), .C(pi1155), .Y(new_n28151_));
  AND3X1   g25715(.A(new_n28151_), .B(new_n28150_), .C(pi0211), .Y(new_n28152_));
  OAI21X1  g25716(.A0(new_n26580_), .A1(new_n12364_), .B0(new_n12463_), .Y(new_n28153_));
  OR3X1    g25717(.A(new_n28153_), .B(new_n27626_), .C(new_n26533_), .Y(new_n28154_));
  OAI21X1  g25718(.A0(new_n28128_), .A1(new_n27787_), .B0(pi1155), .Y(new_n28155_));
  AND3X1   g25719(.A(new_n28155_), .B(new_n28154_), .C(new_n12487_), .Y(new_n28156_));
  INVX1    g25720(.A(new_n28155_), .Y(new_n28157_));
  OR3X1    g25721(.A(new_n26579_), .B(new_n26526_), .C(new_n26522_), .Y(new_n28158_));
  AND2X1   g25722(.A(new_n28158_), .B(new_n12364_), .Y(new_n28159_));
  NOR2X1   g25723(.A(new_n27893_), .B(new_n12487_), .Y(new_n28160_));
  OAI21X1  g25724(.A0(new_n28159_), .A1(new_n28153_), .B0(new_n28160_), .Y(new_n28161_));
  OAI21X1  g25725(.A0(new_n28161_), .A1(new_n28157_), .B0(new_n23173_), .Y(new_n28162_));
  OAI21X1  g25726(.A0(new_n28162_), .A1(new_n28156_), .B0(new_n28127_), .Y(new_n28163_));
  AND2X1   g25727(.A(new_n26589_), .B(new_n12364_), .Y(new_n28164_));
  OR2X1    g25728(.A(new_n28164_), .B(new_n26582_), .Y(new_n28165_));
  NOR3X1   g25729(.A(new_n26522_), .B(new_n26521_), .C(pi1155), .Y(new_n28166_));
  OR3X1    g25730(.A(new_n26544_), .B(new_n26522_), .C(new_n26521_), .Y(new_n28167_));
  OAI21X1  g25731(.A0(new_n28141_), .A1(new_n28167_), .B0(pi1154), .Y(new_n28168_));
  AOI21X1  g25732(.A0(new_n28166_), .A1(new_n28165_), .B0(new_n28168_), .Y(new_n28169_));
  OR3X1    g25733(.A(new_n27565_), .B(new_n27919_), .C(pi1154), .Y(new_n28170_));
  AND2X1   g25734(.A(new_n28170_), .B(new_n12463_), .Y(new_n28171_));
  NOR4X1   g25735(.A(new_n28171_), .B(new_n27565_), .C(new_n26562_), .D(pi1154), .Y(new_n28172_));
  OAI21X1  g25736(.A0(new_n28172_), .A1(new_n28169_), .B0(pi0211), .Y(new_n28173_));
  OAI21X1  g25737(.A0(new_n28165_), .A1(new_n12487_), .B0(new_n28171_), .Y(new_n28174_));
  OR2X1    g25738(.A(new_n27776_), .B(new_n26541_), .Y(new_n28175_));
  AOI21X1  g25739(.A0(new_n26521_), .A1(pi1154), .B0(new_n12463_), .Y(new_n28176_));
  AOI21X1  g25740(.A0(new_n28176_), .A1(new_n28175_), .B0(pi0211), .Y(new_n28177_));
  AOI21X1  g25741(.A0(new_n28177_), .A1(new_n28174_), .B0(new_n28127_), .Y(new_n28178_));
  AOI21X1  g25742(.A0(new_n28178_), .A1(new_n28173_), .B0(pi0219), .Y(new_n28179_));
  OAI21X1  g25743(.A0(new_n28163_), .A1(new_n28152_), .B0(new_n28179_), .Y(new_n28180_));
  AOI21X1  g25744(.A0(new_n28180_), .A1(new_n28145_), .B0(new_n28122_), .Y(new_n28181_));
  AOI21X1  g25745(.A0(new_n27951_), .A1(pi1153), .B0(new_n12463_), .Y(new_n28182_));
  OAI21X1  g25746(.A0(new_n27809_), .A1(pi1153), .B0(new_n28182_), .Y(new_n28183_));
  OAI21X1  g25747(.A0(new_n9445_), .A1(new_n12364_), .B0(new_n12463_), .Y(new_n28184_));
  OR2X1    g25748(.A(new_n28184_), .B(new_n2702_), .Y(new_n28185_));
  AOI21X1  g25749(.A0(new_n28185_), .A1(new_n28183_), .B0(pi1154), .Y(new_n28186_));
  NOR2X1   g25750(.A(new_n27741_), .B(pi1155), .Y(new_n28187_));
  AOI22X1  g25751(.A0(new_n28187_), .A1(new_n27659_), .B0(new_n28182_), .B1(new_n27811_), .Y(new_n28188_));
  OAI21X1  g25752(.A0(new_n28188_), .A1(new_n12487_), .B0(new_n8422_), .Y(new_n28189_));
  NOR4X1   g25753(.A(new_n27640_), .B(new_n25549_), .C(new_n12463_), .D(new_n2702_), .Y(new_n28190_));
  NOR3X1   g25754(.A(new_n25197_), .B(pi0299), .C(pi0199), .Y(new_n28191_));
  NOR4X1   g25755(.A(new_n28191_), .B(new_n28190_), .C(new_n12487_), .D(new_n2702_), .Y(new_n28192_));
  NAND2X1  g25756(.A(new_n25204_), .B(pi1153), .Y(new_n28193_));
  AND2X1   g25757(.A(new_n28193_), .B(new_n27818_), .Y(new_n28194_));
  OAI21X1  g25758(.A0(new_n25659_), .A1(new_n12463_), .B0(new_n28194_), .Y(new_n28195_));
  NAND2X1  g25759(.A(new_n28195_), .B(pi0219), .Y(new_n28196_));
  OAI22X1  g25760(.A0(new_n28196_), .A1(new_n28192_), .B0(new_n28189_), .B1(new_n28186_), .Y(new_n28197_));
  MX2X1    g25761(.A(new_n25199_), .B(new_n24970_), .S0(pi1155), .Y(new_n28198_));
  OR2X1    g25762(.A(new_n28198_), .B(new_n9447_), .Y(new_n28199_));
  NAND3X1  g25763(.A(new_n25212_), .B(new_n24907_), .C(pi1155), .Y(new_n28200_));
  AND3X1   g25764(.A(new_n28200_), .B(pi1154), .C(pi1091), .Y(new_n28201_));
  INVX1    g25765(.A(new_n28194_), .Y(new_n28202_));
  AOI21X1  g25766(.A0(new_n24992_), .A1(new_n12463_), .B0(new_n27809_), .Y(new_n28203_));
  OAI21X1  g25767(.A0(new_n28203_), .A1(new_n28202_), .B0(pi0211), .Y(new_n28204_));
  AOI21X1  g25768(.A0(new_n28201_), .A1(new_n28199_), .B0(new_n28204_), .Y(new_n28205_));
  AOI21X1  g25769(.A0(new_n28197_), .A1(new_n23173_), .B0(new_n28205_), .Y(new_n28206_));
  NOR3X1   g25770(.A(new_n25199_), .B(pi1155), .C(new_n2702_), .Y(new_n28207_));
  NOR3X1   g25771(.A(new_n28207_), .B(new_n28190_), .C(new_n27698_), .Y(new_n28208_));
  AND3X1   g25772(.A(new_n12487_), .B(new_n2933_), .C(pi0200), .Y(new_n28209_));
  NOR3X1   g25773(.A(new_n28209_), .B(new_n24982_), .C(new_n25241_), .Y(new_n28210_));
  AOI21X1  g25774(.A0(new_n28210_), .A1(pi1091), .B0(pi0211), .Y(new_n28211_));
  NOR3X1   g25775(.A(new_n28211_), .B(new_n28208_), .C(pi0219), .Y(new_n28212_));
  AND3X1   g25776(.A(new_n28191_), .B(new_n12463_), .C(pi1091), .Y(new_n28213_));
  OR3X1    g25777(.A(new_n28213_), .B(new_n28190_), .C(new_n12487_), .Y(new_n28214_));
  NAND3X1  g25778(.A(new_n28200_), .B(new_n27952_), .C(pi1154), .Y(new_n28215_));
  AOI21X1  g25779(.A0(new_n28215_), .A1(new_n28214_), .B0(new_n23173_), .Y(new_n28216_));
  OAI21X1  g25780(.A0(new_n24961_), .A1(pi1155), .B0(new_n27818_), .Y(new_n28217_));
  OAI21X1  g25781(.A0(new_n28217_), .A1(new_n25659_), .B0(new_n23173_), .Y(new_n28218_));
  AOI21X1  g25782(.A0(new_n28214_), .A1(pi1154), .B0(new_n28218_), .Y(new_n28219_));
  NOR3X1   g25783(.A(new_n28219_), .B(new_n28216_), .C(new_n8422_), .Y(new_n28220_));
  AND2X1   g25784(.A(new_n27764_), .B(new_n24916_), .Y(new_n28221_));
  OAI21X1  g25785(.A0(new_n28221_), .A1(new_n27794_), .B0(new_n28184_), .Y(new_n28222_));
  AND2X1   g25786(.A(new_n12487_), .B(pi0211), .Y(new_n28223_));
  AOI21X1  g25787(.A0(new_n28223_), .A1(new_n28222_), .B0(pi0267), .Y(new_n28224_));
  OAI21X1  g25788(.A0(new_n28220_), .A1(new_n28212_), .B0(new_n28224_), .Y(new_n28225_));
  OAI21X1  g25789(.A0(new_n28206_), .A1(new_n28127_), .B0(new_n28225_), .Y(new_n28226_));
  AND2X1   g25790(.A(new_n28226_), .B(new_n28122_), .Y(new_n28227_));
  OR2X1    g25791(.A(new_n28227_), .B(po1038), .Y(new_n28228_));
  AND3X1   g25792(.A(new_n27758_), .B(new_n27756_), .C(pi0267), .Y(new_n28229_));
  INVX1    g25793(.A(new_n26516_), .Y(new_n28230_));
  OAI21X1  g25794(.A0(new_n28230_), .A1(pi1091), .B0(new_n28127_), .Y(new_n28231_));
  OAI21X1  g25795(.A0(new_n28231_), .A1(new_n27763_), .B0(new_n28121_), .Y(new_n28232_));
  NAND2X1  g25796(.A(new_n27698_), .B(new_n8422_), .Y(new_n28233_));
  OAI22X1  g25797(.A0(new_n28233_), .A1(new_n24878_), .B0(new_n28129_), .B1(new_n8422_), .Y(new_n28234_));
  NOR3X1   g25798(.A(new_n28121_), .B(pi1091), .C(pi0267), .Y(new_n28235_));
  AOI21X1  g25799(.A0(new_n28234_), .A1(pi1091), .B0(new_n28235_), .Y(new_n28236_));
  OAI21X1  g25800(.A0(new_n28232_), .A1(new_n28229_), .B0(new_n28236_), .Y(new_n28237_));
  AOI21X1  g25801(.A0(new_n28237_), .A1(po1038), .B0(new_n27711_), .Y(new_n28238_));
  OAI21X1  g25802(.A0(new_n28228_), .A1(new_n28181_), .B0(new_n28238_), .Y(new_n28239_));
  MX2X1    g25803(.A(new_n28234_), .B(new_n28127_), .S0(new_n2702_), .Y(new_n28240_));
  AOI21X1  g25804(.A0(new_n28240_), .A1(po1038), .B0(new_n26711_), .Y(new_n28241_));
  OAI21X1  g25805(.A0(new_n28226_), .A1(po1038), .B0(new_n28241_), .Y(new_n28242_));
  AND2X1   g25806(.A(new_n28242_), .B(new_n24814_), .Y(new_n28243_));
  AOI21X1  g25807(.A0(new_n25212_), .A1(new_n24907_), .B0(new_n8422_), .Y(new_n28244_));
  OAI21X1  g25808(.A0(new_n28193_), .A1(pi1155), .B0(new_n12487_), .Y(new_n28245_));
  NOR4X1   g25809(.A(new_n25207_), .B(new_n12463_), .C(pi0299), .D(pi0200), .Y(new_n28246_));
  AOI21X1  g25810(.A0(new_n28245_), .A1(new_n25726_), .B0(new_n28246_), .Y(new_n28247_));
  OAI21X1  g25811(.A0(new_n28247_), .A1(new_n28244_), .B0(pi0211), .Y(new_n28248_));
  AOI21X1  g25812(.A0(pi1154), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n28249_));
  OAI21X1  g25813(.A0(new_n8423_), .A1(pi1155), .B0(new_n25212_), .Y(new_n28250_));
  OAI21X1  g25814(.A0(new_n28250_), .A1(new_n28249_), .B0(new_n24955_), .Y(new_n28251_));
  NAND2X1  g25815(.A(new_n28251_), .B(pi0219), .Y(new_n28252_));
  AOI21X1  g25816(.A0(new_n28210_), .A1(new_n8422_), .B0(pi0211), .Y(new_n28253_));
  AOI21X1  g25817(.A0(new_n28253_), .A1(new_n28252_), .B0(po1038), .Y(new_n28254_));
  OAI21X1  g25818(.A0(new_n28234_), .A1(new_n6489_), .B0(pi0230), .Y(new_n28255_));
  AOI21X1  g25819(.A0(new_n28254_), .A1(new_n28248_), .B0(new_n28255_), .Y(new_n28256_));
  AOI21X1  g25820(.A0(new_n28243_), .A1(new_n28239_), .B0(new_n28256_), .Y(po0424));
  INVX1    g25821(.A(new_n26710_), .Y(new_n28258_));
  INVX1    g25822(.A(new_n26527_), .Y(new_n28259_));
  OAI21X1  g25823(.A0(new_n27561_), .A1(new_n27560_), .B0(pi0219), .Y(new_n28260_));
  INVX1    g25824(.A(new_n28260_), .Y(new_n28261_));
  AOI22X1  g25825(.A0(new_n28261_), .A1(new_n28259_), .B0(new_n27616_), .B1(new_n27586_), .Y(new_n28262_));
  INVX1    g25826(.A(new_n28262_), .Y(new_n28263_));
  AOI21X1  g25827(.A0(new_n27553_), .A1(new_n27552_), .B0(po1038), .Y(new_n28264_));
  INVX1    g25828(.A(new_n28264_), .Y(new_n28265_));
  OAI22X1  g25829(.A0(new_n28265_), .A1(new_n28263_), .B0(new_n27609_), .B1(new_n27572_), .Y(new_n28266_));
  AOI21X1  g25830(.A0(new_n26582_), .A1(new_n8422_), .B0(po1038), .Y(new_n28267_));
  OAI21X1  g25831(.A0(new_n27904_), .A1(new_n8422_), .B0(new_n28267_), .Y(new_n28268_));
  INVX1    g25832(.A(new_n28268_), .Y(new_n28269_));
  AOI21X1  g25833(.A0(new_n27758_), .A1(new_n27608_), .B0(new_n28269_), .Y(new_n28270_));
  INVX1    g25834(.A(new_n28270_), .Y(new_n28271_));
  MX2X1    g25835(.A(new_n28271_), .B(new_n28266_), .S0(new_n25694_), .Y(new_n28272_));
  AND3X1   g25836(.A(new_n27605_), .B(new_n27578_), .C(po1038), .Y(new_n28273_));
  AND2X1   g25837(.A(new_n27756_), .B(po1038), .Y(new_n28274_));
  INVX1    g25838(.A(new_n28274_), .Y(new_n28275_));
  OAI21X1  g25839(.A0(new_n28275_), .A1(new_n27570_), .B0(new_n28273_), .Y(new_n28276_));
  NOR2X1   g25840(.A(new_n26529_), .B(new_n8422_), .Y(new_n28277_));
  OAI21X1  g25841(.A0(new_n28277_), .A1(new_n27597_), .B0(new_n26534_), .Y(new_n28278_));
  OR3X1    g25842(.A(new_n28278_), .B(new_n26579_), .C(po1038), .Y(new_n28279_));
  NAND3X1  g25843(.A(new_n28279_), .B(new_n28276_), .C(new_n25694_), .Y(new_n28280_));
  AND2X1   g25844(.A(new_n28267_), .B(new_n26570_), .Y(new_n28281_));
  NOR3X1   g25845(.A(new_n26568_), .B(new_n6489_), .C(new_n8422_), .Y(new_n28282_));
  NOR3X1   g25846(.A(new_n28282_), .B(new_n28281_), .C(new_n27579_), .Y(new_n28283_));
  AOI21X1  g25847(.A0(new_n28271_), .A1(new_n26694_), .B0(new_n28283_), .Y(new_n28284_));
  AOI21X1  g25848(.A0(new_n28284_), .A1(pi1151), .B0(pi0268), .Y(new_n28285_));
  AOI22X1  g25849(.A0(new_n28285_), .A1(new_n28280_), .B0(new_n28272_), .B1(pi0268), .Y(new_n28286_));
  OR2X1    g25850(.A(new_n28286_), .B(pi1152), .Y(new_n28287_));
  NOR2X1   g25851(.A(new_n27632_), .B(new_n26602_), .Y(new_n28288_));
  OAI21X1  g25852(.A0(new_n28288_), .A1(new_n28262_), .B0(new_n6489_), .Y(new_n28289_));
  NOR2X1   g25853(.A(new_n27618_), .B(new_n26568_), .Y(new_n28290_));
  OAI22X1  g25854(.A0(new_n28290_), .A1(new_n28289_), .B0(new_n28275_), .B1(new_n27572_), .Y(new_n28291_));
  AOI21X1  g25855(.A0(new_n28274_), .A1(new_n27758_), .B0(new_n28269_), .Y(new_n28292_));
  OAI21X1  g25856(.A0(new_n28265_), .A1(new_n26503_), .B0(new_n28292_), .Y(new_n28293_));
  INVX1    g25857(.A(new_n28293_), .Y(new_n28294_));
  OAI21X1  g25858(.A0(new_n28294_), .A1(new_n25694_), .B0(pi0268), .Y(new_n28295_));
  AOI21X1  g25859(.A0(new_n28291_), .A1(new_n25694_), .B0(new_n28295_), .Y(new_n28296_));
  INVX1    g25860(.A(pi0268), .Y(new_n28297_));
  AOI21X1  g25861(.A0(new_n28278_), .A1(new_n27596_), .B0(po1038), .Y(new_n28298_));
  OAI21X1  g25862(.A0(new_n28298_), .A1(new_n28273_), .B0(new_n25694_), .Y(new_n28299_));
  NOR3X1   g25863(.A(new_n26539_), .B(new_n26530_), .C(pi0219), .Y(new_n28300_));
  OAI21X1  g25864(.A0(new_n28300_), .A1(new_n28261_), .B0(new_n6489_), .Y(new_n28301_));
  AND2X1   g25865(.A(new_n27578_), .B(po1038), .Y(new_n28302_));
  OAI21X1  g25866(.A0(new_n27572_), .A1(pi0219), .B0(new_n28302_), .Y(new_n28303_));
  AND3X1   g25867(.A(new_n28303_), .B(new_n28301_), .C(new_n28276_), .Y(new_n28304_));
  OR2X1    g25868(.A(new_n28304_), .B(new_n25694_), .Y(new_n28305_));
  AND3X1   g25869(.A(new_n28305_), .B(new_n28299_), .C(new_n28297_), .Y(new_n28306_));
  OR3X1    g25870(.A(new_n28306_), .B(new_n28296_), .C(new_n25153_), .Y(new_n28307_));
  AOI21X1  g25871(.A0(new_n28307_), .A1(new_n28287_), .B0(new_n26280_), .Y(new_n28308_));
  NAND3X1  g25872(.A(new_n28000_), .B(new_n27578_), .C(po1038), .Y(new_n28309_));
  NOR2X1   g25873(.A(new_n26561_), .B(pi0219), .Y(new_n28310_));
  OR3X1    g25874(.A(new_n28310_), .B(new_n28301_), .C(new_n26556_), .Y(new_n28311_));
  AND2X1   g25875(.A(new_n28311_), .B(new_n28309_), .Y(new_n28312_));
  INVX1    g25876(.A(new_n28312_), .Y(new_n28313_));
  AOI22X1  g25877(.A0(new_n28302_), .A1(new_n27828_), .B0(new_n28263_), .B1(new_n6489_), .Y(new_n28314_));
  OAI21X1  g25878(.A0(new_n28314_), .A1(new_n25694_), .B0(pi1152), .Y(new_n28315_));
  AOI21X1  g25879(.A0(new_n28313_), .A1(new_n25694_), .B0(new_n28315_), .Y(new_n28316_));
  NOR3X1   g25880(.A(new_n27572_), .B(new_n6489_), .C(pi0219), .Y(new_n28317_));
  INVX1    g25881(.A(new_n28289_), .Y(new_n28318_));
  NOR3X1   g25882(.A(new_n28318_), .B(new_n28282_), .C(new_n28317_), .Y(new_n28319_));
  NOR4X1   g25883(.A(new_n28282_), .B(new_n28281_), .C(new_n27579_), .D(pi1151), .Y(new_n28320_));
  OR2X1    g25884(.A(new_n28320_), .B(pi1152), .Y(new_n28321_));
  AOI21X1  g25885(.A0(new_n28319_), .A1(pi1151), .B0(new_n28321_), .Y(new_n28322_));
  OAI21X1  g25886(.A0(new_n28322_), .A1(new_n28316_), .B0(new_n28297_), .Y(new_n28323_));
  AND2X1   g25887(.A(new_n28140_), .B(pi0219), .Y(new_n28324_));
  INVX1    g25888(.A(new_n28324_), .Y(new_n28325_));
  AOI21X1  g25889(.A0(new_n28325_), .A1(new_n27598_), .B0(new_n27593_), .Y(new_n28326_));
  OAI22X1  g25890(.A0(new_n28326_), .A1(po1038), .B0(new_n28275_), .B1(new_n27606_), .Y(new_n28327_));
  NOR2X1   g25891(.A(new_n27632_), .B(po1038), .Y(new_n28328_));
  AOI22X1  g25892(.A0(new_n28328_), .A1(new_n28325_), .B0(new_n28274_), .B1(new_n27571_), .Y(new_n28329_));
  AOI21X1  g25893(.A0(new_n28329_), .A1(new_n25694_), .B0(new_n25153_), .Y(new_n28330_));
  OAI21X1  g25894(.A0(new_n28327_), .A1(new_n25694_), .B0(new_n28330_), .Y(new_n28331_));
  AND2X1   g25895(.A(new_n27600_), .B(new_n6489_), .Y(new_n28332_));
  AOI21X1  g25896(.A0(new_n28332_), .A1(new_n27598_), .B0(new_n27610_), .Y(new_n28333_));
  NAND2X1  g25897(.A(new_n28333_), .B(pi1151), .Y(new_n28334_));
  OR2X1    g25898(.A(new_n28270_), .B(new_n26694_), .Y(new_n28335_));
  AOI21X1  g25899(.A0(new_n28335_), .A1(new_n25694_), .B0(pi1152), .Y(new_n28336_));
  AOI21X1  g25900(.A0(new_n28336_), .A1(new_n28334_), .B0(new_n28297_), .Y(new_n28337_));
  AOI21X1  g25901(.A0(new_n28337_), .A1(new_n28331_), .B0(pi1150), .Y(new_n28338_));
  AOI21X1  g25902(.A0(new_n28338_), .A1(new_n28323_), .B0(new_n28308_), .Y(new_n28339_));
  NAND2X1  g25903(.A(pi1152), .B(pi0268), .Y(new_n28340_));
  MX2X1    g25904(.A(pi0219), .B(pi0199), .S0(new_n11660_), .Y(new_n28341_));
  AOI22X1  g25905(.A0(new_n24916_), .A1(new_n6489_), .B0(new_n22572_), .B1(new_n23173_), .Y(new_n28342_));
  OAI21X1  g25906(.A0(new_n28342_), .A1(new_n25153_), .B0(new_n28341_), .Y(new_n28343_));
  AOI21X1  g25907(.A0(new_n28342_), .A1(new_n25694_), .B0(new_n26280_), .Y(new_n28344_));
  AND2X1   g25908(.A(new_n28344_), .B(new_n28343_), .Y(new_n28345_));
  AOI22X1  g25909(.A0(new_n27674_), .A1(new_n22572_), .B0(new_n24970_), .B1(new_n6489_), .Y(new_n28346_));
  OR3X1    g25910(.A(new_n28346_), .B(new_n25153_), .C(new_n25694_), .Y(new_n28347_));
  NAND2X1  g25911(.A(new_n27521_), .B(new_n25694_), .Y(new_n28348_));
  MX2X1    g25912(.A(new_n8469_), .B(new_n27664_), .S0(po1038), .Y(new_n28349_));
  OR2X1    g25913(.A(new_n28349_), .B(new_n25694_), .Y(new_n28350_));
  AOI21X1  g25914(.A0(new_n28350_), .A1(new_n25153_), .B0(pi1150), .Y(new_n28351_));
  AND3X1   g25915(.A(new_n28351_), .B(new_n28348_), .C(new_n28347_), .Y(new_n28352_));
  AOI21X1  g25916(.A0(new_n28345_), .A1(new_n28340_), .B0(new_n28352_), .Y(new_n28353_));
  AOI21X1  g25917(.A0(new_n28345_), .A1(pi1152), .B0(new_n2702_), .Y(new_n28354_));
  OAI22X1  g25918(.A0(new_n28354_), .A1(new_n28297_), .B0(new_n28353_), .B1(new_n2702_), .Y(new_n28355_));
  AOI21X1  g25919(.A0(new_n28355_), .A1(new_n28258_), .B0(pi0230), .Y(new_n28356_));
  OAI21X1  g25920(.A0(new_n28339_), .A1(new_n28258_), .B0(new_n28356_), .Y(new_n28357_));
  OR3X1    g25921(.A(new_n28352_), .B(new_n28345_), .C(new_n24814_), .Y(new_n28358_));
  AND2X1   g25922(.A(new_n28358_), .B(new_n28357_), .Y(po0425));
  AOI21X1  g25923(.A0(pi1137), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n28360_));
  NAND2X1  g25924(.A(pi1138), .B(pi0199), .Y(new_n28361_));
  AOI21X1  g25925(.A0(pi1136), .A1(new_n7871_), .B0(pi0200), .Y(new_n28362_));
  AOI21X1  g25926(.A0(new_n28362_), .A1(new_n28361_), .B0(new_n28360_), .Y(new_n28363_));
  OR3X1    g25927(.A(new_n4205_), .B(new_n8422_), .C(pi0211), .Y(new_n28364_));
  MX2X1    g25928(.A(new_n4351_), .B(new_n4554_), .S0(new_n23173_), .Y(new_n28365_));
  OAI21X1  g25929(.A0(new_n28365_), .A1(pi0219), .B0(new_n28364_), .Y(new_n28366_));
  MX2X1    g25930(.A(new_n28366_), .B(new_n28363_), .S0(new_n11660_), .Y(new_n28367_));
  AOI22X1  g25931(.A0(new_n28094_), .A1(new_n7937_), .B0(new_n26670_), .B1(pi1137), .Y(new_n28368_));
  NAND3X1  g25932(.A(new_n28368_), .B(new_n11660_), .C(new_n7871_), .Y(new_n28369_));
  OAI21X1  g25933(.A0(new_n28365_), .A1(new_n2702_), .B0(new_n26027_), .Y(new_n28370_));
  OR2X1    g25934(.A(new_n28029_), .B(pi0817), .Y(new_n28371_));
  AOI21X1  g25935(.A0(new_n28029_), .A1(pi0269), .B0(pi1091), .Y(new_n28372_));
  AOI22X1  g25936(.A0(new_n28372_), .A1(new_n28371_), .B0(new_n28370_), .B1(new_n28369_), .Y(new_n28373_));
  AOI21X1  g25937(.A0(new_n28038_), .A1(pi0269), .B0(pi1091), .Y(new_n28374_));
  OAI21X1  g25938(.A0(new_n28038_), .A1(pi0817), .B0(new_n28374_), .Y(new_n28375_));
  AND3X1   g25939(.A(pi1138), .B(pi1091), .C(new_n23173_), .Y(new_n28376_));
  OR2X1    g25940(.A(new_n11660_), .B(new_n8422_), .Y(new_n28377_));
  AND3X1   g25941(.A(pi1138), .B(pi1091), .C(new_n7937_), .Y(new_n28378_));
  OR2X1    g25942(.A(new_n28378_), .B(new_n7871_), .Y(new_n28379_));
  OAI22X1  g25943(.A0(new_n28379_), .A1(new_n22572_), .B0(new_n28377_), .B1(new_n28376_), .Y(new_n28380_));
  AOI21X1  g25944(.A0(new_n28380_), .A1(new_n28375_), .B0(new_n28373_), .Y(new_n28381_));
  MX2X1    g25945(.A(new_n28381_), .B(new_n28367_), .S0(pi0230), .Y(po0426));
  INVX1    g25946(.A(pi0805), .Y(new_n28383_));
  AND2X1   g25947(.A(new_n26501_), .B(new_n28383_), .Y(new_n28384_));
  OAI21X1  g25948(.A0(new_n26501_), .A1(new_n3817_), .B0(new_n2702_), .Y(new_n28385_));
  AND2X1   g25949(.A(pi1141), .B(new_n23173_), .Y(new_n28386_));
  AOI21X1  g25950(.A0(new_n28386_), .A1(new_n27746_), .B0(new_n28377_), .Y(new_n28387_));
  OR2X1    g25951(.A(new_n28032_), .B(pi0200), .Y(new_n28388_));
  AND3X1   g25952(.A(new_n28388_), .B(new_n11660_), .C(pi0199), .Y(new_n28389_));
  OAI22X1  g25953(.A0(new_n28389_), .A1(new_n28387_), .B0(new_n28385_), .B1(new_n28384_), .Y(new_n28390_));
  AND3X1   g25954(.A(new_n26508_), .B(new_n28383_), .C(pi0314), .Y(new_n28391_));
  OAI21X1  g25955(.A0(new_n28028_), .A1(new_n3817_), .B0(new_n2702_), .Y(new_n28392_));
  MX2X1    g25956(.A(new_n3908_), .B(new_n4019_), .S0(new_n23173_), .Y(new_n28393_));
  OR2X1    g25957(.A(new_n28393_), .B(new_n2702_), .Y(new_n28394_));
  AND2X1   g25958(.A(new_n28394_), .B(new_n26027_), .Y(new_n28395_));
  NAND4X1  g25959(.A(new_n5102_), .B(new_n2933_), .C(new_n7871_), .D(new_n2436_), .Y(new_n28396_));
  AND3X1   g25960(.A(pi1140), .B(pi1091), .C(pi0200), .Y(new_n28397_));
  AND3X1   g25961(.A(pi1139), .B(pi1091), .C(new_n7937_), .Y(new_n28398_));
  NOR3X1   g25962(.A(new_n28398_), .B(new_n28397_), .C(new_n28396_), .Y(new_n28399_));
  OAI22X1  g25963(.A0(new_n28399_), .A1(new_n28395_), .B0(new_n28392_), .B1(new_n28391_), .Y(new_n28400_));
  AND3X1   g25964(.A(new_n28400_), .B(new_n28390_), .C(new_n24814_), .Y(new_n28401_));
  INVX1    g25965(.A(new_n28386_), .Y(new_n28402_));
  MX2X1    g25966(.A(new_n28393_), .B(new_n28402_), .S0(pi0219), .Y(new_n28403_));
  OR2X1    g25967(.A(new_n3908_), .B(pi0199), .Y(new_n28404_));
  NAND2X1  g25968(.A(pi1141), .B(pi0199), .Y(new_n28405_));
  AOI21X1  g25969(.A0(pi1139), .A1(new_n7871_), .B0(pi0200), .Y(new_n28406_));
  AOI22X1  g25970(.A0(new_n28406_), .A1(new_n28405_), .B0(new_n28404_), .B1(pi0200), .Y(new_n28407_));
  OAI21X1  g25971(.A0(new_n28407_), .A1(new_n22572_), .B0(pi0230), .Y(new_n28408_));
  AOI21X1  g25972(.A0(new_n28403_), .A1(new_n22572_), .B0(new_n28408_), .Y(new_n28409_));
  OR2X1    g25973(.A(new_n28409_), .B(new_n28401_), .Y(po0427));
  MX2X1    g25974(.A(new_n26695_), .B(new_n26503_), .S0(pi0271), .Y(new_n28411_));
  INVX1    g25975(.A(new_n28411_), .Y(new_n28412_));
  AND2X1   g25976(.A(new_n26509_), .B(new_n2702_), .Y(new_n28413_));
  MX2X1    g25977(.A(new_n28413_), .B(new_n26510_), .S0(new_n26500_), .Y(new_n28414_));
  AND2X1   g25978(.A(pi1146), .B(pi1091), .Y(new_n28415_));
  NOR2X1   g25979(.A(new_n28415_), .B(new_n28414_), .Y(new_n28416_));
  AND2X1   g25980(.A(new_n28415_), .B(new_n23173_), .Y(new_n28417_));
  OR2X1    g25981(.A(new_n28417_), .B(new_n28416_), .Y(new_n28418_));
  AOI21X1  g25982(.A0(new_n26067_), .A1(pi1091), .B0(pi0219), .Y(new_n28419_));
  AOI22X1  g25983(.A0(new_n28419_), .A1(new_n28418_), .B0(new_n28412_), .B1(pi0219), .Y(new_n28420_));
  OR2X1    g25984(.A(new_n25993_), .B(pi0211), .Y(new_n28421_));
  OAI21X1  g25985(.A0(new_n28421_), .A1(new_n27574_), .B0(new_n22572_), .Y(new_n28422_));
  MX2X1    g25986(.A(new_n28416_), .B(new_n28412_), .S0(pi0199), .Y(new_n28423_));
  AND2X1   g25987(.A(pi1145), .B(pi1091), .Y(new_n28424_));
  OR2X1    g25988(.A(new_n28424_), .B(pi0199), .Y(new_n28425_));
  OAI22X1  g25989(.A0(new_n28425_), .A1(new_n28414_), .B0(new_n28411_), .B1(new_n7871_), .Y(new_n28426_));
  AOI21X1  g25990(.A0(new_n26660_), .A1(pi1147), .B0(pi0200), .Y(new_n28427_));
  AOI22X1  g25991(.A0(new_n28427_), .A1(new_n28426_), .B0(new_n28423_), .B1(pi0200), .Y(new_n28428_));
  OAI22X1  g25992(.A0(new_n28428_), .A1(new_n22572_), .B0(new_n28422_), .B1(new_n28420_), .Y(new_n28429_));
  MX2X1    g25993(.A(new_n26106_), .B(new_n25605_), .S0(new_n23173_), .Y(new_n28430_));
  AND2X1   g25994(.A(new_n28430_), .B(new_n8422_), .Y(new_n28431_));
  AOI21X1  g25995(.A0(pi1145), .A1(new_n7871_), .B0(pi0200), .Y(new_n28432_));
  OR3X1    g25996(.A(new_n28432_), .B(new_n26152_), .C(pi0299), .Y(new_n28433_));
  OAI21X1  g25997(.A0(new_n27519_), .A1(new_n25993_), .B0(new_n28433_), .Y(new_n28434_));
  OAI21X1  g25998(.A0(new_n28434_), .A1(new_n28431_), .B0(new_n6489_), .Y(new_n28435_));
  NOR2X1   g25999(.A(new_n26962_), .B(new_n26067_), .Y(new_n28436_));
  AOI21X1  g26000(.A0(new_n28421_), .A1(pi0219), .B0(new_n28436_), .Y(new_n28437_));
  AOI21X1  g26001(.A0(new_n28437_), .A1(po1038), .B0(new_n24814_), .Y(new_n28438_));
  AOI22X1  g26002(.A0(new_n28438_), .A1(new_n28435_), .B0(new_n28429_), .B1(new_n24814_), .Y(po0428));
  OAI21X1  g26003(.A0(new_n28271_), .A1(pi1150), .B0(pi1149), .Y(new_n28440_));
  AOI21X1  g26004(.A0(new_n28294_), .A1(pi1150), .B0(new_n28440_), .Y(new_n28441_));
  INVX1    g26005(.A(new_n28291_), .Y(new_n28442_));
  OAI21X1  g26006(.A0(new_n28266_), .A1(pi1150), .B0(new_n25955_), .Y(new_n28443_));
  AOI21X1  g26007(.A0(new_n28442_), .A1(pi1150), .B0(new_n28443_), .Y(new_n28444_));
  OAI21X1  g26008(.A0(new_n28444_), .A1(new_n28441_), .B0(pi1148), .Y(new_n28445_));
  INVX1    g26009(.A(pi0283), .Y(new_n28446_));
  INVX1    g26010(.A(new_n28329_), .Y(new_n28447_));
  AOI21X1  g26011(.A0(new_n28335_), .A1(new_n26280_), .B0(pi1149), .Y(new_n28448_));
  OAI21X1  g26012(.A0(new_n28447_), .A1(new_n26280_), .B0(new_n28448_), .Y(new_n28449_));
  NOR2X1   g26013(.A(new_n28327_), .B(new_n26280_), .Y(new_n28450_));
  AND2X1   g26014(.A(new_n28333_), .B(new_n26280_), .Y(new_n28451_));
  OR2X1    g26015(.A(new_n28451_), .B(new_n25955_), .Y(new_n28452_));
  OAI21X1  g26016(.A0(new_n28452_), .A1(new_n28450_), .B0(new_n28449_), .Y(new_n28453_));
  AOI21X1  g26017(.A0(new_n28453_), .A1(new_n26084_), .B0(new_n28446_), .Y(new_n28454_));
  INVX1    g26018(.A(pi0272), .Y(new_n28455_));
  INVX1    g26019(.A(new_n28341_), .Y(new_n28456_));
  MX2X1    g26020(.A(new_n9449_), .B(new_n27524_), .S0(po1038), .Y(new_n28457_));
  AOI21X1  g26021(.A0(new_n28457_), .A1(new_n26280_), .B0(new_n28342_), .Y(new_n28458_));
  AOI21X1  g26022(.A0(new_n26280_), .A1(pi1149), .B0(new_n28342_), .Y(new_n28459_));
  OAI22X1  g26023(.A0(new_n28459_), .A1(new_n28456_), .B0(new_n28458_), .B1(pi1149), .Y(new_n28460_));
  AOI21X1  g26024(.A0(new_n28460_), .A1(pi1091), .B0(new_n26084_), .Y(new_n28461_));
  AOI21X1  g26025(.A0(new_n27522_), .A1(pi1150), .B0(pi1149), .Y(new_n28462_));
  INVX1    g26026(.A(new_n28346_), .Y(new_n28463_));
  AOI21X1  g26027(.A0(new_n28463_), .A1(pi1091), .B0(new_n26280_), .Y(new_n28464_));
  OAI22X1  g26028(.A0(new_n27807_), .A1(new_n11660_), .B0(new_n26665_), .B1(po1038), .Y(new_n28465_));
  OAI21X1  g26029(.A0(new_n28465_), .A1(pi1150), .B0(pi1149), .Y(new_n28466_));
  OAI21X1  g26030(.A0(new_n28466_), .A1(new_n28464_), .B0(new_n26084_), .Y(new_n28467_));
  AOI21X1  g26031(.A0(new_n28462_), .A1(pi1091), .B0(new_n28467_), .Y(new_n28468_));
  NOR3X1   g26032(.A(new_n28468_), .B(new_n28461_), .C(pi0283), .Y(new_n28469_));
  OR2X1    g26033(.A(new_n28469_), .B(new_n28455_), .Y(new_n28470_));
  AOI21X1  g26034(.A0(new_n28454_), .A1(new_n28445_), .B0(new_n28470_), .Y(new_n28471_));
  OR2X1    g26035(.A(new_n28304_), .B(new_n26280_), .Y(new_n28472_));
  OR2X1    g26036(.A(new_n28284_), .B(pi1150), .Y(new_n28473_));
  AND3X1   g26037(.A(new_n28473_), .B(new_n28472_), .C(pi1149), .Y(new_n28474_));
  OAI21X1  g26038(.A0(new_n28298_), .A1(new_n28273_), .B0(pi1150), .Y(new_n28475_));
  AOI21X1  g26039(.A0(new_n28279_), .A1(new_n28276_), .B0(pi1150), .Y(new_n28476_));
  NOR2X1   g26040(.A(new_n28476_), .B(pi1149), .Y(new_n28477_));
  AOI21X1  g26041(.A0(new_n28477_), .A1(new_n28475_), .B0(new_n28474_), .Y(new_n28478_));
  INVX1    g26042(.A(new_n28319_), .Y(new_n28479_));
  NAND2X1  g26043(.A(new_n28314_), .B(pi1150), .Y(new_n28480_));
  NAND2X1  g26044(.A(new_n28480_), .B(pi1149), .Y(new_n28481_));
  AOI21X1  g26045(.A0(new_n28479_), .A1(new_n26280_), .B0(new_n28481_), .Y(new_n28482_));
  AND3X1   g26046(.A(new_n28311_), .B(new_n28309_), .C(pi1150), .Y(new_n28483_));
  OAI21X1  g26047(.A0(new_n28283_), .A1(pi1150), .B0(new_n25955_), .Y(new_n28484_));
  OAI21X1  g26048(.A0(new_n28484_), .A1(new_n28483_), .B0(new_n26084_), .Y(new_n28485_));
  OAI22X1  g26049(.A0(new_n28485_), .A1(new_n28482_), .B0(new_n28478_), .B1(new_n26084_), .Y(new_n28486_));
  OR2X1    g26050(.A(new_n11660_), .B(pi0211), .Y(new_n28487_));
  AOI21X1  g26051(.A0(new_n24907_), .A1(new_n6489_), .B0(new_n26027_), .Y(new_n28488_));
  AOI21X1  g26052(.A0(new_n28488_), .A1(new_n28487_), .B0(new_n26280_), .Y(new_n28489_));
  NOR3X1   g26053(.A(new_n28489_), .B(new_n28456_), .C(new_n25955_), .Y(new_n28490_));
  OAI21X1  g26054(.A0(new_n28458_), .A1(pi1149), .B0(pi1148), .Y(new_n28491_));
  NOR3X1   g26055(.A(new_n28491_), .B(new_n28490_), .C(new_n2702_), .Y(new_n28492_));
  OR2X1    g26056(.A(new_n28462_), .B(pi1148), .Y(new_n28493_));
  AND2X1   g26057(.A(new_n28346_), .B(pi1150), .Y(new_n28494_));
  OAI21X1  g26058(.A0(new_n28349_), .A1(pi1150), .B0(pi1149), .Y(new_n28495_));
  OAI21X1  g26059(.A0(new_n28495_), .A1(new_n28494_), .B0(pi1091), .Y(new_n28496_));
  OAI21X1  g26060(.A0(new_n28496_), .A1(new_n28493_), .B0(new_n28446_), .Y(new_n28497_));
  OAI21X1  g26061(.A0(new_n28497_), .A1(new_n28492_), .B0(new_n28455_), .Y(new_n28498_));
  AOI21X1  g26062(.A0(new_n28486_), .A1(pi0283), .B0(new_n28498_), .Y(new_n28499_));
  OR3X1    g26063(.A(new_n28499_), .B(new_n28471_), .C(pi0230), .Y(new_n28500_));
  OR2X1    g26064(.A(new_n28349_), .B(pi1150), .Y(new_n28501_));
  AOI21X1  g26065(.A0(new_n28489_), .A1(new_n28346_), .B0(new_n25955_), .Y(new_n28502_));
  AOI21X1  g26066(.A0(new_n28502_), .A1(new_n28501_), .B0(new_n28493_), .Y(new_n28503_));
  OAI21X1  g26067(.A0(new_n28491_), .A1(new_n28490_), .B0(pi0230), .Y(new_n28504_));
  OR2X1    g26068(.A(new_n28504_), .B(new_n28503_), .Y(new_n28505_));
  AND2X1   g26069(.A(new_n28505_), .B(new_n28500_), .Y(po0429));
  OAI21X1  g26070(.A0(new_n26528_), .A1(pi0273), .B0(new_n26512_), .Y(new_n28507_));
  NAND2X1  g26071(.A(new_n28507_), .B(pi0219), .Y(new_n28508_));
  OR3X1    g26072(.A(new_n26509_), .B(pi1091), .C(new_n26500_), .Y(new_n28509_));
  AOI21X1  g26073(.A0(new_n28509_), .A1(new_n26513_), .B0(new_n28230_), .Y(new_n28510_));
  OR2X1    g26074(.A(new_n28417_), .B(pi0219), .Y(new_n28511_));
  OAI21X1  g26075(.A0(new_n28511_), .A1(new_n28510_), .B0(new_n28508_), .Y(new_n28512_));
  AND2X1   g26076(.A(new_n28415_), .B(new_n7937_), .Y(new_n28513_));
  OR2X1    g26077(.A(new_n28513_), .B(pi0199), .Y(new_n28514_));
  AOI21X1  g26078(.A0(new_n28507_), .A1(pi0199), .B0(pi0299), .Y(new_n28515_));
  OAI21X1  g26079(.A0(new_n28514_), .A1(new_n28510_), .B0(new_n28515_), .Y(new_n28516_));
  OAI21X1  g26080(.A0(new_n28512_), .A1(new_n2933_), .B0(new_n28516_), .Y(new_n28517_));
  OR2X1    g26081(.A(new_n26631_), .B(new_n8468_), .Y(new_n28518_));
  AOI21X1  g26082(.A0(new_n28518_), .A1(pi1091), .B0(new_n28517_), .Y(new_n28519_));
  OR3X1    g26083(.A(new_n27609_), .B(new_n27606_), .C(new_n2702_), .Y(new_n28520_));
  OAI21X1  g26084(.A0(new_n28519_), .A1(po1038), .B0(new_n28520_), .Y(new_n28521_));
  AOI21X1  g26085(.A0(new_n28517_), .A1(new_n26204_), .B0(pi1148), .Y(new_n28522_));
  OR3X1    g26086(.A(new_n2702_), .B(new_n8422_), .C(pi0211), .Y(new_n28523_));
  AOI21X1  g26087(.A0(new_n28523_), .A1(new_n28512_), .B0(new_n2933_), .Y(new_n28524_));
  INVX1    g26088(.A(new_n26661_), .Y(new_n28525_));
  AND2X1   g26089(.A(new_n28423_), .B(pi0200), .Y(new_n28526_));
  OAI21X1  g26090(.A0(new_n28526_), .A1(new_n28525_), .B0(new_n28516_), .Y(new_n28527_));
  OAI21X1  g26091(.A0(new_n28527_), .A1(new_n28524_), .B0(new_n6489_), .Y(new_n28528_));
  OR3X1    g26092(.A(new_n27574_), .B(new_n6489_), .C(pi0211), .Y(new_n28529_));
  AND3X1   g26093(.A(new_n28529_), .B(new_n28528_), .C(pi1148), .Y(new_n28530_));
  OAI22X1  g26094(.A0(new_n28530_), .A1(new_n28522_), .B0(new_n28512_), .B1(new_n6489_), .Y(new_n28531_));
  AOI21X1  g26095(.A0(new_n28521_), .A1(pi1147), .B0(new_n28531_), .Y(new_n28532_));
  OAI21X1  g26096(.A0(new_n26106_), .A1(pi0211), .B0(new_n26027_), .Y(new_n28533_));
  NOR3X1   g26097(.A(pi1146), .B(pi0200), .C(pi0199), .Y(new_n28534_));
  OAI21X1  g26098(.A0(new_n28534_), .A1(new_n28396_), .B0(new_n28533_), .Y(new_n28535_));
  NAND2X1  g26099(.A(new_n26903_), .B(pi1146), .Y(new_n28536_));
  OAI21X1  g26100(.A0(new_n28536_), .A1(new_n28457_), .B0(new_n26084_), .Y(new_n28537_));
  AOI21X1  g26101(.A0(new_n28535_), .A1(pi1147), .B0(new_n28537_), .Y(new_n28538_));
  OR3X1    g26102(.A(new_n11660_), .B(new_n25993_), .C(pi0219), .Y(new_n28539_));
  AOI22X1  g26103(.A0(new_n28539_), .A1(new_n28487_), .B0(new_n7997_), .B1(new_n3140_), .Y(new_n28540_));
  AOI21X1  g26104(.A0(pi1147), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n28541_));
  OR2X1    g26105(.A(new_n28541_), .B(new_n28534_), .Y(new_n28542_));
  OAI21X1  g26106(.A0(new_n28542_), .A1(new_n22572_), .B0(pi1148), .Y(new_n28543_));
  OAI21X1  g26107(.A0(new_n28543_), .A1(new_n28540_), .B0(pi0230), .Y(new_n28544_));
  OAI22X1  g26108(.A0(new_n28544_), .A1(new_n28538_), .B0(new_n28532_), .B1(pi0230), .Y(po0430));
  AOI21X1  g26109(.A0(new_n28029_), .A1(pi0274), .B0(pi1091), .Y(new_n28546_));
  OAI21X1  g26110(.A0(new_n28029_), .A1(pi0659), .B0(new_n28546_), .Y(new_n28547_));
  OAI21X1  g26111(.A0(new_n2439_), .A1(new_n2702_), .B0(new_n28547_), .Y(new_n28548_));
  AND2X1   g26112(.A(new_n28548_), .B(pi0200), .Y(new_n28549_));
  AOI21X1  g26113(.A0(new_n28547_), .A1(new_n28060_), .B0(pi0200), .Y(new_n28550_));
  OR2X1    g26114(.A(new_n28550_), .B(pi0199), .Y(new_n28551_));
  AOI21X1  g26115(.A0(new_n28038_), .A1(pi0274), .B0(pi1091), .Y(new_n28552_));
  OAI21X1  g26116(.A0(new_n28038_), .A1(pi0659), .B0(new_n28552_), .Y(new_n28553_));
  AOI21X1  g26117(.A0(new_n28424_), .A1(new_n7937_), .B0(new_n7871_), .Y(new_n28554_));
  AOI21X1  g26118(.A0(new_n28554_), .A1(new_n28553_), .B0(new_n22572_), .Y(new_n28555_));
  OAI21X1  g26119(.A0(new_n28551_), .A1(new_n28549_), .B0(new_n28555_), .Y(new_n28556_));
  AND2X1   g26120(.A(new_n28548_), .B(pi0211), .Y(new_n28557_));
  AOI21X1  g26121(.A0(new_n28547_), .A1(new_n28060_), .B0(pi0211), .Y(new_n28558_));
  OR3X1    g26122(.A(new_n28558_), .B(new_n28557_), .C(pi0219), .Y(new_n28559_));
  AOI21X1  g26123(.A0(new_n26067_), .A1(pi1091), .B0(new_n8422_), .Y(new_n28560_));
  AOI21X1  g26124(.A0(new_n28560_), .A1(new_n28553_), .B0(new_n11660_), .Y(new_n28561_));
  AOI21X1  g26125(.A0(new_n28561_), .A1(new_n28559_), .B0(pi0230), .Y(new_n28562_));
  AND2X1   g26126(.A(pi1144), .B(pi0211), .Y(new_n28563_));
  NOR3X1   g26127(.A(new_n28563_), .B(new_n24826_), .C(pi0219), .Y(new_n28564_));
  OR2X1    g26128(.A(new_n28564_), .B(new_n26068_), .Y(new_n28565_));
  NAND2X1  g26129(.A(new_n25498_), .B(new_n2933_), .Y(new_n28566_));
  AOI22X1  g26130(.A0(new_n25605_), .A1(new_n23173_), .B0(pi0299), .B1(new_n8422_), .Y(new_n28567_));
  AND2X1   g26131(.A(new_n26157_), .B(new_n24837_), .Y(new_n28568_));
  OAI22X1  g26132(.A0(new_n28568_), .A1(new_n28566_), .B0(new_n28567_), .B1(new_n28564_), .Y(new_n28569_));
  AOI21X1  g26133(.A0(new_n28569_), .A1(new_n6489_), .B0(new_n24814_), .Y(new_n28570_));
  AOI22X1  g26134(.A0(new_n28570_), .A1(new_n28565_), .B0(new_n28562_), .B1(new_n28556_), .Y(po0431));
  AND2X1   g26135(.A(new_n28341_), .B(pi1149), .Y(new_n28572_));
  OAI21X1  g26136(.A0(new_n28342_), .A1(new_n25694_), .B0(new_n28572_), .Y(new_n28573_));
  AOI21X1  g26137(.A0(new_n28349_), .A1(new_n25694_), .B0(new_n26280_), .Y(new_n28574_));
  OAI21X1  g26138(.A0(new_n28346_), .A1(new_n25694_), .B0(new_n28574_), .Y(new_n28575_));
  OR3X1    g26139(.A(new_n27521_), .B(new_n25694_), .C(pi1150), .Y(new_n28576_));
  NAND3X1  g26140(.A(new_n28576_), .B(new_n28575_), .C(new_n25955_), .Y(new_n28577_));
  NAND3X1  g26141(.A(new_n28342_), .B(new_n26280_), .C(pi1149), .Y(new_n28578_));
  AND3X1   g26142(.A(new_n28578_), .B(new_n28577_), .C(new_n28573_), .Y(new_n28579_));
  AND2X1   g26143(.A(pi0283), .B(pi0272), .Y(new_n28580_));
  INVX1    g26144(.A(pi0275), .Y(new_n28581_));
  OR3X1    g26145(.A(new_n28346_), .B(new_n25694_), .C(pi1149), .Y(new_n28582_));
  AND2X1   g26146(.A(new_n28582_), .B(new_n28573_), .Y(new_n28583_));
  OR2X1    g26147(.A(new_n28342_), .B(new_n25955_), .Y(new_n28584_));
  AOI21X1  g26148(.A0(new_n28457_), .A1(new_n25694_), .B0(new_n28584_), .Y(new_n28585_));
  OR2X1    g26149(.A(new_n25694_), .B(pi1149), .Y(new_n28586_));
  OAI21X1  g26150(.A0(new_n28586_), .A1(new_n27521_), .B0(new_n26280_), .Y(new_n28587_));
  OAI22X1  g26151(.A0(new_n28587_), .A1(new_n28585_), .B0(new_n28583_), .B1(new_n26280_), .Y(new_n28588_));
  AND3X1   g26152(.A(new_n25694_), .B(pi1150), .C(new_n25955_), .Y(new_n28589_));
  AOI22X1  g26153(.A0(new_n28589_), .A1(new_n28465_), .B0(new_n28588_), .B1(pi1091), .Y(new_n28590_));
  NOR2X1   g26154(.A(new_n28590_), .B(new_n28581_), .Y(new_n28591_));
  AOI21X1  g26155(.A0(new_n28579_), .A1(pi1091), .B0(pi0275), .Y(new_n28592_));
  OR3X1    g26156(.A(new_n28592_), .B(new_n28591_), .C(new_n28580_), .Y(new_n28593_));
  NAND3X1  g26157(.A(new_n28311_), .B(new_n28309_), .C(new_n26280_), .Y(new_n28594_));
  AND3X1   g26158(.A(new_n28594_), .B(new_n28480_), .C(pi1151), .Y(new_n28595_));
  OAI21X1  g26159(.A0(new_n28283_), .A1(pi1150), .B0(new_n25694_), .Y(new_n28596_));
  AOI21X1  g26160(.A0(new_n28479_), .A1(pi1150), .B0(new_n28596_), .Y(new_n28597_));
  OAI21X1  g26161(.A0(new_n28597_), .A1(new_n28595_), .B0(new_n28581_), .Y(new_n28598_));
  MX2X1    g26162(.A(new_n28447_), .B(new_n28327_), .S0(pi1150), .Y(new_n28599_));
  MX2X1    g26163(.A(new_n28335_), .B(new_n28333_), .S0(pi1150), .Y(new_n28600_));
  AOI21X1  g26164(.A0(new_n28600_), .A1(new_n25694_), .B0(new_n28581_), .Y(new_n28601_));
  OAI21X1  g26165(.A0(new_n28599_), .A1(new_n25694_), .B0(new_n28601_), .Y(new_n28602_));
  AND3X1   g26166(.A(new_n28602_), .B(new_n28598_), .C(new_n25955_), .Y(new_n28603_));
  AOI21X1  g26167(.A0(new_n28266_), .A1(new_n25694_), .B0(pi1150), .Y(new_n28604_));
  OAI21X1  g26168(.A0(new_n28442_), .A1(new_n25694_), .B0(new_n28604_), .Y(new_n28605_));
  AOI21X1  g26169(.A0(new_n28271_), .A1(new_n25694_), .B0(new_n26280_), .Y(new_n28606_));
  OAI21X1  g26170(.A0(new_n28294_), .A1(new_n25694_), .B0(new_n28606_), .Y(new_n28607_));
  AND3X1   g26171(.A(new_n28607_), .B(new_n28605_), .C(pi0275), .Y(new_n28608_));
  OAI21X1  g26172(.A0(new_n28298_), .A1(new_n28273_), .B0(new_n26280_), .Y(new_n28609_));
  AND3X1   g26173(.A(new_n28609_), .B(new_n28472_), .C(pi1151), .Y(new_n28610_));
  OAI21X1  g26174(.A0(new_n28284_), .A1(new_n26280_), .B0(new_n25694_), .Y(new_n28611_));
  OAI21X1  g26175(.A0(new_n28611_), .A1(new_n28476_), .B0(new_n28581_), .Y(new_n28612_));
  OAI21X1  g26176(.A0(new_n28612_), .A1(new_n28610_), .B0(pi1149), .Y(new_n28613_));
  OAI21X1  g26177(.A0(new_n28613_), .A1(new_n28608_), .B0(new_n28580_), .Y(new_n28614_));
  OAI21X1  g26178(.A0(new_n28614_), .A1(new_n28603_), .B0(new_n28593_), .Y(new_n28615_));
  MX2X1    g26179(.A(new_n28615_), .B(new_n28579_), .S0(pi0230), .Y(po0432));
  INVX1    g26180(.A(pi0802), .Y(new_n28617_));
  OAI21X1  g26181(.A0(new_n28029_), .A1(new_n28617_), .B0(new_n3151_), .Y(new_n28618_));
  MX2X1    g26182(.A(new_n3309_), .B(new_n2439_), .S0(new_n23173_), .Y(new_n28619_));
  OAI21X1  g26183(.A0(new_n28619_), .A1(new_n2702_), .B0(new_n26027_), .Y(new_n28620_));
  AND2X1   g26184(.A(new_n28065_), .B(new_n7937_), .Y(new_n28621_));
  AND3X1   g26185(.A(pi1145), .B(pi1091), .C(pi0200), .Y(new_n28622_));
  OR3X1    g26186(.A(new_n28622_), .B(new_n28396_), .C(new_n28621_), .Y(new_n28623_));
  AOI22X1  g26187(.A0(new_n28623_), .A1(new_n28620_), .B0(new_n28618_), .B1(new_n28413_), .Y(new_n28624_));
  OAI21X1  g26188(.A0(new_n28038_), .A1(new_n28617_), .B0(new_n3151_), .Y(new_n28625_));
  OR3X1    g26189(.A(new_n28417_), .B(new_n11660_), .C(new_n8422_), .Y(new_n28626_));
  OR3X1    g26190(.A(new_n28513_), .B(new_n22572_), .C(new_n7871_), .Y(new_n28627_));
  AOI22X1  g26191(.A0(new_n28627_), .A1(new_n28626_), .B0(new_n28625_), .B1(new_n26503_), .Y(new_n28628_));
  OR3X1    g26192(.A(new_n28628_), .B(new_n28624_), .C(pi0230), .Y(new_n28629_));
  OAI21X1  g26193(.A0(new_n2439_), .A1(pi0199), .B0(new_n26793_), .Y(new_n28630_));
  AOI21X1  g26194(.A0(new_n28630_), .A1(new_n26159_), .B0(new_n22572_), .Y(new_n28631_));
  OAI22X1  g26195(.A0(new_n28619_), .A1(pi0219), .B0(new_n24894_), .B1(new_n3140_), .Y(new_n28632_));
  OAI21X1  g26196(.A0(new_n28632_), .A1(new_n11660_), .B0(pi0230), .Y(new_n28633_));
  OAI21X1  g26197(.A0(new_n28633_), .A1(new_n28631_), .B0(new_n28629_), .Y(po0433));
  NAND2X1  g26198(.A(pi1140), .B(pi1091), .Y(new_n28635_));
  AOI21X1  g26199(.A0(new_n28029_), .A1(pi0277), .B0(pi1091), .Y(new_n28636_));
  OAI21X1  g26200(.A0(new_n28029_), .A1(pi0820), .B0(new_n28636_), .Y(new_n28637_));
  AOI21X1  g26201(.A0(new_n28637_), .A1(new_n28635_), .B0(pi0200), .Y(new_n28638_));
  AOI21X1  g26202(.A0(new_n28637_), .A1(new_n28032_), .B0(new_n7937_), .Y(new_n28639_));
  OR3X1    g26203(.A(new_n28639_), .B(new_n28638_), .C(pi0199), .Y(new_n28640_));
  AOI21X1  g26204(.A0(new_n28038_), .A1(pi0277), .B0(pi1091), .Y(new_n28641_));
  OAI21X1  g26205(.A0(new_n28038_), .A1(pi0820), .B0(new_n28641_), .Y(new_n28642_));
  AOI21X1  g26206(.A0(new_n28034_), .A1(new_n7937_), .B0(new_n7871_), .Y(new_n28643_));
  AOI21X1  g26207(.A0(new_n28643_), .A1(new_n28642_), .B0(new_n22572_), .Y(new_n28644_));
  AOI21X1  g26208(.A0(new_n28637_), .A1(new_n28635_), .B0(pi0211), .Y(new_n28645_));
  AOI21X1  g26209(.A0(new_n28637_), .A1(new_n28032_), .B0(new_n23173_), .Y(new_n28646_));
  OR3X1    g26210(.A(new_n28646_), .B(new_n28645_), .C(pi0219), .Y(new_n28647_));
  OAI21X1  g26211(.A0(new_n24820_), .A1(pi0211), .B0(pi0219), .Y(new_n28648_));
  OAI21X1  g26212(.A0(new_n27746_), .A1(new_n8422_), .B0(new_n28648_), .Y(new_n28649_));
  AOI21X1  g26213(.A0(new_n28649_), .A1(new_n28642_), .B0(new_n11660_), .Y(new_n28650_));
  AOI22X1  g26214(.A0(new_n28650_), .A1(new_n28647_), .B0(new_n28644_), .B1(new_n28640_), .Y(new_n28651_));
  AOI21X1  g26215(.A0(pi1140), .A1(new_n23173_), .B0(pi0219), .Y(new_n28652_));
  OAI21X1  g26216(.A0(new_n3759_), .A1(new_n23173_), .B0(new_n28652_), .Y(new_n28653_));
  AOI21X1  g26217(.A0(new_n28653_), .A1(new_n28648_), .B0(new_n11660_), .Y(new_n28654_));
  AOI22X1  g26218(.A0(new_n28404_), .A1(new_n24832_), .B0(new_n28053_), .B1(pi0200), .Y(new_n28655_));
  OAI21X1  g26219(.A0(new_n28655_), .A1(new_n22572_), .B0(pi0230), .Y(new_n28656_));
  OAI22X1  g26220(.A0(new_n28656_), .A1(new_n28654_), .B0(new_n28651_), .B1(pi0230), .Y(po0434));
  INVX1    g26221(.A(pi0278), .Y(po1130));
  OAI21X1  g26222(.A0(new_n28038_), .A1(pi0976), .B0(new_n2702_), .Y(new_n28659_));
  AOI21X1  g26223(.A0(new_n28038_), .A1(po1130), .B0(new_n28659_), .Y(new_n28660_));
  INVX1    g26224(.A(pi1132), .Y(new_n28661_));
  NAND3X1  g26225(.A(new_n26508_), .B(pi0976), .C(pi0314), .Y(new_n28662_));
  AOI21X1  g26226(.A0(new_n28029_), .A1(pi0278), .B0(pi1091), .Y(new_n28663_));
  AOI22X1  g26227(.A0(new_n28663_), .A1(new_n28662_), .B0(new_n28661_), .B1(pi1091), .Y(new_n28664_));
  MX2X1    g26228(.A(new_n28664_), .B(new_n28660_), .S0(pi0199), .Y(new_n28665_));
  OR2X1    g26229(.A(new_n28665_), .B(pi0200), .Y(new_n28666_));
  INVX1    g26230(.A(pi1133), .Y(new_n28667_));
  AOI22X1  g26231(.A0(new_n28663_), .A1(new_n28662_), .B0(new_n28667_), .B1(pi1091), .Y(new_n28668_));
  MX2X1    g26232(.A(new_n28668_), .B(new_n28660_), .S0(pi0199), .Y(new_n28669_));
  OR2X1    g26233(.A(new_n28669_), .B(new_n7937_), .Y(new_n28670_));
  AND2X1   g26234(.A(new_n28670_), .B(new_n2933_), .Y(new_n28671_));
  MX2X1    g26235(.A(pi1132), .B(pi1133), .S0(pi0211), .Y(new_n28672_));
  INVX1    g26236(.A(new_n28672_), .Y(new_n28673_));
  AOI22X1  g26237(.A0(new_n28673_), .A1(pi1091), .B0(new_n28663_), .B1(new_n28662_), .Y(new_n28674_));
  MX2X1    g26238(.A(new_n28674_), .B(new_n28660_), .S0(pi0219), .Y(new_n28675_));
  AOI22X1  g26239(.A0(new_n28675_), .A1(pi0299), .B0(new_n28671_), .B1(new_n28666_), .Y(new_n28676_));
  AOI21X1  g26240(.A0(new_n28675_), .A1(po1038), .B0(pi0230), .Y(new_n28677_));
  OAI21X1  g26241(.A0(new_n28676_), .A1(po1038), .B0(new_n28677_), .Y(new_n28678_));
  AND2X1   g26242(.A(new_n28672_), .B(new_n25796_), .Y(new_n28679_));
  OAI21X1  g26243(.A0(new_n28661_), .A1(pi0199), .B0(new_n7937_), .Y(new_n28680_));
  OAI21X1  g26244(.A0(new_n28667_), .A1(pi0199), .B0(pi0200), .Y(new_n28681_));
  NAND3X1  g26245(.A(new_n28681_), .B(new_n28680_), .C(new_n2933_), .Y(new_n28682_));
  NAND3X1  g26246(.A(new_n28672_), .B(pi0299), .C(new_n8422_), .Y(new_n28683_));
  AOI21X1  g26247(.A0(new_n28683_), .A1(new_n28682_), .B0(po1038), .Y(new_n28684_));
  OR3X1    g26248(.A(new_n28684_), .B(new_n28679_), .C(new_n24814_), .Y(new_n28685_));
  AOI21X1  g26249(.A0(new_n28685_), .A1(new_n28678_), .B0(pi1134), .Y(new_n28686_));
  AOI21X1  g26250(.A0(new_n28673_), .A1(new_n8422_), .B0(new_n25957_), .Y(new_n28687_));
  OR3X1    g26251(.A(pi1132), .B(pi0200), .C(pi0199), .Y(new_n28688_));
  NAND3X1  g26252(.A(new_n28688_), .B(new_n28681_), .C(new_n2933_), .Y(new_n28689_));
  AOI22X1  g26253(.A0(new_n28672_), .A1(new_n24884_), .B0(new_n24893_), .B1(pi0299), .Y(new_n28690_));
  AOI21X1  g26254(.A0(new_n28690_), .A1(new_n28689_), .B0(po1038), .Y(new_n28691_));
  OR3X1    g26255(.A(new_n28691_), .B(new_n28687_), .C(new_n24814_), .Y(new_n28692_));
  OAI21X1  g26256(.A0(new_n28666_), .A1(new_n26660_), .B0(new_n28671_), .Y(new_n28693_));
  AOI22X1  g26257(.A0(new_n28675_), .A1(pi0299), .B0(new_n27746_), .B1(new_n9447_), .Y(new_n28694_));
  AOI21X1  g26258(.A0(new_n28694_), .A1(new_n28693_), .B0(po1038), .Y(new_n28695_));
  NAND2X1  g26259(.A(new_n28677_), .B(new_n28529_), .Y(new_n28696_));
  OAI21X1  g26260(.A0(new_n28696_), .A1(new_n28695_), .B0(new_n28692_), .Y(new_n28697_));
  AOI21X1  g26261(.A0(new_n28697_), .A1(pi1134), .B0(new_n28686_), .Y(po0435));
  INVX1    g26262(.A(new_n26670_), .Y(new_n28699_));
  OAI21X1  g26263(.A0(new_n28038_), .A1(pi0958), .B0(new_n2702_), .Y(new_n28700_));
  AOI21X1  g26264(.A0(new_n28038_), .A1(new_n4626_), .B0(new_n28700_), .Y(new_n28701_));
  AND3X1   g26265(.A(pi1135), .B(pi1091), .C(new_n7937_), .Y(new_n28702_));
  OAI21X1  g26266(.A0(new_n28702_), .A1(new_n28701_), .B0(pi0199), .Y(new_n28703_));
  NAND3X1  g26267(.A(new_n26508_), .B(pi0958), .C(pi0314), .Y(new_n28704_));
  AOI21X1  g26268(.A0(new_n28029_), .A1(pi0279), .B0(pi1091), .Y(new_n28705_));
  AND2X1   g26269(.A(new_n28705_), .B(new_n28704_), .Y(new_n28706_));
  AND3X1   g26270(.A(new_n28667_), .B(pi1091), .C(new_n7937_), .Y(new_n28707_));
  OR3X1    g26271(.A(new_n28707_), .B(new_n28706_), .C(pi0199), .Y(new_n28708_));
  AOI21X1  g26272(.A0(new_n28708_), .A1(new_n28703_), .B0(new_n22572_), .Y(new_n28709_));
  INVX1    g26273(.A(new_n28706_), .Y(new_n28710_));
  OAI21X1  g26274(.A0(new_n28667_), .A1(pi0211), .B0(pi1091), .Y(new_n28711_));
  AOI21X1  g26275(.A0(new_n28711_), .A1(new_n28710_), .B0(pi0219), .Y(new_n28712_));
  OAI21X1  g26276(.A0(new_n27747_), .A1(new_n4622_), .B0(pi0219), .Y(new_n28713_));
  OAI21X1  g26277(.A0(new_n28713_), .A1(new_n28701_), .B0(new_n22572_), .Y(new_n28714_));
  OAI21X1  g26278(.A0(new_n28714_), .A1(new_n28712_), .B0(new_n24814_), .Y(new_n28715_));
  AOI21X1  g26279(.A0(new_n28709_), .A1(new_n28699_), .B0(new_n28715_), .Y(new_n28716_));
  MX2X1    g26280(.A(new_n4622_), .B(new_n28667_), .S0(new_n7871_), .Y(new_n28717_));
  AND3X1   g26281(.A(pi1135), .B(pi0219), .C(new_n23173_), .Y(new_n28718_));
  NOR2X1   g26282(.A(pi1133), .B(pi0211), .Y(new_n28719_));
  NOR2X1   g26283(.A(new_n28719_), .B(pi0219), .Y(new_n28720_));
  AOI21X1  g26284(.A0(new_n28720_), .A1(new_n23173_), .B0(new_n28718_), .Y(new_n28721_));
  OAI22X1  g26285(.A0(new_n28721_), .A1(new_n2933_), .B0(new_n28717_), .B1(new_n24917_), .Y(new_n28722_));
  OAI21X1  g26286(.A0(new_n28721_), .A1(new_n6489_), .B0(pi0230), .Y(new_n28723_));
  AOI21X1  g26287(.A0(new_n28722_), .A1(new_n6489_), .B0(new_n28723_), .Y(new_n28724_));
  OAI21X1  g26288(.A0(new_n28724_), .A1(new_n28716_), .B0(new_n4747_), .Y(new_n28725_));
  NOR3X1   g26289(.A(pi1133), .B(pi0200), .C(pi0199), .Y(new_n28726_));
  AOI21X1  g26290(.A0(pi1135), .A1(new_n7937_), .B0(new_n7871_), .Y(new_n28727_));
  OAI21X1  g26291(.A0(new_n28727_), .A1(new_n28726_), .B0(new_n11660_), .Y(new_n28728_));
  OR3X1    g26292(.A(new_n28720_), .B(new_n28718_), .C(new_n11660_), .Y(new_n28729_));
  AOI21X1  g26293(.A0(new_n28729_), .A1(new_n28728_), .B0(new_n24814_), .Y(new_n28730_));
  NOR4X1   g26294(.A(new_n28719_), .B(new_n11660_), .C(new_n2702_), .D(pi0219), .Y(new_n28731_));
  NOR3X1   g26295(.A(new_n28731_), .B(new_n28715_), .C(new_n28709_), .Y(new_n28732_));
  OAI21X1  g26296(.A0(new_n28732_), .A1(new_n28730_), .B0(pi1134), .Y(new_n28733_));
  AND2X1   g26297(.A(new_n28733_), .B(new_n28725_), .Y(po0436));
  MX2X1    g26298(.A(new_n4554_), .B(new_n4622_), .S0(new_n23173_), .Y(new_n28735_));
  NAND2X1  g26299(.A(new_n28735_), .B(pi1091), .Y(new_n28736_));
  AOI21X1  g26300(.A0(new_n28028_), .A1(pi0914), .B0(pi1091), .Y(new_n28737_));
  OAI21X1  g26301(.A0(new_n28028_), .A1(pi0280), .B0(new_n28737_), .Y(new_n28738_));
  AOI21X1  g26302(.A0(new_n28738_), .A1(new_n28736_), .B0(pi0219), .Y(new_n28739_));
  AOI21X1  g26303(.A0(pi1137), .A1(new_n23173_), .B0(new_n8422_), .Y(new_n28740_));
  OR2X1    g26304(.A(new_n28740_), .B(new_n28071_), .Y(new_n28741_));
  AOI21X1  g26305(.A0(new_n28038_), .A1(pi0280), .B0(pi1091), .Y(new_n28742_));
  OAI21X1  g26306(.A0(new_n28038_), .A1(pi0914), .B0(new_n28742_), .Y(new_n28743_));
  AOI21X1  g26307(.A0(new_n28743_), .A1(new_n28741_), .B0(new_n28739_), .Y(new_n28744_));
  AND3X1   g26308(.A(pi1137), .B(pi1091), .C(new_n7937_), .Y(new_n28745_));
  INVX1    g26309(.A(new_n28745_), .Y(new_n28746_));
  AOI21X1  g26310(.A0(new_n28746_), .A1(new_n28743_), .B0(new_n7871_), .Y(new_n28747_));
  AOI21X1  g26311(.A0(pi1135), .A1(new_n7937_), .B0(new_n2702_), .Y(new_n28748_));
  OAI21X1  g26312(.A0(new_n4554_), .A1(new_n7937_), .B0(new_n28748_), .Y(new_n28749_));
  AND3X1   g26313(.A(new_n28749_), .B(new_n28738_), .C(new_n7871_), .Y(new_n28750_));
  OR2X1    g26314(.A(new_n28750_), .B(new_n22572_), .Y(new_n28751_));
  OAI22X1  g26315(.A0(new_n28751_), .A1(new_n28747_), .B0(new_n28744_), .B1(new_n11660_), .Y(new_n28752_));
  AOI21X1  g26316(.A0(pi1136), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n28753_));
  OAI21X1  g26317(.A0(new_n4622_), .A1(pi0199), .B0(new_n7937_), .Y(new_n28754_));
  AOI21X1  g26318(.A0(pi1137), .A1(pi0199), .B0(new_n28754_), .Y(new_n28755_));
  OR3X1    g26319(.A(new_n28755_), .B(new_n28753_), .C(new_n22572_), .Y(new_n28756_));
  AOI21X1  g26320(.A0(new_n28735_), .A1(new_n8422_), .B0(new_n28740_), .Y(new_n28757_));
  AOI21X1  g26321(.A0(new_n28757_), .A1(new_n22572_), .B0(new_n24814_), .Y(new_n28758_));
  AOI22X1  g26322(.A0(new_n28758_), .A1(new_n28756_), .B0(new_n28752_), .B1(new_n24814_), .Y(po0437));
  AOI21X1  g26323(.A0(pi1138), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n28760_));
  NAND2X1  g26324(.A(pi1139), .B(pi0199), .Y(new_n28761_));
  AOI21X1  g26325(.A0(pi1137), .A1(new_n7871_), .B0(pi0200), .Y(new_n28762_));
  AOI21X1  g26326(.A0(new_n28762_), .A1(new_n28761_), .B0(new_n28760_), .Y(new_n28763_));
  OR3X1    g26327(.A(new_n4019_), .B(new_n8422_), .C(pi0211), .Y(new_n28764_));
  MX2X1    g26328(.A(new_n4205_), .B(new_n4351_), .S0(new_n23173_), .Y(new_n28765_));
  OAI21X1  g26329(.A0(new_n28765_), .A1(pi0219), .B0(new_n28764_), .Y(new_n28766_));
  MX2X1    g26330(.A(new_n28766_), .B(new_n28763_), .S0(new_n11660_), .Y(new_n28767_));
  OR2X1    g26331(.A(new_n28029_), .B(pi0830), .Y(new_n28768_));
  AOI21X1  g26332(.A0(new_n28029_), .A1(pi0281), .B0(pi1091), .Y(new_n28769_));
  OAI21X1  g26333(.A0(new_n28765_), .A1(new_n2702_), .B0(new_n26027_), .Y(new_n28770_));
  AND3X1   g26334(.A(pi1138), .B(pi1091), .C(pi0200), .Y(new_n28771_));
  OR3X1    g26335(.A(new_n28771_), .B(new_n28745_), .C(new_n28396_), .Y(new_n28772_));
  AOI22X1  g26336(.A0(new_n28772_), .A1(new_n28770_), .B0(new_n28769_), .B1(new_n28768_), .Y(new_n28773_));
  AOI21X1  g26337(.A0(new_n28038_), .A1(pi0281), .B0(pi1091), .Y(new_n28774_));
  OAI21X1  g26338(.A0(new_n28038_), .A1(pi0830), .B0(new_n28774_), .Y(new_n28775_));
  AND3X1   g26339(.A(pi1139), .B(pi1091), .C(new_n23173_), .Y(new_n28776_));
  OR2X1    g26340(.A(new_n28398_), .B(new_n7871_), .Y(new_n28777_));
  OAI22X1  g26341(.A0(new_n28777_), .A1(new_n22572_), .B0(new_n28776_), .B1(new_n28377_), .Y(new_n28778_));
  AOI21X1  g26342(.A0(new_n28778_), .A1(new_n28775_), .B0(new_n28773_), .Y(new_n28779_));
  MX2X1    g26343(.A(new_n28779_), .B(new_n28767_), .S0(pi0230), .Y(po0438));
  AOI21X1  g26344(.A0(pi1139), .A1(new_n7871_), .B0(new_n7937_), .Y(new_n28781_));
  NAND2X1  g26345(.A(pi1140), .B(pi0199), .Y(new_n28782_));
  AOI21X1  g26346(.A0(pi1138), .A1(new_n7871_), .B0(pi0200), .Y(new_n28783_));
  AOI21X1  g26347(.A0(new_n28783_), .A1(new_n28782_), .B0(new_n28781_), .Y(new_n28784_));
  OR3X1    g26348(.A(new_n3908_), .B(new_n8422_), .C(pi0211), .Y(new_n28785_));
  MX2X1    g26349(.A(new_n4019_), .B(new_n4205_), .S0(new_n23173_), .Y(new_n28786_));
  OAI21X1  g26350(.A0(new_n28786_), .A1(pi0219), .B0(new_n28785_), .Y(new_n28787_));
  MX2X1    g26351(.A(new_n28787_), .B(new_n28784_), .S0(new_n11660_), .Y(new_n28788_));
  OR2X1    g26352(.A(new_n28029_), .B(pi0836), .Y(new_n28789_));
  AOI21X1  g26353(.A0(new_n28029_), .A1(pi0282), .B0(pi1091), .Y(new_n28790_));
  OAI21X1  g26354(.A0(new_n28786_), .A1(new_n2702_), .B0(new_n26027_), .Y(new_n28791_));
  AND3X1   g26355(.A(pi1139), .B(pi1091), .C(pi0200), .Y(new_n28792_));
  OR3X1    g26356(.A(new_n28792_), .B(new_n28378_), .C(new_n28396_), .Y(new_n28793_));
  AOI22X1  g26357(.A0(new_n28793_), .A1(new_n28791_), .B0(new_n28790_), .B1(new_n28789_), .Y(new_n28794_));
  AOI21X1  g26358(.A0(new_n28038_), .A1(pi0282), .B0(pi1091), .Y(new_n28795_));
  OAI21X1  g26359(.A0(new_n28038_), .A1(pi0836), .B0(new_n28795_), .Y(new_n28796_));
  AND3X1   g26360(.A(pi1140), .B(pi1091), .C(new_n23173_), .Y(new_n28797_));
  OAI21X1  g26361(.A0(new_n28635_), .A1(pi0200), .B0(pi0199), .Y(new_n28798_));
  OAI22X1  g26362(.A0(new_n28798_), .A1(new_n22572_), .B0(new_n28797_), .B1(new_n28377_), .Y(new_n28799_));
  AOI21X1  g26363(.A0(new_n28799_), .A1(new_n28796_), .B0(new_n28794_), .Y(new_n28800_));
  MX2X1    g26364(.A(new_n28800_), .B(new_n28788_), .S0(pi0230), .Y(po0439));
  OR2X1    g26365(.A(new_n28457_), .B(new_n25993_), .Y(new_n28802_));
  AND3X1   g26366(.A(new_n28802_), .B(new_n28463_), .C(pi1149), .Y(new_n28803_));
  OR2X1    g26367(.A(new_n28341_), .B(new_n25993_), .Y(new_n28804_));
  AND3X1   g26368(.A(new_n28804_), .B(new_n28349_), .C(new_n25955_), .Y(new_n28805_));
  OR3X1    g26369(.A(new_n28805_), .B(new_n28803_), .C(new_n26084_), .Y(new_n28806_));
  OAI22X1  g26370(.A0(new_n28457_), .A1(new_n25993_), .B0(new_n27521_), .B1(new_n25955_), .Y(new_n28807_));
  AOI21X1  g26371(.A0(new_n28807_), .A1(new_n26084_), .B0(new_n24814_), .Y(new_n28808_));
  OAI21X1  g26372(.A0(new_n28447_), .A1(pi1147), .B0(new_n26084_), .Y(new_n28809_));
  AOI21X1  g26373(.A0(new_n28442_), .A1(pi1147), .B0(new_n28809_), .Y(new_n28810_));
  NOR2X1   g26374(.A(new_n28327_), .B(pi1147), .Y(new_n28811_));
  OAI21X1  g26375(.A0(new_n28293_), .A1(new_n25993_), .B0(pi1148), .Y(new_n28812_));
  OAI21X1  g26376(.A0(new_n28812_), .A1(new_n28811_), .B0(pi1149), .Y(new_n28813_));
  AOI21X1  g26377(.A0(new_n28335_), .A1(new_n25993_), .B0(pi1148), .Y(new_n28814_));
  OAI21X1  g26378(.A0(new_n28266_), .A1(new_n25993_), .B0(new_n28814_), .Y(new_n28815_));
  NAND2X1  g26379(.A(new_n28333_), .B(new_n25993_), .Y(new_n28816_));
  AOI21X1  g26380(.A0(new_n28270_), .A1(pi1147), .B0(new_n26084_), .Y(new_n28817_));
  AOI21X1  g26381(.A0(new_n28817_), .A1(new_n28816_), .B0(pi1149), .Y(new_n28818_));
  AOI21X1  g26382(.A0(new_n28818_), .A1(new_n28815_), .B0(new_n28446_), .Y(new_n28819_));
  OAI21X1  g26383(.A0(new_n28813_), .A1(new_n28810_), .B0(new_n28819_), .Y(new_n28820_));
  OR3X1    g26384(.A(new_n28298_), .B(new_n28273_), .C(new_n25993_), .Y(new_n28821_));
  NAND3X1  g26385(.A(new_n28311_), .B(new_n28309_), .C(new_n25993_), .Y(new_n28822_));
  AND3X1   g26386(.A(new_n28822_), .B(new_n28821_), .C(pi1149), .Y(new_n28823_));
  AND3X1   g26387(.A(new_n28279_), .B(new_n28276_), .C(pi1147), .Y(new_n28824_));
  OAI21X1  g26388(.A0(new_n28283_), .A1(pi1147), .B0(new_n25955_), .Y(new_n28825_));
  OAI21X1  g26389(.A0(new_n28825_), .A1(new_n28824_), .B0(new_n26084_), .Y(new_n28826_));
  AOI21X1  g26390(.A0(new_n28284_), .A1(pi1147), .B0(pi1149), .Y(new_n28827_));
  OAI21X1  g26391(.A0(new_n28319_), .A1(pi1147), .B0(new_n28827_), .Y(new_n28828_));
  NAND2X1  g26392(.A(new_n28314_), .B(new_n25993_), .Y(new_n28829_));
  AOI21X1  g26393(.A0(new_n28304_), .A1(pi1147), .B0(new_n25955_), .Y(new_n28830_));
  AOI21X1  g26394(.A0(new_n28830_), .A1(new_n28829_), .B0(new_n26084_), .Y(new_n28831_));
  AOI21X1  g26395(.A0(new_n28831_), .A1(new_n28828_), .B0(pi0283), .Y(new_n28832_));
  OAI21X1  g26396(.A0(new_n28826_), .A1(new_n28823_), .B0(new_n28832_), .Y(new_n28833_));
  AND2X1   g26397(.A(new_n28833_), .B(new_n24814_), .Y(new_n28834_));
  AOI22X1  g26398(.A0(new_n28834_), .A1(new_n28820_), .B0(new_n28808_), .B1(new_n28806_), .Y(po0440));
  NAND2X1  g26399(.A(new_n27865_), .B(pi1143), .Y(new_n28836_));
  OAI22X1  g26400(.A0(new_n28836_), .A1(new_n26028_), .B0(new_n27865_), .B1(pi0284), .Y(po0441));
  INVX1    g26401(.A(pi0286), .Y(new_n28838_));
  NOR4X1   g26402(.A(new_n7786_), .B(new_n10077_), .C(new_n3105_), .D(new_n28838_), .Y(new_n28839_));
  AND3X1   g26403(.A(new_n28839_), .B(pi0289), .C(pi0288), .Y(new_n28840_));
  AND2X1   g26404(.A(new_n28840_), .B(pi0285), .Y(new_n28841_));
  NOR2X1   g26405(.A(new_n7786_), .B(new_n3105_), .Y(new_n28842_));
  AOI21X1  g26406(.A0(new_n28842_), .A1(pi0285), .B0(new_n28840_), .Y(new_n28843_));
  OR3X1    g26407(.A(new_n28843_), .B(new_n28841_), .C(po1038), .Y(new_n28844_));
  NAND4X1  g26408(.A(new_n28839_), .B(new_n6489_), .C(pi0289), .D(pi0288), .Y(new_n28845_));
  OR4X1    g26409(.A(new_n10124_), .B(pi0289), .C(pi0288), .D(pi0286), .Y(new_n28846_));
  NAND3X1  g26410(.A(new_n28846_), .B(new_n28845_), .C(pi0285), .Y(new_n28847_));
  AOI21X1  g26411(.A0(new_n28847_), .A1(new_n28844_), .B0(pi0793), .Y(po0442));
  NOR3X1   g26412(.A(pi0289), .B(pi0286), .C(pi0285), .Y(new_n28849_));
  NOR2X1   g26413(.A(new_n28849_), .B(pi0288), .Y(new_n28850_));
  INVX1    g26414(.A(new_n28842_), .Y(new_n28851_));
  AOI21X1  g26415(.A0(new_n28851_), .A1(new_n10077_), .B0(new_n28838_), .Y(new_n28852_));
  NOR3X1   g26416(.A(new_n28842_), .B(new_n10124_), .C(pi0286), .Y(new_n28853_));
  OAI21X1  g26417(.A0(new_n28853_), .A1(new_n28852_), .B0(new_n28850_), .Y(new_n28854_));
  OAI21X1  g26418(.A0(new_n28851_), .A1(new_n10077_), .B0(new_n28838_), .Y(new_n28855_));
  INVX1    g26419(.A(pi0288), .Y(new_n28856_));
  NOR2X1   g26420(.A(new_n28839_), .B(new_n28856_), .Y(new_n28857_));
  AOI21X1  g26421(.A0(new_n28857_), .A1(new_n28855_), .B0(po1038), .Y(new_n28858_));
  INVX1    g26422(.A(pi0793), .Y(new_n28859_));
  NAND3X1  g26423(.A(new_n28850_), .B(new_n6246_), .C(new_n2702_), .Y(new_n28860_));
  AND2X1   g26424(.A(new_n28860_), .B(pi0286), .Y(new_n28861_));
  OAI21X1  g26425(.A0(new_n28860_), .A1(pi0286), .B0(po1038), .Y(new_n28862_));
  OAI21X1  g26426(.A0(new_n28862_), .A1(new_n28861_), .B0(new_n28859_), .Y(new_n28863_));
  AOI21X1  g26427(.A0(new_n28858_), .A1(new_n28854_), .B0(new_n28863_), .Y(po0443));
  AOI21X1  g26428(.A0(pi0457), .A1(new_n7795_), .B0(pi0332), .Y(po0444));
  OAI21X1  g26429(.A0(new_n10077_), .A1(new_n28856_), .B0(new_n28860_), .Y(new_n28866_));
  NOR3X1   g26430(.A(new_n7786_), .B(po1038), .C(new_n3105_), .Y(po0637));
  OAI21X1  g26431(.A0(po0637), .A1(new_n28866_), .B0(new_n28859_), .Y(new_n28868_));
  AOI21X1  g26432(.A0(po0637), .A1(new_n28866_), .B0(new_n28868_), .Y(po0445));
  OR3X1    g26433(.A(new_n28839_), .B(pi0289), .C(new_n28856_), .Y(new_n28870_));
  INVX1    g26434(.A(pi0285), .Y(new_n28871_));
  OR2X1    g26435(.A(pi0289), .B(new_n28871_), .Y(new_n28872_));
  OR4X1    g26436(.A(new_n28872_), .B(new_n28842_), .C(new_n10124_), .D(pi0286), .Y(new_n28873_));
  INVX1    g26437(.A(new_n28853_), .Y(new_n28874_));
  AOI21X1  g26438(.A0(new_n28874_), .A1(pi0289), .B0(pi0288), .Y(new_n28875_));
  AOI21X1  g26439(.A0(new_n28875_), .A1(new_n28873_), .B0(new_n28840_), .Y(new_n28876_));
  AOI21X1  g26440(.A0(new_n28876_), .A1(new_n28870_), .B0(po1038), .Y(new_n28877_));
  AND3X1   g26441(.A(new_n10077_), .B(new_n28856_), .C(new_n28838_), .Y(new_n28878_));
  INVX1    g26442(.A(new_n28878_), .Y(new_n28879_));
  AND2X1   g26443(.A(new_n28879_), .B(pi0289), .Y(new_n28880_));
  OAI21X1  g26444(.A0(new_n28872_), .A1(new_n28879_), .B0(po1038), .Y(new_n28881_));
  OAI21X1  g26445(.A0(new_n28881_), .A1(new_n28880_), .B0(new_n28859_), .Y(new_n28882_));
  NOR2X1   g26446(.A(new_n28882_), .B(new_n28877_), .Y(po0446));
  MX2X1    g26447(.A(pi1048), .B(pi0290), .S0(pi0476), .Y(po0447));
  MX2X1    g26448(.A(pi1049), .B(pi0291), .S0(pi0476), .Y(po0448));
  MX2X1    g26449(.A(pi1084), .B(pi0292), .S0(pi0476), .Y(po0449));
  MX2X1    g26450(.A(pi1059), .B(pi0293), .S0(pi0476), .Y(po0450));
  MX2X1    g26451(.A(pi1072), .B(pi0294), .S0(pi0476), .Y(po0451));
  MX2X1    g26452(.A(pi1053), .B(pi0295), .S0(pi0476), .Y(po0452));
  MX2X1    g26453(.A(pi1037), .B(pi0296), .S0(pi0476), .Y(po0453));
  MX2X1    g26454(.A(pi1044), .B(pi0297), .S0(pi0476), .Y(po0454));
  MX2X1    g26455(.A(pi1044), .B(pi0298), .S0(pi0478), .Y(po0455));
  OR3X1    g26456(.A(new_n2985_), .B(new_n2536_), .C(new_n3091_), .Y(new_n28893_));
  NAND4X1  g26457(.A(new_n9677_), .B(new_n7606_), .C(new_n2497_), .D(new_n3091_), .Y(new_n28894_));
  NAND2X1  g26458(.A(new_n6721_), .B(new_n3088_), .Y(new_n28895_));
  AOI21X1  g26459(.A0(new_n28894_), .A1(new_n28893_), .B0(new_n28895_), .Y(new_n28896_));
  MX2X1    g26460(.A(new_n28896_), .B(new_n8352_), .S0(pi0039), .Y(po0456));
  INVX1    g26461(.A(pi0300), .Y(new_n28898_));
  NAND3X1  g26462(.A(new_n8375_), .B(new_n3127_), .C(pi0057), .Y(new_n28899_));
  NOR2X1   g26463(.A(new_n28899_), .B(pi0312), .Y(new_n28900_));
  AOI21X1  g26464(.A0(new_n28900_), .A1(new_n28898_), .B0(pi0055), .Y(new_n28901_));
  OAI21X1  g26465(.A0(new_n28900_), .A1(new_n28898_), .B0(new_n28901_), .Y(po0457));
  INVX1    g26466(.A(pi0301), .Y(new_n28903_));
  AND2X1   g26467(.A(new_n28901_), .B(new_n28903_), .Y(new_n28904_));
  OR2X1    g26468(.A(new_n28903_), .B(pi0055), .Y(new_n28905_));
  NOR4X1   g26469(.A(new_n28905_), .B(new_n28899_), .C(pi0312), .D(pi0300), .Y(new_n28906_));
  OR2X1    g26470(.A(new_n28906_), .B(new_n28904_), .Y(po0458));
  NOR4X1   g26471(.A(new_n5103_), .B(new_n4770_), .C(new_n2943_), .D(pi0057), .Y(new_n28908_));
  NOR2X1   g26472(.A(pi0223), .B(pi0222), .Y(new_n28909_));
  INVX1    g26473(.A(new_n28909_), .Y(new_n28910_));
  AOI22X1  g26474(.A0(new_n28910_), .A1(pi0937), .B0(new_n3138_), .B1(pi0273), .Y(new_n28911_));
  AND2X1   g26475(.A(new_n28911_), .B(new_n28908_), .Y(new_n28912_));
  NOR3X1   g26476(.A(new_n11660_), .B(new_n10045_), .C(pi0215), .Y(new_n28913_));
  OAI21X1  g26477(.A0(new_n28913_), .A1(new_n28912_), .B0(pi0237), .Y(new_n28914_));
  AOI21X1  g26478(.A0(new_n22572_), .A1(new_n4844_), .B0(new_n28908_), .Y(new_n28915_));
  NAND2X1  g26479(.A(new_n28915_), .B(new_n26084_), .Y(new_n28916_));
  OR4X1    g26480(.A(pi0273), .B(pi0221), .C(new_n2438_), .D(pi0215), .Y(new_n28917_));
  NOR4X1   g26481(.A(new_n2701_), .B(new_n2437_), .C(pi0216), .D(pi0215), .Y(new_n28918_));
  INVX1    g26482(.A(new_n28918_), .Y(new_n28919_));
  OAI21X1  g26483(.A0(new_n28919_), .A1(pi0937), .B0(new_n28917_), .Y(new_n28920_));
  AOI22X1  g26484(.A0(new_n28920_), .A1(new_n22572_), .B0(new_n28912_), .B1(new_n2952_), .Y(new_n28921_));
  AND3X1   g26485(.A(new_n28921_), .B(new_n28916_), .C(new_n28914_), .Y(po0459));
  MX2X1    g26486(.A(pi1049), .B(pi0303), .S0(pi0478), .Y(po0460));
  MX2X1    g26487(.A(pi1048), .B(pi0304), .S0(pi0478), .Y(po0461));
  MX2X1    g26488(.A(pi1084), .B(pi0305), .S0(pi0478), .Y(po0462));
  MX2X1    g26489(.A(pi1059), .B(pi0306), .S0(pi0478), .Y(po0463));
  MX2X1    g26490(.A(pi1053), .B(pi0307), .S0(pi0478), .Y(po0464));
  MX2X1    g26491(.A(pi1037), .B(pi0308), .S0(pi0478), .Y(po0465));
  MX2X1    g26492(.A(pi1072), .B(pi0309), .S0(pi0478), .Y(po0466));
  AND2X1   g26493(.A(new_n28915_), .B(pi1147), .Y(new_n28930_));
  OR4X1    g26494(.A(new_n11660_), .B(new_n4761_), .C(new_n10044_), .D(pi0215), .Y(new_n28931_));
  AOI22X1  g26495(.A0(new_n3152_), .A1(pi0271), .B0(new_n3019_), .B1(pi0934), .Y(new_n28932_));
  INVX1    g26496(.A(pi0934), .Y(new_n28933_));
  AOI22X1  g26497(.A0(new_n3138_), .A1(new_n26500_), .B0(new_n28933_), .B1(pi0222), .Y(new_n28934_));
  AOI21X1  g26498(.A0(new_n28934_), .A1(new_n28908_), .B0(new_n28913_), .Y(new_n28935_));
  OAI21X1  g26499(.A0(new_n28932_), .A1(new_n28931_), .B0(new_n28935_), .Y(new_n28936_));
  OAI21X1  g26500(.A0(new_n28936_), .A1(new_n28930_), .B0(new_n22655_), .Y(new_n28937_));
  NAND3X1  g26501(.A(new_n28932_), .B(new_n22572_), .C(new_n4844_), .Y(new_n28938_));
  INVX1    g26502(.A(new_n28908_), .Y(new_n28939_));
  OAI21X1  g26503(.A0(new_n28934_), .A1(new_n28939_), .B0(pi1147), .Y(new_n28940_));
  AOI21X1  g26504(.A0(new_n11660_), .A1(new_n2990_), .B0(new_n28940_), .Y(new_n28941_));
  OAI21X1  g26505(.A0(new_n28939_), .A1(new_n2951_), .B0(new_n28931_), .Y(new_n28942_));
  AND3X1   g26506(.A(new_n28942_), .B(new_n28936_), .C(new_n25993_), .Y(new_n28943_));
  AOI21X1  g26507(.A0(new_n28941_), .A1(new_n28938_), .B0(new_n28943_), .Y(new_n28944_));
  OAI21X1  g26508(.A0(new_n28944_), .A1(new_n22655_), .B0(new_n28937_), .Y(po0467));
  NOR2X1   g26509(.A(pi0311), .B(pi0055), .Y(new_n28946_));
  MX2X1    g26510(.A(new_n28946_), .B(pi0311), .S0(new_n28906_), .Y(po0468));
  XOR2X1   g26511(.A(new_n28899_), .B(pi0312), .Y(new_n28948_));
  NOR2X1   g26512(.A(new_n28948_), .B(pi0055), .Y(po0469));
  AOI21X1  g26513(.A0(new_n9704_), .A1(po0740), .B0(new_n9441_), .Y(new_n28950_));
  OAI21X1  g26514(.A0(new_n9699_), .A1(new_n7776_), .B0(new_n28950_), .Y(po0634));
  AND2X1   g26515(.A(pi0954), .B(pi0313), .Y(new_n28952_));
  AOI21X1  g26516(.A0(po0634), .A1(po1110), .B0(new_n28952_), .Y(po0470));
  NAND4X1  g26517(.A(new_n6720_), .B(new_n5299_), .C(new_n4982_), .D(new_n3107_), .Y(new_n28954_));
  NAND2X1  g26518(.A(new_n28954_), .B(new_n11099_), .Y(new_n28955_));
  OAI21X1  g26519(.A0(new_n10914_), .A1(new_n2939_), .B0(new_n3251_), .Y(new_n28956_));
  AOI21X1  g26520(.A0(new_n10846_), .A1(new_n2939_), .B0(new_n28956_), .Y(new_n28957_));
  AND3X1   g26521(.A(new_n7607_), .B(new_n3077_), .C(new_n3079_), .Y(new_n28958_));
  OAI21X1  g26522(.A0(new_n28957_), .A1(new_n11401_), .B0(new_n28958_), .Y(new_n28959_));
  NAND2X1  g26523(.A(new_n10337_), .B(new_n10335_), .Y(new_n28960_));
  AOI21X1  g26524(.A0(new_n28959_), .A1(new_n28955_), .B0(new_n28960_), .Y(po0471));
  OR4X1    g26525(.A(new_n7786_), .B(po1038), .C(new_n3105_), .D(pi0340), .Y(new_n28962_));
  MX2X1    g26526(.A(pi1080), .B(pi0315), .S0(new_n28962_), .Y(po0472));
  MX2X1    g26527(.A(pi1047), .B(pi0316), .S0(new_n28962_), .Y(po0473));
  OR4X1    g26528(.A(new_n7786_), .B(po1038), .C(new_n3105_), .D(pi0330), .Y(new_n28965_));
  MX2X1    g26529(.A(pi1078), .B(pi0317), .S0(new_n28965_), .Y(po0474));
  OR4X1    g26530(.A(new_n7786_), .B(po1038), .C(new_n3105_), .D(pi0341), .Y(new_n28967_));
  MX2X1    g26531(.A(pi1074), .B(pi0318), .S0(new_n28967_), .Y(po0475));
  MX2X1    g26532(.A(pi1072), .B(pi0319), .S0(new_n28967_), .Y(po0476));
  MX2X1    g26533(.A(pi1048), .B(pi0320), .S0(new_n28962_), .Y(po0477));
  MX2X1    g26534(.A(pi1058), .B(pi0321), .S0(new_n28962_), .Y(po0478));
  MX2X1    g26535(.A(pi1051), .B(pi0322), .S0(new_n28962_), .Y(po0479));
  MX2X1    g26536(.A(pi1065), .B(pi0323), .S0(new_n28962_), .Y(po0480));
  MX2X1    g26537(.A(pi1086), .B(pi0324), .S0(new_n28967_), .Y(po0481));
  MX2X1    g26538(.A(pi1063), .B(pi0325), .S0(new_n28967_), .Y(po0482));
  MX2X1    g26539(.A(pi1057), .B(pi0326), .S0(new_n28967_), .Y(po0483));
  MX2X1    g26540(.A(pi1040), .B(pi0327), .S0(new_n28962_), .Y(po0484));
  MX2X1    g26541(.A(pi1058), .B(pi0328), .S0(new_n28967_), .Y(po0485));
  MX2X1    g26542(.A(pi1043), .B(pi0329), .S0(new_n28967_), .Y(po0486));
  NOR3X1   g26543(.A(new_n6489_), .B(new_n2759_), .C(new_n5024_), .Y(new_n28980_));
  INVX1    g26544(.A(new_n28980_), .Y(new_n28981_));
  NOR2X1   g26545(.A(new_n2759_), .B(new_n5024_), .Y(new_n28982_));
  NAND2X1  g26546(.A(new_n28982_), .B(new_n6489_), .Y(new_n28983_));
  MX2X1    g26547(.A(pi0330), .B(pi0340), .S0(new_n28842_), .Y(new_n28984_));
  OAI22X1  g26548(.A0(new_n28984_), .A1(new_n28983_), .B0(new_n28981_), .B1(pi0330), .Y(po0487));
  MX2X1    g26549(.A(pi0331), .B(pi0341), .S0(new_n28842_), .Y(new_n28986_));
  OAI22X1  g26550(.A0(new_n28986_), .A1(new_n28983_), .B0(new_n28981_), .B1(pi0331), .Y(po0488));
  NOR3X1   g26551(.A(new_n8179_), .B(new_n8243_), .C(pi0332), .Y(new_n28988_));
  AOI21X1  g26552(.A0(new_n9475_), .A1(new_n8179_), .B0(new_n5898_), .Y(new_n28989_));
  OR2X1    g26553(.A(new_n28989_), .B(pi0070), .Y(new_n28990_));
  AND3X1   g26554(.A(new_n28990_), .B(new_n7216_), .C(pi0332), .Y(new_n28991_));
  OAI21X1  g26555(.A0(new_n28991_), .A1(new_n28988_), .B0(new_n2939_), .Y(new_n28992_));
  AOI21X1  g26556(.A0(new_n7796_), .A1(pi0039), .B0(pi0038), .Y(new_n28993_));
  AOI21X1  g26557(.A0(new_n28993_), .A1(new_n28992_), .B0(new_n24723_), .Y(po0489));
  MX2X1    g26558(.A(pi1040), .B(pi0333), .S0(new_n28967_), .Y(po0490));
  MX2X1    g26559(.A(pi1065), .B(pi0334), .S0(new_n28967_), .Y(po0491));
  MX2X1    g26560(.A(pi1069), .B(pi0335), .S0(new_n28967_), .Y(po0492));
  MX2X1    g26561(.A(pi1070), .B(pi0336), .S0(new_n28965_), .Y(po0493));
  MX2X1    g26562(.A(pi1044), .B(pi0337), .S0(new_n28965_), .Y(po0494));
  MX2X1    g26563(.A(pi1072), .B(pi0338), .S0(new_n28965_), .Y(po0495));
  MX2X1    g26564(.A(pi1086), .B(pi0339), .S0(new_n28965_), .Y(po0496));
  OR2X1    g26565(.A(new_n28842_), .B(pi0340), .Y(new_n29002_));
  NOR3X1   g26566(.A(new_n7786_), .B(new_n3105_), .C(pi0331), .Y(new_n29003_));
  NOR2X1   g26567(.A(new_n29003_), .B(new_n28983_), .Y(new_n29004_));
  AOI22X1  g26568(.A0(new_n29004_), .A1(new_n29002_), .B0(new_n28980_), .B1(pi0340), .Y(po0497));
  OAI21X1  g26569(.A0(po0637), .A1(pi0341), .B0(new_n28965_), .Y(new_n29006_));
  AND2X1   g26570(.A(new_n29006_), .B(new_n28982_), .Y(po0498));
  MX2X1    g26571(.A(pi1049), .B(pi0342), .S0(new_n28962_), .Y(po0499));
  MX2X1    g26572(.A(pi1062), .B(pi0343), .S0(new_n28962_), .Y(po0500));
  MX2X1    g26573(.A(pi1069), .B(pi0344), .S0(new_n28962_), .Y(po0501));
  MX2X1    g26574(.A(pi1039), .B(pi0345), .S0(new_n28962_), .Y(po0502));
  MX2X1    g26575(.A(pi1067), .B(pi0346), .S0(new_n28962_), .Y(po0503));
  MX2X1    g26576(.A(pi1055), .B(pi0347), .S0(new_n28962_), .Y(po0504));
  MX2X1    g26577(.A(pi1087), .B(pi0348), .S0(new_n28962_), .Y(po0505));
  MX2X1    g26578(.A(pi1043), .B(pi0349), .S0(new_n28962_), .Y(po0506));
  MX2X1    g26579(.A(pi1035), .B(pi0350), .S0(new_n28962_), .Y(po0507));
  MX2X1    g26580(.A(pi1079), .B(pi0351), .S0(new_n28962_), .Y(po0508));
  MX2X1    g26581(.A(pi1078), .B(pi0352), .S0(new_n28962_), .Y(po0509));
  MX2X1    g26582(.A(pi1063), .B(pi0353), .S0(new_n28962_), .Y(po0510));
  MX2X1    g26583(.A(pi1045), .B(pi0354), .S0(new_n28962_), .Y(po0511));
  MX2X1    g26584(.A(pi1084), .B(pi0355), .S0(new_n28962_), .Y(po0512));
  MX2X1    g26585(.A(pi1081), .B(pi0356), .S0(new_n28962_), .Y(po0513));
  MX2X1    g26586(.A(pi1076), .B(pi0357), .S0(new_n28962_), .Y(po0514));
  MX2X1    g26587(.A(pi1071), .B(pi0358), .S0(new_n28962_), .Y(po0515));
  MX2X1    g26588(.A(pi1068), .B(pi0359), .S0(new_n28962_), .Y(po0516));
  MX2X1    g26589(.A(pi1042), .B(pi0360), .S0(new_n28962_), .Y(po0517));
  MX2X1    g26590(.A(pi1059), .B(pi0361), .S0(new_n28962_), .Y(po0518));
  MX2X1    g26591(.A(pi1070), .B(pi0362), .S0(new_n28962_), .Y(po0519));
  MX2X1    g26592(.A(pi1049), .B(pi0363), .S0(new_n28965_), .Y(po0520));
  MX2X1    g26593(.A(pi1062), .B(pi0364), .S0(new_n28965_), .Y(po0521));
  MX2X1    g26594(.A(pi1065), .B(pi0365), .S0(new_n28965_), .Y(po0522));
  MX2X1    g26595(.A(pi1069), .B(pi0366), .S0(new_n28965_), .Y(po0523));
  MX2X1    g26596(.A(pi1039), .B(pi0367), .S0(new_n28965_), .Y(po0524));
  MX2X1    g26597(.A(pi1067), .B(pi0368), .S0(new_n28965_), .Y(po0525));
  MX2X1    g26598(.A(pi1080), .B(pi0369), .S0(new_n28965_), .Y(po0526));
  MX2X1    g26599(.A(pi1055), .B(pi0370), .S0(new_n28965_), .Y(po0527));
  MX2X1    g26600(.A(pi1051), .B(pi0371), .S0(new_n28965_), .Y(po0528));
  MX2X1    g26601(.A(pi1048), .B(pi0372), .S0(new_n28965_), .Y(po0529));
  MX2X1    g26602(.A(pi1087), .B(pi0373), .S0(new_n28965_), .Y(po0530));
  MX2X1    g26603(.A(pi1035), .B(pi0374), .S0(new_n28965_), .Y(po0531));
  MX2X1    g26604(.A(pi1047), .B(pi0375), .S0(new_n28965_), .Y(po0532));
  MX2X1    g26605(.A(pi1079), .B(pi0376), .S0(new_n28965_), .Y(po0533));
  MX2X1    g26606(.A(pi1074), .B(pi0377), .S0(new_n28965_), .Y(po0534));
  MX2X1    g26607(.A(pi1063), .B(pi0378), .S0(new_n28965_), .Y(po0535));
  MX2X1    g26608(.A(pi1045), .B(pi0379), .S0(new_n28965_), .Y(po0536));
  MX2X1    g26609(.A(pi1084), .B(pi0380), .S0(new_n28965_), .Y(po0537));
  MX2X1    g26610(.A(pi1081), .B(pi0381), .S0(new_n28965_), .Y(po0538));
  MX2X1    g26611(.A(pi1076), .B(pi0382), .S0(new_n28965_), .Y(po0539));
  MX2X1    g26612(.A(pi1071), .B(pi0383), .S0(new_n28965_), .Y(po0540));
  MX2X1    g26613(.A(pi1068), .B(pi0384), .S0(new_n28965_), .Y(po0541));
  MX2X1    g26614(.A(pi1042), .B(pi0385), .S0(new_n28965_), .Y(po0542));
  MX2X1    g26615(.A(pi1059), .B(pi0386), .S0(new_n28965_), .Y(po0543));
  MX2X1    g26616(.A(pi1053), .B(pi0387), .S0(new_n28965_), .Y(po0544));
  MX2X1    g26617(.A(pi1037), .B(pi0388), .S0(new_n28965_), .Y(po0545));
  MX2X1    g26618(.A(pi1036), .B(pi0389), .S0(new_n28965_), .Y(po0546));
  MX2X1    g26619(.A(pi1049), .B(pi0390), .S0(new_n28967_), .Y(po0547));
  MX2X1    g26620(.A(pi1062), .B(pi0391), .S0(new_n28967_), .Y(po0548));
  MX2X1    g26621(.A(pi1039), .B(pi0392), .S0(new_n28967_), .Y(po0549));
  MX2X1    g26622(.A(pi1067), .B(pi0393), .S0(new_n28967_), .Y(po0550));
  MX2X1    g26623(.A(pi1080), .B(pi0394), .S0(new_n28967_), .Y(po0551));
  MX2X1    g26624(.A(pi1055), .B(pi0395), .S0(new_n28967_), .Y(po0552));
  MX2X1    g26625(.A(pi1051), .B(pi0396), .S0(new_n28967_), .Y(po0553));
  MX2X1    g26626(.A(pi1048), .B(pi0397), .S0(new_n28967_), .Y(po0554));
  MX2X1    g26627(.A(pi1087), .B(pi0398), .S0(new_n28967_), .Y(po0555));
  MX2X1    g26628(.A(pi1047), .B(pi0399), .S0(new_n28967_), .Y(po0556));
  MX2X1    g26629(.A(pi1035), .B(pi0400), .S0(new_n28967_), .Y(po0557));
  MX2X1    g26630(.A(pi1079), .B(pi0401), .S0(new_n28967_), .Y(po0558));
  MX2X1    g26631(.A(pi1078), .B(pi0402), .S0(new_n28967_), .Y(po0559));
  MX2X1    g26632(.A(pi1045), .B(pi0403), .S0(new_n28967_), .Y(po0560));
  MX2X1    g26633(.A(pi1084), .B(pi0404), .S0(new_n28967_), .Y(po0561));
  MX2X1    g26634(.A(pi1081), .B(pi0405), .S0(new_n28967_), .Y(po0562));
  MX2X1    g26635(.A(pi1076), .B(pi0406), .S0(new_n28967_), .Y(po0563));
  MX2X1    g26636(.A(pi1071), .B(pi0407), .S0(new_n28967_), .Y(po0564));
  MX2X1    g26637(.A(pi1068), .B(pi0408), .S0(new_n28967_), .Y(po0565));
  MX2X1    g26638(.A(pi1042), .B(pi0409), .S0(new_n28967_), .Y(po0566));
  MX2X1    g26639(.A(pi1059), .B(pi0410), .S0(new_n28967_), .Y(po0567));
  MX2X1    g26640(.A(pi1053), .B(pi0411), .S0(new_n28967_), .Y(po0568));
  MX2X1    g26641(.A(pi1037), .B(pi0412), .S0(new_n28967_), .Y(po0569));
  MX2X1    g26642(.A(pi1036), .B(pi0413), .S0(new_n28967_), .Y(po0570));
  OR4X1    g26643(.A(new_n7786_), .B(po1038), .C(new_n3105_), .D(pi0331), .Y(new_n29080_));
  MX2X1    g26644(.A(pi1049), .B(pi0414), .S0(new_n29080_), .Y(po0571));
  MX2X1    g26645(.A(pi1062), .B(pi0415), .S0(new_n29080_), .Y(po0572));
  MX2X1    g26646(.A(pi1069), .B(pi0416), .S0(new_n29080_), .Y(po0573));
  MX2X1    g26647(.A(pi1039), .B(pi0417), .S0(new_n29080_), .Y(po0574));
  MX2X1    g26648(.A(pi1067), .B(pi0418), .S0(new_n29080_), .Y(po0575));
  MX2X1    g26649(.A(pi1080), .B(pi0419), .S0(new_n29080_), .Y(po0576));
  MX2X1    g26650(.A(pi1055), .B(pi0420), .S0(new_n29080_), .Y(po0577));
  MX2X1    g26651(.A(pi1051), .B(pi0421), .S0(new_n29080_), .Y(po0578));
  MX2X1    g26652(.A(pi1048), .B(pi0422), .S0(new_n29080_), .Y(po0579));
  MX2X1    g26653(.A(pi1087), .B(pi0423), .S0(new_n29080_), .Y(po0580));
  MX2X1    g26654(.A(pi1047), .B(pi0424), .S0(new_n29080_), .Y(po0581));
  MX2X1    g26655(.A(pi1035), .B(pi0425), .S0(new_n29080_), .Y(po0582));
  MX2X1    g26656(.A(pi1079), .B(pi0426), .S0(new_n29080_), .Y(po0583));
  MX2X1    g26657(.A(pi1078), .B(pi0427), .S0(new_n29080_), .Y(po0584));
  MX2X1    g26658(.A(pi1045), .B(pi0428), .S0(new_n29080_), .Y(po0585));
  MX2X1    g26659(.A(pi1084), .B(pi0429), .S0(new_n29080_), .Y(po0586));
  MX2X1    g26660(.A(pi1076), .B(pi0430), .S0(new_n29080_), .Y(po0587));
  MX2X1    g26661(.A(pi1071), .B(pi0431), .S0(new_n29080_), .Y(po0588));
  MX2X1    g26662(.A(pi1068), .B(pi0432), .S0(new_n29080_), .Y(po0589));
  MX2X1    g26663(.A(pi1042), .B(pi0433), .S0(new_n29080_), .Y(po0590));
  MX2X1    g26664(.A(pi1059), .B(pi0434), .S0(new_n29080_), .Y(po0591));
  MX2X1    g26665(.A(pi1053), .B(pi0435), .S0(new_n29080_), .Y(po0592));
  MX2X1    g26666(.A(pi1037), .B(pi0436), .S0(new_n29080_), .Y(po0593));
  MX2X1    g26667(.A(pi1070), .B(pi0437), .S0(new_n29080_), .Y(po0594));
  MX2X1    g26668(.A(pi1036), .B(pi0438), .S0(new_n29080_), .Y(po0595));
  MX2X1    g26669(.A(pi1057), .B(pi0439), .S0(new_n28965_), .Y(po0596));
  MX2X1    g26670(.A(pi1043), .B(pi0440), .S0(new_n28965_), .Y(po0597));
  MX2X1    g26671(.A(pi1044), .B(pi0441), .S0(new_n28962_), .Y(po0598));
  MX2X1    g26672(.A(pi1058), .B(pi0442), .S0(new_n28965_), .Y(po0599));
  MX2X1    g26673(.A(pi1044), .B(pi0443), .S0(new_n29080_), .Y(po0600));
  MX2X1    g26674(.A(pi1072), .B(pi0444), .S0(new_n29080_), .Y(po0601));
  MX2X1    g26675(.A(pi1081), .B(pi0445), .S0(new_n29080_), .Y(po0602));
  MX2X1    g26676(.A(pi1086), .B(pi0446), .S0(new_n29080_), .Y(po0603));
  MX2X1    g26677(.A(pi1040), .B(pi0447), .S0(new_n28965_), .Y(po0604));
  MX2X1    g26678(.A(pi1074), .B(pi0448), .S0(new_n29080_), .Y(po0605));
  MX2X1    g26679(.A(pi1057), .B(pi0449), .S0(new_n29080_), .Y(po0606));
  MX2X1    g26680(.A(pi1036), .B(pi0450), .S0(new_n28962_), .Y(po0607));
  MX2X1    g26681(.A(pi1063), .B(pi0451), .S0(new_n29080_), .Y(po0608));
  MX2X1    g26682(.A(pi1053), .B(pi0452), .S0(new_n28962_), .Y(po0609));
  MX2X1    g26683(.A(pi1040), .B(pi0453), .S0(new_n29080_), .Y(po0610));
  MX2X1    g26684(.A(pi1043), .B(pi0454), .S0(new_n29080_), .Y(po0611));
  MX2X1    g26685(.A(pi1037), .B(pi0455), .S0(new_n28962_), .Y(po0612));
  MX2X1    g26686(.A(pi1044), .B(pi0456), .S0(new_n28967_), .Y(po0613));
  INVX1    g26687(.A(pi0821), .Y(new_n29124_));
  NAND4X1  g26688(.A(pi0601), .B(pi0600), .C(pi0597), .D(pi0594), .Y(new_n29125_));
  OR3X1    g26689(.A(pi0810), .B(pi0804), .C(pi0595), .Y(new_n29126_));
  INVX1    g26690(.A(pi0804), .Y(new_n29127_));
  INVX1    g26691(.A(pi0596), .Y(new_n29128_));
  INVX1    g26692(.A(pi0599), .Y(new_n29129_));
  AOI21X1  g26693(.A0(pi0810), .A1(new_n29129_), .B0(new_n29128_), .Y(new_n29130_));
  AND2X1   g26694(.A(pi0815), .B(pi0595), .Y(new_n29131_));
  OAI21X1  g26695(.A0(new_n29130_), .A1(new_n29127_), .B0(new_n29131_), .Y(new_n29132_));
  AOI21X1  g26696(.A0(new_n29132_), .A1(new_n29126_), .B0(new_n29125_), .Y(new_n29133_));
  INVX1    g26697(.A(pi0815), .Y(new_n29134_));
  INVX1    g26698(.A(pi0600), .Y(new_n29135_));
  OAI21X1  g26699(.A0(pi0810), .A1(new_n29135_), .B0(pi0804), .Y(new_n29136_));
  NOR2X1   g26700(.A(pi0810), .B(pi0804), .Y(new_n29137_));
  OR2X1    g26701(.A(new_n29137_), .B(pi0601), .Y(new_n29138_));
  AND3X1   g26702(.A(new_n29138_), .B(new_n29136_), .C(new_n29134_), .Y(new_n29139_));
  OAI21X1  g26703(.A0(new_n29139_), .A1(new_n29133_), .B0(pi0605), .Y(new_n29140_));
  NAND3X1  g26704(.A(pi0990), .B(pi0600), .C(pi0594), .Y(new_n29141_));
  OR3X1    g26705(.A(new_n29141_), .B(new_n29136_), .C(pi0815), .Y(new_n29142_));
  AOI21X1  g26706(.A0(new_n29142_), .A1(new_n29140_), .B0(new_n29124_), .Y(po0614));
  MX2X1    g26707(.A(pi1072), .B(pi0458), .S0(new_n28962_), .Y(po0615));
  MX2X1    g26708(.A(pi1058), .B(pi0459), .S0(new_n29080_), .Y(po0616));
  MX2X1    g26709(.A(pi1086), .B(pi0460), .S0(new_n28962_), .Y(po0617));
  MX2X1    g26710(.A(pi1057), .B(pi0461), .S0(new_n28962_), .Y(po0618));
  MX2X1    g26711(.A(pi1074), .B(pi0462), .S0(new_n28962_), .Y(po0619));
  MX2X1    g26712(.A(pi1070), .B(pi0463), .S0(new_n28967_), .Y(po0620));
  MX2X1    g26713(.A(pi1065), .B(pi0464), .S0(new_n29080_), .Y(po0621));
  OR2X1    g26714(.A(new_n4771_), .B(new_n4762_), .Y(new_n29151_));
  AND2X1   g26715(.A(new_n29151_), .B(pi0926), .Y(new_n29152_));
  OAI21X1  g26716(.A0(new_n8437_), .A1(new_n8435_), .B0(new_n26499_), .Y(new_n29153_));
  OAI21X1  g26717(.A0(new_n29151_), .A1(new_n12578_), .B0(new_n29153_), .Y(new_n29154_));
  AOI22X1  g26718(.A0(new_n28909_), .A1(new_n2933_), .B0(new_n4889_), .B1(new_n2437_), .Y(new_n29155_));
  AOI21X1  g26719(.A0(pi1157), .A1(new_n26499_), .B0(new_n29155_), .Y(new_n29156_));
  OAI21X1  g26720(.A0(new_n8455_), .A1(pi0216), .B0(new_n3261_), .Y(new_n29157_));
  AND3X1   g26721(.A(pi1157), .B(pi0926), .C(new_n26499_), .Y(new_n29158_));
  AOI22X1  g26722(.A0(new_n29158_), .A1(new_n29157_), .B0(new_n29156_), .B1(new_n29153_), .Y(new_n29159_));
  OAI21X1  g26723(.A0(new_n29154_), .A1(new_n29152_), .B0(new_n29159_), .Y(new_n29160_));
  AND3X1   g26724(.A(new_n2437_), .B(pi0216), .C(new_n2934_), .Y(new_n29161_));
  AOI21X1  g26725(.A0(new_n29161_), .A1(new_n26499_), .B0(new_n6489_), .Y(new_n29162_));
  AOI22X1  g26726(.A0(new_n28918_), .A1(pi0926), .B0(new_n4845_), .B1(pi1157), .Y(new_n29163_));
  AOI22X1  g26727(.A0(new_n29163_), .A1(new_n29162_), .B0(new_n29160_), .B1(new_n6489_), .Y(po0622));
  OR2X1    g26728(.A(new_n29161_), .B(new_n6489_), .Y(new_n29165_));
  OR4X1    g26729(.A(new_n8437_), .B(new_n8435_), .C(new_n5103_), .D(pi0057), .Y(new_n29166_));
  AND2X1   g26730(.A(new_n29166_), .B(new_n29165_), .Y(new_n29167_));
  MX2X1    g26731(.A(new_n29167_), .B(new_n28942_), .S0(pi0943), .Y(new_n29168_));
  OR2X1    g26732(.A(new_n29168_), .B(pi1151), .Y(new_n29169_));
  OR3X1    g26733(.A(new_n29167_), .B(new_n28915_), .C(pi0943), .Y(new_n29170_));
  MX2X1    g26734(.A(new_n3242_), .B(new_n2990_), .S0(new_n11660_), .Y(new_n29171_));
  AND3X1   g26735(.A(new_n29171_), .B(pi1151), .C(pi0943), .Y(new_n29172_));
  OR2X1    g26736(.A(new_n6489_), .B(new_n3019_), .Y(new_n29173_));
  OAI21X1  g26737(.A0(new_n29155_), .A1(po1038), .B0(new_n29173_), .Y(new_n29174_));
  AOI21X1  g26738(.A0(new_n29174_), .A1(new_n28581_), .B0(new_n29172_), .Y(new_n29175_));
  AND3X1   g26739(.A(new_n29175_), .B(new_n29170_), .C(new_n29169_), .Y(po0623));
  NOR4X1   g26740(.A(new_n27497_), .B(new_n27496_), .C(pi0287), .D(new_n2529_), .Y(new_n29177_));
  AOI21X1  g26741(.A0(new_n29177_), .A1(po0950), .B0(new_n7608_), .Y(new_n29178_));
  NOR3X1   g26742(.A(new_n11774_), .B(new_n8243_), .C(new_n6738_), .Y(new_n29179_));
  OAI21X1  g26743(.A0(new_n9655_), .A1(pi0102), .B0(new_n29179_), .Y(new_n29180_));
  NOR3X1   g26744(.A(new_n29180_), .B(new_n2582_), .C(pi0098), .Y(new_n29181_));
  INVX1    g26745(.A(new_n29181_), .Y(new_n29182_));
  XOR2X1   g26746(.A(new_n29182_), .B(new_n29177_), .Y(new_n29183_));
  MX2X1    g26747(.A(new_n29183_), .B(new_n29182_), .S0(new_n5882_), .Y(new_n29184_));
  NOR2X1   g26748(.A(new_n29184_), .B(new_n5970_), .Y(new_n29185_));
  INVX1    g26749(.A(new_n5970_), .Y(new_n29186_));
  OAI21X1  g26750(.A0(new_n29183_), .A1(new_n29186_), .B0(pi1091), .Y(new_n29187_));
  NOR2X1   g26751(.A(new_n29184_), .B(pi1093), .Y(new_n29188_));
  MX2X1    g26752(.A(new_n29183_), .B(new_n29182_), .S0(new_n5927_), .Y(new_n29189_));
  OAI21X1  g26753(.A0(new_n29189_), .A1(new_n5032_), .B0(new_n2702_), .Y(new_n29190_));
  OAI22X1  g26754(.A0(new_n29190_), .A1(new_n29188_), .B0(new_n29187_), .B1(new_n29185_), .Y(new_n29191_));
  NOR2X1   g26755(.A(new_n28954_), .B(new_n3074_), .Y(new_n29192_));
  AOI21X1  g26756(.A0(new_n29192_), .A1(new_n29191_), .B0(new_n29178_), .Y(po0624));
  NOR4X1   g26757(.A(new_n9483_), .B(new_n7553_), .C(pi0039), .D(new_n2979_), .Y(new_n29194_));
  OAI22X1  g26758(.A0(new_n29194_), .A1(new_n8621_), .B0(new_n8398_), .B1(new_n7629_), .Y(po0625));
  AND2X1   g26759(.A(new_n29151_), .B(pi0942), .Y(new_n29196_));
  OAI21X1  g26760(.A0(new_n8437_), .A1(new_n8435_), .B0(new_n26599_), .Y(new_n29197_));
  OAI21X1  g26761(.A0(new_n29151_), .A1(new_n12555_), .B0(new_n29197_), .Y(new_n29198_));
  AOI21X1  g26762(.A0(pi1156), .A1(new_n26599_), .B0(new_n29155_), .Y(new_n29199_));
  AND3X1   g26763(.A(pi1156), .B(pi0942), .C(new_n26599_), .Y(new_n29200_));
  AOI22X1  g26764(.A0(new_n29200_), .A1(new_n29157_), .B0(new_n29199_), .B1(new_n29197_), .Y(new_n29201_));
  OAI21X1  g26765(.A0(new_n29198_), .A1(new_n29196_), .B0(new_n29201_), .Y(new_n29202_));
  AOI21X1  g26766(.A0(new_n29161_), .A1(new_n26599_), .B0(new_n6489_), .Y(new_n29203_));
  AOI22X1  g26767(.A0(new_n28918_), .A1(pi0942), .B0(new_n4845_), .B1(pi1156), .Y(new_n29204_));
  AOI22X1  g26768(.A0(new_n29204_), .A1(new_n29203_), .B0(new_n29202_), .B1(new_n6489_), .Y(po0626));
  AND2X1   g26769(.A(new_n29151_), .B(pi0925), .Y(new_n29206_));
  OAI21X1  g26770(.A0(new_n8437_), .A1(new_n8435_), .B0(pi0267), .Y(new_n29207_));
  OAI21X1  g26771(.A0(new_n29151_), .A1(new_n12463_), .B0(new_n29207_), .Y(new_n29208_));
  AOI21X1  g26772(.A0(pi1155), .A1(pi0267), .B0(new_n29155_), .Y(new_n29209_));
  AND3X1   g26773(.A(pi1155), .B(pi0925), .C(pi0267), .Y(new_n29210_));
  AOI22X1  g26774(.A0(new_n29210_), .A1(new_n29157_), .B0(new_n29209_), .B1(new_n29207_), .Y(new_n29211_));
  OAI21X1  g26775(.A0(new_n29208_), .A1(new_n29206_), .B0(new_n29211_), .Y(new_n29212_));
  AOI21X1  g26776(.A0(new_n29161_), .A1(pi0267), .B0(new_n6489_), .Y(new_n29213_));
  AOI22X1  g26777(.A0(new_n28918_), .A1(pi0925), .B0(new_n4845_), .B1(pi1155), .Y(new_n29214_));
  AOI22X1  g26778(.A0(new_n29214_), .A1(new_n29213_), .B0(new_n29212_), .B1(new_n6489_), .Y(po0627));
  AND2X1   g26779(.A(new_n29151_), .B(pi0941), .Y(new_n29216_));
  OAI21X1  g26780(.A0(new_n8437_), .A1(new_n8435_), .B0(pi0253), .Y(new_n29217_));
  OAI21X1  g26781(.A0(new_n29151_), .A1(new_n12364_), .B0(new_n29217_), .Y(new_n29218_));
  AOI21X1  g26782(.A0(pi1153), .A1(pi0253), .B0(new_n29155_), .Y(new_n29219_));
  AND3X1   g26783(.A(pi1153), .B(pi0941), .C(pi0253), .Y(new_n29220_));
  AOI22X1  g26784(.A0(new_n29220_), .A1(new_n29157_), .B0(new_n29219_), .B1(new_n29217_), .Y(new_n29221_));
  OAI21X1  g26785(.A0(new_n29218_), .A1(new_n29216_), .B0(new_n29221_), .Y(new_n29222_));
  AOI21X1  g26786(.A0(new_n29161_), .A1(pi0253), .B0(new_n6489_), .Y(new_n29223_));
  AOI22X1  g26787(.A0(new_n28918_), .A1(pi0941), .B0(new_n4845_), .B1(pi1153), .Y(new_n29224_));
  AOI22X1  g26788(.A0(new_n29224_), .A1(new_n29223_), .B0(new_n29222_), .B1(new_n6489_), .Y(po0628));
  AND2X1   g26789(.A(new_n29151_), .B(pi0923), .Y(new_n29226_));
  OAI21X1  g26790(.A0(new_n8437_), .A1(new_n8435_), .B0(pi0254), .Y(new_n29227_));
  OAI21X1  g26791(.A0(new_n29151_), .A1(new_n12487_), .B0(new_n29227_), .Y(new_n29228_));
  AOI21X1  g26792(.A0(pi1154), .A1(pi0254), .B0(new_n29155_), .Y(new_n29229_));
  AND3X1   g26793(.A(pi1154), .B(pi0923), .C(pi0254), .Y(new_n29230_));
  AOI22X1  g26794(.A0(new_n29230_), .A1(new_n29157_), .B0(new_n29229_), .B1(new_n29227_), .Y(new_n29231_));
  OAI21X1  g26795(.A0(new_n29228_), .A1(new_n29226_), .B0(new_n29231_), .Y(new_n29232_));
  AOI21X1  g26796(.A0(new_n29161_), .A1(pi0254), .B0(new_n6489_), .Y(new_n29233_));
  AOI22X1  g26797(.A0(new_n28918_), .A1(pi0923), .B0(new_n4845_), .B1(pi1154), .Y(new_n29234_));
  AOI22X1  g26798(.A0(new_n29234_), .A1(new_n29233_), .B0(new_n29232_), .B1(new_n6489_), .Y(po0629));
  MX2X1    g26799(.A(new_n29167_), .B(new_n28942_), .S0(pi0922), .Y(new_n29236_));
  OR2X1    g26800(.A(new_n29236_), .B(pi1152), .Y(new_n29237_));
  OR3X1    g26801(.A(new_n29167_), .B(new_n28915_), .C(pi0922), .Y(new_n29238_));
  AND3X1   g26802(.A(new_n29171_), .B(pi1152), .C(pi0922), .Y(new_n29239_));
  AOI21X1  g26803(.A0(new_n29174_), .A1(new_n28297_), .B0(new_n29239_), .Y(new_n29240_));
  AND3X1   g26804(.A(new_n29240_), .B(new_n29238_), .C(new_n29237_), .Y(po0630));
  MX2X1    g26805(.A(new_n29167_), .B(new_n28942_), .S0(pi0931), .Y(new_n29242_));
  OR2X1    g26806(.A(new_n29242_), .B(pi1150), .Y(new_n29243_));
  OR3X1    g26807(.A(new_n29167_), .B(new_n28915_), .C(pi0931), .Y(new_n29244_));
  AND3X1   g26808(.A(new_n29171_), .B(pi1150), .C(pi0931), .Y(new_n29245_));
  AOI21X1  g26809(.A0(new_n29174_), .A1(new_n28455_), .B0(new_n29245_), .Y(new_n29246_));
  AND3X1   g26810(.A(new_n29246_), .B(new_n29244_), .C(new_n29243_), .Y(po0631));
  MX2X1    g26811(.A(new_n29167_), .B(new_n28942_), .S0(pi0936), .Y(new_n29248_));
  OR2X1    g26812(.A(new_n29248_), .B(pi1149), .Y(new_n29249_));
  OR3X1    g26813(.A(new_n29167_), .B(new_n28915_), .C(pi0936), .Y(new_n29250_));
  AND3X1   g26814(.A(new_n29171_), .B(pi1149), .C(pi0936), .Y(new_n29251_));
  AOI21X1  g26815(.A0(new_n29174_), .A1(new_n28446_), .B0(new_n29251_), .Y(new_n29252_));
  AND3X1   g26816(.A(new_n29252_), .B(new_n29250_), .C(new_n29249_), .Y(po0632));
  OR4X1    g26817(.A(new_n6489_), .B(pi0219), .C(new_n23173_), .D(new_n2590_), .Y(new_n29254_));
  NAND3X1  g26818(.A(new_n9438_), .B(new_n2595_), .C(new_n2594_), .Y(new_n29255_));
  NOR2X1   g26819(.A(new_n8469_), .B(new_n7601_), .Y(new_n29256_));
  AOI22X1  g26820(.A0(new_n29256_), .A1(new_n7600_), .B0(new_n9437_), .B1(new_n8469_), .Y(new_n29257_));
  NOR4X1   g26821(.A(new_n29257_), .B(new_n29255_), .C(new_n8243_), .D(new_n3105_), .Y(new_n29258_));
  AOI21X1  g26822(.A0(new_n8470_), .A1(pi0071), .B0(new_n29258_), .Y(new_n29259_));
  OAI21X1  g26823(.A0(new_n29259_), .A1(po1038), .B0(new_n29254_), .Y(po0633));
  NOR2X1   g26824(.A(new_n28457_), .B(new_n2590_), .Y(po0635));
  MX2X1    g26825(.A(pi0481), .B(pi0248), .S0(new_n22576_), .Y(po0638));
  MX2X1    g26826(.A(pi0482), .B(pi0249), .S0(new_n22587_), .Y(po0639));
  MX2X1    g26827(.A(pi0483), .B(pi0242), .S0(new_n22658_), .Y(po0640));
  MX2X1    g26828(.A(pi0484), .B(pi0249), .S0(new_n22658_), .Y(po0641));
  MX2X1    g26829(.A(pi0485), .B(pi0234), .S0(new_n23383_), .Y(po0642));
  MX2X1    g26830(.A(pi0486), .B(pi0244), .S0(new_n23383_), .Y(po0643));
  MX2X1    g26831(.A(pi0487), .B(pi0246), .S0(new_n22576_), .Y(po0644));
  INVX1    g26832(.A(pi0488), .Y(new_n29269_));
  MX2X1    g26833(.A(new_n29269_), .B(pi0239), .S0(new_n22576_), .Y(po0645));
  MX2X1    g26834(.A(pi0489), .B(pi0242), .S0(new_n23383_), .Y(po0646));
  MX2X1    g26835(.A(pi0490), .B(pi0241), .S0(new_n22658_), .Y(po0647));
  MX2X1    g26836(.A(pi0491), .B(pi0238), .S0(new_n22658_), .Y(po0648));
  MX2X1    g26837(.A(pi0492), .B(pi0240), .S0(new_n22658_), .Y(po0649));
  MX2X1    g26838(.A(pi0493), .B(pi0244), .S0(new_n22658_), .Y(po0650));
  INVX1    g26839(.A(pi0494), .Y(new_n29276_));
  MX2X1    g26840(.A(new_n29276_), .B(pi0239), .S0(new_n22658_), .Y(po0651));
  MX2X1    g26841(.A(pi0495), .B(pi0235), .S0(new_n22658_), .Y(po0652));
  MX2X1    g26842(.A(pi0496), .B(pi0249), .S0(new_n22652_), .Y(po0653));
  INVX1    g26843(.A(pi0497), .Y(new_n29280_));
  MX2X1    g26844(.A(new_n29280_), .B(pi0239), .S0(new_n22652_), .Y(po0654));
  MX2X1    g26845(.A(pi0498), .B(pi0238), .S0(new_n22587_), .Y(po0655));
  MX2X1    g26846(.A(pi0499), .B(pi0246), .S0(new_n22652_), .Y(po0656));
  MX2X1    g26847(.A(pi0500), .B(pi0241), .S0(new_n22652_), .Y(po0657));
  MX2X1    g26848(.A(pi0501), .B(pi0248), .S0(new_n22652_), .Y(po0658));
  MX2X1    g26849(.A(pi0502), .B(pi0247), .S0(new_n22652_), .Y(po0659));
  MX2X1    g26850(.A(pi0503), .B(pi0245), .S0(new_n22652_), .Y(po0660));
  MX2X1    g26851(.A(pi0504), .B(pi0242), .S0(new_n22648_), .Y(po0661));
  INVX1    g26852(.A(pi0505), .Y(new_n29289_));
  MX2X1    g26853(.A(new_n5197_), .B(new_n5105_), .S0(new_n22572_), .Y(new_n29290_));
  AND3X1   g26854(.A(new_n29290_), .B(new_n22652_), .C(new_n2973_), .Y(new_n29291_));
  OR4X1    g26855(.A(new_n22647_), .B(new_n22646_), .C(new_n22574_), .D(new_n2973_), .Y(new_n29292_));
  OR3X1    g26856(.A(pi0505), .B(new_n22579_), .C(pi0233), .Y(new_n29293_));
  OAI22X1  g26857(.A0(new_n29293_), .A1(new_n29292_), .B0(new_n29291_), .B1(new_n29289_), .Y(po0662));
  MX2X1    g26858(.A(pi0506), .B(pi0241), .S0(new_n22648_), .Y(po0663));
  MX2X1    g26859(.A(pi0507), .B(pi0238), .S0(new_n22648_), .Y(po0664));
  MX2X1    g26860(.A(pi0508), .B(pi0247), .S0(new_n22648_), .Y(po0665));
  MX2X1    g26861(.A(pi0509), .B(pi0245), .S0(new_n22648_), .Y(po0666));
  MX2X1    g26862(.A(pi0510), .B(pi0242), .S0(new_n22576_), .Y(po0667));
  AOI21X1  g26863(.A0(new_n6489_), .A1(new_n5339_), .B0(new_n22575_), .Y(new_n29300_));
  AND2X1   g26864(.A(new_n29300_), .B(new_n2973_), .Y(new_n29301_));
  INVX1    g26865(.A(new_n29301_), .Y(new_n29302_));
  MX2X1    g26866(.A(pi0511), .B(new_n29302_), .S0(new_n22576_), .Y(po0668));
  MX2X1    g26867(.A(pi0512), .B(pi0235), .S0(new_n22576_), .Y(po0669));
  MX2X1    g26868(.A(pi0513), .B(pi0244), .S0(new_n22576_), .Y(po0670));
  MX2X1    g26869(.A(pi0514), .B(pi0245), .S0(new_n22576_), .Y(po0671));
  MX2X1    g26870(.A(pi0515), .B(pi0240), .S0(new_n22576_), .Y(po0672));
  MX2X1    g26871(.A(pi0516), .B(pi0247), .S0(new_n22576_), .Y(po0673));
  MX2X1    g26872(.A(pi0517), .B(pi0238), .S0(new_n22576_), .Y(po0674));
  INVX1    g26873(.A(pi0518), .Y(new_n29310_));
  AND3X1   g26874(.A(new_n29300_), .B(new_n22582_), .C(new_n2973_), .Y(new_n29311_));
  OR4X1    g26875(.A(new_n22575_), .B(new_n22574_), .C(new_n22573_), .D(new_n2973_), .Y(new_n29312_));
  OR3X1    g26876(.A(pi0518), .B(new_n22579_), .C(pi0233), .Y(new_n29313_));
  OAI22X1  g26877(.A0(new_n29313_), .A1(new_n29312_), .B0(new_n29311_), .B1(new_n29310_), .Y(po0675));
  INVX1    g26878(.A(pi0519), .Y(new_n29315_));
  MX2X1    g26879(.A(new_n29315_), .B(pi0239), .S0(new_n22582_), .Y(po0676));
  MX2X1    g26880(.A(pi0520), .B(pi0246), .S0(new_n22582_), .Y(po0677));
  MX2X1    g26881(.A(pi0521), .B(pi0248), .S0(new_n22582_), .Y(po0678));
  MX2X1    g26882(.A(pi0522), .B(pi0238), .S0(new_n22582_), .Y(po0679));
  INVX1    g26883(.A(pi0523), .Y(new_n29320_));
  AND3X1   g26884(.A(new_n29300_), .B(new_n23398_), .C(new_n2973_), .Y(new_n29321_));
  OR3X1    g26885(.A(pi0523), .B(pi0237), .C(new_n22655_), .Y(new_n29322_));
  OAI22X1  g26886(.A0(new_n29322_), .A1(new_n29312_), .B0(new_n29321_), .B1(new_n29320_), .Y(po0680));
  INVX1    g26887(.A(pi0524), .Y(new_n29324_));
  MX2X1    g26888(.A(new_n29324_), .B(pi0239), .S0(new_n23398_), .Y(po0681));
  MX2X1    g26889(.A(pi0525), .B(pi0245), .S0(new_n23398_), .Y(po0682));
  MX2X1    g26890(.A(pi0526), .B(pi0246), .S0(new_n23398_), .Y(po0683));
  MX2X1    g26891(.A(pi0527), .B(pi0247), .S0(new_n23398_), .Y(po0684));
  MX2X1    g26892(.A(pi0528), .B(pi0249), .S0(new_n23398_), .Y(po0685));
  MX2X1    g26893(.A(pi0529), .B(pi0238), .S0(new_n23398_), .Y(po0686));
  MX2X1    g26894(.A(pi0530), .B(pi0240), .S0(new_n23398_), .Y(po0687));
  MX2X1    g26895(.A(pi0531), .B(pi0235), .S0(new_n22587_), .Y(po0688));
  MX2X1    g26896(.A(pi0532), .B(pi0247), .S0(new_n22587_), .Y(po0689));
  MX2X1    g26897(.A(pi0533), .B(pi0235), .S0(new_n22648_), .Y(po0690));
  INVX1    g26898(.A(pi0534), .Y(new_n29335_));
  MX2X1    g26899(.A(new_n29335_), .B(pi0239), .S0(new_n22648_), .Y(po0691));
  MX2X1    g26900(.A(pi0535), .B(pi0240), .S0(new_n22648_), .Y(po0692));
  MX2X1    g26901(.A(pi0536), .B(pi0246), .S0(new_n22648_), .Y(po0693));
  MX2X1    g26902(.A(pi0537), .B(pi0248), .S0(new_n22648_), .Y(po0694));
  MX2X1    g26903(.A(pi0538), .B(pi0249), .S0(new_n22648_), .Y(po0695));
  MX2X1    g26904(.A(pi0539), .B(pi0242), .S0(new_n22652_), .Y(po0696));
  MX2X1    g26905(.A(pi0540), .B(pi0235), .S0(new_n22652_), .Y(po0697));
  MX2X1    g26906(.A(pi0541), .B(pi0244), .S0(new_n22652_), .Y(po0698));
  MX2X1    g26907(.A(pi0542), .B(pi0240), .S0(new_n22652_), .Y(po0699));
  MX2X1    g26908(.A(pi0543), .B(pi0238), .S0(new_n22652_), .Y(po0700));
  INVX1    g26909(.A(pi0544), .Y(new_n29346_));
  AND3X1   g26910(.A(new_n29290_), .B(new_n22658_), .C(new_n2973_), .Y(new_n29347_));
  OR3X1    g26911(.A(pi0544), .B(pi0237), .C(new_n22655_), .Y(new_n29348_));
  OAI22X1  g26912(.A0(new_n29348_), .A1(new_n29292_), .B0(new_n29347_), .B1(new_n29346_), .Y(po0701));
  MX2X1    g26913(.A(pi0545), .B(pi0245), .S0(new_n22658_), .Y(po0702));
  MX2X1    g26914(.A(pi0546), .B(pi0246), .S0(new_n22658_), .Y(po0703));
  MX2X1    g26915(.A(pi0547), .B(pi0247), .S0(new_n22658_), .Y(po0704));
  MX2X1    g26916(.A(pi0548), .B(pi0248), .S0(new_n22658_), .Y(po0705));
  MX2X1    g26917(.A(pi0549), .B(pi0235), .S0(new_n23383_), .Y(po0706));
  INVX1    g26918(.A(pi0550), .Y(new_n29355_));
  MX2X1    g26919(.A(new_n29355_), .B(pi0239), .S0(new_n23383_), .Y(po0707));
  MX2X1    g26920(.A(pi0551), .B(pi0240), .S0(new_n23383_), .Y(po0708));
  MX2X1    g26921(.A(pi0552), .B(pi0247), .S0(new_n23383_), .Y(po0709));
  MX2X1    g26922(.A(pi0553), .B(pi0241), .S0(new_n23383_), .Y(po0710));
  MX2X1    g26923(.A(pi0554), .B(pi0248), .S0(new_n23383_), .Y(po0711));
  MX2X1    g26924(.A(pi0555), .B(pi0249), .S0(new_n23383_), .Y(po0712));
  MX2X1    g26925(.A(pi0556), .B(pi0242), .S0(new_n22587_), .Y(po0713));
  INVX1    g26926(.A(pi0557), .Y(new_n29363_));
  AND3X1   g26927(.A(new_n29290_), .B(new_n22648_), .C(new_n2973_), .Y(new_n29364_));
  OR2X1    g26928(.A(new_n22458_), .B(pi0557), .Y(new_n29365_));
  OAI22X1  g26929(.A0(new_n29365_), .A1(new_n29292_), .B0(new_n29364_), .B1(new_n29363_), .Y(po0714));
  MX2X1    g26930(.A(pi0558), .B(pi0244), .S0(new_n22648_), .Y(po0715));
  MX2X1    g26931(.A(pi0559), .B(pi0241), .S0(new_n22576_), .Y(po0716));
  MX2X1    g26932(.A(pi0560), .B(pi0240), .S0(new_n22587_), .Y(po0717));
  MX2X1    g26933(.A(pi0561), .B(pi0247), .S0(new_n22582_), .Y(po0718));
  MX2X1    g26934(.A(pi0562), .B(pi0241), .S0(new_n22587_), .Y(po0719));
  MX2X1    g26935(.A(pi0563), .B(pi0246), .S0(new_n23383_), .Y(po0720));
  MX2X1    g26936(.A(pi0564), .B(pi0246), .S0(new_n22587_), .Y(po0721));
  MX2X1    g26937(.A(pi0565), .B(pi0248), .S0(new_n22587_), .Y(po0722));
  MX2X1    g26938(.A(pi0566), .B(pi0244), .S0(new_n22587_), .Y(po0723));
  AND2X1   g26939(.A(pi1092), .B(new_n5979_), .Y(new_n29376_));
  NAND3X1  g26940(.A(new_n11979_), .B(new_n2720_), .C(pi0603), .Y(new_n29377_));
  NOR4X1   g26941(.A(new_n29377_), .B(new_n14039_), .C(new_n14034_), .D(new_n12473_), .Y(new_n29378_));
  AND3X1   g26942(.A(new_n5032_), .B(pi1092), .C(new_n5979_), .Y(new_n29379_));
  NOR3X1   g26943(.A(new_n29379_), .B(new_n29378_), .C(pi0789), .Y(new_n29380_));
  AND2X1   g26944(.A(new_n29378_), .B(new_n12509_), .Y(new_n29381_));
  OR2X1    g26945(.A(new_n29381_), .B(new_n29379_), .Y(new_n29382_));
  AOI21X1  g26946(.A0(new_n29378_), .A1(pi0619), .B0(new_n29379_), .Y(new_n29383_));
  OAI21X1  g26947(.A0(new_n29383_), .A1(new_n12510_), .B0(pi0789), .Y(new_n29384_));
  AOI21X1  g26948(.A0(new_n29382_), .A1(new_n12510_), .B0(new_n29384_), .Y(new_n29385_));
  NOR2X1   g26949(.A(new_n29385_), .B(new_n29380_), .Y(new_n29386_));
  INVX1    g26950(.A(new_n29379_), .Y(new_n29387_));
  OR4X1    g26951(.A(new_n13433_), .B(new_n12095_), .C(new_n2725_), .D(new_n5019_), .Y(new_n29388_));
  AND2X1   g26952(.A(new_n29388_), .B(new_n29387_), .Y(new_n29389_));
  OR3X1    g26953(.A(new_n29389_), .B(new_n12513_), .C(new_n12490_), .Y(new_n29390_));
  AOI21X1  g26954(.A0(new_n29385_), .A1(new_n16113_), .B0(new_n29390_), .Y(new_n29391_));
  OAI21X1  g26955(.A0(new_n29391_), .A1(new_n29386_), .B0(new_n12709_), .Y(new_n29392_));
  NOR4X1   g26956(.A(new_n29389_), .B(new_n12531_), .C(new_n12513_), .D(new_n12490_), .Y(new_n29393_));
  AOI21X1  g26957(.A0(new_n29393_), .A1(pi0641), .B0(new_n29379_), .Y(new_n29394_));
  AOI21X1  g26958(.A0(new_n29393_), .A1(new_n12543_), .B0(new_n29379_), .Y(new_n29395_));
  OAI22X1  g26959(.A0(new_n29395_), .A1(new_n14062_), .B0(new_n29394_), .B1(new_n14050_), .Y(new_n29396_));
  AOI21X1  g26960(.A0(new_n29386_), .A1(new_n22865_), .B0(new_n29396_), .Y(new_n29397_));
  OAI21X1  g26961(.A0(new_n29397_), .A1(new_n11765_), .B0(new_n29392_), .Y(new_n29398_));
  MX2X1    g26962(.A(new_n29386_), .B(new_n29379_), .S0(new_n12708_), .Y(new_n29399_));
  NAND2X1  g26963(.A(new_n29399_), .B(new_n12735_), .Y(new_n29400_));
  OR2X1    g26964(.A(new_n29389_), .B(new_n13489_), .Y(new_n29401_));
  OAI21X1  g26965(.A0(new_n29401_), .A1(new_n12554_), .B0(new_n29387_), .Y(new_n29402_));
  AOI21X1  g26966(.A0(new_n29402_), .A1(pi1156), .B0(pi0629), .Y(new_n29403_));
  NAND2X1  g26967(.A(new_n29403_), .B(new_n29400_), .Y(new_n29404_));
  NAND2X1  g26968(.A(new_n29399_), .B(new_n12733_), .Y(new_n29405_));
  OAI21X1  g26969(.A0(new_n29401_), .A1(pi0628), .B0(new_n29387_), .Y(new_n29406_));
  AOI21X1  g26970(.A0(new_n29406_), .A1(new_n12555_), .B0(new_n12561_), .Y(new_n29407_));
  AOI21X1  g26971(.A0(new_n29407_), .A1(new_n29405_), .B0(new_n11764_), .Y(new_n29408_));
  AOI22X1  g26972(.A0(new_n29408_), .A1(new_n29404_), .B0(new_n29398_), .B1(new_n14126_), .Y(new_n29409_));
  MX2X1    g26973(.A(new_n29399_), .B(new_n29379_), .S0(new_n12580_), .Y(new_n29410_));
  AOI21X1  g26974(.A0(new_n29410_), .A1(pi0647), .B0(pi1157), .Y(new_n29411_));
  OAI21X1  g26975(.A0(new_n29409_), .A1(pi0647), .B0(new_n29411_), .Y(new_n29412_));
  OR4X1    g26976(.A(new_n29389_), .B(new_n13508_), .C(new_n13489_), .D(new_n12577_), .Y(new_n29413_));
  NOR2X1   g26977(.A(new_n29379_), .B(new_n12578_), .Y(new_n29414_));
  AOI21X1  g26978(.A0(new_n29414_), .A1(new_n29413_), .B0(pi0630), .Y(new_n29415_));
  AOI21X1  g26979(.A0(new_n29410_), .A1(new_n12577_), .B0(new_n12578_), .Y(new_n29416_));
  OAI21X1  g26980(.A0(new_n29409_), .A1(new_n12577_), .B0(new_n29416_), .Y(new_n29417_));
  OR4X1    g26981(.A(new_n29389_), .B(new_n13508_), .C(new_n13489_), .D(pi0647), .Y(new_n29418_));
  NOR2X1   g26982(.A(new_n29379_), .B(pi1157), .Y(new_n29419_));
  AOI21X1  g26983(.A0(new_n29419_), .A1(new_n29418_), .B0(new_n12592_), .Y(new_n29420_));
  AOI22X1  g26984(.A0(new_n29420_), .A1(new_n29417_), .B0(new_n29415_), .B1(new_n29412_), .Y(new_n29421_));
  MX2X1    g26985(.A(new_n29421_), .B(new_n29409_), .S0(new_n11763_), .Y(new_n29422_));
  NOR4X1   g26986(.A(new_n29389_), .B(new_n13520_), .C(new_n13508_), .D(new_n13489_), .Y(new_n29423_));
  OR2X1    g26987(.A(new_n29423_), .B(new_n29379_), .Y(new_n29424_));
  AOI21X1  g26988(.A0(new_n29424_), .A1(pi0644), .B0(pi0715), .Y(new_n29425_));
  OAI21X1  g26989(.A0(new_n29422_), .A1(pi0644), .B0(new_n29425_), .Y(new_n29426_));
  NAND4X1  g26990(.A(new_n29399_), .B(new_n12605_), .C(new_n14327_), .D(new_n12612_), .Y(new_n29427_));
  NAND3X1  g26991(.A(new_n29427_), .B(new_n29387_), .C(pi0715), .Y(new_n29428_));
  AOI21X1  g26992(.A0(new_n29428_), .A1(new_n29426_), .B0(pi1160), .Y(new_n29429_));
  OAI21X1  g26993(.A0(new_n29424_), .A1(pi0644), .B0(pi0715), .Y(new_n29430_));
  AOI21X1  g26994(.A0(new_n29422_), .A1(pi0644), .B0(new_n29430_), .Y(new_n29431_));
  NAND4X1  g26995(.A(new_n29399_), .B(new_n12605_), .C(new_n14327_), .D(pi0644), .Y(new_n29432_));
  AOI21X1  g26996(.A0(new_n29432_), .A1(new_n29387_), .B0(pi0715), .Y(new_n29433_));
  OR2X1    g26997(.A(new_n29433_), .B(new_n11762_), .Y(new_n29434_));
  OAI21X1  g26998(.A0(new_n29434_), .A1(new_n29431_), .B0(pi0790), .Y(new_n29435_));
  OAI22X1  g26999(.A0(new_n29435_), .A1(new_n29429_), .B0(new_n29422_), .B1(pi0790), .Y(new_n29436_));
  MX2X1    g27000(.A(new_n29436_), .B(new_n29376_), .S0(new_n24814_), .Y(po0724));
  MX2X1    g27001(.A(pi0568), .B(pi0245), .S0(new_n22587_), .Y(po0725));
  INVX1    g27002(.A(pi0569), .Y(new_n29439_));
  MX2X1    g27003(.A(new_n29439_), .B(pi0239), .S0(new_n22587_), .Y(po0726));
  INVX1    g27004(.A(pi0570), .Y(new_n29441_));
  AND3X1   g27005(.A(new_n29300_), .B(new_n22587_), .C(new_n2973_), .Y(new_n29442_));
  OR3X1    g27006(.A(pi0570), .B(pi0237), .C(pi0233), .Y(new_n29443_));
  OAI22X1  g27007(.A0(new_n29443_), .A1(new_n29312_), .B0(new_n29442_), .B1(new_n29441_), .Y(po0727));
  MX2X1    g27008(.A(pi0571), .B(pi0241), .S0(new_n23398_), .Y(po0728));
  MX2X1    g27009(.A(pi0572), .B(pi0244), .S0(new_n23398_), .Y(po0729));
  MX2X1    g27010(.A(pi0573), .B(pi0242), .S0(new_n23398_), .Y(po0730));
  MX2X1    g27011(.A(pi0574), .B(pi0241), .S0(new_n22582_), .Y(po0731));
  MX2X1    g27012(.A(pi0575), .B(pi0235), .S0(new_n23398_), .Y(po0732));
  MX2X1    g27013(.A(pi0576), .B(pi0248), .S0(new_n23398_), .Y(po0733));
  MX2X1    g27014(.A(pi0577), .B(pi0238), .S0(new_n23383_), .Y(po0734));
  MX2X1    g27015(.A(pi0578), .B(pi0249), .S0(new_n22582_), .Y(po0735));
  MX2X1    g27016(.A(pi0579), .B(pi0249), .S0(new_n22576_), .Y(po0736));
  MX2X1    g27017(.A(pi0580), .B(pi0245), .S0(new_n23383_), .Y(po0737));
  MX2X1    g27018(.A(pi0581), .B(pi0235), .S0(new_n22582_), .Y(po0738));
  MX2X1    g27019(.A(pi0582), .B(pi0240), .S0(new_n22582_), .Y(po0739));
  MX2X1    g27020(.A(pi0584), .B(pi0245), .S0(new_n22582_), .Y(po0741));
  MX2X1    g27021(.A(pi0585), .B(pi0244), .S0(new_n22582_), .Y(po0742));
  MX2X1    g27022(.A(pi0586), .B(pi0242), .S0(new_n22582_), .Y(po0743));
  OR4X1    g27023(.A(new_n23093_), .B(new_n14034_), .C(new_n12048_), .D(new_n24814_), .Y(new_n29460_));
  OR4X1    g27024(.A(new_n29460_), .B(new_n16164_), .C(new_n14040_), .D(new_n12708_), .Y(new_n29461_));
  OAI21X1  g27025(.A0(new_n5354_), .A1(pi0230), .B0(new_n29461_), .Y(po0744));
  NAND2X1  g27026(.A(new_n8959_), .B(new_n27864_), .Y(new_n29463_));
  OAI21X1  g27027(.A0(new_n29463_), .A1(pi0591), .B0(new_n28982_), .Y(new_n29464_));
  AOI21X1  g27028(.A0(new_n29463_), .A1(new_n6603_), .B0(new_n29464_), .Y(po0745));
  NAND2X1  g27029(.A(new_n29290_), .B(new_n22589_), .Y(new_n29466_));
  AOI21X1  g27030(.A0(new_n29300_), .A1(new_n22457_), .B0(new_n22655_), .Y(new_n29467_));
  NAND2X1  g27031(.A(new_n29290_), .B(new_n22650_), .Y(new_n29468_));
  AOI21X1  g27032(.A0(new_n29300_), .A1(new_n22578_), .B0(pi0233), .Y(new_n29469_));
  AOI22X1  g27033(.A0(new_n29469_), .A1(new_n29468_), .B0(new_n29467_), .B1(new_n29466_), .Y(new_n29470_));
  NAND2X1  g27034(.A(new_n29290_), .B(new_n22654_), .Y(new_n29471_));
  AOI21X1  g27035(.A0(new_n29300_), .A1(new_n23396_), .B0(new_n22655_), .Y(new_n29472_));
  NAND2X1  g27036(.A(new_n29290_), .B(new_n23381_), .Y(new_n29473_));
  AOI21X1  g27037(.A0(new_n29300_), .A1(new_n22584_), .B0(pi0233), .Y(new_n29474_));
  AOI22X1  g27038(.A0(new_n29474_), .A1(new_n29473_), .B0(new_n29472_), .B1(new_n29471_), .Y(new_n29475_));
  MX2X1    g27039(.A(new_n29475_), .B(new_n29470_), .S0(pi0237), .Y(po0746));
  AND3X1   g27040(.A(new_n8959_), .B(pi0588), .C(new_n27864_), .Y(new_n29477_));
  AOI21X1  g27041(.A0(new_n8959_), .A1(new_n27864_), .B0(new_n6334_), .Y(new_n29478_));
  OR4X1    g27042(.A(new_n29478_), .B(new_n29477_), .C(new_n2759_), .D(new_n5024_), .Y(po0747));
  OAI21X1  g27043(.A0(new_n29463_), .A1(pi0592), .B0(new_n28982_), .Y(new_n29480_));
  AOI21X1  g27044(.A0(new_n29463_), .A1(new_n6069_), .B0(new_n29480_), .Y(po0748));
  OAI21X1  g27045(.A0(new_n29463_), .A1(pi0590), .B0(new_n28982_), .Y(new_n29482_));
  AOI21X1  g27046(.A0(new_n29463_), .A1(new_n6009_), .B0(new_n29482_), .Y(po0749));
  INVX1    g27047(.A(pi0517), .Y(new_n29484_));
  INVX1    g27048(.A(pi0508), .Y(new_n29485_));
  INVX1    g27049(.A(pi0509), .Y(new_n29486_));
  INVX1    g27050(.A(pi0504), .Y(new_n29487_));
  INVX1    g27051(.A(pi0537), .Y(new_n29488_));
  AOI21X1  g27052(.A0(new_n29290_), .A1(new_n2973_), .B0(pi0557), .Y(new_n29489_));
  AOI21X1  g27053(.A0(new_n29290_), .A1(pi0234), .B0(new_n29363_), .Y(new_n29490_));
  XOR2X1   g27054(.A(pi0536), .B(pi0246), .Y(new_n29491_));
  NOR4X1   g27055(.A(new_n29491_), .B(new_n29490_), .C(new_n29489_), .D(pi0538), .Y(new_n29492_));
  INVX1    g27056(.A(pi0538), .Y(new_n29493_));
  NOR4X1   g27057(.A(new_n29491_), .B(new_n29490_), .C(new_n29489_), .D(new_n29493_), .Y(new_n29494_));
  MX2X1    g27058(.A(new_n29492_), .B(new_n29494_), .S0(pi0249), .Y(new_n29495_));
  AOI21X1  g27059(.A0(new_n29495_), .A1(new_n29488_), .B0(pi0248), .Y(new_n29496_));
  AOI21X1  g27060(.A0(new_n29495_), .A1(pi0537), .B0(new_n4000_), .Y(new_n29497_));
  XOR2X1   g27061(.A(pi0506), .B(pi0241), .Y(new_n29498_));
  XOR2X1   g27062(.A(pi0535), .B(pi0240), .Y(new_n29499_));
  NOR4X1   g27063(.A(new_n29499_), .B(new_n29498_), .C(new_n29497_), .D(new_n29496_), .Y(new_n29500_));
  AOI21X1  g27064(.A0(new_n29500_), .A1(pi0534), .B0(pi0239), .Y(new_n29501_));
  AOI21X1  g27065(.A0(new_n29500_), .A1(new_n29335_), .B0(new_n3229_), .Y(new_n29502_));
  OR2X1    g27066(.A(new_n29502_), .B(new_n29501_), .Y(new_n29503_));
  OAI21X1  g27067(.A0(new_n29503_), .A1(new_n29487_), .B0(pi0242), .Y(new_n29504_));
  OAI21X1  g27068(.A0(new_n29503_), .A1(pi0504), .B0(new_n4884_), .Y(new_n29505_));
  NAND3X1  g27069(.A(new_n29505_), .B(new_n29504_), .C(pi0533), .Y(new_n29506_));
  AND2X1   g27070(.A(new_n29506_), .B(pi0235), .Y(new_n29507_));
  INVX1    g27071(.A(pi0533), .Y(new_n29508_));
  AND3X1   g27072(.A(new_n29505_), .B(new_n29504_), .C(new_n29508_), .Y(new_n29509_));
  NOR2X1   g27073(.A(new_n29509_), .B(pi0235), .Y(new_n29510_));
  NOR2X1   g27074(.A(new_n29510_), .B(new_n29507_), .Y(new_n29511_));
  AOI21X1  g27075(.A0(new_n29511_), .A1(pi0558), .B0(new_n4691_), .Y(new_n29512_));
  INVX1    g27076(.A(pi0558), .Y(new_n29513_));
  AOI21X1  g27077(.A0(new_n29511_), .A1(new_n29513_), .B0(pi0244), .Y(new_n29514_));
  OR3X1    g27078(.A(new_n29514_), .B(new_n29512_), .C(new_n29486_), .Y(new_n29515_));
  AND2X1   g27079(.A(new_n29515_), .B(pi0245), .Y(new_n29516_));
  NOR3X1   g27080(.A(new_n29514_), .B(new_n29512_), .C(pi0509), .Y(new_n29517_));
  NOR2X1   g27081(.A(new_n29517_), .B(pi0245), .Y(new_n29518_));
  OR2X1    g27082(.A(new_n29518_), .B(new_n29516_), .Y(new_n29519_));
  OAI21X1  g27083(.A0(new_n29519_), .A1(new_n29485_), .B0(pi0247), .Y(new_n29520_));
  XOR2X1   g27084(.A(pi0481), .B(pi0248), .Y(new_n29521_));
  AND2X1   g27085(.A(new_n29300_), .B(pi0234), .Y(new_n29522_));
  INVX1    g27086(.A(new_n29522_), .Y(new_n29523_));
  XOR2X1   g27087(.A(pi0487), .B(pi0246), .Y(new_n29524_));
  AOI21X1  g27088(.A0(new_n29523_), .A1(pi0511), .B0(new_n29524_), .Y(new_n29525_));
  OAI21X1  g27089(.A0(new_n29301_), .A1(pi0511), .B0(new_n29525_), .Y(new_n29526_));
  XOR2X1   g27090(.A(pi0579), .B(pi0249), .Y(new_n29527_));
  NOR3X1   g27091(.A(new_n29527_), .B(new_n29526_), .C(new_n29521_), .Y(new_n29528_));
  AOI21X1  g27092(.A0(new_n29528_), .A1(pi0559), .B0(new_n3854_), .Y(new_n29529_));
  INVX1    g27093(.A(pi0559), .Y(new_n29530_));
  AOI21X1  g27094(.A0(new_n29528_), .A1(new_n29530_), .B0(pi0241), .Y(new_n29531_));
  NOR2X1   g27095(.A(new_n29531_), .B(new_n29529_), .Y(new_n29532_));
  AOI21X1  g27096(.A0(new_n29532_), .A1(pi0515), .B0(new_n4443_), .Y(new_n29533_));
  INVX1    g27097(.A(pi0515), .Y(new_n29534_));
  INVX1    g27098(.A(new_n29497_), .Y(new_n29535_));
  NOR2X1   g27099(.A(new_n29527_), .B(new_n29526_), .Y(new_n29536_));
  OR2X1    g27100(.A(new_n29536_), .B(pi0579), .Y(new_n29537_));
  NOR2X1   g27101(.A(new_n29492_), .B(pi0249), .Y(new_n29538_));
  OAI21X1  g27102(.A0(new_n29526_), .A1(new_n29538_), .B0(pi0579), .Y(new_n29539_));
  AOI21X1  g27103(.A0(new_n29539_), .A1(new_n29537_), .B0(new_n29495_), .Y(new_n29540_));
  AOI21X1  g27104(.A0(new_n29536_), .A1(pi0537), .B0(pi0248), .Y(new_n29541_));
  OAI21X1  g27105(.A0(new_n29540_), .A1(pi0537), .B0(new_n29541_), .Y(new_n29542_));
  NAND2X1  g27106(.A(new_n29542_), .B(new_n29535_), .Y(new_n29543_));
  INVX1    g27107(.A(new_n29496_), .Y(new_n29544_));
  AOI21X1  g27108(.A0(new_n29536_), .A1(new_n29488_), .B0(new_n4000_), .Y(new_n29545_));
  OAI21X1  g27109(.A0(new_n29540_), .A1(new_n29488_), .B0(new_n29545_), .Y(new_n29546_));
  NAND2X1  g27110(.A(new_n29546_), .B(new_n29544_), .Y(new_n29547_));
  MX2X1    g27111(.A(new_n29543_), .B(new_n29547_), .S0(pi0481), .Y(new_n29548_));
  OR2X1    g27112(.A(new_n29548_), .B(pi0559), .Y(new_n29549_));
  NOR2X1   g27113(.A(new_n29497_), .B(new_n29496_), .Y(new_n29550_));
  AOI21X1  g27114(.A0(new_n29550_), .A1(pi0559), .B0(pi0241), .Y(new_n29551_));
  AOI21X1  g27115(.A0(new_n29551_), .A1(new_n29549_), .B0(new_n29529_), .Y(new_n29552_));
  OR2X1    g27116(.A(new_n29548_), .B(new_n29530_), .Y(new_n29553_));
  AOI21X1  g27117(.A0(new_n29550_), .A1(new_n29530_), .B0(new_n3854_), .Y(new_n29554_));
  AOI21X1  g27118(.A0(new_n29554_), .A1(new_n29553_), .B0(new_n29531_), .Y(new_n29555_));
  MX2X1    g27119(.A(new_n29552_), .B(new_n29555_), .S0(pi0506), .Y(new_n29556_));
  OR3X1    g27120(.A(new_n29498_), .B(new_n29497_), .C(new_n29496_), .Y(new_n29557_));
  OAI21X1  g27121(.A0(new_n29557_), .A1(new_n29534_), .B0(new_n4443_), .Y(new_n29558_));
  AOI21X1  g27122(.A0(new_n29556_), .A1(new_n29534_), .B0(new_n29558_), .Y(new_n29559_));
  NOR2X1   g27123(.A(new_n29559_), .B(new_n29533_), .Y(new_n29560_));
  AOI21X1  g27124(.A0(new_n29532_), .A1(new_n29534_), .B0(pi0240), .Y(new_n29561_));
  OAI21X1  g27125(.A0(new_n29557_), .A1(pi0515), .B0(pi0240), .Y(new_n29562_));
  AOI21X1  g27126(.A0(new_n29556_), .A1(pi0515), .B0(new_n29562_), .Y(new_n29563_));
  NOR2X1   g27127(.A(new_n29563_), .B(new_n29561_), .Y(new_n29564_));
  MX2X1    g27128(.A(new_n29560_), .B(new_n29564_), .S0(pi0535), .Y(new_n29565_));
  OR2X1    g27129(.A(new_n29561_), .B(new_n29533_), .Y(new_n29566_));
  OAI21X1  g27130(.A0(new_n29566_), .A1(new_n29335_), .B0(pi0239), .Y(new_n29567_));
  AOI21X1  g27131(.A0(new_n29565_), .A1(new_n29335_), .B0(new_n29567_), .Y(new_n29568_));
  OAI21X1  g27132(.A0(new_n29568_), .A1(new_n29501_), .B0(new_n29269_), .Y(new_n29569_));
  OAI21X1  g27133(.A0(new_n29566_), .A1(pi0534), .B0(new_n3229_), .Y(new_n29570_));
  AOI21X1  g27134(.A0(new_n29565_), .A1(pi0534), .B0(new_n29570_), .Y(new_n29571_));
  OAI21X1  g27135(.A0(new_n29571_), .A1(new_n29502_), .B0(pi0488), .Y(new_n29572_));
  NAND2X1  g27136(.A(new_n29572_), .B(new_n29569_), .Y(new_n29573_));
  XOR2X1   g27137(.A(pi0488), .B(new_n3229_), .Y(new_n29574_));
  NOR3X1   g27138(.A(new_n29574_), .B(new_n29561_), .C(new_n29533_), .Y(new_n29575_));
  AOI21X1  g27139(.A0(new_n29575_), .A1(pi0504), .B0(pi0242), .Y(new_n29576_));
  OAI21X1  g27140(.A0(new_n29573_), .A1(pi0504), .B0(new_n29576_), .Y(new_n29577_));
  NAND2X1  g27141(.A(new_n29577_), .B(new_n29504_), .Y(new_n29578_));
  AOI21X1  g27142(.A0(new_n29575_), .A1(new_n29487_), .B0(new_n4884_), .Y(new_n29579_));
  OAI21X1  g27143(.A0(new_n29573_), .A1(new_n29487_), .B0(new_n29579_), .Y(new_n29580_));
  NAND2X1  g27144(.A(new_n29580_), .B(new_n29505_), .Y(new_n29581_));
  MX2X1    g27145(.A(new_n29578_), .B(new_n29581_), .S0(pi0510), .Y(new_n29582_));
  OR2X1    g27146(.A(new_n29582_), .B(pi0533), .Y(new_n29583_));
  XOR2X1   g27147(.A(pi0510), .B(pi0242), .Y(new_n29584_));
  NOR4X1   g27148(.A(new_n29584_), .B(new_n29574_), .C(new_n29561_), .D(new_n29533_), .Y(new_n29585_));
  AOI21X1  g27149(.A0(new_n29585_), .A1(pi0533), .B0(pi0235), .Y(new_n29586_));
  AOI21X1  g27150(.A0(new_n29586_), .A1(new_n29583_), .B0(new_n29507_), .Y(new_n29587_));
  OR2X1    g27151(.A(new_n29582_), .B(new_n29508_), .Y(new_n29588_));
  AOI21X1  g27152(.A0(new_n29585_), .A1(new_n29508_), .B0(new_n3373_), .Y(new_n29589_));
  AOI21X1  g27153(.A0(new_n29589_), .A1(new_n29588_), .B0(new_n29510_), .Y(new_n29590_));
  MX2X1    g27154(.A(new_n29587_), .B(new_n29590_), .S0(pi0512), .Y(new_n29591_));
  XOR2X1   g27155(.A(pi0512), .B(new_n3373_), .Y(new_n29592_));
  NAND2X1  g27156(.A(new_n29592_), .B(new_n29585_), .Y(new_n29593_));
  OAI21X1  g27157(.A0(new_n29593_), .A1(new_n29513_), .B0(new_n4691_), .Y(new_n29594_));
  AOI21X1  g27158(.A0(new_n29591_), .A1(new_n29513_), .B0(new_n29594_), .Y(new_n29595_));
  NOR2X1   g27159(.A(new_n29595_), .B(new_n29512_), .Y(new_n29596_));
  OAI21X1  g27160(.A0(new_n29593_), .A1(pi0558), .B0(pi0244), .Y(new_n29597_));
  AOI21X1  g27161(.A0(new_n29591_), .A1(pi0558), .B0(new_n29597_), .Y(new_n29598_));
  NOR2X1   g27162(.A(new_n29598_), .B(new_n29514_), .Y(new_n29599_));
  MX2X1    g27163(.A(new_n29596_), .B(new_n29599_), .S0(pi0513), .Y(new_n29600_));
  XOR2X1   g27164(.A(pi0513), .B(new_n4691_), .Y(new_n29601_));
  NAND3X1  g27165(.A(new_n29601_), .B(new_n29592_), .C(new_n29585_), .Y(new_n29602_));
  OAI21X1  g27166(.A0(new_n29602_), .A1(new_n29486_), .B0(new_n4545_), .Y(new_n29603_));
  AOI21X1  g27167(.A0(new_n29600_), .A1(new_n29486_), .B0(new_n29603_), .Y(new_n29604_));
  OR2X1    g27168(.A(new_n29604_), .B(new_n29516_), .Y(new_n29605_));
  OAI21X1  g27169(.A0(new_n29602_), .A1(pi0509), .B0(pi0245), .Y(new_n29606_));
  AOI21X1  g27170(.A0(new_n29600_), .A1(pi0509), .B0(new_n29606_), .Y(new_n29607_));
  OR2X1    g27171(.A(new_n29607_), .B(new_n29518_), .Y(new_n29608_));
  MX2X1    g27172(.A(new_n29605_), .B(new_n29608_), .S0(pi0514), .Y(new_n29609_));
  XOR2X1   g27173(.A(pi0514), .B(pi0245), .Y(new_n29610_));
  NOR2X1   g27174(.A(new_n29610_), .B(new_n29602_), .Y(new_n29611_));
  AOI21X1  g27175(.A0(new_n29611_), .A1(pi0508), .B0(pi0247), .Y(new_n29612_));
  OAI21X1  g27176(.A0(new_n29609_), .A1(pi0508), .B0(new_n29612_), .Y(new_n29613_));
  NAND2X1  g27177(.A(new_n29613_), .B(new_n29520_), .Y(new_n29614_));
  OAI21X1  g27178(.A0(new_n29519_), .A1(pi0508), .B0(new_n4102_), .Y(new_n29615_));
  AOI21X1  g27179(.A0(new_n29611_), .A1(new_n29485_), .B0(new_n4102_), .Y(new_n29616_));
  OAI21X1  g27180(.A0(new_n29609_), .A1(new_n29485_), .B0(new_n29616_), .Y(new_n29617_));
  NAND2X1  g27181(.A(new_n29617_), .B(new_n29615_), .Y(new_n29618_));
  MX2X1    g27182(.A(new_n29614_), .B(new_n29618_), .S0(pi0516), .Y(new_n29619_));
  OAI21X1  g27183(.A0(new_n29619_), .A1(pi0238), .B0(new_n29484_), .Y(new_n29620_));
  NAND3X1  g27184(.A(new_n29615_), .B(new_n29520_), .C(new_n3551_), .Y(new_n29621_));
  XOR2X1   g27185(.A(pi0516), .B(pi0247), .Y(new_n29622_));
  OR4X1    g27186(.A(new_n29622_), .B(new_n29610_), .C(new_n29602_), .D(new_n3551_), .Y(new_n29623_));
  AND2X1   g27187(.A(new_n29623_), .B(pi0517), .Y(new_n29624_));
  AOI21X1  g27188(.A0(new_n29624_), .A1(new_n29621_), .B0(pi0507), .Y(new_n29625_));
  AND2X1   g27189(.A(new_n29625_), .B(new_n29620_), .Y(new_n29626_));
  OR2X1    g27190(.A(new_n29619_), .B(new_n3551_), .Y(new_n29627_));
  AND3X1   g27191(.A(new_n29615_), .B(new_n29520_), .C(pi0238), .Y(new_n29628_));
  NOR4X1   g27192(.A(new_n29622_), .B(new_n29610_), .C(new_n29602_), .D(pi0238), .Y(new_n29629_));
  OR2X1    g27193(.A(new_n29629_), .B(pi0517), .Y(new_n29630_));
  OAI21X1  g27194(.A0(new_n29630_), .A1(new_n29628_), .B0(pi0507), .Y(new_n29631_));
  AOI21X1  g27195(.A0(new_n29627_), .A1(pi0517), .B0(new_n29631_), .Y(new_n29632_));
  OAI21X1  g27196(.A0(new_n29632_), .A1(new_n29626_), .B0(pi0233), .Y(new_n29633_));
  INVX1    g27197(.A(pi0539), .Y(new_n29634_));
  XOR2X1   g27198(.A(pi0542), .B(new_n4443_), .Y(new_n29635_));
  AOI21X1  g27199(.A0(new_n29290_), .A1(pi0234), .B0(new_n29289_), .Y(new_n29636_));
  AOI21X1  g27200(.A0(new_n29290_), .A1(new_n2973_), .B0(pi0505), .Y(new_n29637_));
  XOR2X1   g27201(.A(pi0501), .B(pi0248), .Y(new_n29638_));
  XOR2X1   g27202(.A(pi0499), .B(pi0246), .Y(new_n29639_));
  XOR2X1   g27203(.A(pi0496), .B(pi0249), .Y(new_n29640_));
  OR3X1    g27204(.A(new_n29640_), .B(new_n29639_), .C(new_n29638_), .Y(new_n29641_));
  XOR2X1   g27205(.A(pi0500), .B(pi0241), .Y(new_n29642_));
  NOR4X1   g27206(.A(new_n29642_), .B(new_n29641_), .C(new_n29637_), .D(new_n29636_), .Y(new_n29643_));
  AND2X1   g27207(.A(new_n29643_), .B(new_n29635_), .Y(new_n29644_));
  AOI21X1  g27208(.A0(new_n29644_), .A1(pi0497), .B0(pi0239), .Y(new_n29645_));
  AOI21X1  g27209(.A0(new_n29644_), .A1(new_n29280_), .B0(new_n3229_), .Y(new_n29646_));
  OR2X1    g27210(.A(new_n29646_), .B(new_n29645_), .Y(new_n29647_));
  OAI21X1  g27211(.A0(new_n29647_), .A1(new_n29634_), .B0(pi0242), .Y(new_n29648_));
  OAI21X1  g27212(.A0(new_n29647_), .A1(pi0539), .B0(new_n4884_), .Y(new_n29649_));
  AND2X1   g27213(.A(new_n29649_), .B(new_n29648_), .Y(new_n29650_));
  AOI21X1  g27214(.A0(new_n29650_), .A1(pi0540), .B0(new_n3373_), .Y(new_n29651_));
  INVX1    g27215(.A(pi0540), .Y(new_n29652_));
  AND3X1   g27216(.A(new_n29649_), .B(new_n29648_), .C(new_n29652_), .Y(new_n29653_));
  NOR2X1   g27217(.A(new_n29653_), .B(pi0235), .Y(new_n29654_));
  XOR2X1   g27218(.A(pi0541), .B(pi0244), .Y(new_n29655_));
  XOR2X1   g27219(.A(pi0503), .B(pi0245), .Y(new_n29656_));
  OR4X1    g27220(.A(new_n29656_), .B(new_n29655_), .C(new_n29654_), .D(new_n29651_), .Y(new_n29657_));
  OAI21X1  g27221(.A0(new_n29657_), .A1(pi0502), .B0(new_n4102_), .Y(new_n29658_));
  OAI21X1  g27222(.A0(pi0561), .A1(pi0247), .B0(new_n29658_), .Y(new_n29659_));
  AOI21X1  g27223(.A0(new_n29300_), .A1(pi0234), .B0(new_n29310_), .Y(new_n29660_));
  XOR2X1   g27224(.A(pi0521), .B(pi0248), .Y(new_n29661_));
  XOR2X1   g27225(.A(pi0520), .B(pi0246), .Y(new_n29662_));
  XOR2X1   g27226(.A(pi0574), .B(pi0241), .Y(new_n29663_));
  XOR2X1   g27227(.A(pi0578), .B(pi0249), .Y(new_n29664_));
  NOR4X1   g27228(.A(new_n29664_), .B(new_n29663_), .C(new_n29662_), .D(new_n29661_), .Y(new_n29665_));
  OAI21X1  g27229(.A0(new_n29301_), .A1(pi0518), .B0(new_n29665_), .Y(new_n29666_));
  NOR2X1   g27230(.A(new_n29666_), .B(new_n29660_), .Y(new_n29667_));
  AOI21X1  g27231(.A0(new_n29667_), .A1(pi0582), .B0(new_n4443_), .Y(new_n29668_));
  INVX1    g27232(.A(pi0582), .Y(new_n29669_));
  AOI21X1  g27233(.A0(new_n29667_), .A1(new_n29669_), .B0(pi0240), .Y(new_n29670_));
  XOR2X1   g27234(.A(pi0519), .B(new_n3229_), .Y(new_n29671_));
  XOR2X1   g27235(.A(pi0586), .B(pi0242), .Y(new_n29672_));
  NOR4X1   g27236(.A(new_n29672_), .B(new_n29671_), .C(new_n29670_), .D(new_n29668_), .Y(new_n29673_));
  XOR2X1   g27237(.A(pi0581), .B(new_n3373_), .Y(new_n29674_));
  AND2X1   g27238(.A(new_n29674_), .B(new_n29673_), .Y(new_n29675_));
  AOI21X1  g27239(.A0(new_n29675_), .A1(pi0585), .B0(new_n4691_), .Y(new_n29676_));
  INVX1    g27240(.A(pi0585), .Y(new_n29677_));
  AOI21X1  g27241(.A0(new_n29675_), .A1(new_n29677_), .B0(pi0244), .Y(new_n29678_));
  NOR2X1   g27242(.A(new_n29678_), .B(new_n29676_), .Y(new_n29679_));
  AOI21X1  g27243(.A0(new_n29679_), .A1(pi0584), .B0(new_n4545_), .Y(new_n29680_));
  INVX1    g27244(.A(pi0584), .Y(new_n29681_));
  INVX1    g27245(.A(new_n29651_), .Y(new_n29682_));
  INVX1    g27246(.A(pi0500), .Y(new_n29683_));
  NAND2X1  g27247(.A(pi0500), .B(pi0241), .Y(new_n29684_));
  OR4X1    g27248(.A(new_n29684_), .B(new_n29641_), .C(new_n29637_), .D(new_n29636_), .Y(new_n29685_));
  OAI21X1  g27249(.A0(new_n29666_), .A1(new_n29660_), .B0(new_n29685_), .Y(new_n29686_));
  AOI21X1  g27250(.A0(new_n29643_), .A1(new_n29683_), .B0(new_n29686_), .Y(new_n29687_));
  OR2X1    g27251(.A(new_n29687_), .B(pi0582), .Y(new_n29688_));
  AOI21X1  g27252(.A0(new_n29643_), .A1(pi0582), .B0(pi0240), .Y(new_n29689_));
  AOI21X1  g27253(.A0(new_n29689_), .A1(new_n29688_), .B0(new_n29668_), .Y(new_n29690_));
  OR2X1    g27254(.A(new_n29687_), .B(new_n29669_), .Y(new_n29691_));
  AOI21X1  g27255(.A0(new_n29643_), .A1(new_n29669_), .B0(new_n4443_), .Y(new_n29692_));
  AOI21X1  g27256(.A0(new_n29692_), .A1(new_n29691_), .B0(new_n29670_), .Y(new_n29693_));
  MX2X1    g27257(.A(new_n29690_), .B(new_n29693_), .S0(pi0542), .Y(new_n29694_));
  OR2X1    g27258(.A(new_n29670_), .B(new_n29668_), .Y(new_n29695_));
  OAI21X1  g27259(.A0(new_n29695_), .A1(new_n29280_), .B0(pi0239), .Y(new_n29696_));
  AOI21X1  g27260(.A0(new_n29694_), .A1(new_n29280_), .B0(new_n29696_), .Y(new_n29697_));
  OAI21X1  g27261(.A0(new_n29697_), .A1(new_n29645_), .B0(new_n29315_), .Y(new_n29698_));
  OAI21X1  g27262(.A0(new_n29695_), .A1(pi0497), .B0(new_n3229_), .Y(new_n29699_));
  AOI21X1  g27263(.A0(new_n29694_), .A1(pi0497), .B0(new_n29699_), .Y(new_n29700_));
  OAI21X1  g27264(.A0(new_n29700_), .A1(new_n29646_), .B0(pi0519), .Y(new_n29701_));
  AND3X1   g27265(.A(new_n29701_), .B(new_n29698_), .C(new_n29634_), .Y(new_n29702_));
  OR3X1    g27266(.A(new_n29671_), .B(new_n29670_), .C(new_n29668_), .Y(new_n29703_));
  OAI21X1  g27267(.A0(new_n29703_), .A1(new_n29634_), .B0(new_n4884_), .Y(new_n29704_));
  OAI21X1  g27268(.A0(new_n29704_), .A1(new_n29702_), .B0(new_n29648_), .Y(new_n29705_));
  AND3X1   g27269(.A(new_n29701_), .B(new_n29698_), .C(pi0539), .Y(new_n29706_));
  OAI21X1  g27270(.A0(new_n29703_), .A1(pi0539), .B0(pi0242), .Y(new_n29707_));
  OAI21X1  g27271(.A0(new_n29707_), .A1(new_n29706_), .B0(new_n29649_), .Y(new_n29708_));
  MX2X1    g27272(.A(new_n29705_), .B(new_n29708_), .S0(pi0586), .Y(new_n29709_));
  AOI21X1  g27273(.A0(new_n29673_), .A1(pi0540), .B0(pi0235), .Y(new_n29710_));
  OAI21X1  g27274(.A0(new_n29709_), .A1(pi0540), .B0(new_n29710_), .Y(new_n29711_));
  NAND2X1  g27275(.A(new_n29711_), .B(new_n29682_), .Y(new_n29712_));
  AOI21X1  g27276(.A0(new_n29673_), .A1(new_n29652_), .B0(new_n3373_), .Y(new_n29713_));
  OAI21X1  g27277(.A0(new_n29709_), .A1(new_n29652_), .B0(new_n29713_), .Y(new_n29714_));
  OAI21X1  g27278(.A0(new_n29653_), .A1(pi0235), .B0(new_n29714_), .Y(new_n29715_));
  MX2X1    g27279(.A(new_n29712_), .B(new_n29715_), .S0(pi0581), .Y(new_n29716_));
  OR2X1    g27280(.A(new_n29716_), .B(pi0585), .Y(new_n29717_));
  NOR2X1   g27281(.A(new_n29654_), .B(new_n29651_), .Y(new_n29718_));
  AOI21X1  g27282(.A0(new_n29718_), .A1(pi0585), .B0(pi0244), .Y(new_n29719_));
  AOI21X1  g27283(.A0(new_n29719_), .A1(new_n29717_), .B0(new_n29676_), .Y(new_n29720_));
  OR2X1    g27284(.A(new_n29716_), .B(new_n29677_), .Y(new_n29721_));
  AOI21X1  g27285(.A0(new_n29718_), .A1(new_n29677_), .B0(new_n4691_), .Y(new_n29722_));
  AOI21X1  g27286(.A0(new_n29722_), .A1(new_n29721_), .B0(new_n29678_), .Y(new_n29723_));
  MX2X1    g27287(.A(new_n29720_), .B(new_n29723_), .S0(pi0541), .Y(new_n29724_));
  OR3X1    g27288(.A(new_n29655_), .B(new_n29654_), .C(new_n29651_), .Y(new_n29725_));
  OAI21X1  g27289(.A0(new_n29725_), .A1(new_n29681_), .B0(new_n4545_), .Y(new_n29726_));
  AOI21X1  g27290(.A0(new_n29724_), .A1(new_n29681_), .B0(new_n29726_), .Y(new_n29727_));
  NOR2X1   g27291(.A(new_n29727_), .B(new_n29680_), .Y(new_n29728_));
  AOI21X1  g27292(.A0(new_n29679_), .A1(new_n29681_), .B0(pi0245), .Y(new_n29729_));
  OAI21X1  g27293(.A0(new_n29725_), .A1(pi0584), .B0(pi0245), .Y(new_n29730_));
  AOI21X1  g27294(.A0(new_n29724_), .A1(pi0584), .B0(new_n29730_), .Y(new_n29731_));
  NOR2X1   g27295(.A(new_n29731_), .B(new_n29729_), .Y(new_n29732_));
  MX2X1    g27296(.A(new_n29728_), .B(new_n29732_), .S0(pi0503), .Y(new_n29733_));
  OR2X1    g27297(.A(new_n29729_), .B(new_n29680_), .Y(new_n29734_));
  AOI21X1  g27298(.A0(new_n29734_), .A1(pi0502), .B0(pi0561), .Y(new_n29735_));
  OAI21X1  g27299(.A0(new_n29733_), .A1(pi0502), .B0(new_n29735_), .Y(new_n29736_));
  INVX1    g27300(.A(pi0561), .Y(new_n29737_));
  INVX1    g27301(.A(pi0502), .Y(new_n29738_));
  OAI21X1  g27302(.A0(new_n29657_), .A1(new_n29738_), .B0(pi0247), .Y(new_n29739_));
  OAI21X1  g27303(.A0(new_n29737_), .A1(new_n4102_), .B0(new_n29739_), .Y(new_n29740_));
  AOI21X1  g27304(.A0(new_n29734_), .A1(new_n29738_), .B0(new_n29737_), .Y(new_n29741_));
  OAI21X1  g27305(.A0(new_n29733_), .A1(new_n29738_), .B0(new_n29741_), .Y(new_n29742_));
  AOI22X1  g27306(.A0(new_n29742_), .A1(new_n29740_), .B0(new_n29736_), .B1(new_n29659_), .Y(new_n29743_));
  AOI21X1  g27307(.A0(new_n29743_), .A1(new_n3551_), .B0(pi0522), .Y(new_n29744_));
  INVX1    g27308(.A(pi0543), .Y(new_n29745_));
  AND3X1   g27309(.A(new_n29739_), .B(new_n29658_), .C(new_n3551_), .Y(new_n29746_));
  XOR2X1   g27310(.A(pi0561), .B(pi0247), .Y(new_n29747_));
  OR3X1    g27311(.A(new_n29747_), .B(new_n29729_), .C(new_n29680_), .Y(new_n29748_));
  OAI21X1  g27312(.A0(new_n29748_), .A1(new_n3551_), .B0(pi0522), .Y(new_n29749_));
  OAI21X1  g27313(.A0(new_n29749_), .A1(new_n29746_), .B0(new_n29745_), .Y(new_n29750_));
  INVX1    g27314(.A(pi0522), .Y(new_n29751_));
  AOI21X1  g27315(.A0(new_n29743_), .A1(pi0238), .B0(new_n29751_), .Y(new_n29752_));
  AND3X1   g27316(.A(new_n29739_), .B(new_n29658_), .C(pi0238), .Y(new_n29753_));
  OAI21X1  g27317(.A0(new_n29748_), .A1(pi0238), .B0(new_n29751_), .Y(new_n29754_));
  OAI21X1  g27318(.A0(new_n29754_), .A1(new_n29753_), .B0(pi0543), .Y(new_n29755_));
  OAI22X1  g27319(.A0(new_n29755_), .A1(new_n29752_), .B0(new_n29750_), .B1(new_n29744_), .Y(new_n29756_));
  AOI21X1  g27320(.A0(new_n29756_), .A1(new_n22655_), .B0(new_n22579_), .Y(new_n29757_));
  INVX1    g27321(.A(pi0491), .Y(new_n29758_));
  INVX1    g27322(.A(pi0529), .Y(new_n29759_));
  INVX1    g27323(.A(pi0547), .Y(new_n29760_));
  INVX1    g27324(.A(pi0483), .Y(new_n29761_));
  XOR2X1   g27325(.A(pi0492), .B(new_n4443_), .Y(new_n29762_));
  XOR2X1   g27326(.A(pi0490), .B(pi0241), .Y(new_n29763_));
  AOI21X1  g27327(.A0(new_n29290_), .A1(new_n2973_), .B0(pi0544), .Y(new_n29764_));
  AOI21X1  g27328(.A0(new_n29290_), .A1(pi0234), .B0(new_n29346_), .Y(new_n29765_));
  XOR2X1   g27329(.A(pi0484), .B(pi0249), .Y(new_n29766_));
  XOR2X1   g27330(.A(pi0546), .B(pi0246), .Y(new_n29767_));
  XOR2X1   g27331(.A(pi0548), .B(pi0248), .Y(new_n29768_));
  OR3X1    g27332(.A(new_n29768_), .B(new_n29767_), .C(new_n29766_), .Y(new_n29769_));
  NOR4X1   g27333(.A(new_n29769_), .B(new_n29765_), .C(new_n29764_), .D(new_n29763_), .Y(new_n29770_));
  AND2X1   g27334(.A(new_n29770_), .B(new_n29762_), .Y(new_n29771_));
  AOI21X1  g27335(.A0(new_n29771_), .A1(pi0494), .B0(pi0239), .Y(new_n29772_));
  AOI21X1  g27336(.A0(new_n29771_), .A1(new_n29276_), .B0(new_n3229_), .Y(new_n29773_));
  OR2X1    g27337(.A(new_n29773_), .B(new_n29772_), .Y(new_n29774_));
  OAI21X1  g27338(.A0(new_n29774_), .A1(new_n29761_), .B0(pi0242), .Y(new_n29775_));
  OAI21X1  g27339(.A0(new_n29774_), .A1(pi0483), .B0(new_n4884_), .Y(new_n29776_));
  AND2X1   g27340(.A(new_n29776_), .B(new_n29775_), .Y(new_n29777_));
  AOI21X1  g27341(.A0(new_n29777_), .A1(pi0495), .B0(new_n3373_), .Y(new_n29778_));
  INVX1    g27342(.A(pi0495), .Y(new_n29779_));
  AND3X1   g27343(.A(new_n29776_), .B(new_n29775_), .C(new_n29779_), .Y(new_n29780_));
  NOR2X1   g27344(.A(new_n29780_), .B(pi0235), .Y(new_n29781_));
  XOR2X1   g27345(.A(pi0493), .B(pi0244), .Y(new_n29782_));
  NOR3X1   g27346(.A(new_n29782_), .B(new_n29781_), .C(new_n29778_), .Y(new_n29783_));
  AOI21X1  g27347(.A0(new_n29783_), .A1(pi0545), .B0(new_n4545_), .Y(new_n29784_));
  INVX1    g27348(.A(pi0545), .Y(new_n29785_));
  AOI21X1  g27349(.A0(new_n29783_), .A1(new_n29785_), .B0(pi0245), .Y(new_n29786_));
  OR3X1    g27350(.A(new_n29786_), .B(new_n29784_), .C(new_n29760_), .Y(new_n29787_));
  AND2X1   g27351(.A(new_n29787_), .B(pi0247), .Y(new_n29788_));
  INVX1    g27352(.A(pi0571), .Y(new_n29789_));
  AOI21X1  g27353(.A0(new_n29300_), .A1(pi0234), .B0(new_n29320_), .Y(new_n29790_));
  AOI21X1  g27354(.A0(new_n29300_), .A1(new_n2973_), .B0(pi0523), .Y(new_n29791_));
  XOR2X1   g27355(.A(pi0528), .B(pi0249), .Y(new_n29792_));
  XOR2X1   g27356(.A(pi0526), .B(pi0246), .Y(new_n29793_));
  XOR2X1   g27357(.A(pi0576), .B(pi0248), .Y(new_n29794_));
  OR3X1    g27358(.A(new_n29794_), .B(new_n29793_), .C(new_n29792_), .Y(new_n29795_));
  OR4X1    g27359(.A(new_n29795_), .B(new_n29791_), .C(new_n29790_), .D(new_n29789_), .Y(new_n29796_));
  OR4X1    g27360(.A(new_n29795_), .B(new_n29791_), .C(new_n29790_), .D(pi0571), .Y(new_n29797_));
  MX2X1    g27361(.A(new_n29797_), .B(new_n29796_), .S0(pi0241), .Y(new_n29798_));
  NOR2X1   g27362(.A(new_n29798_), .B(pi0530), .Y(new_n29799_));
  NOR2X1   g27363(.A(new_n29799_), .B(pi0240), .Y(new_n29800_));
  INVX1    g27364(.A(pi0530), .Y(new_n29801_));
  NOR2X1   g27365(.A(new_n29798_), .B(new_n29801_), .Y(new_n29802_));
  NOR2X1   g27366(.A(new_n29802_), .B(new_n4443_), .Y(new_n29803_));
  XOR2X1   g27367(.A(pi0524), .B(new_n3229_), .Y(new_n29804_));
  XOR2X1   g27368(.A(pi0573), .B(pi0242), .Y(new_n29805_));
  NOR4X1   g27369(.A(new_n29805_), .B(new_n29804_), .C(new_n29803_), .D(new_n29800_), .Y(new_n29806_));
  XOR2X1   g27370(.A(pi0575), .B(new_n3373_), .Y(new_n29807_));
  AND2X1   g27371(.A(new_n29807_), .B(new_n29806_), .Y(new_n29808_));
  AOI21X1  g27372(.A0(new_n29808_), .A1(pi0572), .B0(new_n4691_), .Y(new_n29809_));
  INVX1    g27373(.A(new_n29778_), .Y(new_n29810_));
  AOI21X1  g27374(.A0(new_n29799_), .A1(pi0492), .B0(pi0240), .Y(new_n29811_));
  OR3X1    g27375(.A(new_n29769_), .B(new_n29765_), .C(new_n29764_), .Y(new_n29812_));
  AND2X1   g27376(.A(new_n29812_), .B(new_n3854_), .Y(new_n29813_));
  AOI22X1  g27377(.A0(new_n29813_), .A1(new_n29797_), .B0(new_n29796_), .B1(pi0241), .Y(new_n29814_));
  AND2X1   g27378(.A(new_n29812_), .B(pi0241), .Y(new_n29815_));
  AOI22X1  g27379(.A0(new_n29815_), .A1(new_n29796_), .B0(new_n29797_), .B1(new_n3854_), .Y(new_n29816_));
  MX2X1    g27380(.A(new_n29814_), .B(new_n29816_), .S0(pi0490), .Y(new_n29817_));
  INVX1    g27381(.A(new_n29770_), .Y(new_n29818_));
  AOI21X1  g27382(.A0(new_n29818_), .A1(pi0530), .B0(pi0492), .Y(new_n29819_));
  OAI21X1  g27383(.A0(new_n29817_), .A1(pi0530), .B0(new_n29819_), .Y(new_n29820_));
  INVX1    g27384(.A(pi0492), .Y(new_n29821_));
  AOI21X1  g27385(.A0(new_n29802_), .A1(new_n29821_), .B0(new_n4443_), .Y(new_n29822_));
  AOI21X1  g27386(.A0(new_n29818_), .A1(new_n29801_), .B0(new_n29821_), .Y(new_n29823_));
  OAI21X1  g27387(.A0(new_n29817_), .A1(new_n29801_), .B0(new_n29823_), .Y(new_n29824_));
  AOI22X1  g27388(.A0(new_n29824_), .A1(new_n29822_), .B0(new_n29820_), .B1(new_n29811_), .Y(new_n29825_));
  OR2X1    g27389(.A(new_n29803_), .B(new_n29800_), .Y(new_n29826_));
  OAI21X1  g27390(.A0(new_n29826_), .A1(new_n29276_), .B0(pi0239), .Y(new_n29827_));
  AOI21X1  g27391(.A0(new_n29825_), .A1(new_n29276_), .B0(new_n29827_), .Y(new_n29828_));
  OAI21X1  g27392(.A0(new_n29828_), .A1(new_n29772_), .B0(new_n29324_), .Y(new_n29829_));
  OAI21X1  g27393(.A0(new_n29826_), .A1(pi0494), .B0(new_n3229_), .Y(new_n29830_));
  AOI21X1  g27394(.A0(new_n29825_), .A1(pi0494), .B0(new_n29830_), .Y(new_n29831_));
  OAI21X1  g27395(.A0(new_n29831_), .A1(new_n29773_), .B0(pi0524), .Y(new_n29832_));
  AND3X1   g27396(.A(new_n29832_), .B(new_n29829_), .C(new_n29761_), .Y(new_n29833_));
  OR3X1    g27397(.A(new_n29804_), .B(new_n29803_), .C(new_n29800_), .Y(new_n29834_));
  OAI21X1  g27398(.A0(new_n29834_), .A1(new_n29761_), .B0(new_n4884_), .Y(new_n29835_));
  OAI21X1  g27399(.A0(new_n29835_), .A1(new_n29833_), .B0(new_n29775_), .Y(new_n29836_));
  AND3X1   g27400(.A(new_n29832_), .B(new_n29829_), .C(pi0483), .Y(new_n29837_));
  OAI21X1  g27401(.A0(new_n29834_), .A1(pi0483), .B0(pi0242), .Y(new_n29838_));
  OAI21X1  g27402(.A0(new_n29838_), .A1(new_n29837_), .B0(new_n29776_), .Y(new_n29839_));
  MX2X1    g27403(.A(new_n29836_), .B(new_n29839_), .S0(pi0573), .Y(new_n29840_));
  AOI21X1  g27404(.A0(new_n29806_), .A1(pi0495), .B0(pi0235), .Y(new_n29841_));
  OAI21X1  g27405(.A0(new_n29840_), .A1(pi0495), .B0(new_n29841_), .Y(new_n29842_));
  NAND2X1  g27406(.A(new_n29842_), .B(new_n29810_), .Y(new_n29843_));
  AOI21X1  g27407(.A0(new_n29806_), .A1(new_n29779_), .B0(new_n3373_), .Y(new_n29844_));
  OAI21X1  g27408(.A0(new_n29840_), .A1(new_n29779_), .B0(new_n29844_), .Y(new_n29845_));
  OAI21X1  g27409(.A0(new_n29780_), .A1(pi0235), .B0(new_n29845_), .Y(new_n29846_));
  MX2X1    g27410(.A(new_n29843_), .B(new_n29846_), .S0(pi0575), .Y(new_n29847_));
  OR2X1    g27411(.A(new_n29847_), .B(pi0572), .Y(new_n29848_));
  NOR2X1   g27412(.A(new_n29781_), .B(new_n29778_), .Y(new_n29849_));
  AOI21X1  g27413(.A0(new_n29849_), .A1(pi0572), .B0(pi0244), .Y(new_n29850_));
  AOI21X1  g27414(.A0(new_n29850_), .A1(new_n29848_), .B0(new_n29809_), .Y(new_n29851_));
  INVX1    g27415(.A(pi0572), .Y(new_n29852_));
  AOI21X1  g27416(.A0(new_n29808_), .A1(new_n29852_), .B0(pi0244), .Y(new_n29853_));
  OR2X1    g27417(.A(new_n29847_), .B(new_n29852_), .Y(new_n29854_));
  AOI21X1  g27418(.A0(new_n29849_), .A1(new_n29852_), .B0(new_n4691_), .Y(new_n29855_));
  AOI21X1  g27419(.A0(new_n29855_), .A1(new_n29854_), .B0(new_n29853_), .Y(new_n29856_));
  MX2X1    g27420(.A(new_n29851_), .B(new_n29856_), .S0(pi0493), .Y(new_n29857_));
  OR2X1    g27421(.A(new_n29853_), .B(new_n29809_), .Y(new_n29858_));
  OAI21X1  g27422(.A0(new_n29858_), .A1(new_n29785_), .B0(new_n4545_), .Y(new_n29859_));
  AOI21X1  g27423(.A0(new_n29857_), .A1(new_n29785_), .B0(new_n29859_), .Y(new_n29860_));
  NOR2X1   g27424(.A(new_n29860_), .B(new_n29784_), .Y(new_n29861_));
  OAI21X1  g27425(.A0(new_n29858_), .A1(pi0545), .B0(pi0245), .Y(new_n29862_));
  AOI21X1  g27426(.A0(new_n29857_), .A1(pi0545), .B0(new_n29862_), .Y(new_n29863_));
  NOR2X1   g27427(.A(new_n29863_), .B(new_n29786_), .Y(new_n29864_));
  MX2X1    g27428(.A(new_n29861_), .B(new_n29864_), .S0(pi0525), .Y(new_n29865_));
  XOR2X1   g27429(.A(pi0525), .B(pi0245), .Y(new_n29866_));
  OR3X1    g27430(.A(new_n29866_), .B(new_n29853_), .C(new_n29809_), .Y(new_n29867_));
  OAI21X1  g27431(.A0(new_n29867_), .A1(new_n29760_), .B0(new_n4102_), .Y(new_n29868_));
  AOI21X1  g27432(.A0(new_n29865_), .A1(new_n29760_), .B0(new_n29868_), .Y(new_n29869_));
  OR2X1    g27433(.A(new_n29869_), .B(new_n29788_), .Y(new_n29870_));
  NOR3X1   g27434(.A(new_n29786_), .B(new_n29784_), .C(pi0547), .Y(new_n29871_));
  NOR2X1   g27435(.A(new_n29871_), .B(pi0247), .Y(new_n29872_));
  OAI21X1  g27436(.A0(new_n29867_), .A1(pi0547), .B0(pi0247), .Y(new_n29873_));
  AOI21X1  g27437(.A0(new_n29865_), .A1(pi0547), .B0(new_n29873_), .Y(new_n29874_));
  OR2X1    g27438(.A(new_n29874_), .B(new_n29872_), .Y(new_n29875_));
  MX2X1    g27439(.A(new_n29870_), .B(new_n29875_), .S0(pi0527), .Y(new_n29876_));
  OAI21X1  g27440(.A0(new_n29876_), .A1(pi0238), .B0(new_n29759_), .Y(new_n29877_));
  OR2X1    g27441(.A(new_n29872_), .B(new_n29788_), .Y(new_n29878_));
  XOR2X1   g27442(.A(pi0527), .B(pi0247), .Y(new_n29879_));
  NOR4X1   g27443(.A(new_n29879_), .B(new_n29866_), .C(new_n29853_), .D(new_n29809_), .Y(new_n29880_));
  AOI21X1  g27444(.A0(new_n29880_), .A1(pi0238), .B0(new_n29759_), .Y(new_n29881_));
  OAI21X1  g27445(.A0(new_n29878_), .A1(pi0238), .B0(new_n29881_), .Y(new_n29882_));
  AND3X1   g27446(.A(new_n29882_), .B(new_n29877_), .C(new_n29758_), .Y(new_n29883_));
  OAI21X1  g27447(.A0(new_n29876_), .A1(new_n3551_), .B0(pi0529), .Y(new_n29884_));
  AOI21X1  g27448(.A0(new_n29880_), .A1(new_n3551_), .B0(pi0529), .Y(new_n29885_));
  OAI21X1  g27449(.A0(new_n29878_), .A1(new_n3551_), .B0(new_n29885_), .Y(new_n29886_));
  AND3X1   g27450(.A(new_n29886_), .B(new_n29884_), .C(pi0491), .Y(new_n29887_));
  OAI21X1  g27451(.A0(new_n29887_), .A1(new_n29883_), .B0(pi0233), .Y(new_n29888_));
  INVX1    g27452(.A(pi0486), .Y(new_n29889_));
  INVX1    g27453(.A(pi0549), .Y(new_n29890_));
  INVX1    g27454(.A(pi0489), .Y(new_n29891_));
  INVX1    g27455(.A(pi0485), .Y(new_n29892_));
  AOI21X1  g27456(.A0(new_n29290_), .A1(pi0234), .B0(new_n29892_), .Y(new_n29893_));
  AOI21X1  g27457(.A0(new_n29290_), .A1(new_n2973_), .B0(pi0485), .Y(new_n29894_));
  XOR2X1   g27458(.A(pi0555), .B(pi0249), .Y(new_n29895_));
  XOR2X1   g27459(.A(pi0553), .B(pi0241), .Y(new_n29896_));
  XOR2X1   g27460(.A(pi0551), .B(pi0240), .Y(new_n29897_));
  XOR2X1   g27461(.A(pi0554), .B(pi0248), .Y(new_n29898_));
  XOR2X1   g27462(.A(pi0563), .B(pi0246), .Y(new_n29899_));
  OR3X1    g27463(.A(new_n29899_), .B(new_n29898_), .C(new_n29897_), .Y(new_n29900_));
  OR3X1    g27464(.A(new_n29900_), .B(new_n29896_), .C(new_n29895_), .Y(new_n29901_));
  NOR4X1   g27465(.A(new_n29901_), .B(new_n29894_), .C(new_n29893_), .D(new_n29355_), .Y(new_n29902_));
  NOR4X1   g27466(.A(new_n29901_), .B(new_n29894_), .C(new_n29893_), .D(pi0550), .Y(new_n29903_));
  MX2X1    g27467(.A(new_n29903_), .B(new_n29902_), .S0(new_n3229_), .Y(new_n29904_));
  AOI21X1  g27468(.A0(new_n29904_), .A1(new_n29891_), .B0(pi0242), .Y(new_n29905_));
  AOI21X1  g27469(.A0(new_n29904_), .A1(pi0489), .B0(new_n4884_), .Y(new_n29906_));
  OR2X1    g27470(.A(new_n29906_), .B(new_n29905_), .Y(new_n29907_));
  OAI21X1  g27471(.A0(new_n29907_), .A1(new_n29890_), .B0(pi0235), .Y(new_n29908_));
  OAI21X1  g27472(.A0(new_n29907_), .A1(pi0549), .B0(new_n3373_), .Y(new_n29909_));
  NAND2X1  g27473(.A(new_n29909_), .B(new_n29908_), .Y(new_n29910_));
  OAI21X1  g27474(.A0(new_n29910_), .A1(new_n29889_), .B0(pi0244), .Y(new_n29911_));
  OAI21X1  g27475(.A0(new_n29910_), .A1(pi0486), .B0(new_n4691_), .Y(new_n29912_));
  XOR2X1   g27476(.A(pi0580), .B(new_n4545_), .Y(new_n29913_));
  NAND4X1  g27477(.A(new_n29913_), .B(new_n29912_), .C(new_n29911_), .D(pi0552), .Y(new_n29914_));
  AND2X1   g27478(.A(new_n29914_), .B(pi0247), .Y(new_n29915_));
  INVX1    g27479(.A(pi0552), .Y(new_n29916_));
  NOR2X1   g27480(.A(pi0556), .B(pi0242), .Y(new_n29917_));
  AND2X1   g27481(.A(pi0556), .B(pi0242), .Y(new_n29918_));
  AOI21X1  g27482(.A0(new_n29300_), .A1(new_n2973_), .B0(pi0570), .Y(new_n29919_));
  XOR2X1   g27483(.A(pi0562), .B(pi0241), .Y(new_n29920_));
  INVX1    g27484(.A(pi0482), .Y(new_n29921_));
  AND2X1   g27485(.A(new_n29921_), .B(pi0249), .Y(new_n29922_));
  INVX1    g27486(.A(pi0564), .Y(new_n29923_));
  OAI22X1  g27487(.A0(new_n29923_), .A1(pi0246), .B0(new_n29921_), .B1(pi0249), .Y(new_n29924_));
  NOR4X1   g27488(.A(new_n29924_), .B(new_n29922_), .C(new_n29920_), .D(new_n29919_), .Y(new_n29925_));
  OAI21X1  g27489(.A0(new_n29522_), .A1(new_n29441_), .B0(new_n29925_), .Y(new_n29926_));
  XOR2X1   g27490(.A(pi0565), .B(pi0248), .Y(new_n29927_));
  XOR2X1   g27491(.A(pi0560), .B(pi0240), .Y(new_n29928_));
  AND2X1   g27492(.A(new_n29923_), .B(pi0246), .Y(new_n29929_));
  NOR4X1   g27493(.A(new_n29929_), .B(new_n29928_), .C(new_n29927_), .D(new_n29926_), .Y(new_n29930_));
  INVX1    g27494(.A(pi0560), .Y(new_n29931_));
  NOR4X1   g27495(.A(new_n29929_), .B(new_n29927_), .C(new_n29926_), .D(new_n29931_), .Y(new_n29932_));
  MX2X1    g27496(.A(new_n29932_), .B(new_n29930_), .S0(new_n4443_), .Y(new_n29933_));
  XOR2X1   g27497(.A(pi0569), .B(pi0239), .Y(new_n29934_));
  AND2X1   g27498(.A(new_n29934_), .B(new_n29933_), .Y(new_n29935_));
  OAI21X1  g27499(.A0(new_n29918_), .A1(new_n29917_), .B0(new_n29935_), .Y(new_n29936_));
  XOR2X1   g27500(.A(pi0531), .B(pi0235), .Y(new_n29937_));
  XOR2X1   g27501(.A(pi0566), .B(pi0244), .Y(new_n29938_));
  NOR3X1   g27502(.A(new_n29938_), .B(new_n29937_), .C(new_n29936_), .Y(new_n29939_));
  AOI21X1  g27503(.A0(new_n29939_), .A1(pi0568), .B0(new_n4545_), .Y(new_n29940_));
  OR4X1    g27504(.A(new_n29901_), .B(new_n29894_), .C(new_n29893_), .D(pi0550), .Y(new_n29941_));
  AOI21X1  g27505(.A0(new_n29941_), .A1(pi0239), .B0(new_n29439_), .Y(new_n29942_));
  AND3X1   g27506(.A(new_n29930_), .B(new_n29439_), .C(pi0239), .Y(new_n29943_));
  OR2X1    g27507(.A(new_n29943_), .B(new_n29904_), .Y(new_n29944_));
  AOI21X1  g27508(.A0(new_n29942_), .A1(new_n29933_), .B0(new_n29944_), .Y(new_n29945_));
  AND2X1   g27509(.A(new_n29945_), .B(new_n29891_), .Y(new_n29946_));
  AOI21X1  g27510(.A0(new_n29934_), .A1(new_n29933_), .B0(new_n29891_), .Y(new_n29947_));
  OR2X1    g27511(.A(new_n29947_), .B(pi0556), .Y(new_n29948_));
  OAI22X1  g27512(.A0(new_n29948_), .A1(new_n29946_), .B0(new_n29917_), .B1(new_n29905_), .Y(new_n29949_));
  AND2X1   g27513(.A(new_n29945_), .B(pi0489), .Y(new_n29950_));
  OAI21X1  g27514(.A0(new_n29935_), .A1(pi0489), .B0(pi0556), .Y(new_n29951_));
  OAI22X1  g27515(.A0(new_n29951_), .A1(new_n29950_), .B0(new_n29918_), .B1(new_n29906_), .Y(new_n29952_));
  AND3X1   g27516(.A(new_n29952_), .B(new_n29949_), .C(new_n29890_), .Y(new_n29953_));
  OAI21X1  g27517(.A0(new_n29936_), .A1(new_n29890_), .B0(new_n3373_), .Y(new_n29954_));
  OAI21X1  g27518(.A0(new_n29954_), .A1(new_n29953_), .B0(new_n29908_), .Y(new_n29955_));
  AND3X1   g27519(.A(new_n29952_), .B(new_n29949_), .C(pi0549), .Y(new_n29956_));
  OAI21X1  g27520(.A0(new_n29936_), .A1(pi0549), .B0(pi0235), .Y(new_n29957_));
  OAI21X1  g27521(.A0(new_n29957_), .A1(new_n29956_), .B0(new_n29909_), .Y(new_n29958_));
  MX2X1    g27522(.A(new_n29955_), .B(new_n29958_), .S0(pi0531), .Y(new_n29959_));
  NOR2X1   g27523(.A(new_n29937_), .B(new_n29936_), .Y(new_n29960_));
  AOI21X1  g27524(.A0(new_n29960_), .A1(pi0486), .B0(pi0244), .Y(new_n29961_));
  OAI21X1  g27525(.A0(new_n29959_), .A1(pi0486), .B0(new_n29961_), .Y(new_n29962_));
  NAND2X1  g27526(.A(new_n29962_), .B(new_n29911_), .Y(new_n29963_));
  AOI21X1  g27527(.A0(new_n29960_), .A1(new_n29889_), .B0(new_n4691_), .Y(new_n29964_));
  OAI21X1  g27528(.A0(new_n29959_), .A1(new_n29889_), .B0(new_n29964_), .Y(new_n29965_));
  NAND2X1  g27529(.A(new_n29965_), .B(new_n29912_), .Y(new_n29966_));
  MX2X1    g27530(.A(new_n29963_), .B(new_n29966_), .S0(pi0566), .Y(new_n29967_));
  OR2X1    g27531(.A(new_n29967_), .B(pi0568), .Y(new_n29968_));
  AND2X1   g27532(.A(new_n29912_), .B(new_n29911_), .Y(new_n29969_));
  AOI21X1  g27533(.A0(new_n29969_), .A1(pi0568), .B0(pi0245), .Y(new_n29970_));
  AOI21X1  g27534(.A0(new_n29970_), .A1(new_n29968_), .B0(new_n29940_), .Y(new_n29971_));
  INVX1    g27535(.A(pi0568), .Y(new_n29972_));
  AOI21X1  g27536(.A0(new_n29939_), .A1(new_n29972_), .B0(pi0245), .Y(new_n29973_));
  OR2X1    g27537(.A(new_n29967_), .B(new_n29972_), .Y(new_n29974_));
  AOI21X1  g27538(.A0(new_n29969_), .A1(new_n29972_), .B0(new_n4545_), .Y(new_n29975_));
  AOI21X1  g27539(.A0(new_n29975_), .A1(new_n29974_), .B0(new_n29973_), .Y(new_n29976_));
  MX2X1    g27540(.A(new_n29971_), .B(new_n29976_), .S0(pi0580), .Y(new_n29977_));
  OR2X1    g27541(.A(new_n29973_), .B(new_n29940_), .Y(new_n29978_));
  OAI21X1  g27542(.A0(new_n29978_), .A1(new_n29916_), .B0(new_n4102_), .Y(new_n29979_));
  AOI21X1  g27543(.A0(new_n29977_), .A1(new_n29916_), .B0(new_n29979_), .Y(new_n29980_));
  NOR2X1   g27544(.A(new_n29980_), .B(new_n29915_), .Y(new_n29981_));
  NAND4X1  g27545(.A(new_n29913_), .B(new_n29912_), .C(new_n29911_), .D(new_n29916_), .Y(new_n29982_));
  AND2X1   g27546(.A(new_n29982_), .B(new_n4102_), .Y(new_n29983_));
  OAI21X1  g27547(.A0(new_n29978_), .A1(pi0552), .B0(pi0247), .Y(new_n29984_));
  AOI21X1  g27548(.A0(new_n29977_), .A1(pi0552), .B0(new_n29984_), .Y(new_n29985_));
  NOR2X1   g27549(.A(new_n29985_), .B(new_n29983_), .Y(new_n29986_));
  MX2X1    g27550(.A(new_n29981_), .B(new_n29986_), .S0(pi0532), .Y(new_n29987_));
  AOI21X1  g27551(.A0(new_n29987_), .A1(new_n3551_), .B0(pi0577), .Y(new_n29988_));
  INVX1    g27552(.A(pi0498), .Y(new_n29989_));
  NOR3X1   g27553(.A(new_n29983_), .B(new_n29915_), .C(new_n3551_), .Y(new_n29990_));
  XOR2X1   g27554(.A(pi0532), .B(pi0247), .Y(new_n29991_));
  OR3X1    g27555(.A(new_n29991_), .B(new_n29973_), .C(new_n29940_), .Y(new_n29992_));
  OAI21X1  g27556(.A0(new_n29992_), .A1(pi0238), .B0(pi0577), .Y(new_n29993_));
  OAI21X1  g27557(.A0(new_n29993_), .A1(new_n29990_), .B0(new_n29989_), .Y(new_n29994_));
  INVX1    g27558(.A(pi0577), .Y(new_n29995_));
  AOI21X1  g27559(.A0(new_n29987_), .A1(pi0238), .B0(new_n29995_), .Y(new_n29996_));
  NOR3X1   g27560(.A(new_n29983_), .B(new_n29915_), .C(pi0238), .Y(new_n29997_));
  OAI21X1  g27561(.A0(new_n29992_), .A1(new_n3551_), .B0(new_n29995_), .Y(new_n29998_));
  OAI21X1  g27562(.A0(new_n29998_), .A1(new_n29997_), .B0(pi0498), .Y(new_n29999_));
  OAI22X1  g27563(.A0(new_n29999_), .A1(new_n29996_), .B0(new_n29994_), .B1(new_n29988_), .Y(new_n30000_));
  AOI21X1  g27564(.A0(new_n30000_), .A1(new_n22655_), .B0(pi0237), .Y(new_n30001_));
  AOI22X1  g27565(.A0(new_n30001_), .A1(new_n29888_), .B0(new_n29757_), .B1(new_n29633_), .Y(po0750));
  NOR2X1   g27566(.A(new_n29141_), .B(pi0806), .Y(new_n30003_));
  INVX1    g27567(.A(pi0990), .Y(new_n30004_));
  OR4X1    g27568(.A(new_n30004_), .B(pi0806), .C(new_n29135_), .D(pi0332), .Y(new_n30005_));
  NAND2X1  g27569(.A(pi0594), .B(new_n2444_), .Y(new_n30006_));
  AOI21X1  g27570(.A0(new_n30006_), .A1(new_n30005_), .B0(new_n30003_), .Y(po0751));
  INVX1    g27571(.A(pi0595), .Y(new_n30008_));
  INVX1    g27572(.A(pi0605), .Y(new_n30009_));
  OR3X1    g27573(.A(new_n29125_), .B(pi0806), .C(new_n30009_), .Y(new_n30010_));
  OAI21X1  g27574(.A0(new_n30010_), .A1(new_n30008_), .B0(new_n2444_), .Y(new_n30011_));
  AOI21X1  g27575(.A0(new_n30010_), .A1(new_n30008_), .B0(new_n30011_), .Y(po0752));
  AND2X1   g27576(.A(pi0596), .B(new_n2444_), .Y(new_n30013_));
  NAND4X1  g27577(.A(pi0600), .B(pi0597), .C(pi0595), .D(pi0594), .Y(new_n30014_));
  NOR4X1   g27578(.A(new_n30014_), .B(new_n30004_), .C(pi0806), .D(pi0332), .Y(new_n30015_));
  MX2X1    g27579(.A(new_n30013_), .B(new_n29128_), .S0(new_n30015_), .Y(po0753));
  INVX1    g27580(.A(pi0597), .Y(new_n30017_));
  OAI21X1  g27581(.A0(new_n29141_), .A1(pi0806), .B0(new_n30017_), .Y(new_n30018_));
  OR3X1    g27582(.A(new_n29141_), .B(pi0806), .C(new_n30017_), .Y(new_n30019_));
  AND3X1   g27583(.A(new_n30019_), .B(new_n30018_), .C(new_n2444_), .Y(po0754));
  OR3X1    g27584(.A(new_n5103_), .B(pi0882), .C(pi0057), .Y(new_n30021_));
  OAI21X1  g27585(.A0(new_n30021_), .A1(new_n5362_), .B0(pi0598), .Y(new_n30022_));
  NAND3X1  g27586(.A(new_n5018_), .B(pi0780), .C(pi0740), .Y(new_n30023_));
  NAND2X1  g27587(.A(new_n30023_), .B(new_n30022_), .Y(po0755));
  AND2X1   g27588(.A(new_n30015_), .B(pi0596), .Y(new_n30025_));
  AND2X1   g27589(.A(pi0599), .B(new_n2444_), .Y(new_n30026_));
  MX2X1    g27590(.A(new_n30026_), .B(new_n29129_), .S0(new_n30025_), .Y(po0756));
  INVX1    g27591(.A(pi0806), .Y(new_n30028_));
  AND3X1   g27592(.A(pi0990), .B(new_n30028_), .C(new_n2444_), .Y(new_n30029_));
  AND2X1   g27593(.A(pi0600), .B(new_n2444_), .Y(new_n30030_));
  MX2X1    g27594(.A(new_n30030_), .B(new_n29135_), .S0(new_n30029_), .Y(po0757));
  NOR2X1   g27595(.A(pi0989), .B(pi0806), .Y(new_n30032_));
  OAI21X1  g27596(.A0(new_n30028_), .A1(pi0601), .B0(new_n2444_), .Y(new_n30033_));
  NOR2X1   g27597(.A(new_n30033_), .B(new_n30032_), .Y(po0758));
  NOR3X1   g27598(.A(new_n12737_), .B(new_n12275_), .C(new_n24814_), .Y(new_n30035_));
  AOI21X1  g27599(.A0(pi1160), .A1(pi0715), .B0(new_n12766_), .Y(new_n30036_));
  OAI21X1  g27600(.A0(pi1160), .A1(pi0715), .B0(new_n30036_), .Y(new_n30037_));
  NAND4X1  g27601(.A(new_n30037_), .B(new_n30035_), .C(new_n14140_), .D(new_n13434_), .Y(new_n30038_));
  OAI22X1  g27602(.A0(new_n30038_), .A1(new_n13489_), .B0(new_n5273_), .B1(pi0230), .Y(po0759));
  INVX1    g27603(.A(pi0952), .Y(new_n30040_));
  INVX1    g27604(.A(pi0980), .Y(new_n30041_));
  NAND3X1  g27605(.A(pi1060), .B(pi1038), .C(new_n30041_), .Y(new_n30042_));
  NOR4X1   g27606(.A(new_n30042_), .B(pi1061), .C(new_n30040_), .D(new_n12767_), .Y(po0897));
  NOR2X1   g27607(.A(po0897), .B(pi0603), .Y(new_n30044_));
  OR2X1    g27608(.A(pi1100), .B(new_n12767_), .Y(new_n30045_));
  NOR4X1   g27609(.A(new_n30045_), .B(new_n30042_), .C(pi1061), .D(new_n30040_), .Y(new_n30046_));
  OR2X1    g27610(.A(new_n30046_), .B(pi0966), .Y(new_n30047_));
  OAI21X1  g27611(.A0(pi0872), .A1(pi0871), .B0(pi0966), .Y(new_n30048_));
  OAI21X1  g27612(.A0(new_n30047_), .A1(new_n30044_), .B0(new_n30048_), .Y(po0760));
  NAND2X1  g27613(.A(new_n11863_), .B(pi0823), .Y(new_n30050_));
  NAND3X1  g27614(.A(pi0983), .B(pi0907), .C(new_n2933_), .Y(new_n30051_));
  NAND3X1  g27615(.A(new_n30051_), .B(new_n30050_), .C(pi0604), .Y(new_n30052_));
  OAI21X1  g27616(.A0(new_n30050_), .A1(pi0779), .B0(new_n30052_), .Y(po0761));
  OAI21X1  g27617(.A0(pi0806), .A1(pi0332), .B0(new_n30009_), .Y(new_n30054_));
  AOI21X1  g27618(.A0(new_n30028_), .A1(pi0605), .B0(pi0332), .Y(new_n30055_));
  AND2X1   g27619(.A(new_n30055_), .B(new_n30054_), .Y(po0762));
  MX2X1    g27620(.A(pi0606), .B(pi1104), .S0(po0897), .Y(new_n30057_));
  MX2X1    g27621(.A(new_n30057_), .B(pi0837), .S0(pi0966), .Y(po0763));
  INVX1    g27622(.A(po0897), .Y(new_n30059_));
  INVX1    g27623(.A(pi0966), .Y(new_n30060_));
  OAI21X1  g27624(.A0(new_n30059_), .A1(pi1107), .B0(new_n30060_), .Y(new_n30061_));
  AOI21X1  g27625(.A0(new_n30059_), .A1(new_n22960_), .B0(new_n30061_), .Y(po0764));
  OAI21X1  g27626(.A0(new_n30059_), .A1(pi1116), .B0(new_n30060_), .Y(new_n30063_));
  AOI21X1  g27627(.A0(new_n30059_), .A1(new_n12368_), .B0(new_n30063_), .Y(po0765));
  OAI21X1  g27628(.A0(new_n30059_), .A1(pi1118), .B0(new_n30060_), .Y(new_n30065_));
  AOI21X1  g27629(.A0(new_n30059_), .A1(new_n12462_), .B0(new_n30065_), .Y(po0766));
  INVX1    g27630(.A(pi0610), .Y(new_n30067_));
  OAI21X1  g27631(.A0(new_n30059_), .A1(pi1113), .B0(new_n30060_), .Y(new_n30068_));
  AOI21X1  g27632(.A0(new_n30059_), .A1(new_n30067_), .B0(new_n30068_), .Y(po0767));
  INVX1    g27633(.A(pi0611), .Y(new_n30070_));
  OAI21X1  g27634(.A0(new_n30059_), .A1(pi1114), .B0(new_n30060_), .Y(new_n30071_));
  AOI21X1  g27635(.A0(new_n30059_), .A1(new_n30070_), .B0(new_n30071_), .Y(po0768));
  OAI21X1  g27636(.A0(new_n30059_), .A1(pi1111), .B0(new_n30060_), .Y(new_n30073_));
  AOI21X1  g27637(.A0(new_n30059_), .A1(new_n23370_), .B0(new_n30073_), .Y(po0769));
  INVX1    g27638(.A(pi0613), .Y(new_n30075_));
  OAI21X1  g27639(.A0(new_n30059_), .A1(pi1115), .B0(new_n30060_), .Y(new_n30076_));
  AOI21X1  g27640(.A0(new_n30059_), .A1(new_n30075_), .B0(new_n30076_), .Y(po0770));
  INVX1    g27641(.A(pi0871), .Y(new_n30078_));
  NOR2X1   g27642(.A(po0897), .B(pi0614), .Y(new_n30079_));
  OAI21X1  g27643(.A0(new_n30059_), .A1(pi1102), .B0(new_n30060_), .Y(new_n30080_));
  OAI22X1  g27644(.A0(new_n30080_), .A1(new_n30079_), .B0(new_n30060_), .B1(new_n30078_), .Y(po0771));
  NOR4X1   g27645(.A(new_n5103_), .B(new_n5277_), .C(pi0882), .D(pi0057), .Y(new_n30082_));
  NAND3X1  g27646(.A(new_n5020_), .B(pi0797), .C(pi0779), .Y(new_n30083_));
  OAI21X1  g27647(.A0(new_n30082_), .A1(pi0615), .B0(new_n30083_), .Y(po0772));
  INVX1    g27648(.A(pi0872), .Y(new_n30085_));
  NOR2X1   g27649(.A(po0897), .B(pi0616), .Y(new_n30086_));
  OAI21X1  g27650(.A0(new_n30059_), .A1(pi1101), .B0(new_n30060_), .Y(new_n30087_));
  OAI22X1  g27651(.A0(new_n30087_), .A1(new_n30086_), .B0(new_n30060_), .B1(new_n30085_), .Y(po0773));
  MX2X1    g27652(.A(pi0617), .B(pi1105), .S0(po0897), .Y(new_n30089_));
  MX2X1    g27653(.A(new_n30089_), .B(pi0850), .S0(pi0966), .Y(po0774));
  OAI21X1  g27654(.A0(new_n30059_), .A1(pi1117), .B0(new_n30060_), .Y(new_n30091_));
  AOI21X1  g27655(.A0(new_n30059_), .A1(new_n12486_), .B0(new_n30091_), .Y(po0775));
  OAI21X1  g27656(.A0(new_n30059_), .A1(pi1122), .B0(new_n30060_), .Y(new_n30093_));
  AOI21X1  g27657(.A0(new_n30059_), .A1(new_n12509_), .B0(new_n30093_), .Y(po0776));
  INVX1    g27658(.A(pi0620), .Y(new_n30095_));
  OAI21X1  g27659(.A0(new_n30059_), .A1(pi1112), .B0(new_n30060_), .Y(new_n30096_));
  AOI21X1  g27660(.A0(new_n30059_), .A1(new_n30095_), .B0(new_n30096_), .Y(po0777));
  OAI21X1  g27661(.A0(new_n30059_), .A1(pi1108), .B0(new_n30060_), .Y(new_n30098_));
  AOI21X1  g27662(.A0(new_n30059_), .A1(new_n11963_), .B0(new_n30098_), .Y(po0778));
  OAI21X1  g27663(.A0(new_n30059_), .A1(pi1109), .B0(new_n30060_), .Y(new_n30100_));
  AOI21X1  g27664(.A0(new_n30059_), .A1(new_n23047_), .B0(new_n30100_), .Y(po0779));
  OAI21X1  g27665(.A0(new_n30059_), .A1(pi1106), .B0(new_n30060_), .Y(new_n30102_));
  AOI21X1  g27666(.A0(new_n30059_), .A1(new_n22661_), .B0(new_n30102_), .Y(po0780));
  NAND2X1  g27667(.A(new_n11999_), .B(pi0831), .Y(new_n30104_));
  NAND3X1  g27668(.A(pi0983), .B(pi0947), .C(new_n2933_), .Y(new_n30105_));
  NAND3X1  g27669(.A(new_n30105_), .B(new_n30104_), .C(pi0624), .Y(new_n30106_));
  OAI21X1  g27670(.A0(new_n30104_), .A1(pi0780), .B0(new_n30106_), .Y(po0781));
  INVX1    g27671(.A(pi1054), .Y(new_n30108_));
  NAND3X1  g27672(.A(pi1088), .B(pi1066), .C(new_n30108_), .Y(new_n30109_));
  NOR4X1   g27673(.A(new_n30109_), .B(pi0973), .C(pi0953), .D(new_n12767_), .Y(po0954));
  INVX1    g27674(.A(po0954), .Y(new_n30111_));
  INVX1    g27675(.A(pi0962), .Y(new_n30112_));
  OAI21X1  g27676(.A0(new_n30111_), .A1(pi1116), .B0(new_n30112_), .Y(new_n30113_));
  AOI21X1  g27677(.A0(new_n30111_), .A1(new_n12363_), .B0(new_n30113_), .Y(po0782));
  OAI21X1  g27678(.A0(new_n30059_), .A1(pi1121), .B0(new_n30060_), .Y(new_n30115_));
  AOI21X1  g27679(.A0(new_n30059_), .A1(new_n12542_), .B0(new_n30115_), .Y(po0783));
  OAI21X1  g27680(.A0(new_n30111_), .A1(pi1117), .B0(new_n30112_), .Y(new_n30117_));
  AOI21X1  g27681(.A0(new_n30111_), .A1(new_n12494_), .B0(new_n30117_), .Y(po0784));
  OAI21X1  g27682(.A0(new_n30111_), .A1(pi1119), .B0(new_n30112_), .Y(new_n30119_));
  AOI21X1  g27683(.A0(new_n30111_), .A1(new_n12554_), .B0(new_n30119_), .Y(po0785));
  OAI21X1  g27684(.A0(new_n30059_), .A1(pi1119), .B0(new_n30060_), .Y(new_n30121_));
  AOI21X1  g27685(.A0(new_n30059_), .A1(new_n12561_), .B0(new_n30121_), .Y(po0786));
  OAI21X1  g27686(.A0(new_n30059_), .A1(pi1120), .B0(new_n30060_), .Y(new_n30123_));
  AOI21X1  g27687(.A0(new_n30059_), .A1(new_n12592_), .B0(new_n30123_), .Y(po0787));
  INVX1    g27688(.A(pi1113), .Y(new_n30125_));
  INVX1    g27689(.A(pi0631), .Y(new_n30126_));
  OAI21X1  g27690(.A0(po0954), .A1(new_n30126_), .B0(new_n30112_), .Y(new_n30127_));
  AOI21X1  g27691(.A0(po0954), .A1(new_n30125_), .B0(new_n30127_), .Y(po0788));
  INVX1    g27692(.A(pi1115), .Y(new_n30129_));
  INVX1    g27693(.A(pi0632), .Y(new_n30130_));
  OAI21X1  g27694(.A0(po0954), .A1(new_n30130_), .B0(new_n30112_), .Y(new_n30131_));
  AOI21X1  g27695(.A0(po0954), .A1(new_n30129_), .B0(new_n30131_), .Y(po0789));
  OAI21X1  g27696(.A0(new_n30059_), .A1(pi1110), .B0(new_n30060_), .Y(new_n30133_));
  AOI21X1  g27697(.A0(new_n30059_), .A1(new_n21784_), .B0(new_n30133_), .Y(po0790));
  OAI21X1  g27698(.A0(new_n30111_), .A1(pi1110), .B0(new_n30112_), .Y(new_n30135_));
  AOI21X1  g27699(.A0(new_n30111_), .A1(new_n21904_), .B0(new_n30135_), .Y(po0791));
  INVX1    g27700(.A(pi1112), .Y(new_n30137_));
  INVX1    g27701(.A(pi0635), .Y(new_n30138_));
  OAI21X1  g27702(.A0(po0954), .A1(new_n30138_), .B0(new_n30112_), .Y(new_n30139_));
  AOI21X1  g27703(.A0(po0954), .A1(new_n30137_), .B0(new_n30139_), .Y(po0792));
  OR2X1    g27704(.A(po0897), .B(pi0636), .Y(new_n30141_));
  INVX1    g27705(.A(pi1127), .Y(new_n30142_));
  AOI21X1  g27706(.A0(po0897), .A1(new_n30142_), .B0(pi0966), .Y(new_n30143_));
  AND2X1   g27707(.A(new_n30143_), .B(new_n30141_), .Y(po0793));
  OAI21X1  g27708(.A0(new_n30111_), .A1(pi1105), .B0(new_n30112_), .Y(new_n30145_));
  AOI21X1  g27709(.A0(new_n30111_), .A1(new_n22139_), .B0(new_n30145_), .Y(po0794));
  OAI21X1  g27710(.A0(new_n30111_), .A1(pi1107), .B0(new_n30112_), .Y(new_n30147_));
  AOI21X1  g27711(.A0(new_n30111_), .A1(new_n22966_), .B0(new_n30147_), .Y(po0795));
  OAI21X1  g27712(.A0(new_n30111_), .A1(pi1109), .B0(new_n30112_), .Y(new_n30149_));
  AOI21X1  g27713(.A0(new_n30111_), .A1(new_n23002_), .B0(new_n30149_), .Y(po0796));
  OR2X1    g27714(.A(po0897), .B(pi0640), .Y(new_n30151_));
  INVX1    g27715(.A(pi1128), .Y(new_n30152_));
  AOI21X1  g27716(.A0(po0897), .A1(new_n30152_), .B0(pi0966), .Y(new_n30153_));
  AND2X1   g27717(.A(new_n30153_), .B(new_n30151_), .Y(po0797));
  OAI21X1  g27718(.A0(new_n30111_), .A1(pi1121), .B0(new_n30112_), .Y(new_n30155_));
  AOI21X1  g27719(.A0(new_n30111_), .A1(new_n12543_), .B0(new_n30155_), .Y(po0798));
  OAI21X1  g27720(.A0(new_n30059_), .A1(pi1103), .B0(new_n30060_), .Y(new_n30157_));
  AOI21X1  g27721(.A0(new_n30059_), .A1(new_n5016_), .B0(new_n30157_), .Y(po0799));
  OAI21X1  g27722(.A0(new_n30111_), .A1(pi1104), .B0(new_n30112_), .Y(new_n30159_));
  AOI21X1  g27723(.A0(new_n30111_), .A1(new_n22368_), .B0(new_n30159_), .Y(po0800));
  OAI21X1  g27724(.A0(new_n30059_), .A1(pi1123), .B0(new_n30060_), .Y(new_n30161_));
  AOI21X1  g27725(.A0(new_n30059_), .A1(new_n12612_), .B0(new_n30161_), .Y(po0801));
  OR2X1    g27726(.A(po0897), .B(pi0645), .Y(new_n30163_));
  INVX1    g27727(.A(pi1125), .Y(new_n30164_));
  AOI21X1  g27728(.A0(po0897), .A1(new_n30164_), .B0(pi0966), .Y(new_n30165_));
  AND2X1   g27729(.A(new_n30165_), .B(new_n30163_), .Y(po0802));
  INVX1    g27730(.A(pi1114), .Y(new_n30167_));
  INVX1    g27731(.A(pi0646), .Y(new_n30168_));
  OAI21X1  g27732(.A0(po0954), .A1(new_n30168_), .B0(new_n30112_), .Y(new_n30169_));
  AOI21X1  g27733(.A0(po0954), .A1(new_n30167_), .B0(new_n30169_), .Y(po0803));
  OAI21X1  g27734(.A0(new_n30111_), .A1(pi1120), .B0(new_n30112_), .Y(new_n30171_));
  AOI21X1  g27735(.A0(new_n30111_), .A1(new_n12577_), .B0(new_n30171_), .Y(po0804));
  OAI21X1  g27736(.A0(new_n30111_), .A1(pi1122), .B0(new_n30112_), .Y(new_n30173_));
  AOI21X1  g27737(.A0(new_n30111_), .A1(new_n12517_), .B0(new_n30173_), .Y(po0805));
  INVX1    g27738(.A(pi1126), .Y(new_n30175_));
  INVX1    g27739(.A(pi0649), .Y(new_n30176_));
  OAI21X1  g27740(.A0(po0954), .A1(new_n30176_), .B0(new_n30112_), .Y(new_n30177_));
  AOI21X1  g27741(.A0(po0954), .A1(new_n30175_), .B0(new_n30177_), .Y(po0806));
  INVX1    g27742(.A(pi0650), .Y(new_n30179_));
  OAI21X1  g27743(.A0(po0954), .A1(new_n30179_), .B0(new_n30112_), .Y(new_n30180_));
  AOI21X1  g27744(.A0(po0954), .A1(new_n30142_), .B0(new_n30180_), .Y(po0807));
  OR2X1    g27745(.A(po0897), .B(pi0651), .Y(new_n30182_));
  INVX1    g27746(.A(pi1130), .Y(new_n30183_));
  AOI21X1  g27747(.A0(po0897), .A1(new_n30183_), .B0(pi0966), .Y(new_n30184_));
  AND2X1   g27748(.A(new_n30184_), .B(new_n30182_), .Y(po0808));
  OR2X1    g27749(.A(po0897), .B(pi0652), .Y(new_n30186_));
  INVX1    g27750(.A(pi1131), .Y(new_n30187_));
  AOI21X1  g27751(.A0(po0897), .A1(new_n30187_), .B0(pi0966), .Y(new_n30188_));
  AND2X1   g27752(.A(new_n30188_), .B(new_n30186_), .Y(po0809));
  OR2X1    g27753(.A(po0897), .B(pi0653), .Y(new_n30190_));
  INVX1    g27754(.A(pi1129), .Y(new_n30191_));
  AOI21X1  g27755(.A0(po0897), .A1(new_n30191_), .B0(pi0966), .Y(new_n30192_));
  AND2X1   g27756(.A(new_n30192_), .B(new_n30190_), .Y(po0810));
  INVX1    g27757(.A(pi0654), .Y(new_n30194_));
  OAI21X1  g27758(.A0(po0954), .A1(new_n30194_), .B0(new_n30112_), .Y(new_n30195_));
  AOI21X1  g27759(.A0(po0954), .A1(new_n30183_), .B0(new_n30195_), .Y(po0811));
  INVX1    g27760(.A(pi1124), .Y(new_n30197_));
  INVX1    g27761(.A(pi0655), .Y(new_n30198_));
  OAI21X1  g27762(.A0(po0954), .A1(new_n30198_), .B0(new_n30112_), .Y(new_n30199_));
  AOI21X1  g27763(.A0(po0954), .A1(new_n30197_), .B0(new_n30199_), .Y(po0812));
  OR2X1    g27764(.A(po0897), .B(pi0656), .Y(new_n30201_));
  AOI21X1  g27765(.A0(po0897), .A1(new_n30175_), .B0(pi0966), .Y(new_n30202_));
  AND2X1   g27766(.A(new_n30202_), .B(new_n30201_), .Y(po0813));
  INVX1    g27767(.A(pi0657), .Y(new_n30204_));
  OAI21X1  g27768(.A0(po0954), .A1(new_n30204_), .B0(new_n30112_), .Y(new_n30205_));
  AOI21X1  g27769(.A0(po0954), .A1(new_n30187_), .B0(new_n30205_), .Y(po0814));
  OR2X1    g27770(.A(po0897), .B(pi0658), .Y(new_n30207_));
  AOI21X1  g27771(.A0(po0897), .A1(new_n30197_), .B0(pi0966), .Y(new_n30208_));
  AND2X1   g27772(.A(new_n30208_), .B(new_n30207_), .Y(po0815));
  INVX1    g27773(.A(pi0265), .Y(new_n30210_));
  INVX1    g27774(.A(pi0281), .Y(new_n30211_));
  AND2X1   g27775(.A(pi0992), .B(pi0266), .Y(new_n30212_));
  AND2X1   g27776(.A(new_n30212_), .B(new_n4406_), .Y(new_n30213_));
  AND3X1   g27777(.A(new_n30213_), .B(new_n30211_), .C(new_n4260_), .Y(new_n30214_));
  NOR3X1   g27778(.A(pi0282), .B(pi0277), .C(pi0270), .Y(new_n30215_));
  NAND4X1  g27779(.A(new_n30215_), .B(new_n30214_), .C(new_n30210_), .D(new_n3521_), .Y(new_n30216_));
  XOR2X1   g27780(.A(new_n30216_), .B(pi0274), .Y(po0816));
  OAI21X1  g27781(.A0(new_n30111_), .A1(pi1118), .B0(new_n30112_), .Y(new_n30218_));
  AOI21X1  g27782(.A0(new_n30111_), .A1(new_n12468_), .B0(new_n30218_), .Y(po0817));
  OAI21X1  g27783(.A0(new_n30111_), .A1(pi1101), .B0(new_n30112_), .Y(new_n30220_));
  AOI21X1  g27784(.A0(new_n30111_), .A1(new_n11848_), .B0(new_n30220_), .Y(po0818));
  OAI21X1  g27785(.A0(new_n30111_), .A1(pi1102), .B0(new_n30112_), .Y(new_n30222_));
  AOI21X1  g27786(.A0(new_n30111_), .A1(new_n11849_), .B0(new_n30222_), .Y(po0819));
  NOR2X1   g27787(.A(pi0257), .B(pi0199), .Y(new_n30224_));
  OAI22X1  g27788(.A0(pi1065), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30225_));
  NOR2X1   g27789(.A(new_n30225_), .B(new_n30224_), .Y(new_n30226_));
  AND2X1   g27790(.A(pi0592), .B(new_n6069_), .Y(new_n30227_));
  AND3X1   g27791(.A(new_n6009_), .B(pi0591), .C(pi0334), .Y(new_n30228_));
  AOI21X1  g27792(.A0(new_n30227_), .A1(pi0365), .B0(new_n30228_), .Y(new_n30229_));
  AND3X1   g27793(.A(new_n6009_), .B(new_n6069_), .C(pi0590), .Y(new_n30230_));
  AOI21X1  g27794(.A0(new_n30230_), .A1(pi0323), .B0(pi0588), .Y(new_n30231_));
  OAI21X1  g27795(.A0(new_n30229_), .A1(pi0590), .B0(new_n30231_), .Y(new_n30232_));
  NOR2X1   g27796(.A(pi0224), .B(pi0223), .Y(new_n30233_));
  INVX1    g27797(.A(new_n30233_), .Y(new_n30234_));
  NAND3X1  g27798(.A(new_n6561_), .B(new_n6009_), .C(pi0464), .Y(new_n30235_));
  AOI21X1  g27799(.A0(new_n30235_), .A1(pi0588), .B0(new_n30234_), .Y(new_n30236_));
  AOI21X1  g27800(.A0(new_n30236_), .A1(new_n30232_), .B0(new_n30226_), .Y(new_n30237_));
  NOR3X1   g27801(.A(pi1138), .B(pi1137), .C(pi1134), .Y(new_n30238_));
  INVX1    g27802(.A(new_n30238_), .Y(new_n30239_));
  AOI21X1  g27803(.A0(pi1136), .A1(new_n21904_), .B0(new_n4622_), .Y(new_n30240_));
  OAI21X1  g27804(.A0(pi1136), .A1(pi0784), .B0(new_n30240_), .Y(new_n30241_));
  AOI21X1  g27805(.A0(pi1136), .A1(new_n21784_), .B0(pi1135), .Y(new_n30242_));
  OAI21X1  g27806(.A0(pi1136), .A1(pi0815), .B0(new_n30242_), .Y(new_n30243_));
  AOI21X1  g27807(.A0(new_n30243_), .A1(new_n30241_), .B0(new_n30239_), .Y(new_n30244_));
  NOR2X1   g27808(.A(pi1138), .B(pi1137), .Y(new_n30245_));
  AOI21X1  g27809(.A0(new_n30245_), .A1(pi1135), .B0(new_n4554_), .Y(new_n30246_));
  AND2X1   g27810(.A(new_n30246_), .B(new_n14844_), .Y(new_n30247_));
  AND2X1   g27811(.A(new_n30245_), .B(pi1134), .Y(new_n30248_));
  INVX1    g27812(.A(new_n30248_), .Y(new_n30249_));
  AOI21X1  g27813(.A0(new_n4554_), .A1(pi1135), .B0(new_n30249_), .Y(new_n30250_));
  INVX1    g27814(.A(new_n30250_), .Y(new_n30251_));
  OAI22X1  g27815(.A0(pi1136), .A1(pi0855), .B0(new_n4622_), .B1(pi0700), .Y(new_n30252_));
  NOR3X1   g27816(.A(new_n30252_), .B(new_n30251_), .C(new_n30247_), .Y(new_n30253_));
  OAI21X1  g27817(.A0(new_n30253_), .A1(new_n30244_), .B0(new_n8943_), .Y(new_n30254_));
  OAI21X1  g27818(.A0(new_n30237_), .A1(new_n8943_), .B0(new_n30254_), .Y(po0820));
  INVX1    g27819(.A(new_n30230_), .Y(new_n30256_));
  AND2X1   g27820(.A(pi0591), .B(new_n6334_), .Y(new_n30257_));
  AOI21X1  g27821(.A0(pi0592), .A1(new_n6334_), .B0(pi0588), .Y(new_n30258_));
  INVX1    g27822(.A(new_n30258_), .Y(new_n30259_));
  AOI21X1  g27823(.A0(new_n30257_), .A1(pi0404), .B0(new_n30259_), .Y(new_n30260_));
  AOI21X1  g27824(.A0(new_n6069_), .A1(pi0380), .B0(new_n6009_), .Y(new_n30261_));
  OAI22X1  g27825(.A0(new_n30261_), .A1(new_n30260_), .B0(new_n30256_), .B1(new_n6013_), .Y(new_n30262_));
  OR3X1    g27826(.A(pi0592), .B(pi0591), .C(pi0590), .Y(new_n30263_));
  OAI21X1  g27827(.A0(new_n30263_), .A1(new_n8983_), .B0(pi0588), .Y(new_n30264_));
  AND2X1   g27828(.A(new_n30264_), .B(new_n30233_), .Y(new_n30265_));
  NOR2X1   g27829(.A(pi0292), .B(pi0199), .Y(new_n30266_));
  OAI22X1  g27830(.A0(pi1084), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30267_));
  NOR2X1   g27831(.A(new_n30267_), .B(new_n30266_), .Y(new_n30268_));
  AOI21X1  g27832(.A0(new_n30265_), .A1(new_n30262_), .B0(new_n30268_), .Y(new_n30269_));
  AOI21X1  g27833(.A0(pi1135), .A1(pi0662), .B0(new_n4554_), .Y(new_n30270_));
  OAI21X1  g27834(.A0(pi1135), .A1(new_n11838_), .B0(new_n30270_), .Y(new_n30271_));
  INVX1    g27835(.A(pi0811), .Y(new_n30272_));
  AOI21X1  g27836(.A0(pi1135), .A1(pi0785), .B0(pi1136), .Y(new_n30273_));
  OAI21X1  g27837(.A0(pi1135), .A1(new_n30272_), .B0(new_n30273_), .Y(new_n30274_));
  AOI21X1  g27838(.A0(new_n30274_), .A1(new_n30271_), .B0(pi1134), .Y(new_n30275_));
  OAI21X1  g27839(.A0(new_n4622_), .A1(pi0727), .B0(pi1136), .Y(new_n30276_));
  AOI21X1  g27840(.A0(new_n4622_), .A1(new_n15306_), .B0(new_n30276_), .Y(new_n30277_));
  NOR2X1   g27841(.A(pi1136), .B(pi1135), .Y(new_n30278_));
  INVX1    g27842(.A(new_n30278_), .Y(new_n30279_));
  OAI21X1  g27843(.A0(new_n30279_), .A1(new_n30085_), .B0(pi1134), .Y(new_n30280_));
  NOR3X1   g27844(.A(new_n6713_), .B(pi1138), .C(pi1137), .Y(new_n30281_));
  OAI21X1  g27845(.A0(new_n30280_), .A1(new_n30277_), .B0(new_n30281_), .Y(new_n30282_));
  OAI22X1  g27846(.A0(new_n30282_), .A1(new_n30275_), .B0(new_n30269_), .B1(new_n8943_), .Y(po0821));
  OAI21X1  g27847(.A0(new_n30111_), .A1(pi1108), .B0(new_n30112_), .Y(new_n30284_));
  AOI21X1  g27848(.A0(new_n30111_), .A1(new_n12091_), .B0(new_n30284_), .Y(po0822));
  AOI21X1  g27849(.A0(pi1135), .A1(new_n22966_), .B0(new_n4554_), .Y(new_n30286_));
  OAI21X1  g27850(.A0(pi1135), .A1(pi0607), .B0(new_n30286_), .Y(new_n30287_));
  AOI21X1  g27851(.A0(new_n4622_), .A1(pi0799), .B0(pi1136), .Y(new_n30288_));
  OAI21X1  g27852(.A0(new_n4622_), .A1(pi0790), .B0(new_n30288_), .Y(new_n30289_));
  AOI21X1  g27853(.A0(new_n30289_), .A1(new_n30287_), .B0(new_n30239_), .Y(new_n30290_));
  AND2X1   g27854(.A(new_n30246_), .B(new_n15517_), .Y(new_n30291_));
  OAI22X1  g27855(.A0(pi1136), .A1(pi0873), .B0(new_n4622_), .B1(pi0691), .Y(new_n30292_));
  NOR3X1   g27856(.A(new_n30292_), .B(new_n30291_), .C(new_n30251_), .Y(new_n30293_));
  OAI21X1  g27857(.A0(new_n30293_), .A1(new_n30290_), .B0(new_n8943_), .Y(new_n30294_));
  OR2X1    g27858(.A(pi0297), .B(pi0199), .Y(new_n30295_));
  AOI21X1  g27859(.A0(new_n27850_), .A1(pi0199), .B0(new_n30233_), .Y(new_n30296_));
  AOI21X1  g27860(.A0(new_n30257_), .A1(pi0456), .B0(new_n30259_), .Y(new_n30297_));
  AOI21X1  g27861(.A0(new_n6069_), .A1(pi0337), .B0(new_n6009_), .Y(new_n30298_));
  OAI22X1  g27862(.A0(new_n30298_), .A1(new_n30297_), .B0(new_n30256_), .B1(new_n6609_), .Y(new_n30299_));
  OAI21X1  g27863(.A0(new_n30263_), .A1(new_n8984_), .B0(pi0588), .Y(new_n30300_));
  AND2X1   g27864(.A(new_n30300_), .B(new_n30233_), .Y(new_n30301_));
  AOI22X1  g27865(.A0(new_n30301_), .A1(new_n30299_), .B0(new_n30296_), .B1(new_n30295_), .Y(new_n30302_));
  OAI21X1  g27866(.A0(new_n30302_), .A1(new_n8943_), .B0(new_n30294_), .Y(po0823));
  AOI21X1  g27867(.A0(new_n30257_), .A1(pi0319), .B0(new_n30259_), .Y(new_n30304_));
  AOI21X1  g27868(.A0(new_n6069_), .A1(pi0338), .B0(new_n6009_), .Y(new_n30305_));
  OAI22X1  g27869(.A0(new_n30305_), .A1(new_n30304_), .B0(new_n30256_), .B1(new_n6029_), .Y(new_n30306_));
  OAI21X1  g27870(.A0(new_n30263_), .A1(new_n6520_), .B0(pi0588), .Y(new_n30307_));
  AND2X1   g27871(.A(new_n30307_), .B(new_n30233_), .Y(new_n30308_));
  NOR2X1   g27872(.A(pi0294), .B(pi0199), .Y(new_n30309_));
  OAI22X1  g27873(.A0(pi1072), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30310_));
  NOR2X1   g27874(.A(new_n30310_), .B(new_n30309_), .Y(new_n30311_));
  AOI21X1  g27875(.A0(new_n30308_), .A1(new_n30306_), .B0(new_n30311_), .Y(new_n30312_));
  AOI21X1  g27876(.A0(pi1136), .A1(pi0681), .B0(new_n4622_), .Y(new_n30313_));
  OAI21X1  g27877(.A0(pi1136), .A1(new_n11764_), .B0(new_n30313_), .Y(new_n30314_));
  AOI21X1  g27878(.A0(pi1136), .A1(pi0642), .B0(pi1135), .Y(new_n30315_));
  OAI21X1  g27879(.A0(pi1136), .A1(pi0809), .B0(new_n30315_), .Y(new_n30316_));
  AOI21X1  g27880(.A0(new_n30316_), .A1(new_n30314_), .B0(pi1134), .Y(new_n30317_));
  OAI21X1  g27881(.A0(new_n4622_), .A1(pi0699), .B0(pi1136), .Y(new_n30318_));
  AOI21X1  g27882(.A0(new_n4622_), .A1(new_n15365_), .B0(new_n30318_), .Y(new_n30319_));
  OAI21X1  g27883(.A0(new_n30279_), .A1(new_n30078_), .B0(pi1134), .Y(new_n30320_));
  OAI21X1  g27884(.A0(new_n30320_), .A1(new_n30319_), .B0(new_n30281_), .Y(new_n30321_));
  OAI22X1  g27885(.A0(new_n30321_), .A1(new_n30317_), .B0(new_n30312_), .B1(new_n8943_), .Y(po0824));
  AOI21X1  g27886(.A0(pi1135), .A1(new_n5019_), .B0(new_n4554_), .Y(new_n30323_));
  OAI21X1  g27887(.A0(pi1135), .A1(pi0603), .B0(new_n30323_), .Y(new_n30324_));
  AOI21X1  g27888(.A0(pi1135), .A1(new_n11769_), .B0(pi1136), .Y(new_n30325_));
  OAI21X1  g27889(.A0(pi1135), .A1(pi0981), .B0(new_n30325_), .Y(new_n30326_));
  AOI21X1  g27890(.A0(new_n30326_), .A1(new_n30324_), .B0(new_n30239_), .Y(new_n30327_));
  AND2X1   g27891(.A(new_n30246_), .B(new_n14767_), .Y(new_n30328_));
  OAI22X1  g27892(.A0(pi1136), .A1(pi0837), .B0(new_n4622_), .B1(pi0696), .Y(new_n30329_));
  NOR3X1   g27893(.A(new_n30329_), .B(new_n30328_), .C(new_n30251_), .Y(new_n30330_));
  OAI21X1  g27894(.A0(new_n30330_), .A1(new_n30327_), .B0(new_n8943_), .Y(new_n30331_));
  NOR2X1   g27895(.A(pi0291), .B(pi0199), .Y(new_n30332_));
  OAI22X1  g27896(.A0(pi1049), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30333_));
  NOR2X1   g27897(.A(new_n30333_), .B(new_n30332_), .Y(new_n30334_));
  INVX1    g27898(.A(pi0342), .Y(new_n30335_));
  AOI21X1  g27899(.A0(new_n30257_), .A1(pi0390), .B0(new_n30259_), .Y(new_n30336_));
  AOI21X1  g27900(.A0(new_n6069_), .A1(pi0363), .B0(new_n6009_), .Y(new_n30337_));
  OAI22X1  g27901(.A0(new_n30337_), .A1(new_n30336_), .B0(new_n30256_), .B1(new_n30335_), .Y(new_n30338_));
  OAI21X1  g27902(.A0(new_n30263_), .A1(new_n6530_), .B0(pi0588), .Y(new_n30339_));
  AND2X1   g27903(.A(new_n30339_), .B(new_n30233_), .Y(new_n30340_));
  AOI21X1  g27904(.A0(new_n30340_), .A1(new_n30338_), .B0(new_n30334_), .Y(new_n30341_));
  OAI21X1  g27905(.A0(new_n30341_), .A1(new_n8943_), .B0(new_n30331_), .Y(po0825));
  INVX1    g27906(.A(pi0669), .Y(new_n30343_));
  OAI21X1  g27907(.A0(po0954), .A1(new_n30343_), .B0(new_n30112_), .Y(new_n30344_));
  AOI21X1  g27908(.A0(po0954), .A1(new_n30164_), .B0(new_n30344_), .Y(po0826));
  NOR2X1   g27909(.A(pi0258), .B(pi0199), .Y(new_n30346_));
  OAI22X1  g27910(.A0(pi1062), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30347_));
  NOR2X1   g27911(.A(new_n30347_), .B(new_n30346_), .Y(new_n30348_));
  AND3X1   g27912(.A(new_n6009_), .B(pi0591), .C(pi0391), .Y(new_n30349_));
  AOI21X1  g27913(.A0(new_n30227_), .A1(pi0364), .B0(new_n30349_), .Y(new_n30350_));
  AOI21X1  g27914(.A0(new_n30230_), .A1(pi0343), .B0(pi0588), .Y(new_n30351_));
  OAI21X1  g27915(.A0(new_n30350_), .A1(pi0590), .B0(new_n30351_), .Y(new_n30352_));
  NAND3X1  g27916(.A(new_n6561_), .B(new_n6009_), .C(pi0415), .Y(new_n30353_));
  AOI21X1  g27917(.A0(new_n30353_), .A1(pi0588), .B0(new_n30234_), .Y(new_n30354_));
  AOI21X1  g27918(.A0(new_n30354_), .A1(new_n30352_), .B0(new_n30348_), .Y(new_n30355_));
  AND2X1   g27919(.A(new_n30246_), .B(pi0745), .Y(new_n30356_));
  OAI22X1  g27920(.A0(pi1136), .A1(pi0852), .B0(new_n4622_), .B1(new_n14743_), .Y(new_n30357_));
  NOR3X1   g27921(.A(new_n30357_), .B(new_n30356_), .C(new_n30251_), .Y(new_n30358_));
  AND2X1   g27922(.A(new_n30245_), .B(pi1136), .Y(new_n30359_));
  NAND2X1  g27923(.A(pi1135), .B(pi0695), .Y(new_n30360_));
  AOI21X1  g27924(.A0(new_n4622_), .A1(new_n23370_), .B0(pi1134), .Y(new_n30361_));
  AND3X1   g27925(.A(new_n30361_), .B(new_n30360_), .C(new_n30359_), .Y(new_n30362_));
  OAI21X1  g27926(.A0(new_n30362_), .A1(new_n30358_), .B0(new_n8943_), .Y(new_n30363_));
  OAI21X1  g27927(.A0(new_n30355_), .A1(new_n8943_), .B0(new_n30363_), .Y(po0827));
  NOR2X1   g27928(.A(pi0261), .B(pi0199), .Y(new_n30365_));
  OAI22X1  g27929(.A0(pi1040), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30366_));
  NOR2X1   g27930(.A(new_n30366_), .B(new_n30365_), .Y(new_n30367_));
  AND3X1   g27931(.A(new_n6009_), .B(pi0591), .C(pi0333), .Y(new_n30368_));
  AOI21X1  g27932(.A0(new_n30227_), .A1(pi0447), .B0(new_n30368_), .Y(new_n30369_));
  AOI21X1  g27933(.A0(new_n30230_), .A1(pi0327), .B0(pi0588), .Y(new_n30370_));
  OAI21X1  g27934(.A0(new_n30369_), .A1(pi0590), .B0(new_n30370_), .Y(new_n30371_));
  OAI21X1  g27935(.A0(new_n30263_), .A1(new_n6500_), .B0(pi0588), .Y(new_n30372_));
  AND2X1   g27936(.A(new_n30372_), .B(new_n30233_), .Y(new_n30373_));
  AOI21X1  g27937(.A0(new_n30373_), .A1(new_n30371_), .B0(new_n30367_), .Y(new_n30374_));
  AND2X1   g27938(.A(new_n30246_), .B(pi0741), .Y(new_n30375_));
  OAI22X1  g27939(.A0(pi1136), .A1(pi0865), .B0(new_n4622_), .B1(new_n14956_), .Y(new_n30376_));
  NOR3X1   g27940(.A(new_n30376_), .B(new_n30375_), .C(new_n30251_), .Y(new_n30377_));
  NAND2X1  g27941(.A(pi1135), .B(pi0646), .Y(new_n30378_));
  AOI21X1  g27942(.A0(new_n4622_), .A1(new_n30070_), .B0(pi1134), .Y(new_n30379_));
  AND3X1   g27943(.A(new_n30379_), .B(new_n30378_), .C(new_n30359_), .Y(new_n30380_));
  OAI21X1  g27944(.A0(new_n30380_), .A1(new_n30377_), .B0(new_n8943_), .Y(new_n30381_));
  OAI21X1  g27945(.A0(new_n30374_), .A1(new_n8943_), .B0(new_n30381_), .Y(po0828));
  AOI21X1  g27946(.A0(pi1135), .A1(new_n11848_), .B0(new_n4554_), .Y(new_n30383_));
  OAI21X1  g27947(.A0(pi1135), .A1(pi0616), .B0(new_n30383_), .Y(new_n30384_));
  AOI21X1  g27948(.A0(pi1135), .A1(new_n11767_), .B0(pi1136), .Y(new_n30385_));
  OAI21X1  g27949(.A0(pi1135), .A1(pi0808), .B0(new_n30385_), .Y(new_n30386_));
  AOI21X1  g27950(.A0(new_n30386_), .A1(new_n30384_), .B0(new_n30239_), .Y(new_n30387_));
  AND2X1   g27951(.A(new_n30246_), .B(new_n13836_), .Y(new_n30388_));
  OAI22X1  g27952(.A0(pi1136), .A1(pi0850), .B0(new_n4622_), .B1(pi0736), .Y(new_n30389_));
  NOR3X1   g27953(.A(new_n30389_), .B(new_n30388_), .C(new_n30251_), .Y(new_n30390_));
  OAI21X1  g27954(.A0(new_n30390_), .A1(new_n30387_), .B0(new_n8943_), .Y(new_n30391_));
  NOR2X1   g27955(.A(pi0290), .B(pi0199), .Y(new_n30392_));
  OAI22X1  g27956(.A0(pi1048), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30393_));
  NOR2X1   g27957(.A(new_n30393_), .B(new_n30392_), .Y(new_n30394_));
  INVX1    g27958(.A(pi0320), .Y(new_n30395_));
  AOI21X1  g27959(.A0(new_n30257_), .A1(pi0397), .B0(new_n30259_), .Y(new_n30396_));
  AOI21X1  g27960(.A0(new_n6069_), .A1(pi0372), .B0(new_n6009_), .Y(new_n30397_));
  OAI22X1  g27961(.A0(new_n30397_), .A1(new_n30396_), .B0(new_n30256_), .B1(new_n30395_), .Y(new_n30398_));
  NAND3X1  g27962(.A(new_n6561_), .B(new_n6009_), .C(pi0422), .Y(new_n30399_));
  AOI21X1  g27963(.A0(new_n30399_), .A1(pi0588), .B0(new_n30234_), .Y(new_n30400_));
  AOI21X1  g27964(.A0(new_n30400_), .A1(new_n30398_), .B0(new_n30394_), .Y(new_n30401_));
  OAI21X1  g27965(.A0(new_n30401_), .A1(new_n8943_), .B0(new_n30391_), .Y(po0829));
  AOI21X1  g27966(.A0(pi1135), .A1(new_n22139_), .B0(new_n4554_), .Y(new_n30403_));
  OAI21X1  g27967(.A0(pi1135), .A1(pi0617), .B0(new_n30403_), .Y(new_n30404_));
  AOI21X1  g27968(.A0(new_n4622_), .A1(pi0814), .B0(pi1136), .Y(new_n30405_));
  OAI21X1  g27969(.A0(new_n4622_), .A1(pi0788), .B0(new_n30405_), .Y(new_n30406_));
  AOI21X1  g27970(.A0(new_n30406_), .A1(new_n30404_), .B0(new_n30239_), .Y(new_n30407_));
  AND2X1   g27971(.A(new_n30246_), .B(new_n12774_), .Y(new_n30408_));
  OAI22X1  g27972(.A0(pi1136), .A1(pi0866), .B0(new_n4622_), .B1(pi0706), .Y(new_n30409_));
  NOR3X1   g27973(.A(new_n30409_), .B(new_n30408_), .C(new_n30251_), .Y(new_n30410_));
  OAI21X1  g27974(.A0(new_n30410_), .A1(new_n30407_), .B0(new_n8943_), .Y(new_n30411_));
  OR2X1    g27975(.A(pi0295), .B(pi0199), .Y(new_n30412_));
  AOI21X1  g27976(.A0(new_n27487_), .A1(pi0199), .B0(new_n30233_), .Y(new_n30413_));
  AOI21X1  g27977(.A0(new_n30257_), .A1(pi0411), .B0(new_n30259_), .Y(new_n30414_));
  AOI21X1  g27978(.A0(new_n6069_), .A1(pi0387), .B0(new_n6009_), .Y(new_n30415_));
  OAI22X1  g27979(.A0(new_n30415_), .A1(new_n30414_), .B0(new_n30256_), .B1(new_n6030_), .Y(new_n30416_));
  OAI21X1  g27980(.A0(new_n30263_), .A1(new_n8998_), .B0(pi0588), .Y(new_n30417_));
  AND2X1   g27981(.A(new_n30417_), .B(new_n30233_), .Y(new_n30418_));
  AOI22X1  g27982(.A0(new_n30418_), .A1(new_n30416_), .B0(new_n30413_), .B1(new_n30412_), .Y(new_n30419_));
  OAI21X1  g27983(.A0(new_n30419_), .A1(new_n8943_), .B0(new_n30411_), .Y(po0830));
  NOR2X1   g27984(.A(pi0256), .B(pi0199), .Y(new_n30421_));
  OAI22X1  g27985(.A0(pi1070), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30422_));
  NOR2X1   g27986(.A(new_n30422_), .B(new_n30421_), .Y(new_n30423_));
  AND3X1   g27987(.A(new_n6009_), .B(pi0591), .C(pi0463), .Y(new_n30424_));
  AOI21X1  g27988(.A0(new_n30227_), .A1(pi0336), .B0(new_n30424_), .Y(new_n30425_));
  AOI21X1  g27989(.A0(new_n30230_), .A1(pi0362), .B0(pi0588), .Y(new_n30426_));
  OAI21X1  g27990(.A0(new_n30425_), .A1(pi0590), .B0(new_n30426_), .Y(new_n30427_));
  NAND3X1  g27991(.A(new_n6561_), .B(new_n6009_), .C(pi0437), .Y(new_n30428_));
  AOI21X1  g27992(.A0(new_n30428_), .A1(pi0588), .B0(new_n30234_), .Y(new_n30429_));
  AOI21X1  g27993(.A0(new_n30429_), .A1(new_n30427_), .B0(new_n30423_), .Y(new_n30430_));
  AOI21X1  g27994(.A0(pi1135), .A1(pi0639), .B0(new_n4554_), .Y(new_n30431_));
  OAI21X1  g27995(.A0(pi1135), .A1(new_n23047_), .B0(new_n30431_), .Y(new_n30432_));
  AOI21X1  g27996(.A0(pi1135), .A1(pi0783), .B0(pi1136), .Y(new_n30433_));
  OAI21X1  g27997(.A0(pi1135), .A1(new_n29127_), .B0(new_n30433_), .Y(new_n30434_));
  AOI21X1  g27998(.A0(new_n30434_), .A1(new_n30432_), .B0(pi1134), .Y(new_n30435_));
  OAI21X1  g27999(.A0(new_n4622_), .A1(pi0735), .B0(pi1136), .Y(new_n30436_));
  AOI21X1  g28000(.A0(new_n4622_), .A1(new_n13086_), .B0(new_n30436_), .Y(new_n30437_));
  AND2X1   g28001(.A(new_n30278_), .B(pi0859), .Y(new_n30438_));
  OR2X1    g28002(.A(new_n30438_), .B(new_n4747_), .Y(new_n30439_));
  OAI21X1  g28003(.A0(new_n30439_), .A1(new_n30437_), .B0(new_n30281_), .Y(new_n30440_));
  OAI22X1  g28004(.A0(new_n30440_), .A1(new_n30435_), .B0(new_n30430_), .B1(new_n8943_), .Y(po0831));
  OR2X1    g28005(.A(pi1135), .B(pi0748), .Y(new_n30442_));
  AOI21X1  g28006(.A0(pi1135), .A1(new_n15466_), .B0(new_n4554_), .Y(new_n30443_));
  AOI22X1  g28007(.A0(new_n30443_), .A1(new_n30442_), .B0(new_n30278_), .B1(pi0876), .Y(new_n30444_));
  AND2X1   g28008(.A(new_n30246_), .B(new_n22661_), .Y(new_n30445_));
  AND3X1   g28009(.A(new_n4554_), .B(pi1135), .C(pi0789), .Y(new_n30446_));
  OAI21X1  g28010(.A0(new_n4622_), .A1(pi0710), .B0(pi1136), .Y(new_n30447_));
  OAI21X1  g28011(.A0(pi1135), .A1(pi0803), .B0(new_n30447_), .Y(new_n30448_));
  OAI21X1  g28012(.A0(new_n30448_), .A1(new_n30446_), .B0(new_n30238_), .Y(new_n30449_));
  OAI22X1  g28013(.A0(new_n30449_), .A1(new_n30445_), .B0(new_n30444_), .B1(new_n30249_), .Y(new_n30450_));
  AOI21X1  g28014(.A0(new_n27854_), .A1(pi0199), .B0(new_n30233_), .Y(new_n30451_));
  OAI21X1  g28015(.A0(pi0296), .A1(pi0199), .B0(new_n30451_), .Y(new_n30452_));
  OR3X1    g28016(.A(new_n6069_), .B(pi0590), .C(new_n9273_), .Y(new_n30453_));
  NAND2X1  g28017(.A(new_n30453_), .B(new_n30258_), .Y(new_n30454_));
  INVX1    g28018(.A(pi0388), .Y(new_n30455_));
  OAI21X1  g28019(.A0(pi0591), .A1(new_n30455_), .B0(pi0592), .Y(new_n30456_));
  AOI22X1  g28020(.A0(new_n30456_), .A1(new_n30454_), .B0(new_n30230_), .B1(pi0455), .Y(new_n30457_));
  OAI21X1  g28021(.A0(new_n30263_), .A1(new_n6527_), .B0(pi0588), .Y(new_n30458_));
  NAND2X1  g28022(.A(new_n30458_), .B(new_n30233_), .Y(new_n30459_));
  OAI21X1  g28023(.A0(new_n30459_), .A1(new_n30457_), .B0(new_n30452_), .Y(new_n30460_));
  MX2X1    g28024(.A(new_n30460_), .B(new_n30450_), .S0(new_n8943_), .Y(po0832));
  AOI21X1  g28025(.A0(pi1135), .A1(new_n22368_), .B0(new_n4554_), .Y(new_n30462_));
  OAI21X1  g28026(.A0(pi1135), .A1(pi0606), .B0(new_n30462_), .Y(new_n30463_));
  AOI21X1  g28027(.A0(new_n4622_), .A1(pi0812), .B0(pi1136), .Y(new_n30464_));
  OAI21X1  g28028(.A0(new_n4622_), .A1(pi0787), .B0(new_n30464_), .Y(new_n30465_));
  AOI21X1  g28029(.A0(new_n30465_), .A1(new_n30463_), .B0(new_n30239_), .Y(new_n30466_));
  AND2X1   g28030(.A(new_n30246_), .B(new_n15416_), .Y(new_n30467_));
  OAI22X1  g28031(.A0(pi1136), .A1(pi0881), .B0(new_n4622_), .B1(pi0729), .Y(new_n30468_));
  NOR3X1   g28032(.A(new_n30468_), .B(new_n30467_), .C(new_n30251_), .Y(new_n30469_));
  OAI21X1  g28033(.A0(new_n30469_), .A1(new_n30466_), .B0(new_n8943_), .Y(new_n30470_));
  NOR2X1   g28034(.A(pi0293), .B(pi0199), .Y(new_n30471_));
  OAI22X1  g28035(.A0(pi1059), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30472_));
  NOR2X1   g28036(.A(new_n30472_), .B(new_n30471_), .Y(new_n30473_));
  AOI21X1  g28037(.A0(new_n30257_), .A1(pi0410), .B0(new_n30259_), .Y(new_n30474_));
  AOI21X1  g28038(.A0(new_n6069_), .A1(pi0386), .B0(new_n6009_), .Y(new_n30475_));
  OAI22X1  g28039(.A0(new_n30475_), .A1(new_n30474_), .B0(new_n30256_), .B1(new_n6018_), .Y(new_n30476_));
  NAND3X1  g28040(.A(new_n6561_), .B(new_n6009_), .C(pi0434), .Y(new_n30477_));
  AOI21X1  g28041(.A0(new_n30477_), .A1(pi0588), .B0(new_n30234_), .Y(new_n30478_));
  AOI21X1  g28042(.A0(new_n30478_), .A1(new_n30476_), .B0(new_n30473_), .Y(new_n30479_));
  OAI21X1  g28043(.A0(new_n30479_), .A1(new_n8943_), .B0(new_n30470_), .Y(po0833));
  NOR2X1   g28044(.A(pi0259), .B(pi0199), .Y(new_n30481_));
  OAI22X1  g28045(.A0(pi1069), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30482_));
  NOR2X1   g28046(.A(new_n30482_), .B(new_n30481_), .Y(new_n30483_));
  AND3X1   g28047(.A(new_n6009_), .B(pi0591), .C(pi0335), .Y(new_n30484_));
  AOI21X1  g28048(.A0(new_n30227_), .A1(pi0366), .B0(new_n30484_), .Y(new_n30485_));
  AOI21X1  g28049(.A0(new_n30230_), .A1(pi0344), .B0(pi0588), .Y(new_n30486_));
  OAI21X1  g28050(.A0(new_n30485_), .A1(pi0590), .B0(new_n30486_), .Y(new_n30487_));
  OAI21X1  g28051(.A0(new_n30263_), .A1(new_n6504_), .B0(pi0588), .Y(new_n30488_));
  AND2X1   g28052(.A(new_n30488_), .B(new_n30233_), .Y(new_n30489_));
  AOI21X1  g28053(.A0(new_n30489_), .A1(new_n30487_), .B0(new_n30483_), .Y(new_n30490_));
  AND2X1   g28054(.A(new_n30246_), .B(pi0742), .Y(new_n30491_));
  OAI22X1  g28055(.A0(pi1136), .A1(pi0870), .B0(new_n4622_), .B1(new_n14896_), .Y(new_n30492_));
  NOR3X1   g28056(.A(new_n30492_), .B(new_n30491_), .C(new_n30251_), .Y(new_n30493_));
  NAND2X1  g28057(.A(pi1135), .B(pi0635), .Y(new_n30494_));
  AOI21X1  g28058(.A0(new_n4622_), .A1(new_n30095_), .B0(pi1134), .Y(new_n30495_));
  AND3X1   g28059(.A(new_n30495_), .B(new_n30494_), .C(new_n30359_), .Y(new_n30496_));
  OAI21X1  g28060(.A0(new_n30496_), .A1(new_n30493_), .B0(new_n8943_), .Y(new_n30497_));
  OAI21X1  g28061(.A0(new_n30490_), .A1(new_n8943_), .B0(new_n30497_), .Y(po0834));
  NOR2X1   g28062(.A(pi0260), .B(pi0199), .Y(new_n30499_));
  OAI22X1  g28063(.A0(pi1067), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30500_));
  NOR2X1   g28064(.A(new_n30500_), .B(new_n30499_), .Y(new_n30501_));
  AND3X1   g28065(.A(new_n6009_), .B(pi0591), .C(pi0393), .Y(new_n30502_));
  AOI21X1  g28066(.A0(new_n30227_), .A1(pi0368), .B0(new_n30502_), .Y(new_n30503_));
  AOI21X1  g28067(.A0(new_n30230_), .A1(pi0346), .B0(pi0588), .Y(new_n30504_));
  OAI21X1  g28068(.A0(new_n30503_), .A1(pi0590), .B0(new_n30504_), .Y(new_n30505_));
  NAND3X1  g28069(.A(new_n6561_), .B(new_n6009_), .C(pi0418), .Y(new_n30506_));
  AOI21X1  g28070(.A0(new_n30506_), .A1(pi0588), .B0(new_n30234_), .Y(new_n30507_));
  AOI21X1  g28071(.A0(new_n30507_), .A1(new_n30505_), .B0(new_n30501_), .Y(new_n30508_));
  AND2X1   g28072(.A(new_n30246_), .B(pi0760), .Y(new_n30509_));
  OAI22X1  g28073(.A0(pi1136), .A1(pi0856), .B0(new_n4622_), .B1(new_n14997_), .Y(new_n30510_));
  NOR3X1   g28074(.A(new_n30510_), .B(new_n30509_), .C(new_n30251_), .Y(new_n30511_));
  NAND2X1  g28075(.A(pi1135), .B(pi0632), .Y(new_n30512_));
  AOI21X1  g28076(.A0(new_n4622_), .A1(new_n30075_), .B0(pi1134), .Y(new_n30513_));
  AND3X1   g28077(.A(new_n30513_), .B(new_n30512_), .C(new_n30359_), .Y(new_n30514_));
  OAI21X1  g28078(.A0(new_n30514_), .A1(new_n30511_), .B0(new_n8943_), .Y(new_n30515_));
  OAI21X1  g28079(.A0(new_n30508_), .A1(new_n8943_), .B0(new_n30515_), .Y(po0835));
  NOR2X1   g28080(.A(pi0255), .B(pi0199), .Y(new_n30517_));
  OAI22X1  g28081(.A0(pi1036), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30518_));
  NOR2X1   g28082(.A(new_n30518_), .B(new_n30517_), .Y(new_n30519_));
  AND3X1   g28083(.A(new_n6009_), .B(pi0591), .C(pi0413), .Y(new_n30520_));
  AOI21X1  g28084(.A0(new_n30227_), .A1(pi0389), .B0(new_n30520_), .Y(new_n30521_));
  AOI21X1  g28085(.A0(new_n30230_), .A1(pi0450), .B0(pi0588), .Y(new_n30522_));
  OAI21X1  g28086(.A0(new_n30521_), .A1(pi0590), .B0(new_n30522_), .Y(new_n30523_));
  NAND3X1  g28087(.A(new_n6561_), .B(new_n6009_), .C(pi0438), .Y(new_n30524_));
  AOI21X1  g28088(.A0(new_n30524_), .A1(pi0588), .B0(new_n30234_), .Y(new_n30525_));
  AOI21X1  g28089(.A0(new_n30525_), .A1(new_n30523_), .B0(new_n30519_), .Y(new_n30526_));
  AOI21X1  g28090(.A0(pi1136), .A1(new_n12091_), .B0(new_n4622_), .Y(new_n30527_));
  OAI21X1  g28091(.A0(pi1136), .A1(pi0791), .B0(new_n30527_), .Y(new_n30528_));
  AOI21X1  g28092(.A0(pi1136), .A1(new_n11963_), .B0(pi1135), .Y(new_n30529_));
  OAI21X1  g28093(.A0(pi1136), .A1(pi0810), .B0(new_n30529_), .Y(new_n30530_));
  AOI21X1  g28094(.A0(new_n30530_), .A1(new_n30528_), .B0(new_n30239_), .Y(new_n30531_));
  AND2X1   g28095(.A(new_n30246_), .B(new_n15571_), .Y(new_n30532_));
  OAI22X1  g28096(.A0(pi1136), .A1(pi0874), .B0(new_n4622_), .B1(pi0690), .Y(new_n30533_));
  NOR3X1   g28097(.A(new_n30533_), .B(new_n30532_), .C(new_n30251_), .Y(new_n30534_));
  OAI21X1  g28098(.A0(new_n30534_), .A1(new_n30531_), .B0(new_n8943_), .Y(new_n30535_));
  OAI21X1  g28099(.A0(new_n30526_), .A1(new_n8943_), .B0(new_n30535_), .Y(po0836));
  OAI21X1  g28100(.A0(new_n30111_), .A1(pi1100), .B0(new_n30112_), .Y(new_n30537_));
  AOI21X1  g28101(.A0(new_n30111_), .A1(new_n5019_), .B0(new_n30537_), .Y(po0837));
  OAI21X1  g28102(.A0(new_n30111_), .A1(pi1103), .B0(new_n30112_), .Y(new_n30539_));
  AOI21X1  g28103(.A0(new_n30111_), .A1(new_n11859_), .B0(new_n30539_), .Y(po0838));
  NOR2X1   g28104(.A(pi0251), .B(pi0199), .Y(new_n30541_));
  OAI22X1  g28105(.A0(pi1039), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30542_));
  NOR2X1   g28106(.A(new_n30542_), .B(new_n30541_), .Y(new_n30543_));
  AND3X1   g28107(.A(new_n6009_), .B(pi0591), .C(pi0392), .Y(new_n30544_));
  AOI21X1  g28108(.A0(new_n30227_), .A1(pi0367), .B0(new_n30544_), .Y(new_n30545_));
  AOI21X1  g28109(.A0(new_n30230_), .A1(pi0345), .B0(pi0588), .Y(new_n30546_));
  OAI21X1  g28110(.A0(new_n30545_), .A1(pi0590), .B0(new_n30546_), .Y(new_n30547_));
  NAND3X1  g28111(.A(new_n6561_), .B(new_n6009_), .C(pi0417), .Y(new_n30548_));
  AOI21X1  g28112(.A0(new_n30548_), .A1(pi0588), .B0(new_n30234_), .Y(new_n30549_));
  AOI21X1  g28113(.A0(new_n30549_), .A1(new_n30547_), .B0(new_n30543_), .Y(new_n30550_));
  AND2X1   g28114(.A(new_n30246_), .B(pi0757), .Y(new_n30551_));
  OAI22X1  g28115(.A0(pi1136), .A1(pi0848), .B0(new_n4622_), .B1(new_n14935_), .Y(new_n30552_));
  NOR3X1   g28116(.A(new_n30552_), .B(new_n30551_), .C(new_n30251_), .Y(new_n30553_));
  NAND2X1  g28117(.A(pi1135), .B(pi0631), .Y(new_n30554_));
  AOI21X1  g28118(.A0(new_n4622_), .A1(new_n30067_), .B0(pi1134), .Y(new_n30555_));
  AND3X1   g28119(.A(new_n30555_), .B(new_n30554_), .C(new_n30359_), .Y(new_n30556_));
  OAI21X1  g28120(.A0(new_n30556_), .A1(new_n30553_), .B0(new_n8943_), .Y(new_n30557_));
  OAI21X1  g28121(.A0(new_n30550_), .A1(new_n8943_), .B0(new_n30557_), .Y(po0839));
  INVX1    g28122(.A(pi0953), .Y(new_n30559_));
  NOR4X1   g28123(.A(new_n30109_), .B(pi0973), .C(new_n30559_), .D(new_n12767_), .Y(po0980));
  INVX1    g28124(.A(pi0684), .Y(new_n30561_));
  OAI21X1  g28125(.A0(po0980), .A1(new_n30561_), .B0(new_n30112_), .Y(new_n30562_));
  AOI21X1  g28126(.A0(po0980), .A1(new_n30183_), .B0(new_n30562_), .Y(po0841));
  INVX1    g28127(.A(new_n27852_), .Y(new_n30564_));
  AND2X1   g28128(.A(pi0592), .B(new_n6334_), .Y(new_n30565_));
  AND2X1   g28129(.A(new_n6009_), .B(pi0590), .Y(new_n30566_));
  AOI22X1  g28130(.A0(new_n30566_), .A1(pi0357), .B0(new_n30565_), .B1(pi0382), .Y(new_n30567_));
  OR4X1    g28131(.A(pi0592), .B(new_n6069_), .C(pi0590), .D(new_n6195_), .Y(new_n30568_));
  OAI21X1  g28132(.A0(new_n30567_), .A1(pi0591), .B0(new_n30568_), .Y(new_n30569_));
  OR2X1    g28133(.A(pi0590), .B(new_n6603_), .Y(new_n30570_));
  NOR4X1   g28134(.A(new_n30570_), .B(pi0592), .C(pi0591), .D(new_n6550_), .Y(new_n30571_));
  AOI21X1  g28135(.A0(new_n30569_), .A1(new_n6603_), .B0(new_n30571_), .Y(new_n30572_));
  OAI22X1  g28136(.A0(pi1076), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30573_));
  OAI22X1  g28137(.A0(new_n30573_), .A1(new_n30564_), .B0(new_n30572_), .B1(new_n30234_), .Y(new_n30574_));
  NAND2X1  g28138(.A(new_n4622_), .B(pi0744), .Y(new_n30575_));
  AOI21X1  g28139(.A0(pi1135), .A1(pi0728), .B0(new_n4554_), .Y(new_n30576_));
  AOI22X1  g28140(.A0(new_n30576_), .A1(new_n30575_), .B0(new_n30278_), .B1(pi0860), .Y(new_n30577_));
  OAI21X1  g28141(.A0(new_n30245_), .A1(new_n4554_), .B0(new_n4747_), .Y(new_n30578_));
  OR2X1    g28142(.A(pi1135), .B(pi0652), .Y(new_n30579_));
  AOI21X1  g28143(.A0(pi1135), .A1(pi0657), .B0(new_n4554_), .Y(new_n30580_));
  AND3X1   g28144(.A(new_n30278_), .B(new_n30245_), .C(pi0813), .Y(new_n30581_));
  AOI21X1  g28145(.A0(new_n30580_), .A1(new_n30579_), .B0(new_n30581_), .Y(new_n30582_));
  OAI22X1  g28146(.A0(new_n30582_), .A1(new_n30578_), .B0(new_n30577_), .B1(new_n30249_), .Y(new_n30583_));
  MX2X1    g28147(.A(new_n30583_), .B(new_n30574_), .S0(new_n6713_), .Y(po0842));
  OAI21X1  g28148(.A0(po0980), .A1(new_n14935_), .B0(new_n30112_), .Y(new_n30585_));
  AOI21X1  g28149(.A0(po0980), .A1(new_n30125_), .B0(new_n30585_), .Y(po0843));
  INVX1    g28150(.A(po0980), .Y(new_n30587_));
  OAI21X1  g28151(.A0(new_n30587_), .A1(pi1127), .B0(new_n30112_), .Y(new_n30588_));
  AOI21X1  g28152(.A0(new_n30587_), .A1(new_n13538_), .B0(new_n30588_), .Y(po0844));
  OAI21X1  g28153(.A0(po0980), .A1(new_n14997_), .B0(new_n30112_), .Y(new_n30590_));
  AOI21X1  g28154(.A0(po0980), .A1(new_n30129_), .B0(new_n30590_), .Y(po0845));
  AOI22X1  g28155(.A0(new_n30566_), .A1(pi0351), .B0(new_n30565_), .B1(pi0376), .Y(new_n30592_));
  NAND4X1  g28156(.A(new_n6009_), .B(pi0591), .C(new_n6334_), .D(pi0401), .Y(new_n30593_));
  OAI21X1  g28157(.A0(new_n30592_), .A1(pi0591), .B0(new_n30593_), .Y(new_n30594_));
  NOR4X1   g28158(.A(new_n30570_), .B(pi0592), .C(pi0591), .D(new_n6553_), .Y(new_n30595_));
  AOI21X1  g28159(.A0(new_n30594_), .A1(new_n6603_), .B0(new_n30595_), .Y(new_n30596_));
  NOR2X1   g28160(.A(new_n27840_), .B(pi0199), .Y(new_n30597_));
  OAI22X1  g28161(.A0(pi1079), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30598_));
  OAI22X1  g28162(.A0(new_n30598_), .A1(new_n30597_), .B0(new_n30596_), .B1(new_n30234_), .Y(new_n30599_));
  OR2X1    g28163(.A(pi1135), .B(pi0658), .Y(new_n30600_));
  AOI21X1  g28164(.A0(pi1135), .A1(pi0655), .B0(new_n4554_), .Y(new_n30601_));
  AOI22X1  g28165(.A0(new_n30601_), .A1(new_n30600_), .B0(new_n30278_), .B1(pi0798), .Y(new_n30602_));
  AND2X1   g28166(.A(new_n30246_), .B(pi0752), .Y(new_n30603_));
  OAI22X1  g28167(.A0(pi1136), .A1(pi0843), .B0(new_n4622_), .B1(pi0703), .Y(new_n30604_));
  OR3X1    g28168(.A(new_n30604_), .B(new_n30603_), .C(new_n30251_), .Y(new_n30605_));
  OAI21X1  g28169(.A0(new_n30602_), .A1(new_n30239_), .B0(new_n30605_), .Y(new_n30606_));
  MX2X1    g28170(.A(new_n30606_), .B(new_n30599_), .S0(new_n6713_), .Y(po0846));
  OAI21X1  g28171(.A0(new_n30587_), .A1(pi1108), .B0(new_n30112_), .Y(new_n30608_));
  AOI21X1  g28172(.A0(new_n30587_), .A1(new_n15565_), .B0(new_n30608_), .Y(po0847));
  OAI21X1  g28173(.A0(new_n30587_), .A1(pi1107), .B0(new_n30112_), .Y(new_n30610_));
  AOI21X1  g28174(.A0(new_n30587_), .A1(new_n15513_), .B0(new_n30610_), .Y(po0848));
  AND3X1   g28175(.A(new_n6009_), .B(pi0590), .C(pi0352), .Y(new_n30612_));
  AND3X1   g28176(.A(pi0592), .B(new_n6334_), .C(pi0317), .Y(new_n30613_));
  OAI21X1  g28177(.A0(new_n30613_), .A1(new_n30612_), .B0(new_n6069_), .Y(new_n30614_));
  NAND4X1  g28178(.A(new_n6009_), .B(pi0591), .C(new_n6334_), .D(pi0402), .Y(new_n30615_));
  AOI21X1  g28179(.A0(new_n30615_), .A1(new_n30614_), .B0(pi0588), .Y(new_n30616_));
  NOR4X1   g28180(.A(new_n30570_), .B(pi0592), .C(pi0591), .D(new_n6496_), .Y(new_n30617_));
  OAI21X1  g28181(.A0(new_n30617_), .A1(new_n30616_), .B0(new_n30233_), .Y(new_n30618_));
  NOR2X1   g28182(.A(new_n27844_), .B(pi0199), .Y(new_n30619_));
  OAI22X1  g28183(.A0(pi1078), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30620_));
  OR2X1    g28184(.A(new_n30620_), .B(new_n30619_), .Y(new_n30621_));
  AOI21X1  g28185(.A0(new_n30621_), .A1(new_n30618_), .B0(new_n8943_), .Y(new_n30622_));
  INVX1    g28186(.A(new_n30281_), .Y(new_n30623_));
  AOI21X1  g28187(.A0(new_n4622_), .A1(pi0770), .B0(new_n4554_), .Y(new_n30624_));
  OAI21X1  g28188(.A0(new_n4622_), .A1(pi0726), .B0(new_n30624_), .Y(new_n30625_));
  AOI21X1  g28189(.A0(new_n30278_), .A1(pi0844), .B0(new_n4747_), .Y(new_n30626_));
  AND2X1   g28190(.A(new_n30626_), .B(new_n30625_), .Y(new_n30627_));
  OR2X1    g28191(.A(pi1135), .B(pi0656), .Y(new_n30628_));
  AOI21X1  g28192(.A0(pi1135), .A1(pi0649), .B0(new_n4554_), .Y(new_n30629_));
  INVX1    g28193(.A(pi0801), .Y(new_n30630_));
  OAI21X1  g28194(.A0(new_n30279_), .A1(new_n30630_), .B0(new_n4747_), .Y(new_n30631_));
  AOI21X1  g28195(.A0(new_n30629_), .A1(new_n30628_), .B0(new_n30631_), .Y(new_n30632_));
  NOR3X1   g28196(.A(new_n30632_), .B(new_n30627_), .C(new_n30623_), .Y(new_n30633_));
  OR2X1    g28197(.A(new_n30633_), .B(new_n30622_), .Y(po0849));
  INVX1    g28198(.A(pi0693), .Y(new_n30635_));
  OAI21X1  g28199(.A0(po0954), .A1(new_n30635_), .B0(new_n30112_), .Y(new_n30636_));
  AOI21X1  g28200(.A0(po0954), .A1(new_n30191_), .B0(new_n30636_), .Y(po0850));
  INVX1    g28201(.A(pi0694), .Y(new_n30638_));
  OAI21X1  g28202(.A0(po0980), .A1(new_n30638_), .B0(new_n30112_), .Y(new_n30639_));
  AOI21X1  g28203(.A0(po0980), .A1(new_n30152_), .B0(new_n30639_), .Y(po0851));
  INVX1    g28204(.A(pi1111), .Y(new_n30641_));
  OAI21X1  g28205(.A0(po0954), .A1(new_n23366_), .B0(new_n30112_), .Y(new_n30642_));
  AOI21X1  g28206(.A0(po0954), .A1(new_n30641_), .B0(new_n30642_), .Y(po0852));
  OAI21X1  g28207(.A0(new_n30587_), .A1(pi1100), .B0(new_n30112_), .Y(new_n30644_));
  AOI21X1  g28208(.A0(new_n30587_), .A1(new_n14807_), .B0(new_n30644_), .Y(po0853));
  INVX1    g28209(.A(pi0697), .Y(new_n30646_));
  OAI21X1  g28210(.A0(po0980), .A1(new_n30646_), .B0(new_n30112_), .Y(new_n30647_));
  AOI21X1  g28211(.A0(po0980), .A1(new_n30191_), .B0(new_n30647_), .Y(po0854));
  INVX1    g28212(.A(pi1116), .Y(new_n30649_));
  OAI21X1  g28213(.A0(po0980), .A1(new_n14359_), .B0(new_n30112_), .Y(new_n30650_));
  AOI21X1  g28214(.A0(po0980), .A1(new_n30649_), .B0(new_n30650_), .Y(po0855));
  OAI21X1  g28215(.A0(new_n30587_), .A1(pi1103), .B0(new_n30112_), .Y(new_n30652_));
  AOI21X1  g28216(.A0(new_n30587_), .A1(new_n15361_), .B0(new_n30652_), .Y(po0856));
  OAI21X1  g28217(.A0(new_n30587_), .A1(pi1110), .B0(new_n30112_), .Y(new_n30654_));
  AOI21X1  g28218(.A0(new_n30587_), .A1(new_n14840_), .B0(new_n30654_), .Y(po0857));
  INVX1    g28219(.A(pi1123), .Y(new_n30656_));
  OAI21X1  g28220(.A0(po0980), .A1(new_n14697_), .B0(new_n30112_), .Y(new_n30657_));
  AOI21X1  g28221(.A0(po0980), .A1(new_n30656_), .B0(new_n30657_), .Y(po0858));
  INVX1    g28222(.A(pi1117), .Y(new_n30659_));
  OAI21X1  g28223(.A0(po0980), .A1(new_n15025_), .B0(new_n30112_), .Y(new_n30660_));
  AOI21X1  g28224(.A0(po0980), .A1(new_n30659_), .B0(new_n30660_), .Y(po0859));
  OAI21X1  g28225(.A0(new_n30587_), .A1(pi1124), .B0(new_n30112_), .Y(new_n30662_));
  AOI21X1  g28226(.A0(new_n30587_), .A1(new_n15229_), .B0(new_n30662_), .Y(po0860));
  OAI21X1  g28227(.A0(po0980), .A1(new_n14896_), .B0(new_n30112_), .Y(new_n30664_));
  AOI21X1  g28228(.A0(po0980), .A1(new_n30137_), .B0(new_n30664_), .Y(po0861));
  OAI21X1  g28229(.A0(new_n30587_), .A1(pi1125), .B0(new_n30112_), .Y(new_n30666_));
  AOI21X1  g28230(.A0(new_n30587_), .A1(new_n15335_), .B0(new_n30666_), .Y(po0862));
  OAI21X1  g28231(.A0(new_n30587_), .A1(pi1105), .B0(new_n30112_), .Y(new_n30668_));
  AOI21X1  g28232(.A0(new_n30587_), .A1(new_n12805_), .B0(new_n30668_), .Y(po0863));
  INVX1    g28233(.A(new_n30227_), .Y(new_n30670_));
  OR3X1    g28234(.A(pi0592), .B(new_n6069_), .C(new_n6167_), .Y(new_n30671_));
  OAI21X1  g28235(.A0(new_n30670_), .A1(new_n6077_), .B0(new_n30671_), .Y(new_n30672_));
  AOI22X1  g28236(.A0(new_n30672_), .A1(new_n6334_), .B0(new_n30230_), .B1(pi0347), .Y(new_n30673_));
  NOR3X1   g28237(.A(pi0588), .B(pi0224), .C(pi0223), .Y(new_n30674_));
  INVX1    g28238(.A(new_n30674_), .Y(new_n30675_));
  MX2X1    g28239(.A(pi0304), .B(pi1048), .S0(pi0200), .Y(new_n30676_));
  OR2X1    g28240(.A(new_n30676_), .B(pi0199), .Y(new_n30677_));
  INVX1    g28241(.A(pi1055), .Y(new_n30678_));
  AOI21X1  g28242(.A0(new_n30678_), .A1(pi0199), .B0(new_n30233_), .Y(new_n30679_));
  NAND2X1  g28243(.A(pi0588), .B(pi0420), .Y(new_n30680_));
  NOR4X1   g28244(.A(new_n30680_), .B(new_n30263_), .C(pi0224), .D(pi0223), .Y(new_n30681_));
  AOI21X1  g28245(.A0(new_n30679_), .A1(new_n30677_), .B0(new_n30681_), .Y(new_n30682_));
  OAI21X1  g28246(.A0(new_n30675_), .A1(new_n30673_), .B0(new_n30682_), .Y(new_n30683_));
  INVX1    g28247(.A(new_n30359_), .Y(new_n30684_));
  AOI21X1  g28248(.A0(new_n4622_), .A1(new_n12486_), .B0(pi1134), .Y(new_n30685_));
  OAI21X1  g28249(.A0(new_n4622_), .A1(pi0627), .B0(new_n30685_), .Y(new_n30686_));
  AND2X1   g28250(.A(new_n30246_), .B(pi0753), .Y(new_n30687_));
  OAI22X1  g28251(.A0(pi1136), .A1(pi0847), .B0(new_n4622_), .B1(new_n15025_), .Y(new_n30688_));
  OR3X1    g28252(.A(new_n30688_), .B(new_n30687_), .C(new_n30251_), .Y(new_n30689_));
  OAI21X1  g28253(.A0(new_n30686_), .A1(new_n30684_), .B0(new_n30689_), .Y(new_n30690_));
  MX2X1    g28254(.A(new_n30690_), .B(new_n30683_), .S0(new_n6713_), .Y(po0864));
  NAND4X1  g28255(.A(new_n30233_), .B(pi0592), .C(new_n6069_), .D(pi0442), .Y(new_n30692_));
  NAND4X1  g28256(.A(new_n30233_), .B(new_n6009_), .C(pi0591), .D(pi0328), .Y(new_n30693_));
  AOI21X1  g28257(.A0(new_n30693_), .A1(new_n30692_), .B0(pi0590), .Y(new_n30694_));
  AND3X1   g28258(.A(new_n30230_), .B(new_n30233_), .C(pi0321), .Y(new_n30695_));
  OAI21X1  g28259(.A0(new_n30695_), .A1(new_n30694_), .B0(new_n6603_), .Y(new_n30696_));
  MX2X1    g28260(.A(pi0305), .B(pi1084), .S0(pi0200), .Y(new_n30697_));
  NOR2X1   g28261(.A(new_n30697_), .B(pi0199), .Y(new_n30698_));
  OAI22X1  g28262(.A0(pi1058), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30699_));
  OR2X1    g28263(.A(new_n30699_), .B(new_n30698_), .Y(new_n30700_));
  INVX1    g28264(.A(pi0459), .Y(new_n30701_));
  OR4X1    g28265(.A(pi0592), .B(pi0591), .C(pi0224), .D(pi0223), .Y(new_n30702_));
  OR4X1    g28266(.A(new_n30702_), .B(pi0590), .C(new_n6603_), .D(new_n30701_), .Y(new_n30703_));
  AND3X1   g28267(.A(new_n30703_), .B(new_n30700_), .C(new_n6713_), .Y(new_n30704_));
  NAND2X1  g28268(.A(new_n30246_), .B(pi0754), .Y(new_n30705_));
  OR2X1    g28269(.A(pi1136), .B(new_n4622_), .Y(new_n30706_));
  AND2X1   g28270(.A(new_n30706_), .B(new_n30245_), .Y(new_n30707_));
  OAI21X1  g28271(.A0(pi1136), .A1(pi0857), .B0(pi1134), .Y(new_n30708_));
  AOI21X1  g28272(.A0(pi1135), .A1(pi0709), .B0(new_n30708_), .Y(new_n30709_));
  NAND3X1  g28273(.A(new_n30709_), .B(new_n30707_), .C(new_n30705_), .Y(new_n30710_));
  OAI21X1  g28274(.A0(new_n4622_), .A1(pi0660), .B0(new_n4747_), .Y(new_n30711_));
  AOI21X1  g28275(.A0(new_n4622_), .A1(new_n12462_), .B0(new_n30711_), .Y(new_n30712_));
  AOI21X1  g28276(.A0(new_n30712_), .A1(new_n30359_), .B0(new_n6713_), .Y(new_n30713_));
  AOI22X1  g28277(.A0(new_n30713_), .A1(new_n30710_), .B0(new_n30704_), .B1(new_n30696_), .Y(po0865));
  INVX1    g28278(.A(pi1118), .Y(new_n30715_));
  OAI21X1  g28279(.A0(po0980), .A1(new_n15056_), .B0(new_n30112_), .Y(new_n30716_));
  AOI21X1  g28280(.A0(po0980), .A1(new_n30715_), .B0(new_n30716_), .Y(po0866));
  OAI21X1  g28281(.A0(new_n30111_), .A1(pi1106), .B0(new_n30112_), .Y(new_n30718_));
  AOI21X1  g28282(.A0(new_n30111_), .A1(new_n22697_), .B0(new_n30718_), .Y(po0867));
  NAND3X1  g28283(.A(new_n6009_), .B(pi0591), .C(pi0398), .Y(new_n30720_));
  OAI21X1  g28284(.A0(new_n30670_), .A1(new_n6075_), .B0(new_n30720_), .Y(new_n30721_));
  AOI22X1  g28285(.A0(new_n30721_), .A1(new_n6334_), .B0(new_n30230_), .B1(pi0348), .Y(new_n30722_));
  MX2X1    g28286(.A(pi0306), .B(pi1059), .S0(pi0200), .Y(new_n30723_));
  OR2X1    g28287(.A(new_n30723_), .B(pi0199), .Y(new_n30724_));
  INVX1    g28288(.A(pi1087), .Y(new_n30725_));
  AOI21X1  g28289(.A0(new_n30725_), .A1(pi0199), .B0(new_n30233_), .Y(new_n30726_));
  NAND2X1  g28290(.A(pi0588), .B(pi0423), .Y(new_n30727_));
  NOR4X1   g28291(.A(new_n30727_), .B(new_n30263_), .C(pi0224), .D(pi0223), .Y(new_n30728_));
  AOI21X1  g28292(.A0(new_n30726_), .A1(new_n30724_), .B0(new_n30728_), .Y(new_n30729_));
  OAI21X1  g28293(.A0(new_n30722_), .A1(new_n30675_), .B0(new_n30729_), .Y(new_n30730_));
  AOI21X1  g28294(.A0(new_n4622_), .A1(new_n12592_), .B0(pi1134), .Y(new_n30731_));
  OAI21X1  g28295(.A0(new_n4622_), .A1(pi0647), .B0(new_n30731_), .Y(new_n30732_));
  AND2X1   g28296(.A(new_n30246_), .B(pi0755), .Y(new_n30733_));
  OAI22X1  g28297(.A0(pi1136), .A1(pi0858), .B0(new_n4622_), .B1(new_n14667_), .Y(new_n30734_));
  OR3X1    g28298(.A(new_n30734_), .B(new_n30733_), .C(new_n30251_), .Y(new_n30735_));
  OAI21X1  g28299(.A0(new_n30732_), .A1(new_n30684_), .B0(new_n30735_), .Y(new_n30736_));
  MX2X1    g28300(.A(new_n30736_), .B(new_n30730_), .S0(new_n6713_), .Y(po0868));
  NAND2X1  g28301(.A(new_n30246_), .B(pi0751), .Y(new_n30738_));
  OAI21X1  g28302(.A0(pi1136), .A1(pi0842), .B0(pi1134), .Y(new_n30739_));
  AOI21X1  g28303(.A0(pi1135), .A1(pi0701), .B0(new_n30739_), .Y(new_n30740_));
  AND3X1   g28304(.A(new_n30740_), .B(new_n30706_), .C(new_n30245_), .Y(new_n30741_));
  OAI21X1  g28305(.A0(pi1135), .A1(pi0644), .B0(new_n4747_), .Y(new_n30742_));
  AOI21X1  g28306(.A0(pi1135), .A1(new_n12608_), .B0(new_n30742_), .Y(new_n30743_));
  AOI22X1  g28307(.A0(new_n30743_), .A1(new_n30359_), .B0(new_n30741_), .B1(new_n30738_), .Y(new_n30744_));
  AND3X1   g28308(.A(new_n6009_), .B(pi0591), .C(pi0400), .Y(new_n30745_));
  AOI21X1  g28309(.A0(new_n30227_), .A1(pi0374), .B0(new_n30745_), .Y(new_n30746_));
  OAI22X1  g28310(.A0(new_n30746_), .A1(pi0590), .B0(new_n30256_), .B1(new_n6007_), .Y(new_n30747_));
  OR2X1    g28311(.A(pi0592), .B(pi0591), .Y(new_n30748_));
  NAND3X1  g28312(.A(new_n6334_), .B(pi0588), .C(pi0425), .Y(new_n30749_));
  OAI21X1  g28313(.A0(new_n30749_), .A1(new_n30748_), .B0(new_n30233_), .Y(new_n30750_));
  AOI21X1  g28314(.A0(new_n30747_), .A1(new_n6603_), .B0(new_n30750_), .Y(new_n30751_));
  AND2X1   g28315(.A(new_n8055_), .B(pi0298), .Y(new_n30752_));
  OR3X1    g28316(.A(new_n27850_), .B(new_n7937_), .C(pi0199), .Y(new_n30753_));
  AOI21X1  g28317(.A0(pi1035), .A1(pi0199), .B0(new_n30233_), .Y(new_n30754_));
  NAND2X1  g28318(.A(new_n30754_), .B(new_n30753_), .Y(new_n30755_));
  OAI21X1  g28319(.A0(new_n30755_), .A1(new_n30752_), .B0(new_n6713_), .Y(new_n30756_));
  OAI22X1  g28320(.A0(new_n30756_), .A1(new_n30751_), .B0(new_n30744_), .B1(new_n6713_), .Y(po0869));
  NAND3X1  g28321(.A(new_n6009_), .B(pi0591), .C(pi0396), .Y(new_n30758_));
  OAI21X1  g28322(.A0(new_n30670_), .A1(new_n6076_), .B0(new_n30758_), .Y(new_n30759_));
  AOI22X1  g28323(.A0(new_n30759_), .A1(new_n6334_), .B0(new_n30230_), .B1(pi0322), .Y(new_n30760_));
  MX2X1    g28324(.A(pi0309), .B(pi1072), .S0(pi0200), .Y(new_n30761_));
  OR2X1    g28325(.A(new_n30761_), .B(pi0199), .Y(new_n30762_));
  INVX1    g28326(.A(pi1051), .Y(new_n30763_));
  AOI21X1  g28327(.A0(new_n30763_), .A1(pi0199), .B0(new_n30233_), .Y(new_n30764_));
  NAND2X1  g28328(.A(pi0588), .B(pi0421), .Y(new_n30765_));
  NOR4X1   g28329(.A(new_n30765_), .B(new_n30263_), .C(pi0224), .D(pi0223), .Y(new_n30766_));
  AOI21X1  g28330(.A0(new_n30764_), .A1(new_n30762_), .B0(new_n30766_), .Y(new_n30767_));
  OAI21X1  g28331(.A0(new_n30760_), .A1(new_n30675_), .B0(new_n30767_), .Y(new_n30768_));
  AOI21X1  g28332(.A0(new_n4622_), .A1(new_n12561_), .B0(pi1134), .Y(new_n30769_));
  OAI21X1  g28333(.A0(new_n4622_), .A1(pi0628), .B0(new_n30769_), .Y(new_n30770_));
  AND2X1   g28334(.A(new_n30246_), .B(pi0756), .Y(new_n30771_));
  OAI22X1  g28335(.A0(pi1136), .A1(pi0854), .B0(new_n4622_), .B1(new_n15095_), .Y(new_n30772_));
  OR3X1    g28336(.A(new_n30772_), .B(new_n30771_), .C(new_n30251_), .Y(new_n30773_));
  OAI21X1  g28337(.A0(new_n30770_), .A1(new_n30684_), .B0(new_n30773_), .Y(new_n30774_));
  MX2X1    g28338(.A(new_n30774_), .B(new_n30768_), .S0(new_n6713_), .Y(po0870));
  AOI22X1  g28339(.A0(new_n30566_), .A1(pi0461), .B0(new_n30565_), .B1(pi0439), .Y(new_n30776_));
  NAND4X1  g28340(.A(new_n6009_), .B(pi0591), .C(new_n6334_), .D(pi0326), .Y(new_n30777_));
  OAI21X1  g28341(.A0(new_n30776_), .A1(pi0591), .B0(new_n30777_), .Y(new_n30778_));
  NOR4X1   g28342(.A(new_n30748_), .B(pi0590), .C(new_n6603_), .D(new_n6492_), .Y(new_n30779_));
  AOI21X1  g28343(.A0(new_n30778_), .A1(new_n6603_), .B0(new_n30779_), .Y(new_n30780_));
  OAI22X1  g28344(.A0(pi1057), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30781_));
  OAI22X1  g28345(.A0(new_n30781_), .A1(new_n27490_), .B0(new_n30780_), .B1(new_n30234_), .Y(new_n30782_));
  NAND2X1  g28346(.A(new_n4622_), .B(pi0762), .Y(new_n30783_));
  AOI21X1  g28347(.A0(pi1135), .A1(pi0697), .B0(new_n4554_), .Y(new_n30784_));
  AOI22X1  g28348(.A0(new_n30784_), .A1(new_n30783_), .B0(new_n30278_), .B1(pi0867), .Y(new_n30785_));
  OR2X1    g28349(.A(pi1135), .B(pi0653), .Y(new_n30786_));
  AOI21X1  g28350(.A0(pi1135), .A1(pi0693), .B0(new_n4554_), .Y(new_n30787_));
  AND3X1   g28351(.A(new_n30278_), .B(new_n30245_), .C(pi0816), .Y(new_n30788_));
  AOI21X1  g28352(.A0(new_n30787_), .A1(new_n30786_), .B0(new_n30788_), .Y(new_n30789_));
  OAI22X1  g28353(.A0(new_n30789_), .A1(new_n30578_), .B0(new_n30785_), .B1(new_n30249_), .Y(new_n30790_));
  MX2X1    g28354(.A(new_n30790_), .B(new_n30782_), .S0(new_n6713_), .Y(po0871));
  OAI21X1  g28355(.A0(new_n30111_), .A1(pi1123), .B0(new_n30112_), .Y(new_n30792_));
  AOI21X1  g28356(.A0(new_n30111_), .A1(new_n12608_), .B0(new_n30792_), .Y(po0872));
  NAND4X1  g28357(.A(new_n30233_), .B(pi0592), .C(new_n6069_), .D(pi0440), .Y(new_n30794_));
  NAND4X1  g28358(.A(new_n30233_), .B(new_n6009_), .C(pi0591), .D(pi0329), .Y(new_n30795_));
  AOI21X1  g28359(.A0(new_n30795_), .A1(new_n30794_), .B0(pi0590), .Y(new_n30796_));
  AND3X1   g28360(.A(new_n30230_), .B(new_n30233_), .C(pi0349), .Y(new_n30797_));
  OAI21X1  g28361(.A0(new_n30797_), .A1(new_n30796_), .B0(new_n6603_), .Y(new_n30798_));
  MX2X1    g28362(.A(pi0307), .B(pi1053), .S0(pi0200), .Y(new_n30799_));
  NOR2X1   g28363(.A(new_n30799_), .B(pi0199), .Y(new_n30800_));
  OAI22X1  g28364(.A0(pi1043), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30801_));
  OR2X1    g28365(.A(new_n30801_), .B(new_n30800_), .Y(new_n30802_));
  INVX1    g28366(.A(pi0454), .Y(new_n30803_));
  OR4X1    g28367(.A(new_n30702_), .B(pi0590), .C(new_n6603_), .D(new_n30803_), .Y(new_n30804_));
  AND3X1   g28368(.A(new_n30804_), .B(new_n30802_), .C(new_n6713_), .Y(new_n30805_));
  NAND2X1  g28369(.A(new_n30246_), .B(pi0761), .Y(new_n30806_));
  OAI21X1  g28370(.A0(pi1136), .A1(pi0845), .B0(pi1134), .Y(new_n30807_));
  AOI21X1  g28371(.A0(pi1135), .A1(pi0738), .B0(new_n30807_), .Y(new_n30808_));
  NAND3X1  g28372(.A(new_n30808_), .B(new_n30806_), .C(new_n30707_), .Y(new_n30809_));
  OAI21X1  g28373(.A0(new_n4622_), .A1(pi0641), .B0(new_n4747_), .Y(new_n30810_));
  AOI21X1  g28374(.A0(new_n4622_), .A1(new_n12542_), .B0(new_n30810_), .Y(new_n30811_));
  AOI21X1  g28375(.A0(new_n30811_), .A1(new_n30359_), .B0(new_n6713_), .Y(new_n30812_));
  AOI22X1  g28376(.A0(new_n30812_), .A1(new_n30809_), .B0(new_n30805_), .B1(new_n30798_), .Y(po0873));
  NAND2X1  g28377(.A(pi0591), .B(pi0318), .Y(new_n30814_));
  NAND2X1  g28378(.A(new_n6101_), .B(new_n6069_), .Y(new_n30815_));
  OAI21X1  g28379(.A0(new_n30814_), .A1(pi0592), .B0(new_n30815_), .Y(new_n30816_));
  AOI22X1  g28380(.A0(new_n30816_), .A1(new_n6334_), .B0(new_n30230_), .B1(pi0462), .Y(new_n30817_));
  OR2X1    g28381(.A(new_n27842_), .B(pi0199), .Y(new_n30818_));
  INVX1    g28382(.A(pi1074), .Y(new_n30819_));
  AOI21X1  g28383(.A0(new_n30819_), .A1(pi0199), .B0(new_n30233_), .Y(new_n30820_));
  NOR4X1   g28384(.A(new_n30263_), .B(new_n30234_), .C(new_n6603_), .D(new_n6491_), .Y(new_n30821_));
  AOI21X1  g28385(.A0(new_n30820_), .A1(new_n30818_), .B0(new_n30821_), .Y(new_n30822_));
  OAI21X1  g28386(.A0(new_n30817_), .A1(new_n30675_), .B0(new_n30822_), .Y(new_n30823_));
  AND2X1   g28387(.A(new_n30246_), .B(pi0768), .Y(new_n30824_));
  OAI21X1  g28388(.A0(pi1136), .A1(pi0839), .B0(pi1134), .Y(new_n30825_));
  AOI21X1  g28389(.A0(pi1135), .A1(new_n15335_), .B0(new_n30825_), .Y(new_n30826_));
  NAND3X1  g28390(.A(new_n30826_), .B(new_n30706_), .C(new_n30245_), .Y(new_n30827_));
  OR2X1    g28391(.A(pi1135), .B(pi0645), .Y(new_n30828_));
  AOI21X1  g28392(.A0(pi1135), .A1(pi0669), .B0(new_n4554_), .Y(new_n30829_));
  AOI22X1  g28393(.A0(new_n30829_), .A1(new_n30828_), .B0(new_n30278_), .B1(pi0800), .Y(new_n30830_));
  OAI22X1  g28394(.A0(new_n30830_), .A1(new_n30239_), .B0(new_n30827_), .B1(new_n30824_), .Y(new_n30831_));
  MX2X1    g28395(.A(new_n30831_), .B(new_n30823_), .S0(new_n6713_), .Y(po0874));
  NAND4X1  g28396(.A(new_n30233_), .B(pi0592), .C(new_n6069_), .D(pi0369), .Y(new_n30833_));
  NAND4X1  g28397(.A(new_n30233_), .B(new_n6009_), .C(pi0591), .D(pi0394), .Y(new_n30834_));
  AOI21X1  g28398(.A0(new_n30834_), .A1(new_n30833_), .B0(pi0590), .Y(new_n30835_));
  AND3X1   g28399(.A(new_n30230_), .B(new_n30233_), .C(pi0315), .Y(new_n30836_));
  OAI21X1  g28400(.A0(new_n30836_), .A1(new_n30835_), .B0(new_n6603_), .Y(new_n30837_));
  MX2X1    g28401(.A(pi0303), .B(pi1049), .S0(pi0200), .Y(new_n30838_));
  NOR2X1   g28402(.A(new_n30838_), .B(pi0199), .Y(new_n30839_));
  OAI22X1  g28403(.A0(pi1080), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30840_));
  OR2X1    g28404(.A(new_n30840_), .B(new_n30839_), .Y(new_n30841_));
  INVX1    g28405(.A(pi0419), .Y(new_n30842_));
  OR4X1    g28406(.A(new_n30702_), .B(pi0590), .C(new_n6603_), .D(new_n30842_), .Y(new_n30843_));
  AND3X1   g28407(.A(new_n30843_), .B(new_n30841_), .C(new_n6713_), .Y(new_n30844_));
  NAND2X1  g28408(.A(new_n30246_), .B(pi0767), .Y(new_n30845_));
  OAI21X1  g28409(.A0(pi1136), .A1(pi0853), .B0(pi1134), .Y(new_n30846_));
  AOI21X1  g28410(.A0(pi1135), .A1(pi0698), .B0(new_n30846_), .Y(new_n30847_));
  NAND3X1  g28411(.A(new_n30847_), .B(new_n30845_), .C(new_n30707_), .Y(new_n30848_));
  OAI21X1  g28412(.A0(new_n4622_), .A1(pi0625), .B0(new_n4747_), .Y(new_n30849_));
  AOI21X1  g28413(.A0(new_n4622_), .A1(new_n12368_), .B0(new_n30849_), .Y(new_n30850_));
  AOI21X1  g28414(.A0(new_n30850_), .A1(new_n30359_), .B0(new_n6713_), .Y(new_n30851_));
  AOI22X1  g28415(.A0(new_n30851_), .A1(new_n30848_), .B0(new_n30844_), .B1(new_n30837_), .Y(po0875));
  NAND3X1  g28416(.A(new_n6009_), .B(pi0591), .C(pi0325), .Y(new_n30853_));
  OAI21X1  g28417(.A0(new_n30670_), .A1(new_n6105_), .B0(new_n30853_), .Y(new_n30854_));
  AOI22X1  g28418(.A0(new_n30854_), .A1(new_n6334_), .B0(new_n30230_), .B1(pi0353), .Y(new_n30855_));
  OR2X1    g28419(.A(new_n27846_), .B(pi0199), .Y(new_n30856_));
  INVX1    g28420(.A(pi1063), .Y(new_n30857_));
  AOI21X1  g28421(.A0(new_n30857_), .A1(pi0199), .B0(new_n30233_), .Y(new_n30858_));
  NAND2X1  g28422(.A(pi0588), .B(pi0451), .Y(new_n30859_));
  NOR4X1   g28423(.A(new_n30859_), .B(new_n30263_), .C(pi0224), .D(pi0223), .Y(new_n30860_));
  AOI21X1  g28424(.A0(new_n30858_), .A1(new_n30856_), .B0(new_n30860_), .Y(new_n30861_));
  OAI21X1  g28425(.A0(new_n30855_), .A1(new_n30675_), .B0(new_n30861_), .Y(new_n30862_));
  AND2X1   g28426(.A(new_n30246_), .B(pi0774), .Y(new_n30863_));
  OAI21X1  g28427(.A0(pi1136), .A1(pi0868), .B0(pi1134), .Y(new_n30864_));
  AOI21X1  g28428(.A0(pi1135), .A1(new_n13538_), .B0(new_n30864_), .Y(new_n30865_));
  NAND3X1  g28429(.A(new_n30865_), .B(new_n30706_), .C(new_n30245_), .Y(new_n30866_));
  OR2X1    g28430(.A(pi1135), .B(pi0636), .Y(new_n30867_));
  AOI21X1  g28431(.A0(pi1135), .A1(pi0650), .B0(new_n4554_), .Y(new_n30868_));
  AOI22X1  g28432(.A0(new_n30868_), .A1(new_n30867_), .B0(new_n30278_), .B1(pi0807), .Y(new_n30869_));
  OAI22X1  g28433(.A0(new_n30869_), .A1(new_n30239_), .B0(new_n30866_), .B1(new_n30863_), .Y(new_n30870_));
  MX2X1    g28434(.A(new_n30870_), .B(new_n30862_), .S0(new_n6713_), .Y(po0876));
  INVX1    g28435(.A(new_n27856_), .Y(new_n30872_));
  AOI22X1  g28436(.A0(new_n30566_), .A1(pi0356), .B0(new_n30565_), .B1(pi0381), .Y(new_n30873_));
  NAND4X1  g28437(.A(new_n6009_), .B(pi0591), .C(new_n6334_), .D(pi0405), .Y(new_n30874_));
  OAI21X1  g28438(.A0(new_n30873_), .A1(pi0591), .B0(new_n30874_), .Y(new_n30875_));
  NOR4X1   g28439(.A(new_n30748_), .B(pi0590), .C(new_n6603_), .D(new_n6557_), .Y(new_n30876_));
  AOI21X1  g28440(.A0(new_n30875_), .A1(new_n6603_), .B0(new_n30876_), .Y(new_n30877_));
  OAI22X1  g28441(.A0(pi1081), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30878_));
  OAI22X1  g28442(.A0(new_n30878_), .A1(new_n30872_), .B0(new_n30877_), .B1(new_n30234_), .Y(new_n30879_));
  NAND2X1  g28443(.A(new_n4622_), .B(pi0750), .Y(new_n30880_));
  AOI21X1  g28444(.A0(pi1135), .A1(pi0684), .B0(new_n4554_), .Y(new_n30881_));
  AOI22X1  g28445(.A0(new_n30881_), .A1(new_n30880_), .B0(new_n30278_), .B1(pi0880), .Y(new_n30882_));
  OR2X1    g28446(.A(pi1135), .B(pi0651), .Y(new_n30883_));
  AOI21X1  g28447(.A0(pi1135), .A1(pi0654), .B0(new_n4554_), .Y(new_n30884_));
  AND3X1   g28448(.A(new_n30278_), .B(new_n30245_), .C(pi0794), .Y(new_n30885_));
  AOI21X1  g28449(.A0(new_n30884_), .A1(new_n30883_), .B0(new_n30885_), .Y(new_n30886_));
  OAI22X1  g28450(.A0(new_n30886_), .A1(new_n30578_), .B0(new_n30882_), .B1(new_n30249_), .Y(new_n30887_));
  MX2X1    g28451(.A(new_n30887_), .B(new_n30879_), .S0(new_n6713_), .Y(po0877));
  INVX1    g28452(.A(pi0795), .Y(new_n30889_));
  AND3X1   g28453(.A(pi0773), .B(pi0769), .C(pi0747), .Y(new_n30890_));
  OAI21X1  g28454(.A0(new_n30890_), .A1(pi0721), .B0(pi0775), .Y(new_n30891_));
  AOI21X1  g28455(.A0(new_n30890_), .A1(pi0721), .B0(new_n30891_), .Y(new_n30892_));
  INVX1    g28456(.A(pi0721), .Y(new_n30893_));
  INVX1    g28457(.A(pi0813), .Y(new_n30894_));
  XOR2X1   g28458(.A(pi0801), .B(pi0773), .Y(new_n30895_));
  XOR2X1   g28459(.A(pi0800), .B(pi0771), .Y(new_n30896_));
  XOR2X1   g28460(.A(pi0794), .B(pi0769), .Y(new_n30897_));
  INVX1    g28461(.A(new_n30897_), .Y(new_n30898_));
  INVX1    g28462(.A(pi0747), .Y(new_n30899_));
  INVX1    g28463(.A(pi0807), .Y(new_n30900_));
  XOR2X1   g28464(.A(pi0798), .B(pi0765), .Y(new_n30901_));
  NOR3X1   g28465(.A(new_n30901_), .B(new_n30900_), .C(new_n30899_), .Y(new_n30902_));
  NOR3X1   g28466(.A(new_n30901_), .B(pi0807), .C(pi0747), .Y(new_n30903_));
  OR2X1    g28467(.A(new_n30903_), .B(new_n30902_), .Y(new_n30904_));
  AND2X1   g28468(.A(new_n30904_), .B(new_n30898_), .Y(new_n30905_));
  INVX1    g28469(.A(new_n30905_), .Y(new_n30906_));
  OR3X1    g28470(.A(new_n30906_), .B(new_n30896_), .C(new_n30895_), .Y(new_n30907_));
  NOR3X1   g28471(.A(new_n30907_), .B(new_n30894_), .C(new_n30893_), .Y(new_n30908_));
  NOR3X1   g28472(.A(new_n30901_), .B(new_n30896_), .C(new_n30900_), .Y(new_n30909_));
  INVX1    g28473(.A(pi0794), .Y(new_n30910_));
  NOR4X1   g28474(.A(pi0813), .B(new_n30630_), .C(new_n30910_), .D(pi0721), .Y(new_n30911_));
  AND2X1   g28475(.A(new_n30911_), .B(new_n30909_), .Y(new_n30912_));
  OAI21X1  g28476(.A0(new_n30912_), .A1(new_n30908_), .B0(pi0816), .Y(new_n30913_));
  AOI21X1  g28477(.A0(new_n30913_), .A1(new_n30892_), .B0(new_n30889_), .Y(new_n30914_));
  INVX1    g28478(.A(pi0945), .Y(new_n30915_));
  AND3X1   g28479(.A(pi0988), .B(new_n30915_), .C(pi0731), .Y(new_n30916_));
  INVX1    g28480(.A(pi0775), .Y(new_n30917_));
  AND2X1   g28481(.A(new_n30917_), .B(pi0721), .Y(new_n30918_));
  OAI21X1  g28482(.A0(new_n30918_), .A1(new_n30892_), .B0(new_n30916_), .Y(new_n30919_));
  XOR2X1   g28483(.A(pi0816), .B(pi0775), .Y(new_n30920_));
  OR4X1    g28484(.A(new_n30920_), .B(new_n30907_), .C(new_n30894_), .D(new_n30893_), .Y(new_n30921_));
  XOR2X1   g28485(.A(pi0795), .B(pi0731), .Y(new_n30922_));
  OR2X1    g28486(.A(new_n30922_), .B(new_n30921_), .Y(new_n30923_));
  NOR2X1   g28487(.A(new_n30916_), .B(new_n30893_), .Y(new_n30924_));
  AOI22X1  g28488(.A0(new_n30924_), .A1(new_n30923_), .B0(new_n30921_), .B1(new_n30918_), .Y(new_n30925_));
  OAI21X1  g28489(.A0(new_n30919_), .A1(new_n30914_), .B0(new_n30925_), .Y(po0878));
  AND3X1   g28490(.A(new_n6009_), .B(pi0591), .C(pi0403), .Y(new_n30927_));
  AOI21X1  g28491(.A0(new_n30227_), .A1(pi0379), .B0(new_n30927_), .Y(new_n30928_));
  OAI22X1  g28492(.A0(new_n30928_), .A1(pi0590), .B0(new_n30256_), .B1(new_n9057_), .Y(new_n30929_));
  NOR2X1   g28493(.A(new_n27848_), .B(pi0199), .Y(new_n30930_));
  OAI22X1  g28494(.A0(pi1045), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30931_));
  OR4X1    g28495(.A(new_n30263_), .B(new_n30234_), .C(new_n6603_), .D(new_n6497_), .Y(new_n30932_));
  OAI21X1  g28496(.A0(new_n30931_), .A1(new_n30930_), .B0(new_n30932_), .Y(new_n30933_));
  AOI21X1  g28497(.A0(new_n30929_), .A1(new_n30674_), .B0(new_n30933_), .Y(new_n30934_));
  NOR2X1   g28498(.A(pi1134), .B(pi0795), .Y(new_n30935_));
  OAI21X1  g28499(.A0(new_n4747_), .A1(pi0851), .B0(new_n4554_), .Y(new_n30936_));
  NOR2X1   g28500(.A(pi1134), .B(pi0640), .Y(new_n30937_));
  AND2X1   g28501(.A(pi1134), .B(pi0776), .Y(new_n30938_));
  OR3X1    g28502(.A(new_n30938_), .B(new_n30937_), .C(new_n4554_), .Y(new_n30939_));
  OAI21X1  g28503(.A0(new_n30936_), .A1(new_n30935_), .B0(new_n30939_), .Y(new_n30940_));
  INVX1    g28504(.A(pi0732), .Y(new_n30941_));
  AND2X1   g28505(.A(pi1136), .B(pi1135), .Y(new_n30942_));
  OAI21X1  g28506(.A0(pi1134), .A1(new_n30941_), .B0(new_n30942_), .Y(new_n30943_));
  AOI21X1  g28507(.A0(pi1134), .A1(pi0694), .B0(new_n30943_), .Y(new_n30944_));
  AOI21X1  g28508(.A0(new_n30940_), .A1(new_n4622_), .B0(new_n30944_), .Y(new_n30945_));
  OAI22X1  g28509(.A0(new_n30945_), .A1(new_n30623_), .B0(new_n30934_), .B1(new_n8943_), .Y(po0879));
  OAI21X1  g28510(.A0(po0980), .A1(new_n14743_), .B0(new_n30112_), .Y(new_n30947_));
  AOI21X1  g28511(.A0(po0980), .A1(new_n30641_), .B0(new_n30947_), .Y(po0880));
  OAI21X1  g28512(.A0(po0980), .A1(new_n14956_), .B0(new_n30112_), .Y(new_n30949_));
  AOI21X1  g28513(.A0(po0980), .A1(new_n30167_), .B0(new_n30949_), .Y(po0881));
  INVX1    g28514(.A(pi1120), .Y(new_n30951_));
  OAI21X1  g28515(.A0(po0980), .A1(new_n14667_), .B0(new_n30112_), .Y(new_n30952_));
  AOI21X1  g28516(.A0(po0980), .A1(new_n30951_), .B0(new_n30952_), .Y(po0882));
  OAI21X1  g28517(.A0(new_n30587_), .A1(pi1126), .B0(new_n30112_), .Y(new_n30954_));
  AOI21X1  g28518(.A0(new_n30587_), .A1(new_n14500_), .B0(new_n30954_), .Y(po0883));
  OAI21X1  g28519(.A0(new_n30587_), .A1(pi1102), .B0(new_n30112_), .Y(new_n30956_));
  AOI21X1  g28520(.A0(new_n30587_), .A1(new_n15292_), .B0(new_n30956_), .Y(po0884));
  INVX1    g28521(.A(pi0728), .Y(new_n30958_));
  OAI21X1  g28522(.A0(po0980), .A1(new_n30958_), .B0(new_n30112_), .Y(new_n30959_));
  AOI21X1  g28523(.A0(po0980), .A1(new_n30187_), .B0(new_n30959_), .Y(po0885));
  OAI21X1  g28524(.A0(new_n30587_), .A1(pi1104), .B0(new_n30112_), .Y(new_n30961_));
  AOI21X1  g28525(.A0(new_n30587_), .A1(new_n15412_), .B0(new_n30961_), .Y(po0886));
  OAI21X1  g28526(.A0(new_n30587_), .A1(pi1106), .B0(new_n30112_), .Y(new_n30963_));
  AOI21X1  g28527(.A0(new_n30587_), .A1(new_n15466_), .B0(new_n30963_), .Y(po0887));
  NAND2X1  g28528(.A(pi0773), .B(pi0747), .Y(new_n30965_));
  XOR2X1   g28529(.A(pi0813), .B(pi0721), .Y(new_n30966_));
  NOR4X1   g28530(.A(new_n30966_), .B(new_n30920_), .C(new_n30907_), .D(new_n30889_), .Y(new_n30967_));
  INVX1    g28531(.A(new_n30967_), .Y(new_n30968_));
  NAND2X1  g28532(.A(new_n30968_), .B(new_n30965_), .Y(new_n30969_));
  INVX1    g28533(.A(pi0731), .Y(new_n30970_));
  NOR2X1   g28534(.A(new_n30967_), .B(new_n30970_), .Y(new_n30971_));
  INVX1    g28535(.A(new_n30971_), .Y(new_n30972_));
  AND2X1   g28536(.A(pi0988), .B(new_n30915_), .Y(new_n30973_));
  OR2X1    g28537(.A(new_n30966_), .B(new_n30920_), .Y(new_n30974_));
  NOR4X1   g28538(.A(new_n30974_), .B(new_n30897_), .C(new_n30630_), .D(pi0795), .Y(new_n30975_));
  AOI21X1  g28539(.A0(new_n30975_), .A1(new_n30909_), .B0(new_n30965_), .Y(new_n30976_));
  OAI21X1  g28540(.A0(new_n30976_), .A1(pi0731), .B0(new_n30973_), .Y(new_n30977_));
  AOI22X1  g28541(.A0(new_n30977_), .A1(new_n30972_), .B0(new_n30969_), .B1(new_n30916_), .Y(po0888));
  OAI21X1  g28542(.A0(po0954), .A1(new_n30941_), .B0(new_n30112_), .Y(new_n30979_));
  AOI21X1  g28543(.A0(po0954), .A1(new_n30152_), .B0(new_n30979_), .Y(po0889));
  NAND4X1  g28544(.A(new_n30233_), .B(pi0592), .C(new_n6069_), .D(pi0375), .Y(new_n30981_));
  NAND4X1  g28545(.A(new_n30233_), .B(new_n6009_), .C(pi0591), .D(pi0399), .Y(new_n30982_));
  AOI21X1  g28546(.A0(new_n30982_), .A1(new_n30981_), .B0(pi0590), .Y(new_n30983_));
  AND3X1   g28547(.A(new_n30230_), .B(new_n30233_), .C(pi0316), .Y(new_n30984_));
  OAI21X1  g28548(.A0(new_n30984_), .A1(new_n30983_), .B0(new_n6603_), .Y(new_n30985_));
  MX2X1    g28549(.A(pi0308), .B(pi1037), .S0(pi0200), .Y(new_n30986_));
  NOR2X1   g28550(.A(new_n30986_), .B(pi0199), .Y(new_n30987_));
  OAI22X1  g28551(.A0(pi1047), .A1(new_n7871_), .B0(pi0224), .B1(pi0223), .Y(new_n30988_));
  OR2X1    g28552(.A(new_n30988_), .B(new_n30987_), .Y(new_n30989_));
  INVX1    g28553(.A(pi0424), .Y(new_n30990_));
  OR4X1    g28554(.A(new_n30702_), .B(pi0590), .C(new_n6603_), .D(new_n30990_), .Y(new_n30991_));
  AND3X1   g28555(.A(new_n30991_), .B(new_n30989_), .C(new_n6713_), .Y(new_n30992_));
  NAND2X1  g28556(.A(new_n30246_), .B(pi0777), .Y(new_n30993_));
  OAI21X1  g28557(.A0(pi1136), .A1(pi0838), .B0(pi1134), .Y(new_n30994_));
  AOI21X1  g28558(.A0(pi1135), .A1(pi0737), .B0(new_n30994_), .Y(new_n30995_));
  NAND3X1  g28559(.A(new_n30995_), .B(new_n30993_), .C(new_n30707_), .Y(new_n30996_));
  OAI21X1  g28560(.A0(new_n4622_), .A1(pi0648), .B0(new_n4747_), .Y(new_n30997_));
  AOI21X1  g28561(.A0(new_n4622_), .A1(new_n12509_), .B0(new_n30997_), .Y(new_n30998_));
  AOI21X1  g28562(.A0(new_n30998_), .A1(new_n30359_), .B0(new_n6713_), .Y(new_n30999_));
  AOI22X1  g28563(.A0(new_n30999_), .A1(new_n30996_), .B0(new_n30992_), .B1(new_n30985_), .Y(po0890));
  INVX1    g28564(.A(pi1119), .Y(new_n31001_));
  OAI21X1  g28565(.A0(po0980), .A1(new_n15095_), .B0(new_n30112_), .Y(new_n31002_));
  AOI21X1  g28566(.A0(po0980), .A1(new_n31001_), .B0(new_n31002_), .Y(po0891));
  OAI21X1  g28567(.A0(new_n30587_), .A1(pi1109), .B0(new_n30112_), .Y(new_n31004_));
  AOI21X1  g28568(.A0(new_n30587_), .A1(new_n13171_), .B0(new_n31004_), .Y(po0892));
  OAI21X1  g28569(.A0(new_n30587_), .A1(pi1101), .B0(new_n30112_), .Y(new_n31006_));
  AOI21X1  g28570(.A0(new_n30587_), .A1(new_n13832_), .B0(new_n31006_), .Y(po0893));
  INVX1    g28571(.A(pi1122), .Y(new_n31008_));
  OAI21X1  g28572(.A0(po0980), .A1(new_n15220_), .B0(new_n30112_), .Y(new_n31009_));
  AOI21X1  g28573(.A0(po0980), .A1(new_n31008_), .B0(new_n31009_), .Y(po0894));
  INVX1    g28574(.A(pi1121), .Y(new_n31011_));
  OAI21X1  g28575(.A0(po0980), .A1(new_n11771_), .B0(new_n30112_), .Y(new_n31012_));
  AOI21X1  g28576(.A0(po0980), .A1(new_n31011_), .B0(new_n31012_), .Y(po0895));
  NOR4X1   g28577(.A(new_n30042_), .B(pi1061), .C(pi0952), .D(new_n12767_), .Y(po0988));
  AND2X1   g28578(.A(po0988), .B(pi1108), .Y(new_n31015_));
  OAI21X1  g28579(.A0(po0988), .A1(new_n15571_), .B0(new_n30060_), .Y(new_n31016_));
  OR2X1    g28580(.A(new_n31016_), .B(new_n31015_), .Y(po0896));
  AOI21X1  g28581(.A0(po0988), .A1(pi1114), .B0(pi0966), .Y(new_n31018_));
  OAI21X1  g28582(.A0(po0988), .A1(pi0741), .B0(new_n31018_), .Y(po0898));
  AOI21X1  g28583(.A0(po0988), .A1(pi1112), .B0(pi0966), .Y(new_n31020_));
  OAI21X1  g28584(.A0(po0988), .A1(pi0742), .B0(new_n31020_), .Y(po0899));
  AND2X1   g28585(.A(po0988), .B(pi1109), .Y(new_n31022_));
  OAI21X1  g28586(.A0(po0988), .A1(new_n13086_), .B0(new_n30060_), .Y(new_n31023_));
  OR2X1    g28587(.A(new_n31023_), .B(new_n31022_), .Y(po0900));
  AOI21X1  g28588(.A0(po0988), .A1(pi1131), .B0(pi0966), .Y(new_n31025_));
  OAI21X1  g28589(.A0(po0988), .A1(pi0744), .B0(new_n31025_), .Y(po0901));
  AOI21X1  g28590(.A0(po0988), .A1(pi1111), .B0(pi0966), .Y(new_n31027_));
  OAI21X1  g28591(.A0(po0988), .A1(pi0745), .B0(new_n31027_), .Y(po0902));
  AND2X1   g28592(.A(po0988), .B(pi1104), .Y(new_n31029_));
  OAI21X1  g28593(.A0(po0988), .A1(new_n15416_), .B0(new_n30060_), .Y(new_n31030_));
  OR2X1    g28594(.A(new_n31030_), .B(new_n31029_), .Y(po0903));
  NOR4X1   g28595(.A(new_n30901_), .B(pi0807), .C(new_n30630_), .D(pi0747), .Y(new_n31032_));
  AND3X1   g28596(.A(pi0988), .B(new_n30915_), .C(pi0773), .Y(new_n31033_));
  NOR4X1   g28597(.A(new_n31033_), .B(new_n30901_), .C(new_n30895_), .D(new_n30900_), .Y(new_n31034_));
  OR2X1    g28598(.A(new_n31034_), .B(new_n31032_), .Y(new_n31035_));
  OR3X1    g28599(.A(new_n30966_), .B(new_n30922_), .C(new_n30920_), .Y(new_n31036_));
  NOR3X1   g28600(.A(new_n31036_), .B(new_n30897_), .C(new_n30896_), .Y(new_n31037_));
  INVX1    g28601(.A(pi0988), .Y(new_n31038_));
  OR3X1    g28602(.A(new_n30965_), .B(new_n31038_), .C(pi0945), .Y(new_n31039_));
  OAI21X1  g28603(.A0(new_n31033_), .A1(pi0747), .B0(new_n31039_), .Y(new_n31040_));
  AOI21X1  g28604(.A0(new_n31037_), .A1(new_n31035_), .B0(new_n31040_), .Y(po0904));
  AND2X1   g28605(.A(po0988), .B(pi1106), .Y(new_n31042_));
  OAI21X1  g28606(.A0(po0988), .A1(new_n15462_), .B0(new_n30060_), .Y(new_n31043_));
  OR2X1    g28607(.A(new_n31043_), .B(new_n31042_), .Y(po0905));
  AND2X1   g28608(.A(po0988), .B(pi1105), .Y(new_n31045_));
  OAI21X1  g28609(.A0(po0988), .A1(new_n12774_), .B0(new_n30060_), .Y(new_n31046_));
  OR2X1    g28610(.A(new_n31046_), .B(new_n31045_), .Y(po0906));
  AOI21X1  g28611(.A0(po0988), .A1(pi1130), .B0(pi0966), .Y(new_n31048_));
  OAI21X1  g28612(.A0(po0988), .A1(pi0750), .B0(new_n31048_), .Y(po0907));
  AOI21X1  g28613(.A0(po0988), .A1(pi1123), .B0(pi0966), .Y(new_n31050_));
  OAI21X1  g28614(.A0(po0988), .A1(pi0751), .B0(new_n31050_), .Y(po0908));
  AOI21X1  g28615(.A0(po0988), .A1(pi1124), .B0(pi0966), .Y(new_n31052_));
  OAI21X1  g28616(.A0(po0988), .A1(pi0752), .B0(new_n31052_), .Y(po0909));
  AOI21X1  g28617(.A0(po0988), .A1(pi1117), .B0(pi0966), .Y(new_n31054_));
  OAI21X1  g28618(.A0(po0988), .A1(pi0753), .B0(new_n31054_), .Y(po0910));
  AOI21X1  g28619(.A0(po0988), .A1(pi1118), .B0(pi0966), .Y(new_n31056_));
  OAI21X1  g28620(.A0(po0988), .A1(pi0754), .B0(new_n31056_), .Y(po0911));
  AOI21X1  g28621(.A0(po0988), .A1(pi1120), .B0(pi0966), .Y(new_n31058_));
  OAI21X1  g28622(.A0(po0988), .A1(pi0755), .B0(new_n31058_), .Y(po0912));
  AOI21X1  g28623(.A0(po0988), .A1(pi1119), .B0(pi0966), .Y(new_n31060_));
  OAI21X1  g28624(.A0(po0988), .A1(pi0756), .B0(new_n31060_), .Y(po0913));
  AOI21X1  g28625(.A0(po0988), .A1(pi1113), .B0(pi0966), .Y(new_n31062_));
  OAI21X1  g28626(.A0(po0988), .A1(pi0757), .B0(new_n31062_), .Y(po0914));
  AND2X1   g28627(.A(po0988), .B(pi1101), .Y(new_n31064_));
  OAI21X1  g28628(.A0(po0988), .A1(new_n13836_), .B0(new_n30060_), .Y(new_n31065_));
  OR2X1    g28629(.A(new_n31065_), .B(new_n31064_), .Y(po0915));
  NOR2X1   g28630(.A(po0988), .B(pi0759), .Y(new_n31067_));
  NOR4X1   g28631(.A(new_n30045_), .B(new_n30042_), .C(pi1061), .D(pi0952), .Y(new_n31068_));
  OAI21X1  g28632(.A0(new_n31068_), .A1(new_n31067_), .B0(new_n30060_), .Y(po0916));
  AOI21X1  g28633(.A0(po0988), .A1(pi1115), .B0(pi0966), .Y(new_n31070_));
  OAI21X1  g28634(.A0(po0988), .A1(pi0760), .B0(new_n31070_), .Y(po0917));
  AOI21X1  g28635(.A0(po0988), .A1(pi1121), .B0(pi0966), .Y(new_n31072_));
  OAI21X1  g28636(.A0(po0988), .A1(pi0761), .B0(new_n31072_), .Y(po0918));
  AOI21X1  g28637(.A0(po0988), .A1(pi1129), .B0(pi0966), .Y(new_n31074_));
  OAI21X1  g28638(.A0(po0988), .A1(pi0762), .B0(new_n31074_), .Y(po0919));
  INVX1    g28639(.A(pi1103), .Y(new_n31076_));
  INVX1    g28640(.A(po0988), .Y(new_n31077_));
  AOI21X1  g28641(.A0(new_n31077_), .A1(pi0763), .B0(pi0966), .Y(new_n31078_));
  OAI21X1  g28642(.A0(new_n31077_), .A1(new_n31076_), .B0(new_n31078_), .Y(po0920));
  INVX1    g28643(.A(pi1107), .Y(new_n31080_));
  AOI21X1  g28644(.A0(new_n31077_), .A1(pi0764), .B0(pi0966), .Y(new_n31081_));
  OAI21X1  g28645(.A0(new_n31077_), .A1(new_n31080_), .B0(new_n31081_), .Y(po0921));
  INVX1    g28646(.A(pi0765), .Y(new_n31083_));
  NOR4X1   g28647(.A(new_n31036_), .B(new_n30906_), .C(new_n30896_), .D(new_n30895_), .Y(po0978));
  OR2X1    g28648(.A(po0978), .B(new_n31083_), .Y(new_n31085_));
  AND2X1   g28649(.A(new_n31085_), .B(pi0945), .Y(new_n31086_));
  AOI21X1  g28650(.A0(new_n30894_), .A1(new_n30893_), .B0(new_n30908_), .Y(new_n31087_));
  NOR2X1   g28651(.A(new_n30906_), .B(new_n30896_), .Y(new_n31088_));
  OR2X1    g28652(.A(pi0801), .B(pi0773), .Y(new_n31089_));
  NAND2X1  g28653(.A(pi0801), .B(pi0773), .Y(new_n31090_));
  AND2X1   g28654(.A(pi0800), .B(pi0771), .Y(new_n31091_));
  AND2X1   g28655(.A(pi0794), .B(pi0769), .Y(new_n31092_));
  NOR4X1   g28656(.A(new_n30902_), .B(new_n31092_), .C(new_n31091_), .D(pi0765), .Y(new_n31093_));
  OAI21X1  g28657(.A0(new_n31093_), .A1(new_n31089_), .B0(new_n31090_), .Y(new_n31094_));
  AOI21X1  g28658(.A0(new_n31094_), .A1(new_n31088_), .B0(pi0721), .Y(new_n31095_));
  OR4X1    g28659(.A(new_n31095_), .B(new_n31087_), .C(pi0816), .D(pi0775), .Y(new_n31096_));
  AND2X1   g28660(.A(pi0816), .B(pi0775), .Y(new_n31097_));
  NOR4X1   g28661(.A(new_n30966_), .B(new_n30906_), .C(new_n30896_), .D(new_n30895_), .Y(new_n31098_));
  AOI21X1  g28662(.A0(new_n31098_), .A1(new_n31097_), .B0(pi0765), .Y(new_n31099_));
  NAND2X1  g28663(.A(new_n31099_), .B(new_n31096_), .Y(new_n31100_));
  AOI21X1  g28664(.A0(new_n31100_), .A1(new_n30889_), .B0(pi0731), .Y(new_n31101_));
  NOR3X1   g28665(.A(new_n31100_), .B(pi0795), .C(pi0731), .Y(new_n31102_));
  OAI22X1  g28666(.A0(new_n31102_), .A1(new_n31083_), .B0(new_n31101_), .B1(new_n30971_), .Y(new_n31103_));
  AOI21X1  g28667(.A0(new_n31103_), .A1(new_n30915_), .B0(new_n31086_), .Y(po0922));
  INVX1    g28668(.A(pi1110), .Y(new_n31105_));
  AOI21X1  g28669(.A0(new_n31077_), .A1(pi0766), .B0(pi0966), .Y(new_n31106_));
  OAI21X1  g28670(.A0(new_n31077_), .A1(new_n31105_), .B0(new_n31106_), .Y(po0923));
  AOI21X1  g28671(.A0(po0988), .A1(pi1116), .B0(pi0966), .Y(new_n31108_));
  OAI21X1  g28672(.A0(po0988), .A1(pi0767), .B0(new_n31108_), .Y(po0924));
  AOI21X1  g28673(.A0(po0988), .A1(pi1125), .B0(pi0966), .Y(new_n31110_));
  OAI21X1  g28674(.A0(po0988), .A1(pi0768), .B0(new_n31110_), .Y(po0925));
  AND2X1   g28675(.A(new_n31098_), .B(new_n31097_), .Y(new_n31112_));
  NOR4X1   g28676(.A(new_n30974_), .B(new_n30896_), .C(new_n30895_), .D(new_n30910_), .Y(new_n31113_));
  AND3X1   g28677(.A(new_n31113_), .B(new_n30904_), .C(new_n30917_), .Y(new_n31114_));
  OAI21X1  g28678(.A0(new_n31114_), .A1(new_n31112_), .B0(pi0795), .Y(new_n31115_));
  AND3X1   g28679(.A(pi0775), .B(pi0773), .C(pi0747), .Y(new_n31116_));
  XOR2X1   g28680(.A(new_n31116_), .B(pi0769), .Y(new_n31117_));
  AND3X1   g28681(.A(new_n31117_), .B(new_n31115_), .C(new_n30916_), .Y(new_n31118_));
  INVX1    g28682(.A(pi0769), .Y(new_n31119_));
  INVX1    g28683(.A(new_n30922_), .Y(new_n31120_));
  AND3X1   g28684(.A(new_n31113_), .B(new_n31120_), .C(new_n30904_), .Y(new_n31121_));
  NOR3X1   g28685(.A(new_n31121_), .B(new_n30916_), .C(new_n31119_), .Y(new_n31122_));
  OR2X1    g28686(.A(new_n31122_), .B(new_n31118_), .Y(po0926));
  AOI21X1  g28687(.A0(po0988), .A1(pi1126), .B0(pi0966), .Y(new_n31124_));
  OAI21X1  g28688(.A0(po0988), .A1(pi0770), .B0(new_n31124_), .Y(po0927));
  INVX1    g28689(.A(new_n31098_), .Y(new_n31126_));
  NOR2X1   g28690(.A(pi0795), .B(pi0731), .Y(new_n31127_));
  NOR3X1   g28691(.A(new_n31095_), .B(pi0816), .C(pi0775), .Y(new_n31128_));
  OAI21X1  g28692(.A0(new_n31128_), .A1(new_n31097_), .B0(new_n31127_), .Y(new_n31129_));
  NOR3X1   g28693(.A(new_n30920_), .B(new_n30889_), .C(new_n30970_), .Y(new_n31130_));
  INVX1    g28694(.A(new_n31130_), .Y(new_n31131_));
  AOI21X1  g28695(.A0(new_n31131_), .A1(new_n31129_), .B0(new_n31126_), .Y(po0963));
  NAND2X1  g28696(.A(pi0987), .B(new_n30915_), .Y(new_n31133_));
  NAND2X1  g28697(.A(pi0945), .B(pi0771), .Y(new_n31134_));
  OAI22X1  g28698(.A0(new_n31134_), .A1(po0978), .B0(new_n31133_), .B1(po0963), .Y(po0928));
  AND2X1   g28699(.A(po0988), .B(pi1102), .Y(new_n31136_));
  OAI21X1  g28700(.A0(po0988), .A1(new_n15306_), .B0(new_n30060_), .Y(new_n31137_));
  OR2X1    g28701(.A(new_n31137_), .B(new_n31136_), .Y(po0929));
  NAND3X1  g28702(.A(po0963), .B(new_n31088_), .C(new_n30630_), .Y(new_n31139_));
  NAND2X1  g28703(.A(new_n31139_), .B(new_n30973_), .Y(new_n31140_));
  AND2X1   g28704(.A(new_n31036_), .B(pi0801), .Y(new_n31141_));
  OAI21X1  g28705(.A0(new_n31141_), .A1(new_n30907_), .B0(pi0773), .Y(new_n31142_));
  AOI21X1  g28706(.A0(new_n31142_), .A1(new_n31140_), .B0(new_n31033_), .Y(po0930));
  AOI21X1  g28707(.A0(po0988), .A1(pi1127), .B0(pi0966), .Y(new_n31144_));
  OAI21X1  g28708(.A0(po0988), .A1(pi0774), .B0(new_n31144_), .Y(po0931));
  OR2X1    g28709(.A(po0978), .B(new_n30917_), .Y(new_n31146_));
  AND2X1   g28710(.A(new_n30915_), .B(pi0731), .Y(new_n31147_));
  NAND4X1  g28711(.A(pi0773), .B(pi0771), .C(pi0765), .D(pi0747), .Y(new_n31148_));
  NAND2X1  g28712(.A(pi0800), .B(pi0795), .Y(new_n31149_));
  NOR4X1   g28713(.A(new_n31149_), .B(new_n30966_), .C(pi0816), .D(new_n30630_), .Y(new_n31150_));
  AOI21X1  g28714(.A0(new_n31150_), .A1(new_n30905_), .B0(new_n31148_), .Y(new_n31151_));
  OAI21X1  g28715(.A0(new_n31151_), .A1(pi0775), .B0(new_n31147_), .Y(new_n31152_));
  NAND2X1  g28716(.A(new_n31148_), .B(new_n30968_), .Y(new_n31153_));
  AND3X1   g28717(.A(new_n30915_), .B(pi0775), .C(pi0731), .Y(new_n31154_));
  AOI22X1  g28718(.A0(new_n31154_), .A1(new_n31153_), .B0(new_n31152_), .B1(new_n31146_), .Y(po0932));
  AOI21X1  g28719(.A0(po0988), .A1(pi1128), .B0(pi0966), .Y(new_n31156_));
  OAI21X1  g28720(.A0(po0988), .A1(pi0776), .B0(new_n31156_), .Y(po0933));
  AOI21X1  g28721(.A0(po0988), .A1(pi1122), .B0(pi0966), .Y(new_n31158_));
  OAI21X1  g28722(.A0(po0988), .A1(pi0777), .B0(new_n31158_), .Y(po0934));
  NOR2X1   g28723(.A(pi1083), .B(pi1046), .Y(new_n31160_));
  NAND4X1  g28724(.A(new_n31160_), .B(pi1085), .C(pi0956), .D(pi0832), .Y(new_n31161_));
  OR2X1    g28725(.A(new_n31161_), .B(pi0968), .Y(new_n31162_));
  MX2X1    g28726(.A(pi1100), .B(pi0778), .S0(new_n31162_), .Y(po0935));
  OAI21X1  g28727(.A0(new_n30021_), .A1(new_n5277_), .B0(pi0779), .Y(po0936));
  OAI21X1  g28728(.A0(new_n30021_), .A1(new_n5362_), .B0(pi0780), .Y(po0937));
  MX2X1    g28729(.A(pi1101), .B(pi0781), .S0(new_n31162_), .Y(po0938));
  AOI22X1  g28730(.A0(new_n5222_), .A1(new_n5026_), .B0(pi0983), .B1(new_n2933_), .Y(new_n31167_));
  NAND2X1  g28731(.A(new_n31167_), .B(new_n30021_), .Y(po0939));
  MX2X1    g28732(.A(pi1109), .B(pi0783), .S0(new_n31162_), .Y(po0940));
  MX2X1    g28733(.A(pi1110), .B(pi0784), .S0(new_n31162_), .Y(po0941));
  MX2X1    g28734(.A(pi1102), .B(pi0785), .S0(new_n31162_), .Y(po0942));
  MX2X1    g28735(.A(new_n7648_), .B(new_n5777_), .S0(po1110), .Y(po0943));
  MX2X1    g28736(.A(pi1104), .B(pi0787), .S0(new_n31162_), .Y(po0944));
  MX2X1    g28737(.A(pi1105), .B(pi0788), .S0(new_n31162_), .Y(po0945));
  MX2X1    g28738(.A(pi1106), .B(pi0789), .S0(new_n31162_), .Y(po0946));
  MX2X1    g28739(.A(pi1107), .B(pi0790), .S0(new_n31162_), .Y(po0947));
  MX2X1    g28740(.A(pi1108), .B(pi0791), .S0(new_n31162_), .Y(po0948));
  MX2X1    g28741(.A(pi1103), .B(pi0792), .S0(new_n31162_), .Y(po0949));
  AND2X1   g28742(.A(pi0956), .B(pi0832), .Y(new_n31179_));
  NAND4X1  g28743(.A(new_n31160_), .B(new_n31179_), .C(pi1085), .D(pi0968), .Y(new_n31180_));
  MX2X1    g28744(.A(pi1130), .B(pi0794), .S0(new_n31180_), .Y(po0951));
  MX2X1    g28745(.A(pi1128), .B(pi0795), .S0(new_n31180_), .Y(po0952));
  NAND2X1  g28746(.A(pi0279), .B(pi0278), .Y(new_n31183_));
  NOR4X1   g28747(.A(new_n31183_), .B(pi0280), .C(pi0269), .D(new_n4470_), .Y(new_n31184_));
  AND3X1   g28748(.A(new_n31184_), .B(new_n30215_), .C(new_n30211_), .Y(new_n31185_));
  XOR2X1   g28749(.A(new_n31185_), .B(new_n3521_), .Y(po0953));
  MX2X1    g28750(.A(pi1124), .B(pi0798), .S0(new_n31180_), .Y(po0955));
  INVX1    g28751(.A(pi0799), .Y(new_n31188_));
  MX2X1    g28752(.A(pi1107), .B(new_n31188_), .S0(new_n31180_), .Y(po0956));
  MX2X1    g28753(.A(pi1125), .B(pi0800), .S0(new_n31180_), .Y(po0957));
  MX2X1    g28754(.A(pi1126), .B(pi0801), .S0(new_n31180_), .Y(po0958));
  AND3X1   g28755(.A(new_n30215_), .B(new_n30214_), .C(new_n3521_), .Y(new_n31192_));
  AND3X1   g28756(.A(new_n31192_), .B(new_n3313_), .C(new_n30210_), .Y(po0959));
  INVX1    g28757(.A(pi0803), .Y(new_n31194_));
  MX2X1    g28758(.A(pi1106), .B(new_n31194_), .S0(new_n31180_), .Y(po0960));
  MX2X1    g28759(.A(pi1109), .B(pi0804), .S0(new_n31180_), .Y(po0961));
  NAND4X1  g28760(.A(new_n30213_), .B(new_n3963_), .C(new_n30211_), .D(new_n4260_), .Y(new_n31197_));
  XOR2X1   g28761(.A(new_n31197_), .B(pi0270), .Y(po0962));
  MX2X1    g28762(.A(pi1127), .B(pi0807), .S0(new_n31180_), .Y(po0964));
  MX2X1    g28763(.A(pi1101), .B(pi0808), .S0(new_n31180_), .Y(po0965));
  INVX1    g28764(.A(pi0809), .Y(new_n31201_));
  MX2X1    g28765(.A(pi1103), .B(new_n31201_), .S0(new_n31180_), .Y(po0966));
  MX2X1    g28766(.A(pi1108), .B(pi0810), .S0(new_n31180_), .Y(po0967));
  MX2X1    g28767(.A(pi1102), .B(pi0811), .S0(new_n31180_), .Y(po0968));
  INVX1    g28768(.A(pi0812), .Y(new_n31205_));
  MX2X1    g28769(.A(pi1104), .B(new_n31205_), .S0(new_n31180_), .Y(po0969));
  MX2X1    g28770(.A(pi1131), .B(pi0813), .S0(new_n31180_), .Y(po0970));
  INVX1    g28771(.A(pi0814), .Y(new_n31208_));
  MX2X1    g28772(.A(pi1105), .B(new_n31208_), .S0(new_n31180_), .Y(po0971));
  MX2X1    g28773(.A(pi1110), .B(pi0815), .S0(new_n31180_), .Y(po0972));
  MX2X1    g28774(.A(pi1129), .B(pi0816), .S0(new_n31180_), .Y(po0973));
  XOR2X1   g28775(.A(new_n30213_), .B(new_n4260_), .Y(po0974));
  OAI21X1  g28776(.A0(new_n10215_), .A1(new_n8943_), .B0(new_n10076_), .Y(po0975));
  XOR2X1   g28777(.A(new_n31192_), .B(new_n30210_), .Y(po0976));
  OR2X1    g28778(.A(new_n31197_), .B(pi0270), .Y(new_n31215_));
  AOI22X1  g28779(.A0(new_n31215_), .A1(pi0277), .B0(new_n30215_), .B1(new_n30214_), .Y(po0977));
  NOR2X1   g28780(.A(pi0893), .B(pi0811), .Y(po0979));
  OAI22X1  g28781(.A0(new_n7555_), .A1(pi0982), .B0(new_n8943_), .B1(new_n5968_), .Y(new_n31218_));
  AND2X1   g28782(.A(new_n31218_), .B(new_n5225_), .Y(po0981));
  AND2X1   g28783(.A(new_n2990_), .B(pi0123), .Y(new_n31220_));
  INVX1    g28784(.A(new_n31220_), .Y(new_n31221_));
  OAI22X1  g28785(.A0(new_n2991_), .A1(new_n27864_), .B0(pi1131), .B1(pi1127), .Y(new_n31222_));
  OAI21X1  g28786(.A0(new_n31221_), .A1(pi0825), .B0(new_n31222_), .Y(new_n31223_));
  AOI21X1  g28787(.A0(new_n2990_), .A1(pi0123), .B0(new_n30142_), .Y(new_n31224_));
  NAND2X1  g28788(.A(new_n31224_), .B(pi1131), .Y(new_n31225_));
  NAND2X1  g28789(.A(new_n31225_), .B(new_n31223_), .Y(new_n31226_));
  XOR2X1   g28790(.A(pi1130), .B(new_n30197_), .Y(new_n31227_));
  XOR2X1   g28791(.A(pi1129), .B(pi1128), .Y(new_n31228_));
  XOR2X1   g28792(.A(pi1126), .B(pi1125), .Y(new_n31229_));
  XOR2X1   g28793(.A(new_n31229_), .B(new_n31228_), .Y(new_n31230_));
  XOR2X1   g28794(.A(new_n31230_), .B(new_n31227_), .Y(new_n31231_));
  INVX1    g28795(.A(pi0825), .Y(po1147));
  OAI21X1  g28796(.A0(new_n31221_), .A1(po1147), .B0(new_n31222_), .Y(new_n31233_));
  AOI21X1  g28797(.A0(new_n31224_), .A1(pi1131), .B0(new_n31231_), .Y(new_n31234_));
  AOI22X1  g28798(.A0(new_n31234_), .A1(new_n31233_), .B0(new_n31231_), .B1(new_n31226_), .Y(po0982));
  OAI22X1  g28799(.A0(new_n2991_), .A1(new_n27864_), .B0(pi1123), .B1(pi1122), .Y(new_n31236_));
  OAI21X1  g28800(.A0(new_n31221_), .A1(pi0826), .B0(new_n31236_), .Y(new_n31237_));
  AOI21X1  g28801(.A0(new_n2990_), .A1(pi0123), .B0(new_n31008_), .Y(new_n31238_));
  NAND2X1  g28802(.A(new_n31238_), .B(pi1123), .Y(new_n31239_));
  NAND2X1  g28803(.A(new_n31239_), .B(new_n31237_), .Y(new_n31240_));
  XOR2X1   g28804(.A(pi1119), .B(new_n30715_), .Y(new_n31241_));
  XOR2X1   g28805(.A(pi1121), .B(pi1120), .Y(new_n31242_));
  XOR2X1   g28806(.A(pi1117), .B(pi1116), .Y(new_n31243_));
  XOR2X1   g28807(.A(new_n31243_), .B(new_n31242_), .Y(new_n31244_));
  XOR2X1   g28808(.A(new_n31244_), .B(new_n31241_), .Y(new_n31245_));
  INVX1    g28809(.A(pi0826), .Y(po1148));
  OAI21X1  g28810(.A0(new_n31221_), .A1(po1148), .B0(new_n31236_), .Y(new_n31247_));
  AOI21X1  g28811(.A0(new_n31238_), .A1(pi1123), .B0(new_n31245_), .Y(new_n31248_));
  AOI22X1  g28812(.A0(new_n31248_), .A1(new_n31247_), .B0(new_n31245_), .B1(new_n31240_), .Y(po0983));
  OAI22X1  g28813(.A0(new_n2991_), .A1(new_n27864_), .B0(pi1107), .B1(pi1100), .Y(new_n31250_));
  OAI21X1  g28814(.A0(new_n31221_), .A1(pi0827), .B0(new_n31250_), .Y(new_n31251_));
  AOI21X1  g28815(.A0(new_n2990_), .A1(pi0123), .B0(new_n31080_), .Y(new_n31252_));
  NAND2X1  g28816(.A(new_n31252_), .B(pi1100), .Y(new_n31253_));
  NAND2X1  g28817(.A(new_n31253_), .B(new_n31251_), .Y(new_n31254_));
  XOR2X1   g28818(.A(pi1105), .B(new_n31076_), .Y(new_n31255_));
  XOR2X1   g28819(.A(pi1102), .B(pi1101), .Y(new_n31256_));
  XOR2X1   g28820(.A(pi1106), .B(pi1104), .Y(new_n31257_));
  XOR2X1   g28821(.A(new_n31257_), .B(new_n31256_), .Y(new_n31258_));
  XOR2X1   g28822(.A(new_n31258_), .B(new_n31255_), .Y(new_n31259_));
  INVX1    g28823(.A(pi0827), .Y(po1178));
  OAI21X1  g28824(.A0(new_n31221_), .A1(po1178), .B0(new_n31250_), .Y(new_n31261_));
  AOI21X1  g28825(.A0(new_n31252_), .A1(pi1100), .B0(new_n31259_), .Y(new_n31262_));
  AOI22X1  g28826(.A0(new_n31262_), .A1(new_n31261_), .B0(new_n31259_), .B1(new_n31254_), .Y(po0984));
  OAI22X1  g28827(.A0(new_n2991_), .A1(new_n27864_), .B0(pi1115), .B1(pi1114), .Y(new_n31264_));
  OAI21X1  g28828(.A0(new_n31221_), .A1(pi0828), .B0(new_n31264_), .Y(new_n31265_));
  AOI21X1  g28829(.A0(new_n2990_), .A1(pi0123), .B0(new_n30167_), .Y(new_n31266_));
  NAND2X1  g28830(.A(new_n31266_), .B(pi1115), .Y(new_n31267_));
  NAND2X1  g28831(.A(new_n31267_), .B(new_n31265_), .Y(new_n31268_));
  XOR2X1   g28832(.A(pi1111), .B(new_n31105_), .Y(new_n31269_));
  XOR2X1   g28833(.A(pi1113), .B(pi1112), .Y(new_n31270_));
  XOR2X1   g28834(.A(pi1109), .B(pi1108), .Y(new_n31271_));
  XOR2X1   g28835(.A(new_n31271_), .B(new_n31270_), .Y(new_n31272_));
  XOR2X1   g28836(.A(new_n31272_), .B(new_n31269_), .Y(new_n31273_));
  INVX1    g28837(.A(pi0828), .Y(po1182));
  OAI21X1  g28838(.A0(new_n31221_), .A1(po1182), .B0(new_n31264_), .Y(new_n31275_));
  AOI21X1  g28839(.A0(new_n31266_), .A1(pi1115), .B0(new_n31273_), .Y(new_n31276_));
  AOI22X1  g28840(.A0(new_n31276_), .A1(new_n31275_), .B0(new_n31273_), .B1(new_n31268_), .Y(po0985));
  NAND2X1  g28841(.A(new_n6713_), .B(new_n2759_), .Y(new_n31278_));
  AOI21X1  g28842(.A0(new_n31278_), .A1(pi0951), .B0(new_n5024_), .Y(po0986));
  XOR2X1   g28843(.A(new_n31184_), .B(new_n30211_), .Y(po0987));
  NOR4X1   g28844(.A(new_n6717_), .B(new_n6715_), .C(new_n2702_), .D(pi0832), .Y(po0989));
  OAI22X1  g28845(.A0(new_n10098_), .A1(new_n5024_), .B0(new_n2720_), .B1(new_n2701_), .Y(po0990));
  AND3X1   g28846(.A(pi1093), .B(pi1092), .C(pi0946), .Y(po0991));
  XOR2X1   g28847(.A(new_n30214_), .B(new_n3963_), .Y(po0992));
  MX2X1    g28848(.A(pi1049), .B(pi0837), .S0(pi0955), .Y(po0993));
  MX2X1    g28849(.A(pi1047), .B(pi0838), .S0(pi0955), .Y(po0994));
  MX2X1    g28850(.A(pi1074), .B(pi0839), .S0(pi0955), .Y(po0995));
  MX2X1    g28851(.A(pi0840), .B(pi1196), .S0(new_n2720_), .Y(po0996));
  AND3X1   g28852(.A(new_n6787_), .B(new_n6783_), .C(new_n7298_), .Y(po0997));
  MX2X1    g28853(.A(pi1035), .B(pi0842), .S0(pi0955), .Y(po0998));
  MX2X1    g28854(.A(pi1079), .B(pi0843), .S0(pi0955), .Y(po0999));
  MX2X1    g28855(.A(pi1078), .B(pi0844), .S0(pi0955), .Y(po1000));
  MX2X1    g28856(.A(pi1043), .B(pi0845), .S0(pi0955), .Y(po1001));
  MX2X1    g28857(.A(pi0846), .B(pi1134), .S0(new_n27865_), .Y(po1002));
  MX2X1    g28858(.A(pi1055), .B(pi0847), .S0(pi0955), .Y(po1003));
  MX2X1    g28859(.A(pi1039), .B(pi0848), .S0(pi0955), .Y(po1004));
  MX2X1    g28860(.A(pi0849), .B(pi1198), .S0(new_n2720_), .Y(po1005));
  MX2X1    g28861(.A(pi1048), .B(pi0850), .S0(pi0955), .Y(po1006));
  MX2X1    g28862(.A(pi1045), .B(pi0851), .S0(pi0955), .Y(po1007));
  MX2X1    g28863(.A(pi1062), .B(pi0852), .S0(pi0955), .Y(po1008));
  MX2X1    g28864(.A(pi1080), .B(pi0853), .S0(pi0955), .Y(po1009));
  MX2X1    g28865(.A(pi1051), .B(pi0854), .S0(pi0955), .Y(po1010));
  MX2X1    g28866(.A(pi1065), .B(pi0855), .S0(pi0955), .Y(po1011));
  MX2X1    g28867(.A(pi1067), .B(pi0856), .S0(pi0955), .Y(po1012));
  MX2X1    g28868(.A(pi1058), .B(pi0857), .S0(pi0955), .Y(po1013));
  MX2X1    g28869(.A(pi1087), .B(pi0858), .S0(pi0955), .Y(po1014));
  MX2X1    g28870(.A(pi1070), .B(pi0859), .S0(pi0955), .Y(po1015));
  MX2X1    g28871(.A(pi1076), .B(pi0860), .S0(pi0955), .Y(po1016));
  MX2X1    g28872(.A(new_n3759_), .B(new_n3716_), .S0(new_n5032_), .Y(new_n31309_));
  NOR2X1   g28873(.A(pi1141), .B(pi0123), .Y(new_n31310_));
  OAI21X1  g28874(.A0(pi0861), .A1(new_n27864_), .B0(pi0228), .Y(new_n31311_));
  OAI22X1  g28875(.A0(new_n31311_), .A1(new_n31310_), .B0(new_n31309_), .B1(pi0228), .Y(po1017));
  MX2X1    g28876(.A(pi0862), .B(pi1139), .S0(new_n27865_), .Y(po1018));
  MX2X1    g28877(.A(pi0863), .B(pi1199), .S0(new_n2720_), .Y(po1019));
  MX2X1    g28878(.A(pi0864), .B(pi1197), .S0(new_n2720_), .Y(po1020));
  MX2X1    g28879(.A(pi1040), .B(pi0865), .S0(pi0955), .Y(po1021));
  MX2X1    g28880(.A(pi1053), .B(pi0866), .S0(pi0955), .Y(po1022));
  MX2X1    g28881(.A(pi1057), .B(pi0867), .S0(pi0955), .Y(po1023));
  MX2X1    g28882(.A(pi1063), .B(pi0868), .S0(pi0955), .Y(po1024));
  MX2X1    g28883(.A(new_n3908_), .B(new_n3866_), .S0(new_n5032_), .Y(new_n31320_));
  NOR2X1   g28884(.A(pi1140), .B(pi0123), .Y(new_n31321_));
  OAI21X1  g28885(.A0(pi0869), .A1(new_n27864_), .B0(pi0228), .Y(new_n31322_));
  OAI22X1  g28886(.A0(new_n31322_), .A1(new_n31321_), .B0(new_n31320_), .B1(pi0228), .Y(po1025));
  MX2X1    g28887(.A(pi1069), .B(pi0870), .S0(pi0955), .Y(po1026));
  MX2X1    g28888(.A(pi1072), .B(pi0871), .S0(pi0955), .Y(po1027));
  MX2X1    g28889(.A(pi1084), .B(pi0872), .S0(pi0955), .Y(po1028));
  MX2X1    g28890(.A(pi1044), .B(pi0873), .S0(pi0955), .Y(po1029));
  MX2X1    g28891(.A(pi1036), .B(pi0874), .S0(pi0955), .Y(po1030));
  MX2X1    g28892(.A(new_n4554_), .B(new_n4453_), .S0(new_n5032_), .Y(new_n31329_));
  OR2X1    g28893(.A(new_n4554_), .B(pi0123), .Y(new_n31330_));
  AOI21X1  g28894(.A0(pi0875), .A1(pi0123), .B0(new_n2793_), .Y(new_n31331_));
  AOI22X1  g28895(.A0(new_n31331_), .A1(new_n31330_), .B0(new_n31329_), .B1(new_n2793_), .Y(po1031));
  MX2X1    g28896(.A(pi1037), .B(pi0876), .S0(pi0955), .Y(po1032));
  MX2X1    g28897(.A(new_n4205_), .B(new_n4163_), .S0(new_n5032_), .Y(new_n31334_));
  NOR2X1   g28898(.A(pi1138), .B(pi0123), .Y(new_n31335_));
  OAI21X1  g28899(.A0(pi0877), .A1(new_n27864_), .B0(pi0228), .Y(new_n31336_));
  OAI22X1  g28900(.A0(new_n31336_), .A1(new_n31335_), .B0(new_n31334_), .B1(pi0228), .Y(po1033));
  MX2X1    g28901(.A(new_n4351_), .B(new_n4309_), .S0(new_n5032_), .Y(new_n31338_));
  NOR2X1   g28902(.A(pi1137), .B(pi0123), .Y(new_n31339_));
  OAI21X1  g28903(.A0(pi0878), .A1(new_n27864_), .B0(pi0228), .Y(new_n31340_));
  OAI22X1  g28904(.A0(new_n31340_), .A1(new_n31339_), .B0(new_n31338_), .B1(pi0228), .Y(po1034));
  MX2X1    g28905(.A(new_n4622_), .B(new_n4605_), .S0(new_n5032_), .Y(new_n31342_));
  NOR2X1   g28906(.A(pi1135), .B(pi0123), .Y(new_n31343_));
  OAI21X1  g28907(.A0(pi0879), .A1(new_n27864_), .B0(pi0228), .Y(new_n31344_));
  OAI22X1  g28908(.A0(new_n31344_), .A1(new_n31343_), .B0(new_n31342_), .B1(pi0228), .Y(po1035));
  MX2X1    g28909(.A(pi1081), .B(pi0880), .S0(pi0955), .Y(po1036));
  MX2X1    g28910(.A(pi1059), .B(pi0881), .S0(pi0955), .Y(po1037));
  INVX1    g28911(.A(pi0883), .Y(po1163));
  MX2X1    g28912(.A(pi1107), .B(po1163), .S0(new_n31220_), .Y(po1039));
  INVX1    g28913(.A(pi0884), .Y(po1180));
  MX2X1    g28914(.A(pi1124), .B(po1180), .S0(new_n31220_), .Y(po1040));
  INVX1    g28915(.A(pi0885), .Y(po1172));
  MX2X1    g28916(.A(pi1125), .B(po1172), .S0(new_n31220_), .Y(po1041));
  INVX1    g28917(.A(pi0886), .Y(po1166));
  MX2X1    g28918(.A(pi1109), .B(po1166), .S0(new_n31220_), .Y(po1042));
  INVX1    g28919(.A(pi0887), .Y(po1179));
  MX2X1    g28920(.A(pi1100), .B(po1179), .S0(new_n31220_), .Y(po1043));
  INVX1    g28921(.A(pi0888), .Y(po1164));
  MX2X1    g28922(.A(pi1120), .B(po1164), .S0(new_n31220_), .Y(po1044));
  INVX1    g28923(.A(pi0889), .Y(po1170));
  MX2X1    g28924(.A(pi1103), .B(po1170), .S0(new_n31220_), .Y(po1045));
  INVX1    g28925(.A(pi0890), .Y(po1153));
  MX2X1    g28926(.A(pi1126), .B(po1153), .S0(new_n31220_), .Y(po1046));
  INVX1    g28927(.A(pi0891), .Y(po1160));
  MX2X1    g28928(.A(pi1116), .B(po1160), .S0(new_n31220_), .Y(po1047));
  INVX1    g28929(.A(pi0892), .Y(po1183));
  MX2X1    g28930(.A(pi1101), .B(po1183), .S0(new_n31220_), .Y(po1048));
  INVX1    g28931(.A(pi0894), .Y(po1150));
  MX2X1    g28932(.A(pi1119), .B(po1150), .S0(new_n31220_), .Y(po1050));
  INVX1    g28933(.A(pi0895), .Y(po1168));
  MX2X1    g28934(.A(pi1113), .B(po1168), .S0(new_n31220_), .Y(po1051));
  INVX1    g28935(.A(pi0896), .Y(po1156));
  MX2X1    g28936(.A(pi1118), .B(po1156), .S0(new_n31220_), .Y(po1052));
  INVX1    g28937(.A(pi0898), .Y(po1176));
  MX2X1    g28938(.A(pi1129), .B(po1176), .S0(new_n31220_), .Y(po1054));
  INVX1    g28939(.A(pi0899), .Y(po1174));
  MX2X1    g28940(.A(pi1115), .B(po1174), .S0(new_n31220_), .Y(po1055));
  INVX1    g28941(.A(pi0900), .Y(po1171));
  MX2X1    g28942(.A(pi1110), .B(po1171), .S0(new_n31220_), .Y(po1056));
  INVX1    g28943(.A(pi0902), .Y(po1161));
  MX2X1    g28944(.A(pi1111), .B(po1161), .S0(new_n31220_), .Y(po1058));
  INVX1    g28945(.A(pi0903), .Y(po1162));
  MX2X1    g28946(.A(pi1121), .B(po1162), .S0(new_n31220_), .Y(po1059));
  INVX1    g28947(.A(pi0904), .Y(po1173));
  MX2X1    g28948(.A(pi1127), .B(po1173), .S0(new_n31220_), .Y(po1060));
  INVX1    g28949(.A(pi0905), .Y(po1151));
  MX2X1    g28950(.A(pi1131), .B(po1151), .S0(new_n31220_), .Y(po1061));
  INVX1    g28951(.A(pi0906), .Y(po1155));
  MX2X1    g28952(.A(pi1128), .B(po1155), .S0(new_n31220_), .Y(po1062));
  NOR2X1   g28953(.A(pi0979), .B(pi0624), .Y(new_n31390_));
  OAI21X1  g28954(.A0(new_n5026_), .A1(pi0598), .B0(pi0782), .Y(new_n31391_));
  OR2X1    g28955(.A(new_n31391_), .B(new_n31390_), .Y(new_n31392_));
  INVX1    g28956(.A(pi0782), .Y(new_n31393_));
  INVX1    g28957(.A(pi0615), .Y(new_n31394_));
  MX2X1    g28958(.A(new_n31394_), .B(pi0604), .S0(new_n5026_), .Y(new_n31395_));
  MX2X1    g28959(.A(new_n31395_), .B(pi0907), .S0(new_n31393_), .Y(new_n31396_));
  AND2X1   g28960(.A(new_n31396_), .B(new_n31392_), .Y(po1063));
  INVX1    g28961(.A(pi0908), .Y(po1159));
  MX2X1    g28962(.A(pi1122), .B(po1159), .S0(new_n31220_), .Y(po1064));
  INVX1    g28963(.A(pi0909), .Y(po1157));
  MX2X1    g28964(.A(pi1105), .B(po1157), .S0(new_n31220_), .Y(po1065));
  INVX1    g28965(.A(pi0910), .Y(po1181));
  MX2X1    g28966(.A(pi1117), .B(po1181), .S0(new_n31220_), .Y(po1066));
  INVX1    g28967(.A(pi0911), .Y(po1158));
  MX2X1    g28968(.A(pi1130), .B(po1158), .S0(new_n31220_), .Y(po1067));
  INVX1    g28969(.A(pi0912), .Y(po1167));
  MX2X1    g28970(.A(pi1114), .B(po1167), .S0(new_n31220_), .Y(po1068));
  INVX1    g28971(.A(pi0913), .Y(po1149));
  MX2X1    g28972(.A(pi1106), .B(po1149), .S0(new_n31220_), .Y(po1069));
  XOR2X1   g28973(.A(new_n30212_), .B(new_n4406_), .Y(po1070));
  INVX1    g28974(.A(pi0915), .Y(po1146));
  MX2X1    g28975(.A(pi1108), .B(po1146), .S0(new_n31220_), .Y(po1071));
  INVX1    g28976(.A(pi0916), .Y(po1169));
  MX2X1    g28977(.A(pi1123), .B(po1169), .S0(new_n31220_), .Y(po1072));
  INVX1    g28978(.A(pi0917), .Y(po1177));
  MX2X1    g28979(.A(pi1112), .B(po1177), .S0(new_n31220_), .Y(po1073));
  INVX1    g28980(.A(pi0918), .Y(po1175));
  MX2X1    g28981(.A(pi1104), .B(po1175), .S0(new_n31220_), .Y(po1074));
  INVX1    g28982(.A(pi0919), .Y(po1165));
  MX2X1    g28983(.A(pi1102), .B(po1165), .S0(new_n31220_), .Y(po1075));
  MX2X1    g28984(.A(pi0920), .B(pi1139), .S0(pi1093), .Y(po1076));
  MX2X1    g28985(.A(pi0921), .B(pi1140), .S0(pi1093), .Y(po1077));
  MX2X1    g28986(.A(pi0922), .B(pi1152), .S0(pi1093), .Y(po1078));
  MX2X1    g28987(.A(pi0923), .B(pi1154), .S0(pi1093), .Y(po1079));
  INVX1    g28988(.A(pi0311), .Y(new_n31425_));
  NOR4X1   g28989(.A(pi0312), .B(new_n31425_), .C(new_n28903_), .D(pi0300), .Y(po1080));
  MX2X1    g28990(.A(pi0925), .B(pi1155), .S0(pi1093), .Y(po1081));
  MX2X1    g28991(.A(pi0926), .B(pi1157), .S0(pi1093), .Y(po1082));
  MX2X1    g28992(.A(pi0927), .B(pi1145), .S0(pi1093), .Y(po1083));
  MX2X1    g28993(.A(pi0928), .B(pi1136), .S0(pi1093), .Y(po1084));
  MX2X1    g28994(.A(pi0929), .B(pi1144), .S0(pi1093), .Y(po1085));
  MX2X1    g28995(.A(pi0930), .B(pi1134), .S0(pi1093), .Y(po1086));
  MX2X1    g28996(.A(pi0931), .B(pi1150), .S0(pi1093), .Y(po1087));
  MX2X1    g28997(.A(pi0932), .B(pi1142), .S0(pi1093), .Y(po1088));
  MX2X1    g28998(.A(pi0933), .B(pi1137), .S0(pi1093), .Y(po1089));
  MX2X1    g28999(.A(pi0934), .B(pi1147), .S0(pi1093), .Y(po1090));
  MX2X1    g29000(.A(pi0935), .B(pi1141), .S0(pi1093), .Y(po1091));
  MX2X1    g29001(.A(pi0936), .B(pi1149), .S0(pi1093), .Y(po1092));
  MX2X1    g29002(.A(pi0937), .B(pi1148), .S0(pi1093), .Y(po1093));
  MX2X1    g29003(.A(pi0938), .B(pi1135), .S0(pi1093), .Y(po1094));
  MX2X1    g29004(.A(pi0939), .B(pi1146), .S0(pi1093), .Y(po1095));
  MX2X1    g29005(.A(pi0940), .B(pi1138), .S0(pi1093), .Y(po1096));
  MX2X1    g29006(.A(pi0941), .B(pi1153), .S0(pi1093), .Y(po1097));
  MX2X1    g29007(.A(pi0942), .B(pi1156), .S0(pi1093), .Y(po1098));
  MX2X1    g29008(.A(pi0943), .B(pi1151), .S0(pi1093), .Y(po1099));
  MX2X1    g29009(.A(pi0944), .B(pi1143), .S0(pi1093), .Y(po1100));
  AND3X1   g29010(.A(pi1093), .B(pi1092), .C(pi0230), .Y(po1102));
  OAI22X1  g29011(.A0(new_n31391_), .A1(new_n31390_), .B0(new_n5362_), .B1(pi0782), .Y(po1103));
  XOR2X1   g29012(.A(pi0992), .B(pi0266), .Y(po1104));
  INVX1    g29013(.A(pi0313), .Y(new_n31450_));
  MX2X1    g29014(.A(pi0949), .B(new_n31450_), .S0(po1110), .Y(po1105));
  NOR3X1   g29015(.A(new_n5967_), .B(new_n5024_), .C(new_n5237_), .Y(po1107));
  OAI21X1  g29016(.A0(new_n5024_), .A1(new_n2758_), .B0(new_n10074_), .Y(po1112));
  AND2X1   g29017(.A(pi0960), .B(new_n31393_), .Y(po1115));
  AND2X1   g29018(.A(pi0961), .B(new_n24814_), .Y(po1116));
  AND2X1   g29019(.A(pi0963), .B(new_n31393_), .Y(po1118));
  AND2X1   g29020(.A(pi0967), .B(new_n24814_), .Y(po1122));
  AND2X1   g29021(.A(pi0969), .B(new_n24814_), .Y(po1124));
  AND2X1   g29022(.A(pi0970), .B(new_n31393_), .Y(po1125));
  AND2X1   g29023(.A(pi0971), .B(new_n24814_), .Y(po1126));
  AND2X1   g29024(.A(pi0972), .B(new_n31393_), .Y(po1127));
  AND2X1   g29025(.A(pi0974), .B(new_n24814_), .Y(po1128));
  AND2X1   g29026(.A(pi0975), .B(new_n31393_), .Y(po1129));
  AND2X1   g29027(.A(pi0977), .B(new_n24814_), .Y(po1131));
  AND2X1   g29028(.A(pi0978), .B(new_n31393_), .Y(po1132));
  OR2X1    g29029(.A(new_n31394_), .B(pi0598), .Y(po1133));
  AND2X1   g29030(.A(pi1092), .B(pi0824), .Y(po1135));
  OR2X1    g29031(.A(pi0624), .B(pi0604), .Y(po1137));
  ONE      g29032(.Y(po0166));
  BUFX1    g29033(.A(pi0668), .Y(po0000));
  BUFX1    g29034(.A(pi0672), .Y(po0001));
  BUFX1    g29035(.A(pi0664), .Y(po0002));
  BUFX1    g29036(.A(pi0667), .Y(po0003));
  BUFX1    g29037(.A(pi0676), .Y(po0004));
  BUFX1    g29038(.A(pi0673), .Y(po0005));
  BUFX1    g29039(.A(pi0675), .Y(po0006));
  BUFX1    g29040(.A(pi0666), .Y(po0007));
  BUFX1    g29041(.A(pi0679), .Y(po0008));
  BUFX1    g29042(.A(pi0674), .Y(po0009));
  BUFX1    g29043(.A(pi0663), .Y(po0010));
  BUFX1    g29044(.A(pi0670), .Y(po0011));
  BUFX1    g29045(.A(pi0677), .Y(po0012));
  BUFX1    g29046(.A(pi0682), .Y(po0013));
  BUFX1    g29047(.A(pi0671), .Y(po0014));
  BUFX1    g29048(.A(pi0678), .Y(po0015));
  BUFX1    g29049(.A(pi0718), .Y(po0016));
  BUFX1    g29050(.A(pi0707), .Y(po0017));
  BUFX1    g29051(.A(pi0708), .Y(po0018));
  BUFX1    g29052(.A(pi0713), .Y(po0019));
  BUFX1    g29053(.A(pi0711), .Y(po0020));
  BUFX1    g29054(.A(pi0716), .Y(po0021));
  BUFX1    g29055(.A(pi0733), .Y(po0022));
  BUFX1    g29056(.A(pi0712), .Y(po0023));
  BUFX1    g29057(.A(pi0689), .Y(po0024));
  BUFX1    g29058(.A(pi0717), .Y(po0025));
  BUFX1    g29059(.A(pi0692), .Y(po0026));
  BUFX1    g29060(.A(pi0719), .Y(po0027));
  BUFX1    g29061(.A(pi0722), .Y(po0028));
  BUFX1    g29062(.A(pi0714), .Y(po0029));
  BUFX1    g29063(.A(pi0720), .Y(po0030));
  BUFX1    g29064(.A(pi0685), .Y(po0031));
  BUFX1    g29065(.A(pi0837), .Y(po0032));
  BUFX1    g29066(.A(pi0850), .Y(po0033));
  BUFX1    g29067(.A(pi0872), .Y(po0034));
  BUFX1    g29068(.A(pi0871), .Y(po0035));
  BUFX1    g29069(.A(pi0881), .Y(po0036));
  BUFX1    g29070(.A(pi0866), .Y(po0037));
  BUFX1    g29071(.A(pi0876), .Y(po0038));
  BUFX1    g29072(.A(pi0873), .Y(po0039));
  BUFX1    g29073(.A(pi0874), .Y(po0040));
  BUFX1    g29074(.A(pi0859), .Y(po0041));
  BUFX1    g29075(.A(pi0855), .Y(po0042));
  BUFX1    g29076(.A(pi0852), .Y(po0043));
  BUFX1    g29077(.A(pi0870), .Y(po0044));
  BUFX1    g29078(.A(pi0848), .Y(po0045));
  BUFX1    g29079(.A(pi0865), .Y(po0046));
  BUFX1    g29080(.A(pi0856), .Y(po0047));
  BUFX1    g29081(.A(pi0853), .Y(po0048));
  BUFX1    g29082(.A(pi0847), .Y(po0049));
  BUFX1    g29083(.A(pi0857), .Y(po0050));
  BUFX1    g29084(.A(pi0854), .Y(po0051));
  BUFX1    g29085(.A(pi0858), .Y(po0052));
  BUFX1    g29086(.A(pi0845), .Y(po0053));
  BUFX1    g29087(.A(pi0838), .Y(po0054));
  BUFX1    g29088(.A(pi0842), .Y(po0055));
  BUFX1    g29089(.A(pi0843), .Y(po0056));
  BUFX1    g29090(.A(pi0839), .Y(po0057));
  BUFX1    g29091(.A(pi0844), .Y(po0058));
  BUFX1    g29092(.A(pi0868), .Y(po0059));
  BUFX1    g29093(.A(pi0851), .Y(po0060));
  BUFX1    g29094(.A(pi0867), .Y(po0061));
  BUFX1    g29095(.A(pi0880), .Y(po0062));
  BUFX1    g29096(.A(pi0860), .Y(po0063));
  BUFX1    g29097(.A(pi1030), .Y(po0064));
  BUFX1    g29098(.A(pi1034), .Y(po0065));
  BUFX1    g29099(.A(pi1015), .Y(po0066));
  BUFX1    g29100(.A(pi1020), .Y(po0067));
  BUFX1    g29101(.A(pi1025), .Y(po0068));
  BUFX1    g29102(.A(pi1005), .Y(po0069));
  BUFX1    g29103(.A(pi0996), .Y(po0070));
  BUFX1    g29104(.A(pi1012), .Y(po0071));
  BUFX1    g29105(.A(pi0993), .Y(po0072));
  BUFX1    g29106(.A(pi1016), .Y(po0073));
  BUFX1    g29107(.A(pi1021), .Y(po0074));
  BUFX1    g29108(.A(pi1010), .Y(po0075));
  BUFX1    g29109(.A(pi1027), .Y(po0076));
  BUFX1    g29110(.A(pi1018), .Y(po0077));
  BUFX1    g29111(.A(pi1017), .Y(po0078));
  BUFX1    g29112(.A(pi1024), .Y(po0079));
  BUFX1    g29113(.A(pi1009), .Y(po0080));
  BUFX1    g29114(.A(pi1032), .Y(po0081));
  BUFX1    g29115(.A(pi1003), .Y(po0082));
  BUFX1    g29116(.A(pi0997), .Y(po0083));
  BUFX1    g29117(.A(pi1013), .Y(po0084));
  BUFX1    g29118(.A(pi1011), .Y(po0085));
  BUFX1    g29119(.A(pi1008), .Y(po0086));
  BUFX1    g29120(.A(pi1019), .Y(po0087));
  BUFX1    g29121(.A(pi1031), .Y(po0088));
  BUFX1    g29122(.A(pi1022), .Y(po0089));
  BUFX1    g29123(.A(pi1000), .Y(po0090));
  BUFX1    g29124(.A(pi1023), .Y(po0091));
  BUFX1    g29125(.A(pi1002), .Y(po0092));
  BUFX1    g29126(.A(pi1026), .Y(po0093));
  BUFX1    g29127(.A(pi1006), .Y(po0094));
  BUFX1    g29128(.A(pi0998), .Y(po0095));
  BUFX1    g29129(.A(pi0031), .Y(po0096));
  BUFX1    g29130(.A(pi0080), .Y(po0097));
  BUFX1    g29131(.A(pi0893), .Y(po0098));
  BUFX1    g29132(.A(pi0467), .Y(po0099));
  BUFX1    g29133(.A(pi0078), .Y(po0100));
  BUFX1    g29134(.A(pi0112), .Y(po0101));
  BUFX1    g29135(.A(pi0013), .Y(po0102));
  BUFX1    g29136(.A(pi0025), .Y(po0103));
  BUFX1    g29137(.A(pi0226), .Y(po0104));
  BUFX1    g29138(.A(pi0127), .Y(po0105));
  BUFX1    g29139(.A(pi0822), .Y(po0106));
  BUFX1    g29140(.A(pi0808), .Y(po0107));
  BUFX1    g29141(.A(pi0227), .Y(po0108));
  BUFX1    g29142(.A(pi0477), .Y(po0109));
  BUFX1    g29143(.A(pi0834), .Y(po0110));
  BUFX1    g29144(.A(pi0229), .Y(po0111));
  BUFX1    g29145(.A(pi0012), .Y(po0112));
  BUFX1    g29146(.A(pi0011), .Y(po0113));
  BUFX1    g29147(.A(pi0010), .Y(po0114));
  BUFX1    g29148(.A(pi0009), .Y(po0115));
  BUFX1    g29149(.A(pi0008), .Y(po0116));
  BUFX1    g29150(.A(pi0007), .Y(po0117));
  BUFX1    g29151(.A(pi0006), .Y(po0118));
  BUFX1    g29152(.A(pi0005), .Y(po0119));
  BUFX1    g29153(.A(pi0004), .Y(po0120));
  BUFX1    g29154(.A(pi0003), .Y(po0121));
  BUFX1    g29155(.A(pi0000), .Y(po0122));
  BUFX1    g29156(.A(pi0002), .Y(po0123));
  BUFX1    g29157(.A(pi0001), .Y(po0124));
  BUFX1    g29158(.A(pi0310), .Y(po0125));
  BUFX1    g29159(.A(pi0302), .Y(po0126));
  BUFX1    g29160(.A(pi0475), .Y(po0127));
  BUFX1    g29161(.A(pi0474), .Y(po0128));
  BUFX1    g29162(.A(pi0466), .Y(po0129));
  BUFX1    g29163(.A(pi0473), .Y(po0130));
  BUFX1    g29164(.A(pi0471), .Y(po0131));
  BUFX1    g29165(.A(pi0472), .Y(po0132));
  BUFX1    g29166(.A(pi0470), .Y(po0133));
  BUFX1    g29167(.A(pi0469), .Y(po0134));
  BUFX1    g29168(.A(pi0465), .Y(po0135));
  BUFX1    g29169(.A(pi1028), .Y(po0136));
  BUFX1    g29170(.A(pi1033), .Y(po0137));
  BUFX1    g29171(.A(pi0995), .Y(po0138));
  BUFX1    g29172(.A(pi0994), .Y(po0139));
  BUFX1    g29173(.A(pi0028), .Y(po0140));
  BUFX1    g29174(.A(pi0027), .Y(po0141));
  BUFX1    g29175(.A(pi0026), .Y(po0142));
  BUFX1    g29176(.A(pi0029), .Y(po0143));
  BUFX1    g29177(.A(pi0015), .Y(po0144));
  BUFX1    g29178(.A(pi0014), .Y(po0145));
  BUFX1    g29179(.A(pi0021), .Y(po0146));
  BUFX1    g29180(.A(pi0020), .Y(po0147));
  BUFX1    g29181(.A(pi0019), .Y(po0148));
  BUFX1    g29182(.A(pi0018), .Y(po0149));
  BUFX1    g29183(.A(pi0017), .Y(po0150));
  BUFX1    g29184(.A(pi0016), .Y(po0151));
  BUFX1    g29185(.A(pi1096), .Y(po0152));
  BUFX1    g29186(.A(pi0228), .Y(po0168));
  BUFX1    g29187(.A(pi0022), .Y(po0169));
  BUFX1    g29188(.A(pi1089), .Y(po0179));
  BUFX1    g29189(.A(pi0023), .Y(po0180));
  MX2X1    g29190(.A(new_n5099_), .B(new_n4978_), .S0(pi0057), .Y(po0181));
  BUFX1    g29191(.A(pi0037), .Y(po0188));
  BUFX1    g29192(.A(pi0117), .Y(po0263));
  BUFX1    g29193(.A(pi0131), .Y(po0285));
  BUFX1    g29194(.A(pi0232), .Y(po0386));
  BUFX1    g29195(.A(pi0236), .Y(po0388));
  BUFX1    g29196(.A(pi0583), .Y(po0636));
  BUFX1    g29197(.A(pi0067), .Y(po1053));
  BUFX1    g29198(.A(pi1134), .Y(po1108));
  BUFX1    g29199(.A(pi0964), .Y(po1109));
  BUFX1    g29200(.A(pi0965), .Y(po1111));
  BUFX1    g29201(.A(pi0991), .Y(po1113));
  BUFX1    g29202(.A(pi0985), .Y(po1114));
  BUFX1    g29203(.A(pi1014), .Y(po1117));
  BUFX1    g29204(.A(pi1029), .Y(po1119));
  BUFX1    g29205(.A(pi1004), .Y(po1120));
  BUFX1    g29206(.A(pi1007), .Y(po1121));
  BUFX1    g29207(.A(pi1135), .Y(po1123));
  BUFX1    g29208(.A(pi1064), .Y(po1134));
  BUFX1    g29209(.A(pi0299), .Y(po1136));
  BUFX1    g29210(.A(pi1075), .Y(po1138));
  BUFX1    g29211(.A(pi1052), .Y(po1139));
  BUFX1    g29212(.A(pi0771), .Y(po1140));
  BUFX1    g29213(.A(pi0765), .Y(po1141));
  BUFX1    g29214(.A(pi0605), .Y(po1142));
  BUFX1    g29215(.A(pi0601), .Y(po1143));
  BUFX1    g29216(.A(pi0278), .Y(po1144));
  BUFX1    g29217(.A(pi0279), .Y(po1145));
  BUFX1    g29218(.A(pi1095), .Y(po1152));
  BUFX1    g29219(.A(pi1094), .Y(po1154));
  BUFX1    g29220(.A(pi1187), .Y(po1184));
  BUFX1    g29221(.A(pi1172), .Y(po1185));
  BUFX1    g29222(.A(pi1170), .Y(po1186));
  BUFX1    g29223(.A(pi1138), .Y(po1187));
  BUFX1    g29224(.A(pi1177), .Y(po1188));
  BUFX1    g29225(.A(pi1178), .Y(po1189));
  BUFX1    g29226(.A(pi0863), .Y(po1190));
  BUFX1    g29227(.A(pi1203), .Y(po1191));
  BUFX1    g29228(.A(pi1185), .Y(po1192));
  BUFX1    g29229(.A(pi1171), .Y(po1193));
  BUFX1    g29230(.A(pi1192), .Y(po1194));
  BUFX1    g29231(.A(pi1137), .Y(po1195));
  BUFX1    g29232(.A(pi1186), .Y(po1196));
  BUFX1    g29233(.A(pi1165), .Y(po1197));
  BUFX1    g29234(.A(pi1164), .Y(po1198));
  BUFX1    g29235(.A(pi1098), .Y(po1199));
  BUFX1    g29236(.A(pi1183), .Y(po1200));
  BUFX1    g29237(.A(pi0230), .Y(po1201));
  BUFX1    g29238(.A(pi1169), .Y(po1202));
  BUFX1    g29239(.A(pi1136), .Y(po1203));
  BUFX1    g29240(.A(pi1181), .Y(po1204));
  BUFX1    g29241(.A(pi0849), .Y(po1205));
  BUFX1    g29242(.A(pi1193), .Y(po1206));
  BUFX1    g29243(.A(pi1182), .Y(po1207));
  BUFX1    g29244(.A(pi1168), .Y(po1208));
  BUFX1    g29245(.A(pi1175), .Y(po1209));
  BUFX1    g29246(.A(pi1191), .Y(po1210));
  BUFX1    g29247(.A(pi1099), .Y(po1211));
  BUFX1    g29248(.A(pi1174), .Y(po1212));
  BUFX1    g29249(.A(pi1179), .Y(po1213));
  BUFX1    g29250(.A(pi1202), .Y(po1214));
  BUFX1    g29251(.A(pi1176), .Y(po1215));
  BUFX1    g29252(.A(pi1173), .Y(po1216));
  BUFX1    g29253(.A(pi1201), .Y(po1217));
  BUFX1    g29254(.A(pi1167), .Y(po1218));
  BUFX1    g29255(.A(pi0840), .Y(po1219));
  BUFX1    g29256(.A(pi1189), .Y(po1220));
  BUFX1    g29257(.A(pi1195), .Y(po1221));
  BUFX1    g29258(.A(pi0864), .Y(po1222));
  BUFX1    g29259(.A(pi1190), .Y(po1223));
  BUFX1    g29260(.A(pi1188), .Y(po1224));
  BUFX1    g29261(.A(pi1180), .Y(po1225));
  BUFX1    g29262(.A(pi1194), .Y(po1226));
  BUFX1    g29263(.A(pi1097), .Y(po1227));
  BUFX1    g29264(.A(pi1166), .Y(po1228));
  BUFX1    g29265(.A(pi1200), .Y(po1229));
  BUFX1    g29266(.A(pi1184), .Y(po1230));
endmodule


