// Benchmark "top" written by ABC on Mon Sep 21 03:42:41 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ;
  output \sin[0] , \sin[1] , \sin[2] , \sin[3] , \sin[4] , \sin[5] , \sin[6] ,
    \sin[7] , \sin[8] , \sin[9] , \sin[10] , \sin[11] , \sin[12] ,
    \sin[13] , \sin[14] , \sin[15] , \sin[16] , \sin[17] , \sin[18] ,
    \sin[19] , \sin[20] , \sin[21] , \sin[22] , \sin[23] , \sin[24] ;
  wire new_n50_, new_n51_, new_n52_, new_n53_, new_n54_, new_n55_, new_n56_,
    new_n57_, new_n58_, new_n59_, new_n60_, new_n61_, new_n62_, new_n63_,
    new_n64_, new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_,
    new_n71_, new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_,
    new_n78_, new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_,
    new_n85_, new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_,
    new_n92_, new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_,
    new_n99_, new_n100_, new_n101_, new_n102_, new_n103_, new_n104_,
    new_n105_, new_n106_, new_n107_, new_n108_, new_n109_, new_n110_,
    new_n111_, new_n112_, new_n113_, new_n114_, new_n115_, new_n116_,
    new_n117_, new_n118_, new_n119_, new_n120_, new_n121_, new_n122_,
    new_n123_, new_n124_, new_n125_, new_n126_, new_n127_, new_n128_,
    new_n129_, new_n130_, new_n131_, new_n132_, new_n133_, new_n134_,
    new_n135_, new_n136_, new_n137_, new_n138_, new_n139_, new_n140_,
    new_n141_, new_n142_, new_n143_, new_n144_, new_n145_, new_n146_,
    new_n147_, new_n148_, new_n149_, new_n150_, new_n151_, new_n152_,
    new_n153_, new_n154_, new_n155_, new_n156_, new_n157_, new_n158_,
    new_n159_, new_n160_, new_n161_, new_n162_, new_n163_, new_n164_,
    new_n165_, new_n166_, new_n167_, new_n168_, new_n169_, new_n170_,
    new_n171_, new_n172_, new_n173_, new_n174_, new_n175_, new_n176_,
    new_n177_, new_n178_, new_n179_, new_n180_, new_n181_, new_n182_,
    new_n183_, new_n184_, new_n185_, new_n186_, new_n187_, new_n188_,
    new_n189_, new_n190_, new_n191_, new_n192_, new_n193_, new_n194_,
    new_n195_, new_n196_, new_n197_, new_n198_, new_n199_, new_n200_,
    new_n201_, new_n202_, new_n203_, new_n204_, new_n205_, new_n206_,
    new_n207_, new_n208_, new_n209_, new_n210_, new_n211_, new_n212_,
    new_n213_, new_n214_, new_n215_, new_n216_, new_n217_, new_n218_,
    new_n219_, new_n220_, new_n221_, new_n222_, new_n223_, new_n224_,
    new_n225_, new_n226_, new_n227_, new_n228_, new_n229_, new_n230_,
    new_n231_, new_n232_, new_n233_, new_n234_, new_n235_, new_n236_,
    new_n237_, new_n238_, new_n239_, new_n240_, new_n241_, new_n242_,
    new_n243_, new_n244_, new_n245_, new_n246_, new_n247_, new_n248_,
    new_n249_, new_n250_, new_n251_, new_n252_, new_n253_, new_n254_,
    new_n255_, new_n256_, new_n257_, new_n258_, new_n259_, new_n260_,
    new_n261_, new_n262_, new_n263_, new_n264_, new_n265_, new_n266_,
    new_n267_, new_n268_, new_n269_, new_n270_, new_n271_, new_n272_,
    new_n273_, new_n274_, new_n275_, new_n276_, new_n277_, new_n278_,
    new_n279_, new_n280_, new_n281_, new_n282_, new_n283_, new_n284_,
    new_n285_, new_n286_, new_n287_, new_n288_, new_n289_, new_n290_,
    new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n325_, new_n326_,
    new_n327_, new_n328_, new_n329_, new_n330_, new_n331_, new_n332_,
    new_n333_, new_n334_, new_n335_, new_n336_, new_n337_, new_n338_,
    new_n339_, new_n340_, new_n341_, new_n342_, new_n343_, new_n344_,
    new_n345_, new_n346_, new_n347_, new_n348_, new_n349_, new_n350_,
    new_n351_, new_n352_, new_n353_, new_n354_, new_n355_, new_n356_,
    new_n357_, new_n358_, new_n359_, new_n360_, new_n361_, new_n362_,
    new_n363_, new_n364_, new_n365_, new_n366_, new_n367_, new_n368_,
    new_n369_, new_n370_, new_n371_, new_n372_, new_n373_, new_n374_,
    new_n375_, new_n376_, new_n377_, new_n378_, new_n379_, new_n380_,
    new_n381_, new_n382_, new_n383_, new_n384_, new_n385_, new_n386_,
    new_n387_, new_n388_, new_n389_, new_n390_, new_n391_, new_n392_,
    new_n393_, new_n394_, new_n395_, new_n396_, new_n397_, new_n398_,
    new_n399_, new_n400_, new_n401_, new_n402_, new_n403_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n408_, new_n409_, new_n410_,
    new_n411_, new_n412_, new_n413_, new_n414_, new_n415_, new_n416_,
    new_n417_, new_n418_, new_n419_, new_n420_, new_n421_, new_n422_,
    new_n423_, new_n424_, new_n425_, new_n426_, new_n427_, new_n428_,
    new_n429_, new_n430_, new_n431_, new_n432_, new_n433_, new_n434_,
    new_n435_, new_n436_, new_n437_, new_n438_, new_n439_, new_n440_,
    new_n441_, new_n442_, new_n443_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n448_, new_n449_, new_n450_, new_n451_, new_n452_,
    new_n453_, new_n454_, new_n455_, new_n456_, new_n457_, new_n458_,
    new_n459_, new_n460_, new_n461_, new_n462_, new_n463_, new_n464_,
    new_n465_, new_n466_, new_n467_, new_n468_, new_n469_, new_n470_,
    new_n471_, new_n472_, new_n473_, new_n474_, new_n475_, new_n476_,
    new_n477_, new_n478_, new_n479_, new_n480_, new_n481_, new_n482_,
    new_n483_, new_n484_, new_n485_, new_n486_, new_n487_, new_n488_,
    new_n489_, new_n490_, new_n491_, new_n492_, new_n493_, new_n494_,
    new_n495_, new_n496_, new_n497_, new_n498_, new_n499_, new_n500_,
    new_n501_, new_n502_, new_n503_, new_n504_, new_n505_, new_n506_,
    new_n507_, new_n508_, new_n509_, new_n510_, new_n511_, new_n512_,
    new_n513_, new_n514_, new_n515_, new_n516_, new_n517_, new_n518_,
    new_n519_, new_n520_, new_n521_, new_n522_, new_n523_, new_n524_,
    new_n525_, new_n526_, new_n527_, new_n528_, new_n529_, new_n530_,
    new_n531_, new_n532_, new_n533_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n551_, new_n552_, new_n553_, new_n554_,
    new_n555_, new_n556_, new_n557_, new_n558_, new_n559_, new_n560_,
    new_n561_, new_n562_, new_n563_, new_n564_, new_n565_, new_n566_,
    new_n567_, new_n568_, new_n569_, new_n570_, new_n571_, new_n572_,
    new_n573_, new_n574_, new_n575_, new_n576_, new_n577_, new_n578_,
    new_n579_, new_n580_, new_n581_, new_n582_, new_n583_, new_n584_,
    new_n585_, new_n586_, new_n587_, new_n588_, new_n589_, new_n590_,
    new_n591_, new_n592_, new_n593_, new_n594_, new_n595_, new_n596_,
    new_n597_, new_n598_, new_n599_, new_n600_, new_n601_, new_n602_,
    new_n603_, new_n604_, new_n605_, new_n606_, new_n607_, new_n608_,
    new_n609_, new_n610_, new_n611_, new_n612_, new_n613_, new_n614_,
    new_n615_, new_n616_, new_n617_, new_n618_, new_n619_, new_n620_,
    new_n621_, new_n622_, new_n623_, new_n624_, new_n625_, new_n626_,
    new_n627_, new_n628_, new_n629_, new_n630_, new_n631_, new_n632_,
    new_n633_, new_n634_, new_n635_, new_n636_, new_n637_, new_n638_,
    new_n639_, new_n640_, new_n641_, new_n642_, new_n643_, new_n644_,
    new_n645_, new_n646_, new_n647_, new_n648_, new_n649_, new_n650_,
    new_n651_, new_n652_, new_n653_, new_n654_, new_n655_, new_n656_,
    new_n657_, new_n658_, new_n659_, new_n660_, new_n661_, new_n662_,
    new_n663_, new_n664_, new_n665_, new_n666_, new_n667_, new_n668_,
    new_n669_, new_n670_, new_n671_, new_n672_, new_n673_, new_n674_,
    new_n675_, new_n676_, new_n677_, new_n678_, new_n679_, new_n680_,
    new_n681_, new_n682_, new_n683_, new_n684_, new_n685_, new_n686_,
    new_n687_, new_n688_, new_n689_, new_n690_, new_n691_, new_n692_,
    new_n693_, new_n694_, new_n695_, new_n696_, new_n697_, new_n698_,
    new_n699_, new_n700_, new_n701_, new_n702_, new_n703_, new_n704_,
    new_n705_, new_n706_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n718_, new_n719_, new_n720_, new_n721_, new_n722_,
    new_n723_, new_n724_, new_n725_, new_n726_, new_n727_, new_n728_,
    new_n729_, new_n730_, new_n731_, new_n732_, new_n733_, new_n734_,
    new_n735_, new_n736_, new_n737_, new_n738_, new_n739_, new_n740_,
    new_n741_, new_n742_, new_n743_, new_n744_, new_n745_, new_n746_,
    new_n747_, new_n748_, new_n749_, new_n750_, new_n751_, new_n752_,
    new_n753_, new_n754_, new_n755_, new_n756_, new_n757_, new_n758_,
    new_n759_, new_n760_, new_n761_, new_n762_, new_n763_, new_n764_,
    new_n765_, new_n766_, new_n767_, new_n768_, new_n769_, new_n770_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n782_,
    new_n783_, new_n784_, new_n785_, new_n786_, new_n787_, new_n788_,
    new_n789_, new_n790_, new_n791_, new_n792_, new_n793_, new_n794_,
    new_n795_, new_n796_, new_n797_, new_n798_, new_n799_, new_n800_,
    new_n801_, new_n802_, new_n803_, new_n804_, new_n805_, new_n806_,
    new_n807_, new_n808_, new_n809_, new_n810_, new_n811_, new_n812_,
    new_n813_, new_n814_, new_n815_, new_n816_, new_n817_, new_n818_,
    new_n819_, new_n820_, new_n821_, new_n822_, new_n823_, new_n824_,
    new_n825_, new_n826_, new_n827_, new_n828_, new_n829_, new_n830_,
    new_n831_, new_n832_, new_n833_, new_n834_, new_n835_, new_n836_,
    new_n837_, new_n838_, new_n839_, new_n840_, new_n841_, new_n842_,
    new_n843_, new_n844_, new_n845_, new_n846_, new_n847_, new_n848_,
    new_n849_, new_n850_, new_n851_, new_n852_, new_n853_, new_n854_,
    new_n855_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n868_, new_n869_, new_n870_, new_n871_, new_n872_,
    new_n873_, new_n874_, new_n875_, new_n876_, new_n877_, new_n878_,
    new_n879_, new_n880_, new_n881_, new_n882_, new_n883_, new_n884_,
    new_n885_, new_n886_, new_n887_, new_n888_, new_n889_, new_n890_,
    new_n891_, new_n892_, new_n893_, new_n894_, new_n895_, new_n896_,
    new_n897_, new_n898_, new_n899_, new_n900_, new_n901_, new_n902_,
    new_n903_, new_n904_, new_n905_, new_n906_, new_n907_, new_n908_,
    new_n909_, new_n910_, new_n911_, new_n912_, new_n913_, new_n914_,
    new_n915_, new_n916_, new_n917_, new_n918_, new_n919_, new_n920_,
    new_n921_, new_n922_, new_n923_, new_n924_, new_n925_, new_n926_,
    new_n927_, new_n928_, new_n929_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n938_,
    new_n939_, new_n940_, new_n941_, new_n942_, new_n943_, new_n944_,
    new_n945_, new_n946_, new_n947_, new_n948_, new_n949_, new_n950_,
    new_n951_, new_n952_, new_n953_, new_n954_, new_n955_, new_n956_,
    new_n957_, new_n958_, new_n959_, new_n960_, new_n961_, new_n962_,
    new_n963_, new_n964_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n971_, new_n972_, new_n973_, new_n974_,
    new_n975_, new_n976_, new_n977_, new_n978_, new_n979_, new_n980_,
    new_n981_, new_n982_, new_n983_, new_n984_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n991_, new_n992_,
    new_n993_, new_n994_, new_n995_, new_n996_, new_n997_, new_n998_,
    new_n999_, new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_,
    new_n1005_, new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_,
    new_n1011_, new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_,
    new_n1017_, new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_,
    new_n1035_, new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_,
    new_n1041_, new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_,
    new_n1047_, new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_,
    new_n1053_, new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_,
    new_n1059_, new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_,
    new_n1065_, new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_,
    new_n1071_, new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_,
    new_n1077_, new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_,
    new_n1083_, new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_,
    new_n1089_, new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_,
    new_n1095_, new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_,
    new_n1101_, new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_,
    new_n1107_, new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_,
    new_n1113_, new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_,
    new_n1119_, new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_,
    new_n1125_, new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_,
    new_n1131_, new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_,
    new_n1137_, new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_,
    new_n1143_, new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_,
    new_n1149_, new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_,
    new_n1155_, new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_,
    new_n1161_, new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_,
    new_n1167_, new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_,
    new_n1173_, new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_,
    new_n1179_, new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_,
    new_n1185_, new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_,
    new_n1191_, new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_,
    new_n1197_, new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_,
    new_n1203_, new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_,
    new_n1209_, new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_,
    new_n1215_, new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_,
    new_n1221_, new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_,
    new_n1227_, new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_,
    new_n1233_, new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_,
    new_n1239_, new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_,
    new_n1245_, new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_,
    new_n1251_, new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_,
    new_n1257_, new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_,
    new_n1263_, new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_,
    new_n1269_, new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_,
    new_n1275_, new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_,
    new_n1281_, new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_,
    new_n1287_, new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_,
    new_n1293_, new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_,
    new_n1299_, new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_,
    new_n1305_, new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_,
    new_n1311_, new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_,
    new_n1317_, new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_,
    new_n1323_, new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_,
    new_n1329_, new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_,
    new_n1335_, new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_,
    new_n1341_, new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_,
    new_n1347_, new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_,
    new_n1353_, new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_,
    new_n1359_, new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_,
    new_n1365_, new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_,
    new_n1371_, new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_,
    new_n1377_, new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_,
    new_n1383_, new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_,
    new_n1389_, new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_,
    new_n1395_, new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_,
    new_n1401_, new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_,
    new_n1407_, new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_,
    new_n1413_, new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_,
    new_n1419_, new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_,
    new_n1425_, new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_,
    new_n1431_, new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_,
    new_n1437_, new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_,
    new_n1443_, new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_,
    new_n1449_, new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_,
    new_n1455_, new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_,
    new_n1461_, new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_,
    new_n1467_, new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_,
    new_n1473_, new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_,
    new_n1479_, new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_,
    new_n1485_, new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_,
    new_n1491_, new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_,
    new_n1497_, new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_,
    new_n1503_, new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_,
    new_n1509_, new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_,
    new_n1515_, new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_,
    new_n1521_, new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_,
    new_n1527_, new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_,
    new_n1533_, new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_,
    new_n1539_, new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_,
    new_n1545_, new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_,
    new_n1551_, new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_,
    new_n1557_, new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_,
    new_n1563_, new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_,
    new_n1569_, new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_,
    new_n1575_, new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_,
    new_n1581_, new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_,
    new_n1587_, new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_,
    new_n1593_, new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_,
    new_n1599_, new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_,
    new_n1605_, new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_,
    new_n1611_, new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_,
    new_n1617_, new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_,
    new_n1623_, new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_,
    new_n1629_, new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_,
    new_n1635_, new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_,
    new_n1641_, new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_,
    new_n1647_, new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_,
    new_n1653_, new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_,
    new_n1659_, new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_,
    new_n1665_, new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_,
    new_n1671_, new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_,
    new_n1677_, new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_,
    new_n1683_, new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_,
    new_n1689_, new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_,
    new_n1695_, new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_,
    new_n1701_, new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_,
    new_n1707_, new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_,
    new_n1713_, new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_,
    new_n1719_, new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_,
    new_n1725_, new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_,
    new_n1731_, new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_,
    new_n1737_, new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_,
    new_n1743_, new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_,
    new_n1749_, new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_,
    new_n1755_, new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_,
    new_n1761_, new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_,
    new_n1767_, new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_,
    new_n1773_, new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_,
    new_n1779_, new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_,
    new_n1785_, new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_,
    new_n1791_, new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_,
    new_n1797_, new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_,
    new_n1803_, new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_,
    new_n1809_, new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_,
    new_n1815_, new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_,
    new_n1821_, new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_,
    new_n1827_, new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_,
    new_n1833_, new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_,
    new_n1839_, new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_,
    new_n1845_, new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_,
    new_n1851_, new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_,
    new_n1857_, new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_,
    new_n1863_, new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_,
    new_n1869_, new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_,
    new_n1875_, new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_,
    new_n1881_, new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_,
    new_n1887_, new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_,
    new_n1893_, new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_,
    new_n1899_, new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_,
    new_n1905_, new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_,
    new_n1911_, new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_,
    new_n1917_, new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_,
    new_n1923_, new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_,
    new_n1929_, new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_,
    new_n1935_, new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_,
    new_n1941_, new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_,
    new_n1947_, new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_,
    new_n1953_, new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_,
    new_n1959_, new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_,
    new_n1965_, new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_,
    new_n1971_, new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_,
    new_n1977_, new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_,
    new_n1983_, new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_,
    new_n1989_, new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_,
    new_n1995_, new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_,
    new_n2001_, new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_,
    new_n2007_, new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_,
    new_n2013_, new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_,
    new_n2019_, new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_,
    new_n2025_, new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_,
    new_n2031_, new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_,
    new_n2037_, new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_,
    new_n2043_, new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_,
    new_n2049_, new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_,
    new_n2055_, new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_,
    new_n2061_, new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_,
    new_n2067_, new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_,
    new_n2073_, new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_,
    new_n2079_, new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_,
    new_n2085_, new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_,
    new_n2091_, new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_,
    new_n2097_, new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_,
    new_n2103_, new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_,
    new_n2109_, new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_,
    new_n2115_, new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_,
    new_n2121_, new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_,
    new_n2127_, new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_,
    new_n2133_, new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_,
    new_n2139_, new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_,
    new_n2145_, new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_,
    new_n2151_, new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_,
    new_n2157_, new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_,
    new_n2163_, new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_,
    new_n2169_, new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_,
    new_n2175_, new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_,
    new_n2181_, new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_,
    new_n2187_, new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_,
    new_n2193_, new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_,
    new_n2199_, new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_,
    new_n2205_, new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_,
    new_n2211_, new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_,
    new_n2217_, new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_,
    new_n2223_, new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_,
    new_n2229_, new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_,
    new_n2235_, new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_,
    new_n2241_, new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_,
    new_n2247_, new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_,
    new_n2253_, new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_,
    new_n2259_, new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_,
    new_n2265_, new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_,
    new_n2271_, new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_,
    new_n2277_, new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_,
    new_n2283_, new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_,
    new_n2289_, new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_,
    new_n2295_, new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_,
    new_n2301_, new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_,
    new_n2307_, new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_,
    new_n2313_, new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_,
    new_n2319_, new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_,
    new_n2325_, new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_,
    new_n2331_, new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_,
    new_n2337_, new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_,
    new_n2343_, new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_,
    new_n2349_, new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_,
    new_n2355_, new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_,
    new_n2361_, new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_,
    new_n2367_, new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_,
    new_n2373_, new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_,
    new_n2379_, new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_,
    new_n2385_, new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_,
    new_n2391_, new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_,
    new_n2397_, new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_,
    new_n2403_, new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_,
    new_n2409_, new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_,
    new_n2415_, new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_,
    new_n2421_, new_n2422_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_,
    new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_, new_n2512_,
    new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_, new_n2518_,
    new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_, new_n2524_,
    new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_, new_n2530_,
    new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_, new_n2536_,
    new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_, new_n2542_,
    new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_, new_n2548_,
    new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_, new_n2554_,
    new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_, new_n2560_,
    new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_, new_n2566_,
    new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_, new_n2572_,
    new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_, new_n2578_,
    new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_, new_n2585_,
    new_n2586_, new_n2587_, new_n2588_, new_n2589_, new_n2590_, new_n2591_,
    new_n2592_, new_n2593_, new_n2594_, new_n2595_, new_n2596_, new_n2597_,
    new_n2598_, new_n2599_, new_n2600_, new_n2601_, new_n2602_, new_n2603_,
    new_n2604_, new_n2605_, new_n2606_, new_n2607_, new_n2608_, new_n2609_,
    new_n2610_, new_n2611_, new_n2612_, new_n2613_, new_n2614_, new_n2615_,
    new_n2616_, new_n2617_, new_n2618_, new_n2619_, new_n2620_, new_n2621_,
    new_n2622_, new_n2623_, new_n2624_, new_n2625_, new_n2626_, new_n2627_,
    new_n2628_, new_n2629_, new_n2630_, new_n2631_, new_n2632_, new_n2633_,
    new_n2634_, new_n2635_, new_n2636_, new_n2637_, new_n2638_, new_n2639_,
    new_n2640_, new_n2641_, new_n2642_, new_n2643_, new_n2644_, new_n2645_,
    new_n2646_, new_n2647_, new_n2648_, new_n2650_, new_n2651_, new_n2652_,
    new_n2653_, new_n2654_, new_n2655_, new_n2656_, new_n2657_, new_n2658_,
    new_n2659_, new_n2660_, new_n2661_, new_n2662_, new_n2663_, new_n2664_,
    new_n2665_, new_n2666_, new_n2667_, new_n2668_, new_n2669_, new_n2670_,
    new_n2671_, new_n2672_, new_n2673_, new_n2674_, new_n2675_, new_n2676_,
    new_n2677_, new_n2678_, new_n2679_, new_n2680_, new_n2681_, new_n2682_,
    new_n2683_, new_n2684_, new_n2685_, new_n2686_, new_n2687_, new_n2688_,
    new_n2689_, new_n2690_, new_n2691_, new_n2692_, new_n2693_, new_n2694_,
    new_n2695_, new_n2696_, new_n2697_, new_n2698_, new_n2699_, new_n2700_,
    new_n2701_, new_n2702_, new_n2703_, new_n2704_, new_n2705_, new_n2706_,
    new_n2707_, new_n2708_, new_n2709_, new_n2710_, new_n2712_, new_n2713_,
    new_n2714_, new_n2715_, new_n2716_, new_n2717_, new_n2718_, new_n2719_,
    new_n2720_, new_n2721_, new_n2722_, new_n2723_, new_n2724_, new_n2725_,
    new_n2726_, new_n2727_, new_n2728_, new_n2729_, new_n2730_, new_n2731_,
    new_n2732_, new_n2733_, new_n2734_, new_n2735_, new_n2736_, new_n2737_,
    new_n2738_, new_n2739_, new_n2740_, new_n2741_, new_n2742_, new_n2743_,
    new_n2744_, new_n2745_, new_n2746_, new_n2747_, new_n2748_, new_n2749_,
    new_n2750_, new_n2751_, new_n2752_, new_n2753_, new_n2754_, new_n2755_,
    new_n2756_, new_n2757_, new_n2758_, new_n2759_, new_n2760_, new_n2761_,
    new_n2762_, new_n2763_, new_n2764_, new_n2765_, new_n2766_, new_n2767_,
    new_n2768_, new_n2769_, new_n2770_, new_n2771_, new_n2772_, new_n2773_,
    new_n2774_, new_n2775_, new_n2776_, new_n2778_, new_n2779_, new_n2780_,
    new_n2781_, new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_,
    new_n2787_, new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_,
    new_n2793_, new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_,
    new_n2799_, new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_,
    new_n2805_, new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_,
    new_n2811_, new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_,
    new_n2817_, new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_,
    new_n2823_, new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_,
    new_n2829_, new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_,
    new_n2835_, new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_,
    new_n2841_, new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_,
    new_n2847_, new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2908_,
    new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_, new_n2914_,
    new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_, new_n2920_,
    new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_, new_n2926_,
    new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_, new_n2932_,
    new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_, new_n2938_,
    new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_, new_n2944_,
    new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_, new_n2950_,
    new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_, new_n2956_,
    new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_, new_n2962_,
    new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_, new_n2968_,
    new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_, new_n2975_,
    new_n2976_, new_n2977_, new_n2978_, new_n2979_, new_n2980_, new_n2981_,
    new_n2982_, new_n2983_, new_n2984_, new_n2985_, new_n2986_, new_n2987_,
    new_n2988_, new_n2989_, new_n2990_, new_n2991_, new_n2992_, new_n2993_,
    new_n2994_, new_n2995_, new_n2996_, new_n2997_, new_n2998_, new_n2999_,
    new_n3000_, new_n3001_, new_n3002_, new_n3003_, new_n3004_, new_n3005_,
    new_n3006_, new_n3007_, new_n3008_, new_n3009_, new_n3010_, new_n3011_,
    new_n3012_, new_n3013_, new_n3014_, new_n3015_, new_n3016_, new_n3017_,
    new_n3018_, new_n3019_, new_n3020_, new_n3021_, new_n3022_, new_n3023_,
    new_n3024_, new_n3025_, new_n3026_, new_n3027_, new_n3028_, new_n3029_,
    new_n3031_, new_n3032_, new_n3033_, new_n3034_, new_n3035_, new_n3036_,
    new_n3037_, new_n3038_, new_n3039_, new_n3040_, new_n3041_, new_n3042_,
    new_n3043_, new_n3044_, new_n3045_, new_n3046_, new_n3047_, new_n3048_,
    new_n3049_, new_n3050_, new_n3051_, new_n3052_, new_n3053_, new_n3054_,
    new_n3055_, new_n3056_, new_n3057_, new_n3058_, new_n3059_, new_n3060_,
    new_n3061_, new_n3062_, new_n3063_, new_n3064_, new_n3065_, new_n3066_,
    new_n3067_, new_n3068_, new_n3069_, new_n3070_, new_n3071_, new_n3072_,
    new_n3073_, new_n3074_, new_n3075_, new_n3076_, new_n3077_, new_n3078_,
    new_n3079_, new_n3080_, new_n3081_, new_n3082_, new_n3083_, new_n3084_,
    new_n3085_, new_n3086_, new_n3088_, new_n3089_, new_n3090_, new_n3091_,
    new_n3092_, new_n3093_, new_n3094_, new_n3095_, new_n3096_, new_n3097_,
    new_n3098_, new_n3099_, new_n3100_, new_n3101_, new_n3102_, new_n3103_,
    new_n3104_, new_n3105_, new_n3106_, new_n3107_, new_n3108_, new_n3109_,
    new_n3110_, new_n3111_, new_n3112_, new_n3113_, new_n3114_, new_n3115_,
    new_n3116_, new_n3117_, new_n3118_, new_n3119_, new_n3120_, new_n3121_,
    new_n3122_, new_n3123_, new_n3124_, new_n3125_, new_n3126_, new_n3127_,
    new_n3128_, new_n3129_, new_n3131_, new_n3132_, new_n3133_, new_n3134_,
    new_n3135_, new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_,
    new_n3141_, new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_,
    new_n3147_, new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_,
    new_n3153_, new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_,
    new_n3159_, new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_,
    new_n3165_, new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_,
    new_n3171_, new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_,
    new_n3177_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3230_, new_n3231_, new_n3232_,
    new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_, new_n3238_,
    new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_, new_n3244_,
    new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_, new_n3250_,
    new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_, new_n3256_,
    new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_, new_n3262_,
    new_n3263_, new_n3265_, new_n3266_, new_n3267_, new_n3268_, new_n3269_,
    new_n3270_, new_n3271_, new_n3272_, new_n3273_, new_n3274_, new_n3275_,
    new_n3276_, new_n3277_, new_n3278_, new_n3279_, new_n3280_, new_n3281_,
    new_n3282_, new_n3283_, new_n3284_, new_n3285_, new_n3286_, new_n3287_,
    new_n3288_, new_n3289_, new_n3290_, new_n3291_, new_n3292_, new_n3293_,
    new_n3294_, new_n3295_, new_n3296_, new_n3297_, new_n3298_, new_n3299_,
    new_n3301_, new_n3302_, new_n3303_, new_n3304_, new_n3305_, new_n3306_,
    new_n3307_, new_n3308_, new_n3309_, new_n3310_, new_n3311_, new_n3312_,
    new_n3313_, new_n3314_, new_n3315_, new_n3316_, new_n3317_, new_n3318_,
    new_n3319_, new_n3320_, new_n3321_, new_n3322_, new_n3323_, new_n3324_,
    new_n3325_, new_n3326_, new_n3327_, new_n3328_, new_n3329_, new_n3330_,
    new_n3331_, new_n3332_, new_n3333_, new_n3334_, new_n3335_, new_n3336_,
    new_n3337_, new_n3338_, new_n3339_, new_n3340_, new_n3341_, new_n3342_,
    new_n3343_, new_n3344_, new_n3345_, new_n3346_, new_n3347_, new_n3349_,
    new_n3350_, new_n3351_, new_n3352_, new_n3353_, new_n3354_, new_n3355_,
    new_n3356_, new_n3357_, new_n3358_, new_n3359_, new_n3361_, new_n3362_,
    new_n3363_, new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_,
    new_n3369_, new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_,
    new_n3375_, new_n3376_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3388_,
    new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_, new_n3394_,
    new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_, new_n3400_,
    new_n3401_, new_n3402_, new_n3403_, new_n3405_, new_n3406_, new_n3407_,
    new_n3408_, new_n3409_, new_n3410_, new_n3412_, new_n3413_, new_n3414_,
    new_n3415_, new_n3416_, new_n3417_, new_n3418_, new_n3419_, new_n3421_,
    new_n3422_, new_n3423_, new_n3424_, new_n3425_, new_n3426_, new_n3428_,
    new_n3429_, new_n3430_, new_n3431_, new_n3432_;
  INVX1    g0000(.A(\a[22] ), .Y(new_n50_));
  OR4X1    g0001(.A(\a[3] ), .B(\a[2] ), .C(\a[1] ), .D(\a[0] ), .Y(new_n51_));
  OR4X1    g0002(.A(new_n51_), .B(\a[6] ), .C(\a[5] ), .D(\a[4] ), .Y(new_n52_));
  OR4X1    g0003(.A(new_n52_), .B(\a[9] ), .C(\a[8] ), .D(\a[7] ), .Y(new_n53_));
  OR4X1    g0004(.A(new_n53_), .B(\a[12] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n54_));
  OR4X1    g0005(.A(new_n54_), .B(\a[15] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n55_));
  OR4X1    g0006(.A(new_n55_), .B(\a[18] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n56_));
  AND2X1   g0007(.A(new_n56_), .B(new_n50_), .Y(new_n57_));
  XOR2X1   g0008(.A(new_n57_), .B(\a[19] ), .Y(new_n58_));
  INVX1    g0009(.A(\a[16] ), .Y(new_n59_));
  INVX1    g0010(.A(\a[17] ), .Y(new_n60_));
  NOR4X1   g0011(.A(new_n54_), .B(\a[15] ), .C(\a[14] ), .D(\a[13] ), .Y(new_n61_));
  NAND3X1  g0012(.A(new_n61_), .B(new_n60_), .C(new_n59_), .Y(new_n62_));
  NAND2X1  g0013(.A(new_n62_), .B(\a[18] ), .Y(new_n63_));
  AOI22X1  g0014(.A0(new_n63_), .A1(new_n57_), .B0(\a[22] ), .B1(\a[18] ), .Y(new_n64_));
  AOI21X1  g0015(.A0(new_n61_), .A1(new_n59_), .B0(\a[22] ), .Y(new_n65_));
  XOR2X1   g0016(.A(new_n65_), .B(new_n60_), .Y(new_n66_));
  AND2X1   g0017(.A(new_n55_), .B(new_n50_), .Y(new_n67_));
  XOR2X1   g0018(.A(new_n67_), .B(\a[16] ), .Y(new_n68_));
  AND2X1   g0019(.A(new_n68_), .B(new_n66_), .Y(new_n69_));
  NAND3X1  g0020(.A(new_n69_), .B(new_n64_), .C(new_n58_), .Y(new_n70_));
  INVX1    g0021(.A(\a[21] ), .Y(new_n71_));
  INVX1    g0022(.A(\a[19] ), .Y(new_n72_));
  INVX1    g0023(.A(\a[20] ), .Y(new_n73_));
  NOR4X1   g0024(.A(new_n55_), .B(\a[18] ), .C(\a[17] ), .D(\a[16] ), .Y(new_n74_));
  NAND3X1  g0025(.A(new_n74_), .B(new_n73_), .C(new_n72_), .Y(new_n75_));
  AND2X1   g0026(.A(new_n75_), .B(\a[21] ), .Y(new_n76_));
  OAI21X1  g0027(.A0(new_n75_), .A1(\a[21] ), .B0(new_n50_), .Y(new_n77_));
  OAI22X1  g0028(.A0(new_n77_), .A1(new_n76_), .B0(new_n50_), .B1(new_n71_), .Y(new_n78_));
  AND2X1   g0029(.A(\a[22] ), .B(\a[20] ), .Y(new_n79_));
  NOR3X1   g0030(.A(new_n56_), .B(\a[20] ), .C(\a[19] ), .Y(new_n80_));
  AOI21X1  g0031(.A0(new_n74_), .A1(new_n72_), .B0(new_n73_), .Y(new_n81_));
  NOR3X1   g0032(.A(new_n81_), .B(new_n80_), .C(\a[22] ), .Y(new_n82_));
  OR2X1    g0033(.A(new_n82_), .B(new_n79_), .Y(new_n83_));
  AND2X1   g0034(.A(\a[22] ), .B(\a[15] ), .Y(new_n84_));
  INVX1    g0035(.A(\a[13] ), .Y(new_n85_));
  INVX1    g0036(.A(\a[14] ), .Y(new_n86_));
  NOR4X1   g0037(.A(new_n53_), .B(\a[12] ), .C(\a[11] ), .D(\a[10] ), .Y(new_n87_));
  NAND3X1  g0038(.A(new_n87_), .B(new_n86_), .C(new_n85_), .Y(new_n88_));
  NAND2X1  g0039(.A(new_n88_), .B(\a[15] ), .Y(new_n89_));
  AOI21X1  g0040(.A0(new_n89_), .A1(new_n67_), .B0(new_n84_), .Y(new_n90_));
  NOR4X1   g0041(.A(new_n90_), .B(new_n83_), .C(new_n78_), .D(new_n70_), .Y(new_n91_));
  NOR2X1   g0042(.A(new_n82_), .B(new_n79_), .Y(new_n92_));
  XOR2X1   g0043(.A(new_n65_), .B(\a[17] ), .Y(new_n93_));
  XOR2X1   g0044(.A(new_n67_), .B(new_n59_), .Y(new_n94_));
  AND2X1   g0045(.A(new_n94_), .B(new_n93_), .Y(new_n95_));
  NAND3X1  g0046(.A(new_n95_), .B(new_n64_), .C(new_n58_), .Y(new_n96_));
  NOR4X1   g0047(.A(new_n96_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n97_));
  NOR2X1   g0048(.A(new_n97_), .B(new_n91_), .Y(new_n98_));
  OR2X1    g0049(.A(new_n80_), .B(new_n71_), .Y(new_n99_));
  AOI21X1  g0050(.A0(new_n80_), .A1(new_n71_), .B0(\a[22] ), .Y(new_n100_));
  AOI22X1  g0051(.A0(new_n100_), .A1(new_n99_), .B0(\a[22] ), .B1(\a[21] ), .Y(new_n101_));
  OR2X1    g0052(.A(new_n74_), .B(\a[22] ), .Y(new_n102_));
  NAND2X1  g0053(.A(\a[22] ), .B(\a[18] ), .Y(new_n103_));
  AND2X1   g0054(.A(new_n62_), .B(\a[18] ), .Y(new_n104_));
  OAI21X1  g0055(.A0(new_n104_), .A1(new_n102_), .B0(new_n103_), .Y(new_n105_));
  NAND3X1  g0056(.A(new_n69_), .B(new_n105_), .C(new_n58_), .Y(new_n106_));
  NOR4X1   g0057(.A(new_n106_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n107_));
  INVX1    g0058(.A(new_n90_), .Y(new_n108_));
  NAND3X1  g0059(.A(new_n95_), .B(new_n105_), .C(new_n58_), .Y(new_n109_));
  NOR4X1   g0060(.A(new_n109_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n110_));
  AND2X1   g0061(.A(new_n68_), .B(new_n93_), .Y(new_n111_));
  NAND3X1  g0062(.A(new_n111_), .B(new_n64_), .C(new_n58_), .Y(new_n112_));
  NOR4X1   g0063(.A(new_n112_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n113_));
  AND2X1   g0064(.A(new_n94_), .B(new_n66_), .Y(new_n114_));
  NAND3X1  g0065(.A(new_n114_), .B(new_n64_), .C(new_n58_), .Y(new_n115_));
  NOR4X1   g0066(.A(new_n115_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n116_));
  NOR4X1   g0067(.A(new_n116_), .B(new_n113_), .C(new_n110_), .D(new_n107_), .Y(new_n117_));
  AND2X1   g0068(.A(new_n117_), .B(new_n98_), .Y(new_n118_));
  XOR2X1   g0069(.A(new_n57_), .B(new_n72_), .Y(new_n119_));
  NAND3X1  g0070(.A(new_n111_), .B(new_n64_), .C(new_n119_), .Y(new_n120_));
  NOR4X1   g0071(.A(new_n120_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n121_));
  NAND3X1  g0072(.A(new_n95_), .B(new_n105_), .C(new_n119_), .Y(new_n122_));
  NOR4X1   g0073(.A(new_n122_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n123_));
  NAND3X1  g0074(.A(new_n69_), .B(new_n105_), .C(new_n119_), .Y(new_n124_));
  NOR4X1   g0075(.A(new_n124_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n125_));
  NAND3X1  g0076(.A(new_n69_), .B(new_n64_), .C(new_n119_), .Y(new_n126_));
  NOR4X1   g0077(.A(new_n126_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n127_));
  OR4X1    g0078(.A(new_n127_), .B(new_n125_), .C(new_n123_), .D(new_n121_), .Y(new_n128_));
  NAND3X1  g0079(.A(new_n114_), .B(new_n105_), .C(new_n119_), .Y(new_n129_));
  NOR4X1   g0080(.A(new_n129_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n130_));
  NOR4X1   g0081(.A(new_n96_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n131_));
  NOR4X1   g0082(.A(new_n124_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n132_));
  NAND3X1  g0083(.A(new_n114_), .B(new_n105_), .C(new_n58_), .Y(new_n133_));
  NOR4X1   g0084(.A(new_n133_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n134_));
  OR4X1    g0085(.A(new_n134_), .B(new_n132_), .C(new_n131_), .D(new_n130_), .Y(new_n135_));
  NOR4X1   g0086(.A(new_n120_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n136_));
  NOR4X1   g0087(.A(new_n109_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n137_));
  OR2X1    g0088(.A(new_n137_), .B(new_n136_), .Y(new_n138_));
  NOR4X1   g0089(.A(new_n120_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n139_));
  NAND3X1  g0090(.A(new_n95_), .B(new_n64_), .C(new_n119_), .Y(new_n140_));
  NOR4X1   g0091(.A(new_n140_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n141_));
  OR2X1    g0092(.A(new_n141_), .B(new_n139_), .Y(new_n142_));
  NOR4X1   g0093(.A(new_n142_), .B(new_n138_), .C(new_n135_), .D(new_n128_), .Y(new_n143_));
  NAND2X1  g0094(.A(new_n143_), .B(new_n118_), .Y(new_n144_));
  NOR4X1   g0095(.A(new_n124_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n145_));
  NAND3X1  g0096(.A(new_n111_), .B(new_n105_), .C(new_n58_), .Y(new_n146_));
  NOR4X1   g0097(.A(new_n146_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n147_));
  NAND3X1  g0098(.A(new_n114_), .B(new_n64_), .C(new_n119_), .Y(new_n148_));
  NOR4X1   g0099(.A(new_n148_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n149_));
  NOR4X1   g0100(.A(new_n148_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n150_));
  OR4X1    g0101(.A(new_n150_), .B(new_n149_), .C(new_n147_), .D(new_n145_), .Y(new_n151_));
  NOR2X1   g0102(.A(new_n151_), .B(new_n144_), .Y(new_n152_));
  INVX1    g0103(.A(new_n152_), .Y(new_n153_));
  OR4X1    g0104(.A(new_n112_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n154_));
  NOR4X1   g0105(.A(new_n129_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n155_));
  INVX1    g0106(.A(new_n155_), .Y(new_n156_));
  NOR4X1   g0107(.A(new_n146_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n157_));
  NOR4X1   g0108(.A(new_n96_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n158_));
  NOR4X1   g0109(.A(new_n126_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n159_));
  NOR3X1   g0110(.A(new_n159_), .B(new_n158_), .C(new_n157_), .Y(new_n160_));
  NAND3X1  g0111(.A(new_n160_), .B(new_n156_), .C(new_n154_), .Y(new_n161_));
  NOR4X1   g0112(.A(new_n148_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n162_));
  NOR4X1   g0113(.A(new_n112_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n163_));
  NOR4X1   g0114(.A(new_n133_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n164_));
  NOR4X1   g0115(.A(new_n106_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n165_));
  OR4X1    g0116(.A(new_n165_), .B(new_n164_), .C(new_n163_), .D(new_n162_), .Y(new_n166_));
  NOR4X1   g0117(.A(new_n129_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n167_));
  NOR4X1   g0118(.A(new_n133_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n168_));
  NOR4X1   g0119(.A(new_n112_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n169_));
  NOR4X1   g0120(.A(new_n90_), .B(new_n92_), .C(new_n78_), .D(new_n70_), .Y(new_n170_));
  OR4X1    g0121(.A(new_n170_), .B(new_n169_), .C(new_n168_), .D(new_n167_), .Y(new_n171_));
  NOR4X1   g0122(.A(new_n133_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n172_));
  NOR4X1   g0123(.A(new_n120_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n173_));
  NOR4X1   g0124(.A(new_n106_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n174_));
  NOR4X1   g0125(.A(new_n112_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n175_));
  OR4X1    g0126(.A(new_n175_), .B(new_n174_), .C(new_n173_), .D(new_n172_), .Y(new_n176_));
  OR4X1    g0127(.A(new_n176_), .B(new_n171_), .C(new_n166_), .D(new_n161_), .Y(new_n177_));
  NAND3X1  g0128(.A(new_n111_), .B(new_n105_), .C(new_n119_), .Y(new_n178_));
  NOR4X1   g0129(.A(new_n178_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n179_));
  NOR4X1   g0130(.A(new_n109_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n180_));
  OR2X1    g0131(.A(new_n180_), .B(new_n179_), .Y(new_n181_));
  NOR4X1   g0132(.A(new_n109_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n182_));
  NOR4X1   g0133(.A(new_n124_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n183_));
  NOR4X1   g0134(.A(new_n96_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n184_));
  NOR4X1   g0135(.A(new_n112_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n185_));
  OR2X1    g0136(.A(new_n185_), .B(new_n184_), .Y(new_n186_));
  OR4X1    g0137(.A(new_n186_), .B(new_n183_), .C(new_n182_), .D(new_n181_), .Y(new_n187_));
  NOR4X1   g0138(.A(new_n178_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n188_));
  NOR4X1   g0139(.A(new_n90_), .B(new_n92_), .C(new_n101_), .D(new_n70_), .Y(new_n189_));
  NOR4X1   g0140(.A(new_n178_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n190_));
  OR2X1    g0141(.A(new_n190_), .B(new_n189_), .Y(new_n191_));
  NOR4X1   g0142(.A(new_n109_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n192_));
  NOR4X1   g0143(.A(new_n106_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n193_));
  OR2X1    g0144(.A(new_n193_), .B(new_n192_), .Y(new_n194_));
  NOR4X1   g0145(.A(new_n108_), .B(new_n92_), .C(new_n101_), .D(new_n70_), .Y(new_n195_));
  NOR4X1   g0146(.A(new_n122_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n196_));
  NOR4X1   g0147(.A(new_n122_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n197_));
  NOR4X1   g0148(.A(new_n109_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n198_));
  OR4X1    g0149(.A(new_n198_), .B(new_n197_), .C(new_n196_), .D(new_n195_), .Y(new_n199_));
  OR4X1    g0150(.A(new_n199_), .B(new_n194_), .C(new_n191_), .D(new_n188_), .Y(new_n200_));
  OR2X1    g0151(.A(new_n200_), .B(new_n187_), .Y(new_n201_));
  NOR4X1   g0152(.A(new_n109_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n202_));
  NOR4X1   g0153(.A(new_n133_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n203_));
  NOR4X1   g0154(.A(new_n115_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n204_));
  NOR4X1   g0155(.A(new_n129_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n205_));
  OR4X1    g0156(.A(new_n205_), .B(new_n204_), .C(new_n203_), .D(new_n202_), .Y(new_n206_));
  NOR4X1   g0157(.A(new_n126_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n207_));
  NOR4X1   g0158(.A(new_n146_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n208_));
  OR2X1    g0159(.A(new_n208_), .B(new_n207_), .Y(new_n209_));
  NOR4X1   g0160(.A(new_n115_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n210_));
  NOR4X1   g0161(.A(new_n126_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n211_));
  OR2X1    g0162(.A(new_n211_), .B(new_n210_), .Y(new_n212_));
  NOR4X1   g0163(.A(new_n124_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n213_));
  NOR4X1   g0164(.A(new_n140_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n214_));
  OR4X1    g0165(.A(new_n122_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n215_));
  INVX1    g0166(.A(new_n215_), .Y(new_n216_));
  NOR3X1   g0167(.A(new_n216_), .B(new_n214_), .C(new_n213_), .Y(new_n217_));
  INVX1    g0168(.A(new_n217_), .Y(new_n218_));
  NOR4X1   g0169(.A(new_n109_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n219_));
  NOR4X1   g0170(.A(new_n90_), .B(new_n83_), .C(new_n101_), .D(new_n70_), .Y(new_n220_));
  NOR4X1   g0171(.A(new_n96_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n221_));
  OR4X1    g0172(.A(new_n221_), .B(new_n220_), .C(new_n219_), .D(new_n218_), .Y(new_n222_));
  OR4X1    g0173(.A(new_n222_), .B(new_n212_), .C(new_n209_), .D(new_n206_), .Y(new_n223_));
  NOR4X1   g0174(.A(new_n223_), .B(new_n201_), .C(new_n177_), .D(new_n153_), .Y(new_n224_));
  INVX1    g0175(.A(new_n224_), .Y(new_n225_));
  INVX1    g0176(.A(\a[5] ), .Y(new_n226_));
  NOR2X1   g0177(.A(new_n51_), .B(\a[4] ), .Y(new_n227_));
  NOR2X1   g0178(.A(new_n227_), .B(\a[22] ), .Y(new_n228_));
  XOR2X1   g0179(.A(new_n228_), .B(new_n226_), .Y(new_n229_));
  INVX1    g0180(.A(new_n229_), .Y(new_n230_));
  AND2X1   g0181(.A(new_n51_), .B(\a[4] ), .Y(new_n231_));
  NOR3X1   g0182(.A(new_n231_), .B(new_n227_), .C(\a[22] ), .Y(new_n232_));
  AOI21X1  g0183(.A0(\a[22] ), .A1(\a[4] ), .B0(new_n232_), .Y(new_n233_));
  XOR2X1   g0184(.A(new_n233_), .B(new_n230_), .Y(new_n234_));
  NOR3X1   g0185(.A(\a[2] ), .B(\a[1] ), .C(\a[0] ), .Y(new_n235_));
  NOR2X1   g0186(.A(new_n235_), .B(\a[22] ), .Y(new_n236_));
  INVX1    g0187(.A(new_n236_), .Y(new_n237_));
  XOR2X1   g0188(.A(new_n237_), .B(\a[3] ), .Y(new_n238_));
  INVX1    g0189(.A(\a[2] ), .Y(new_n239_));
  INVX1    g0190(.A(\a[0] ), .Y(new_n240_));
  INVX1    g0191(.A(\a[1] ), .Y(new_n241_));
  AOI21X1  g0192(.A0(new_n241_), .A1(new_n240_), .B0(new_n239_), .Y(new_n242_));
  OAI22X1  g0193(.A0(new_n242_), .A1(new_n237_), .B0(new_n50_), .B1(new_n239_), .Y(new_n243_));
  XOR2X1   g0194(.A(new_n243_), .B(new_n238_), .Y(new_n244_));
  NOR2X1   g0195(.A(new_n244_), .B(new_n234_), .Y(new_n245_));
  OR2X1    g0196(.A(new_n183_), .B(new_n182_), .Y(new_n246_));
  NOR4X1   g0197(.A(new_n120_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n247_));
  NOR4X1   g0198(.A(new_n106_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n248_));
  NOR4X1   g0199(.A(new_n108_), .B(new_n92_), .C(new_n78_), .D(new_n70_), .Y(new_n249_));
  NOR4X1   g0200(.A(new_n249_), .B(new_n248_), .C(new_n247_), .D(new_n164_), .Y(new_n250_));
  NOR4X1   g0201(.A(new_n126_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n251_));
  NOR4X1   g0202(.A(new_n122_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n252_));
  NOR4X1   g0203(.A(new_n126_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n253_));
  NOR3X1   g0204(.A(new_n253_), .B(new_n252_), .C(new_n251_), .Y(new_n254_));
  NOR4X1   g0205(.A(new_n140_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n255_));
  NOR4X1   g0206(.A(new_n148_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n256_));
  NOR3X1   g0207(.A(new_n256_), .B(new_n255_), .C(new_n110_), .Y(new_n257_));
  NAND3X1  g0208(.A(new_n257_), .B(new_n254_), .C(new_n250_), .Y(new_n258_));
  NOR4X1   g0209(.A(new_n129_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n259_));
  OR2X1    g0210(.A(new_n259_), .B(new_n127_), .Y(new_n260_));
  NOR4X1   g0211(.A(new_n106_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n261_));
  NOR4X1   g0212(.A(new_n146_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n262_));
  OR4X1    g0213(.A(new_n262_), .B(new_n261_), .C(new_n260_), .D(new_n116_), .Y(new_n263_));
  NOR4X1   g0214(.A(new_n178_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n264_));
  NOR4X1   g0215(.A(new_n96_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n265_));
  OR4X1    g0216(.A(new_n265_), .B(new_n264_), .C(new_n157_), .D(new_n147_), .Y(new_n266_));
  OR4X1    g0217(.A(new_n266_), .B(new_n263_), .C(new_n258_), .D(new_n246_), .Y(new_n267_));
  OR2X1    g0218(.A(new_n169_), .B(new_n139_), .Y(new_n268_));
  NOR4X1   g0219(.A(new_n148_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n269_));
  OR2X1    g0220(.A(new_n269_), .B(new_n137_), .Y(new_n270_));
  NOR4X1   g0221(.A(new_n146_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n271_));
  NOR4X1   g0222(.A(new_n148_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n272_));
  OR2X1    g0223(.A(new_n272_), .B(new_n271_), .Y(new_n273_));
  OR4X1    g0224(.A(new_n273_), .B(new_n270_), .C(new_n268_), .D(new_n194_), .Y(new_n274_));
  OR4X1    g0225(.A(new_n109_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n275_));
  OR4X1    g0226(.A(new_n140_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n276_));
  NAND3X1  g0227(.A(new_n276_), .B(new_n275_), .C(new_n215_), .Y(new_n277_));
  OR4X1    g0228(.A(new_n126_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n278_));
  INVX1    g0229(.A(new_n278_), .Y(new_n279_));
  NOR4X1   g0230(.A(new_n133_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n280_));
  NOR4X1   g0231(.A(new_n140_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n281_));
  OR4X1    g0232(.A(new_n281_), .B(new_n280_), .C(new_n279_), .D(new_n277_), .Y(new_n282_));
  NOR4X1   g0233(.A(new_n126_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n283_));
  OR4X1    g0234(.A(new_n283_), .B(new_n220_), .C(new_n175_), .D(new_n131_), .Y(new_n284_));
  OR4X1    g0235(.A(new_n106_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n285_));
  INVX1    g0236(.A(new_n203_), .Y(new_n286_));
  NOR4X1   g0237(.A(new_n133_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n287_));
  INVX1    g0238(.A(new_n287_), .Y(new_n288_));
  NAND3X1  g0239(.A(new_n288_), .B(new_n286_), .C(new_n285_), .Y(new_n289_));
  OR4X1    g0240(.A(new_n289_), .B(new_n284_), .C(new_n282_), .D(new_n274_), .Y(new_n290_));
  OR2X1    g0241(.A(new_n196_), .B(new_n195_), .Y(new_n291_));
  NOR4X1   g0242(.A(new_n115_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n292_));
  NOR4X1   g0243(.A(new_n122_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n293_));
  NOR4X1   g0244(.A(new_n122_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n294_));
  OR4X1    g0245(.A(new_n294_), .B(new_n293_), .C(new_n292_), .D(new_n123_), .Y(new_n295_));
  OR2X1    g0246(.A(new_n202_), .B(new_n130_), .Y(new_n296_));
  OR2X1    g0247(.A(new_n189_), .B(new_n162_), .Y(new_n297_));
  OR4X1    g0248(.A(new_n297_), .B(new_n296_), .C(new_n295_), .D(new_n291_), .Y(new_n298_));
  OR4X1    g0249(.A(new_n90_), .B(new_n92_), .C(new_n78_), .D(new_n70_), .Y(new_n299_));
  OR4X1    g0250(.A(new_n112_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n300_));
  OR4X1    g0251(.A(new_n120_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n301_));
  NAND3X1  g0252(.A(new_n301_), .B(new_n300_), .C(new_n299_), .Y(new_n302_));
  NOR4X1   g0253(.A(new_n96_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n303_));
  NOR4X1   g0254(.A(new_n178_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n304_));
  NOR4X1   g0255(.A(new_n129_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n305_));
  OR4X1    g0256(.A(new_n305_), .B(new_n304_), .C(new_n303_), .D(new_n136_), .Y(new_n306_));
  OR4X1    g0257(.A(new_n306_), .B(new_n302_), .C(new_n180_), .D(new_n134_), .Y(new_n307_));
  NOR4X1   g0258(.A(new_n307_), .B(new_n298_), .C(new_n290_), .D(new_n267_), .Y(new_n308_));
  INVX1    g0259(.A(\a[11] ), .Y(new_n309_));
  NOR2X1   g0260(.A(new_n53_), .B(\a[10] ), .Y(new_n310_));
  NOR2X1   g0261(.A(new_n310_), .B(\a[22] ), .Y(new_n311_));
  XOR2X1   g0262(.A(new_n311_), .B(new_n309_), .Y(new_n312_));
  INVX1    g0263(.A(new_n312_), .Y(new_n313_));
  NOR4X1   g0264(.A(new_n133_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n314_));
  NOR4X1   g0265(.A(new_n106_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n315_));
  OR2X1    g0266(.A(new_n315_), .B(new_n314_), .Y(new_n316_));
  NOR4X1   g0267(.A(new_n124_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n317_));
  OR4X1    g0268(.A(new_n317_), .B(new_n269_), .C(new_n167_), .D(new_n137_), .Y(new_n318_));
  OR2X1    g0269(.A(new_n155_), .B(new_n132_), .Y(new_n319_));
  OR2X1    g0270(.A(new_n319_), .B(new_n162_), .Y(new_n320_));
  NOR4X1   g0271(.A(new_n146_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n321_));
  NOR4X1   g0272(.A(new_n146_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n322_));
  OR4X1    g0273(.A(new_n322_), .B(new_n321_), .C(new_n248_), .D(new_n202_), .Y(new_n323_));
  OR4X1    g0274(.A(new_n323_), .B(new_n320_), .C(new_n318_), .D(new_n316_), .Y(new_n324_));
  NOR4X1   g0275(.A(new_n112_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n325_));
  OR4X1    g0276(.A(new_n325_), .B(new_n287_), .C(new_n265_), .D(new_n169_), .Y(new_n326_));
  OR2X1    g0277(.A(new_n203_), .B(new_n149_), .Y(new_n327_));
  OR2X1    g0278(.A(new_n327_), .B(new_n256_), .Y(new_n328_));
  NOR4X1   g0279(.A(new_n120_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n329_));
  NOR4X1   g0280(.A(new_n140_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n330_));
  OR2X1    g0281(.A(new_n330_), .B(new_n329_), .Y(new_n331_));
  NOR4X1   g0282(.A(new_n146_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n332_));
  NAND3X1  g0283(.A(new_n108_), .B(new_n92_), .C(new_n78_), .Y(new_n333_));
  AOI21X1  g0284(.A0(new_n140_), .A1(new_n126_), .B0(new_n333_), .Y(new_n334_));
  OR4X1    g0285(.A(new_n334_), .B(new_n332_), .C(new_n331_), .D(new_n252_), .Y(new_n335_));
  NOR4X1   g0286(.A(new_n112_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n336_));
  NOR4X1   g0287(.A(new_n112_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n337_));
  OR4X1    g0288(.A(new_n106_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n338_));
  OR4X1    g0289(.A(new_n133_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n339_));
  OR4X1    g0290(.A(new_n106_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n340_));
  NAND3X1  g0291(.A(new_n340_), .B(new_n339_), .C(new_n338_), .Y(new_n341_));
  OR4X1    g0292(.A(new_n341_), .B(new_n337_), .C(new_n182_), .D(new_n336_), .Y(new_n342_));
  OR2X1    g0293(.A(new_n192_), .B(new_n147_), .Y(new_n343_));
  OR4X1    g0294(.A(new_n343_), .B(new_n247_), .C(new_n207_), .D(new_n97_), .Y(new_n344_));
  OR4X1    g0295(.A(new_n344_), .B(new_n342_), .C(new_n335_), .D(new_n328_), .Y(new_n345_));
  NOR4X1   g0296(.A(new_n96_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n346_));
  NOR4X1   g0297(.A(new_n108_), .B(new_n83_), .C(new_n78_), .D(new_n70_), .Y(new_n347_));
  NOR4X1   g0298(.A(new_n115_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n348_));
  OR4X1    g0299(.A(new_n348_), .B(new_n347_), .C(new_n346_), .D(new_n91_), .Y(new_n349_));
  NOR4X1   g0300(.A(new_n349_), .B(new_n345_), .C(new_n326_), .D(new_n324_), .Y(new_n350_));
  NOR2X1   g0301(.A(new_n317_), .B(new_n167_), .Y(new_n351_));
  INVX1    g0302(.A(new_n351_), .Y(new_n352_));
  INVX1    g0303(.A(new_n293_), .Y(new_n353_));
  INVX1    g0304(.A(new_n304_), .Y(new_n354_));
  OR4X1    g0305(.A(new_n124_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n355_));
  NAND3X1  g0306(.A(new_n355_), .B(new_n354_), .C(new_n353_), .Y(new_n356_));
  NOR4X1   g0307(.A(new_n122_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n357_));
  NOR4X1   g0308(.A(new_n178_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n358_));
  OR4X1    g0309(.A(new_n358_), .B(new_n204_), .C(new_n170_), .D(new_n131_), .Y(new_n359_));
  OR4X1    g0310(.A(new_n359_), .B(new_n357_), .C(new_n292_), .D(new_n249_), .Y(new_n360_));
  OR4X1    g0311(.A(new_n360_), .B(new_n356_), .C(new_n319_), .D(new_n352_), .Y(new_n361_));
  OR2X1    g0312(.A(new_n251_), .B(new_n205_), .Y(new_n362_));
  NOR4X1   g0313(.A(new_n120_), .B(new_n108_), .C(new_n92_), .D(new_n78_), .Y(new_n363_));
  OR4X1    g0314(.A(new_n363_), .B(new_n362_), .C(new_n281_), .D(new_n253_), .Y(new_n364_));
  OR4X1    g0315(.A(new_n364_), .B(new_n305_), .C(new_n214_), .D(new_n136_), .Y(new_n365_));
  NOR4X1   g0316(.A(new_n365_), .B(new_n361_), .C(new_n345_), .D(new_n183_), .Y(new_n366_));
  XOR2X1   g0317(.A(new_n366_), .B(new_n350_), .Y(new_n367_));
  INVX1    g0318(.A(new_n367_), .Y(new_n368_));
  OR4X1    g0319(.A(new_n185_), .B(new_n184_), .C(new_n173_), .D(new_n172_), .Y(new_n369_));
  OR4X1    g0320(.A(new_n369_), .B(new_n221_), .C(new_n121_), .D(new_n107_), .Y(new_n370_));
  NOR3X1   g0321(.A(new_n370_), .B(new_n261_), .C(new_n134_), .Y(new_n371_));
  NOR4X1   g0322(.A(new_n108_), .B(new_n83_), .C(new_n101_), .D(new_n70_), .Y(new_n372_));
  NOR4X1   g0323(.A(new_n372_), .B(new_n259_), .C(new_n188_), .D(new_n123_), .Y(new_n373_));
  INVX1    g0324(.A(new_n373_), .Y(new_n374_));
  OR4X1    g0325(.A(new_n178_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n375_));
  OR4X1    g0326(.A(new_n115_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n376_));
  OR4X1    g0327(.A(new_n115_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n377_));
  NAND3X1  g0328(.A(new_n377_), .B(new_n376_), .C(new_n375_), .Y(new_n378_));
  NOR4X1   g0329(.A(new_n129_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n379_));
  NOR4X1   g0330(.A(new_n379_), .B(new_n378_), .C(new_n374_), .D(new_n220_), .Y(new_n380_));
  OR4X1    g0331(.A(new_n193_), .B(new_n165_), .C(new_n150_), .D(new_n127_), .Y(new_n381_));
  OR2X1    g0332(.A(new_n272_), .B(new_n208_), .Y(new_n382_));
  NOR4X1   g0333(.A(new_n382_), .B(new_n381_), .C(new_n219_), .D(new_n189_), .Y(new_n383_));
  NAND3X1  g0334(.A(new_n383_), .B(new_n380_), .C(new_n371_), .Y(new_n384_));
  NOR4X1   g0335(.A(new_n115_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n385_));
  OR4X1    g0336(.A(new_n385_), .B(new_n303_), .C(new_n163_), .D(new_n158_), .Y(new_n386_));
  OR2X1    g0337(.A(new_n213_), .B(new_n175_), .Y(new_n387_));
  NOR4X1   g0338(.A(new_n178_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n388_));
  OR2X1    g0339(.A(new_n388_), .B(new_n125_), .Y(new_n389_));
  OR4X1    g0340(.A(new_n389_), .B(new_n387_), .C(new_n291_), .D(new_n116_), .Y(new_n390_));
  OR4X1    g0341(.A(new_n390_), .B(new_n386_), .C(new_n264_), .D(new_n216_), .Y(new_n391_));
  INVX1    g0342(.A(new_n164_), .Y(new_n392_));
  OR4X1    g0343(.A(new_n109_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n393_));
  NOR4X1   g0344(.A(new_n271_), .B(new_n168_), .C(new_n113_), .D(new_n110_), .Y(new_n394_));
  NAND3X1  g0345(.A(new_n394_), .B(new_n393_), .C(new_n392_), .Y(new_n395_));
  OR2X1    g0346(.A(new_n180_), .B(new_n159_), .Y(new_n396_));
  NOR4X1   g0347(.A(new_n140_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n397_));
  NOR4X1   g0348(.A(new_n140_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n398_));
  OR4X1    g0349(.A(new_n398_), .B(new_n397_), .C(new_n262_), .D(new_n157_), .Y(new_n399_));
  OR4X1    g0350(.A(new_n399_), .B(new_n396_), .C(new_n395_), .D(new_n391_), .Y(new_n400_));
  NOR2X1   g0351(.A(new_n400_), .B(new_n384_), .Y(new_n401_));
  INVX1    g0352(.A(new_n401_), .Y(new_n402_));
  AOI21X1  g0353(.A0(new_n366_), .A1(new_n350_), .B0(new_n402_), .Y(new_n403_));
  NOR2X1   g0354(.A(new_n403_), .B(new_n368_), .Y(new_n404_));
  NOR2X1   g0355(.A(new_n366_), .B(new_n350_), .Y(new_n405_));
  NOR2X1   g0356(.A(new_n405_), .B(new_n401_), .Y(new_n406_));
  NOR2X1   g0357(.A(new_n406_), .B(new_n368_), .Y(new_n407_));
  MX2X1    g0358(.A(new_n407_), .B(new_n404_), .S0(new_n313_), .Y(new_n408_));
  AND2X1   g0359(.A(\a[22] ), .B(\a[10] ), .Y(new_n409_));
  AND2X1   g0360(.A(new_n53_), .B(\a[10] ), .Y(new_n410_));
  NOR3X1   g0361(.A(new_n410_), .B(new_n310_), .C(\a[22] ), .Y(new_n411_));
  NOR2X1   g0362(.A(new_n411_), .B(new_n409_), .Y(new_n412_));
  INVX1    g0363(.A(new_n412_), .Y(new_n413_));
  NOR3X1   g0364(.A(new_n413_), .B(new_n406_), .C(new_n367_), .Y(new_n414_));
  NOR3X1   g0365(.A(new_n412_), .B(new_n403_), .C(new_n367_), .Y(new_n415_));
  OR2X1    g0366(.A(new_n188_), .B(new_n116_), .Y(new_n416_));
  OR4X1    g0367(.A(new_n303_), .B(new_n252_), .C(new_n183_), .D(new_n134_), .Y(new_n417_));
  NOR2X1   g0368(.A(new_n417_), .B(new_n416_), .Y(new_n418_));
  OR2X1    g0369(.A(new_n248_), .B(new_n147_), .Y(new_n419_));
  OR2X1    g0370(.A(new_n292_), .B(new_n197_), .Y(new_n420_));
  NOR4X1   g0371(.A(new_n420_), .B(new_n419_), .C(new_n192_), .D(new_n173_), .Y(new_n421_));
  OR4X1    g0372(.A(new_n129_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n422_));
  OR4X1    g0373(.A(new_n124_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n423_));
  OR4X1    g0374(.A(new_n129_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n424_));
  NAND3X1  g0375(.A(new_n424_), .B(new_n423_), .C(new_n422_), .Y(new_n425_));
  NOR4X1   g0376(.A(new_n178_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n426_));
  NOR4X1   g0377(.A(new_n426_), .B(new_n425_), .C(new_n347_), .D(new_n210_), .Y(new_n427_));
  NAND3X1  g0378(.A(new_n427_), .B(new_n421_), .C(new_n418_), .Y(new_n428_));
  OR2X1    g0379(.A(new_n385_), .B(new_n137_), .Y(new_n429_));
  NOR4X1   g0380(.A(new_n115_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n430_));
  OR4X1    g0381(.A(new_n430_), .B(new_n293_), .C(new_n253_), .D(new_n249_), .Y(new_n431_));
  OR2X1    g0382(.A(new_n431_), .B(new_n429_), .Y(new_n432_));
  OR2X1    g0383(.A(new_n202_), .B(new_n195_), .Y(new_n433_));
  OR4X1    g0384(.A(new_n358_), .B(new_n280_), .C(new_n214_), .D(new_n141_), .Y(new_n434_));
  OR2X1    g0385(.A(new_n434_), .B(new_n433_), .Y(new_n435_));
  OR4X1    g0386(.A(new_n435_), .B(new_n432_), .C(new_n320_), .D(new_n284_), .Y(new_n436_));
  NOR4X1   g0387(.A(new_n140_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n437_));
  OR2X1    g0388(.A(new_n207_), .B(new_n107_), .Y(new_n438_));
  OR4X1    g0389(.A(new_n148_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n439_));
  OR4X1    g0390(.A(new_n122_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n440_));
  OR4X1    g0391(.A(new_n129_), .B(new_n90_), .C(new_n92_), .D(new_n101_), .Y(new_n441_));
  NAND3X1  g0392(.A(new_n441_), .B(new_n440_), .C(new_n439_), .Y(new_n442_));
  OR4X1    g0393(.A(new_n259_), .B(new_n198_), .C(new_n139_), .D(new_n110_), .Y(new_n443_));
  OR4X1    g0394(.A(new_n443_), .B(new_n442_), .C(new_n438_), .D(new_n437_), .Y(new_n444_));
  OR4X1    g0395(.A(new_n346_), .B(new_n305_), .C(new_n287_), .D(new_n272_), .Y(new_n445_));
  NOR4X1   g0396(.A(new_n148_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n446_));
  OR4X1    g0397(.A(new_n446_), .B(new_n174_), .C(new_n127_), .D(new_n121_), .Y(new_n447_));
  OR2X1    g0398(.A(new_n190_), .B(new_n169_), .Y(new_n448_));
  OR4X1    g0399(.A(new_n388_), .B(new_n363_), .C(new_n322_), .D(new_n337_), .Y(new_n449_));
  OR4X1    g0400(.A(new_n449_), .B(new_n448_), .C(new_n447_), .D(new_n445_), .Y(new_n450_));
  NOR4X1   g0401(.A(new_n450_), .B(new_n444_), .C(new_n436_), .D(new_n428_), .Y(new_n451_));
  OR2X1    g0402(.A(new_n363_), .B(new_n204_), .Y(new_n452_));
  OR2X1    g0403(.A(new_n271_), .B(new_n147_), .Y(new_n453_));
  OR4X1    g0404(.A(new_n453_), .B(new_n452_), .C(new_n389_), .D(new_n277_), .Y(new_n454_));
  OR2X1    g0405(.A(new_n287_), .B(new_n163_), .Y(new_n455_));
  OR4X1    g0406(.A(new_n455_), .B(new_n446_), .C(new_n303_), .D(new_n127_), .Y(new_n456_));
  NOR3X1   g0407(.A(new_n426_), .B(new_n325_), .C(new_n141_), .Y(new_n457_));
  NOR4X1   g0408(.A(new_n256_), .B(new_n193_), .C(new_n192_), .D(new_n174_), .Y(new_n458_));
  NAND2X1  g0409(.A(new_n458_), .B(new_n457_), .Y(new_n459_));
  OR4X1    g0410(.A(new_n358_), .B(new_n253_), .C(new_n172_), .D(new_n157_), .Y(new_n460_));
  OR2X1    g0411(.A(new_n357_), .B(new_n203_), .Y(new_n461_));
  OR4X1    g0412(.A(new_n461_), .B(new_n460_), .C(new_n185_), .D(new_n179_), .Y(new_n462_));
  OR4X1    g0413(.A(new_n462_), .B(new_n459_), .C(new_n456_), .D(new_n454_), .Y(new_n463_));
  OR4X1    g0414(.A(new_n146_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n464_));
  OR4X1    g0415(.A(new_n120_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n465_));
  NAND2X1  g0416(.A(new_n465_), .B(new_n464_), .Y(new_n466_));
  OR4X1    g0417(.A(new_n466_), .B(new_n378_), .C(new_n221_), .D(new_n131_), .Y(new_n467_));
  OR4X1    g0418(.A(new_n108_), .B(new_n92_), .C(new_n78_), .D(new_n70_), .Y(new_n468_));
  NOR3X1   g0419(.A(new_n372_), .B(new_n183_), .C(new_n121_), .Y(new_n469_));
  NOR2X1   g0420(.A(new_n264_), .B(new_n195_), .Y(new_n470_));
  NAND4X1  g0421(.A(new_n470_), .B(new_n469_), .C(new_n468_), .D(new_n285_), .Y(new_n471_));
  OR2X1    g0422(.A(new_n139_), .B(new_n136_), .Y(new_n472_));
  OR2X1    g0423(.A(new_n472_), .B(new_n322_), .Y(new_n473_));
  OR4X1    g0424(.A(new_n348_), .B(new_n347_), .C(new_n332_), .D(new_n330_), .Y(new_n474_));
  OR4X1    g0425(.A(new_n474_), .B(new_n473_), .C(new_n471_), .D(new_n467_), .Y(new_n475_));
  NOR3X1   g0426(.A(new_n430_), .B(new_n379_), .C(new_n180_), .Y(new_n476_));
  NOR3X1   g0427(.A(new_n175_), .B(new_n155_), .C(new_n123_), .Y(new_n477_));
  NOR3X1   g0428(.A(new_n262_), .B(new_n336_), .C(new_n137_), .Y(new_n478_));
  NAND3X1  g0429(.A(new_n478_), .B(new_n477_), .C(new_n476_), .Y(new_n479_));
  OR4X1    g0430(.A(new_n198_), .B(new_n167_), .C(new_n158_), .D(new_n150_), .Y(new_n480_));
  OR4X1    g0431(.A(new_n480_), .B(new_n314_), .C(new_n283_), .D(new_n134_), .Y(new_n481_));
  OR4X1    g0432(.A(new_n437_), .B(new_n255_), .C(new_n211_), .D(new_n208_), .Y(new_n482_));
  NOR4X1   g0433(.A(new_n148_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n483_));
  OR2X1    g0434(.A(new_n483_), .B(new_n220_), .Y(new_n484_));
  OR4X1    g0435(.A(new_n484_), .B(new_n482_), .C(new_n481_), .D(new_n362_), .Y(new_n485_));
  OR4X1    g0436(.A(new_n485_), .B(new_n479_), .C(new_n475_), .D(new_n463_), .Y(new_n486_));
  NOR4X1   g0437(.A(new_n348_), .B(new_n347_), .C(new_n332_), .D(new_n330_), .Y(new_n487_));
  NOR4X1   g0438(.A(new_n106_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n488_));
  NOR4X1   g0439(.A(new_n488_), .B(new_n219_), .C(new_n168_), .D(new_n157_), .Y(new_n489_));
  NOR3X1   g0440(.A(new_n398_), .B(new_n123_), .C(new_n91_), .Y(new_n490_));
  NAND3X1  g0441(.A(new_n490_), .B(new_n489_), .C(new_n487_), .Y(new_n491_));
  INVX1    g0442(.A(new_n110_), .Y(new_n492_));
  NOR4X1   g0443(.A(new_n208_), .B(new_n207_), .C(new_n165_), .D(new_n162_), .Y(new_n493_));
  NAND3X1  g0444(.A(new_n493_), .B(new_n338_), .C(new_n492_), .Y(new_n494_));
  OR4X1    g0445(.A(new_n430_), .B(new_n426_), .C(new_n385_), .D(new_n164_), .Y(new_n495_));
  OR4X1    g0446(.A(new_n495_), .B(new_n494_), .C(new_n491_), .D(new_n263_), .Y(new_n496_));
  NAND2X1  g0447(.A(new_n440_), .B(new_n154_), .Y(new_n497_));
  OR4X1    g0448(.A(new_n497_), .B(new_n169_), .C(new_n163_), .D(new_n155_), .Y(new_n498_));
  OR4X1    g0449(.A(new_n317_), .B(new_n252_), .C(new_n179_), .D(new_n113_), .Y(new_n499_));
  OR4X1    g0450(.A(new_n499_), .B(new_n379_), .C(new_n397_), .D(new_n270_), .Y(new_n500_));
  OR4X1    g0451(.A(new_n108_), .B(new_n83_), .C(new_n101_), .D(new_n70_), .Y(new_n501_));
  NAND3X1  g0452(.A(new_n501_), .B(new_n464_), .C(new_n468_), .Y(new_n502_));
  OR4X1    g0453(.A(new_n502_), .B(new_n500_), .C(new_n498_), .D(new_n291_), .Y(new_n503_));
  OR4X1    g0454(.A(new_n96_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n504_));
  NAND3X1  g0455(.A(new_n504_), .B(new_n376_), .C(new_n393_), .Y(new_n505_));
  OR4X1    g0456(.A(new_n363_), .B(new_n264_), .C(new_n256_), .D(new_n193_), .Y(new_n506_));
  OR4X1    g0457(.A(new_n506_), .B(new_n505_), .C(new_n322_), .D(new_n265_), .Y(new_n507_));
  OR4X1    g0458(.A(new_n507_), .B(new_n503_), .C(new_n496_), .D(new_n307_), .Y(new_n508_));
  AOI21X1  g0459(.A0(new_n508_), .A1(new_n486_), .B0(new_n451_), .Y(new_n509_));
  INVX1    g0460(.A(\a[7] ), .Y(new_n510_));
  AND2X1   g0461(.A(new_n52_), .B(new_n50_), .Y(new_n511_));
  XOR2X1   g0462(.A(new_n511_), .B(new_n510_), .Y(new_n512_));
  NOR3X1   g0463(.A(new_n512_), .B(new_n509_), .C(new_n401_), .Y(new_n513_));
  OAI21X1  g0464(.A0(new_n512_), .A1(new_n401_), .B0(new_n509_), .Y(new_n514_));
  AND2X1   g0465(.A(\a[22] ), .B(\a[8] ), .Y(new_n515_));
  NOR3X1   g0466(.A(new_n52_), .B(\a[8] ), .C(\a[7] ), .Y(new_n516_));
  NOR2X1   g0467(.A(new_n516_), .B(\a[22] ), .Y(new_n517_));
  OAI21X1  g0468(.A0(new_n52_), .A1(\a[7] ), .B0(\a[8] ), .Y(new_n518_));
  AOI21X1  g0469(.A0(new_n518_), .A1(new_n517_), .B0(new_n515_), .Y(new_n519_));
  NOR2X1   g0470(.A(new_n519_), .B(new_n401_), .Y(new_n520_));
  AOI21X1  g0471(.A0(new_n520_), .A1(new_n514_), .B0(new_n513_), .Y(new_n521_));
  OR4X1    g0472(.A(new_n521_), .B(new_n415_), .C(new_n414_), .D(new_n408_), .Y(new_n522_));
  AOI21X1  g0473(.A0(new_n87_), .A1(new_n85_), .B0(new_n86_), .Y(new_n523_));
  NAND2X1  g0474(.A(new_n88_), .B(new_n50_), .Y(new_n524_));
  OAI22X1  g0475(.A0(new_n524_), .A1(new_n523_), .B0(new_n50_), .B1(new_n86_), .Y(new_n525_));
  OR4X1    g0476(.A(new_n450_), .B(new_n444_), .C(new_n436_), .D(new_n428_), .Y(new_n526_));
  NOR4X1   g0477(.A(new_n124_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n527_));
  OR4X1    g0478(.A(new_n527_), .B(new_n304_), .C(new_n259_), .D(new_n132_), .Y(new_n528_));
  OR2X1    g0479(.A(new_n358_), .B(new_n131_), .Y(new_n529_));
  OR2X1    g0480(.A(new_n219_), .B(new_n173_), .Y(new_n530_));
  OR4X1    g0481(.A(new_n530_), .B(new_n396_), .C(new_n529_), .D(new_n186_), .Y(new_n531_));
  OR2X1    g0482(.A(new_n531_), .B(new_n528_), .Y(new_n532_));
  OR4X1    g0483(.A(new_n532_), .B(new_n500_), .C(new_n430_), .D(new_n262_), .Y(new_n533_));
  OR4X1    g0484(.A(new_n363_), .B(new_n303_), .C(new_n261_), .D(new_n121_), .Y(new_n534_));
  INVX1    g0485(.A(new_n221_), .Y(new_n535_));
  INVX1    g0486(.A(new_n330_), .Y(new_n536_));
  INVX1    g0487(.A(new_n398_), .Y(new_n537_));
  NAND3X1  g0488(.A(new_n537_), .B(new_n536_), .C(new_n535_), .Y(new_n538_));
  OR4X1    g0489(.A(new_n332_), .B(new_n172_), .C(new_n170_), .D(new_n91_), .Y(new_n539_));
  OR2X1    g0490(.A(new_n189_), .B(new_n168_), .Y(new_n540_));
  OR2X1    g0491(.A(new_n540_), .B(new_n147_), .Y(new_n541_));
  OR4X1    g0492(.A(new_n541_), .B(new_n539_), .C(new_n538_), .D(new_n289_), .Y(new_n542_));
  OR4X1    g0493(.A(new_n542_), .B(new_n534_), .C(new_n202_), .D(new_n198_), .Y(new_n543_));
  OR4X1    g0494(.A(new_n140_), .B(new_n90_), .C(new_n92_), .D(new_n78_), .Y(new_n544_));
  OR4X1    g0495(.A(new_n346_), .B(new_n211_), .C(new_n183_), .D(new_n182_), .Y(new_n545_));
  OR2X1    g0496(.A(new_n437_), .B(new_n145_), .Y(new_n546_));
  NAND2X1  g0497(.A(new_n465_), .B(new_n278_), .Y(new_n547_));
  NOR3X1   g0498(.A(new_n547_), .B(new_n546_), .C(new_n545_), .Y(new_n548_));
  NAND3X1  g0499(.A(new_n548_), .B(new_n339_), .C(new_n544_), .Y(new_n549_));
  OR4X1    g0500(.A(new_n372_), .B(new_n205_), .C(new_n157_), .D(new_n107_), .Y(new_n550_));
  NOR4X1   g0501(.A(new_n115_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n551_));
  OR4X1    g0502(.A(new_n551_), .B(new_n220_), .C(new_n193_), .D(new_n164_), .Y(new_n552_));
  OR4X1    g0503(.A(new_n315_), .B(new_n174_), .C(new_n139_), .D(new_n110_), .Y(new_n553_));
  OR4X1    g0504(.A(new_n325_), .B(new_n283_), .C(new_n281_), .D(new_n162_), .Y(new_n554_));
  OR4X1    g0505(.A(new_n554_), .B(new_n553_), .C(new_n552_), .D(new_n550_), .Y(new_n555_));
  NOR4X1   g0506(.A(new_n555_), .B(new_n549_), .C(new_n543_), .D(new_n533_), .Y(new_n556_));
  XOR2X1   g0507(.A(new_n556_), .B(new_n526_), .Y(new_n557_));
  OR2X1    g0508(.A(new_n305_), .B(new_n116_), .Y(new_n558_));
  OR4X1    g0509(.A(new_n106_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n559_));
  OR4X1    g0510(.A(new_n106_), .B(new_n108_), .C(new_n83_), .D(new_n101_), .Y(new_n560_));
  OR4X1    g0511(.A(new_n112_), .B(new_n90_), .C(new_n83_), .D(new_n78_), .Y(new_n561_));
  NAND3X1  g0512(.A(new_n561_), .B(new_n560_), .C(new_n559_), .Y(new_n562_));
  OR4X1    g0513(.A(new_n562_), .B(new_n255_), .C(new_n252_), .D(new_n219_), .Y(new_n563_));
  OR2X1    g0514(.A(new_n221_), .B(new_n113_), .Y(new_n564_));
  OR2X1    g0515(.A(new_n564_), .B(new_n262_), .Y(new_n565_));
  NOR3X1   g0516(.A(new_n565_), .B(new_n563_), .C(new_n473_), .Y(new_n566_));
  INVX1    g0517(.A(new_n566_), .Y(new_n567_));
  OR2X1    g0518(.A(new_n294_), .B(new_n141_), .Y(new_n568_));
  OR4X1    g0519(.A(new_n568_), .B(new_n321_), .C(new_n213_), .D(new_n125_), .Y(new_n569_));
  OR4X1    g0520(.A(new_n569_), .B(new_n567_), .C(new_n171_), .D(new_n166_), .Y(new_n570_));
  OR2X1    g0521(.A(new_n332_), .B(new_n292_), .Y(new_n571_));
  OR2X1    g0522(.A(new_n571_), .B(new_n269_), .Y(new_n572_));
  OR4X1    g0523(.A(new_n488_), .B(new_n317_), .C(new_n247_), .D(new_n134_), .Y(new_n573_));
  OAI21X1  g0524(.A0(new_n133_), .A1(new_n333_), .B0(new_n465_), .Y(new_n574_));
  OR4X1    g0525(.A(new_n574_), .B(new_n573_), .C(new_n572_), .D(new_n426_), .Y(new_n575_));
  OR2X1    g0526(.A(new_n205_), .B(new_n157_), .Y(new_n576_));
  OR4X1    g0527(.A(new_n576_), .B(new_n265_), .C(new_n249_), .D(new_n204_), .Y(new_n577_));
  NOR3X1   g0528(.A(new_n430_), .B(new_n158_), .C(new_n110_), .Y(new_n578_));
  NOR2X1   g0529(.A(new_n132_), .B(new_n131_), .Y(new_n579_));
  NAND2X1  g0530(.A(new_n579_), .B(new_n578_), .Y(new_n580_));
  NOR4X1   g0531(.A(new_n385_), .B(new_n329_), .C(new_n287_), .D(new_n147_), .Y(new_n581_));
  NAND2X1  g0532(.A(new_n581_), .B(new_n477_), .Y(new_n582_));
  OR4X1    g0533(.A(new_n582_), .B(new_n580_), .C(new_n577_), .D(new_n575_), .Y(new_n583_));
  OR4X1    g0534(.A(new_n583_), .B(new_n570_), .C(new_n558_), .D(new_n201_), .Y(new_n584_));
  AOI21X1  g0535(.A0(new_n556_), .A1(new_n451_), .B0(new_n584_), .Y(new_n585_));
  NOR2X1   g0536(.A(new_n585_), .B(new_n557_), .Y(new_n586_));
  OR2X1    g0537(.A(new_n556_), .B(new_n451_), .Y(new_n587_));
  AOI21X1  g0538(.A0(new_n587_), .A1(new_n584_), .B0(new_n557_), .Y(new_n588_));
  MX2X1    g0539(.A(new_n588_), .B(new_n586_), .S0(new_n525_), .Y(new_n589_));
  AND2X1   g0540(.A(new_n54_), .B(new_n50_), .Y(new_n590_));
  XOR2X1   g0541(.A(new_n590_), .B(new_n85_), .Y(new_n591_));
  INVX1    g0542(.A(new_n557_), .Y(new_n592_));
  AND2X1   g0543(.A(new_n587_), .B(new_n584_), .Y(new_n593_));
  NOR2X1   g0544(.A(new_n593_), .B(new_n592_), .Y(new_n594_));
  NOR2X1   g0545(.A(new_n585_), .B(new_n592_), .Y(new_n595_));
  MX2X1    g0546(.A(new_n595_), .B(new_n594_), .S0(new_n591_), .Y(new_n596_));
  NOR2X1   g0547(.A(new_n596_), .B(new_n589_), .Y(new_n597_));
  NAND2X1  g0548(.A(\a[22] ), .B(\a[12] ), .Y(new_n598_));
  INVX1    g0549(.A(\a[12] ), .Y(new_n599_));
  NOR3X1   g0550(.A(new_n53_), .B(\a[11] ), .C(\a[10] ), .Y(new_n600_));
  OAI21X1  g0551(.A0(new_n600_), .A1(new_n599_), .B0(new_n590_), .Y(new_n601_));
  AND2X1   g0552(.A(new_n601_), .B(new_n598_), .Y(new_n602_));
  OR2X1    g0553(.A(new_n314_), .B(new_n247_), .Y(new_n603_));
  OR4X1    g0554(.A(new_n129_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n604_));
  INVX1    g0555(.A(new_n604_), .Y(new_n605_));
  OR4X1    g0556(.A(new_n605_), .B(new_n256_), .C(new_n155_), .D(new_n145_), .Y(new_n606_));
  OR2X1    g0557(.A(new_n204_), .B(new_n127_), .Y(new_n607_));
  OR2X1    g0558(.A(new_n607_), .B(new_n385_), .Y(new_n608_));
  OR4X1    g0559(.A(new_n213_), .B(new_n190_), .C(new_n170_), .D(new_n150_), .Y(new_n609_));
  OR4X1    g0560(.A(new_n609_), .B(new_n608_), .C(new_n606_), .D(new_n603_), .Y(new_n610_));
  OR4X1    g0561(.A(new_n322_), .B(new_n197_), .C(new_n193_), .D(new_n125_), .Y(new_n611_));
  OR2X1    g0562(.A(new_n279_), .B(new_n121_), .Y(new_n612_));
  OR4X1    g0563(.A(new_n612_), .B(new_n611_), .C(new_n538_), .D(new_n209_), .Y(new_n613_));
  OR4X1    g0564(.A(new_n357_), .B(new_n437_), .C(new_n164_), .D(new_n157_), .Y(new_n614_));
  OR4X1    g0565(.A(new_n614_), .B(new_n273_), .C(new_n249_), .D(new_n165_), .Y(new_n615_));
  INVX1    g0566(.A(new_n355_), .Y(new_n616_));
  OR4X1    g0567(.A(new_n426_), .B(new_n321_), .C(new_n168_), .D(new_n167_), .Y(new_n617_));
  OR2X1    g0568(.A(new_n248_), .B(new_n149_), .Y(new_n618_));
  OR4X1    g0569(.A(new_n618_), .B(new_n617_), .C(new_n616_), .D(new_n329_), .Y(new_n619_));
  OR4X1    g0570(.A(new_n619_), .B(new_n615_), .C(new_n416_), .D(new_n315_), .Y(new_n620_));
  OR2X1    g0571(.A(new_n620_), .B(new_n613_), .Y(new_n621_));
  NOR4X1   g0572(.A(new_n621_), .B(new_n610_), .C(new_n533_), .D(new_n298_), .Y(new_n622_));
  XOR2X1   g0573(.A(new_n622_), .B(new_n584_), .Y(new_n623_));
  INVX1    g0574(.A(new_n350_), .Y(new_n624_));
  NOR4X1   g0575(.A(new_n583_), .B(new_n570_), .C(new_n558_), .D(new_n201_), .Y(new_n625_));
  AOI21X1  g0576(.A0(new_n622_), .A1(new_n625_), .B0(new_n624_), .Y(new_n626_));
  NOR2X1   g0577(.A(new_n626_), .B(new_n623_), .Y(new_n627_));
  INVX1    g0578(.A(new_n622_), .Y(new_n628_));
  AOI21X1  g0579(.A0(new_n628_), .A1(new_n584_), .B0(new_n350_), .Y(new_n629_));
  NOR2X1   g0580(.A(new_n629_), .B(new_n623_), .Y(new_n630_));
  MX2X1    g0581(.A(new_n627_), .B(new_n630_), .S0(new_n602_), .Y(new_n631_));
  INVX1    g0582(.A(new_n623_), .Y(new_n632_));
  NOR2X1   g0583(.A(new_n629_), .B(new_n632_), .Y(new_n633_));
  NOR2X1   g0584(.A(new_n626_), .B(new_n632_), .Y(new_n634_));
  MX2X1    g0585(.A(new_n634_), .B(new_n633_), .S0(new_n312_), .Y(new_n635_));
  NOR2X1   g0586(.A(new_n635_), .B(new_n631_), .Y(new_n636_));
  MX2X1    g0587(.A(new_n407_), .B(new_n404_), .S0(new_n413_), .Y(new_n637_));
  OR2X1    g0588(.A(new_n406_), .B(new_n367_), .Y(new_n638_));
  INVX1    g0589(.A(new_n638_), .Y(new_n639_));
  NOR2X1   g0590(.A(new_n403_), .B(new_n367_), .Y(new_n640_));
  XOR2X1   g0591(.A(new_n517_), .B(\a[9] ), .Y(new_n641_));
  INVX1    g0592(.A(new_n641_), .Y(new_n642_));
  MX2X1    g0593(.A(new_n640_), .B(new_n639_), .S0(new_n642_), .Y(new_n643_));
  INVX1    g0594(.A(new_n597_), .Y(new_n644_));
  XOR2X1   g0595(.A(new_n636_), .B(new_n644_), .Y(new_n645_));
  NOR3X1   g0596(.A(new_n645_), .B(new_n643_), .C(new_n637_), .Y(new_n646_));
  AOI21X1  g0597(.A0(new_n636_), .A1(new_n597_), .B0(new_n646_), .Y(new_n647_));
  NOR3X1   g0598(.A(new_n415_), .B(new_n414_), .C(new_n408_), .Y(new_n648_));
  XOR2X1   g0599(.A(new_n521_), .B(new_n648_), .Y(new_n649_));
  OAI21X1  g0600(.A0(new_n649_), .A1(new_n647_), .B0(new_n522_), .Y(new_n650_));
  NOR2X1   g0601(.A(new_n642_), .B(new_n401_), .Y(new_n651_));
  INVX1    g0602(.A(new_n651_), .Y(new_n652_));
  XOR2X1   g0603(.A(new_n652_), .B(new_n593_), .Y(new_n653_));
  NOR2X1   g0604(.A(new_n412_), .B(new_n401_), .Y(new_n654_));
  XOR2X1   g0605(.A(new_n654_), .B(new_n653_), .Y(new_n655_));
  AND2X1   g0606(.A(new_n655_), .B(new_n650_), .Y(new_n656_));
  XOR2X1   g0607(.A(new_n655_), .B(new_n650_), .Y(new_n657_));
  AOI22X1  g0608(.A0(new_n587_), .A1(new_n584_), .B0(new_n557_), .B1(new_n525_), .Y(new_n658_));
  AOI21X1  g0609(.A0(new_n595_), .A1(new_n525_), .B0(new_n658_), .Y(new_n659_));
  AND2X1   g0610(.A(new_n659_), .B(new_n652_), .Y(new_n660_));
  MX2X1    g0611(.A(new_n627_), .B(new_n630_), .S0(new_n591_), .Y(new_n661_));
  MX2X1    g0612(.A(new_n634_), .B(new_n633_), .S0(new_n602_), .Y(new_n662_));
  NOR2X1   g0613(.A(new_n662_), .B(new_n661_), .Y(new_n663_));
  XOR2X1   g0614(.A(new_n659_), .B(new_n652_), .Y(new_n664_));
  AND2X1   g0615(.A(new_n664_), .B(new_n663_), .Y(new_n665_));
  OR2X1    g0616(.A(new_n665_), .B(new_n660_), .Y(new_n666_));
  MX2X1    g0617(.A(new_n630_), .B(new_n627_), .S0(new_n525_), .Y(new_n667_));
  MX2X1    g0618(.A(new_n634_), .B(new_n633_), .S0(new_n591_), .Y(new_n668_));
  MX2X1    g0619(.A(new_n404_), .B(new_n407_), .S0(new_n602_), .Y(new_n669_));
  MX2X1    g0620(.A(new_n640_), .B(new_n639_), .S0(new_n312_), .Y(new_n670_));
  NOR4X1   g0621(.A(new_n670_), .B(new_n669_), .C(new_n668_), .D(new_n667_), .Y(new_n671_));
  INVX1    g0622(.A(new_n671_), .Y(new_n672_));
  OAI22X1  g0623(.A0(new_n670_), .A1(new_n669_), .B0(new_n668_), .B1(new_n667_), .Y(new_n673_));
  AND2X1   g0624(.A(new_n673_), .B(new_n672_), .Y(new_n674_));
  XOR2X1   g0625(.A(new_n674_), .B(new_n666_), .Y(new_n675_));
  AOI21X1  g0626(.A0(new_n675_), .A1(new_n657_), .B0(new_n656_), .Y(new_n676_));
  NOR2X1   g0627(.A(new_n652_), .B(new_n593_), .Y(new_n677_));
  AOI21X1  g0628(.A0(new_n654_), .A1(new_n653_), .B0(new_n677_), .Y(new_n678_));
  AOI21X1  g0629(.A0(new_n673_), .A1(new_n666_), .B0(new_n671_), .Y(new_n679_));
  XOR2X1   g0630(.A(new_n679_), .B(new_n678_), .Y(new_n680_));
  INVX1    g0631(.A(new_n680_), .Y(new_n681_));
  MX2X1    g0632(.A(new_n404_), .B(new_n407_), .S0(new_n591_), .Y(new_n682_));
  MX2X1    g0633(.A(new_n640_), .B(new_n639_), .S0(new_n602_), .Y(new_n683_));
  NOR2X1   g0634(.A(new_n683_), .B(new_n682_), .Y(new_n684_));
  NOR2X1   g0635(.A(new_n401_), .B(new_n312_), .Y(new_n685_));
  INVX1    g0636(.A(new_n685_), .Y(new_n686_));
  AOI21X1  g0637(.A0(new_n623_), .A1(new_n525_), .B0(new_n629_), .Y(new_n687_));
  AOI21X1  g0638(.A0(new_n634_), .A1(new_n525_), .B0(new_n687_), .Y(new_n688_));
  XOR2X1   g0639(.A(new_n688_), .B(new_n686_), .Y(new_n689_));
  XOR2X1   g0640(.A(new_n689_), .B(new_n684_), .Y(new_n690_));
  XOR2X1   g0641(.A(new_n690_), .B(new_n681_), .Y(new_n691_));
  XOR2X1   g0642(.A(new_n691_), .B(new_n676_), .Y(new_n692_));
  INVX1    g0643(.A(new_n692_), .Y(new_n693_));
  MX2X1    g0644(.A(new_n630_), .B(new_n627_), .S0(new_n313_), .Y(new_n694_));
  MX2X1    g0645(.A(new_n633_), .B(new_n634_), .S0(new_n413_), .Y(new_n695_));
  MX2X1    g0646(.A(new_n404_), .B(new_n407_), .S0(new_n642_), .Y(new_n696_));
  MX2X1    g0647(.A(new_n640_), .B(new_n639_), .S0(new_n519_), .Y(new_n697_));
  NOR4X1   g0648(.A(new_n697_), .B(new_n696_), .C(new_n695_), .D(new_n694_), .Y(new_n698_));
  NOR4X1   g0649(.A(new_n485_), .B(new_n479_), .C(new_n475_), .D(new_n463_), .Y(new_n699_));
  OR4X1    g0650(.A(new_n90_), .B(new_n83_), .C(new_n78_), .D(new_n70_), .Y(new_n700_));
  AND2X1   g0651(.A(new_n441_), .B(new_n276_), .Y(new_n701_));
  NOR2X1   g0652(.A(new_n551_), .B(new_n196_), .Y(new_n702_));
  NAND4X1  g0653(.A(new_n702_), .B(new_n604_), .C(new_n701_), .D(new_n700_), .Y(new_n703_));
  OR4X1    g0654(.A(new_n483_), .B(new_n220_), .C(new_n198_), .D(new_n174_), .Y(new_n704_));
  OR4X1    g0655(.A(new_n704_), .B(new_n426_), .C(new_n214_), .D(new_n173_), .Y(new_n705_));
  OR4X1    g0656(.A(new_n303_), .B(new_n205_), .C(new_n158_), .D(new_n137_), .Y(new_n706_));
  OR4X1    g0657(.A(new_n706_), .B(new_n337_), .C(new_n336_), .D(new_n97_), .Y(new_n707_));
  OR4X1    g0658(.A(new_n707_), .B(new_n705_), .C(new_n703_), .D(new_n569_), .Y(new_n708_));
  OR4X1    g0659(.A(new_n372_), .B(new_n325_), .C(new_n292_), .D(new_n280_), .Y(new_n709_));
  OR4X1    g0660(.A(new_n190_), .B(new_n168_), .C(new_n167_), .D(new_n155_), .Y(new_n710_));
  OR4X1    g0661(.A(new_n710_), .B(new_n709_), .C(new_n546_), .D(new_n461_), .Y(new_n711_));
  OR2X1    g0662(.A(new_n348_), .B(new_n281_), .Y(new_n712_));
  OR4X1    g0663(.A(new_n446_), .B(new_n165_), .C(new_n150_), .D(new_n134_), .Y(new_n713_));
  OR4X1    g0664(.A(new_n713_), .B(new_n712_), .C(new_n358_), .D(new_n331_), .Y(new_n714_));
  NOR4X1   g0665(.A(new_n714_), .B(new_n711_), .C(new_n708_), .D(new_n267_), .Y(new_n715_));
  OR4X1    g0666(.A(new_n426_), .B(new_n372_), .C(new_n283_), .D(new_n252_), .Y(new_n716_));
  OR2X1    g0667(.A(new_n159_), .B(new_n150_), .Y(new_n717_));
  OR4X1    g0668(.A(new_n717_), .B(new_n716_), .C(new_n455_), .D(new_n273_), .Y(new_n718_));
  OR4X1    g0669(.A(new_n211_), .B(new_n179_), .C(new_n175_), .D(new_n130_), .Y(new_n719_));
  OR2X1    g0670(.A(new_n483_), .B(new_n551_), .Y(new_n720_));
  OR4X1    g0671(.A(new_n720_), .B(new_n562_), .C(new_n505_), .D(new_n446_), .Y(new_n721_));
  OR4X1    g0672(.A(new_n721_), .B(new_n719_), .C(new_n718_), .D(new_n319_), .Y(new_n722_));
  NOR3X1   g0673(.A(new_n315_), .B(new_n188_), .C(new_n116_), .Y(new_n723_));
  NOR3X1   g0674(.A(new_n527_), .B(new_n363_), .C(new_n149_), .Y(new_n724_));
  NAND3X1  g0675(.A(new_n724_), .B(new_n723_), .C(new_n476_), .Y(new_n725_));
  OR2X1    g0676(.A(new_n220_), .B(new_n164_), .Y(new_n726_));
  NAND2X1  g0677(.A(new_n604_), .B(new_n700_), .Y(new_n727_));
  OR2X1    g0678(.A(new_n262_), .B(new_n123_), .Y(new_n728_));
  OR4X1    g0679(.A(new_n728_), .B(new_n727_), .C(new_n726_), .D(new_n334_), .Y(new_n729_));
  OR4X1    g0680(.A(new_n219_), .B(new_n184_), .C(new_n170_), .D(new_n157_), .Y(new_n730_));
  OR2X1    g0681(.A(new_n730_), .B(new_n389_), .Y(new_n731_));
  OR4X1    g0682(.A(new_n731_), .B(new_n729_), .C(new_n725_), .D(new_n707_), .Y(new_n732_));
  OR4X1    g0683(.A(new_n259_), .B(new_n213_), .C(new_n203_), .D(new_n192_), .Y(new_n733_));
  OR4X1    g0684(.A(new_n341_), .B(new_n251_), .C(new_n185_), .D(new_n121_), .Y(new_n734_));
  NOR4X1   g0685(.A(new_n305_), .B(new_n304_), .C(new_n281_), .D(new_n269_), .Y(new_n735_));
  NAND3X1  g0686(.A(new_n735_), .B(new_n355_), .C(new_n301_), .Y(new_n736_));
  OR4X1    g0687(.A(new_n419_), .B(new_n358_), .C(new_n291_), .D(new_n131_), .Y(new_n737_));
  OR4X1    g0688(.A(new_n737_), .B(new_n736_), .C(new_n734_), .D(new_n733_), .Y(new_n738_));
  NOR3X1   g0689(.A(new_n738_), .B(new_n732_), .C(new_n722_), .Y(new_n739_));
  AND2X1   g0690(.A(new_n715_), .B(new_n699_), .Y(new_n740_));
  OR4X1    g0691(.A(new_n730_), .B(new_n729_), .C(new_n707_), .D(new_n389_), .Y(new_n741_));
  OR4X1    g0692(.A(new_n738_), .B(new_n741_), .C(new_n725_), .D(new_n722_), .Y(new_n742_));
  NOR3X1   g0693(.A(new_n742_), .B(new_n715_), .C(new_n699_), .Y(new_n743_));
  INVX1    g0694(.A(new_n743_), .Y(new_n744_));
  NAND2X1  g0695(.A(\a[22] ), .B(\a[6] ), .Y(new_n745_));
  INVX1    g0696(.A(\a[6] ), .Y(new_n746_));
  NOR3X1   g0697(.A(new_n51_), .B(\a[5] ), .C(\a[4] ), .Y(new_n747_));
  OAI21X1  g0698(.A0(new_n747_), .A1(new_n746_), .B0(new_n511_), .Y(new_n748_));
  AND2X1   g0699(.A(new_n748_), .B(new_n745_), .Y(new_n749_));
  NOR2X1   g0700(.A(new_n749_), .B(new_n401_), .Y(new_n750_));
  AOI21X1  g0701(.A0(new_n750_), .A1(new_n744_), .B0(new_n740_), .Y(new_n751_));
  INVX1    g0702(.A(new_n751_), .Y(new_n752_));
  OAI22X1  g0703(.A0(new_n697_), .A1(new_n696_), .B0(new_n695_), .B1(new_n694_), .Y(new_n753_));
  AOI21X1  g0704(.A0(new_n753_), .A1(new_n752_), .B0(new_n698_), .Y(new_n754_));
  NOR2X1   g0705(.A(new_n512_), .B(new_n401_), .Y(new_n755_));
  INVX1    g0706(.A(new_n755_), .Y(new_n756_));
  NOR4X1   g0707(.A(new_n507_), .B(new_n503_), .C(new_n496_), .D(new_n307_), .Y(new_n757_));
  XOR2X1   g0708(.A(new_n757_), .B(new_n699_), .Y(new_n758_));
  AOI21X1  g0709(.A0(new_n757_), .A1(new_n699_), .B0(new_n526_), .Y(new_n759_));
  NOR2X1   g0710(.A(new_n759_), .B(new_n758_), .Y(new_n760_));
  XOR2X1   g0711(.A(new_n757_), .B(new_n486_), .Y(new_n761_));
  AOI21X1  g0712(.A0(new_n761_), .A1(new_n525_), .B0(new_n509_), .Y(new_n762_));
  AOI21X1  g0713(.A0(new_n760_), .A1(new_n525_), .B0(new_n762_), .Y(new_n763_));
  AND2X1   g0714(.A(new_n763_), .B(new_n756_), .Y(new_n764_));
  MX2X1    g0715(.A(new_n586_), .B(new_n588_), .S0(new_n591_), .Y(new_n765_));
  MX2X1    g0716(.A(new_n595_), .B(new_n594_), .S0(new_n602_), .Y(new_n766_));
  NOR2X1   g0717(.A(new_n766_), .B(new_n765_), .Y(new_n767_));
  XOR2X1   g0718(.A(new_n763_), .B(new_n756_), .Y(new_n768_));
  AOI21X1  g0719(.A0(new_n768_), .A1(new_n767_), .B0(new_n764_), .Y(new_n769_));
  OR2X1    g0720(.A(new_n769_), .B(new_n754_), .Y(new_n770_));
  XOR2X1   g0721(.A(new_n769_), .B(new_n754_), .Y(new_n771_));
  INVX1    g0722(.A(new_n771_), .Y(new_n772_));
  XOR2X1   g0723(.A(new_n755_), .B(new_n509_), .Y(new_n773_));
  XOR2X1   g0724(.A(new_n520_), .B(new_n773_), .Y(new_n774_));
  OAI21X1  g0725(.A0(new_n774_), .A1(new_n772_), .B0(new_n770_), .Y(new_n775_));
  XOR2X1   g0726(.A(new_n664_), .B(new_n663_), .Y(new_n776_));
  NAND2X1  g0727(.A(new_n776_), .B(new_n775_), .Y(new_n777_));
  XOR2X1   g0728(.A(new_n649_), .B(new_n647_), .Y(new_n778_));
  INVX1    g0729(.A(new_n778_), .Y(new_n779_));
  NOR2X1   g0730(.A(new_n776_), .B(new_n775_), .Y(new_n780_));
  OAI21X1  g0731(.A0(new_n780_), .A1(new_n779_), .B0(new_n777_), .Y(new_n781_));
  XOR2X1   g0732(.A(new_n675_), .B(new_n657_), .Y(new_n782_));
  AND2X1   g0733(.A(new_n782_), .B(new_n781_), .Y(new_n783_));
  XOR2X1   g0734(.A(new_n776_), .B(new_n775_), .Y(new_n784_));
  XOR2X1   g0735(.A(new_n784_), .B(new_n779_), .Y(new_n785_));
  MX2X1    g0736(.A(new_n630_), .B(new_n627_), .S0(new_n413_), .Y(new_n786_));
  MX2X1    g0737(.A(new_n634_), .B(new_n633_), .S0(new_n642_), .Y(new_n787_));
  NOR2X1   g0738(.A(new_n787_), .B(new_n786_), .Y(new_n788_));
  MX2X1    g0739(.A(new_n404_), .B(new_n407_), .S0(new_n519_), .Y(new_n789_));
  INVX1    g0740(.A(new_n512_), .Y(new_n790_));
  MX2X1    g0741(.A(new_n639_), .B(new_n640_), .S0(new_n790_), .Y(new_n791_));
  NOR2X1   g0742(.A(new_n791_), .B(new_n789_), .Y(new_n792_));
  INVX1    g0743(.A(new_n525_), .Y(new_n793_));
  NOR2X1   g0744(.A(new_n761_), .B(new_n509_), .Y(new_n794_));
  NOR2X1   g0745(.A(new_n759_), .B(new_n761_), .Y(new_n795_));
  MX2X1    g0746(.A(new_n795_), .B(new_n794_), .S0(new_n793_), .Y(new_n796_));
  NOR2X1   g0747(.A(new_n758_), .B(new_n509_), .Y(new_n797_));
  MX2X1    g0748(.A(new_n760_), .B(new_n797_), .S0(new_n591_), .Y(new_n798_));
  OR2X1    g0749(.A(new_n798_), .B(new_n796_), .Y(new_n799_));
  INVX1    g0750(.A(new_n792_), .Y(new_n800_));
  XOR2X1   g0751(.A(new_n800_), .B(new_n788_), .Y(new_n801_));
  NOR2X1   g0752(.A(new_n801_), .B(new_n799_), .Y(new_n802_));
  AOI21X1  g0753(.A0(new_n792_), .A1(new_n788_), .B0(new_n802_), .Y(new_n803_));
  INVX1    g0754(.A(new_n803_), .Y(new_n804_));
  XOR2X1   g0755(.A(new_n768_), .B(new_n767_), .Y(new_n805_));
  AND2X1   g0756(.A(new_n805_), .B(new_n804_), .Y(new_n806_));
  XOR2X1   g0757(.A(new_n805_), .B(new_n803_), .Y(new_n807_));
  INVX1    g0758(.A(new_n807_), .Y(new_n808_));
  INVX1    g0759(.A(new_n698_), .Y(new_n809_));
  AND2X1   g0760(.A(new_n753_), .B(new_n809_), .Y(new_n810_));
  XOR2X1   g0761(.A(new_n810_), .B(new_n752_), .Y(new_n811_));
  AOI21X1  g0762(.A0(new_n811_), .A1(new_n808_), .B0(new_n806_), .Y(new_n812_));
  NOR2X1   g0763(.A(new_n643_), .B(new_n637_), .Y(new_n813_));
  XOR2X1   g0764(.A(new_n645_), .B(new_n813_), .Y(new_n814_));
  NOR2X1   g0765(.A(new_n814_), .B(new_n812_), .Y(new_n815_));
  XOR2X1   g0766(.A(new_n814_), .B(new_n812_), .Y(new_n816_));
  XOR2X1   g0767(.A(new_n774_), .B(new_n771_), .Y(new_n817_));
  INVX1    g0768(.A(new_n817_), .Y(new_n818_));
  AOI21X1  g0769(.A0(new_n818_), .A1(new_n816_), .B0(new_n815_), .Y(new_n819_));
  OR2X1    g0770(.A(new_n819_), .B(new_n785_), .Y(new_n820_));
  INVX1    g0771(.A(new_n785_), .Y(new_n821_));
  XOR2X1   g0772(.A(new_n819_), .B(new_n821_), .Y(new_n822_));
  MX2X1    g0773(.A(new_n586_), .B(new_n588_), .S0(new_n602_), .Y(new_n823_));
  MX2X1    g0774(.A(new_n595_), .B(new_n594_), .S0(new_n312_), .Y(new_n824_));
  OR4X1    g0775(.A(new_n749_), .B(new_n743_), .C(new_n740_), .D(new_n401_), .Y(new_n825_));
  AOI22X1  g0776(.A0(new_n751_), .A1(new_n744_), .B0(new_n825_), .B1(new_n750_), .Y(new_n826_));
  NOR3X1   g0777(.A(new_n826_), .B(new_n824_), .C(new_n823_), .Y(new_n827_));
  NOR3X1   g0778(.A(new_n715_), .B(new_n401_), .C(new_n229_), .Y(new_n828_));
  OR4X1    g0779(.A(new_n714_), .B(new_n711_), .C(new_n708_), .D(new_n267_), .Y(new_n829_));
  XOR2X1   g0780(.A(new_n739_), .B(new_n829_), .Y(new_n830_));
  OAI21X1  g0781(.A0(new_n742_), .A1(new_n829_), .B0(new_n699_), .Y(new_n831_));
  NAND3X1  g0782(.A(new_n831_), .B(new_n830_), .C(new_n525_), .Y(new_n832_));
  OAI21X1  g0783(.A0(new_n739_), .A1(new_n715_), .B0(new_n486_), .Y(new_n833_));
  XOR2X1   g0784(.A(new_n739_), .B(new_n715_), .Y(new_n834_));
  OAI21X1  g0785(.A0(new_n834_), .A1(new_n793_), .B0(new_n833_), .Y(new_n835_));
  AND2X1   g0786(.A(new_n835_), .B(new_n832_), .Y(new_n836_));
  AOI21X1  g0787(.A0(new_n402_), .A1(new_n230_), .B0(new_n829_), .Y(new_n837_));
  INVX1    g0788(.A(new_n837_), .Y(new_n838_));
  AOI21X1  g0789(.A0(new_n838_), .A1(new_n836_), .B0(new_n828_), .Y(new_n839_));
  INVX1    g0790(.A(new_n839_), .Y(new_n840_));
  OR2X1    g0791(.A(new_n824_), .B(new_n823_), .Y(new_n841_));
  XOR2X1   g0792(.A(new_n826_), .B(new_n841_), .Y(new_n842_));
  AOI21X1  g0793(.A0(new_n842_), .A1(new_n840_), .B0(new_n827_), .Y(new_n843_));
  MX2X1    g0794(.A(new_n795_), .B(new_n794_), .S0(new_n591_), .Y(new_n844_));
  MX2X1    g0795(.A(new_n760_), .B(new_n797_), .S0(new_n602_), .Y(new_n845_));
  OR2X1    g0796(.A(new_n845_), .B(new_n844_), .Y(new_n846_));
  MX2X1    g0797(.A(new_n588_), .B(new_n586_), .S0(new_n313_), .Y(new_n847_));
  MX2X1    g0798(.A(new_n594_), .B(new_n595_), .S0(new_n413_), .Y(new_n848_));
  NOR3X1   g0799(.A(new_n848_), .B(new_n847_), .C(new_n846_), .Y(new_n849_));
  MX2X1    g0800(.A(new_n627_), .B(new_n630_), .S0(new_n642_), .Y(new_n850_));
  MX2X1    g0801(.A(new_n634_), .B(new_n633_), .S0(new_n519_), .Y(new_n851_));
  NOR2X1   g0802(.A(new_n848_), .B(new_n847_), .Y(new_n852_));
  XOR2X1   g0803(.A(new_n852_), .B(new_n846_), .Y(new_n853_));
  NOR3X1   g0804(.A(new_n853_), .B(new_n851_), .C(new_n850_), .Y(new_n854_));
  OR2X1    g0805(.A(new_n854_), .B(new_n849_), .Y(new_n855_));
  XOR2X1   g0806(.A(new_n801_), .B(new_n799_), .Y(new_n856_));
  AND2X1   g0807(.A(new_n856_), .B(new_n855_), .Y(new_n857_));
  MX2X1    g0808(.A(new_n407_), .B(new_n404_), .S0(new_n790_), .Y(new_n858_));
  MX2X1    g0809(.A(new_n640_), .B(new_n639_), .S0(new_n749_), .Y(new_n859_));
  NOR2X1   g0810(.A(new_n859_), .B(new_n858_), .Y(new_n860_));
  NOR3X1   g0811(.A(new_n715_), .B(new_n401_), .C(new_n233_), .Y(new_n861_));
  AOI21X1  g0812(.A0(new_n742_), .A1(new_n829_), .B0(new_n699_), .Y(new_n862_));
  NOR2X1   g0813(.A(new_n830_), .B(new_n862_), .Y(new_n863_));
  AOI21X1  g0814(.A0(new_n739_), .A1(new_n715_), .B0(new_n486_), .Y(new_n864_));
  NOR2X1   g0815(.A(new_n864_), .B(new_n830_), .Y(new_n865_));
  MX2X1    g0816(.A(new_n865_), .B(new_n863_), .S0(new_n793_), .Y(new_n866_));
  NOR2X1   g0817(.A(new_n864_), .B(new_n834_), .Y(new_n867_));
  NOR2X1   g0818(.A(new_n834_), .B(new_n862_), .Y(new_n868_));
  MX2X1    g0819(.A(new_n867_), .B(new_n868_), .S0(new_n591_), .Y(new_n869_));
  NOR2X1   g0820(.A(new_n401_), .B(new_n233_), .Y(new_n870_));
  XOR2X1   g0821(.A(new_n870_), .B(new_n715_), .Y(new_n871_));
  NOR3X1   g0822(.A(new_n871_), .B(new_n869_), .C(new_n866_), .Y(new_n872_));
  OAI21X1  g0823(.A0(new_n872_), .A1(new_n861_), .B0(new_n860_), .Y(new_n873_));
  NOR2X1   g0824(.A(new_n869_), .B(new_n866_), .Y(new_n874_));
  NOR2X1   g0825(.A(new_n870_), .B(new_n829_), .Y(new_n875_));
  INVX1    g0826(.A(new_n875_), .Y(new_n876_));
  AOI21X1  g0827(.A0(new_n876_), .A1(new_n874_), .B0(new_n861_), .Y(new_n877_));
  XOR2X1   g0828(.A(new_n877_), .B(new_n860_), .Y(new_n878_));
  MX2X1    g0829(.A(new_n588_), .B(new_n586_), .S0(new_n413_), .Y(new_n879_));
  MX2X1    g0830(.A(new_n595_), .B(new_n594_), .S0(new_n642_), .Y(new_n880_));
  MX2X1    g0831(.A(new_n795_), .B(new_n794_), .S0(new_n602_), .Y(new_n881_));
  MX2X1    g0832(.A(new_n797_), .B(new_n760_), .S0(new_n313_), .Y(new_n882_));
  OR2X1    g0833(.A(new_n882_), .B(new_n881_), .Y(new_n883_));
  NOR3X1   g0834(.A(new_n883_), .B(new_n880_), .C(new_n879_), .Y(new_n884_));
  MX2X1    g0835(.A(new_n627_), .B(new_n630_), .S0(new_n519_), .Y(new_n885_));
  MX2X1    g0836(.A(new_n633_), .B(new_n634_), .S0(new_n790_), .Y(new_n886_));
  NOR2X1   g0837(.A(new_n880_), .B(new_n879_), .Y(new_n887_));
  XOR2X1   g0838(.A(new_n883_), .B(new_n887_), .Y(new_n888_));
  NOR3X1   g0839(.A(new_n888_), .B(new_n886_), .C(new_n885_), .Y(new_n889_));
  NOR2X1   g0840(.A(new_n889_), .B(new_n884_), .Y(new_n890_));
  OAI21X1  g0841(.A0(new_n890_), .A1(new_n878_), .B0(new_n873_), .Y(new_n891_));
  XOR2X1   g0842(.A(new_n856_), .B(new_n855_), .Y(new_n892_));
  AOI21X1  g0843(.A0(new_n892_), .A1(new_n891_), .B0(new_n857_), .Y(new_n893_));
  NOR2X1   g0844(.A(new_n893_), .B(new_n843_), .Y(new_n894_));
  XOR2X1   g0845(.A(new_n893_), .B(new_n843_), .Y(new_n895_));
  XOR2X1   g0846(.A(new_n811_), .B(new_n808_), .Y(new_n896_));
  AOI21X1  g0847(.A0(new_n896_), .A1(new_n895_), .B0(new_n894_), .Y(new_n897_));
  XOR2X1   g0848(.A(new_n817_), .B(new_n816_), .Y(new_n898_));
  NOR2X1   g0849(.A(new_n898_), .B(new_n897_), .Y(new_n899_));
  XOR2X1   g0850(.A(new_n896_), .B(new_n895_), .Y(new_n900_));
  OR2X1    g0851(.A(new_n837_), .B(new_n828_), .Y(new_n901_));
  AOI22X1  g0852(.A0(new_n839_), .A1(new_n838_), .B0(new_n901_), .B1(new_n836_), .Y(new_n902_));
  NOR2X1   g0853(.A(new_n851_), .B(new_n850_), .Y(new_n903_));
  XOR2X1   g0854(.A(new_n853_), .B(new_n903_), .Y(new_n904_));
  OR2X1    g0855(.A(new_n904_), .B(new_n902_), .Y(new_n905_));
  INVX1    g0856(.A(new_n902_), .Y(new_n906_));
  XOR2X1   g0857(.A(new_n904_), .B(new_n906_), .Y(new_n907_));
  MX2X1    g0858(.A(new_n404_), .B(new_n407_), .S0(new_n749_), .Y(new_n908_));
  MX2X1    g0859(.A(new_n640_), .B(new_n639_), .S0(new_n229_), .Y(new_n909_));
  NOR2X1   g0860(.A(new_n401_), .B(new_n238_), .Y(new_n910_));
  OR4X1    g0861(.A(new_n248_), .B(new_n210_), .C(new_n198_), .D(new_n149_), .Y(new_n911_));
  NOR4X1   g0862(.A(new_n911_), .B(new_n396_), .C(new_n150_), .D(new_n136_), .Y(new_n912_));
  NOR3X1   g0863(.A(new_n363_), .B(new_n303_), .C(new_n123_), .Y(new_n913_));
  NOR4X1   g0864(.A(new_n573_), .B(new_n385_), .C(new_n321_), .D(new_n261_), .Y(new_n914_));
  NAND3X1  g0865(.A(new_n914_), .B(new_n913_), .C(new_n912_), .Y(new_n915_));
  OR4X1    g0866(.A(new_n126_), .B(new_n108_), .C(new_n83_), .D(new_n78_), .Y(new_n916_));
  NAND3X1  g0867(.A(new_n604_), .B(new_n355_), .C(new_n916_), .Y(new_n917_));
  OR4X1    g0868(.A(new_n213_), .B(new_n205_), .C(new_n168_), .D(new_n145_), .Y(new_n918_));
  OR4X1    g0869(.A(new_n918_), .B(new_n917_), .C(new_n370_), .D(new_n296_), .Y(new_n919_));
  NOR4X1   g0870(.A(new_n426_), .B(new_n437_), .C(new_n332_), .D(new_n255_), .Y(new_n920_));
  NOR4X1   g0871(.A(new_n220_), .B(new_n163_), .C(new_n147_), .D(new_n125_), .Y(new_n921_));
  NAND4X1  g0872(.A(new_n921_), .B(new_n920_), .C(new_n465_), .D(new_n278_), .Y(new_n922_));
  OR4X1    g0873(.A(new_n148_), .B(new_n90_), .C(new_n83_), .D(new_n101_), .Y(new_n923_));
  NAND3X1  g0874(.A(new_n301_), .B(new_n923_), .C(new_n468_), .Y(new_n924_));
  OR4X1    g0875(.A(new_n483_), .B(new_n314_), .C(new_n269_), .D(new_n131_), .Y(new_n925_));
  OR4X1    g0876(.A(new_n925_), .B(new_n924_), .C(new_n179_), .D(new_n162_), .Y(new_n926_));
  NOR4X1   g0877(.A(new_n926_), .B(new_n922_), .C(new_n919_), .D(new_n915_), .Y(new_n927_));
  AOI21X1  g0878(.A0(new_n927_), .A1(new_n525_), .B0(new_n715_), .Y(new_n928_));
  AND2X1   g0879(.A(new_n928_), .B(new_n910_), .Y(new_n929_));
  MX2X1    g0880(.A(new_n865_), .B(new_n863_), .S0(new_n591_), .Y(new_n930_));
  MX2X1    g0881(.A(new_n867_), .B(new_n868_), .S0(new_n602_), .Y(new_n931_));
  NOR2X1   g0882(.A(new_n931_), .B(new_n930_), .Y(new_n932_));
  XOR2X1   g0883(.A(new_n928_), .B(new_n910_), .Y(new_n933_));
  AOI21X1  g0884(.A0(new_n933_), .A1(new_n932_), .B0(new_n929_), .Y(new_n934_));
  NOR3X1   g0885(.A(new_n934_), .B(new_n909_), .C(new_n908_), .Y(new_n935_));
  NOR2X1   g0886(.A(new_n909_), .B(new_n908_), .Y(new_n936_));
  XOR2X1   g0887(.A(new_n934_), .B(new_n936_), .Y(new_n937_));
  MX2X1    g0888(.A(new_n586_), .B(new_n588_), .S0(new_n642_), .Y(new_n938_));
  MX2X1    g0889(.A(new_n595_), .B(new_n594_), .S0(new_n519_), .Y(new_n939_));
  MX2X1    g0890(.A(new_n795_), .B(new_n794_), .S0(new_n312_), .Y(new_n940_));
  MX2X1    g0891(.A(new_n797_), .B(new_n760_), .S0(new_n413_), .Y(new_n941_));
  OR2X1    g0892(.A(new_n941_), .B(new_n940_), .Y(new_n942_));
  NOR3X1   g0893(.A(new_n942_), .B(new_n939_), .C(new_n938_), .Y(new_n943_));
  MX2X1    g0894(.A(new_n630_), .B(new_n627_), .S0(new_n790_), .Y(new_n944_));
  MX2X1    g0895(.A(new_n634_), .B(new_n633_), .S0(new_n749_), .Y(new_n945_));
  NOR2X1   g0896(.A(new_n939_), .B(new_n938_), .Y(new_n946_));
  XOR2X1   g0897(.A(new_n942_), .B(new_n946_), .Y(new_n947_));
  NOR3X1   g0898(.A(new_n947_), .B(new_n945_), .C(new_n944_), .Y(new_n948_));
  NOR2X1   g0899(.A(new_n948_), .B(new_n943_), .Y(new_n949_));
  NOR2X1   g0900(.A(new_n949_), .B(new_n937_), .Y(new_n950_));
  NOR2X1   g0901(.A(new_n950_), .B(new_n935_), .Y(new_n951_));
  OAI21X1  g0902(.A0(new_n951_), .A1(new_n907_), .B0(new_n905_), .Y(new_n952_));
  XOR2X1   g0903(.A(new_n842_), .B(new_n840_), .Y(new_n953_));
  AND2X1   g0904(.A(new_n953_), .B(new_n952_), .Y(new_n954_));
  XOR2X1   g0905(.A(new_n953_), .B(new_n952_), .Y(new_n955_));
  XOR2X1   g0906(.A(new_n892_), .B(new_n891_), .Y(new_n956_));
  AND2X1   g0907(.A(new_n956_), .B(new_n955_), .Y(new_n957_));
  OAI21X1  g0908(.A0(new_n957_), .A1(new_n954_), .B0(new_n900_), .Y(new_n958_));
  AOI21X1  g0909(.A0(new_n956_), .A1(new_n955_), .B0(new_n954_), .Y(new_n959_));
  XOR2X1   g0910(.A(new_n959_), .B(new_n900_), .Y(new_n960_));
  OR4X1    g0911(.A(new_n926_), .B(new_n922_), .C(new_n919_), .D(new_n915_), .Y(new_n961_));
  NAND3X1  g0912(.A(new_n961_), .B(new_n829_), .C(new_n525_), .Y(new_n962_));
  NAND3X1  g0913(.A(new_n961_), .B(new_n715_), .C(new_n793_), .Y(new_n963_));
  INVX1    g0914(.A(new_n591_), .Y(new_n964_));
  OAI21X1  g0915(.A0(new_n715_), .A1(new_n964_), .B0(new_n927_), .Y(new_n965_));
  NAND3X1  g0916(.A(new_n965_), .B(new_n963_), .C(new_n962_), .Y(new_n966_));
  INVX1    g0917(.A(new_n238_), .Y(new_n967_));
  AOI21X1  g0918(.A0(new_n367_), .A1(new_n967_), .B0(new_n406_), .Y(new_n968_));
  AOI21X1  g0919(.A0(new_n404_), .A1(new_n967_), .B0(new_n968_), .Y(new_n969_));
  NAND2X1  g0920(.A(new_n969_), .B(new_n406_), .Y(new_n970_));
  MX2X1    g0921(.A(new_n407_), .B(new_n404_), .S0(new_n230_), .Y(new_n971_));
  MX2X1    g0922(.A(new_n640_), .B(new_n639_), .S0(new_n233_), .Y(new_n972_));
  NOR4X1   g0923(.A(new_n972_), .B(new_n971_), .C(new_n970_), .D(new_n966_), .Y(new_n973_));
  MX2X1    g0924(.A(new_n794_), .B(new_n795_), .S0(new_n413_), .Y(new_n974_));
  MX2X1    g0925(.A(new_n760_), .B(new_n797_), .S0(new_n642_), .Y(new_n975_));
  NOR2X1   g0926(.A(new_n975_), .B(new_n974_), .Y(new_n976_));
  INVX1    g0927(.A(new_n976_), .Y(new_n977_));
  MX2X1    g0928(.A(new_n586_), .B(new_n588_), .S0(new_n519_), .Y(new_n978_));
  MX2X1    g0929(.A(new_n594_), .B(new_n595_), .S0(new_n790_), .Y(new_n979_));
  OR2X1    g0930(.A(new_n979_), .B(new_n978_), .Y(new_n980_));
  MX2X1    g0931(.A(new_n627_), .B(new_n630_), .S0(new_n749_), .Y(new_n981_));
  MX2X1    g0932(.A(new_n634_), .B(new_n633_), .S0(new_n229_), .Y(new_n982_));
  NOR2X1   g0933(.A(new_n982_), .B(new_n981_), .Y(new_n983_));
  XOR2X1   g0934(.A(new_n983_), .B(new_n980_), .Y(new_n984_));
  OR4X1    g0935(.A(new_n982_), .B(new_n981_), .C(new_n979_), .D(new_n978_), .Y(new_n985_));
  OAI21X1  g0936(.A0(new_n984_), .A1(new_n977_), .B0(new_n985_), .Y(new_n986_));
  OAI22X1  g0937(.A0(new_n972_), .A1(new_n971_), .B0(new_n970_), .B1(new_n966_), .Y(new_n987_));
  AOI21X1  g0938(.A0(new_n987_), .A1(new_n986_), .B0(new_n973_), .Y(new_n988_));
  INVX1    g0939(.A(new_n988_), .Y(new_n989_));
  AOI22X1  g0940(.A0(new_n877_), .A1(new_n876_), .B0(new_n871_), .B1(new_n874_), .Y(new_n990_));
  XOR2X1   g0941(.A(new_n990_), .B(new_n989_), .Y(new_n991_));
  NOR2X1   g0942(.A(new_n886_), .B(new_n885_), .Y(new_n992_));
  XOR2X1   g0943(.A(new_n888_), .B(new_n992_), .Y(new_n993_));
  OR2X1    g0944(.A(new_n990_), .B(new_n988_), .Y(new_n994_));
  OAI21X1  g0945(.A0(new_n993_), .A1(new_n991_), .B0(new_n994_), .Y(new_n995_));
  XOR2X1   g0946(.A(new_n890_), .B(new_n878_), .Y(new_n996_));
  AND2X1   g0947(.A(new_n996_), .B(new_n995_), .Y(new_n997_));
  XOR2X1   g0948(.A(new_n951_), .B(new_n907_), .Y(new_n998_));
  XOR2X1   g0949(.A(new_n996_), .B(new_n995_), .Y(new_n999_));
  AND2X1   g0950(.A(new_n999_), .B(new_n998_), .Y(new_n1000_));
  OR2X1    g0951(.A(new_n1000_), .B(new_n997_), .Y(new_n1001_));
  XOR2X1   g0952(.A(new_n956_), .B(new_n955_), .Y(new_n1002_));
  AND2X1   g0953(.A(new_n1002_), .B(new_n1001_), .Y(new_n1003_));
  MX2X1    g0954(.A(new_n865_), .B(new_n863_), .S0(new_n602_), .Y(new_n1004_));
  MX2X1    g0955(.A(new_n868_), .B(new_n867_), .S0(new_n313_), .Y(new_n1005_));
  OR2X1    g0956(.A(new_n1005_), .B(new_n1004_), .Y(new_n1006_));
  MX2X1    g0957(.A(new_n404_), .B(new_n407_), .S0(new_n233_), .Y(new_n1007_));
  MX2X1    g0958(.A(new_n640_), .B(new_n639_), .S0(new_n238_), .Y(new_n1008_));
  NOR3X1   g0959(.A(new_n1008_), .B(new_n1007_), .C(new_n1006_), .Y(new_n1009_));
  OAI21X1  g0960(.A0(new_n1008_), .A1(new_n1007_), .B0(new_n1006_), .Y(new_n1010_));
  XOR2X1   g0961(.A(new_n970_), .B(new_n966_), .Y(new_n1011_));
  AOI21X1  g0962(.A0(new_n1011_), .A1(new_n1010_), .B0(new_n1009_), .Y(new_n1012_));
  INVX1    g0963(.A(new_n1012_), .Y(new_n1013_));
  XOR2X1   g0964(.A(new_n933_), .B(new_n932_), .Y(new_n1014_));
  NAND2X1  g0965(.A(new_n1014_), .B(new_n1013_), .Y(new_n1015_));
  XOR2X1   g0966(.A(new_n1014_), .B(new_n1012_), .Y(new_n1016_));
  NOR2X1   g0967(.A(new_n945_), .B(new_n944_), .Y(new_n1017_));
  XOR2X1   g0968(.A(new_n947_), .B(new_n1017_), .Y(new_n1018_));
  OAI21X1  g0969(.A0(new_n1018_), .A1(new_n1016_), .B0(new_n1015_), .Y(new_n1019_));
  XOR2X1   g0970(.A(new_n949_), .B(new_n937_), .Y(new_n1020_));
  AND2X1   g0971(.A(new_n1020_), .B(new_n1019_), .Y(new_n1021_));
  XOR2X1   g0972(.A(new_n1020_), .B(new_n1019_), .Y(new_n1022_));
  XOR2X1   g0973(.A(new_n993_), .B(new_n991_), .Y(new_n1023_));
  AOI21X1  g0974(.A0(new_n1023_), .A1(new_n1022_), .B0(new_n1021_), .Y(new_n1024_));
  INVX1    g0975(.A(new_n1024_), .Y(new_n1025_));
  XOR2X1   g0976(.A(new_n999_), .B(new_n998_), .Y(new_n1026_));
  NAND2X1  g0977(.A(new_n1026_), .B(new_n1025_), .Y(new_n1027_));
  NOR3X1   g0978(.A(new_n927_), .B(new_n715_), .C(new_n602_), .Y(new_n1028_));
  INVX1    g0979(.A(new_n602_), .Y(new_n1029_));
  NOR3X1   g0980(.A(new_n927_), .B(new_n829_), .C(new_n1029_), .Y(new_n1030_));
  AOI21X1  g0981(.A0(new_n829_), .A1(new_n312_), .B0(new_n961_), .Y(new_n1031_));
  NOR3X1   g0982(.A(new_n1031_), .B(new_n1030_), .C(new_n1028_), .Y(new_n1032_));
  AOI21X1  g0983(.A0(new_n628_), .A1(new_n584_), .B0(new_n350_), .Y(new_n1033_));
  OAI21X1  g0984(.A0(new_n629_), .A1(new_n967_), .B0(new_n1033_), .Y(new_n1034_));
  AOI21X1  g0985(.A0(new_n627_), .A1(new_n967_), .B0(new_n1034_), .Y(new_n1035_));
  NAND2X1  g0986(.A(new_n1035_), .B(new_n1032_), .Y(new_n1036_));
  MX2X1    g0987(.A(new_n795_), .B(new_n794_), .S0(new_n642_), .Y(new_n1037_));
  MX2X1    g0988(.A(new_n760_), .B(new_n797_), .S0(new_n519_), .Y(new_n1038_));
  NOR2X1   g0989(.A(new_n1038_), .B(new_n1037_), .Y(new_n1039_));
  INVX1    g0990(.A(new_n1039_), .Y(new_n1040_));
  MX2X1    g0991(.A(new_n588_), .B(new_n586_), .S0(new_n790_), .Y(new_n1041_));
  MX2X1    g0992(.A(new_n595_), .B(new_n594_), .S0(new_n749_), .Y(new_n1042_));
  NOR2X1   g0993(.A(new_n1042_), .B(new_n1041_), .Y(new_n1043_));
  XOR2X1   g0994(.A(new_n1043_), .B(new_n1040_), .Y(new_n1044_));
  OR4X1    g0995(.A(new_n1042_), .B(new_n1041_), .C(new_n1038_), .D(new_n1037_), .Y(new_n1045_));
  OAI21X1  g0996(.A0(new_n1044_), .A1(new_n1036_), .B0(new_n1045_), .Y(new_n1046_));
  MX2X1    g0997(.A(new_n630_), .B(new_n627_), .S0(new_n230_), .Y(new_n1047_));
  MX2X1    g0998(.A(new_n634_), .B(new_n633_), .S0(new_n233_), .Y(new_n1048_));
  NOR2X1   g0999(.A(new_n1048_), .B(new_n1047_), .Y(new_n1049_));
  NOR3X1   g1000(.A(new_n927_), .B(new_n715_), .C(new_n591_), .Y(new_n1050_));
  NOR3X1   g1001(.A(new_n927_), .B(new_n829_), .C(new_n964_), .Y(new_n1051_));
  AOI21X1  g1002(.A0(new_n829_), .A1(new_n602_), .B0(new_n961_), .Y(new_n1052_));
  NOR3X1   g1003(.A(new_n1052_), .B(new_n1051_), .C(new_n1050_), .Y(new_n1053_));
  MX2X1    g1004(.A(new_n865_), .B(new_n863_), .S0(new_n312_), .Y(new_n1054_));
  MX2X1    g1005(.A(new_n868_), .B(new_n867_), .S0(new_n413_), .Y(new_n1055_));
  NOR2X1   g1006(.A(new_n1055_), .B(new_n1054_), .Y(new_n1056_));
  XOR2X1   g1007(.A(new_n1056_), .B(new_n1053_), .Y(new_n1057_));
  AND2X1   g1008(.A(new_n1057_), .B(new_n1049_), .Y(new_n1058_));
  AND2X1   g1009(.A(new_n1056_), .B(new_n1053_), .Y(new_n1059_));
  OAI21X1  g1010(.A0(new_n1059_), .A1(new_n1058_), .B0(new_n1046_), .Y(new_n1060_));
  AOI21X1  g1011(.A0(new_n1057_), .A1(new_n1049_), .B0(new_n1059_), .Y(new_n1061_));
  XOR2X1   g1012(.A(new_n1061_), .B(new_n1046_), .Y(new_n1062_));
  XOR2X1   g1013(.A(new_n984_), .B(new_n976_), .Y(new_n1063_));
  OAI21X1  g1014(.A0(new_n1063_), .A1(new_n1062_), .B0(new_n1060_), .Y(new_n1064_));
  INVX1    g1015(.A(new_n973_), .Y(new_n1065_));
  AND2X1   g1016(.A(new_n987_), .B(new_n1065_), .Y(new_n1066_));
  XOR2X1   g1017(.A(new_n1066_), .B(new_n986_), .Y(new_n1067_));
  AND2X1   g1018(.A(new_n1067_), .B(new_n1064_), .Y(new_n1068_));
  XOR2X1   g1019(.A(new_n1018_), .B(new_n1016_), .Y(new_n1069_));
  XOR2X1   g1020(.A(new_n1067_), .B(new_n1064_), .Y(new_n1070_));
  AOI21X1  g1021(.A0(new_n1070_), .A1(new_n1069_), .B0(new_n1068_), .Y(new_n1071_));
  INVX1    g1022(.A(new_n1071_), .Y(new_n1072_));
  XOR2X1   g1023(.A(new_n1023_), .B(new_n1022_), .Y(new_n1073_));
  AND2X1   g1024(.A(new_n1073_), .B(new_n1072_), .Y(new_n1074_));
  MX2X1    g1025(.A(new_n795_), .B(new_n794_), .S0(new_n519_), .Y(new_n1075_));
  MX2X1    g1026(.A(new_n797_), .B(new_n760_), .S0(new_n790_), .Y(new_n1076_));
  OR2X1    g1027(.A(new_n1076_), .B(new_n1075_), .Y(new_n1077_));
  MX2X1    g1028(.A(new_n863_), .B(new_n865_), .S0(new_n413_), .Y(new_n1078_));
  MX2X1    g1029(.A(new_n867_), .B(new_n868_), .S0(new_n642_), .Y(new_n1079_));
  OR2X1    g1030(.A(new_n1079_), .B(new_n1078_), .Y(new_n1080_));
  MX2X1    g1031(.A(new_n586_), .B(new_n588_), .S0(new_n749_), .Y(new_n1081_));
  MX2X1    g1032(.A(new_n595_), .B(new_n594_), .S0(new_n229_), .Y(new_n1082_));
  NOR2X1   g1033(.A(new_n1082_), .B(new_n1081_), .Y(new_n1083_));
  XOR2X1   g1034(.A(new_n1083_), .B(new_n1080_), .Y(new_n1084_));
  OR4X1    g1035(.A(new_n1082_), .B(new_n1081_), .C(new_n1079_), .D(new_n1078_), .Y(new_n1085_));
  OAI21X1  g1036(.A0(new_n1084_), .A1(new_n1077_), .B0(new_n1085_), .Y(new_n1086_));
  XOR2X1   g1037(.A(new_n969_), .B(new_n406_), .Y(new_n1087_));
  AND2X1   g1038(.A(new_n1087_), .B(new_n1086_), .Y(new_n1088_));
  XOR2X1   g1039(.A(new_n1087_), .B(new_n1086_), .Y(new_n1089_));
  XOR2X1   g1040(.A(new_n1044_), .B(new_n1036_), .Y(new_n1090_));
  AOI21X1  g1041(.A0(new_n1090_), .A1(new_n1089_), .B0(new_n1088_), .Y(new_n1091_));
  INVX1    g1042(.A(new_n1009_), .Y(new_n1092_));
  NAND3X1  g1043(.A(new_n1011_), .B(new_n1010_), .C(new_n1092_), .Y(new_n1093_));
  AOI22X1  g1044(.A0(new_n1012_), .A1(new_n1010_), .B0(new_n1093_), .B1(new_n1011_), .Y(new_n1094_));
  INVX1    g1045(.A(new_n1094_), .Y(new_n1095_));
  XOR2X1   g1046(.A(new_n1095_), .B(new_n1091_), .Y(new_n1096_));
  INVX1    g1047(.A(new_n1063_), .Y(new_n1097_));
  XOR2X1   g1048(.A(new_n1097_), .B(new_n1062_), .Y(new_n1098_));
  OR2X1    g1049(.A(new_n1094_), .B(new_n1091_), .Y(new_n1099_));
  OAI21X1  g1050(.A0(new_n1098_), .A1(new_n1096_), .B0(new_n1099_), .Y(new_n1100_));
  XOR2X1   g1051(.A(new_n1070_), .B(new_n1069_), .Y(new_n1101_));
  AND2X1   g1052(.A(new_n1101_), .B(new_n1100_), .Y(new_n1102_));
  INVX1    g1053(.A(new_n1102_), .Y(new_n1103_));
  NOR3X1   g1054(.A(new_n927_), .B(new_n715_), .C(new_n312_), .Y(new_n1104_));
  NOR3X1   g1055(.A(new_n927_), .B(new_n829_), .C(new_n313_), .Y(new_n1105_));
  AOI21X1  g1056(.A0(new_n829_), .A1(new_n412_), .B0(new_n961_), .Y(new_n1106_));
  NOR3X1   g1057(.A(new_n1106_), .B(new_n1105_), .C(new_n1104_), .Y(new_n1107_));
  MX2X1    g1058(.A(new_n865_), .B(new_n863_), .S0(new_n642_), .Y(new_n1108_));
  MX2X1    g1059(.A(new_n867_), .B(new_n868_), .S0(new_n519_), .Y(new_n1109_));
  NOR2X1   g1060(.A(new_n1109_), .B(new_n1108_), .Y(new_n1110_));
  MX2X1    g1061(.A(new_n794_), .B(new_n795_), .S0(new_n790_), .Y(new_n1111_));
  MX2X1    g1062(.A(new_n760_), .B(new_n797_), .S0(new_n749_), .Y(new_n1112_));
  NOR2X1   g1063(.A(new_n1112_), .B(new_n1111_), .Y(new_n1113_));
  INVX1    g1064(.A(new_n1113_), .Y(new_n1114_));
  INVX1    g1065(.A(new_n1107_), .Y(new_n1115_));
  XOR2X1   g1066(.A(new_n1110_), .B(new_n1115_), .Y(new_n1116_));
  NOR2X1   g1067(.A(new_n1116_), .B(new_n1114_), .Y(new_n1117_));
  AOI21X1  g1068(.A0(new_n1110_), .A1(new_n1107_), .B0(new_n1117_), .Y(new_n1118_));
  MX2X1    g1069(.A(new_n627_), .B(new_n630_), .S0(new_n233_), .Y(new_n1119_));
  MX2X1    g1070(.A(new_n634_), .B(new_n633_), .S0(new_n238_), .Y(new_n1120_));
  NOR2X1   g1071(.A(new_n1120_), .B(new_n1119_), .Y(new_n1121_));
  XOR2X1   g1072(.A(new_n1035_), .B(new_n1032_), .Y(new_n1122_));
  INVX1    g1073(.A(new_n1122_), .Y(new_n1123_));
  XOR2X1   g1074(.A(new_n1123_), .B(new_n1121_), .Y(new_n1124_));
  NAND2X1  g1075(.A(new_n1122_), .B(new_n1121_), .Y(new_n1125_));
  OAI21X1  g1076(.A0(new_n1124_), .A1(new_n1118_), .B0(new_n1125_), .Y(new_n1126_));
  XOR2X1   g1077(.A(new_n1057_), .B(new_n1049_), .Y(new_n1127_));
  AND2X1   g1078(.A(new_n1127_), .B(new_n1126_), .Y(new_n1128_));
  XOR2X1   g1079(.A(new_n1090_), .B(new_n1089_), .Y(new_n1129_));
  XOR2X1   g1080(.A(new_n1127_), .B(new_n1126_), .Y(new_n1130_));
  AOI21X1  g1081(.A0(new_n1130_), .A1(new_n1129_), .B0(new_n1128_), .Y(new_n1131_));
  MX2X1    g1082(.A(new_n586_), .B(new_n588_), .S0(new_n233_), .Y(new_n1132_));
  MX2X1    g1083(.A(new_n595_), .B(new_n594_), .S0(new_n238_), .Y(new_n1133_));
  OR2X1    g1084(.A(new_n1133_), .B(new_n1132_), .Y(new_n1134_));
  MX2X1    g1085(.A(new_n865_), .B(new_n863_), .S0(new_n519_), .Y(new_n1135_));
  MX2X1    g1086(.A(new_n868_), .B(new_n867_), .S0(new_n790_), .Y(new_n1136_));
  OR2X1    g1087(.A(new_n1136_), .B(new_n1135_), .Y(new_n1137_));
  MX2X1    g1088(.A(new_n795_), .B(new_n794_), .S0(new_n749_), .Y(new_n1138_));
  MX2X1    g1089(.A(new_n797_), .B(new_n760_), .S0(new_n230_), .Y(new_n1139_));
  NOR2X1   g1090(.A(new_n1139_), .B(new_n1138_), .Y(new_n1140_));
  XOR2X1   g1091(.A(new_n1140_), .B(new_n1137_), .Y(new_n1141_));
  OR4X1    g1092(.A(new_n1139_), .B(new_n1138_), .C(new_n1136_), .D(new_n1135_), .Y(new_n1142_));
  OAI21X1  g1093(.A0(new_n1141_), .A1(new_n1134_), .B0(new_n1142_), .Y(new_n1143_));
  XOR2X1   g1094(.A(new_n1116_), .B(new_n1114_), .Y(new_n1144_));
  AND2X1   g1095(.A(new_n1144_), .B(new_n1143_), .Y(new_n1145_));
  MX2X1    g1096(.A(new_n588_), .B(new_n586_), .S0(new_n230_), .Y(new_n1146_));
  MX2X1    g1097(.A(new_n595_), .B(new_n594_), .S0(new_n233_), .Y(new_n1147_));
  NOR2X1   g1098(.A(new_n1147_), .B(new_n1146_), .Y(new_n1148_));
  NAND3X1  g1099(.A(new_n961_), .B(new_n829_), .C(new_n413_), .Y(new_n1149_));
  NAND3X1  g1100(.A(new_n961_), .B(new_n715_), .C(new_n412_), .Y(new_n1150_));
  OAI21X1  g1101(.A0(new_n715_), .A1(new_n641_), .B0(new_n927_), .Y(new_n1151_));
  NAND3X1  g1102(.A(new_n1151_), .B(new_n1150_), .C(new_n1149_), .Y(new_n1152_));
  AOI21X1  g1103(.A0(new_n592_), .A1(new_n967_), .B0(new_n593_), .Y(new_n1153_));
  AOI21X1  g1104(.A0(new_n586_), .A1(new_n967_), .B0(new_n1153_), .Y(new_n1154_));
  NAND2X1  g1105(.A(new_n1154_), .B(new_n593_), .Y(new_n1155_));
  NOR2X1   g1106(.A(new_n1155_), .B(new_n1152_), .Y(new_n1156_));
  XOR2X1   g1107(.A(new_n1156_), .B(new_n1148_), .Y(new_n1157_));
  NOR2X1   g1108(.A(new_n623_), .B(new_n238_), .Y(new_n1158_));
  XOR2X1   g1109(.A(new_n1158_), .B(new_n1157_), .Y(new_n1159_));
  XOR2X1   g1110(.A(new_n1144_), .B(new_n1143_), .Y(new_n1160_));
  AOI21X1  g1111(.A0(new_n1160_), .A1(new_n1159_), .B0(new_n1145_), .Y(new_n1161_));
  INVX1    g1112(.A(new_n1161_), .Y(new_n1162_));
  NOR3X1   g1113(.A(new_n927_), .B(new_n715_), .C(new_n519_), .Y(new_n1163_));
  INVX1    g1114(.A(new_n519_), .Y(new_n1164_));
  NOR3X1   g1115(.A(new_n927_), .B(new_n829_), .C(new_n1164_), .Y(new_n1165_));
  AOI21X1  g1116(.A0(new_n829_), .A1(new_n512_), .B0(new_n961_), .Y(new_n1166_));
  OR2X1    g1117(.A(new_n1166_), .B(new_n1165_), .Y(new_n1167_));
  NOR3X1   g1118(.A(new_n759_), .B(new_n761_), .C(new_n238_), .Y(new_n1168_));
  AOI21X1  g1119(.A0(new_n508_), .A1(new_n486_), .B0(new_n451_), .Y(new_n1169_));
  OAI21X1  g1120(.A0(new_n509_), .A1(new_n967_), .B0(new_n1169_), .Y(new_n1170_));
  OR4X1    g1121(.A(new_n1170_), .B(new_n1168_), .C(new_n1167_), .D(new_n1163_), .Y(new_n1171_));
  INVX1    g1122(.A(new_n1171_), .Y(new_n1172_));
  XOR2X1   g1123(.A(new_n1154_), .B(new_n593_), .Y(new_n1173_));
  NAND2X1  g1124(.A(new_n1173_), .B(new_n1172_), .Y(new_n1174_));
  MX2X1    g1125(.A(new_n865_), .B(new_n863_), .S0(new_n749_), .Y(new_n1175_));
  MX2X1    g1126(.A(new_n868_), .B(new_n867_), .S0(new_n230_), .Y(new_n1176_));
  MX2X1    g1127(.A(new_n795_), .B(new_n794_), .S0(new_n233_), .Y(new_n1177_));
  MX2X1    g1128(.A(new_n760_), .B(new_n797_), .S0(new_n238_), .Y(new_n1178_));
  NOR4X1   g1129(.A(new_n1178_), .B(new_n1177_), .C(new_n1176_), .D(new_n1175_), .Y(new_n1179_));
  OAI22X1  g1130(.A0(new_n1178_), .A1(new_n1177_), .B0(new_n1176_), .B1(new_n1175_), .Y(new_n1180_));
  NOR3X1   g1131(.A(new_n1166_), .B(new_n1165_), .C(new_n1163_), .Y(new_n1181_));
  NOR2X1   g1132(.A(new_n1170_), .B(new_n1168_), .Y(new_n1182_));
  XOR2X1   g1133(.A(new_n1182_), .B(new_n1181_), .Y(new_n1183_));
  AOI21X1  g1134(.A0(new_n1183_), .A1(new_n1180_), .B0(new_n1179_), .Y(new_n1184_));
  XOR2X1   g1135(.A(new_n1173_), .B(new_n1171_), .Y(new_n1185_));
  OAI21X1  g1136(.A0(new_n1185_), .A1(new_n1184_), .B0(new_n1174_), .Y(new_n1186_));
  INVX1    g1137(.A(new_n1186_), .Y(new_n1187_));
  NOR3X1   g1138(.A(new_n864_), .B(new_n830_), .C(new_n238_), .Y(new_n1188_));
  AOI21X1  g1139(.A0(new_n834_), .A1(new_n967_), .B0(new_n862_), .Y(new_n1189_));
  OAI21X1  g1140(.A0(new_n1189_), .A1(new_n1188_), .B0(new_n833_), .Y(new_n1190_));
  NAND3X1  g1141(.A(new_n831_), .B(new_n834_), .C(new_n967_), .Y(new_n1191_));
  OAI21X1  g1142(.A0(new_n830_), .A1(new_n238_), .B0(new_n833_), .Y(new_n1192_));
  NAND3X1  g1143(.A(new_n1192_), .B(new_n1191_), .C(new_n862_), .Y(new_n1193_));
  AOI21X1  g1144(.A0(new_n829_), .A1(new_n233_), .B0(new_n961_), .Y(new_n1194_));
  NOR3X1   g1145(.A(new_n927_), .B(new_n715_), .C(new_n229_), .Y(new_n1195_));
  NOR3X1   g1146(.A(new_n927_), .B(new_n829_), .C(new_n230_), .Y(new_n1196_));
  NOR3X1   g1147(.A(new_n1196_), .B(new_n1195_), .C(new_n1194_), .Y(new_n1197_));
  NOR2X1   g1148(.A(new_n927_), .B(new_n233_), .Y(new_n1198_));
  NOR3X1   g1149(.A(new_n1198_), .B(new_n715_), .C(new_n967_), .Y(new_n1199_));
  OR2X1    g1150(.A(new_n1199_), .B(new_n1197_), .Y(new_n1200_));
  NAND3X1  g1151(.A(new_n1200_), .B(new_n1193_), .C(new_n1190_), .Y(new_n1201_));
  NAND2X1  g1152(.A(new_n1199_), .B(new_n1197_), .Y(new_n1202_));
  INVX1    g1153(.A(new_n749_), .Y(new_n1203_));
  NAND3X1  g1154(.A(new_n961_), .B(new_n1203_), .C(new_n829_), .Y(new_n1204_));
  NAND3X1  g1155(.A(new_n961_), .B(new_n749_), .C(new_n715_), .Y(new_n1205_));
  OAI21X1  g1156(.A0(new_n715_), .A1(new_n230_), .B0(new_n927_), .Y(new_n1206_));
  AND2X1   g1157(.A(new_n1206_), .B(new_n1205_), .Y(new_n1207_));
  AND2X1   g1158(.A(new_n1207_), .B(new_n1204_), .Y(new_n1208_));
  XOR2X1   g1159(.A(new_n1208_), .B(new_n1193_), .Y(new_n1209_));
  NAND3X1  g1160(.A(new_n1209_), .B(new_n1202_), .C(new_n1201_), .Y(new_n1210_));
  MX2X1    g1161(.A(new_n865_), .B(new_n863_), .S0(new_n233_), .Y(new_n1211_));
  MX2X1    g1162(.A(new_n867_), .B(new_n868_), .S0(new_n238_), .Y(new_n1212_));
  NOR2X1   g1163(.A(new_n1212_), .B(new_n1211_), .Y(new_n1213_));
  AOI21X1  g1164(.A0(new_n1202_), .A1(new_n1201_), .B0(new_n1209_), .Y(new_n1214_));
  AOI21X1  g1165(.A0(new_n1213_), .A1(new_n1210_), .B0(new_n1214_), .Y(new_n1215_));
  NOR2X1   g1166(.A(new_n761_), .B(new_n238_), .Y(new_n1216_));
  INVX1    g1167(.A(new_n1216_), .Y(new_n1217_));
  NAND3X1  g1168(.A(new_n1206_), .B(new_n1205_), .C(new_n1204_), .Y(new_n1218_));
  NOR4X1   g1169(.A(new_n1218_), .B(new_n1189_), .C(new_n1188_), .D(new_n833_), .Y(new_n1219_));
  NAND3X1  g1170(.A(new_n961_), .B(new_n829_), .C(new_n790_), .Y(new_n1220_));
  NAND3X1  g1171(.A(new_n961_), .B(new_n715_), .C(new_n512_), .Y(new_n1221_));
  OAI21X1  g1172(.A0(new_n1203_), .A1(new_n715_), .B0(new_n927_), .Y(new_n1222_));
  NAND3X1  g1173(.A(new_n1222_), .B(new_n1221_), .C(new_n1220_), .Y(new_n1223_));
  MX2X1    g1174(.A(new_n865_), .B(new_n863_), .S0(new_n229_), .Y(new_n1224_));
  MX2X1    g1175(.A(new_n867_), .B(new_n868_), .S0(new_n233_), .Y(new_n1225_));
  NOR2X1   g1176(.A(new_n1225_), .B(new_n1224_), .Y(new_n1226_));
  XOR2X1   g1177(.A(new_n1226_), .B(new_n1223_), .Y(new_n1227_));
  XOR2X1   g1178(.A(new_n1227_), .B(new_n1219_), .Y(new_n1228_));
  AOI21X1  g1179(.A0(new_n1217_), .A1(new_n1215_), .B0(new_n1228_), .Y(new_n1229_));
  AOI21X1  g1180(.A0(new_n1192_), .A1(new_n1191_), .B0(new_n862_), .Y(new_n1230_));
  NOR3X1   g1181(.A(new_n1189_), .B(new_n1188_), .C(new_n833_), .Y(new_n1231_));
  NOR2X1   g1182(.A(new_n1199_), .B(new_n1197_), .Y(new_n1232_));
  NOR3X1   g1183(.A(new_n1232_), .B(new_n1231_), .C(new_n1230_), .Y(new_n1233_));
  AND2X1   g1184(.A(new_n1199_), .B(new_n1197_), .Y(new_n1234_));
  XOR2X1   g1185(.A(new_n1208_), .B(new_n1231_), .Y(new_n1235_));
  NOR3X1   g1186(.A(new_n1235_), .B(new_n1234_), .C(new_n1233_), .Y(new_n1236_));
  OR2X1    g1187(.A(new_n1212_), .B(new_n1211_), .Y(new_n1237_));
  OAI21X1  g1188(.A0(new_n1234_), .A1(new_n1233_), .B0(new_n1235_), .Y(new_n1238_));
  OAI21X1  g1189(.A0(new_n1237_), .A1(new_n1236_), .B0(new_n1238_), .Y(new_n1239_));
  AND2X1   g1190(.A(new_n1216_), .B(new_n1239_), .Y(new_n1240_));
  OR4X1    g1191(.A(new_n1178_), .B(new_n1177_), .C(new_n1176_), .D(new_n1175_), .Y(new_n1241_));
  NAND3X1  g1192(.A(new_n1183_), .B(new_n1180_), .C(new_n1241_), .Y(new_n1242_));
  AND2X1   g1193(.A(new_n1242_), .B(new_n1183_), .Y(new_n1243_));
  AND2X1   g1194(.A(new_n1184_), .B(new_n1180_), .Y(new_n1244_));
  OR2X1    g1195(.A(new_n1244_), .B(new_n1243_), .Y(new_n1245_));
  NOR3X1   g1196(.A(new_n1245_), .B(new_n1240_), .C(new_n1229_), .Y(new_n1246_));
  INVX1    g1197(.A(new_n1219_), .Y(new_n1247_));
  NAND4X1  g1198(.A(new_n1226_), .B(new_n1222_), .C(new_n1221_), .D(new_n1220_), .Y(new_n1248_));
  OAI21X1  g1199(.A0(new_n1227_), .A1(new_n1247_), .B0(new_n1248_), .Y(new_n1249_));
  INVX1    g1200(.A(new_n1249_), .Y(new_n1250_));
  OAI21X1  g1201(.A0(new_n1240_), .A1(new_n1229_), .B0(new_n1245_), .Y(new_n1251_));
  OAI21X1  g1202(.A0(new_n1250_), .A1(new_n1246_), .B0(new_n1251_), .Y(new_n1252_));
  XOR2X1   g1203(.A(new_n1185_), .B(new_n1184_), .Y(new_n1253_));
  MX2X1    g1204(.A(new_n795_), .B(new_n794_), .S0(new_n229_), .Y(new_n1254_));
  MX2X1    g1205(.A(new_n760_), .B(new_n797_), .S0(new_n233_), .Y(new_n1255_));
  NOR2X1   g1206(.A(new_n1255_), .B(new_n1254_), .Y(new_n1256_));
  MX2X1    g1207(.A(new_n863_), .B(new_n865_), .S0(new_n790_), .Y(new_n1257_));
  MX2X1    g1208(.A(new_n867_), .B(new_n868_), .S0(new_n749_), .Y(new_n1258_));
  NOR2X1   g1209(.A(new_n1258_), .B(new_n1257_), .Y(new_n1259_));
  NOR3X1   g1210(.A(new_n927_), .B(new_n715_), .C(new_n642_), .Y(new_n1260_));
  NOR3X1   g1211(.A(new_n927_), .B(new_n829_), .C(new_n641_), .Y(new_n1261_));
  AOI21X1  g1212(.A0(new_n829_), .A1(new_n519_), .B0(new_n961_), .Y(new_n1262_));
  NOR3X1   g1213(.A(new_n1262_), .B(new_n1261_), .C(new_n1260_), .Y(new_n1263_));
  XOR2X1   g1214(.A(new_n1263_), .B(new_n1259_), .Y(new_n1264_));
  XOR2X1   g1215(.A(new_n1264_), .B(new_n1256_), .Y(new_n1265_));
  OAI21X1  g1216(.A0(new_n1253_), .A1(new_n1252_), .B0(new_n1265_), .Y(new_n1266_));
  NAND2X1  g1217(.A(new_n1253_), .B(new_n1252_), .Y(new_n1267_));
  AOI21X1  g1218(.A0(new_n1267_), .A1(new_n1266_), .B0(new_n1187_), .Y(new_n1268_));
  NAND3X1  g1219(.A(new_n1267_), .B(new_n1266_), .C(new_n1187_), .Y(new_n1269_));
  XOR2X1   g1220(.A(new_n1141_), .B(new_n1134_), .Y(new_n1270_));
  AND2X1   g1221(.A(new_n1154_), .B(new_n593_), .Y(new_n1271_));
  XOR2X1   g1222(.A(new_n1271_), .B(new_n1152_), .Y(new_n1272_));
  AND2X1   g1223(.A(new_n1263_), .B(new_n1259_), .Y(new_n1273_));
  AOI21X1  g1224(.A0(new_n1264_), .A1(new_n1256_), .B0(new_n1273_), .Y(new_n1274_));
  XOR2X1   g1225(.A(new_n1274_), .B(new_n1272_), .Y(new_n1275_));
  XOR2X1   g1226(.A(new_n1275_), .B(new_n1270_), .Y(new_n1276_));
  AOI21X1  g1227(.A0(new_n1276_), .A1(new_n1269_), .B0(new_n1268_), .Y(new_n1277_));
  OR2X1    g1228(.A(new_n1274_), .B(new_n1272_), .Y(new_n1278_));
  AND2X1   g1229(.A(new_n1275_), .B(new_n1270_), .Y(new_n1279_));
  INVX1    g1230(.A(new_n1279_), .Y(new_n1280_));
  AND2X1   g1231(.A(new_n1280_), .B(new_n1278_), .Y(new_n1281_));
  NOR2X1   g1232(.A(new_n1281_), .B(new_n1277_), .Y(new_n1282_));
  XOR2X1   g1233(.A(new_n1160_), .B(new_n1159_), .Y(new_n1283_));
  INVX1    g1234(.A(new_n1283_), .Y(new_n1284_));
  AOI21X1  g1235(.A0(new_n1281_), .A1(new_n1277_), .B0(new_n1284_), .Y(new_n1285_));
  NOR3X1   g1236(.A(new_n1285_), .B(new_n1282_), .C(new_n1162_), .Y(new_n1286_));
  AND2X1   g1237(.A(new_n1158_), .B(new_n1157_), .Y(new_n1287_));
  NOR4X1   g1238(.A(new_n1155_), .B(new_n1152_), .C(new_n1147_), .D(new_n1146_), .Y(new_n1288_));
  OR2X1    g1239(.A(new_n1288_), .B(new_n1287_), .Y(new_n1289_));
  XOR2X1   g1240(.A(new_n1084_), .B(new_n1077_), .Y(new_n1290_));
  XOR2X1   g1241(.A(new_n1290_), .B(new_n1289_), .Y(new_n1291_));
  XOR2X1   g1242(.A(new_n1124_), .B(new_n1118_), .Y(new_n1292_));
  XOR2X1   g1243(.A(new_n1292_), .B(new_n1291_), .Y(new_n1293_));
  INVX1    g1244(.A(new_n1293_), .Y(new_n1294_));
  OAI21X1  g1245(.A0(new_n1285_), .A1(new_n1282_), .B0(new_n1162_), .Y(new_n1295_));
  OAI21X1  g1246(.A0(new_n1294_), .A1(new_n1286_), .B0(new_n1295_), .Y(new_n1296_));
  AND2X1   g1247(.A(new_n1292_), .B(new_n1291_), .Y(new_n1297_));
  AOI21X1  g1248(.A0(new_n1290_), .A1(new_n1289_), .B0(new_n1297_), .Y(new_n1298_));
  INVX1    g1249(.A(new_n1298_), .Y(new_n1299_));
  NAND2X1  g1250(.A(new_n1299_), .B(new_n1296_), .Y(new_n1300_));
  INVX1    g1251(.A(new_n1126_), .Y(new_n1301_));
  XOR2X1   g1252(.A(new_n1127_), .B(new_n1301_), .Y(new_n1302_));
  XOR2X1   g1253(.A(new_n1302_), .B(new_n1129_), .Y(new_n1303_));
  INVX1    g1254(.A(new_n1303_), .Y(new_n1304_));
  OAI21X1  g1255(.A0(new_n1299_), .A1(new_n1296_), .B0(new_n1304_), .Y(new_n1305_));
  NAND3X1  g1256(.A(new_n1305_), .B(new_n1300_), .C(new_n1131_), .Y(new_n1306_));
  XOR2X1   g1257(.A(new_n1098_), .B(new_n1096_), .Y(new_n1307_));
  AOI21X1  g1258(.A0(new_n1305_), .A1(new_n1300_), .B0(new_n1131_), .Y(new_n1308_));
  AOI21X1  g1259(.A0(new_n1307_), .A1(new_n1306_), .B0(new_n1308_), .Y(new_n1309_));
  XOR2X1   g1260(.A(new_n1101_), .B(new_n1100_), .Y(new_n1310_));
  INVX1    g1261(.A(new_n1310_), .Y(new_n1311_));
  OAI21X1  g1262(.A0(new_n1311_), .A1(new_n1309_), .B0(new_n1103_), .Y(new_n1312_));
  XOR2X1   g1263(.A(new_n1073_), .B(new_n1072_), .Y(new_n1313_));
  AOI21X1  g1264(.A0(new_n1313_), .A1(new_n1312_), .B0(new_n1074_), .Y(new_n1314_));
  XOR2X1   g1265(.A(new_n1026_), .B(new_n1025_), .Y(new_n1315_));
  INVX1    g1266(.A(new_n1315_), .Y(new_n1316_));
  OAI21X1  g1267(.A0(new_n1316_), .A1(new_n1314_), .B0(new_n1027_), .Y(new_n1317_));
  XOR2X1   g1268(.A(new_n1002_), .B(new_n1001_), .Y(new_n1318_));
  AOI21X1  g1269(.A0(new_n1318_), .A1(new_n1317_), .B0(new_n1003_), .Y(new_n1319_));
  OAI21X1  g1270(.A0(new_n1319_), .A1(new_n960_), .B0(new_n958_), .Y(new_n1320_));
  XOR2X1   g1271(.A(new_n898_), .B(new_n897_), .Y(new_n1321_));
  AOI21X1  g1272(.A0(new_n1321_), .A1(new_n1320_), .B0(new_n899_), .Y(new_n1322_));
  OAI21X1  g1273(.A0(new_n1322_), .A1(new_n822_), .B0(new_n820_), .Y(new_n1323_));
  XOR2X1   g1274(.A(new_n782_), .B(new_n781_), .Y(new_n1324_));
  AOI21X1  g1275(.A0(new_n1324_), .A1(new_n1323_), .B0(new_n783_), .Y(new_n1325_));
  OR2X1    g1276(.A(new_n1325_), .B(new_n693_), .Y(new_n1326_));
  OAI21X1  g1277(.A0(new_n691_), .A1(new_n676_), .B0(new_n1326_), .Y(new_n1327_));
  NOR2X1   g1278(.A(new_n679_), .B(new_n678_), .Y(new_n1328_));
  AOI21X1  g1279(.A0(new_n690_), .A1(new_n680_), .B0(new_n1328_), .Y(new_n1329_));
  INVX1    g1280(.A(new_n1329_), .Y(new_n1330_));
  MX2X1    g1281(.A(new_n407_), .B(new_n404_), .S0(new_n525_), .Y(new_n1331_));
  MX2X1    g1282(.A(new_n640_), .B(new_n639_), .S0(new_n591_), .Y(new_n1332_));
  OR2X1    g1283(.A(new_n1332_), .B(new_n1331_), .Y(new_n1333_));
  AND2X1   g1284(.A(new_n688_), .B(new_n686_), .Y(new_n1334_));
  AOI21X1  g1285(.A0(new_n689_), .A1(new_n684_), .B0(new_n1334_), .Y(new_n1335_));
  XOR2X1   g1286(.A(new_n1335_), .B(new_n1333_), .Y(new_n1336_));
  XOR2X1   g1287(.A(new_n686_), .B(new_n629_), .Y(new_n1337_));
  NOR2X1   g1288(.A(new_n602_), .B(new_n401_), .Y(new_n1338_));
  XOR2X1   g1289(.A(new_n1338_), .B(new_n1337_), .Y(new_n1339_));
  XOR2X1   g1290(.A(new_n1339_), .B(new_n1336_), .Y(new_n1340_));
  XOR2X1   g1291(.A(new_n1340_), .B(new_n1330_), .Y(new_n1341_));
  XOR2X1   g1292(.A(new_n1341_), .B(new_n1327_), .Y(new_n1342_));
  OR2X1    g1293(.A(new_n1342_), .B(new_n308_), .Y(new_n1343_));
  OR4X1    g1294(.A(new_n256_), .B(new_n203_), .C(new_n183_), .D(new_n174_), .Y(new_n1344_));
  OR4X1    g1295(.A(new_n1344_), .B(new_n337_), .C(new_n207_), .D(new_n141_), .Y(new_n1345_));
  OR4X1    g1296(.A(new_n283_), .B(new_n261_), .C(new_n220_), .D(new_n113_), .Y(new_n1346_));
  NOR4X1   g1297(.A(new_n1346_), .B(new_n1345_), .C(new_n609_), .D(new_n577_), .Y(new_n1347_));
  OR2X1    g1298(.A(new_n398_), .B(new_n208_), .Y(new_n1348_));
  OR2X1    g1299(.A(new_n1348_), .B(new_n317_), .Y(new_n1349_));
  OR4X1    g1300(.A(new_n262_), .B(new_n214_), .C(new_n125_), .D(new_n107_), .Y(new_n1350_));
  OR2X1    g1301(.A(new_n189_), .B(new_n121_), .Y(new_n1351_));
  OR2X1    g1302(.A(new_n1351_), .B(new_n348_), .Y(new_n1352_));
  OR4X1    g1303(.A(new_n616_), .B(new_n210_), .C(new_n198_), .D(new_n192_), .Y(new_n1353_));
  OR4X1    g1304(.A(new_n1353_), .B(new_n1352_), .C(new_n1350_), .D(new_n1349_), .Y(new_n1354_));
  OR4X1    g1305(.A(new_n580_), .B(new_n546_), .C(new_n273_), .D(new_n138_), .Y(new_n1355_));
  NOR2X1   g1306(.A(new_n1355_), .B(new_n1354_), .Y(new_n1356_));
  NOR3X1   g1307(.A(new_n388_), .B(new_n357_), .C(new_n347_), .Y(new_n1357_));
  INVX1    g1308(.A(new_n1357_), .Y(new_n1358_));
  OR2X1    g1309(.A(new_n322_), .B(new_n168_), .Y(new_n1359_));
  OR2X1    g1310(.A(new_n1359_), .B(new_n293_), .Y(new_n1360_));
  OR4X1    g1311(.A(new_n1360_), .B(new_n551_), .C(new_n294_), .D(new_n397_), .Y(new_n1361_));
  OR4X1    g1312(.A(new_n618_), .B(new_n315_), .C(new_n314_), .D(new_n181_), .Y(new_n1362_));
  NOR4X1   g1313(.A(new_n1362_), .B(new_n1361_), .C(new_n1358_), .D(new_n582_), .Y(new_n1363_));
  NAND3X1  g1314(.A(new_n1363_), .B(new_n1356_), .C(new_n1347_), .Y(new_n1364_));
  INVX1    g1315(.A(new_n1364_), .Y(new_n1365_));
  XOR2X1   g1316(.A(new_n1325_), .B(new_n693_), .Y(new_n1366_));
  NOR2X1   g1317(.A(new_n1366_), .B(new_n1365_), .Y(new_n1367_));
  OR2X1    g1318(.A(new_n185_), .B(new_n130_), .Y(new_n1368_));
  OR4X1    g1319(.A(new_n1368_), .B(new_n1355_), .C(new_n1354_), .D(new_n325_), .Y(new_n1369_));
  OR2X1    g1320(.A(new_n385_), .B(new_n163_), .Y(new_n1370_));
  OR4X1    g1321(.A(new_n251_), .B(new_n219_), .C(new_n195_), .D(new_n173_), .Y(new_n1371_));
  OR4X1    g1322(.A(new_n605_), .B(new_n341_), .C(new_n321_), .D(new_n305_), .Y(new_n1372_));
  OR4X1    g1323(.A(new_n1372_), .B(new_n1371_), .C(new_n1360_), .D(new_n1370_), .Y(new_n1373_));
  INVX1    g1324(.A(new_n255_), .Y(new_n1374_));
  NAND4X1  g1325(.A(new_n501_), .B(new_n354_), .C(new_n278_), .D(new_n1374_), .Y(new_n1375_));
  OR4X1    g1326(.A(new_n1375_), .B(new_n539_), .C(new_n196_), .D(new_n183_), .Y(new_n1376_));
  OR4X1    g1327(.A(new_n484_), .B(new_n260_), .C(new_n175_), .D(new_n165_), .Y(new_n1377_));
  NOR3X1   g1328(.A(new_n426_), .B(new_n337_), .C(new_n139_), .Y(new_n1378_));
  INVX1    g1329(.A(new_n1378_), .Y(new_n1379_));
  INVX1    g1330(.A(new_n913_), .Y(new_n1380_));
  OR4X1    g1331(.A(new_n1380_), .B(new_n388_), .C(new_n329_), .D(new_n247_), .Y(new_n1381_));
  OR4X1    g1332(.A(new_n1381_), .B(new_n1379_), .C(new_n1377_), .D(new_n1376_), .Y(new_n1382_));
  NOR3X1   g1333(.A(new_n1382_), .B(new_n1373_), .C(new_n1369_), .Y(new_n1383_));
  XOR2X1   g1334(.A(new_n1324_), .B(new_n1323_), .Y(new_n1384_));
  OR2X1    g1335(.A(new_n1384_), .B(new_n1383_), .Y(new_n1385_));
  OR2X1    g1336(.A(new_n527_), .B(new_n202_), .Y(new_n1386_));
  OR2X1    g1337(.A(new_n385_), .B(new_n332_), .Y(new_n1387_));
  NAND2X1  g1338(.A(new_n300_), .B(new_n278_), .Y(new_n1388_));
  OR2X1    g1339(.A(new_n346_), .B(new_n221_), .Y(new_n1389_));
  OR4X1    g1340(.A(new_n1389_), .B(new_n727_), .C(new_n618_), .D(new_n291_), .Y(new_n1390_));
  OR4X1    g1341(.A(new_n1390_), .B(new_n1388_), .C(new_n1387_), .D(new_n481_), .Y(new_n1391_));
  OR2X1    g1342(.A(new_n182_), .B(new_n145_), .Y(new_n1392_));
  NOR4X1   g1343(.A(new_n1392_), .B(new_n265_), .C(new_n132_), .D(new_n116_), .Y(new_n1393_));
  OR2X1    g1344(.A(new_n220_), .B(new_n113_), .Y(new_n1394_));
  OR4X1    g1345(.A(new_n304_), .B(new_n188_), .C(new_n136_), .D(new_n131_), .Y(new_n1395_));
  NOR4X1   g1346(.A(new_n1395_), .B(new_n1394_), .C(new_n169_), .D(new_n162_), .Y(new_n1396_));
  NOR4X1   g1347(.A(new_n398_), .B(new_n347_), .C(new_n292_), .D(new_n259_), .Y(new_n1397_));
  NOR4X1   g1348(.A(new_n488_), .B(new_n280_), .C(new_n159_), .D(new_n121_), .Y(new_n1398_));
  NAND4X1  g1349(.A(new_n1398_), .B(new_n1397_), .C(new_n1396_), .D(new_n1393_), .Y(new_n1399_));
  NOR4X1   g1350(.A(new_n1399_), .B(new_n1391_), .C(new_n1386_), .D(new_n463_), .Y(new_n1400_));
  XOR2X1   g1351(.A(new_n1322_), .B(new_n822_), .Y(new_n1401_));
  NOR2X1   g1352(.A(new_n1401_), .B(new_n1400_), .Y(new_n1402_));
  NOR4X1   g1353(.A(new_n446_), .B(new_n356_), .C(new_n283_), .D(new_n149_), .Y(new_n1403_));
  INVX1    g1354(.A(new_n1403_), .Y(new_n1404_));
  OR4X1    g1355(.A(new_n188_), .B(new_n182_), .C(new_n180_), .D(new_n159_), .Y(new_n1405_));
  OR4X1    g1356(.A(new_n1405_), .B(new_n603_), .C(new_n467_), .D(new_n389_), .Y(new_n1406_));
  INVX1    g1357(.A(new_n470_), .Y(new_n1407_));
  OR4X1    g1358(.A(new_n527_), .B(new_n265_), .C(new_n204_), .D(new_n170_), .Y(new_n1408_));
  NOR4X1   g1359(.A(new_n1408_), .B(new_n1407_), .C(new_n461_), .D(new_n425_), .Y(new_n1409_));
  INVX1    g1360(.A(new_n1409_), .Y(new_n1410_));
  NOR3X1   g1361(.A(new_n252_), .B(new_n202_), .C(new_n141_), .Y(new_n1411_));
  NOR4X1   g1362(.A(new_n706_), .B(new_n253_), .C(new_n185_), .D(new_n132_), .Y(new_n1412_));
  NAND2X1  g1363(.A(new_n1412_), .B(new_n1411_), .Y(new_n1413_));
  OR4X1    g1364(.A(new_n1413_), .B(new_n1410_), .C(new_n1406_), .D(new_n1404_), .Y(new_n1414_));
  NOR4X1   g1365(.A(new_n1414_), .B(new_n494_), .C(new_n491_), .D(new_n263_), .Y(new_n1415_));
  XOR2X1   g1366(.A(new_n1321_), .B(new_n1320_), .Y(new_n1416_));
  OR2X1    g1367(.A(new_n1416_), .B(new_n1415_), .Y(new_n1417_));
  OR4X1    g1368(.A(new_n346_), .B(new_n330_), .C(new_n321_), .D(new_n221_), .Y(new_n1418_));
  OR4X1    g1369(.A(new_n198_), .B(new_n182_), .C(new_n163_), .D(new_n91_), .Y(new_n1419_));
  OR2X1    g1370(.A(new_n1419_), .B(new_n296_), .Y(new_n1420_));
  NOR4X1   g1371(.A(new_n1420_), .B(new_n1418_), .C(new_n736_), .D(new_n580_), .Y(new_n1421_));
  NOR3X1   g1372(.A(new_n303_), .B(new_n180_), .C(new_n179_), .Y(new_n1422_));
  NAND2X1  g1373(.A(new_n1422_), .B(new_n1421_), .Y(new_n1423_));
  NOR3X1   g1374(.A(new_n488_), .B(new_n294_), .C(new_n208_), .Y(new_n1424_));
  OR4X1    g1375(.A(new_n317_), .B(new_n264_), .C(new_n252_), .D(new_n249_), .Y(new_n1425_));
  OR2X1    g1376(.A(new_n159_), .B(new_n139_), .Y(new_n1426_));
  NOR4X1   g1377(.A(new_n1426_), .B(new_n1425_), .C(new_n173_), .D(new_n155_), .Y(new_n1427_));
  NAND4X1  g1378(.A(new_n1427_), .B(new_n1424_), .C(new_n458_), .D(new_n457_), .Y(new_n1428_));
  OR4X1    g1379(.A(new_n388_), .B(new_n271_), .C(new_n261_), .D(new_n255_), .Y(new_n1429_));
  NOR4X1   g1380(.A(new_n1429_), .B(new_n291_), .C(new_n137_), .D(new_n97_), .Y(new_n1430_));
  NOR4X1   g1381(.A(new_n332_), .B(new_n262_), .C(new_n248_), .D(new_n125_), .Y(new_n1431_));
  OR4X1    g1382(.A(new_n337_), .B(new_n175_), .C(new_n157_), .D(new_n336_), .Y(new_n1432_));
  NOR2X1   g1383(.A(new_n1432_), .B(new_n420_), .Y(new_n1433_));
  NAND3X1  g1384(.A(new_n1433_), .B(new_n1431_), .C(new_n1430_), .Y(new_n1434_));
  NOR3X1   g1385(.A(new_n1434_), .B(new_n1428_), .C(new_n1423_), .Y(new_n1435_));
  XOR2X1   g1386(.A(new_n1319_), .B(new_n960_), .Y(new_n1436_));
  NOR2X1   g1387(.A(new_n1436_), .B(new_n1435_), .Y(new_n1437_));
  AND2X1   g1388(.A(new_n923_), .B(new_n338_), .Y(new_n1438_));
  NOR4X1   g1389(.A(new_n527_), .B(new_n329_), .C(new_n204_), .D(new_n91_), .Y(new_n1439_));
  NAND2X1  g1390(.A(new_n1439_), .B(new_n1438_), .Y(new_n1440_));
  OR4X1    g1391(.A(new_n1440_), .B(new_n1358_), .C(new_n565_), .D(new_n374_), .Y(new_n1441_));
  INVX1    g1392(.A(new_n489_), .Y(new_n1442_));
  OR4X1    g1393(.A(new_n325_), .B(new_n211_), .C(new_n136_), .D(new_n116_), .Y(new_n1443_));
  OR4X1    g1394(.A(new_n1443_), .B(new_n551_), .C(new_n314_), .D(new_n294_), .Y(new_n1444_));
  OR2X1    g1395(.A(new_n1444_), .B(new_n1442_), .Y(new_n1445_));
  OR4X1    g1396(.A(new_n321_), .B(new_n292_), .C(new_n205_), .D(new_n97_), .Y(new_n1446_));
  OR4X1    g1397(.A(new_n1446_), .B(new_n382_), .C(new_n317_), .D(new_n167_), .Y(new_n1447_));
  OR4X1    g1398(.A(new_n574_), .B(new_n246_), .C(new_n121_), .D(new_n110_), .Y(new_n1448_));
  OR2X1    g1399(.A(new_n1448_), .B(new_n1447_), .Y(new_n1449_));
  NOR4X1   g1400(.A(new_n1449_), .B(new_n1445_), .C(new_n1441_), .D(new_n436_), .Y(new_n1450_));
  XOR2X1   g1401(.A(new_n1318_), .B(new_n1317_), .Y(new_n1451_));
  OR2X1    g1402(.A(new_n1451_), .B(new_n1450_), .Y(new_n1452_));
  NOR4X1   g1403(.A(new_n305_), .B(new_n281_), .C(new_n248_), .D(new_n91_), .Y(new_n1453_));
  NAND3X1  g1404(.A(new_n1453_), .B(new_n1378_), .C(new_n487_), .Y(new_n1454_));
  NAND2X1  g1405(.A(new_n604_), .B(new_n1374_), .Y(new_n1455_));
  OR4X1    g1406(.A(new_n1455_), .B(new_n315_), .C(new_n251_), .D(new_n203_), .Y(new_n1456_));
  OR2X1    g1407(.A(new_n488_), .B(new_n325_), .Y(new_n1457_));
  OR4X1    g1408(.A(new_n1457_), .B(new_n322_), .C(new_n296_), .D(new_n265_), .Y(new_n1458_));
  OR4X1    g1409(.A(new_n1458_), .B(new_n1456_), .C(new_n1454_), .D(new_n1404_), .Y(new_n1459_));
  OR2X1    g1410(.A(new_n372_), .B(new_n107_), .Y(new_n1460_));
  OR2X1    g1411(.A(new_n430_), .B(new_n358_), .Y(new_n1461_));
  OR4X1    g1412(.A(new_n1461_), .B(new_n1460_), .C(new_n385_), .D(new_n163_), .Y(new_n1462_));
  OR4X1    g1413(.A(new_n483_), .B(new_n220_), .C(new_n150_), .D(new_n141_), .Y(new_n1463_));
  OR4X1    g1414(.A(new_n1463_), .B(new_n398_), .C(new_n329_), .D(new_n210_), .Y(new_n1464_));
  OR4X1    g1415(.A(new_n1464_), .B(new_n1462_), .C(new_n1447_), .D(new_n263_), .Y(new_n1465_));
  NOR4X1   g1416(.A(new_n1465_), .B(new_n1459_), .C(new_n454_), .D(new_n201_), .Y(new_n1466_));
  XOR2X1   g1417(.A(new_n1316_), .B(new_n1314_), .Y(new_n1467_));
  NOR2X1   g1418(.A(new_n1467_), .B(new_n1466_), .Y(new_n1468_));
  INVX1    g1419(.A(new_n702_), .Y(new_n1469_));
  OR2X1    g1420(.A(new_n197_), .B(new_n165_), .Y(new_n1470_));
  NOR4X1   g1421(.A(new_n1470_), .B(new_n616_), .C(new_n330_), .D(new_n271_), .Y(new_n1471_));
  INVX1    g1422(.A(new_n1471_), .Y(new_n1472_));
  OR4X1    g1423(.A(new_n332_), .B(new_n294_), .C(new_n185_), .D(new_n113_), .Y(new_n1473_));
  OR2X1    g1424(.A(new_n247_), .B(new_n179_), .Y(new_n1474_));
  OR4X1    g1425(.A(new_n1474_), .B(new_n426_), .C(new_n305_), .D(new_n279_), .Y(new_n1475_));
  NOR4X1   g1426(.A(new_n1475_), .B(new_n1473_), .C(new_n1472_), .D(new_n1469_), .Y(new_n1476_));
  OR4X1    g1427(.A(new_n488_), .B(new_n325_), .C(new_n270_), .D(new_n209_), .Y(new_n1477_));
  OR4X1    g1428(.A(new_n385_), .B(new_n347_), .C(new_n304_), .D(new_n97_), .Y(new_n1478_));
  OR4X1    g1429(.A(new_n220_), .B(new_n213_), .C(new_n189_), .D(new_n158_), .Y(new_n1479_));
  NOR4X1   g1430(.A(new_n1479_), .B(new_n1478_), .C(new_n1477_), .D(new_n553_), .Y(new_n1480_));
  NAND3X1  g1431(.A(new_n1480_), .B(new_n1476_), .C(new_n1409_), .Y(new_n1481_));
  INVX1    g1432(.A(new_n1131_), .Y(new_n1482_));
  AND2X1   g1433(.A(new_n1299_), .B(new_n1296_), .Y(new_n1483_));
  OR2X1    g1434(.A(new_n1281_), .B(new_n1277_), .Y(new_n1484_));
  XOR2X1   g1435(.A(new_n1227_), .B(new_n1247_), .Y(new_n1485_));
  OAI21X1  g1436(.A0(new_n1216_), .A1(new_n1239_), .B0(new_n1485_), .Y(new_n1486_));
  OR2X1    g1437(.A(new_n1217_), .B(new_n1215_), .Y(new_n1487_));
  AOI22X1  g1438(.A0(new_n1184_), .A1(new_n1180_), .B0(new_n1242_), .B1(new_n1183_), .Y(new_n1488_));
  NAND3X1  g1439(.A(new_n1488_), .B(new_n1487_), .C(new_n1486_), .Y(new_n1489_));
  AOI21X1  g1440(.A0(new_n1487_), .A1(new_n1486_), .B0(new_n1488_), .Y(new_n1490_));
  AOI21X1  g1441(.A0(new_n1249_), .A1(new_n1489_), .B0(new_n1490_), .Y(new_n1491_));
  XOR2X1   g1442(.A(new_n1173_), .B(new_n1172_), .Y(new_n1492_));
  XOR2X1   g1443(.A(new_n1492_), .B(new_n1184_), .Y(new_n1493_));
  INVX1    g1444(.A(new_n1265_), .Y(new_n1494_));
  AOI21X1  g1445(.A0(new_n1493_), .A1(new_n1491_), .B0(new_n1494_), .Y(new_n1495_));
  AND2X1   g1446(.A(new_n1253_), .B(new_n1252_), .Y(new_n1496_));
  OAI21X1  g1447(.A0(new_n1496_), .A1(new_n1495_), .B0(new_n1186_), .Y(new_n1497_));
  NOR3X1   g1448(.A(new_n1496_), .B(new_n1495_), .C(new_n1186_), .Y(new_n1498_));
  INVX1    g1449(.A(new_n1276_), .Y(new_n1499_));
  OAI21X1  g1450(.A0(new_n1499_), .A1(new_n1498_), .B0(new_n1497_), .Y(new_n1500_));
  NAND2X1  g1451(.A(new_n1280_), .B(new_n1278_), .Y(new_n1501_));
  OAI21X1  g1452(.A0(new_n1501_), .A1(new_n1500_), .B0(new_n1283_), .Y(new_n1502_));
  NAND3X1  g1453(.A(new_n1502_), .B(new_n1484_), .C(new_n1161_), .Y(new_n1503_));
  AOI21X1  g1454(.A0(new_n1502_), .A1(new_n1484_), .B0(new_n1161_), .Y(new_n1504_));
  AOI21X1  g1455(.A0(new_n1293_), .A1(new_n1503_), .B0(new_n1504_), .Y(new_n1505_));
  AOI21X1  g1456(.A0(new_n1298_), .A1(new_n1505_), .B0(new_n1303_), .Y(new_n1506_));
  NOR3X1   g1457(.A(new_n1506_), .B(new_n1483_), .C(new_n1482_), .Y(new_n1507_));
  INVX1    g1458(.A(new_n1307_), .Y(new_n1508_));
  OAI21X1  g1459(.A0(new_n1506_), .A1(new_n1483_), .B0(new_n1482_), .Y(new_n1509_));
  OAI21X1  g1460(.A0(new_n1508_), .A1(new_n1507_), .B0(new_n1509_), .Y(new_n1510_));
  AOI21X1  g1461(.A0(new_n1310_), .A1(new_n1510_), .B0(new_n1102_), .Y(new_n1511_));
  XOR2X1   g1462(.A(new_n1313_), .B(new_n1511_), .Y(new_n1512_));
  NAND2X1  g1463(.A(new_n1512_), .B(new_n1481_), .Y(new_n1513_));
  NOR2X1   g1464(.A(new_n1512_), .B(new_n1481_), .Y(new_n1514_));
  XOR2X1   g1465(.A(new_n1310_), .B(new_n1510_), .Y(new_n1515_));
  OR2X1    g1466(.A(new_n213_), .B(new_n150_), .Y(new_n1516_));
  INVX1    g1467(.A(new_n254_), .Y(new_n1517_));
  OR4X1    g1468(.A(new_n1353_), .B(new_n1442_), .C(new_n320_), .D(new_n1517_), .Y(new_n1518_));
  OR2X1    g1469(.A(new_n280_), .B(new_n269_), .Y(new_n1519_));
  OR2X1    g1470(.A(new_n1519_), .B(new_n272_), .Y(new_n1520_));
  OR4X1    g1471(.A(new_n420_), .B(new_n294_), .C(new_n179_), .D(new_n141_), .Y(new_n1521_));
  OR4X1    g1472(.A(new_n1521_), .B(new_n1520_), .C(new_n1518_), .D(new_n1516_), .Y(new_n1522_));
  INVX1    g1473(.A(new_n250_), .Y(new_n1523_));
  OR4X1    g1474(.A(new_n437_), .B(new_n284_), .C(new_n207_), .D(new_n107_), .Y(new_n1524_));
  OR4X1    g1475(.A(new_n202_), .B(new_n158_), .C(new_n336_), .D(new_n130_), .Y(new_n1525_));
  OR4X1    g1476(.A(new_n1525_), .B(new_n605_), .C(new_n281_), .D(new_n261_), .Y(new_n1526_));
  OR4X1    g1477(.A(new_n1526_), .B(new_n1524_), .C(new_n456_), .D(new_n1523_), .Y(new_n1527_));
  NOR3X1   g1478(.A(new_n1527_), .B(new_n1522_), .C(new_n1441_), .Y(new_n1528_));
  AND2X1   g1479(.A(new_n1528_), .B(new_n1515_), .Y(new_n1529_));
  OAI21X1  g1480(.A0(new_n1529_), .A1(new_n1514_), .B0(new_n1513_), .Y(new_n1530_));
  NAND2X1  g1481(.A(new_n1467_), .B(new_n1466_), .Y(new_n1531_));
  AOI21X1  g1482(.A0(new_n1531_), .A1(new_n1530_), .B0(new_n1468_), .Y(new_n1532_));
  AND2X1   g1483(.A(new_n1451_), .B(new_n1450_), .Y(new_n1533_));
  OAI21X1  g1484(.A0(new_n1533_), .A1(new_n1532_), .B0(new_n1452_), .Y(new_n1534_));
  XOR2X1   g1485(.A(new_n1436_), .B(new_n1435_), .Y(new_n1535_));
  AOI21X1  g1486(.A0(new_n1535_), .A1(new_n1534_), .B0(new_n1437_), .Y(new_n1536_));
  AND2X1   g1487(.A(new_n1416_), .B(new_n1415_), .Y(new_n1537_));
  OAI21X1  g1488(.A0(new_n1537_), .A1(new_n1536_), .B0(new_n1417_), .Y(new_n1538_));
  XOR2X1   g1489(.A(new_n1401_), .B(new_n1400_), .Y(new_n1539_));
  AOI21X1  g1490(.A0(new_n1539_), .A1(new_n1538_), .B0(new_n1402_), .Y(new_n1540_));
  AND2X1   g1491(.A(new_n1384_), .B(new_n1383_), .Y(new_n1541_));
  OAI21X1  g1492(.A0(new_n1541_), .A1(new_n1540_), .B0(new_n1385_), .Y(new_n1542_));
  XOR2X1   g1493(.A(new_n1366_), .B(new_n1365_), .Y(new_n1543_));
  AOI21X1  g1494(.A0(new_n1543_), .A1(new_n1542_), .B0(new_n1367_), .Y(new_n1544_));
  AND2X1   g1495(.A(new_n1342_), .B(new_n308_), .Y(new_n1545_));
  OAI21X1  g1496(.A0(new_n1545_), .A1(new_n1544_), .B0(new_n1343_), .Y(new_n1546_));
  OR2X1    g1497(.A(new_n449_), .B(new_n448_), .Y(new_n1547_));
  OR4X1    g1498(.A(new_n551_), .B(new_n264_), .C(new_n216_), .D(new_n193_), .Y(new_n1548_));
  OR4X1    g1499(.A(new_n1548_), .B(new_n186_), .C(new_n167_), .D(new_n130_), .Y(new_n1549_));
  OR4X1    g1500(.A(new_n398_), .B(new_n358_), .C(new_n321_), .D(new_n116_), .Y(new_n1550_));
  OR4X1    g1501(.A(new_n1550_), .B(new_n1549_), .C(new_n1352_), .D(new_n1547_), .Y(new_n1551_));
  OR2X1    g1502(.A(new_n317_), .B(new_n314_), .Y(new_n1552_));
  OR4X1    g1503(.A(new_n1552_), .B(new_n527_), .C(new_n281_), .D(new_n207_), .Y(new_n1553_));
  INVX1    g1504(.A(new_n283_), .Y(new_n1554_));
  NAND3X1  g1505(.A(new_n465_), .B(new_n1554_), .C(new_n492_), .Y(new_n1555_));
  OR4X1    g1506(.A(new_n214_), .B(new_n175_), .C(new_n336_), .D(new_n134_), .Y(new_n1556_));
  NOR4X1   g1507(.A(new_n1556_), .B(new_n1555_), .C(new_n1553_), .D(new_n419_), .Y(new_n1557_));
  INVX1    g1508(.A(new_n1557_), .Y(new_n1558_));
  NOR4X1   g1509(.A(new_n1558_), .B(new_n1551_), .C(new_n1522_), .D(new_n1376_), .Y(new_n1559_));
  NOR2X1   g1510(.A(new_n1335_), .B(new_n1333_), .Y(new_n1560_));
  AOI21X1  g1511(.A0(new_n1339_), .A1(new_n1336_), .B0(new_n1560_), .Y(new_n1561_));
  NOR2X1   g1512(.A(new_n686_), .B(new_n629_), .Y(new_n1562_));
  AOI21X1  g1513(.A0(new_n1338_), .A1(new_n1337_), .B0(new_n1562_), .Y(new_n1563_));
  NOR3X1   g1514(.A(new_n793_), .B(new_n403_), .C(new_n367_), .Y(new_n1564_));
  OAI22X1  g1515(.A0(new_n793_), .A1(new_n367_), .B0(new_n405_), .B1(new_n401_), .Y(new_n1565_));
  INVX1    g1516(.A(new_n1565_), .Y(new_n1566_));
  NOR2X1   g1517(.A(new_n591_), .B(new_n401_), .Y(new_n1567_));
  NOR3X1   g1518(.A(new_n1567_), .B(new_n1566_), .C(new_n1564_), .Y(new_n1568_));
  NOR2X1   g1519(.A(new_n1566_), .B(new_n1564_), .Y(new_n1569_));
  NOR3X1   g1520(.A(new_n1569_), .B(new_n591_), .C(new_n401_), .Y(new_n1570_));
  NOR3X1   g1521(.A(new_n1570_), .B(new_n1568_), .C(new_n1563_), .Y(new_n1571_));
  INVX1    g1522(.A(new_n1570_), .Y(new_n1572_));
  INVX1    g1523(.A(new_n1563_), .Y(new_n1573_));
  AOI21X1  g1524(.A0(new_n1572_), .A1(new_n1573_), .B0(new_n1568_), .Y(new_n1574_));
  NAND2X1  g1525(.A(new_n1574_), .B(new_n1572_), .Y(new_n1575_));
  OAI21X1  g1526(.A0(new_n1571_), .A1(new_n1563_), .B0(new_n1575_), .Y(new_n1576_));
  XOR2X1   g1527(.A(new_n1576_), .B(new_n1561_), .Y(new_n1577_));
  INVX1    g1528(.A(new_n1577_), .Y(new_n1578_));
  NAND2X1  g1529(.A(new_n1340_), .B(new_n1330_), .Y(new_n1579_));
  NAND2X1  g1530(.A(new_n1341_), .B(new_n1327_), .Y(new_n1580_));
  NAND2X1  g1531(.A(new_n1580_), .B(new_n1579_), .Y(new_n1581_));
  XOR2X1   g1532(.A(new_n1581_), .B(new_n1578_), .Y(new_n1582_));
  XOR2X1   g1533(.A(new_n1582_), .B(new_n1559_), .Y(new_n1583_));
  XOR2X1   g1534(.A(new_n1583_), .B(new_n1546_), .Y(new_n1584_));
  INVX1    g1535(.A(new_n1584_), .Y(new_n1585_));
  NOR2X1   g1536(.A(new_n1582_), .B(new_n1559_), .Y(new_n1586_));
  AOI21X1  g1537(.A0(new_n1583_), .A1(new_n1546_), .B0(new_n1586_), .Y(new_n1587_));
  OR4X1    g1538(.A(new_n213_), .B(new_n211_), .C(new_n210_), .D(new_n189_), .Y(new_n1588_));
  OR4X1    g1539(.A(new_n446_), .B(new_n332_), .C(new_n252_), .D(new_n184_), .Y(new_n1589_));
  OR4X1    g1540(.A(new_n1589_), .B(new_n603_), .C(new_n483_), .D(new_n220_), .Y(new_n1590_));
  OR4X1    g1541(.A(new_n1349_), .B(new_n527_), .C(new_n264_), .D(new_n169_), .Y(new_n1591_));
  OR4X1    g1542(.A(new_n120_), .B(new_n108_), .C(new_n92_), .D(new_n101_), .Y(new_n1592_));
  NOR3X1   g1543(.A(new_n385_), .B(new_n551_), .C(new_n251_), .Y(new_n1593_));
  NAND3X1  g1544(.A(new_n1593_), .B(new_n1592_), .C(new_n392_), .Y(new_n1594_));
  OR4X1    g1545(.A(new_n1594_), .B(new_n1591_), .C(new_n1590_), .D(new_n1588_), .Y(new_n1595_));
  NOR4X1   g1546(.A(new_n1595_), .B(new_n1423_), .C(new_n711_), .D(new_n454_), .Y(new_n1596_));
  XOR2X1   g1547(.A(new_n591_), .B(new_n525_), .Y(new_n1597_));
  AOI21X1  g1548(.A0(new_n1597_), .A1(new_n405_), .B0(new_n401_), .Y(new_n1598_));
  OAI21X1  g1549(.A0(new_n1597_), .A1(new_n405_), .B0(new_n1598_), .Y(new_n1599_));
  OAI21X1  g1550(.A0(new_n1570_), .A1(new_n1568_), .B0(new_n1573_), .Y(new_n1600_));
  AOI21X1  g1551(.A0(new_n1575_), .A1(new_n1600_), .B0(new_n1561_), .Y(new_n1601_));
  AOI21X1  g1552(.A0(new_n1581_), .A1(new_n1578_), .B0(new_n1601_), .Y(new_n1602_));
  XOR2X1   g1553(.A(new_n1602_), .B(new_n1574_), .Y(new_n1603_));
  XOR2X1   g1554(.A(new_n1603_), .B(new_n1599_), .Y(new_n1604_));
  XOR2X1   g1555(.A(new_n1604_), .B(new_n1596_), .Y(new_n1605_));
  OR2X1    g1556(.A(new_n1605_), .B(new_n1587_), .Y(new_n1606_));
  OR2X1    g1557(.A(new_n1604_), .B(new_n1596_), .Y(new_n1607_));
  NAND2X1  g1558(.A(new_n1604_), .B(new_n1596_), .Y(new_n1608_));
  NAND3X1  g1559(.A(new_n1608_), .B(new_n1607_), .C(new_n1587_), .Y(new_n1609_));
  AOI21X1  g1560(.A0(new_n1609_), .A1(new_n1606_), .B0(new_n1585_), .Y(new_n1610_));
  XOR2X1   g1561(.A(new_n1342_), .B(new_n308_), .Y(new_n1611_));
  OR2X1    g1562(.A(new_n1611_), .B(new_n1544_), .Y(new_n1612_));
  OAI21X1  g1563(.A0(new_n1546_), .A1(new_n1545_), .B0(new_n1612_), .Y(new_n1613_));
  NAND2X1  g1564(.A(new_n1613_), .B(new_n1584_), .Y(new_n1614_));
  XOR2X1   g1565(.A(new_n1543_), .B(new_n1542_), .Y(new_n1615_));
  AND2X1   g1566(.A(new_n1615_), .B(new_n1613_), .Y(new_n1616_));
  XOR2X1   g1567(.A(new_n1384_), .B(new_n1383_), .Y(new_n1617_));
  OAI22X1  g1568(.A0(new_n1542_), .A1(new_n1541_), .B0(new_n1617_), .B1(new_n1540_), .Y(new_n1618_));
  NAND2X1  g1569(.A(new_n1618_), .B(new_n1615_), .Y(new_n1619_));
  XOR2X1   g1570(.A(new_n1539_), .B(new_n1538_), .Y(new_n1620_));
  AND2X1   g1571(.A(new_n1620_), .B(new_n1618_), .Y(new_n1621_));
  XOR2X1   g1572(.A(new_n1416_), .B(new_n1415_), .Y(new_n1622_));
  OAI22X1  g1573(.A0(new_n1538_), .A1(new_n1537_), .B0(new_n1622_), .B1(new_n1536_), .Y(new_n1623_));
  NAND2X1  g1574(.A(new_n1623_), .B(new_n1620_), .Y(new_n1624_));
  OR2X1    g1575(.A(new_n1622_), .B(new_n1536_), .Y(new_n1625_));
  NAND2X1  g1576(.A(new_n1416_), .B(new_n1415_), .Y(new_n1626_));
  NAND3X1  g1577(.A(new_n1626_), .B(new_n1536_), .C(new_n1417_), .Y(new_n1627_));
  NOR2X1   g1578(.A(new_n1451_), .B(new_n1450_), .Y(new_n1628_));
  OR2X1    g1579(.A(new_n1467_), .B(new_n1466_), .Y(new_n1629_));
  AND2X1   g1580(.A(new_n1512_), .B(new_n1481_), .Y(new_n1630_));
  OR2X1    g1581(.A(new_n1512_), .B(new_n1481_), .Y(new_n1631_));
  NAND2X1  g1582(.A(new_n1528_), .B(new_n1515_), .Y(new_n1632_));
  AOI21X1  g1583(.A0(new_n1632_), .A1(new_n1631_), .B0(new_n1630_), .Y(new_n1633_));
  AND2X1   g1584(.A(new_n1467_), .B(new_n1466_), .Y(new_n1634_));
  OAI21X1  g1585(.A0(new_n1634_), .A1(new_n1633_), .B0(new_n1629_), .Y(new_n1635_));
  XOR2X1   g1586(.A(new_n1451_), .B(new_n1450_), .Y(new_n1636_));
  AOI21X1  g1587(.A0(new_n1636_), .A1(new_n1635_), .B0(new_n1628_), .Y(new_n1637_));
  XOR2X1   g1588(.A(new_n1535_), .B(new_n1637_), .Y(new_n1638_));
  AOI21X1  g1589(.A0(new_n1627_), .A1(new_n1625_), .B0(new_n1638_), .Y(new_n1639_));
  XOR2X1   g1590(.A(new_n1636_), .B(new_n1532_), .Y(new_n1640_));
  OR2X1    g1591(.A(new_n1640_), .B(new_n1638_), .Y(new_n1641_));
  XOR2X1   g1592(.A(new_n1636_), .B(new_n1635_), .Y(new_n1642_));
  XOR2X1   g1593(.A(new_n1467_), .B(new_n1466_), .Y(new_n1643_));
  OAI22X1  g1594(.A0(new_n1635_), .A1(new_n1634_), .B0(new_n1643_), .B1(new_n1633_), .Y(new_n1644_));
  AND2X1   g1595(.A(new_n1644_), .B(new_n1642_), .Y(new_n1645_));
  NOR2X1   g1596(.A(new_n1643_), .B(new_n1633_), .Y(new_n1646_));
  AOI21X1  g1597(.A0(new_n1532_), .A1(new_n1531_), .B0(new_n1646_), .Y(new_n1647_));
  OAI21X1  g1598(.A0(new_n1514_), .A1(new_n1630_), .B0(new_n1632_), .Y(new_n1648_));
  NAND3X1  g1599(.A(new_n1529_), .B(new_n1631_), .C(new_n1513_), .Y(new_n1649_));
  AND2X1   g1600(.A(new_n1649_), .B(new_n1648_), .Y(new_n1650_));
  XOR2X1   g1601(.A(new_n1528_), .B(new_n1515_), .Y(new_n1651_));
  AOI21X1  g1602(.A0(new_n1651_), .A1(new_n1647_), .B0(new_n1650_), .Y(new_n1652_));
  OR2X1    g1603(.A(new_n1644_), .B(new_n1642_), .Y(new_n1653_));
  AOI21X1  g1604(.A0(new_n1653_), .A1(new_n1652_), .B0(new_n1645_), .Y(new_n1654_));
  AND2X1   g1605(.A(new_n1640_), .B(new_n1638_), .Y(new_n1655_));
  OAI21X1  g1606(.A0(new_n1655_), .A1(new_n1654_), .B0(new_n1641_), .Y(new_n1656_));
  INVX1    g1607(.A(new_n1638_), .Y(new_n1657_));
  XOR2X1   g1608(.A(new_n1657_), .B(new_n1623_), .Y(new_n1658_));
  AOI21X1  g1609(.A0(new_n1658_), .A1(new_n1656_), .B0(new_n1639_), .Y(new_n1659_));
  XOR2X1   g1610(.A(new_n1623_), .B(new_n1620_), .Y(new_n1660_));
  INVX1    g1611(.A(new_n1660_), .Y(new_n1661_));
  OAI21X1  g1612(.A0(new_n1661_), .A1(new_n1659_), .B0(new_n1624_), .Y(new_n1662_));
  XOR2X1   g1613(.A(new_n1620_), .B(new_n1618_), .Y(new_n1663_));
  AOI21X1  g1614(.A0(new_n1663_), .A1(new_n1662_), .B0(new_n1621_), .Y(new_n1664_));
  XOR2X1   g1615(.A(new_n1618_), .B(new_n1615_), .Y(new_n1665_));
  INVX1    g1616(.A(new_n1665_), .Y(new_n1666_));
  OAI21X1  g1617(.A0(new_n1666_), .A1(new_n1664_), .B0(new_n1619_), .Y(new_n1667_));
  XOR2X1   g1618(.A(new_n1615_), .B(new_n1613_), .Y(new_n1668_));
  AOI21X1  g1619(.A0(new_n1668_), .A1(new_n1667_), .B0(new_n1616_), .Y(new_n1669_));
  XOR2X1   g1620(.A(new_n1613_), .B(new_n1584_), .Y(new_n1670_));
  INVX1    g1621(.A(new_n1670_), .Y(new_n1671_));
  OAI21X1  g1622(.A0(new_n1671_), .A1(new_n1669_), .B0(new_n1614_), .Y(new_n1672_));
  AND2X1   g1623(.A(new_n1609_), .B(new_n1606_), .Y(new_n1673_));
  XOR2X1   g1624(.A(new_n1673_), .B(new_n1585_), .Y(new_n1674_));
  AOI21X1  g1625(.A0(new_n1674_), .A1(new_n1672_), .B0(new_n1610_), .Y(new_n1675_));
  NAND2X1  g1626(.A(new_n1609_), .B(new_n1606_), .Y(new_n1676_));
  AND2X1   g1627(.A(new_n1604_), .B(new_n1596_), .Y(new_n1677_));
  OAI21X1  g1628(.A0(new_n1677_), .A1(new_n1587_), .B0(new_n1607_), .Y(new_n1678_));
  NOR3X1   g1629(.A(new_n611_), .B(new_n538_), .C(new_n209_), .Y(new_n1679_));
  NOR4X1   g1630(.A(new_n316_), .B(new_n262_), .C(new_n246_), .D(new_n336_), .Y(new_n1680_));
  NOR4X1   g1631(.A(new_n426_), .B(new_n372_), .C(new_n294_), .D(new_n91_), .Y(new_n1681_));
  NAND4X1  g1632(.A(new_n1681_), .B(new_n1680_), .C(new_n1679_), .D(new_n254_), .Y(new_n1682_));
  OR2X1    g1633(.A(new_n346_), .B(new_n113_), .Y(new_n1683_));
  OR4X1    g1634(.A(new_n1683_), .B(new_n259_), .C(new_n173_), .D(new_n163_), .Y(new_n1684_));
  OR2X1    g1635(.A(new_n1684_), .B(new_n541_), .Y(new_n1685_));
  NOR4X1   g1636(.A(new_n1685_), .B(new_n1682_), .C(new_n1410_), .D(new_n915_), .Y(new_n1686_));
  INVX1    g1637(.A(new_n1686_), .Y(new_n1687_));
  XOR2X1   g1638(.A(new_n1687_), .B(new_n1678_), .Y(new_n1688_));
  XOR2X1   g1639(.A(new_n1688_), .B(new_n1676_), .Y(new_n1689_));
  XOR2X1   g1640(.A(new_n1689_), .B(new_n1675_), .Y(new_n1690_));
  INVX1    g1641(.A(new_n244_), .Y(new_n1691_));
  XOR2X1   g1642(.A(new_n967_), .B(new_n233_), .Y(new_n1692_));
  NOR2X1   g1643(.A(new_n1692_), .B(new_n1691_), .Y(new_n1693_));
  INVX1    g1644(.A(new_n1693_), .Y(new_n1694_));
  XOR2X1   g1645(.A(new_n1686_), .B(new_n1678_), .Y(new_n1695_));
  AND2X1   g1646(.A(new_n1691_), .B(new_n234_), .Y(new_n1696_));
  INVX1    g1647(.A(new_n1692_), .Y(new_n1697_));
  OR2X1    g1648(.A(new_n1691_), .B(new_n234_), .Y(new_n1698_));
  NOR2X1   g1649(.A(new_n1698_), .B(new_n1697_), .Y(new_n1699_));
  AOI22X1  g1650(.A0(new_n1699_), .A1(new_n1584_), .B0(new_n1696_), .B1(new_n1695_), .Y(new_n1700_));
  OAI21X1  g1651(.A0(new_n1694_), .A1(new_n1673_), .B0(new_n1700_), .Y(new_n1701_));
  AOI21X1  g1652(.A0(new_n1690_), .A1(new_n245_), .B0(new_n1701_), .Y(new_n1702_));
  XOR2X1   g1653(.A(new_n1702_), .B(new_n230_), .Y(new_n1703_));
  XOR2X1   g1654(.A(new_n602_), .B(new_n313_), .Y(new_n1704_));
  OAI21X1  g1655(.A0(new_n1704_), .A1(new_n1651_), .B0(new_n525_), .Y(new_n1705_));
  XOR2X1   g1656(.A(new_n1651_), .B(new_n1650_), .Y(new_n1706_));
  NOR2X1   g1657(.A(new_n1704_), .B(new_n1597_), .Y(new_n1707_));
  XOR2X1   g1658(.A(new_n602_), .B(new_n964_), .Y(new_n1708_));
  INVX1    g1659(.A(new_n1708_), .Y(new_n1709_));
  AND2X1   g1660(.A(new_n1709_), .B(new_n1704_), .Y(new_n1710_));
  INVX1    g1661(.A(new_n1710_), .Y(new_n1711_));
  INVX1    g1662(.A(new_n1597_), .Y(new_n1712_));
  NOR2X1   g1663(.A(new_n1704_), .B(new_n1712_), .Y(new_n1713_));
  INVX1    g1664(.A(new_n1713_), .Y(new_n1714_));
  OAI22X1  g1665(.A0(new_n1714_), .A1(new_n1650_), .B0(new_n1711_), .B1(new_n1651_), .Y(new_n1715_));
  AOI21X1  g1666(.A0(new_n1707_), .A1(new_n1706_), .B0(new_n1715_), .Y(new_n1716_));
  XOR2X1   g1667(.A(new_n1716_), .B(new_n525_), .Y(new_n1717_));
  XOR2X1   g1668(.A(new_n1717_), .B(new_n1705_), .Y(new_n1718_));
  XOR2X1   g1669(.A(new_n641_), .B(new_n519_), .Y(new_n1719_));
  XOR2X1   g1670(.A(new_n413_), .B(new_n312_), .Y(new_n1720_));
  NOR2X1   g1671(.A(new_n1720_), .B(new_n1719_), .Y(new_n1721_));
  INVX1    g1672(.A(new_n1721_), .Y(new_n1722_));
  INVX1    g1673(.A(new_n1719_), .Y(new_n1723_));
  AND2X1   g1674(.A(new_n1720_), .B(new_n1723_), .Y(new_n1724_));
  XOR2X1   g1675(.A(new_n641_), .B(new_n412_), .Y(new_n1725_));
  INVX1    g1676(.A(new_n1725_), .Y(new_n1726_));
  NOR3X1   g1677(.A(new_n1726_), .B(new_n1720_), .C(new_n1723_), .Y(new_n1727_));
  INVX1    g1678(.A(new_n1727_), .Y(new_n1728_));
  NOR2X1   g1679(.A(new_n1725_), .B(new_n1723_), .Y(new_n1729_));
  INVX1    g1680(.A(new_n1729_), .Y(new_n1730_));
  OAI22X1  g1681(.A0(new_n1730_), .A1(new_n1640_), .B0(new_n1728_), .B1(new_n1647_), .Y(new_n1731_));
  AOI21X1  g1682(.A0(new_n1724_), .A1(new_n1657_), .B0(new_n1731_), .Y(new_n1732_));
  NAND2X1  g1683(.A(new_n1644_), .B(new_n1642_), .Y(new_n1733_));
  NAND2X1  g1684(.A(new_n1649_), .B(new_n1648_), .Y(new_n1734_));
  INVX1    g1685(.A(new_n1651_), .Y(new_n1735_));
  OAI21X1  g1686(.A0(new_n1735_), .A1(new_n1644_), .B0(new_n1734_), .Y(new_n1736_));
  NOR2X1   g1687(.A(new_n1644_), .B(new_n1642_), .Y(new_n1737_));
  OAI21X1  g1688(.A0(new_n1737_), .A1(new_n1736_), .B0(new_n1733_), .Y(new_n1738_));
  XOR2X1   g1689(.A(new_n1642_), .B(new_n1638_), .Y(new_n1739_));
  AND2X1   g1690(.A(new_n1739_), .B(new_n1738_), .Y(new_n1740_));
  NOR2X1   g1691(.A(new_n1640_), .B(new_n1638_), .Y(new_n1741_));
  NOR3X1   g1692(.A(new_n1655_), .B(new_n1738_), .C(new_n1741_), .Y(new_n1742_));
  NOR2X1   g1693(.A(new_n1742_), .B(new_n1740_), .Y(new_n1743_));
  OAI21X1  g1694(.A0(new_n1743_), .A1(new_n1722_), .B0(new_n1732_), .Y(new_n1744_));
  XOR2X1   g1695(.A(new_n1744_), .B(new_n313_), .Y(new_n1745_));
  NAND2X1  g1696(.A(new_n1745_), .B(new_n1718_), .Y(new_n1746_));
  NOR2X1   g1697(.A(new_n1704_), .B(new_n1651_), .Y(new_n1747_));
  NOR2X1   g1698(.A(new_n1719_), .B(new_n1651_), .Y(new_n1748_));
  NOR2X1   g1699(.A(new_n1748_), .B(new_n312_), .Y(new_n1749_));
  INVX1    g1700(.A(new_n1724_), .Y(new_n1750_));
  OAI22X1  g1701(.A0(new_n1730_), .A1(new_n1651_), .B0(new_n1750_), .B1(new_n1650_), .Y(new_n1751_));
  AOI21X1  g1702(.A0(new_n1721_), .A1(new_n1706_), .B0(new_n1751_), .Y(new_n1752_));
  XOR2X1   g1703(.A(new_n1752_), .B(new_n312_), .Y(new_n1753_));
  AND2X1   g1704(.A(new_n1753_), .B(new_n1749_), .Y(new_n1754_));
  OAI22X1  g1705(.A0(new_n1730_), .A1(new_n1650_), .B0(new_n1728_), .B1(new_n1651_), .Y(new_n1755_));
  AOI21X1  g1706(.A0(new_n1724_), .A1(new_n1644_), .B0(new_n1755_), .Y(new_n1756_));
  NAND2X1  g1707(.A(new_n1651_), .B(new_n1734_), .Y(new_n1757_));
  XOR2X1   g1708(.A(new_n1757_), .B(new_n1644_), .Y(new_n1758_));
  OAI21X1  g1709(.A0(new_n1758_), .A1(new_n1722_), .B0(new_n1756_), .Y(new_n1759_));
  XOR2X1   g1710(.A(new_n1759_), .B(new_n313_), .Y(new_n1760_));
  NAND3X1  g1711(.A(new_n1760_), .B(new_n1754_), .C(new_n1747_), .Y(new_n1761_));
  NAND2X1  g1712(.A(new_n1760_), .B(new_n1754_), .Y(new_n1762_));
  XOR2X1   g1713(.A(new_n1762_), .B(new_n1747_), .Y(new_n1763_));
  XOR2X1   g1714(.A(new_n1644_), .B(new_n1642_), .Y(new_n1764_));
  NOR2X1   g1715(.A(new_n1764_), .B(new_n1736_), .Y(new_n1765_));
  NOR3X1   g1716(.A(new_n1737_), .B(new_n1652_), .C(new_n1645_), .Y(new_n1766_));
  OR2X1    g1717(.A(new_n1766_), .B(new_n1765_), .Y(new_n1767_));
  AOI22X1  g1718(.A0(new_n1729_), .A1(new_n1644_), .B0(new_n1727_), .B1(new_n1734_), .Y(new_n1768_));
  OAI21X1  g1719(.A0(new_n1750_), .A1(new_n1640_), .B0(new_n1768_), .Y(new_n1769_));
  AOI21X1  g1720(.A0(new_n1767_), .A1(new_n1721_), .B0(new_n1769_), .Y(new_n1770_));
  XOR2X1   g1721(.A(new_n1770_), .B(new_n312_), .Y(new_n1771_));
  INVX1    g1722(.A(new_n1771_), .Y(new_n1772_));
  OAI21X1  g1723(.A0(new_n1772_), .A1(new_n1763_), .B0(new_n1761_), .Y(new_n1773_));
  XOR2X1   g1724(.A(new_n1745_), .B(new_n1718_), .Y(new_n1774_));
  NAND2X1  g1725(.A(new_n1774_), .B(new_n1773_), .Y(new_n1775_));
  NAND2X1  g1726(.A(new_n1775_), .B(new_n1746_), .Y(new_n1776_));
  XOR2X1   g1727(.A(new_n1658_), .B(new_n1656_), .Y(new_n1777_));
  AND2X1   g1728(.A(new_n1627_), .B(new_n1625_), .Y(new_n1778_));
  AOI22X1  g1729(.A0(new_n1729_), .A1(new_n1657_), .B0(new_n1727_), .B1(new_n1642_), .Y(new_n1779_));
  OAI21X1  g1730(.A0(new_n1750_), .A1(new_n1778_), .B0(new_n1779_), .Y(new_n1780_));
  AOI21X1  g1731(.A0(new_n1777_), .A1(new_n1721_), .B0(new_n1780_), .Y(new_n1781_));
  XOR2X1   g1732(.A(new_n1781_), .B(new_n312_), .Y(new_n1782_));
  NOR2X1   g1733(.A(new_n1717_), .B(new_n1705_), .Y(new_n1783_));
  INVX1    g1734(.A(new_n1707_), .Y(new_n1784_));
  NAND3X1  g1735(.A(new_n1708_), .B(new_n1704_), .C(new_n1712_), .Y(new_n1785_));
  OAI22X1  g1736(.A0(new_n1785_), .A1(new_n1651_), .B0(new_n1711_), .B1(new_n1650_), .Y(new_n1786_));
  AOI21X1  g1737(.A0(new_n1713_), .A1(new_n1644_), .B0(new_n1786_), .Y(new_n1787_));
  OAI21X1  g1738(.A0(new_n1758_), .A1(new_n1784_), .B0(new_n1787_), .Y(new_n1788_));
  XOR2X1   g1739(.A(new_n1788_), .B(new_n525_), .Y(new_n1789_));
  XOR2X1   g1740(.A(new_n1789_), .B(new_n1783_), .Y(new_n1790_));
  XOR2X1   g1741(.A(new_n1790_), .B(new_n1782_), .Y(new_n1791_));
  XOR2X1   g1742(.A(new_n1791_), .B(new_n1776_), .Y(new_n1792_));
  XOR2X1   g1743(.A(new_n749_), .B(new_n230_), .Y(new_n1793_));
  XOR2X1   g1744(.A(new_n749_), .B(new_n790_), .Y(new_n1794_));
  INVX1    g1745(.A(new_n1794_), .Y(new_n1795_));
  AND2X1   g1746(.A(new_n1795_), .B(new_n1793_), .Y(new_n1796_));
  INVX1    g1747(.A(new_n1615_), .Y(new_n1797_));
  INVX1    g1748(.A(new_n1620_), .Y(new_n1798_));
  INVX1    g1749(.A(new_n1793_), .Y(new_n1799_));
  XOR2X1   g1750(.A(new_n519_), .B(new_n790_), .Y(new_n1800_));
  AND2X1   g1751(.A(new_n1800_), .B(new_n1799_), .Y(new_n1801_));
  INVX1    g1752(.A(new_n1801_), .Y(new_n1802_));
  NAND2X1  g1753(.A(new_n1794_), .B(new_n1793_), .Y(new_n1803_));
  NOR2X1   g1754(.A(new_n1803_), .B(new_n1800_), .Y(new_n1804_));
  INVX1    g1755(.A(new_n1804_), .Y(new_n1805_));
  OAI22X1  g1756(.A0(new_n1805_), .A1(new_n1798_), .B0(new_n1802_), .B1(new_n1797_), .Y(new_n1806_));
  AOI21X1  g1757(.A0(new_n1796_), .A1(new_n1618_), .B0(new_n1806_), .Y(new_n1807_));
  XOR2X1   g1758(.A(new_n1665_), .B(new_n1664_), .Y(new_n1808_));
  NOR2X1   g1759(.A(new_n1800_), .B(new_n1793_), .Y(new_n1809_));
  INVX1    g1760(.A(new_n1809_), .Y(new_n1810_));
  OAI21X1  g1761(.A0(new_n1810_), .A1(new_n1808_), .B0(new_n1807_), .Y(new_n1811_));
  XOR2X1   g1762(.A(new_n1811_), .B(new_n1164_), .Y(new_n1812_));
  NAND2X1  g1763(.A(new_n1812_), .B(new_n1792_), .Y(new_n1813_));
  XOR2X1   g1764(.A(new_n1663_), .B(new_n1662_), .Y(new_n1814_));
  INVX1    g1765(.A(new_n1618_), .Y(new_n1815_));
  AOI22X1  g1766(.A0(new_n1804_), .A1(new_n1623_), .B0(new_n1796_), .B1(new_n1620_), .Y(new_n1816_));
  OAI21X1  g1767(.A0(new_n1802_), .A1(new_n1815_), .B0(new_n1816_), .Y(new_n1817_));
  AOI21X1  g1768(.A0(new_n1814_), .A1(new_n1809_), .B0(new_n1817_), .Y(new_n1818_));
  XOR2X1   g1769(.A(new_n1818_), .B(new_n519_), .Y(new_n1819_));
  XOR2X1   g1770(.A(new_n1774_), .B(new_n1773_), .Y(new_n1820_));
  AND2X1   g1771(.A(new_n1820_), .B(new_n1819_), .Y(new_n1821_));
  XOR2X1   g1772(.A(new_n1771_), .B(new_n1763_), .Y(new_n1822_));
  INVX1    g1773(.A(new_n1822_), .Y(new_n1823_));
  INVX1    g1774(.A(new_n1796_), .Y(new_n1824_));
  OAI22X1  g1775(.A0(new_n1805_), .A1(new_n1638_), .B0(new_n1824_), .B1(new_n1778_), .Y(new_n1825_));
  AOI21X1  g1776(.A0(new_n1801_), .A1(new_n1620_), .B0(new_n1825_), .Y(new_n1826_));
  XOR2X1   g1777(.A(new_n1660_), .B(new_n1659_), .Y(new_n1827_));
  OAI21X1  g1778(.A0(new_n1827_), .A1(new_n1810_), .B0(new_n1826_), .Y(new_n1828_));
  XOR2X1   g1779(.A(new_n1828_), .B(new_n1164_), .Y(new_n1829_));
  NAND2X1  g1780(.A(new_n1829_), .B(new_n1823_), .Y(new_n1830_));
  AOI22X1  g1781(.A0(new_n1804_), .A1(new_n1642_), .B0(new_n1796_), .B1(new_n1657_), .Y(new_n1831_));
  OAI21X1  g1782(.A0(new_n1802_), .A1(new_n1778_), .B0(new_n1831_), .Y(new_n1832_));
  AOI21X1  g1783(.A0(new_n1809_), .A1(new_n1777_), .B0(new_n1832_), .Y(new_n1833_));
  XOR2X1   g1784(.A(new_n1833_), .B(new_n1164_), .Y(new_n1834_));
  INVX1    g1785(.A(new_n1834_), .Y(new_n1835_));
  XOR2X1   g1786(.A(new_n1760_), .B(new_n1754_), .Y(new_n1836_));
  XOR2X1   g1787(.A(new_n1753_), .B(new_n1749_), .Y(new_n1837_));
  OAI22X1  g1788(.A0(new_n1805_), .A1(new_n1647_), .B0(new_n1824_), .B1(new_n1640_), .Y(new_n1838_));
  AOI21X1  g1789(.A0(new_n1801_), .A1(new_n1657_), .B0(new_n1838_), .Y(new_n1839_));
  OAI21X1  g1790(.A0(new_n1810_), .A1(new_n1743_), .B0(new_n1839_), .Y(new_n1840_));
  XOR2X1   g1791(.A(new_n1840_), .B(new_n1164_), .Y(new_n1841_));
  NAND2X1  g1792(.A(new_n1841_), .B(new_n1837_), .Y(new_n1842_));
  OAI22X1  g1793(.A0(new_n1802_), .A1(new_n1650_), .B0(new_n1824_), .B1(new_n1651_), .Y(new_n1843_));
  AOI21X1  g1794(.A0(new_n1809_), .A1(new_n1706_), .B0(new_n1843_), .Y(new_n1844_));
  XOR2X1   g1795(.A(new_n1844_), .B(new_n1164_), .Y(new_n1845_));
  NOR2X1   g1796(.A(new_n1793_), .B(new_n1651_), .Y(new_n1846_));
  OAI22X1  g1797(.A0(new_n1805_), .A1(new_n1651_), .B0(new_n1824_), .B1(new_n1650_), .Y(new_n1847_));
  AOI21X1  g1798(.A0(new_n1801_), .A1(new_n1644_), .B0(new_n1847_), .Y(new_n1848_));
  OAI21X1  g1799(.A0(new_n1810_), .A1(new_n1758_), .B0(new_n1848_), .Y(new_n1849_));
  NOR4X1   g1800(.A(new_n1849_), .B(new_n1846_), .C(new_n1845_), .D(new_n519_), .Y(new_n1850_));
  AND2X1   g1801(.A(new_n1850_), .B(new_n1748_), .Y(new_n1851_));
  INVX1    g1802(.A(new_n1851_), .Y(new_n1852_));
  OR2X1    g1803(.A(new_n1719_), .B(new_n1651_), .Y(new_n1853_));
  XOR2X1   g1804(.A(new_n1850_), .B(new_n1853_), .Y(new_n1854_));
  AOI22X1  g1805(.A0(new_n1804_), .A1(new_n1734_), .B0(new_n1796_), .B1(new_n1644_), .Y(new_n1855_));
  OAI21X1  g1806(.A0(new_n1802_), .A1(new_n1640_), .B0(new_n1855_), .Y(new_n1856_));
  AOI21X1  g1807(.A0(new_n1809_), .A1(new_n1767_), .B0(new_n1856_), .Y(new_n1857_));
  XOR2X1   g1808(.A(new_n1857_), .B(new_n1164_), .Y(new_n1858_));
  OAI21X1  g1809(.A0(new_n1858_), .A1(new_n1854_), .B0(new_n1852_), .Y(new_n1859_));
  XOR2X1   g1810(.A(new_n1841_), .B(new_n1837_), .Y(new_n1860_));
  NAND2X1  g1811(.A(new_n1860_), .B(new_n1859_), .Y(new_n1861_));
  XOR2X1   g1812(.A(new_n1836_), .B(new_n1834_), .Y(new_n1862_));
  AOI21X1  g1813(.A0(new_n1861_), .A1(new_n1842_), .B0(new_n1862_), .Y(new_n1863_));
  AOI21X1  g1814(.A0(new_n1836_), .A1(new_n1835_), .B0(new_n1863_), .Y(new_n1864_));
  XOR2X1   g1815(.A(new_n1829_), .B(new_n1822_), .Y(new_n1865_));
  OAI21X1  g1816(.A0(new_n1865_), .A1(new_n1864_), .B0(new_n1830_), .Y(new_n1866_));
  XOR2X1   g1817(.A(new_n1820_), .B(new_n1819_), .Y(new_n1867_));
  AOI21X1  g1818(.A0(new_n1867_), .A1(new_n1866_), .B0(new_n1821_), .Y(new_n1868_));
  INVX1    g1819(.A(new_n1812_), .Y(new_n1869_));
  XOR2X1   g1820(.A(new_n1869_), .B(new_n1792_), .Y(new_n1870_));
  OAI21X1  g1821(.A0(new_n1870_), .A1(new_n1868_), .B0(new_n1813_), .Y(new_n1871_));
  XOR2X1   g1822(.A(new_n1661_), .B(new_n1659_), .Y(new_n1872_));
  AOI22X1  g1823(.A0(new_n1729_), .A1(new_n1623_), .B0(new_n1727_), .B1(new_n1657_), .Y(new_n1873_));
  OAI21X1  g1824(.A0(new_n1750_), .A1(new_n1798_), .B0(new_n1873_), .Y(new_n1874_));
  AOI21X1  g1825(.A0(new_n1872_), .A1(new_n1721_), .B0(new_n1874_), .Y(new_n1875_));
  XOR2X1   g1826(.A(new_n1875_), .B(new_n312_), .Y(new_n1876_));
  INVX1    g1827(.A(new_n1785_), .Y(new_n1877_));
  AOI22X1  g1828(.A0(new_n1877_), .A1(new_n1734_), .B0(new_n1710_), .B1(new_n1644_), .Y(new_n1878_));
  OAI21X1  g1829(.A0(new_n1714_), .A1(new_n1640_), .B0(new_n1878_), .Y(new_n1879_));
  AOI21X1  g1830(.A0(new_n1767_), .A1(new_n1707_), .B0(new_n1879_), .Y(new_n1880_));
  XOR2X1   g1831(.A(new_n1880_), .B(new_n793_), .Y(new_n1881_));
  NOR4X1   g1832(.A(new_n1788_), .B(new_n1717_), .C(new_n1747_), .D(new_n793_), .Y(new_n1882_));
  NOR2X1   g1833(.A(new_n1651_), .B(new_n793_), .Y(new_n1883_));
  OR2X1    g1834(.A(new_n1883_), .B(new_n1882_), .Y(new_n1884_));
  XOR2X1   g1835(.A(new_n1883_), .B(new_n1882_), .Y(new_n1885_));
  INVX1    g1836(.A(new_n1885_), .Y(new_n1886_));
  AND2X1   g1837(.A(new_n1883_), .B(new_n1882_), .Y(new_n1887_));
  AOI21X1  g1838(.A0(new_n1885_), .A1(new_n1881_), .B0(new_n1887_), .Y(new_n1888_));
  AOI22X1  g1839(.A0(new_n1888_), .A1(new_n1884_), .B0(new_n1886_), .B1(new_n1881_), .Y(new_n1889_));
  XOR2X1   g1840(.A(new_n1889_), .B(new_n1876_), .Y(new_n1890_));
  AND2X1   g1841(.A(new_n1790_), .B(new_n1782_), .Y(new_n1891_));
  AOI21X1  g1842(.A0(new_n1791_), .A1(new_n1776_), .B0(new_n1891_), .Y(new_n1892_));
  XOR2X1   g1843(.A(new_n1892_), .B(new_n1890_), .Y(new_n1893_));
  XOR2X1   g1844(.A(new_n1797_), .B(new_n1613_), .Y(new_n1894_));
  XOR2X1   g1845(.A(new_n1894_), .B(new_n1667_), .Y(new_n1895_));
  OAI22X1  g1846(.A0(new_n1805_), .A1(new_n1815_), .B0(new_n1824_), .B1(new_n1797_), .Y(new_n1896_));
  AOI21X1  g1847(.A0(new_n1801_), .A1(new_n1613_), .B0(new_n1896_), .Y(new_n1897_));
  OAI21X1  g1848(.A0(new_n1895_), .A1(new_n1810_), .B0(new_n1897_), .Y(new_n1898_));
  XOR2X1   g1849(.A(new_n1898_), .B(new_n1164_), .Y(new_n1899_));
  XOR2X1   g1850(.A(new_n1899_), .B(new_n1893_), .Y(new_n1900_));
  INVX1    g1851(.A(new_n1900_), .Y(new_n1901_));
  XOR2X1   g1852(.A(new_n1901_), .B(new_n1871_), .Y(new_n1902_));
  XOR2X1   g1853(.A(new_n1902_), .B(new_n1703_), .Y(new_n1903_));
  XOR2X1   g1854(.A(new_n1870_), .B(new_n1868_), .Y(new_n1904_));
  XOR2X1   g1855(.A(new_n1674_), .B(new_n1672_), .Y(new_n1905_));
  INVX1    g1856(.A(new_n1696_), .Y(new_n1906_));
  AOI22X1  g1857(.A0(new_n1699_), .A1(new_n1613_), .B0(new_n1693_), .B1(new_n1584_), .Y(new_n1907_));
  OAI21X1  g1858(.A0(new_n1906_), .A1(new_n1673_), .B0(new_n1907_), .Y(new_n1908_));
  AOI21X1  g1859(.A0(new_n1905_), .A1(new_n245_), .B0(new_n1908_), .Y(new_n1909_));
  XOR2X1   g1860(.A(new_n1909_), .B(new_n229_), .Y(new_n1910_));
  NAND2X1  g1861(.A(new_n1910_), .B(new_n1904_), .Y(new_n1911_));
  XOR2X1   g1862(.A(new_n1909_), .B(new_n230_), .Y(new_n1912_));
  XOR2X1   g1863(.A(new_n1912_), .B(new_n1904_), .Y(new_n1913_));
  XOR2X1   g1864(.A(new_n1867_), .B(new_n1866_), .Y(new_n1914_));
  INVX1    g1865(.A(new_n245_), .Y(new_n1915_));
  INVX1    g1866(.A(new_n1699_), .Y(new_n1916_));
  OAI22X1  g1867(.A0(new_n1916_), .A1(new_n1797_), .B0(new_n1906_), .B1(new_n1585_), .Y(new_n1917_));
  AOI21X1  g1868(.A0(new_n1693_), .A1(new_n1613_), .B0(new_n1917_), .Y(new_n1918_));
  XOR2X1   g1869(.A(new_n1670_), .B(new_n1669_), .Y(new_n1919_));
  OAI21X1  g1870(.A0(new_n1919_), .A1(new_n1915_), .B0(new_n1918_), .Y(new_n1920_));
  XOR2X1   g1871(.A(new_n1920_), .B(new_n230_), .Y(new_n1921_));
  AND2X1   g1872(.A(new_n1921_), .B(new_n1914_), .Y(new_n1922_));
  XOR2X1   g1873(.A(new_n1865_), .B(new_n1864_), .Y(new_n1923_));
  OAI22X1  g1874(.A0(new_n1916_), .A1(new_n1815_), .B0(new_n1694_), .B1(new_n1797_), .Y(new_n1924_));
  AOI21X1  g1875(.A0(new_n1696_), .A1(new_n1613_), .B0(new_n1924_), .Y(new_n1925_));
  OAI21X1  g1876(.A0(new_n1895_), .A1(new_n1915_), .B0(new_n1925_), .Y(new_n1926_));
  XOR2X1   g1877(.A(new_n1926_), .B(new_n230_), .Y(new_n1927_));
  NAND2X1  g1878(.A(new_n1927_), .B(new_n1923_), .Y(new_n1928_));
  INVX1    g1879(.A(new_n1928_), .Y(new_n1929_));
  AND2X1   g1880(.A(new_n1861_), .B(new_n1842_), .Y(new_n1930_));
  XOR2X1   g1881(.A(new_n1862_), .B(new_n1930_), .Y(new_n1931_));
  OAI22X1  g1882(.A0(new_n1916_), .A1(new_n1798_), .B0(new_n1906_), .B1(new_n1797_), .Y(new_n1932_));
  AOI21X1  g1883(.A0(new_n1693_), .A1(new_n1618_), .B0(new_n1932_), .Y(new_n1933_));
  OAI21X1  g1884(.A0(new_n1808_), .A1(new_n1915_), .B0(new_n1933_), .Y(new_n1934_));
  XOR2X1   g1885(.A(new_n1934_), .B(new_n230_), .Y(new_n1935_));
  NAND2X1  g1886(.A(new_n1935_), .B(new_n1931_), .Y(new_n1936_));
  AOI22X1  g1887(.A0(new_n1699_), .A1(new_n1623_), .B0(new_n1693_), .B1(new_n1620_), .Y(new_n1937_));
  OAI21X1  g1888(.A0(new_n1906_), .A1(new_n1815_), .B0(new_n1937_), .Y(new_n1938_));
  AOI21X1  g1889(.A0(new_n1814_), .A1(new_n245_), .B0(new_n1938_), .Y(new_n1939_));
  XOR2X1   g1890(.A(new_n1939_), .B(new_n229_), .Y(new_n1940_));
  XOR2X1   g1891(.A(new_n1860_), .B(new_n1859_), .Y(new_n1941_));
  AND2X1   g1892(.A(new_n1941_), .B(new_n1940_), .Y(new_n1942_));
  XOR2X1   g1893(.A(new_n1858_), .B(new_n1854_), .Y(new_n1943_));
  OAI22X1  g1894(.A0(new_n1916_), .A1(new_n1638_), .B0(new_n1694_), .B1(new_n1778_), .Y(new_n1944_));
  AOI21X1  g1895(.A0(new_n1696_), .A1(new_n1620_), .B0(new_n1944_), .Y(new_n1945_));
  OAI21X1  g1896(.A0(new_n1827_), .A1(new_n1915_), .B0(new_n1945_), .Y(new_n1946_));
  XOR2X1   g1897(.A(new_n1946_), .B(new_n230_), .Y(new_n1947_));
  AND2X1   g1898(.A(new_n1947_), .B(new_n1943_), .Y(new_n1948_));
  AOI22X1  g1899(.A0(new_n1699_), .A1(new_n1642_), .B0(new_n1693_), .B1(new_n1657_), .Y(new_n1949_));
  OAI21X1  g1900(.A0(new_n1906_), .A1(new_n1778_), .B0(new_n1949_), .Y(new_n1950_));
  AOI21X1  g1901(.A0(new_n1777_), .A1(new_n245_), .B0(new_n1950_), .Y(new_n1951_));
  XOR2X1   g1902(.A(new_n1951_), .B(new_n229_), .Y(new_n1952_));
  OAI21X1  g1903(.A0(new_n1793_), .A1(new_n1651_), .B0(new_n1164_), .Y(new_n1953_));
  NOR2X1   g1904(.A(new_n1953_), .B(new_n1845_), .Y(new_n1954_));
  XOR2X1   g1905(.A(new_n1849_), .B(new_n1164_), .Y(new_n1955_));
  XOR2X1   g1906(.A(new_n1955_), .B(new_n1954_), .Y(new_n1956_));
  NAND2X1  g1907(.A(new_n1956_), .B(new_n1952_), .Y(new_n1957_));
  XOR2X1   g1908(.A(new_n1953_), .B(new_n1845_), .Y(new_n1958_));
  OAI22X1  g1909(.A0(new_n1916_), .A1(new_n1647_), .B0(new_n1694_), .B1(new_n1640_), .Y(new_n1959_));
  AOI21X1  g1910(.A0(new_n1696_), .A1(new_n1657_), .B0(new_n1959_), .Y(new_n1960_));
  OAI21X1  g1911(.A0(new_n1743_), .A1(new_n1915_), .B0(new_n1960_), .Y(new_n1961_));
  XOR2X1   g1912(.A(new_n1961_), .B(new_n230_), .Y(new_n1962_));
  NAND2X1  g1913(.A(new_n1962_), .B(new_n1958_), .Y(new_n1963_));
  NOR2X1   g1914(.A(new_n1651_), .B(new_n244_), .Y(new_n1964_));
  NOR2X1   g1915(.A(new_n1964_), .B(new_n229_), .Y(new_n1965_));
  OAI22X1  g1916(.A0(new_n1906_), .A1(new_n1650_), .B0(new_n1694_), .B1(new_n1651_), .Y(new_n1966_));
  AOI21X1  g1917(.A0(new_n1706_), .A1(new_n245_), .B0(new_n1966_), .Y(new_n1967_));
  XOR2X1   g1918(.A(new_n1967_), .B(new_n229_), .Y(new_n1968_));
  AND2X1   g1919(.A(new_n1968_), .B(new_n1965_), .Y(new_n1969_));
  OAI22X1  g1920(.A0(new_n1916_), .A1(new_n1651_), .B0(new_n1694_), .B1(new_n1650_), .Y(new_n1970_));
  AOI21X1  g1921(.A0(new_n1696_), .A1(new_n1644_), .B0(new_n1970_), .Y(new_n1971_));
  OAI21X1  g1922(.A0(new_n1758_), .A1(new_n1915_), .B0(new_n1971_), .Y(new_n1972_));
  XOR2X1   g1923(.A(new_n1972_), .B(new_n230_), .Y(new_n1973_));
  NAND3X1  g1924(.A(new_n1973_), .B(new_n1969_), .C(new_n1846_), .Y(new_n1974_));
  AND2X1   g1925(.A(new_n1973_), .B(new_n1969_), .Y(new_n1975_));
  XOR2X1   g1926(.A(new_n1975_), .B(new_n1846_), .Y(new_n1976_));
  AOI22X1  g1927(.A0(new_n1699_), .A1(new_n1734_), .B0(new_n1693_), .B1(new_n1644_), .Y(new_n1977_));
  OAI21X1  g1928(.A0(new_n1906_), .A1(new_n1640_), .B0(new_n1977_), .Y(new_n1978_));
  AOI21X1  g1929(.A0(new_n1767_), .A1(new_n245_), .B0(new_n1978_), .Y(new_n1979_));
  XOR2X1   g1930(.A(new_n1979_), .B(new_n229_), .Y(new_n1980_));
  NAND2X1  g1931(.A(new_n1980_), .B(new_n1976_), .Y(new_n1981_));
  NAND2X1  g1932(.A(new_n1981_), .B(new_n1974_), .Y(new_n1982_));
  XOR2X1   g1933(.A(new_n1962_), .B(new_n1958_), .Y(new_n1983_));
  NAND2X1  g1934(.A(new_n1983_), .B(new_n1982_), .Y(new_n1984_));
  NAND2X1  g1935(.A(new_n1984_), .B(new_n1963_), .Y(new_n1985_));
  XOR2X1   g1936(.A(new_n1956_), .B(new_n1952_), .Y(new_n1986_));
  NAND2X1  g1937(.A(new_n1986_), .B(new_n1985_), .Y(new_n1987_));
  INVX1    g1938(.A(new_n1943_), .Y(new_n1988_));
  XOR2X1   g1939(.A(new_n1947_), .B(new_n1988_), .Y(new_n1989_));
  AOI21X1  g1940(.A0(new_n1987_), .A1(new_n1957_), .B0(new_n1989_), .Y(new_n1990_));
  OR2X1    g1941(.A(new_n1990_), .B(new_n1948_), .Y(new_n1991_));
  XOR2X1   g1942(.A(new_n1941_), .B(new_n1940_), .Y(new_n1992_));
  AOI21X1  g1943(.A0(new_n1992_), .A1(new_n1991_), .B0(new_n1942_), .Y(new_n1993_));
  XOR2X1   g1944(.A(new_n1935_), .B(new_n1931_), .Y(new_n1994_));
  INVX1    g1945(.A(new_n1994_), .Y(new_n1995_));
  OR2X1    g1946(.A(new_n1995_), .B(new_n1993_), .Y(new_n1996_));
  INVX1    g1947(.A(new_n1927_), .Y(new_n1997_));
  XOR2X1   g1948(.A(new_n1997_), .B(new_n1923_), .Y(new_n1998_));
  AOI21X1  g1949(.A0(new_n1996_), .A1(new_n1936_), .B0(new_n1998_), .Y(new_n1999_));
  OR2X1    g1950(.A(new_n1999_), .B(new_n1929_), .Y(new_n2000_));
  XOR2X1   g1951(.A(new_n1921_), .B(new_n1914_), .Y(new_n2001_));
  AOI21X1  g1952(.A0(new_n2001_), .A1(new_n2000_), .B0(new_n1922_), .Y(new_n2002_));
  OAI21X1  g1953(.A0(new_n2002_), .A1(new_n1913_), .B0(new_n1911_), .Y(new_n2003_));
  XOR2X1   g1954(.A(new_n2003_), .B(new_n1903_), .Y(new_n2004_));
  AND2X1   g1955(.A(new_n50_), .B(\a[0] ), .Y(new_n2005_));
  XOR2X1   g1956(.A(new_n2005_), .B(new_n241_), .Y(new_n2006_));
  XOR2X1   g1957(.A(new_n2006_), .B(new_n243_), .Y(new_n2007_));
  NOR2X1   g1958(.A(new_n2007_), .B(new_n240_), .Y(new_n2008_));
  INVX1    g1959(.A(new_n2008_), .Y(new_n2009_));
  AND2X1   g1960(.A(new_n2007_), .B(\a[0] ), .Y(new_n2010_));
  OR4X1    g1961(.A(new_n483_), .B(new_n358_), .C(new_n280_), .D(new_n211_), .Y(new_n2011_));
  OR2X1    g1962(.A(new_n147_), .B(new_n139_), .Y(new_n2012_));
  OR4X1    g1963(.A(new_n2012_), .B(new_n1455_), .C(new_n547_), .D(new_n497_), .Y(new_n2013_));
  OR2X1    g1964(.A(new_n2013_), .B(new_n2011_), .Y(new_n2014_));
  OR4X1    g1965(.A(new_n2014_), .B(new_n1404_), .C(new_n1345_), .D(new_n324_), .Y(new_n2015_));
  NOR2X1   g1966(.A(new_n2015_), .B(new_n384_), .Y(new_n2016_));
  INVX1    g1967(.A(new_n2016_), .Y(new_n2017_));
  OR4X1    g1968(.A(new_n527_), .B(new_n551_), .C(new_n437_), .D(new_n193_), .Y(new_n2018_));
  OR4X1    g1969(.A(new_n330_), .B(new_n337_), .C(new_n281_), .D(new_n272_), .Y(new_n2019_));
  OR4X1    g1970(.A(new_n2019_), .B(new_n348_), .C(new_n189_), .D(new_n121_), .Y(new_n2020_));
  OR2X1    g1971(.A(new_n204_), .B(new_n202_), .Y(new_n2021_));
  OR4X1    g1972(.A(new_n314_), .B(new_n251_), .C(new_n149_), .D(new_n110_), .Y(new_n2022_));
  OR2X1    g1973(.A(new_n2022_), .B(new_n2021_), .Y(new_n2023_));
  NOR4X1   g1974(.A(new_n2023_), .B(new_n2020_), .C(new_n2018_), .D(new_n161_), .Y(new_n2024_));
  INVX1    g1975(.A(new_n2024_), .Y(new_n2025_));
  NOR4X1   g1976(.A(new_n616_), .B(new_n315_), .C(new_n256_), .D(new_n113_), .Y(new_n2026_));
  NAND3X1  g1977(.A(new_n2026_), .B(new_n1424_), .C(new_n217_), .Y(new_n2027_));
  OR4X1    g1978(.A(new_n184_), .B(new_n172_), .C(new_n165_), .D(new_n123_), .Y(new_n2028_));
  OR4X1    g1979(.A(new_n2028_), .B(new_n431_), .C(new_n429_), .D(new_n181_), .Y(new_n2029_));
  OR4X1    g1980(.A(new_n2029_), .B(new_n2027_), .C(new_n2025_), .D(new_n428_), .Y(new_n2030_));
  NOR4X1   g1981(.A(new_n2030_), .B(new_n2017_), .C(new_n1687_), .D(new_n1678_), .Y(new_n2031_));
  OR2X1    g1982(.A(new_n264_), .B(new_n216_), .Y(new_n2032_));
  OR2X1    g1983(.A(new_n379_), .B(new_n189_), .Y(new_n2033_));
  OR4X1    g1984(.A(new_n2033_), .B(new_n2032_), .C(new_n332_), .D(new_n252_), .Y(new_n2034_));
  OR4X1    g1985(.A(new_n733_), .B(new_n388_), .C(new_n196_), .D(new_n125_), .Y(new_n2035_));
  OR4X1    g1986(.A(new_n2035_), .B(new_n2034_), .C(new_n395_), .D(new_n342_), .Y(new_n2036_));
  OR4X1    g1987(.A(new_n370_), .B(new_n324_), .C(new_n261_), .D(new_n134_), .Y(new_n2037_));
  NOR3X1   g1988(.A(new_n2037_), .B(new_n2036_), .C(new_n365_), .Y(new_n2038_));
  XOR2X1   g1989(.A(new_n2038_), .B(new_n2031_), .Y(new_n2039_));
  INVX1    g1990(.A(new_n2039_), .Y(new_n2040_));
  NOR3X1   g1991(.A(new_n239_), .B(\a[1] ), .C(\a[0] ), .Y(new_n2041_));
  INVX1    g1992(.A(new_n2041_), .Y(new_n2042_));
  NOR2X1   g1993(.A(new_n1687_), .B(new_n1678_), .Y(new_n2043_));
  XOR2X1   g1994(.A(new_n2030_), .B(new_n2043_), .Y(new_n2044_));
  INVX1    g1995(.A(new_n2044_), .Y(new_n2045_));
  NOR3X1   g1996(.A(new_n2030_), .B(new_n1687_), .C(new_n1678_), .Y(new_n2046_));
  XOR2X1   g1997(.A(new_n2046_), .B(new_n2016_), .Y(new_n2047_));
  AND2X1   g1998(.A(\a[1] ), .B(new_n240_), .Y(new_n2048_));
  INVX1    g1999(.A(new_n2048_), .Y(new_n2049_));
  OAI22X1  g2000(.A0(new_n2049_), .A1(new_n2047_), .B0(new_n2045_), .B1(new_n2042_), .Y(new_n2050_));
  AOI21X1  g2001(.A0(new_n2040_), .A1(new_n2010_), .B0(new_n2050_), .Y(new_n2051_));
  INVX1    g2002(.A(new_n2047_), .Y(new_n2052_));
  NAND2X1  g2003(.A(new_n2052_), .B(new_n2044_), .Y(new_n2053_));
  AND2X1   g2004(.A(new_n2044_), .B(new_n1695_), .Y(new_n2054_));
  NAND2X1  g2005(.A(new_n1695_), .B(new_n1676_), .Y(new_n2055_));
  OAI21X1  g2006(.A0(new_n1689_), .A1(new_n1675_), .B0(new_n2055_), .Y(new_n2056_));
  XOR2X1   g2007(.A(new_n2044_), .B(new_n1695_), .Y(new_n2057_));
  AOI21X1  g2008(.A0(new_n2057_), .A1(new_n2056_), .B0(new_n2054_), .Y(new_n2058_));
  XOR2X1   g2009(.A(new_n2047_), .B(new_n2044_), .Y(new_n2059_));
  OAI21X1  g2010(.A0(new_n2059_), .A1(new_n2058_), .B0(new_n2053_), .Y(new_n2060_));
  XOR2X1   g2011(.A(new_n2047_), .B(new_n2039_), .Y(new_n2061_));
  INVX1    g2012(.A(new_n2061_), .Y(new_n2062_));
  XOR2X1   g2013(.A(new_n2062_), .B(new_n2060_), .Y(new_n2063_));
  OAI21X1  g2014(.A0(new_n2063_), .A1(new_n2009_), .B0(new_n2051_), .Y(new_n2064_));
  XOR2X1   g2015(.A(new_n2064_), .B(new_n243_), .Y(new_n2065_));
  AND2X1   g2016(.A(new_n2065_), .B(new_n2004_), .Y(new_n2066_));
  XOR2X1   g2017(.A(new_n2002_), .B(new_n1913_), .Y(new_n2067_));
  OAI22X1  g2018(.A0(new_n2049_), .A1(new_n2045_), .B0(new_n2042_), .B1(new_n1688_), .Y(new_n2068_));
  AOI21X1  g2019(.A0(new_n2052_), .A1(new_n2010_), .B0(new_n2068_), .Y(new_n2069_));
  INVX1    g2020(.A(new_n2059_), .Y(new_n2070_));
  XOR2X1   g2021(.A(new_n2070_), .B(new_n2058_), .Y(new_n2071_));
  OAI21X1  g2022(.A0(new_n2071_), .A1(new_n2009_), .B0(new_n2069_), .Y(new_n2072_));
  XOR2X1   g2023(.A(new_n2072_), .B(new_n243_), .Y(new_n2073_));
  NAND2X1  g2024(.A(new_n2073_), .B(new_n2067_), .Y(new_n2074_));
  XOR2X1   g2025(.A(new_n2057_), .B(new_n2056_), .Y(new_n2075_));
  INVX1    g2026(.A(new_n2010_), .Y(new_n2076_));
  AOI22X1  g2027(.A0(new_n2048_), .A1(new_n1695_), .B0(new_n2041_), .B1(new_n1676_), .Y(new_n2077_));
  OAI21X1  g2028(.A0(new_n2045_), .A1(new_n2076_), .B0(new_n2077_), .Y(new_n2078_));
  AOI21X1  g2029(.A0(new_n2075_), .A1(new_n2008_), .B0(new_n2078_), .Y(new_n2079_));
  XOR2X1   g2030(.A(new_n2079_), .B(new_n243_), .Y(new_n2080_));
  INVX1    g2031(.A(new_n243_), .Y(new_n2081_));
  OAI21X1  g2032(.A0(new_n1766_), .A1(new_n1765_), .B0(new_n2008_), .Y(new_n2082_));
  NOR2X1   g2033(.A(new_n2076_), .B(new_n1640_), .Y(new_n2083_));
  OAI22X1  g2034(.A0(new_n2049_), .A1(new_n1647_), .B0(new_n2042_), .B1(new_n1650_), .Y(new_n2084_));
  NOR2X1   g2035(.A(new_n2084_), .B(new_n2083_), .Y(new_n2085_));
  NAND3X1  g2036(.A(new_n2085_), .B(new_n2082_), .C(new_n2081_), .Y(new_n2086_));
  AOI22X1  g2037(.A0(new_n2048_), .A1(new_n1734_), .B0(new_n2041_), .B1(new_n1735_), .Y(new_n2087_));
  OAI21X1  g2038(.A0(new_n2076_), .A1(new_n1647_), .B0(new_n2087_), .Y(new_n2088_));
  AND2X1   g2039(.A(new_n2088_), .B(new_n243_), .Y(new_n2089_));
  NOR3X1   g2040(.A(new_n2007_), .B(new_n2081_), .C(new_n240_), .Y(new_n2090_));
  INVX1    g2041(.A(new_n2090_), .Y(new_n2091_));
  NOR2X1   g2042(.A(new_n2091_), .B(new_n1758_), .Y(new_n2092_));
  AND2X1   g2043(.A(new_n2090_), .B(new_n1706_), .Y(new_n2093_));
  OAI21X1  g2044(.A0(new_n1651_), .A1(new_n240_), .B0(new_n243_), .Y(new_n2094_));
  AOI21X1  g2045(.A0(new_n2048_), .A1(new_n1735_), .B0(new_n2094_), .Y(new_n2095_));
  OAI21X1  g2046(.A0(new_n2076_), .A1(new_n1650_), .B0(new_n2095_), .Y(new_n2096_));
  OR2X1    g2047(.A(new_n2096_), .B(new_n2093_), .Y(new_n2097_));
  NOR3X1   g2048(.A(new_n2097_), .B(new_n2092_), .C(new_n2089_), .Y(new_n2098_));
  OR2X1    g2049(.A(new_n2098_), .B(new_n1964_), .Y(new_n2099_));
  OR2X1    g2050(.A(new_n1764_), .B(new_n1736_), .Y(new_n2100_));
  NAND3X1  g2051(.A(new_n1653_), .B(new_n1736_), .C(new_n1733_), .Y(new_n2101_));
  AOI21X1  g2052(.A0(new_n2101_), .A1(new_n2100_), .B0(new_n2009_), .Y(new_n2102_));
  OR2X1    g2053(.A(new_n2084_), .B(new_n2083_), .Y(new_n2103_));
  OAI21X1  g2054(.A0(new_n2103_), .A1(new_n2102_), .B0(new_n243_), .Y(new_n2104_));
  NAND3X1  g2055(.A(new_n2104_), .B(new_n2099_), .C(new_n2086_), .Y(new_n2105_));
  INVX1    g2056(.A(new_n1964_), .Y(new_n2106_));
  NOR4X1   g2057(.A(new_n2097_), .B(new_n2092_), .C(new_n2089_), .D(new_n2106_), .Y(new_n2107_));
  INVX1    g2058(.A(new_n2107_), .Y(new_n2108_));
  XOR2X1   g2059(.A(new_n1968_), .B(new_n1965_), .Y(new_n2109_));
  INVX1    g2060(.A(new_n2109_), .Y(new_n2110_));
  NAND3X1  g2061(.A(new_n2110_), .B(new_n2108_), .C(new_n2105_), .Y(new_n2111_));
  AOI22X1  g2062(.A0(new_n2048_), .A1(new_n1642_), .B0(new_n2041_), .B1(new_n1644_), .Y(new_n2112_));
  OAI21X1  g2063(.A0(new_n2076_), .A1(new_n1638_), .B0(new_n2112_), .Y(new_n2113_));
  NOR2X1   g2064(.A(new_n2113_), .B(new_n243_), .Y(new_n2114_));
  OAI21X1  g2065(.A0(new_n2009_), .A1(new_n1743_), .B0(new_n2114_), .Y(new_n2115_));
  OR2X1    g2066(.A(new_n1742_), .B(new_n1740_), .Y(new_n2116_));
  AOI22X1  g2067(.A0(new_n2113_), .A1(new_n243_), .B0(new_n2090_), .B1(new_n2116_), .Y(new_n2117_));
  AND2X1   g2068(.A(new_n2117_), .B(new_n2115_), .Y(new_n2118_));
  AOI21X1  g2069(.A0(new_n2108_), .A1(new_n2105_), .B0(new_n2110_), .Y(new_n2119_));
  AOI21X1  g2070(.A0(new_n2118_), .A1(new_n2111_), .B0(new_n2119_), .Y(new_n2120_));
  AOI22X1  g2071(.A0(new_n2048_), .A1(new_n1657_), .B0(new_n2041_), .B1(new_n1642_), .Y(new_n2121_));
  OAI21X1  g2072(.A0(new_n2076_), .A1(new_n1778_), .B0(new_n2121_), .Y(new_n2122_));
  AOI21X1  g2073(.A0(new_n2008_), .A1(new_n1777_), .B0(new_n2122_), .Y(new_n2123_));
  XOR2X1   g2074(.A(new_n2123_), .B(new_n243_), .Y(new_n2124_));
  XOR2X1   g2075(.A(new_n1973_), .B(new_n1969_), .Y(new_n2125_));
  INVX1    g2076(.A(new_n2125_), .Y(new_n2126_));
  AOI21X1  g2077(.A0(new_n2124_), .A1(new_n2120_), .B0(new_n2126_), .Y(new_n2127_));
  NOR3X1   g2078(.A(new_n2103_), .B(new_n2102_), .C(new_n243_), .Y(new_n2128_));
  NOR2X1   g2079(.A(new_n2098_), .B(new_n1964_), .Y(new_n2129_));
  AOI21X1  g2080(.A0(new_n2085_), .A1(new_n2082_), .B0(new_n2081_), .Y(new_n2130_));
  NOR3X1   g2081(.A(new_n2130_), .B(new_n2129_), .C(new_n2128_), .Y(new_n2131_));
  NOR3X1   g2082(.A(new_n2109_), .B(new_n2107_), .C(new_n2131_), .Y(new_n2132_));
  NAND2X1  g2083(.A(new_n2117_), .B(new_n2115_), .Y(new_n2133_));
  OAI21X1  g2084(.A0(new_n2107_), .A1(new_n2131_), .B0(new_n2109_), .Y(new_n2134_));
  OAI21X1  g2085(.A0(new_n2133_), .A1(new_n2132_), .B0(new_n2134_), .Y(new_n2135_));
  XOR2X1   g2086(.A(new_n2123_), .B(new_n2081_), .Y(new_n2136_));
  AND2X1   g2087(.A(new_n2136_), .B(new_n2135_), .Y(new_n2137_));
  XOR2X1   g2088(.A(new_n1980_), .B(new_n1976_), .Y(new_n2138_));
  NOR3X1   g2089(.A(new_n2138_), .B(new_n2137_), .C(new_n2127_), .Y(new_n2139_));
  OAI22X1  g2090(.A0(new_n2049_), .A1(new_n1778_), .B0(new_n2042_), .B1(new_n1638_), .Y(new_n2140_));
  AOI21X1  g2091(.A0(new_n2010_), .A1(new_n1620_), .B0(new_n2140_), .Y(new_n2141_));
  NAND2X1  g2092(.A(new_n2141_), .B(new_n2081_), .Y(new_n2142_));
  AOI21X1  g2093(.A0(new_n2008_), .A1(new_n1872_), .B0(new_n2142_), .Y(new_n2143_));
  OAI22X1  g2094(.A0(new_n2141_), .A1(new_n2081_), .B0(new_n2091_), .B1(new_n1827_), .Y(new_n2144_));
  OR2X1    g2095(.A(new_n2144_), .B(new_n2143_), .Y(new_n2145_));
  OAI21X1  g2096(.A0(new_n2137_), .A1(new_n2127_), .B0(new_n2138_), .Y(new_n2146_));
  OAI21X1  g2097(.A0(new_n2145_), .A1(new_n2139_), .B0(new_n2146_), .Y(new_n2147_));
  AOI22X1  g2098(.A0(new_n2048_), .A1(new_n1620_), .B0(new_n2041_), .B1(new_n1623_), .Y(new_n2148_));
  OAI21X1  g2099(.A0(new_n2076_), .A1(new_n1815_), .B0(new_n2148_), .Y(new_n2149_));
  AOI21X1  g2100(.A0(new_n2008_), .A1(new_n1814_), .B0(new_n2149_), .Y(new_n2150_));
  XOR2X1   g2101(.A(new_n2150_), .B(new_n2081_), .Y(new_n2151_));
  XOR2X1   g2102(.A(new_n1983_), .B(new_n1982_), .Y(new_n2152_));
  OAI21X1  g2103(.A0(new_n2151_), .A1(new_n2147_), .B0(new_n2152_), .Y(new_n2153_));
  OAI21X1  g2104(.A0(new_n2136_), .A1(new_n2135_), .B0(new_n2125_), .Y(new_n2154_));
  NAND2X1  g2105(.A(new_n2136_), .B(new_n2135_), .Y(new_n2155_));
  INVX1    g2106(.A(new_n2138_), .Y(new_n2156_));
  NAND3X1  g2107(.A(new_n2156_), .B(new_n2155_), .C(new_n2154_), .Y(new_n2157_));
  NOR2X1   g2108(.A(new_n2144_), .B(new_n2143_), .Y(new_n2158_));
  AOI21X1  g2109(.A0(new_n2155_), .A1(new_n2154_), .B0(new_n2156_), .Y(new_n2159_));
  AOI21X1  g2110(.A0(new_n2158_), .A1(new_n2157_), .B0(new_n2159_), .Y(new_n2160_));
  XOR2X1   g2111(.A(new_n2150_), .B(new_n243_), .Y(new_n2161_));
  OR2X1    g2112(.A(new_n2161_), .B(new_n2160_), .Y(new_n2162_));
  AND2X1   g2113(.A(new_n1984_), .B(new_n1963_), .Y(new_n2163_));
  XOR2X1   g2114(.A(new_n1986_), .B(new_n2163_), .Y(new_n2164_));
  NAND3X1  g2115(.A(new_n2164_), .B(new_n2162_), .C(new_n2153_), .Y(new_n2165_));
  OR2X1    g2116(.A(new_n2009_), .B(new_n1808_), .Y(new_n2166_));
  OAI22X1  g2117(.A0(new_n2042_), .A1(new_n1798_), .B0(new_n2076_), .B1(new_n1797_), .Y(new_n2167_));
  AOI21X1  g2118(.A0(new_n2048_), .A1(new_n1618_), .B0(new_n2167_), .Y(new_n2168_));
  AND2X1   g2119(.A(new_n2168_), .B(new_n2081_), .Y(new_n2169_));
  OAI22X1  g2120(.A0(new_n2168_), .A1(new_n2081_), .B0(new_n2091_), .B1(new_n1808_), .Y(new_n2170_));
  AOI21X1  g2121(.A0(new_n2169_), .A1(new_n2166_), .B0(new_n2170_), .Y(new_n2171_));
  AOI21X1  g2122(.A0(new_n2162_), .A1(new_n2153_), .B0(new_n2164_), .Y(new_n2172_));
  AOI21X1  g2123(.A0(new_n2171_), .A1(new_n2165_), .B0(new_n2172_), .Y(new_n2173_));
  NAND2X1  g2124(.A(new_n1987_), .B(new_n1957_), .Y(new_n2174_));
  XOR2X1   g2125(.A(new_n1989_), .B(new_n2174_), .Y(new_n2175_));
  AND2X1   g2126(.A(new_n2010_), .B(new_n1613_), .Y(new_n2176_));
  OAI22X1  g2127(.A0(new_n2049_), .A1(new_n1797_), .B0(new_n2042_), .B1(new_n1815_), .Y(new_n2177_));
  NOR3X1   g2128(.A(new_n2177_), .B(new_n2176_), .C(new_n243_), .Y(new_n2178_));
  OAI21X1  g2129(.A0(new_n2009_), .A1(new_n1895_), .B0(new_n2178_), .Y(new_n2179_));
  XOR2X1   g2130(.A(new_n1668_), .B(new_n1667_), .Y(new_n2180_));
  OR2X1    g2131(.A(new_n2177_), .B(new_n2176_), .Y(new_n2181_));
  AOI22X1  g2132(.A0(new_n2181_), .A1(new_n243_), .B0(new_n2090_), .B1(new_n2180_), .Y(new_n2182_));
  NAND2X1  g2133(.A(new_n2182_), .B(new_n2179_), .Y(new_n2183_));
  AOI21X1  g2134(.A0(new_n2175_), .A1(new_n2173_), .B0(new_n2183_), .Y(new_n2184_));
  INVX1    g2135(.A(new_n2152_), .Y(new_n2185_));
  AOI21X1  g2136(.A0(new_n2161_), .A1(new_n2160_), .B0(new_n2185_), .Y(new_n2186_));
  NOR2X1   g2137(.A(new_n2161_), .B(new_n2160_), .Y(new_n2187_));
  XOR2X1   g2138(.A(new_n1986_), .B(new_n1985_), .Y(new_n2188_));
  NOR3X1   g2139(.A(new_n2188_), .B(new_n2187_), .C(new_n2186_), .Y(new_n2189_));
  INVX1    g2140(.A(new_n2171_), .Y(new_n2190_));
  OAI21X1  g2141(.A0(new_n2187_), .A1(new_n2186_), .B0(new_n2188_), .Y(new_n2191_));
  OAI21X1  g2142(.A0(new_n2190_), .A1(new_n2189_), .B0(new_n2191_), .Y(new_n2192_));
  AND2X1   g2143(.A(new_n1987_), .B(new_n1957_), .Y(new_n2193_));
  XOR2X1   g2144(.A(new_n1989_), .B(new_n2193_), .Y(new_n2194_));
  AND2X1   g2145(.A(new_n2194_), .B(new_n2192_), .Y(new_n2195_));
  XOR2X1   g2146(.A(new_n1992_), .B(new_n1991_), .Y(new_n2196_));
  NOR3X1   g2147(.A(new_n2196_), .B(new_n2195_), .C(new_n2184_), .Y(new_n2197_));
  INVX1    g2148(.A(new_n1613_), .Y(new_n2198_));
  AOI22X1  g2149(.A0(new_n2041_), .A1(new_n1615_), .B0(new_n2010_), .B1(new_n1584_), .Y(new_n2199_));
  OAI21X1  g2150(.A0(new_n2049_), .A1(new_n2198_), .B0(new_n2199_), .Y(new_n2200_));
  NOR2X1   g2151(.A(new_n2200_), .B(new_n243_), .Y(new_n2201_));
  OAI21X1  g2152(.A0(new_n2009_), .A1(new_n1919_), .B0(new_n2201_), .Y(new_n2202_));
  NOR2X1   g2153(.A(new_n2091_), .B(new_n1919_), .Y(new_n2203_));
  AOI21X1  g2154(.A0(new_n2200_), .A1(new_n243_), .B0(new_n2203_), .Y(new_n2204_));
  NAND2X1  g2155(.A(new_n2204_), .B(new_n2202_), .Y(new_n2205_));
  OAI21X1  g2156(.A0(new_n2195_), .A1(new_n2184_), .B0(new_n2196_), .Y(new_n2206_));
  OAI21X1  g2157(.A0(new_n2205_), .A1(new_n2197_), .B0(new_n2206_), .Y(new_n2207_));
  XOR2X1   g2158(.A(new_n1995_), .B(new_n1993_), .Y(new_n2208_));
  AOI22X1  g2159(.A0(new_n2048_), .A1(new_n1584_), .B0(new_n2041_), .B1(new_n1613_), .Y(new_n2209_));
  OAI21X1  g2160(.A0(new_n2076_), .A1(new_n1673_), .B0(new_n2209_), .Y(new_n2210_));
  AOI21X1  g2161(.A0(new_n2008_), .A1(new_n1905_), .B0(new_n2210_), .Y(new_n2211_));
  XOR2X1   g2162(.A(new_n2211_), .B(new_n2081_), .Y(new_n2212_));
  AOI21X1  g2163(.A0(new_n2208_), .A1(new_n2207_), .B0(new_n2212_), .Y(new_n2213_));
  AND2X1   g2164(.A(new_n2182_), .B(new_n2179_), .Y(new_n2214_));
  OAI21X1  g2165(.A0(new_n2194_), .A1(new_n2192_), .B0(new_n2214_), .Y(new_n2215_));
  NAND2X1  g2166(.A(new_n2194_), .B(new_n2192_), .Y(new_n2216_));
  NOR2X1   g2167(.A(new_n1990_), .B(new_n1948_), .Y(new_n2217_));
  XOR2X1   g2168(.A(new_n1992_), .B(new_n2217_), .Y(new_n2218_));
  NAND3X1  g2169(.A(new_n2218_), .B(new_n2216_), .C(new_n2215_), .Y(new_n2219_));
  AND2X1   g2170(.A(new_n2204_), .B(new_n2202_), .Y(new_n2220_));
  AOI21X1  g2171(.A0(new_n2216_), .A1(new_n2215_), .B0(new_n2218_), .Y(new_n2221_));
  AOI21X1  g2172(.A0(new_n2220_), .A1(new_n2219_), .B0(new_n2221_), .Y(new_n2222_));
  INVX1    g2173(.A(new_n2208_), .Y(new_n2223_));
  AND2X1   g2174(.A(new_n2223_), .B(new_n2222_), .Y(new_n2224_));
  OAI21X1  g2175(.A0(new_n1995_), .A1(new_n1993_), .B0(new_n1936_), .Y(new_n2225_));
  XOR2X1   g2176(.A(new_n1998_), .B(new_n2225_), .Y(new_n2226_));
  OAI21X1  g2177(.A0(new_n2224_), .A1(new_n2213_), .B0(new_n2226_), .Y(new_n2227_));
  AOI22X1  g2178(.A0(new_n2041_), .A1(new_n1584_), .B0(new_n2010_), .B1(new_n1695_), .Y(new_n2228_));
  OAI21X1  g2179(.A0(new_n2049_), .A1(new_n1673_), .B0(new_n2228_), .Y(new_n2229_));
  AOI21X1  g2180(.A0(new_n2008_), .A1(new_n1690_), .B0(new_n2229_), .Y(new_n2230_));
  XOR2X1   g2181(.A(new_n2230_), .B(new_n2081_), .Y(new_n2231_));
  NOR3X1   g2182(.A(new_n2226_), .B(new_n2224_), .C(new_n2213_), .Y(new_n2232_));
  AOI21X1  g2183(.A0(new_n2231_), .A1(new_n2227_), .B0(new_n2232_), .Y(new_n2233_));
  XOR2X1   g2184(.A(new_n2001_), .B(new_n2000_), .Y(new_n2234_));
  INVX1    g2185(.A(new_n2234_), .Y(new_n2235_));
  AOI21X1  g2186(.A0(new_n2233_), .A1(new_n2080_), .B0(new_n2235_), .Y(new_n2236_));
  NOR2X1   g2187(.A(new_n2233_), .B(new_n2080_), .Y(new_n2237_));
  XOR2X1   g2188(.A(new_n2073_), .B(new_n2067_), .Y(new_n2238_));
  OAI21X1  g2189(.A0(new_n2237_), .A1(new_n2236_), .B0(new_n2238_), .Y(new_n2239_));
  XOR2X1   g2190(.A(new_n2064_), .B(new_n2081_), .Y(new_n2240_));
  XOR2X1   g2191(.A(new_n2240_), .B(new_n2004_), .Y(new_n2241_));
  AOI21X1  g2192(.A0(new_n2239_), .A1(new_n2074_), .B0(new_n2241_), .Y(new_n2242_));
  NOR2X1   g2193(.A(new_n1902_), .B(new_n1703_), .Y(new_n2243_));
  AOI21X1  g2194(.A0(new_n2003_), .A1(new_n1903_), .B0(new_n2243_), .Y(new_n2244_));
  AOI22X1  g2195(.A0(new_n1699_), .A1(new_n1676_), .B0(new_n1693_), .B1(new_n1695_), .Y(new_n2245_));
  OAI21X1  g2196(.A0(new_n2045_), .A1(new_n1906_), .B0(new_n2245_), .Y(new_n2246_));
  AOI21X1  g2197(.A0(new_n2075_), .A1(new_n245_), .B0(new_n2246_), .Y(new_n2247_));
  XOR2X1   g2198(.A(new_n2247_), .B(new_n230_), .Y(new_n2248_));
  AND2X1   g2199(.A(new_n1899_), .B(new_n1893_), .Y(new_n2249_));
  AOI21X1  g2200(.A0(new_n1900_), .A1(new_n1871_), .B0(new_n2249_), .Y(new_n2250_));
  INVX1    g2201(.A(new_n1876_), .Y(new_n2251_));
  OR2X1    g2202(.A(new_n1892_), .B(new_n1890_), .Y(new_n2252_));
  OAI21X1  g2203(.A0(new_n1889_), .A1(new_n2251_), .B0(new_n2252_), .Y(new_n2253_));
  AOI22X1  g2204(.A0(new_n1729_), .A1(new_n1620_), .B0(new_n1727_), .B1(new_n1623_), .Y(new_n2254_));
  OAI21X1  g2205(.A0(new_n1750_), .A1(new_n1815_), .B0(new_n2254_), .Y(new_n2255_));
  AOI21X1  g2206(.A0(new_n1814_), .A1(new_n1721_), .B0(new_n2255_), .Y(new_n2256_));
  XOR2X1   g2207(.A(new_n2256_), .B(new_n313_), .Y(new_n2257_));
  INVX1    g2208(.A(new_n1888_), .Y(new_n2258_));
  AOI21X1  g2209(.A0(new_n1649_), .A1(new_n1648_), .B0(new_n793_), .Y(new_n2259_));
  AOI22X1  g2210(.A0(new_n1877_), .A1(new_n1644_), .B0(new_n1710_), .B1(new_n1642_), .Y(new_n2260_));
  OAI21X1  g2211(.A0(new_n1714_), .A1(new_n1638_), .B0(new_n2260_), .Y(new_n2261_));
  AOI21X1  g2212(.A0(new_n2116_), .A1(new_n1707_), .B0(new_n2261_), .Y(new_n2262_));
  NAND3X1  g2213(.A(new_n2262_), .B(new_n1734_), .C(new_n525_), .Y(new_n2263_));
  XOR2X1   g2214(.A(new_n2262_), .B(new_n793_), .Y(new_n2264_));
  OAI21X1  g2215(.A0(new_n2264_), .A1(new_n2259_), .B0(new_n2263_), .Y(new_n2265_));
  XOR2X1   g2216(.A(new_n2265_), .B(new_n2258_), .Y(new_n2266_));
  XOR2X1   g2217(.A(new_n2266_), .B(new_n2257_), .Y(new_n2267_));
  XOR2X1   g2218(.A(new_n2267_), .B(new_n2253_), .Y(new_n2268_));
  INVX1    g2219(.A(new_n2268_), .Y(new_n2269_));
  OAI22X1  g2220(.A0(new_n1805_), .A1(new_n1797_), .B0(new_n1802_), .B1(new_n1585_), .Y(new_n2270_));
  AOI21X1  g2221(.A0(new_n1796_), .A1(new_n1613_), .B0(new_n2270_), .Y(new_n2271_));
  OAI21X1  g2222(.A0(new_n1919_), .A1(new_n1810_), .B0(new_n2271_), .Y(new_n2272_));
  XOR2X1   g2223(.A(new_n2272_), .B(new_n1164_), .Y(new_n2273_));
  XOR2X1   g2224(.A(new_n2273_), .B(new_n2269_), .Y(new_n2274_));
  XOR2X1   g2225(.A(new_n2274_), .B(new_n2250_), .Y(new_n2275_));
  XOR2X1   g2226(.A(new_n2275_), .B(new_n2248_), .Y(new_n2276_));
  XOR2X1   g2227(.A(new_n2276_), .B(new_n2244_), .Y(new_n2277_));
  INVX1    g2228(.A(new_n380_), .Y(new_n2278_));
  OR4X1    g2229(.A(new_n2278_), .B(new_n360_), .C(new_n356_), .D(new_n324_), .Y(new_n2279_));
  OR2X1    g2230(.A(new_n252_), .B(new_n183_), .Y(new_n2280_));
  OR2X1    g2231(.A(new_n2280_), .B(new_n365_), .Y(new_n2281_));
  OR4X1    g2232(.A(new_n391_), .B(new_n173_), .C(new_n121_), .D(new_n97_), .Y(new_n2282_));
  NOR3X1   g2233(.A(new_n2282_), .B(new_n2281_), .C(new_n2279_), .Y(new_n2283_));
  INVX1    g2234(.A(new_n2283_), .Y(new_n2284_));
  AND2X1   g2235(.A(new_n2038_), .B(new_n2031_), .Y(new_n2285_));
  XOR2X1   g2236(.A(new_n2285_), .B(new_n2284_), .Y(new_n2286_));
  OAI22X1  g2237(.A0(new_n2049_), .A1(new_n2039_), .B0(new_n2047_), .B1(new_n2042_), .Y(new_n2287_));
  AOI21X1  g2238(.A0(new_n2286_), .A1(new_n2010_), .B0(new_n2287_), .Y(new_n2288_));
  NOR2X1   g2239(.A(new_n2047_), .B(new_n2039_), .Y(new_n2289_));
  AOI21X1  g2240(.A0(new_n2061_), .A1(new_n2060_), .B0(new_n2289_), .Y(new_n2290_));
  XOR2X1   g2241(.A(new_n2286_), .B(new_n2040_), .Y(new_n2291_));
  XOR2X1   g2242(.A(new_n2291_), .B(new_n2290_), .Y(new_n2292_));
  OAI21X1  g2243(.A0(new_n2292_), .A1(new_n2009_), .B0(new_n2288_), .Y(new_n2293_));
  XOR2X1   g2244(.A(new_n2293_), .B(new_n243_), .Y(new_n2294_));
  XOR2X1   g2245(.A(new_n2294_), .B(new_n2277_), .Y(new_n2295_));
  OAI21X1  g2246(.A0(new_n2242_), .A1(new_n2066_), .B0(new_n2295_), .Y(new_n2296_));
  NAND2X1  g2247(.A(new_n2065_), .B(new_n2004_), .Y(new_n2297_));
  AND2X1   g2248(.A(new_n2073_), .B(new_n2067_), .Y(new_n2298_));
  XOR2X1   g2249(.A(new_n2079_), .B(new_n2081_), .Y(new_n2299_));
  XOR2X1   g2250(.A(new_n2211_), .B(new_n243_), .Y(new_n2300_));
  OAI21X1  g2251(.A0(new_n2223_), .A1(new_n2222_), .B0(new_n2300_), .Y(new_n2301_));
  NAND2X1  g2252(.A(new_n2223_), .B(new_n2222_), .Y(new_n2302_));
  INVX1    g2253(.A(new_n2226_), .Y(new_n2303_));
  AOI21X1  g2254(.A0(new_n2302_), .A1(new_n2301_), .B0(new_n2303_), .Y(new_n2304_));
  XOR2X1   g2255(.A(new_n2230_), .B(new_n243_), .Y(new_n2305_));
  NAND3X1  g2256(.A(new_n2303_), .B(new_n2302_), .C(new_n2301_), .Y(new_n2306_));
  OAI21X1  g2257(.A0(new_n2305_), .A1(new_n2304_), .B0(new_n2306_), .Y(new_n2307_));
  OAI21X1  g2258(.A0(new_n2307_), .A1(new_n2299_), .B0(new_n2234_), .Y(new_n2308_));
  OR2X1    g2259(.A(new_n2233_), .B(new_n2080_), .Y(new_n2309_));
  XOR2X1   g2260(.A(new_n2072_), .B(new_n2081_), .Y(new_n2310_));
  XOR2X1   g2261(.A(new_n2310_), .B(new_n2067_), .Y(new_n2311_));
  AOI21X1  g2262(.A0(new_n2309_), .A1(new_n2308_), .B0(new_n2311_), .Y(new_n2312_));
  XOR2X1   g2263(.A(new_n2065_), .B(new_n2004_), .Y(new_n2313_));
  OAI21X1  g2264(.A0(new_n2312_), .A1(new_n2298_), .B0(new_n2313_), .Y(new_n2314_));
  XOR2X1   g2265(.A(new_n2293_), .B(new_n2081_), .Y(new_n2315_));
  XOR2X1   g2266(.A(new_n2315_), .B(new_n2277_), .Y(new_n2316_));
  NAND3X1  g2267(.A(new_n2316_), .B(new_n2314_), .C(new_n2297_), .Y(new_n2317_));
  NAND3X1  g2268(.A(new_n2317_), .B(new_n2296_), .C(new_n225_), .Y(new_n2318_));
  OR4X1    g2269(.A(new_n347_), .B(new_n208_), .C(new_n132_), .D(new_n130_), .Y(new_n2319_));
  OR4X1    g2270(.A(new_n1418_), .B(new_n322_), .C(new_n255_), .D(new_n253_), .Y(new_n2320_));
  OR4X1    g2271(.A(new_n2320_), .B(new_n2319_), .C(new_n729_), .D(new_n529_), .Y(new_n2321_));
  NOR4X1   g2272(.A(new_n2321_), .B(new_n553_), .C(new_n292_), .D(new_n261_), .Y(new_n2322_));
  OR2X1    g2273(.A(new_n204_), .B(new_n179_), .Y(new_n2323_));
  OR4X1    g2274(.A(new_n2323_), .B(new_n325_), .C(new_n293_), .D(new_n283_), .Y(new_n2324_));
  OR4X1    g2275(.A(new_n388_), .B(new_n305_), .C(new_n184_), .D(new_n172_), .Y(new_n2325_));
  OR4X1    g2276(.A(new_n202_), .B(new_n198_), .C(new_n195_), .D(new_n192_), .Y(new_n2326_));
  OR4X1    g2277(.A(new_n2326_), .B(new_n2325_), .C(new_n2324_), .D(new_n1460_), .Y(new_n2327_));
  OR4X1    g2278(.A(new_n280_), .B(new_n264_), .C(new_n256_), .D(new_n207_), .Y(new_n2328_));
  OR4X1    g2279(.A(new_n2328_), .B(new_n260_), .C(new_n190_), .D(new_n182_), .Y(new_n2329_));
  OR4X1    g2280(.A(new_n2329_), .B(new_n314_), .C(new_n287_), .D(new_n251_), .Y(new_n2330_));
  NOR4X1   g2281(.A(new_n2330_), .B(new_n2327_), .C(new_n1473_), .D(new_n1469_), .Y(new_n2331_));
  AND2X1   g2282(.A(new_n2331_), .B(new_n2322_), .Y(new_n2332_));
  NAND3X1  g2283(.A(new_n2241_), .B(new_n2239_), .C(new_n2074_), .Y(new_n2333_));
  NOR3X1   g2284(.A(new_n2238_), .B(new_n2237_), .C(new_n2236_), .Y(new_n2334_));
  NOR3X1   g2285(.A(new_n1594_), .B(new_n190_), .C(new_n180_), .Y(new_n2335_));
  NAND2X1  g2286(.A(new_n2335_), .B(new_n548_), .Y(new_n2336_));
  OR4X1    g2287(.A(new_n315_), .B(new_n269_), .C(new_n249_), .D(new_n193_), .Y(new_n2337_));
  NOR3X1   g2288(.A(new_n2337_), .B(new_n1379_), .C(new_n2032_), .Y(new_n2338_));
  AND2X1   g2289(.A(new_n2338_), .B(new_n1396_), .Y(new_n2339_));
  NOR4X1   g2290(.A(new_n1461_), .B(new_n1457_), .C(new_n603_), .D(new_n331_), .Y(new_n2340_));
  OR4X1    g2291(.A(new_n184_), .B(new_n163_), .C(new_n134_), .D(new_n121_), .Y(new_n2341_));
  NOR4X1   g2292(.A(new_n2341_), .B(new_n357_), .C(new_n397_), .D(new_n272_), .Y(new_n2342_));
  NAND4X1  g2293(.A(new_n2342_), .B(new_n2340_), .C(new_n2339_), .D(new_n1430_), .Y(new_n2343_));
  NOR2X1   g2294(.A(new_n2343_), .B(new_n2336_), .Y(new_n2344_));
  NOR3X1   g2295(.A(new_n2344_), .B(new_n2334_), .C(new_n2312_), .Y(new_n2345_));
  AOI21X1  g2296(.A0(new_n2333_), .A1(new_n2314_), .B0(new_n2345_), .Y(new_n2346_));
  NAND3X1  g2297(.A(new_n2345_), .B(new_n2333_), .C(new_n2314_), .Y(new_n2347_));
  OAI21X1  g2298(.A0(new_n2346_), .A1(new_n2332_), .B0(new_n2347_), .Y(new_n2348_));
  AOI21X1  g2299(.A0(new_n2317_), .A1(new_n2296_), .B0(new_n224_), .Y(new_n2349_));
  AOI21X1  g2300(.A0(new_n2314_), .A1(new_n2297_), .B0(new_n2316_), .Y(new_n2350_));
  NOR3X1   g2301(.A(new_n2295_), .B(new_n2242_), .C(new_n2066_), .Y(new_n2351_));
  NOR3X1   g2302(.A(new_n2351_), .B(new_n2350_), .C(new_n225_), .Y(new_n2352_));
  OAI21X1  g2303(.A0(new_n2352_), .A1(new_n2349_), .B0(new_n2348_), .Y(new_n2353_));
  AND2X1   g2304(.A(new_n2353_), .B(new_n2318_), .Y(new_n2354_));
  NAND2X1  g2305(.A(new_n2286_), .B(new_n2040_), .Y(new_n2355_));
  INVX1    g2306(.A(new_n2291_), .Y(new_n2356_));
  OAI21X1  g2307(.A0(new_n2356_), .A1(new_n2290_), .B0(new_n2355_), .Y(new_n2357_));
  NAND3X1  g2308(.A(new_n2283_), .B(new_n2038_), .C(new_n2031_), .Y(new_n2358_));
  OR4X1    g2309(.A(new_n388_), .B(new_n347_), .C(new_n303_), .D(new_n265_), .Y(new_n2359_));
  OAI21X1  g2310(.A0(new_n333_), .A1(new_n70_), .B0(new_n215_), .Y(new_n2360_));
  OR4X1    g2311(.A(new_n2360_), .B(new_n2359_), .C(new_n574_), .D(new_n142_), .Y(new_n2361_));
  OR4X1    g2312(.A(new_n145_), .B(new_n134_), .C(new_n127_), .D(new_n91_), .Y(new_n2362_));
  OR4X1    g2313(.A(new_n605_), .B(new_n255_), .C(new_n197_), .D(new_n167_), .Y(new_n2363_));
  NOR3X1   g2314(.A(new_n348_), .B(new_n294_), .C(new_n397_), .Y(new_n2364_));
  NAND2X1  g2315(.A(new_n2364_), .B(new_n578_), .Y(new_n2365_));
  OR4X1    g2316(.A(new_n2365_), .B(new_n2363_), .C(new_n2362_), .D(new_n1591_), .Y(new_n2366_));
  NOR3X1   g2317(.A(new_n2366_), .B(new_n2361_), .C(new_n722_), .Y(new_n2367_));
  XOR2X1   g2318(.A(new_n2367_), .B(new_n2358_), .Y(new_n2368_));
  XOR2X1   g2319(.A(new_n2368_), .B(new_n2286_), .Y(new_n2369_));
  XOR2X1   g2320(.A(new_n2369_), .B(new_n2357_), .Y(new_n2370_));
  INVX1    g2321(.A(new_n2368_), .Y(new_n2371_));
  AOI22X1  g2322(.A0(new_n2286_), .A1(new_n2048_), .B0(new_n2041_), .B1(new_n2040_), .Y(new_n2372_));
  OAI21X1  g2323(.A0(new_n2371_), .A1(new_n2076_), .B0(new_n2372_), .Y(new_n2373_));
  AOI21X1  g2324(.A0(new_n2370_), .A1(new_n2008_), .B0(new_n2373_), .Y(new_n2374_));
  XOR2X1   g2325(.A(new_n2374_), .B(new_n243_), .Y(new_n2375_));
  XOR2X1   g2326(.A(new_n2247_), .B(new_n229_), .Y(new_n2376_));
  NAND2X1  g2327(.A(new_n2275_), .B(new_n2376_), .Y(new_n2377_));
  OAI21X1  g2328(.A0(new_n2276_), .A1(new_n2244_), .B0(new_n2377_), .Y(new_n2378_));
  AOI22X1  g2329(.A0(new_n1804_), .A1(new_n1613_), .B0(new_n1796_), .B1(new_n1584_), .Y(new_n2379_));
  OAI21X1  g2330(.A0(new_n1802_), .A1(new_n1673_), .B0(new_n2379_), .Y(new_n2380_));
  AOI21X1  g2331(.A0(new_n1905_), .A1(new_n1809_), .B0(new_n2380_), .Y(new_n2381_));
  XOR2X1   g2332(.A(new_n2381_), .B(new_n519_), .Y(new_n2382_));
  NOR2X1   g2333(.A(new_n2266_), .B(new_n2257_), .Y(new_n2383_));
  AOI21X1  g2334(.A0(new_n2267_), .A1(new_n2253_), .B0(new_n2383_), .Y(new_n2384_));
  OAI21X1  g2335(.A0(new_n2265_), .A1(new_n1888_), .B0(new_n2263_), .Y(new_n2385_));
  AOI22X1  g2336(.A0(new_n1877_), .A1(new_n1642_), .B0(new_n1710_), .B1(new_n1657_), .Y(new_n2386_));
  OAI21X1  g2337(.A0(new_n1714_), .A1(new_n1778_), .B0(new_n2386_), .Y(new_n2387_));
  AOI21X1  g2338(.A0(new_n1777_), .A1(new_n1707_), .B0(new_n2387_), .Y(new_n2388_));
  OR2X1    g2339(.A(new_n1644_), .B(new_n793_), .Y(new_n2389_));
  XOR2X1   g2340(.A(new_n2389_), .B(new_n2388_), .Y(new_n2390_));
  XOR2X1   g2341(.A(new_n2390_), .B(new_n2385_), .Y(new_n2391_));
  OAI22X1  g2342(.A0(new_n1728_), .A1(new_n1798_), .B0(new_n1750_), .B1(new_n1797_), .Y(new_n2392_));
  AOI21X1  g2343(.A0(new_n1729_), .A1(new_n1618_), .B0(new_n2392_), .Y(new_n2393_));
  OAI21X1  g2344(.A0(new_n1808_), .A1(new_n1722_), .B0(new_n2393_), .Y(new_n2394_));
  XOR2X1   g2345(.A(new_n2394_), .B(new_n313_), .Y(new_n2395_));
  XOR2X1   g2346(.A(new_n2395_), .B(new_n2391_), .Y(new_n2396_));
  XOR2X1   g2347(.A(new_n2396_), .B(new_n2384_), .Y(new_n2397_));
  XOR2X1   g2348(.A(new_n2397_), .B(new_n2382_), .Y(new_n2398_));
  NOR2X1   g2349(.A(new_n2274_), .B(new_n2250_), .Y(new_n2399_));
  AOI21X1  g2350(.A0(new_n2273_), .A1(new_n2268_), .B0(new_n2399_), .Y(new_n2400_));
  XOR2X1   g2351(.A(new_n2400_), .B(new_n2398_), .Y(new_n2401_));
  INVX1    g2352(.A(new_n2401_), .Y(new_n2402_));
  OAI22X1  g2353(.A0(new_n2045_), .A1(new_n1694_), .B0(new_n1916_), .B1(new_n1688_), .Y(new_n2403_));
  AOI21X1  g2354(.A0(new_n2052_), .A1(new_n1696_), .B0(new_n2403_), .Y(new_n2404_));
  OAI21X1  g2355(.A0(new_n2071_), .A1(new_n1915_), .B0(new_n2404_), .Y(new_n2405_));
  XOR2X1   g2356(.A(new_n2405_), .B(new_n230_), .Y(new_n2406_));
  XOR2X1   g2357(.A(new_n2406_), .B(new_n2402_), .Y(new_n2407_));
  XOR2X1   g2358(.A(new_n2407_), .B(new_n2378_), .Y(new_n2408_));
  XOR2X1   g2359(.A(new_n2408_), .B(new_n2375_), .Y(new_n2409_));
  NAND2X1  g2360(.A(new_n2294_), .B(new_n2277_), .Y(new_n2410_));
  AND2X1   g2361(.A(new_n2296_), .B(new_n2410_), .Y(new_n2411_));
  XOR2X1   g2362(.A(new_n2411_), .B(new_n2409_), .Y(new_n2412_));
  INVX1    g2363(.A(new_n213_), .Y(new_n2413_));
  NAND4X1  g2364(.A(new_n257_), .B(new_n215_), .C(new_n544_), .D(new_n2413_), .Y(new_n2414_));
  OR2X1    g2365(.A(new_n208_), .B(new_n183_), .Y(new_n2415_));
  OR4X1    g2366(.A(new_n2415_), .B(new_n1460_), .C(new_n446_), .D(new_n142_), .Y(new_n2416_));
  OR4X1    g2367(.A(new_n2416_), .B(new_n2414_), .C(new_n1380_), .D(new_n615_), .Y(new_n2417_));
  NOR4X1   g2368(.A(new_n2417_), .B(new_n1391_), .C(new_n532_), .D(new_n500_), .Y(new_n2418_));
  XOR2X1   g2369(.A(new_n2418_), .B(new_n2412_), .Y(new_n2419_));
  XOR2X1   g2370(.A(new_n2419_), .B(new_n2354_), .Y(new_n2420_));
  NOR2X1   g2371(.A(new_n2352_), .B(new_n2349_), .Y(new_n2421_));
  XOR2X1   g2372(.A(new_n2421_), .B(new_n2348_), .Y(new_n2422_));
  XOR2X1   g2373(.A(new_n2422_), .B(new_n2420_), .Y(\sin[0] ));
  NOR2X1   g2374(.A(new_n2422_), .B(new_n2420_), .Y(new_n2424_));
  AND2X1   g2375(.A(new_n2418_), .B(new_n2412_), .Y(new_n2425_));
  OR2X1    g2376(.A(new_n2418_), .B(new_n2412_), .Y(new_n2426_));
  OAI21X1  g2377(.A0(new_n2425_), .A1(new_n2354_), .B0(new_n2426_), .Y(new_n2427_));
  AND2X1   g2378(.A(new_n2368_), .B(new_n2286_), .Y(new_n2428_));
  AOI21X1  g2379(.A0(new_n2369_), .A1(new_n2357_), .B0(new_n2428_), .Y(new_n2429_));
  NAND4X1  g2380(.A(new_n2367_), .B(new_n2283_), .C(new_n2038_), .D(new_n2031_), .Y(new_n2430_));
  OR4X1    g2381(.A(new_n205_), .B(new_n174_), .C(new_n170_), .D(new_n169_), .Y(new_n2431_));
  OR4X1    g2382(.A(new_n2431_), .B(new_n1461_), .C(new_n420_), .D(new_n138_), .Y(new_n2432_));
  OR4X1    g2383(.A(new_n527_), .B(new_n321_), .C(new_n287_), .D(new_n253_), .Y(new_n2433_));
  NOR4X1   g2384(.A(new_n2433_), .B(new_n568_), .C(new_n497_), .D(new_n452_), .Y(new_n2434_));
  NAND4X1  g2385(.A(new_n2434_), .B(new_n548_), .C(new_n339_), .D(new_n544_), .Y(new_n2435_));
  OR4X1    g2386(.A(new_n2435_), .B(new_n2432_), .C(new_n926_), .D(new_n344_), .Y(new_n2436_));
  NOR2X1   g2387(.A(new_n2436_), .B(new_n1459_), .Y(new_n2437_));
  XOR2X1   g2388(.A(new_n2437_), .B(new_n2430_), .Y(new_n2438_));
  XOR2X1   g2389(.A(new_n2438_), .B(new_n2368_), .Y(new_n2439_));
  INVX1    g2390(.A(new_n2439_), .Y(new_n2440_));
  XOR2X1   g2391(.A(new_n2440_), .B(new_n2429_), .Y(new_n2441_));
  INVX1    g2392(.A(new_n2438_), .Y(new_n2442_));
  AOI22X1  g2393(.A0(new_n2368_), .A1(new_n2048_), .B0(new_n2286_), .B1(new_n2041_), .Y(new_n2443_));
  OAI21X1  g2394(.A0(new_n2442_), .A1(new_n2076_), .B0(new_n2443_), .Y(new_n2444_));
  AOI21X1  g2395(.A0(new_n2441_), .A1(new_n2008_), .B0(new_n2444_), .Y(new_n2445_));
  XOR2X1   g2396(.A(new_n2445_), .B(new_n243_), .Y(new_n2446_));
  NAND2X1  g2397(.A(new_n2406_), .B(new_n2401_), .Y(new_n2447_));
  XOR2X1   g2398(.A(new_n2406_), .B(new_n2401_), .Y(new_n2448_));
  NAND2X1  g2399(.A(new_n2448_), .B(new_n2378_), .Y(new_n2449_));
  NAND2X1  g2400(.A(new_n2449_), .B(new_n2447_), .Y(new_n2450_));
  AOI22X1  g2401(.A0(new_n1804_), .A1(new_n1584_), .B0(new_n1801_), .B1(new_n1695_), .Y(new_n2451_));
  OAI21X1  g2402(.A0(new_n1824_), .A1(new_n1673_), .B0(new_n2451_), .Y(new_n2452_));
  AOI21X1  g2403(.A0(new_n1809_), .A1(new_n1690_), .B0(new_n2452_), .Y(new_n2453_));
  XOR2X1   g2404(.A(new_n2453_), .B(new_n519_), .Y(new_n2454_));
  AND2X1   g2405(.A(new_n2395_), .B(new_n2391_), .Y(new_n2455_));
  INVX1    g2406(.A(new_n2455_), .Y(new_n2456_));
  INVX1    g2407(.A(new_n2396_), .Y(new_n2457_));
  OAI21X1  g2408(.A0(new_n2457_), .A1(new_n2384_), .B0(new_n2456_), .Y(new_n2458_));
  NAND2X1  g2409(.A(new_n2390_), .B(new_n2385_), .Y(new_n2459_));
  NAND3X1  g2410(.A(new_n2388_), .B(new_n1644_), .C(new_n525_), .Y(new_n2460_));
  NAND2X1  g2411(.A(new_n2460_), .B(new_n2459_), .Y(new_n2461_));
  OAI22X1  g2412(.A0(new_n1785_), .A1(new_n1638_), .B0(new_n1711_), .B1(new_n1778_), .Y(new_n2462_));
  AOI21X1  g2413(.A0(new_n1713_), .A1(new_n1620_), .B0(new_n2462_), .Y(new_n2463_));
  OAI21X1  g2414(.A0(new_n1827_), .A1(new_n1784_), .B0(new_n2463_), .Y(new_n2464_));
  AND2X1   g2415(.A(new_n1640_), .B(new_n525_), .Y(new_n2465_));
  XOR2X1   g2416(.A(new_n2465_), .B(new_n2464_), .Y(new_n2466_));
  XOR2X1   g2417(.A(new_n2466_), .B(new_n2461_), .Y(new_n2467_));
  OAI22X1  g2418(.A0(new_n1730_), .A1(new_n1797_), .B0(new_n1728_), .B1(new_n1815_), .Y(new_n2468_));
  AOI21X1  g2419(.A0(new_n1724_), .A1(new_n1613_), .B0(new_n2468_), .Y(new_n2469_));
  OAI21X1  g2420(.A0(new_n1895_), .A1(new_n1722_), .B0(new_n2469_), .Y(new_n2470_));
  XOR2X1   g2421(.A(new_n2470_), .B(new_n313_), .Y(new_n2471_));
  XOR2X1   g2422(.A(new_n2471_), .B(new_n2467_), .Y(new_n2472_));
  INVX1    g2423(.A(new_n2472_), .Y(new_n2473_));
  XOR2X1   g2424(.A(new_n2473_), .B(new_n2458_), .Y(new_n2474_));
  XOR2X1   g2425(.A(new_n2474_), .B(new_n2454_), .Y(new_n2475_));
  XOR2X1   g2426(.A(new_n2381_), .B(new_n1164_), .Y(new_n2476_));
  OR2X1    g2427(.A(new_n2397_), .B(new_n2476_), .Y(new_n2477_));
  OAI21X1  g2428(.A0(new_n2400_), .A1(new_n2398_), .B0(new_n2477_), .Y(new_n2478_));
  XOR2X1   g2429(.A(new_n2478_), .B(new_n2475_), .Y(new_n2479_));
  OAI22X1  g2430(.A0(new_n2047_), .A1(new_n1694_), .B0(new_n2045_), .B1(new_n1916_), .Y(new_n2480_));
  AOI21X1  g2431(.A0(new_n2040_), .A1(new_n1696_), .B0(new_n2480_), .Y(new_n2481_));
  OAI21X1  g2432(.A0(new_n2063_), .A1(new_n1915_), .B0(new_n2481_), .Y(new_n2482_));
  XOR2X1   g2433(.A(new_n2482_), .B(new_n230_), .Y(new_n2483_));
  XOR2X1   g2434(.A(new_n2483_), .B(new_n2479_), .Y(new_n2484_));
  XOR2X1   g2435(.A(new_n2484_), .B(new_n2450_), .Y(new_n2485_));
  XOR2X1   g2436(.A(new_n2485_), .B(new_n2446_), .Y(new_n2486_));
  OR2X1    g2437(.A(new_n2408_), .B(new_n2375_), .Y(new_n2487_));
  AND2X1   g2438(.A(new_n2294_), .B(new_n2277_), .Y(new_n2488_));
  OAI21X1  g2439(.A0(new_n2350_), .A1(new_n2488_), .B0(new_n2409_), .Y(new_n2489_));
  AND2X1   g2440(.A(new_n2489_), .B(new_n2487_), .Y(new_n2490_));
  XOR2X1   g2441(.A(new_n2490_), .B(new_n2486_), .Y(new_n2491_));
  OR2X1    g2442(.A(new_n188_), .B(new_n182_), .Y(new_n2492_));
  OR2X1    g2443(.A(new_n205_), .B(new_n180_), .Y(new_n2493_));
  OR4X1    g2444(.A(new_n2493_), .B(new_n2492_), .C(new_n420_), .D(new_n273_), .Y(new_n2494_));
  NOR4X1   g2445(.A(new_n527_), .B(new_n551_), .C(new_n437_), .D(new_n193_), .Y(new_n2495_));
  NOR4X1   g2446(.A(new_n347_), .B(new_n264_), .C(new_n164_), .D(new_n155_), .Y(new_n2496_));
  NOR4X1   g2447(.A(new_n379_), .B(new_n616_), .C(new_n211_), .D(new_n196_), .Y(new_n2497_));
  NAND4X1  g2448(.A(new_n2497_), .B(new_n2496_), .C(new_n2495_), .D(new_n217_), .Y(new_n2498_));
  NOR4X1   g2449(.A(new_n2498_), .B(new_n2494_), .C(new_n1373_), .D(new_n144_), .Y(new_n2499_));
  XOR2X1   g2450(.A(new_n2499_), .B(new_n2491_), .Y(new_n2500_));
  XOR2X1   g2451(.A(new_n2500_), .B(new_n2427_), .Y(new_n2501_));
  XOR2X1   g2452(.A(new_n2501_), .B(new_n2424_), .Y(new_n2502_));
  XOR2X1   g2453(.A(\a[23] ), .B(new_n50_), .Y(new_n2503_));
  INVX1    g2454(.A(new_n2503_), .Y(new_n2504_));
  AND2X1   g2455(.A(new_n2504_), .B(\sin[0] ), .Y(new_n2505_));
  XOR2X1   g2456(.A(new_n2505_), .B(new_n2502_), .Y(\sin[1] ));
  NAND2X1  g2457(.A(new_n2501_), .B(new_n2424_), .Y(new_n2507_));
  NAND2X1  g2458(.A(new_n2353_), .B(new_n2318_), .Y(new_n2508_));
  NOR2X1   g2459(.A(new_n2418_), .B(new_n2412_), .Y(new_n2509_));
  AOI21X1  g2460(.A0(new_n2419_), .A1(new_n2508_), .B0(new_n2509_), .Y(new_n2510_));
  AND2X1   g2461(.A(new_n2499_), .B(new_n2491_), .Y(new_n2511_));
  OR2X1    g2462(.A(new_n2499_), .B(new_n2491_), .Y(new_n2512_));
  OAI21X1  g2463(.A0(new_n2511_), .A1(new_n2510_), .B0(new_n2512_), .Y(new_n2513_));
  OR4X1    g2464(.A(new_n446_), .B(new_n219_), .C(new_n197_), .D(new_n184_), .Y(new_n2514_));
  OR4X1    g2465(.A(new_n2514_), .B(new_n259_), .C(new_n192_), .D(new_n116_), .Y(new_n2515_));
  OR4X1    g2466(.A(new_n527_), .B(new_n388_), .C(new_n292_), .D(new_n182_), .Y(new_n2516_));
  OR4X1    g2467(.A(new_n608_), .B(new_n358_), .C(new_n293_), .D(new_n279_), .Y(new_n2517_));
  OR4X1    g2468(.A(new_n2517_), .B(new_n2516_), .C(new_n272_), .D(new_n208_), .Y(new_n2518_));
  NOR3X1   g2469(.A(new_n2518_), .B(new_n2515_), .C(new_n543_), .Y(new_n2519_));
  AND2X1   g2470(.A(new_n2519_), .B(new_n2339_), .Y(new_n2520_));
  INVX1    g2471(.A(new_n2520_), .Y(new_n2521_));
  NOR2X1   g2472(.A(new_n2485_), .B(new_n2446_), .Y(new_n2522_));
  XOR2X1   g2473(.A(new_n2445_), .B(new_n2081_), .Y(new_n2523_));
  XOR2X1   g2474(.A(new_n2485_), .B(new_n2523_), .Y(new_n2524_));
  AOI21X1  g2475(.A0(new_n2489_), .A1(new_n2487_), .B0(new_n2524_), .Y(new_n2525_));
  OR2X1    g2476(.A(new_n2525_), .B(new_n2522_), .Y(new_n2526_));
  AND2X1   g2477(.A(new_n2369_), .B(new_n2357_), .Y(new_n2527_));
  OAI21X1  g2478(.A0(new_n2527_), .A1(new_n2428_), .B0(new_n2439_), .Y(new_n2528_));
  AOI21X1  g2479(.A0(new_n2429_), .A1(new_n2371_), .B0(new_n2442_), .Y(new_n2529_));
  AOI21X1  g2480(.A0(new_n2528_), .A1(new_n2442_), .B0(new_n2529_), .Y(new_n2530_));
  OAI22X1  g2481(.A0(new_n2442_), .A1(new_n2049_), .B0(new_n2371_), .B1(new_n2042_), .Y(new_n2531_));
  AOI21X1  g2482(.A0(new_n2530_), .A1(new_n2008_), .B0(new_n2531_), .Y(new_n2532_));
  XOR2X1   g2483(.A(new_n2532_), .B(new_n2081_), .Y(new_n2533_));
  INVX1    g2484(.A(new_n2479_), .Y(new_n2534_));
  AND2X1   g2485(.A(new_n2483_), .B(new_n2534_), .Y(new_n2535_));
  AOI21X1  g2486(.A0(new_n2449_), .A1(new_n2447_), .B0(new_n2484_), .Y(new_n2536_));
  NOR2X1   g2487(.A(new_n2536_), .B(new_n2535_), .Y(new_n2537_));
  AOI22X1  g2488(.A0(new_n1804_), .A1(new_n1676_), .B0(new_n1796_), .B1(new_n1695_), .Y(new_n2538_));
  OAI21X1  g2489(.A0(new_n2045_), .A1(new_n1802_), .B0(new_n2538_), .Y(new_n2539_));
  AOI21X1  g2490(.A0(new_n2075_), .A1(new_n1809_), .B0(new_n2539_), .Y(new_n2540_));
  XOR2X1   g2491(.A(new_n2540_), .B(new_n1164_), .Y(new_n2541_));
  AND2X1   g2492(.A(new_n2471_), .B(new_n2467_), .Y(new_n2542_));
  AOI21X1  g2493(.A0(new_n2472_), .A1(new_n2458_), .B0(new_n2542_), .Y(new_n2543_));
  NOR3X1   g2494(.A(new_n2464_), .B(new_n1640_), .C(new_n793_), .Y(new_n2544_));
  AOI21X1  g2495(.A0(new_n2466_), .A1(new_n2461_), .B0(new_n2544_), .Y(new_n2545_));
  AOI22X1  g2496(.A0(new_n1877_), .A1(new_n1623_), .B0(new_n1710_), .B1(new_n1620_), .Y(new_n2546_));
  OAI21X1  g2497(.A0(new_n1714_), .A1(new_n1815_), .B0(new_n2546_), .Y(new_n2547_));
  AOI21X1  g2498(.A0(new_n1814_), .A1(new_n1707_), .B0(new_n2547_), .Y(new_n2548_));
  AND2X1   g2499(.A(new_n1638_), .B(new_n525_), .Y(new_n2549_));
  XOR2X1   g2500(.A(new_n2549_), .B(new_n2548_), .Y(new_n2550_));
  INVX1    g2501(.A(new_n2550_), .Y(new_n2551_));
  XOR2X1   g2502(.A(new_n2551_), .B(new_n2545_), .Y(new_n2552_));
  OAI22X1  g2503(.A0(new_n1728_), .A1(new_n1797_), .B0(new_n1750_), .B1(new_n1585_), .Y(new_n2553_));
  AOI21X1  g2504(.A0(new_n1729_), .A1(new_n1613_), .B0(new_n2553_), .Y(new_n2554_));
  OAI21X1  g2505(.A0(new_n1919_), .A1(new_n1722_), .B0(new_n2554_), .Y(new_n2555_));
  XOR2X1   g2506(.A(new_n2555_), .B(new_n313_), .Y(new_n2556_));
  XOR2X1   g2507(.A(new_n2556_), .B(new_n2552_), .Y(new_n2557_));
  XOR2X1   g2508(.A(new_n2557_), .B(new_n2543_), .Y(new_n2558_));
  XOR2X1   g2509(.A(new_n2558_), .B(new_n2541_), .Y(new_n2559_));
  INVX1    g2510(.A(new_n2454_), .Y(new_n2560_));
  NOR2X1   g2511(.A(new_n2474_), .B(new_n2560_), .Y(new_n2561_));
  INVX1    g2512(.A(new_n2475_), .Y(new_n2562_));
  AOI21X1  g2513(.A0(new_n2478_), .A1(new_n2562_), .B0(new_n2561_), .Y(new_n2563_));
  XOR2X1   g2514(.A(new_n2563_), .B(new_n2559_), .Y(new_n2564_));
  OAI22X1  g2515(.A0(new_n2047_), .A1(new_n1916_), .B0(new_n2039_), .B1(new_n1694_), .Y(new_n2565_));
  AOI21X1  g2516(.A0(new_n2286_), .A1(new_n1696_), .B0(new_n2565_), .Y(new_n2566_));
  OAI21X1  g2517(.A0(new_n2292_), .A1(new_n1915_), .B0(new_n2566_), .Y(new_n2567_));
  XOR2X1   g2518(.A(new_n2567_), .B(new_n230_), .Y(new_n2568_));
  XOR2X1   g2519(.A(new_n2568_), .B(new_n2564_), .Y(new_n2569_));
  XOR2X1   g2520(.A(new_n2569_), .B(new_n2537_), .Y(new_n2570_));
  XOR2X1   g2521(.A(new_n2570_), .B(new_n2533_), .Y(new_n2571_));
  XOR2X1   g2522(.A(new_n2571_), .B(new_n2526_), .Y(new_n2572_));
  XOR2X1   g2523(.A(new_n2572_), .B(new_n2521_), .Y(new_n2573_));
  NAND2X1  g2524(.A(new_n2573_), .B(new_n2513_), .Y(new_n2574_));
  NOR2X1   g2525(.A(new_n2499_), .B(new_n2491_), .Y(new_n2575_));
  AOI21X1  g2526(.A0(new_n2500_), .A1(new_n2427_), .B0(new_n2575_), .Y(new_n2576_));
  OR2X1    g2527(.A(new_n2572_), .B(new_n2520_), .Y(new_n2577_));
  NAND2X1  g2528(.A(new_n2572_), .B(new_n2520_), .Y(new_n2578_));
  NAND3X1  g2529(.A(new_n2578_), .B(new_n2577_), .C(new_n2576_), .Y(new_n2579_));
  AND2X1   g2530(.A(new_n2579_), .B(new_n2574_), .Y(new_n2580_));
  XOR2X1   g2531(.A(new_n2580_), .B(new_n2507_), .Y(new_n2581_));
  OR2X1    g2532(.A(new_n2502_), .B(\sin[0] ), .Y(new_n2582_));
  AND2X1   g2533(.A(new_n2582_), .B(new_n2504_), .Y(new_n2583_));
  XOR2X1   g2534(.A(new_n2583_), .B(new_n2581_), .Y(\sin[2] ));
  AOI21X1  g2535(.A0(new_n2579_), .A1(new_n2574_), .B0(new_n2507_), .Y(new_n2585_));
  NOR2X1   g2536(.A(new_n2572_), .B(new_n2520_), .Y(new_n2586_));
  AOI21X1  g2537(.A0(new_n2578_), .A1(new_n2513_), .B0(new_n2586_), .Y(new_n2587_));
  NOR4X1   g2538(.A(new_n2324_), .B(new_n580_), .C(new_n447_), .D(new_n445_), .Y(new_n2588_));
  INVX1    g2539(.A(new_n478_), .Y(new_n2589_));
  OR4X1    g2540(.A(new_n2492_), .B(new_n2032_), .C(new_n203_), .D(new_n164_), .Y(new_n2590_));
  OR4X1    g2541(.A(new_n330_), .B(new_n397_), .C(new_n211_), .D(new_n141_), .Y(new_n2591_));
  NOR4X1   g2542(.A(new_n2591_), .B(new_n2590_), .C(new_n1376_), .D(new_n2589_), .Y(new_n2592_));
  NAND2X1  g2543(.A(new_n2592_), .B(new_n2588_), .Y(new_n2593_));
  NOR2X1   g2544(.A(new_n2593_), .B(new_n915_), .Y(new_n2594_));
  XOR2X1   g2545(.A(new_n2532_), .B(new_n243_), .Y(new_n2595_));
  OR2X1    g2546(.A(new_n2570_), .B(new_n2595_), .Y(new_n2596_));
  XOR2X1   g2547(.A(new_n2570_), .B(new_n2595_), .Y(new_n2597_));
  OAI21X1  g2548(.A0(new_n2525_), .A1(new_n2522_), .B0(new_n2597_), .Y(new_n2598_));
  AND2X1   g2549(.A(new_n2598_), .B(new_n2596_), .Y(new_n2599_));
  NAND2X1  g2550(.A(new_n2568_), .B(new_n2564_), .Y(new_n2600_));
  OAI21X1  g2551(.A0(new_n2536_), .A1(new_n2535_), .B0(new_n2569_), .Y(new_n2601_));
  AND2X1   g2552(.A(new_n2601_), .B(new_n2600_), .Y(new_n2602_));
  AOI22X1  g2553(.A0(new_n2529_), .A1(new_n2008_), .B0(new_n2438_), .B1(new_n2041_), .Y(new_n2603_));
  XOR2X1   g2554(.A(new_n2603_), .B(new_n2081_), .Y(new_n2604_));
  INVX1    g2555(.A(new_n2071_), .Y(new_n2605_));
  AOI22X1  g2556(.A0(new_n2044_), .A1(new_n1796_), .B0(new_n1804_), .B1(new_n1695_), .Y(new_n2606_));
  OAI21X1  g2557(.A0(new_n2047_), .A1(new_n1802_), .B0(new_n2606_), .Y(new_n2607_));
  AOI21X1  g2558(.A0(new_n2605_), .A1(new_n1809_), .B0(new_n2607_), .Y(new_n2608_));
  XOR2X1   g2559(.A(new_n2608_), .B(new_n1164_), .Y(new_n2609_));
  INVX1    g2560(.A(new_n2556_), .Y(new_n2610_));
  OR2X1    g2561(.A(new_n2610_), .B(new_n2552_), .Y(new_n2611_));
  OAI21X1  g2562(.A0(new_n2557_), .A1(new_n2543_), .B0(new_n2611_), .Y(new_n2612_));
  INVX1    g2563(.A(new_n2612_), .Y(new_n2613_));
  NAND3X1  g2564(.A(new_n2548_), .B(new_n1657_), .C(new_n525_), .Y(new_n2614_));
  OAI21X1  g2565(.A0(new_n2550_), .A1(new_n2545_), .B0(new_n2614_), .Y(new_n2615_));
  OAI22X1  g2566(.A0(new_n1785_), .A1(new_n1798_), .B0(new_n1714_), .B1(new_n1797_), .Y(new_n2616_));
  AOI21X1  g2567(.A0(new_n1710_), .A1(new_n1618_), .B0(new_n2616_), .Y(new_n2617_));
  OAI21X1  g2568(.A0(new_n1808_), .A1(new_n1784_), .B0(new_n2617_), .Y(new_n2618_));
  NOR2X1   g2569(.A(new_n1623_), .B(new_n793_), .Y(new_n2619_));
  XOR2X1   g2570(.A(new_n2619_), .B(new_n2618_), .Y(new_n2620_));
  XOR2X1   g2571(.A(new_n2620_), .B(new_n2615_), .Y(new_n2621_));
  INVX1    g2572(.A(new_n1905_), .Y(new_n2622_));
  OAI22X1  g2573(.A0(new_n1730_), .A1(new_n1585_), .B0(new_n1728_), .B1(new_n2198_), .Y(new_n2623_));
  AOI21X1  g2574(.A0(new_n1724_), .A1(new_n1676_), .B0(new_n2623_), .Y(new_n2624_));
  OAI21X1  g2575(.A0(new_n2622_), .A1(new_n1722_), .B0(new_n2624_), .Y(new_n2625_));
  XOR2X1   g2576(.A(new_n2625_), .B(new_n313_), .Y(new_n2626_));
  INVX1    g2577(.A(new_n2626_), .Y(new_n2627_));
  XOR2X1   g2578(.A(new_n2627_), .B(new_n2621_), .Y(new_n2628_));
  XOR2X1   g2579(.A(new_n2628_), .B(new_n2613_), .Y(new_n2629_));
  XOR2X1   g2580(.A(new_n2629_), .B(new_n2609_), .Y(new_n2630_));
  INVX1    g2581(.A(new_n2557_), .Y(new_n2631_));
  XOR2X1   g2582(.A(new_n2631_), .B(new_n2543_), .Y(new_n2632_));
  OR2X1    g2583(.A(new_n2632_), .B(new_n2541_), .Y(new_n2633_));
  OAI21X1  g2584(.A0(new_n2563_), .A1(new_n2559_), .B0(new_n2633_), .Y(new_n2634_));
  XOR2X1   g2585(.A(new_n2634_), .B(new_n2630_), .Y(new_n2635_));
  AOI22X1  g2586(.A0(new_n2286_), .A1(new_n1693_), .B0(new_n2040_), .B1(new_n1699_), .Y(new_n2636_));
  OAI21X1  g2587(.A0(new_n2371_), .A1(new_n1906_), .B0(new_n2636_), .Y(new_n2637_));
  AOI21X1  g2588(.A0(new_n2370_), .A1(new_n245_), .B0(new_n2637_), .Y(new_n2638_));
  XOR2X1   g2589(.A(new_n2638_), .B(new_n230_), .Y(new_n2639_));
  XOR2X1   g2590(.A(new_n2639_), .B(new_n2635_), .Y(new_n2640_));
  XOR2X1   g2591(.A(new_n2640_), .B(new_n2604_), .Y(new_n2641_));
  XOR2X1   g2592(.A(new_n2641_), .B(new_n2602_), .Y(new_n2642_));
  XOR2X1   g2593(.A(new_n2642_), .B(new_n2599_), .Y(new_n2643_));
  XOR2X1   g2594(.A(new_n2643_), .B(new_n2594_), .Y(new_n2644_));
  XOR2X1   g2595(.A(new_n2644_), .B(new_n2587_), .Y(new_n2645_));
  INVX1    g2596(.A(new_n2645_), .Y(new_n2646_));
  XOR2X1   g2597(.A(new_n2646_), .B(new_n2585_), .Y(new_n2647_));
  OAI21X1  g2598(.A0(new_n2582_), .A1(new_n2581_), .B0(new_n2504_), .Y(new_n2648_));
  XOR2X1   g2599(.A(new_n2648_), .B(new_n2647_), .Y(\sin[3] ));
  AND2X1   g2600(.A(new_n2645_), .B(new_n2585_), .Y(new_n2650_));
  INVX1    g2601(.A(new_n2594_), .Y(new_n2651_));
  NAND2X1  g2602(.A(new_n2643_), .B(new_n2651_), .Y(new_n2652_));
  OAI21X1  g2603(.A0(new_n2644_), .A1(new_n2587_), .B0(new_n2652_), .Y(new_n2653_));
  NOR2X1   g2604(.A(new_n168_), .B(new_n159_), .Y(new_n2654_));
  NOR4X1   g2605(.A(new_n446_), .B(new_n437_), .C(new_n184_), .D(new_n145_), .Y(new_n2655_));
  NAND3X1  g2606(.A(new_n2655_), .B(new_n2654_), .C(new_n465_), .Y(new_n2656_));
  OR4X1    g2607(.A(new_n2656_), .B(new_n1455_), .C(new_n618_), .D(new_n362_), .Y(new_n2657_));
  NOR3X1   g2608(.A(new_n2657_), .B(new_n507_), .C(new_n436_), .Y(new_n2658_));
  AND2X1   g2609(.A(new_n2658_), .B(new_n1476_), .Y(new_n2659_));
  NAND2X1  g2610(.A(new_n2601_), .B(new_n2600_), .Y(new_n2660_));
  AND2X1   g2611(.A(new_n2641_), .B(new_n2660_), .Y(new_n2661_));
  AOI21X1  g2612(.A0(new_n2598_), .A1(new_n2596_), .B0(new_n2642_), .Y(new_n2662_));
  OR2X1    g2613(.A(new_n2662_), .B(new_n2661_), .Y(new_n2663_));
  OR2X1    g2614(.A(new_n2639_), .B(new_n2635_), .Y(new_n2664_));
  NAND2X1  g2615(.A(new_n2640_), .B(new_n2604_), .Y(new_n2665_));
  NAND2X1  g2616(.A(new_n2665_), .B(new_n2664_), .Y(new_n2666_));
  XOR2X1   g2617(.A(new_n2628_), .B(new_n2612_), .Y(new_n2667_));
  NOR2X1   g2618(.A(new_n2667_), .B(new_n2609_), .Y(new_n2668_));
  OR2X1    g2619(.A(new_n2563_), .B(new_n2559_), .Y(new_n2669_));
  AOI21X1  g2620(.A0(new_n2669_), .A1(new_n2633_), .B0(new_n2630_), .Y(new_n2670_));
  OR2X1    g2621(.A(new_n2670_), .B(new_n2668_), .Y(new_n2671_));
  NAND2X1  g2622(.A(new_n2626_), .B(new_n2621_), .Y(new_n2672_));
  OAI21X1  g2623(.A0(new_n2628_), .A1(new_n2613_), .B0(new_n2672_), .Y(new_n2673_));
  AOI22X1  g2624(.A0(new_n1877_), .A1(new_n1618_), .B0(new_n1710_), .B1(new_n1615_), .Y(new_n2674_));
  OAI21X1  g2625(.A0(new_n1714_), .A1(new_n2198_), .B0(new_n2674_), .Y(new_n2675_));
  AOI21X1  g2626(.A0(new_n2180_), .A1(new_n1707_), .B0(new_n2675_), .Y(new_n2676_));
  XOR2X1   g2627(.A(new_n2676_), .B(new_n525_), .Y(new_n2677_));
  NAND3X1  g2628(.A(new_n1620_), .B(new_n525_), .C(new_n243_), .Y(new_n2678_));
  AND2X1   g2629(.A(new_n1620_), .B(new_n525_), .Y(new_n2679_));
  OAI21X1  g2630(.A0(new_n2679_), .A1(new_n243_), .B0(new_n2678_), .Y(new_n2680_));
  XOR2X1   g2631(.A(new_n2680_), .B(new_n2677_), .Y(new_n2681_));
  NOR3X1   g2632(.A(new_n2618_), .B(new_n1778_), .C(new_n793_), .Y(new_n2682_));
  AOI21X1  g2633(.A0(new_n2620_), .A1(new_n2615_), .B0(new_n2682_), .Y(new_n2683_));
  XOR2X1   g2634(.A(new_n2683_), .B(new_n2681_), .Y(new_n2684_));
  AOI22X1  g2635(.A0(new_n1727_), .A1(new_n1584_), .B0(new_n1724_), .B1(new_n1695_), .Y(new_n2685_));
  OAI21X1  g2636(.A0(new_n1730_), .A1(new_n1673_), .B0(new_n2685_), .Y(new_n2686_));
  AOI21X1  g2637(.A0(new_n1721_), .A1(new_n1690_), .B0(new_n2686_), .Y(new_n2687_));
  XOR2X1   g2638(.A(new_n2687_), .B(new_n312_), .Y(new_n2688_));
  XOR2X1   g2639(.A(new_n2688_), .B(new_n2684_), .Y(new_n2689_));
  XOR2X1   g2640(.A(new_n2689_), .B(new_n2673_), .Y(new_n2690_));
  INVX1    g2641(.A(new_n2063_), .Y(new_n2691_));
  AOI22X1  g2642(.A0(new_n2052_), .A1(new_n1796_), .B0(new_n2044_), .B1(new_n1804_), .Y(new_n2692_));
  OAI21X1  g2643(.A0(new_n2039_), .A1(new_n1802_), .B0(new_n2692_), .Y(new_n2693_));
  AOI21X1  g2644(.A0(new_n2691_), .A1(new_n1809_), .B0(new_n2693_), .Y(new_n2694_));
  XOR2X1   g2645(.A(new_n2694_), .B(new_n1164_), .Y(new_n2695_));
  XOR2X1   g2646(.A(new_n2695_), .B(new_n2690_), .Y(new_n2696_));
  XOR2X1   g2647(.A(new_n2696_), .B(new_n2671_), .Y(new_n2697_));
  AOI22X1  g2648(.A0(new_n2368_), .A1(new_n1693_), .B0(new_n2286_), .B1(new_n1699_), .Y(new_n2698_));
  OAI21X1  g2649(.A0(new_n2442_), .A1(new_n1906_), .B0(new_n2698_), .Y(new_n2699_));
  AOI21X1  g2650(.A0(new_n2441_), .A1(new_n245_), .B0(new_n2699_), .Y(new_n2700_));
  XOR2X1   g2651(.A(new_n2700_), .B(new_n229_), .Y(new_n2701_));
  XOR2X1   g2652(.A(new_n2701_), .B(new_n2697_), .Y(new_n2702_));
  XOR2X1   g2653(.A(new_n2702_), .B(new_n2666_), .Y(new_n2703_));
  XOR2X1   g2654(.A(new_n2703_), .B(new_n2663_), .Y(new_n2704_));
  XOR2X1   g2655(.A(new_n2704_), .B(new_n2659_), .Y(new_n2705_));
  XOR2X1   g2656(.A(new_n2705_), .B(new_n2653_), .Y(new_n2706_));
  XOR2X1   g2657(.A(new_n2706_), .B(new_n2650_), .Y(new_n2707_));
  NOR2X1   g2658(.A(new_n2582_), .B(new_n2581_), .Y(new_n2708_));
  AND2X1   g2659(.A(new_n2708_), .B(new_n2647_), .Y(new_n2709_));
  OR2X1    g2660(.A(new_n2709_), .B(new_n2503_), .Y(new_n2710_));
  XOR2X1   g2661(.A(new_n2710_), .B(new_n2707_), .Y(\sin[4] ));
  INVX1    g2662(.A(new_n2659_), .Y(new_n2712_));
  XOR2X1   g2663(.A(new_n2704_), .B(new_n2712_), .Y(new_n2713_));
  XOR2X1   g2664(.A(new_n2713_), .B(new_n2653_), .Y(new_n2714_));
  AND2X1   g2665(.A(new_n2714_), .B(new_n2650_), .Y(new_n2715_));
  AND2X1   g2666(.A(new_n2704_), .B(new_n2712_), .Y(new_n2716_));
  AOI21X1  g2667(.A0(new_n2713_), .A1(new_n2653_), .B0(new_n2716_), .Y(new_n2717_));
  NOR2X1   g2668(.A(new_n2432_), .B(new_n344_), .Y(new_n2718_));
  NOR3X1   g2669(.A(new_n305_), .B(new_n397_), .C(new_n248_), .Y(new_n2719_));
  NOR4X1   g2670(.A(new_n372_), .B(new_n261_), .C(new_n168_), .D(new_n139_), .Y(new_n2720_));
  NAND3X1  g2671(.A(new_n2720_), .B(new_n2719_), .C(new_n2497_), .Y(new_n2721_));
  INVX1    g2672(.A(new_n2721_), .Y(new_n2722_));
  OR4X1    g2673(.A(new_n388_), .B(new_n173_), .C(new_n172_), .D(new_n125_), .Y(new_n2723_));
  NOR3X1   g2674(.A(new_n2723_), .B(new_n1389_), .C(new_n726_), .Y(new_n2724_));
  AND2X1   g2675(.A(new_n2724_), .B(new_n1393_), .Y(new_n2725_));
  NAND4X1  g2676(.A(new_n2725_), .B(new_n2722_), .C(new_n2718_), .D(new_n2024_), .Y(new_n2726_));
  AND2X1   g2677(.A(new_n2702_), .B(new_n2666_), .Y(new_n2727_));
  INVX1    g2678(.A(new_n2727_), .Y(new_n2728_));
  OAI21X1  g2679(.A0(new_n2662_), .A1(new_n2661_), .B0(new_n2703_), .Y(new_n2729_));
  NAND2X1  g2680(.A(new_n2729_), .B(new_n2728_), .Y(new_n2730_));
  OAI21X1  g2681(.A0(new_n2670_), .A1(new_n2668_), .B0(new_n2696_), .Y(new_n2731_));
  NAND2X1  g2682(.A(new_n2701_), .B(new_n2697_), .Y(new_n2732_));
  NAND2X1  g2683(.A(new_n2732_), .B(new_n2731_), .Y(new_n2733_));
  INVX1    g2684(.A(new_n2673_), .Y(new_n2734_));
  OR2X1    g2685(.A(new_n2695_), .B(new_n2690_), .Y(new_n2735_));
  OAI21X1  g2686(.A0(new_n2689_), .A1(new_n2734_), .B0(new_n2735_), .Y(new_n2736_));
  INVX1    g2687(.A(new_n2292_), .Y(new_n2737_));
  INVX1    g2688(.A(new_n2286_), .Y(new_n2738_));
  AOI22X1  g2689(.A0(new_n2052_), .A1(new_n1804_), .B0(new_n2040_), .B1(new_n1796_), .Y(new_n2739_));
  OAI21X1  g2690(.A0(new_n2738_), .A1(new_n1802_), .B0(new_n2739_), .Y(new_n2740_));
  AOI21X1  g2691(.A0(new_n2737_), .A1(new_n1809_), .B0(new_n2740_), .Y(new_n2741_));
  XOR2X1   g2692(.A(new_n2741_), .B(new_n1164_), .Y(new_n2742_));
  INVX1    g2693(.A(new_n2684_), .Y(new_n2743_));
  INVX1    g2694(.A(new_n2681_), .Y(new_n2744_));
  NOR2X1   g2695(.A(new_n2683_), .B(new_n2744_), .Y(new_n2745_));
  AOI21X1  g2696(.A0(new_n2688_), .A1(new_n2743_), .B0(new_n2745_), .Y(new_n2746_));
  OR2X1    g2697(.A(new_n2680_), .B(new_n2677_), .Y(new_n2747_));
  AND2X1   g2698(.A(new_n2747_), .B(new_n2678_), .Y(new_n2748_));
  NAND3X1  g2699(.A(new_n1618_), .B(new_n525_), .C(new_n243_), .Y(new_n2749_));
  AND2X1   g2700(.A(new_n1618_), .B(new_n525_), .Y(new_n2750_));
  OAI21X1  g2701(.A0(new_n2750_), .A1(new_n243_), .B0(new_n2749_), .Y(new_n2751_));
  XOR2X1   g2702(.A(new_n2751_), .B(new_n2748_), .Y(new_n2752_));
  OAI22X1  g2703(.A0(new_n1785_), .A1(new_n1797_), .B0(new_n1714_), .B1(new_n1585_), .Y(new_n2753_));
  AOI21X1  g2704(.A0(new_n1710_), .A1(new_n1613_), .B0(new_n2753_), .Y(new_n2754_));
  OAI21X1  g2705(.A0(new_n1919_), .A1(new_n1784_), .B0(new_n2754_), .Y(new_n2755_));
  XOR2X1   g2706(.A(new_n2755_), .B(new_n525_), .Y(new_n2756_));
  XOR2X1   g2707(.A(new_n2756_), .B(new_n2752_), .Y(new_n2757_));
  AOI22X1  g2708(.A0(new_n1729_), .A1(new_n1695_), .B0(new_n1727_), .B1(new_n1676_), .Y(new_n2758_));
  OAI21X1  g2709(.A0(new_n2045_), .A1(new_n1750_), .B0(new_n2758_), .Y(new_n2759_));
  AOI21X1  g2710(.A0(new_n2075_), .A1(new_n1721_), .B0(new_n2759_), .Y(new_n2760_));
  XOR2X1   g2711(.A(new_n2760_), .B(new_n312_), .Y(new_n2761_));
  XOR2X1   g2712(.A(new_n2761_), .B(new_n2757_), .Y(new_n2762_));
  XOR2X1   g2713(.A(new_n2762_), .B(new_n2746_), .Y(new_n2763_));
  XOR2X1   g2714(.A(new_n2763_), .B(new_n2742_), .Y(new_n2764_));
  XOR2X1   g2715(.A(new_n2764_), .B(new_n2736_), .Y(new_n2765_));
  OAI22X1  g2716(.A0(new_n2442_), .A1(new_n1694_), .B0(new_n2371_), .B1(new_n1916_), .Y(new_n2766_));
  AOI21X1  g2717(.A0(new_n2530_), .A1(new_n245_), .B0(new_n2766_), .Y(new_n2767_));
  XOR2X1   g2718(.A(new_n2767_), .B(new_n229_), .Y(new_n2768_));
  XOR2X1   g2719(.A(new_n2768_), .B(new_n2765_), .Y(new_n2769_));
  XOR2X1   g2720(.A(new_n2769_), .B(new_n2733_), .Y(new_n2770_));
  XOR2X1   g2721(.A(new_n2770_), .B(new_n2730_), .Y(new_n2771_));
  XOR2X1   g2722(.A(new_n2771_), .B(new_n2726_), .Y(new_n2772_));
  XOR2X1   g2723(.A(new_n2772_), .B(new_n2717_), .Y(new_n2773_));
  XOR2X1   g2724(.A(new_n2773_), .B(new_n2715_), .Y(new_n2774_));
  AND2X1   g2725(.A(new_n2709_), .B(new_n2707_), .Y(new_n2775_));
  OR2X1    g2726(.A(new_n2775_), .B(new_n2503_), .Y(new_n2776_));
  XOR2X1   g2727(.A(new_n2776_), .B(new_n2774_), .Y(\sin[5] ));
  INVX1    g2728(.A(new_n2726_), .Y(new_n2778_));
  XOR2X1   g2729(.A(new_n2771_), .B(new_n2778_), .Y(new_n2779_));
  XOR2X1   g2730(.A(new_n2779_), .B(new_n2717_), .Y(new_n2780_));
  AND2X1   g2731(.A(new_n2780_), .B(new_n2715_), .Y(new_n2781_));
  NAND2X1  g2732(.A(new_n2771_), .B(new_n2726_), .Y(new_n2782_));
  OAI21X1  g2733(.A0(new_n2779_), .A1(new_n2717_), .B0(new_n2782_), .Y(new_n2783_));
  OR4X1    g2734(.A(new_n1389_), .B(new_n452_), .C(new_n304_), .D(new_n181_), .Y(new_n2784_));
  OR4X1    g2735(.A(new_n2492_), .B(new_n497_), .C(new_n551_), .D(new_n196_), .Y(new_n2785_));
  NOR4X1   g2736(.A(new_n2785_), .B(new_n2784_), .C(new_n1456_), .D(new_n572_), .Y(new_n2786_));
  INVX1    g2737(.A(new_n2786_), .Y(new_n2787_));
  NOR4X1   g2738(.A(new_n385_), .B(new_n337_), .C(new_n170_), .D(new_n162_), .Y(new_n2788_));
  NOR2X1   g2739(.A(new_n322_), .B(new_n265_), .Y(new_n2789_));
  INVX1    g2740(.A(new_n2789_), .Y(new_n2790_));
  NOR4X1   g2741(.A(new_n2033_), .B(new_n2790_), .C(new_n184_), .D(new_n183_), .Y(new_n2791_));
  NAND3X1  g2742(.A(new_n2791_), .B(new_n2788_), .C(new_n1471_), .Y(new_n2792_));
  NOR3X1   g2743(.A(new_n2792_), .B(new_n2787_), .C(new_n153_), .Y(new_n2793_));
  AND2X1   g2744(.A(new_n2769_), .B(new_n2733_), .Y(new_n2794_));
  INVX1    g2745(.A(new_n2794_), .Y(new_n2795_));
  INVX1    g2746(.A(new_n2661_), .Y(new_n2796_));
  NOR2X1   g2747(.A(new_n2570_), .B(new_n2595_), .Y(new_n2797_));
  OR2X1    g2748(.A(new_n2485_), .B(new_n2446_), .Y(new_n2798_));
  NOR2X1   g2749(.A(new_n2408_), .B(new_n2375_), .Y(new_n2799_));
  XOR2X1   g2750(.A(new_n2374_), .B(new_n2081_), .Y(new_n2800_));
  XOR2X1   g2751(.A(new_n2408_), .B(new_n2800_), .Y(new_n2801_));
  AOI21X1  g2752(.A0(new_n2296_), .A1(new_n2410_), .B0(new_n2801_), .Y(new_n2802_));
  OAI21X1  g2753(.A0(new_n2802_), .A1(new_n2799_), .B0(new_n2486_), .Y(new_n2803_));
  AOI21X1  g2754(.A0(new_n2803_), .A1(new_n2798_), .B0(new_n2571_), .Y(new_n2804_));
  XOR2X1   g2755(.A(new_n2641_), .B(new_n2660_), .Y(new_n2805_));
  OAI21X1  g2756(.A0(new_n2804_), .A1(new_n2797_), .B0(new_n2805_), .Y(new_n2806_));
  AND2X1   g2757(.A(new_n2665_), .B(new_n2664_), .Y(new_n2807_));
  XOR2X1   g2758(.A(new_n2702_), .B(new_n2807_), .Y(new_n2808_));
  AOI21X1  g2759(.A0(new_n2806_), .A1(new_n2796_), .B0(new_n2808_), .Y(new_n2809_));
  OAI21X1  g2760(.A0(new_n2809_), .A1(new_n2727_), .B0(new_n2770_), .Y(new_n2810_));
  NAND2X1  g2761(.A(new_n2810_), .B(new_n2795_), .Y(new_n2811_));
  AND2X1   g2762(.A(new_n2764_), .B(new_n2736_), .Y(new_n2812_));
  AOI21X1  g2763(.A0(new_n2768_), .A1(new_n2765_), .B0(new_n2812_), .Y(new_n2813_));
  INVX1    g2764(.A(new_n2813_), .Y(new_n2814_));
  INVX1    g2765(.A(new_n2746_), .Y(new_n2815_));
  NOR2X1   g2766(.A(new_n2763_), .B(new_n2742_), .Y(new_n2816_));
  AOI21X1  g2767(.A0(new_n2762_), .A1(new_n2815_), .B0(new_n2816_), .Y(new_n2817_));
  AOI22X1  g2768(.A0(new_n2529_), .A1(new_n245_), .B0(new_n2438_), .B1(new_n1699_), .Y(new_n2818_));
  XOR2X1   g2769(.A(new_n2818_), .B(new_n230_), .Y(new_n2819_));
  XOR2X1   g2770(.A(new_n2819_), .B(new_n2817_), .Y(new_n2820_));
  AOI22X1  g2771(.A0(new_n2286_), .A1(new_n1796_), .B0(new_n2040_), .B1(new_n1804_), .Y(new_n2821_));
  OAI21X1  g2772(.A0(new_n2371_), .A1(new_n1802_), .B0(new_n2821_), .Y(new_n2822_));
  AOI21X1  g2773(.A0(new_n2370_), .A1(new_n1809_), .B0(new_n2822_), .Y(new_n2823_));
  XOR2X1   g2774(.A(new_n2823_), .B(new_n1164_), .Y(new_n2824_));
  AND2X1   g2775(.A(new_n2756_), .B(new_n2752_), .Y(new_n2825_));
  AOI21X1  g2776(.A0(new_n2761_), .A1(new_n2757_), .B0(new_n2825_), .Y(new_n2826_));
  OR2X1    g2777(.A(new_n2751_), .B(new_n2748_), .Y(new_n2827_));
  AND2X1   g2778(.A(new_n2827_), .B(new_n2749_), .Y(new_n2828_));
  NAND3X1  g2779(.A(new_n1615_), .B(new_n525_), .C(new_n243_), .Y(new_n2829_));
  AND2X1   g2780(.A(new_n1615_), .B(new_n525_), .Y(new_n2830_));
  OAI21X1  g2781(.A0(new_n2830_), .A1(new_n243_), .B0(new_n2829_), .Y(new_n2831_));
  XOR2X1   g2782(.A(new_n2831_), .B(new_n2828_), .Y(new_n2832_));
  OAI22X1  g2783(.A0(new_n1785_), .A1(new_n2198_), .B0(new_n1711_), .B1(new_n1585_), .Y(new_n2833_));
  AOI21X1  g2784(.A0(new_n1713_), .A1(new_n1676_), .B0(new_n2833_), .Y(new_n2834_));
  OAI21X1  g2785(.A0(new_n2622_), .A1(new_n1784_), .B0(new_n2834_), .Y(new_n2835_));
  XOR2X1   g2786(.A(new_n2835_), .B(new_n525_), .Y(new_n2836_));
  XOR2X1   g2787(.A(new_n2836_), .B(new_n2832_), .Y(new_n2837_));
  AOI22X1  g2788(.A0(new_n2044_), .A1(new_n1729_), .B0(new_n1727_), .B1(new_n1695_), .Y(new_n2838_));
  OAI21X1  g2789(.A0(new_n2047_), .A1(new_n1750_), .B0(new_n2838_), .Y(new_n2839_));
  AOI21X1  g2790(.A0(new_n2605_), .A1(new_n1721_), .B0(new_n2839_), .Y(new_n2840_));
  XOR2X1   g2791(.A(new_n2840_), .B(new_n312_), .Y(new_n2841_));
  XOR2X1   g2792(.A(new_n2841_), .B(new_n2837_), .Y(new_n2842_));
  XOR2X1   g2793(.A(new_n2842_), .B(new_n2826_), .Y(new_n2843_));
  XOR2X1   g2794(.A(new_n2843_), .B(new_n2824_), .Y(new_n2844_));
  XOR2X1   g2795(.A(new_n2844_), .B(new_n2820_), .Y(new_n2845_));
  XOR2X1   g2796(.A(new_n2845_), .B(new_n2814_), .Y(new_n2846_));
  XOR2X1   g2797(.A(new_n2846_), .B(new_n2811_), .Y(new_n2847_));
  XOR2X1   g2798(.A(new_n2847_), .B(new_n2793_), .Y(new_n2848_));
  XOR2X1   g2799(.A(new_n2848_), .B(new_n2783_), .Y(new_n2849_));
  XOR2X1   g2800(.A(new_n2849_), .B(new_n2781_), .Y(new_n2850_));
  AND2X1   g2801(.A(new_n2775_), .B(new_n2774_), .Y(new_n2851_));
  OR2X1    g2802(.A(new_n2851_), .B(new_n2503_), .Y(new_n2852_));
  XOR2X1   g2803(.A(new_n2852_), .B(new_n2850_), .Y(\sin[6] ));
  INVX1    g2804(.A(new_n2793_), .Y(new_n2854_));
  XOR2X1   g2805(.A(new_n2847_), .B(new_n2854_), .Y(new_n2855_));
  XOR2X1   g2806(.A(new_n2855_), .B(new_n2783_), .Y(new_n2856_));
  AND2X1   g2807(.A(new_n2856_), .B(new_n2781_), .Y(new_n2857_));
  AND2X1   g2808(.A(new_n2847_), .B(new_n2854_), .Y(new_n2858_));
  AOI21X1  g2809(.A0(new_n2855_), .A1(new_n2783_), .B0(new_n2858_), .Y(new_n2859_));
  NOR2X1   g2810(.A(new_n2819_), .B(new_n2817_), .Y(new_n2860_));
  AOI21X1  g2811(.A0(new_n2844_), .A1(new_n2820_), .B0(new_n2860_), .Y(new_n2861_));
  INVX1    g2812(.A(new_n2826_), .Y(new_n2862_));
  AND2X1   g2813(.A(new_n2842_), .B(new_n2862_), .Y(new_n2863_));
  INVX1    g2814(.A(new_n2863_), .Y(new_n2864_));
  OAI21X1  g2815(.A0(new_n2843_), .A1(new_n2824_), .B0(new_n2864_), .Y(new_n2865_));
  AOI22X1  g2816(.A0(new_n2368_), .A1(new_n1796_), .B0(new_n2286_), .B1(new_n1804_), .Y(new_n2866_));
  OAI21X1  g2817(.A0(new_n2442_), .A1(new_n1802_), .B0(new_n2866_), .Y(new_n2867_));
  AOI21X1  g2818(.A0(new_n2441_), .A1(new_n1809_), .B0(new_n2867_), .Y(new_n2868_));
  XOR2X1   g2819(.A(new_n2868_), .B(new_n519_), .Y(new_n2869_));
  XOR2X1   g2820(.A(new_n2869_), .B(new_n2865_), .Y(new_n2870_));
  AND2X1   g2821(.A(new_n2836_), .B(new_n2832_), .Y(new_n2871_));
  AOI21X1  g2822(.A0(new_n2841_), .A1(new_n2837_), .B0(new_n2871_), .Y(new_n2872_));
  OAI21X1  g2823(.A0(new_n2831_), .A1(new_n2828_), .B0(new_n2829_), .Y(new_n2873_));
  AOI22X1  g2824(.A0(new_n1877_), .A1(new_n1584_), .B0(new_n1713_), .B1(new_n1695_), .Y(new_n2874_));
  OAI21X1  g2825(.A0(new_n1711_), .A1(new_n1673_), .B0(new_n2874_), .Y(new_n2875_));
  AOI21X1  g2826(.A0(new_n1707_), .A1(new_n1690_), .B0(new_n2875_), .Y(new_n2876_));
  XOR2X1   g2827(.A(new_n2876_), .B(new_n525_), .Y(new_n2877_));
  AND2X1   g2828(.A(new_n1613_), .B(new_n525_), .Y(new_n2878_));
  XOR2X1   g2829(.A(new_n2081_), .B(new_n229_), .Y(new_n2879_));
  XOR2X1   g2830(.A(new_n2879_), .B(new_n2878_), .Y(new_n2880_));
  XOR2X1   g2831(.A(new_n2880_), .B(new_n2877_), .Y(new_n2881_));
  XOR2X1   g2832(.A(new_n2881_), .B(new_n2873_), .Y(new_n2882_));
  INVX1    g2833(.A(new_n2882_), .Y(new_n2883_));
  OAI22X1  g2834(.A0(new_n2047_), .A1(new_n1730_), .B0(new_n2045_), .B1(new_n1728_), .Y(new_n2884_));
  AOI21X1  g2835(.A0(new_n2040_), .A1(new_n1724_), .B0(new_n2884_), .Y(new_n2885_));
  OAI21X1  g2836(.A0(new_n2063_), .A1(new_n1722_), .B0(new_n2885_), .Y(new_n2886_));
  XOR2X1   g2837(.A(new_n2886_), .B(new_n313_), .Y(new_n2887_));
  XOR2X1   g2838(.A(new_n2887_), .B(new_n2883_), .Y(new_n2888_));
  XOR2X1   g2839(.A(new_n2888_), .B(new_n2872_), .Y(new_n2889_));
  XOR2X1   g2840(.A(new_n2889_), .B(new_n2870_), .Y(new_n2890_));
  XOR2X1   g2841(.A(new_n2890_), .B(new_n2861_), .Y(new_n2891_));
  AND2X1   g2842(.A(new_n2845_), .B(new_n2814_), .Y(new_n2892_));
  INVX1    g2843(.A(new_n2846_), .Y(new_n2893_));
  AOI21X1  g2844(.A0(new_n2810_), .A1(new_n2795_), .B0(new_n2893_), .Y(new_n2894_));
  NOR2X1   g2845(.A(new_n2894_), .B(new_n2892_), .Y(new_n2895_));
  XOR2X1   g2846(.A(new_n2895_), .B(new_n2891_), .Y(new_n2896_));
  OR4X1    g2847(.A(new_n264_), .B(new_n253_), .C(new_n252_), .D(new_n195_), .Y(new_n2897_));
  OR4X1    g2848(.A(new_n2897_), .B(new_n547_), .C(new_n219_), .D(new_n190_), .Y(new_n2898_));
  NOR4X1   g2849(.A(new_n347_), .B(new_n169_), .C(new_n159_), .D(new_n134_), .Y(new_n2899_));
  NAND2X1  g2850(.A(new_n2899_), .B(new_n2719_), .Y(new_n2900_));
  NOR4X1   g2851(.A(new_n2900_), .B(new_n2898_), .C(new_n2787_), .D(new_n1369_), .Y(new_n2901_));
  XOR2X1   g2852(.A(new_n2901_), .B(new_n2896_), .Y(new_n2902_));
  XOR2X1   g2853(.A(new_n2902_), .B(new_n2859_), .Y(new_n2903_));
  XOR2X1   g2854(.A(new_n2903_), .B(new_n2857_), .Y(new_n2904_));
  AND2X1   g2855(.A(new_n2851_), .B(new_n2850_), .Y(new_n2905_));
  OR2X1    g2856(.A(new_n2905_), .B(new_n2503_), .Y(new_n2906_));
  XOR2X1   g2857(.A(new_n2906_), .B(new_n2904_), .Y(\sin[7] ));
  OAI21X1  g2858(.A0(new_n2573_), .A1(new_n2576_), .B0(new_n2577_), .Y(new_n2908_));
  AND2X1   g2859(.A(new_n2643_), .B(new_n2651_), .Y(new_n2909_));
  XOR2X1   g2860(.A(new_n2643_), .B(new_n2651_), .Y(new_n2910_));
  AOI21X1  g2861(.A0(new_n2910_), .A1(new_n2908_), .B0(new_n2909_), .Y(new_n2911_));
  NAND2X1  g2862(.A(new_n2704_), .B(new_n2712_), .Y(new_n2912_));
  OAI21X1  g2863(.A0(new_n2705_), .A1(new_n2911_), .B0(new_n2912_), .Y(new_n2913_));
  AND2X1   g2864(.A(new_n2771_), .B(new_n2726_), .Y(new_n2914_));
  AOI21X1  g2865(.A0(new_n2772_), .A1(new_n2913_), .B0(new_n2914_), .Y(new_n2915_));
  NAND2X1  g2866(.A(new_n2847_), .B(new_n2854_), .Y(new_n2916_));
  OAI21X1  g2867(.A0(new_n2848_), .A1(new_n2915_), .B0(new_n2916_), .Y(new_n2917_));
  XOR2X1   g2868(.A(new_n2902_), .B(new_n2917_), .Y(new_n2918_));
  AND2X1   g2869(.A(new_n2918_), .B(new_n2857_), .Y(new_n2919_));
  NOR2X1   g2870(.A(new_n2901_), .B(new_n2896_), .Y(new_n2920_));
  AOI21X1  g2871(.A0(new_n2902_), .A1(new_n2917_), .B0(new_n2920_), .Y(new_n2921_));
  NOR3X1   g2872(.A(new_n256_), .B(new_n125_), .C(new_n107_), .Y(new_n2922_));
  NOR4X1   g2873(.A(new_n203_), .B(new_n175_), .C(new_n145_), .D(new_n121_), .Y(new_n2923_));
  NAND3X1  g2874(.A(new_n2923_), .B(new_n2922_), .C(new_n701_), .Y(new_n2924_));
  OR4X1    g2875(.A(new_n2924_), .B(new_n1520_), .C(new_n213_), .D(new_n150_), .Y(new_n2925_));
  NOR2X1   g2876(.A(new_n2925_), .B(new_n201_), .Y(new_n2926_));
  OR4X1    g2877(.A(new_n527_), .B(new_n216_), .C(new_n210_), .D(new_n97_), .Y(new_n2927_));
  OR4X1    g2878(.A(new_n2927_), .B(new_n616_), .C(new_n265_), .D(new_n259_), .Y(new_n2928_));
  NAND4X1  g2879(.A(new_n1411_), .B(new_n301_), .C(new_n300_), .D(new_n299_), .Y(new_n2929_));
  NOR3X1   g2880(.A(new_n2929_), .B(new_n2928_), .C(new_n498_), .Y(new_n2930_));
  NAND3X1  g2881(.A(new_n2930_), .B(new_n2926_), .C(new_n2322_), .Y(new_n2931_));
  OAI21X1  g2882(.A0(new_n2894_), .A1(new_n2892_), .B0(new_n2891_), .Y(new_n2932_));
  NOR2X1   g2883(.A(new_n2890_), .B(new_n2861_), .Y(new_n2933_));
  INVX1    g2884(.A(new_n2933_), .Y(new_n2934_));
  NAND2X1  g2885(.A(new_n2934_), .B(new_n2932_), .Y(new_n2935_));
  AND2X1   g2886(.A(new_n2869_), .B(new_n2865_), .Y(new_n2936_));
  INVX1    g2887(.A(new_n2936_), .Y(new_n2937_));
  INVX1    g2888(.A(new_n2870_), .Y(new_n2938_));
  OAI21X1  g2889(.A0(new_n2889_), .A1(new_n2938_), .B0(new_n2937_), .Y(new_n2939_));
  OAI22X1  g2890(.A0(new_n2442_), .A1(new_n1824_), .B0(new_n2371_), .B1(new_n1805_), .Y(new_n2940_));
  AOI21X1  g2891(.A0(new_n2530_), .A1(new_n1809_), .B0(new_n2940_), .Y(new_n2941_));
  XOR2X1   g2892(.A(new_n2941_), .B(new_n519_), .Y(new_n2942_));
  NAND2X1  g2893(.A(new_n2887_), .B(new_n2883_), .Y(new_n2943_));
  XOR2X1   g2894(.A(new_n2887_), .B(new_n2882_), .Y(new_n2944_));
  OAI21X1  g2895(.A0(new_n2944_), .A1(new_n2872_), .B0(new_n2943_), .Y(new_n2945_));
  INVX1    g2896(.A(new_n2873_), .Y(new_n2946_));
  INVX1    g2897(.A(new_n2877_), .Y(new_n2947_));
  NAND2X1  g2898(.A(new_n2880_), .B(new_n2947_), .Y(new_n2948_));
  OAI21X1  g2899(.A0(new_n2881_), .A1(new_n2946_), .B0(new_n2948_), .Y(new_n2949_));
  AND2X1   g2900(.A(new_n1584_), .B(new_n525_), .Y(new_n2950_));
  AND2X1   g2901(.A(new_n2081_), .B(new_n229_), .Y(new_n2951_));
  AOI21X1  g2902(.A0(new_n2879_), .A1(new_n2878_), .B0(new_n2951_), .Y(new_n2952_));
  XOR2X1   g2903(.A(new_n2952_), .B(new_n2950_), .Y(new_n2953_));
  AOI22X1  g2904(.A0(new_n1877_), .A1(new_n1676_), .B0(new_n1710_), .B1(new_n1695_), .Y(new_n2954_));
  OAI21X1  g2905(.A0(new_n2045_), .A1(new_n1714_), .B0(new_n2954_), .Y(new_n2955_));
  AOI21X1  g2906(.A0(new_n2075_), .A1(new_n1707_), .B0(new_n2955_), .Y(new_n2956_));
  XOR2X1   g2907(.A(new_n2956_), .B(new_n793_), .Y(new_n2957_));
  XOR2X1   g2908(.A(new_n2957_), .B(new_n2953_), .Y(new_n2958_));
  XOR2X1   g2909(.A(new_n2958_), .B(new_n2949_), .Y(new_n2959_));
  AOI22X1  g2910(.A0(new_n2052_), .A1(new_n1727_), .B0(new_n2040_), .B1(new_n1729_), .Y(new_n2960_));
  OAI21X1  g2911(.A0(new_n2738_), .A1(new_n1750_), .B0(new_n2960_), .Y(new_n2961_));
  AOI21X1  g2912(.A0(new_n2737_), .A1(new_n1721_), .B0(new_n2961_), .Y(new_n2962_));
  XOR2X1   g2913(.A(new_n2962_), .B(new_n312_), .Y(new_n2963_));
  XOR2X1   g2914(.A(new_n2963_), .B(new_n2959_), .Y(new_n2964_));
  XOR2X1   g2915(.A(new_n2964_), .B(new_n2945_), .Y(new_n2965_));
  XOR2X1   g2916(.A(new_n2965_), .B(new_n2942_), .Y(new_n2966_));
  XOR2X1   g2917(.A(new_n2966_), .B(new_n2939_), .Y(new_n2967_));
  XOR2X1   g2918(.A(new_n2967_), .B(new_n2935_), .Y(new_n2968_));
  XOR2X1   g2919(.A(new_n2968_), .B(new_n2931_), .Y(new_n2969_));
  XOR2X1   g2920(.A(new_n2969_), .B(new_n2921_), .Y(new_n2970_));
  XOR2X1   g2921(.A(new_n2970_), .B(new_n2919_), .Y(new_n2971_));
  AND2X1   g2922(.A(new_n2905_), .B(new_n2904_), .Y(new_n2972_));
  OR2X1    g2923(.A(new_n2972_), .B(new_n2503_), .Y(new_n2973_));
  XOR2X1   g2924(.A(new_n2973_), .B(new_n2971_), .Y(\sin[8] ));
  OR2X1    g2925(.A(new_n2901_), .B(new_n2896_), .Y(new_n2975_));
  AND2X1   g2926(.A(new_n2901_), .B(new_n2896_), .Y(new_n2976_));
  OAI21X1  g2927(.A0(new_n2976_), .A1(new_n2859_), .B0(new_n2975_), .Y(new_n2977_));
  XOR2X1   g2928(.A(new_n2969_), .B(new_n2977_), .Y(new_n2978_));
  AND2X1   g2929(.A(new_n2978_), .B(new_n2919_), .Y(new_n2979_));
  AND2X1   g2930(.A(new_n2968_), .B(new_n2931_), .Y(new_n2980_));
  AOI21X1  g2931(.A0(new_n2969_), .A1(new_n2977_), .B0(new_n2980_), .Y(new_n2981_));
  OR4X1    g2932(.A(new_n198_), .B(new_n136_), .C(new_n131_), .D(new_n107_), .Y(new_n2982_));
  NOR3X1   g2933(.A(new_n2982_), .B(new_n2033_), .C(new_n547_), .Y(new_n2983_));
  NOR4X1   g2934(.A(new_n2018_), .B(new_n385_), .C(new_n269_), .D(new_n264_), .Y(new_n2984_));
  NAND3X1  g2935(.A(new_n2984_), .B(new_n2983_), .C(new_n418_), .Y(new_n2985_));
  NOR3X1   g2936(.A(new_n2985_), .B(new_n1459_), .C(new_n177_), .Y(new_n2986_));
  INVX1    g2937(.A(new_n2986_), .Y(new_n2987_));
  AND2X1   g2938(.A(new_n2964_), .B(new_n2945_), .Y(new_n2988_));
  AOI21X1  g2939(.A0(new_n2965_), .A1(new_n2942_), .B0(new_n2988_), .Y(new_n2989_));
  NOR2X1   g2940(.A(new_n2952_), .B(new_n2950_), .Y(new_n2990_));
  AOI21X1  g2941(.A0(new_n2957_), .A1(new_n2953_), .B0(new_n2990_), .Y(new_n2991_));
  INVX1    g2942(.A(new_n2991_), .Y(new_n2992_));
  AOI22X1  g2943(.A0(new_n2044_), .A1(new_n1710_), .B0(new_n1877_), .B1(new_n1695_), .Y(new_n2993_));
  OAI21X1  g2944(.A0(new_n2047_), .A1(new_n1714_), .B0(new_n2993_), .Y(new_n2994_));
  AOI21X1  g2945(.A0(new_n2605_), .A1(new_n1707_), .B0(new_n2994_), .Y(new_n2995_));
  XOR2X1   g2946(.A(new_n2995_), .B(new_n793_), .Y(new_n2996_));
  AND2X1   g2947(.A(new_n1674_), .B(new_n525_), .Y(new_n2997_));
  XOR2X1   g2948(.A(new_n2997_), .B(new_n2996_), .Y(new_n2998_));
  XOR2X1   g2949(.A(new_n2998_), .B(new_n2992_), .Y(new_n2999_));
  AOI22X1  g2950(.A0(new_n2286_), .A1(new_n1729_), .B0(new_n2040_), .B1(new_n1727_), .Y(new_n3000_));
  OAI21X1  g2951(.A0(new_n2371_), .A1(new_n1750_), .B0(new_n3000_), .Y(new_n3001_));
  AOI21X1  g2952(.A0(new_n2370_), .A1(new_n1721_), .B0(new_n3001_), .Y(new_n3002_));
  XOR2X1   g2953(.A(new_n3002_), .B(new_n312_), .Y(new_n3003_));
  XOR2X1   g2954(.A(new_n3003_), .B(new_n2999_), .Y(new_n3004_));
  AND2X1   g2955(.A(new_n2958_), .B(new_n2949_), .Y(new_n3005_));
  AOI21X1  g2956(.A0(new_n2963_), .A1(new_n2959_), .B0(new_n3005_), .Y(new_n3006_));
  AOI22X1  g2957(.A0(new_n2529_), .A1(new_n1809_), .B0(new_n2438_), .B1(new_n1804_), .Y(new_n3007_));
  XOR2X1   g2958(.A(new_n3007_), .B(new_n1164_), .Y(new_n3008_));
  XOR2X1   g2959(.A(new_n3008_), .B(new_n3006_), .Y(new_n3009_));
  XOR2X1   g2960(.A(new_n3009_), .B(new_n3004_), .Y(new_n3010_));
  XOR2X1   g2961(.A(new_n3010_), .B(new_n2989_), .Y(new_n3011_));
  INVX1    g2962(.A(new_n3011_), .Y(new_n3012_));
  AND2X1   g2963(.A(new_n2966_), .B(new_n2939_), .Y(new_n3013_));
  INVX1    g2964(.A(new_n3013_), .Y(new_n3014_));
  INVX1    g2965(.A(new_n2892_), .Y(new_n3015_));
  AND2X1   g2966(.A(new_n2732_), .B(new_n2731_), .Y(new_n3016_));
  XOR2X1   g2967(.A(new_n2769_), .B(new_n3016_), .Y(new_n3017_));
  AOI21X1  g2968(.A0(new_n2729_), .A1(new_n2728_), .B0(new_n3017_), .Y(new_n3018_));
  OAI21X1  g2969(.A0(new_n3018_), .A1(new_n2794_), .B0(new_n2846_), .Y(new_n3019_));
  INVX1    g2970(.A(new_n2891_), .Y(new_n3020_));
  AOI21X1  g2971(.A0(new_n3019_), .A1(new_n3015_), .B0(new_n3020_), .Y(new_n3021_));
  OAI21X1  g2972(.A0(new_n2933_), .A1(new_n3021_), .B0(new_n2967_), .Y(new_n3022_));
  AND2X1   g2973(.A(new_n3022_), .B(new_n3014_), .Y(new_n3023_));
  XOR2X1   g2974(.A(new_n3023_), .B(new_n3012_), .Y(new_n3024_));
  XOR2X1   g2975(.A(new_n3024_), .B(new_n2987_), .Y(new_n3025_));
  XOR2X1   g2976(.A(new_n3025_), .B(new_n2981_), .Y(new_n3026_));
  XOR2X1   g2977(.A(new_n3026_), .B(new_n2979_), .Y(new_n3027_));
  AND2X1   g2978(.A(new_n2972_), .B(new_n2971_), .Y(new_n3028_));
  OR2X1    g2979(.A(new_n3028_), .B(new_n2503_), .Y(new_n3029_));
  XOR2X1   g2980(.A(new_n3029_), .B(new_n3027_), .Y(\sin[9] ));
  NOR2X1   g2981(.A(new_n2968_), .B(new_n2931_), .Y(new_n3031_));
  NAND2X1  g2982(.A(new_n2968_), .B(new_n2931_), .Y(new_n3032_));
  OAI21X1  g2983(.A0(new_n3031_), .A1(new_n2921_), .B0(new_n3032_), .Y(new_n3033_));
  XOR2X1   g2984(.A(new_n3025_), .B(new_n3033_), .Y(new_n3034_));
  AND2X1   g2985(.A(new_n3034_), .B(new_n2979_), .Y(new_n3035_));
  AND2X1   g2986(.A(new_n3024_), .B(new_n2987_), .Y(new_n3036_));
  AOI21X1  g2987(.A0(new_n3025_), .A1(new_n3033_), .B0(new_n3036_), .Y(new_n3037_));
  NOR3X1   g2988(.A(new_n2033_), .B(new_n529_), .C(new_n212_), .Y(new_n3038_));
  NOR3X1   g2989(.A(new_n363_), .B(new_n271_), .C(new_n158_), .Y(new_n3039_));
  NOR4X1   g2990(.A(new_n497_), .B(new_n319_), .C(new_n163_), .D(new_n162_), .Y(new_n3040_));
  NAND4X1  g2991(.A(new_n3040_), .B(new_n3039_), .C(new_n3038_), .D(new_n217_), .Y(new_n3041_));
  NOR4X1   g2992(.A(new_n3041_), .B(new_n2327_), .C(new_n613_), .D(new_n267_), .Y(new_n3042_));
  INVX1    g2993(.A(new_n3042_), .Y(new_n3043_));
  INVX1    g2994(.A(new_n2967_), .Y(new_n3044_));
  AOI21X1  g2995(.A0(new_n2934_), .A1(new_n2932_), .B0(new_n3044_), .Y(new_n3045_));
  OAI21X1  g2996(.A0(new_n3045_), .A1(new_n3013_), .B0(new_n3011_), .Y(new_n3046_));
  NOR2X1   g2997(.A(new_n3010_), .B(new_n2989_), .Y(new_n3047_));
  INVX1    g2998(.A(new_n3047_), .Y(new_n3048_));
  NAND2X1  g2999(.A(new_n3048_), .B(new_n3046_), .Y(new_n3049_));
  INVX1    g3000(.A(new_n3004_), .Y(new_n3050_));
  NOR2X1   g3001(.A(new_n3008_), .B(new_n3006_), .Y(new_n3051_));
  AOI21X1  g3002(.A0(new_n3009_), .A1(new_n3050_), .B0(new_n3051_), .Y(new_n3052_));
  INVX1    g3003(.A(new_n3052_), .Y(new_n3053_));
  INVX1    g3004(.A(new_n2999_), .Y(new_n3054_));
  NOR2X1   g3005(.A(new_n2998_), .B(new_n2991_), .Y(new_n3055_));
  AOI21X1  g3006(.A0(new_n3003_), .A1(new_n3054_), .B0(new_n3055_), .Y(new_n3056_));
  AOI22X1  g3007(.A0(new_n2368_), .A1(new_n1729_), .B0(new_n2286_), .B1(new_n1727_), .Y(new_n3057_));
  OAI21X1  g3008(.A0(new_n2442_), .A1(new_n1750_), .B0(new_n3057_), .Y(new_n3058_));
  AOI21X1  g3009(.A0(new_n2441_), .A1(new_n1721_), .B0(new_n3058_), .Y(new_n3059_));
  XOR2X1   g3010(.A(new_n3059_), .B(new_n312_), .Y(new_n3060_));
  NAND2X1  g3011(.A(new_n3060_), .B(new_n3056_), .Y(new_n3061_));
  INVX1    g3012(.A(new_n2997_), .Y(new_n3062_));
  NOR2X1   g3013(.A(new_n1584_), .B(new_n793_), .Y(new_n3063_));
  AOI22X1  g3014(.A0(new_n3063_), .A1(new_n1676_), .B0(new_n3062_), .B1(new_n2996_), .Y(new_n3064_));
  NOR3X1   g3015(.A(new_n1688_), .B(new_n793_), .C(new_n1164_), .Y(new_n3065_));
  AOI21X1  g3016(.A0(new_n1695_), .A1(new_n525_), .B0(new_n519_), .Y(new_n3066_));
  OR4X1    g3017(.A(new_n3066_), .B(new_n3065_), .C(new_n1585_), .D(new_n793_), .Y(new_n3067_));
  NOR3X1   g3018(.A(new_n3066_), .B(new_n3065_), .C(new_n2950_), .Y(new_n3068_));
  AOI21X1  g3019(.A0(new_n3067_), .A1(new_n2950_), .B0(new_n3068_), .Y(new_n3069_));
  XOR2X1   g3020(.A(new_n3069_), .B(new_n3064_), .Y(new_n3070_));
  AOI22X1  g3021(.A0(new_n2052_), .A1(new_n1710_), .B0(new_n2044_), .B1(new_n1877_), .Y(new_n3071_));
  OAI21X1  g3022(.A0(new_n2039_), .A1(new_n1714_), .B0(new_n3071_), .Y(new_n3072_));
  AOI21X1  g3023(.A0(new_n2691_), .A1(new_n1707_), .B0(new_n3072_), .Y(new_n3073_));
  XOR2X1   g3024(.A(new_n3073_), .B(new_n525_), .Y(new_n3074_));
  XOR2X1   g3025(.A(new_n3074_), .B(new_n3070_), .Y(new_n3075_));
  OR2X1    g3026(.A(new_n3060_), .B(new_n3056_), .Y(new_n3076_));
  AOI21X1  g3027(.A0(new_n3061_), .A1(new_n3076_), .B0(new_n3075_), .Y(new_n3077_));
  AND2X1   g3028(.A(new_n3076_), .B(new_n3075_), .Y(new_n3078_));
  AOI21X1  g3029(.A0(new_n3078_), .A1(new_n3061_), .B0(new_n3077_), .Y(new_n3079_));
  XOR2X1   g3030(.A(new_n3079_), .B(new_n3053_), .Y(new_n3080_));
  XOR2X1   g3031(.A(new_n3080_), .B(new_n3049_), .Y(new_n3081_));
  XOR2X1   g3032(.A(new_n3081_), .B(new_n3043_), .Y(new_n3082_));
  XOR2X1   g3033(.A(new_n3082_), .B(new_n3037_), .Y(new_n3083_));
  XOR2X1   g3034(.A(new_n3083_), .B(new_n3035_), .Y(new_n3084_));
  AND2X1   g3035(.A(new_n3028_), .B(new_n3027_), .Y(new_n3085_));
  OR2X1    g3036(.A(new_n3085_), .B(new_n2503_), .Y(new_n3086_));
  XOR2X1   g3037(.A(new_n3086_), .B(new_n3084_), .Y(\sin[10] ));
  NAND2X1  g3038(.A(new_n3024_), .B(new_n2987_), .Y(new_n3088_));
  XOR2X1   g3039(.A(new_n3024_), .B(new_n2986_), .Y(new_n3089_));
  OAI21X1  g3040(.A0(new_n3089_), .A1(new_n2981_), .B0(new_n3088_), .Y(new_n3090_));
  XOR2X1   g3041(.A(new_n3082_), .B(new_n3090_), .Y(new_n3091_));
  AND2X1   g3042(.A(new_n3091_), .B(new_n3035_), .Y(new_n3092_));
  AND2X1   g3043(.A(new_n3081_), .B(new_n3043_), .Y(new_n3093_));
  AOI21X1  g3044(.A0(new_n3082_), .A1(new_n3090_), .B0(new_n3093_), .Y(new_n3094_));
  OR4X1    g3045(.A(new_n505_), .B(new_n551_), .C(new_n287_), .D(new_n163_), .Y(new_n3095_));
  OR4X1    g3046(.A(new_n3095_), .B(new_n2361_), .C(new_n364_), .D(new_n342_), .Y(new_n3096_));
  NOR4X1   g3047(.A(new_n3096_), .B(new_n610_), .C(new_n533_), .D(new_n298_), .Y(new_n3097_));
  INVX1    g3048(.A(new_n3097_), .Y(new_n3098_));
  AND2X1   g3049(.A(new_n3079_), .B(new_n3053_), .Y(new_n3099_));
  INVX1    g3050(.A(new_n3080_), .Y(new_n3100_));
  AOI21X1  g3051(.A0(new_n3048_), .A1(new_n3046_), .B0(new_n3100_), .Y(new_n3101_));
  OR2X1    g3052(.A(new_n3101_), .B(new_n3099_), .Y(new_n3102_));
  INVX1    g3053(.A(new_n3056_), .Y(new_n3103_));
  AOI21X1  g3054(.A0(new_n3060_), .A1(new_n3103_), .B0(new_n3077_), .Y(new_n3104_));
  INVX1    g3055(.A(new_n3104_), .Y(new_n3105_));
  OR2X1    g3056(.A(new_n3069_), .B(new_n3064_), .Y(new_n3106_));
  INVX1    g3057(.A(new_n3070_), .Y(new_n3107_));
  OAI21X1  g3058(.A0(new_n3074_), .A1(new_n3107_), .B0(new_n3106_), .Y(new_n3108_));
  INVX1    g3059(.A(new_n3065_), .Y(new_n3109_));
  AND2X1   g3060(.A(new_n3067_), .B(new_n3109_), .Y(new_n3110_));
  AND2X1   g3061(.A(new_n2044_), .B(new_n525_), .Y(new_n3111_));
  XOR2X1   g3062(.A(new_n3111_), .B(new_n3110_), .Y(new_n3112_));
  OAI22X1  g3063(.A0(new_n2047_), .A1(new_n1785_), .B0(new_n2039_), .B1(new_n1711_), .Y(new_n3113_));
  AOI21X1  g3064(.A0(new_n2286_), .A1(new_n1713_), .B0(new_n3113_), .Y(new_n3114_));
  OAI21X1  g3065(.A0(new_n2292_), .A1(new_n1784_), .B0(new_n3114_), .Y(new_n3115_));
  XOR2X1   g3066(.A(new_n3115_), .B(new_n525_), .Y(new_n3116_));
  XOR2X1   g3067(.A(new_n3116_), .B(new_n3112_), .Y(new_n3117_));
  XOR2X1   g3068(.A(new_n3117_), .B(new_n3108_), .Y(new_n3118_));
  OAI22X1  g3069(.A0(new_n2442_), .A1(new_n1730_), .B0(new_n2371_), .B1(new_n1728_), .Y(new_n3119_));
  AOI21X1  g3070(.A0(new_n2530_), .A1(new_n1721_), .B0(new_n3119_), .Y(new_n3120_));
  XOR2X1   g3071(.A(new_n3120_), .B(new_n312_), .Y(new_n3121_));
  XOR2X1   g3072(.A(new_n3121_), .B(new_n3118_), .Y(new_n3122_));
  XOR2X1   g3073(.A(new_n3122_), .B(new_n3105_), .Y(new_n3123_));
  XOR2X1   g3074(.A(new_n3123_), .B(new_n3102_), .Y(new_n3124_));
  XOR2X1   g3075(.A(new_n3124_), .B(new_n3098_), .Y(new_n3125_));
  XOR2X1   g3076(.A(new_n3125_), .B(new_n3094_), .Y(new_n3126_));
  XOR2X1   g3077(.A(new_n3126_), .B(new_n3092_), .Y(new_n3127_));
  AND2X1   g3078(.A(new_n3085_), .B(new_n3084_), .Y(new_n3128_));
  OR2X1    g3079(.A(new_n3128_), .B(new_n2503_), .Y(new_n3129_));
  XOR2X1   g3080(.A(new_n3129_), .B(new_n3127_), .Y(\sin[11] ));
  NAND2X1  g3081(.A(new_n3081_), .B(new_n3043_), .Y(new_n3131_));
  XOR2X1   g3082(.A(new_n3081_), .B(new_n3042_), .Y(new_n3132_));
  OAI21X1  g3083(.A0(new_n3132_), .A1(new_n3037_), .B0(new_n3131_), .Y(new_n3133_));
  XOR2X1   g3084(.A(new_n3125_), .B(new_n3133_), .Y(new_n3134_));
  AND2X1   g3085(.A(new_n3134_), .B(new_n3092_), .Y(new_n3135_));
  AND2X1   g3086(.A(new_n3124_), .B(new_n3098_), .Y(new_n3136_));
  AOI21X1  g3087(.A0(new_n3125_), .A1(new_n3133_), .B0(new_n3136_), .Y(new_n3137_));
  OR4X1    g3088(.A(new_n1426_), .B(new_n195_), .C(new_n189_), .D(new_n145_), .Y(new_n3138_));
  OR2X1    g3089(.A(new_n172_), .B(new_n167_), .Y(new_n3139_));
  OR4X1    g3090(.A(new_n3139_), .B(new_n251_), .C(new_n216_), .D(new_n136_), .Y(new_n3140_));
  NOR4X1   g3091(.A(new_n3140_), .B(new_n3138_), .C(new_n2515_), .D(new_n2589_), .Y(new_n3141_));
  NAND3X1  g3092(.A(new_n3141_), .B(new_n1421_), .C(new_n1347_), .Y(new_n3142_));
  AND2X1   g3093(.A(new_n3122_), .B(new_n3105_), .Y(new_n3143_));
  INVX1    g3094(.A(new_n3099_), .Y(new_n3144_));
  AOI21X1  g3095(.A0(new_n3022_), .A1(new_n3014_), .B0(new_n3012_), .Y(new_n3145_));
  OAI21X1  g3096(.A0(new_n3047_), .A1(new_n3145_), .B0(new_n3080_), .Y(new_n3146_));
  INVX1    g3097(.A(new_n3123_), .Y(new_n3147_));
  AOI21X1  g3098(.A0(new_n3146_), .A1(new_n3144_), .B0(new_n3147_), .Y(new_n3148_));
  OR2X1    g3099(.A(new_n3148_), .B(new_n3143_), .Y(new_n3149_));
  AND2X1   g3100(.A(new_n3117_), .B(new_n3108_), .Y(new_n3150_));
  AOI21X1  g3101(.A0(new_n3121_), .A1(new_n3118_), .B0(new_n3150_), .Y(new_n3151_));
  AOI22X1  g3102(.A0(new_n2529_), .A1(new_n1721_), .B0(new_n2438_), .B1(new_n1727_), .Y(new_n3152_));
  XOR2X1   g3103(.A(new_n3152_), .B(new_n313_), .Y(new_n3153_));
  AOI22X1  g3104(.A0(new_n2286_), .A1(new_n1710_), .B0(new_n2040_), .B1(new_n1877_), .Y(new_n3154_));
  OAI21X1  g3105(.A0(new_n2371_), .A1(new_n1714_), .B0(new_n3154_), .Y(new_n3155_));
  AOI21X1  g3106(.A0(new_n2370_), .A1(new_n1707_), .B0(new_n3155_), .Y(new_n3156_));
  XOR2X1   g3107(.A(new_n3156_), .B(new_n525_), .Y(new_n3157_));
  XOR2X1   g3108(.A(new_n3157_), .B(new_n3153_), .Y(new_n3158_));
  AOI21X1  g3109(.A0(new_n3067_), .A1(new_n3109_), .B0(new_n3111_), .Y(new_n3159_));
  AOI21X1  g3110(.A0(new_n3116_), .A1(new_n3112_), .B0(new_n3159_), .Y(new_n3160_));
  NOR3X1   g3111(.A(new_n2047_), .B(new_n2044_), .C(new_n793_), .Y(new_n3161_));
  NOR3X1   g3112(.A(new_n2052_), .B(new_n2045_), .C(new_n793_), .Y(new_n3162_));
  NOR2X1   g3113(.A(new_n3162_), .B(new_n3161_), .Y(new_n3163_));
  INVX1    g3114(.A(new_n3160_), .Y(new_n3164_));
  INVX1    g3115(.A(new_n3161_), .Y(new_n3165_));
  AOI21X1  g3116(.A0(new_n3165_), .A1(new_n3164_), .B0(new_n3162_), .Y(new_n3166_));
  INVX1    g3117(.A(new_n3166_), .Y(new_n3167_));
  OAI22X1  g3118(.A0(new_n3167_), .A1(new_n3161_), .B0(new_n3163_), .B1(new_n3160_), .Y(new_n3168_));
  INVX1    g3119(.A(new_n3168_), .Y(new_n3169_));
  XOR2X1   g3120(.A(new_n3169_), .B(new_n3158_), .Y(new_n3170_));
  XOR2X1   g3121(.A(new_n3170_), .B(new_n3151_), .Y(new_n3171_));
  XOR2X1   g3122(.A(new_n3171_), .B(new_n3149_), .Y(new_n3172_));
  XOR2X1   g3123(.A(new_n3172_), .B(new_n3142_), .Y(new_n3173_));
  XOR2X1   g3124(.A(new_n3173_), .B(new_n3137_), .Y(new_n3174_));
  XOR2X1   g3125(.A(new_n3174_), .B(new_n3135_), .Y(new_n3175_));
  NAND3X1  g3126(.A(new_n3127_), .B(new_n3085_), .C(new_n3084_), .Y(new_n3176_));
  NAND2X1  g3127(.A(new_n3176_), .B(new_n2504_), .Y(new_n3177_));
  XOR2X1   g3128(.A(new_n3177_), .B(new_n3175_), .Y(\sin[12] ));
  NAND2X1  g3129(.A(new_n3124_), .B(new_n3098_), .Y(new_n3179_));
  XOR2X1   g3130(.A(new_n3124_), .B(new_n3097_), .Y(new_n3180_));
  OAI21X1  g3131(.A0(new_n3180_), .A1(new_n3094_), .B0(new_n3179_), .Y(new_n3181_));
  XOR2X1   g3132(.A(new_n3173_), .B(new_n3181_), .Y(new_n3182_));
  NAND2X1  g3133(.A(new_n3182_), .B(new_n3135_), .Y(new_n3183_));
  NOR2X1   g3134(.A(new_n3172_), .B(new_n3142_), .Y(new_n3184_));
  NAND2X1  g3135(.A(new_n3172_), .B(new_n3142_), .Y(new_n3185_));
  OAI21X1  g3136(.A0(new_n3184_), .A1(new_n3137_), .B0(new_n3185_), .Y(new_n3186_));
  OR4X1    g3137(.A(new_n710_), .B(new_n546_), .C(new_n357_), .D(new_n203_), .Y(new_n3187_));
  NOR2X1   g3138(.A(new_n205_), .B(new_n159_), .Y(new_n3188_));
  NOR3X1   g3139(.A(new_n329_), .B(new_n262_), .C(new_n208_), .Y(new_n3189_));
  AND2X1   g3140(.A(new_n3189_), .B(new_n3188_), .Y(new_n3190_));
  OR4X1    g3141(.A(new_n210_), .B(new_n192_), .C(new_n170_), .D(new_n157_), .Y(new_n3191_));
  NOR3X1   g3142(.A(new_n3191_), .B(new_n260_), .C(new_n181_), .Y(new_n3192_));
  NOR3X1   g3143(.A(new_n430_), .B(new_n287_), .C(new_n247_), .Y(new_n3193_));
  NAND4X1  g3144(.A(new_n3193_), .B(new_n3192_), .C(new_n3190_), .D(new_n2497_), .Y(new_n3194_));
  NOR3X1   g3145(.A(new_n3194_), .B(new_n3187_), .C(new_n709_), .Y(new_n3195_));
  NAND3X1  g3146(.A(new_n3195_), .B(new_n2339_), .C(new_n1557_), .Y(new_n3196_));
  INVX1    g3147(.A(new_n3196_), .Y(new_n3197_));
  NOR2X1   g3148(.A(new_n3170_), .B(new_n3151_), .Y(new_n3198_));
  INVX1    g3149(.A(new_n3143_), .Y(new_n3199_));
  OAI21X1  g3150(.A0(new_n3101_), .A1(new_n3099_), .B0(new_n3123_), .Y(new_n3200_));
  INVX1    g3151(.A(new_n3171_), .Y(new_n3201_));
  AOI21X1  g3152(.A0(new_n3200_), .A1(new_n3199_), .B0(new_n3201_), .Y(new_n3202_));
  OR2X1    g3153(.A(new_n3202_), .B(new_n3198_), .Y(new_n3203_));
  AOI22X1  g3154(.A0(new_n2368_), .A1(new_n1710_), .B0(new_n2286_), .B1(new_n1877_), .Y(new_n3204_));
  OAI21X1  g3155(.A0(new_n2442_), .A1(new_n1714_), .B0(new_n3204_), .Y(new_n3205_));
  AOI21X1  g3156(.A0(new_n2441_), .A1(new_n1707_), .B0(new_n3205_), .Y(new_n3206_));
  XOR2X1   g3157(.A(new_n3206_), .B(new_n525_), .Y(new_n3207_));
  NOR2X1   g3158(.A(new_n2047_), .B(new_n793_), .Y(new_n3208_));
  XOR2X1   g3159(.A(new_n3208_), .B(new_n312_), .Y(new_n3209_));
  NOR2X1   g3160(.A(new_n2039_), .B(new_n793_), .Y(new_n3210_));
  XOR2X1   g3161(.A(new_n3210_), .B(new_n3209_), .Y(new_n3211_));
  XOR2X1   g3162(.A(new_n3211_), .B(new_n3207_), .Y(new_n3212_));
  XOR2X1   g3163(.A(new_n3212_), .B(new_n3167_), .Y(new_n3213_));
  NOR2X1   g3164(.A(new_n3157_), .B(new_n3153_), .Y(new_n3214_));
  AOI21X1  g3165(.A0(new_n3168_), .A1(new_n3158_), .B0(new_n3214_), .Y(new_n3215_));
  XOR2X1   g3166(.A(new_n3215_), .B(new_n3213_), .Y(new_n3216_));
  XOR2X1   g3167(.A(new_n3216_), .B(new_n3203_), .Y(new_n3217_));
  XOR2X1   g3168(.A(new_n3217_), .B(new_n3197_), .Y(new_n3218_));
  NAND2X1  g3169(.A(new_n3218_), .B(new_n3186_), .Y(new_n3219_));
  AND2X1   g3170(.A(new_n3172_), .B(new_n3142_), .Y(new_n3220_));
  AOI21X1  g3171(.A0(new_n3173_), .A1(new_n3181_), .B0(new_n3220_), .Y(new_n3221_));
  NAND2X1  g3172(.A(new_n3217_), .B(new_n3196_), .Y(new_n3222_));
  OR2X1    g3173(.A(new_n3217_), .B(new_n3196_), .Y(new_n3223_));
  NAND3X1  g3174(.A(new_n3223_), .B(new_n3222_), .C(new_n3221_), .Y(new_n3224_));
  AND2X1   g3175(.A(new_n3224_), .B(new_n3219_), .Y(new_n3225_));
  XOR2X1   g3176(.A(new_n3225_), .B(new_n3183_), .Y(new_n3226_));
  NAND3X1  g3177(.A(new_n3175_), .B(new_n3128_), .C(new_n3127_), .Y(new_n3227_));
  AND2X1   g3178(.A(new_n3227_), .B(new_n2504_), .Y(new_n3228_));
  XOR2X1   g3179(.A(new_n3228_), .B(new_n3226_), .Y(\sin[13] ));
  AOI21X1  g3180(.A0(new_n3224_), .A1(new_n3219_), .B0(new_n3183_), .Y(new_n3230_));
  OAI21X1  g3181(.A0(new_n3218_), .A1(new_n3221_), .B0(new_n3222_), .Y(new_n3231_));
  OR4X1    g3182(.A(new_n317_), .B(new_n167_), .C(new_n159_), .D(new_n139_), .Y(new_n3232_));
  OR4X1    g3183(.A(new_n430_), .B(new_n379_), .C(new_n358_), .D(new_n189_), .Y(new_n3233_));
  OR4X1    g3184(.A(new_n551_), .B(new_n221_), .C(new_n188_), .D(new_n165_), .Y(new_n3234_));
  OR4X1    g3185(.A(new_n3234_), .B(new_n330_), .C(new_n293_), .D(new_n247_), .Y(new_n3235_));
  OR4X1    g3186(.A(new_n3235_), .B(new_n3233_), .C(new_n3232_), .D(new_n263_), .Y(new_n3236_));
  NOR4X1   g3187(.A(new_n3236_), .B(new_n1522_), .C(new_n922_), .D(new_n307_), .Y(new_n3237_));
  INVX1    g3188(.A(new_n3237_), .Y(new_n3238_));
  NOR2X1   g3189(.A(new_n3215_), .B(new_n3213_), .Y(new_n3239_));
  INVX1    g3190(.A(new_n3198_), .Y(new_n3240_));
  OAI21X1  g3191(.A0(new_n3148_), .A1(new_n3143_), .B0(new_n3171_), .Y(new_n3241_));
  INVX1    g3192(.A(new_n3216_), .Y(new_n3242_));
  AOI21X1  g3193(.A0(new_n3241_), .A1(new_n3240_), .B0(new_n3242_), .Y(new_n3243_));
  OR2X1    g3194(.A(new_n3243_), .B(new_n3239_), .Y(new_n3244_));
  INVX1    g3195(.A(new_n3207_), .Y(new_n3245_));
  NOR2X1   g3196(.A(new_n3212_), .B(new_n3166_), .Y(new_n3246_));
  AOI21X1  g3197(.A0(new_n3211_), .A1(new_n3245_), .B0(new_n3246_), .Y(new_n3247_));
  INVX1    g3198(.A(new_n3247_), .Y(new_n3248_));
  AND2X1   g3199(.A(new_n2286_), .B(new_n525_), .Y(new_n3249_));
  NOR3X1   g3200(.A(new_n2047_), .B(new_n793_), .C(new_n313_), .Y(new_n3250_));
  AOI21X1  g3201(.A0(new_n3210_), .A1(new_n3209_), .B0(new_n3250_), .Y(new_n3251_));
  XOR2X1   g3202(.A(new_n3251_), .B(new_n3249_), .Y(new_n3252_));
  OAI22X1  g3203(.A0(new_n2442_), .A1(new_n1711_), .B0(new_n2371_), .B1(new_n1785_), .Y(new_n3253_));
  AOI21X1  g3204(.A0(new_n2530_), .A1(new_n1707_), .B0(new_n3253_), .Y(new_n3254_));
  XOR2X1   g3205(.A(new_n3254_), .B(new_n793_), .Y(new_n3255_));
  XOR2X1   g3206(.A(new_n3255_), .B(new_n3252_), .Y(new_n3256_));
  XOR2X1   g3207(.A(new_n3256_), .B(new_n3248_), .Y(new_n3257_));
  XOR2X1   g3208(.A(new_n3257_), .B(new_n3244_), .Y(new_n3258_));
  XOR2X1   g3209(.A(new_n3258_), .B(new_n3238_), .Y(new_n3259_));
  XOR2X1   g3210(.A(new_n3259_), .B(new_n3231_), .Y(new_n3260_));
  INVX1    g3211(.A(new_n3260_), .Y(new_n3261_));
  XOR2X1   g3212(.A(new_n3261_), .B(new_n3230_), .Y(new_n3262_));
  OAI21X1  g3213(.A0(new_n3227_), .A1(new_n3226_), .B0(new_n2504_), .Y(new_n3263_));
  XOR2X1   g3214(.A(new_n3263_), .B(new_n3262_), .Y(\sin[14] ));
  AND2X1   g3215(.A(new_n3260_), .B(new_n3230_), .Y(new_n3265_));
  AND2X1   g3216(.A(new_n3217_), .B(new_n3196_), .Y(new_n3266_));
  AOI21X1  g3217(.A0(new_n3223_), .A1(new_n3186_), .B0(new_n3266_), .Y(new_n3267_));
  NAND2X1  g3218(.A(new_n3258_), .B(new_n3238_), .Y(new_n3268_));
  XOR2X1   g3219(.A(new_n3258_), .B(new_n3237_), .Y(new_n3269_));
  OAI21X1  g3220(.A0(new_n3269_), .A1(new_n3267_), .B0(new_n3268_), .Y(new_n3270_));
  OR4X1    g3221(.A(new_n732_), .B(new_n398_), .C(new_n385_), .D(new_n207_), .Y(new_n3271_));
  OR4X1    g3222(.A(new_n293_), .B(new_n283_), .C(new_n269_), .D(new_n110_), .Y(new_n3272_));
  OR4X1    g3223(.A(new_n603_), .B(new_n2790_), .C(new_n221_), .D(new_n132_), .Y(new_n3273_));
  OR4X1    g3224(.A(new_n3273_), .B(new_n3272_), .C(new_n3140_), .D(new_n714_), .Y(new_n3274_));
  NOR3X1   g3225(.A(new_n3274_), .B(new_n3271_), .C(new_n1428_), .Y(new_n3275_));
  AOI22X1  g3226(.A0(new_n2529_), .A1(new_n1707_), .B0(new_n2438_), .B1(new_n1877_), .Y(new_n3276_));
  XOR2X1   g3227(.A(new_n3276_), .B(new_n525_), .Y(new_n3277_));
  AND2X1   g3228(.A(new_n2369_), .B(new_n525_), .Y(new_n3278_));
  XOR2X1   g3229(.A(new_n3278_), .B(new_n3277_), .Y(new_n3279_));
  INVX1    g3230(.A(new_n3279_), .Y(new_n3280_));
  NOR2X1   g3231(.A(new_n3251_), .B(new_n3249_), .Y(new_n3281_));
  AOI21X1  g3232(.A0(new_n3255_), .A1(new_n3252_), .B0(new_n3281_), .Y(new_n3282_));
  XOR2X1   g3233(.A(new_n3282_), .B(new_n3280_), .Y(new_n3283_));
  INVX1    g3234(.A(new_n3283_), .Y(new_n3284_));
  AND2X1   g3235(.A(new_n3256_), .B(new_n3248_), .Y(new_n3285_));
  INVX1    g3236(.A(new_n3285_), .Y(new_n3286_));
  OAI21X1  g3237(.A0(new_n3243_), .A1(new_n3239_), .B0(new_n3257_), .Y(new_n3287_));
  AND2X1   g3238(.A(new_n3287_), .B(new_n3286_), .Y(new_n3288_));
  XOR2X1   g3239(.A(new_n3288_), .B(new_n3284_), .Y(new_n3289_));
  XOR2X1   g3240(.A(new_n3289_), .B(new_n3275_), .Y(new_n3290_));
  AND2X1   g3241(.A(new_n3290_), .B(new_n3270_), .Y(new_n3291_));
  INVX1    g3242(.A(new_n3275_), .Y(new_n3292_));
  AND2X1   g3243(.A(new_n3289_), .B(new_n3292_), .Y(new_n3293_));
  NOR2X1   g3244(.A(new_n3289_), .B(new_n3292_), .Y(new_n3294_));
  NOR3X1   g3245(.A(new_n3294_), .B(new_n3293_), .C(new_n3270_), .Y(new_n3295_));
  OR2X1    g3246(.A(new_n3295_), .B(new_n3291_), .Y(new_n3296_));
  XOR2X1   g3247(.A(new_n3296_), .B(new_n3265_), .Y(new_n3297_));
  NOR2X1   g3248(.A(new_n3227_), .B(new_n3226_), .Y(new_n3298_));
  AOI21X1  g3249(.A0(new_n3298_), .A1(new_n3262_), .B0(new_n2503_), .Y(new_n3299_));
  XOR2X1   g3250(.A(new_n3299_), .B(new_n3297_), .Y(\sin[15] ));
  OAI21X1  g3251(.A0(new_n3295_), .A1(new_n3291_), .B0(new_n3265_), .Y(new_n3301_));
  AND2X1   g3252(.A(new_n3258_), .B(new_n3238_), .Y(new_n3302_));
  AOI21X1  g3253(.A0(new_n3259_), .A1(new_n3231_), .B0(new_n3302_), .Y(new_n3303_));
  NAND2X1  g3254(.A(new_n3289_), .B(new_n3292_), .Y(new_n3304_));
  OAI21X1  g3255(.A0(new_n3294_), .A1(new_n3303_), .B0(new_n3304_), .Y(new_n3305_));
  OR4X1    g3256(.A(new_n249_), .B(new_n165_), .C(new_n155_), .D(new_n132_), .Y(new_n3306_));
  OR4X1    g3257(.A(new_n3306_), .B(new_n315_), .C(new_n337_), .D(new_n213_), .Y(new_n3307_));
  NAND4X1  g3258(.A(new_n3189_), .B(new_n3188_), .C(new_n117_), .D(new_n98_), .Y(new_n3308_));
  OR4X1    g3259(.A(new_n3308_), .B(new_n3307_), .C(new_n1359_), .D(new_n293_), .Y(new_n3309_));
  NOR4X1   g3260(.A(new_n3309_), .B(new_n2336_), .C(new_n1386_), .D(new_n463_), .Y(new_n3310_));
  INVX1    g3261(.A(new_n3310_), .Y(new_n3311_));
  NOR2X1   g3262(.A(new_n3282_), .B(new_n3280_), .Y(new_n3312_));
  INVX1    g3263(.A(new_n3312_), .Y(new_n3313_));
  INVX1    g3264(.A(new_n3239_), .Y(new_n3314_));
  OAI21X1  g3265(.A0(new_n3202_), .A1(new_n3198_), .B0(new_n3216_), .Y(new_n3315_));
  INVX1    g3266(.A(new_n3257_), .Y(new_n3316_));
  AOI21X1  g3267(.A0(new_n3315_), .A1(new_n3314_), .B0(new_n3316_), .Y(new_n3317_));
  OAI21X1  g3268(.A0(new_n3317_), .A1(new_n3285_), .B0(new_n3283_), .Y(new_n3318_));
  NAND3X1  g3269(.A(new_n2368_), .B(new_n2738_), .C(new_n525_), .Y(new_n3319_));
  OAI21X1  g3270(.A0(new_n3278_), .A1(new_n3277_), .B0(new_n3319_), .Y(new_n3320_));
  AOI21X1  g3271(.A0(new_n3318_), .A1(new_n3313_), .B0(new_n3320_), .Y(new_n3321_));
  AOI21X1  g3272(.A0(new_n3287_), .A1(new_n3286_), .B0(new_n3284_), .Y(new_n3322_));
  INVX1    g3273(.A(new_n3320_), .Y(new_n3323_));
  NOR3X1   g3274(.A(new_n3323_), .B(new_n3322_), .C(new_n3312_), .Y(new_n3324_));
  NAND2X1  g3275(.A(new_n3249_), .B(new_n2442_), .Y(new_n3325_));
  AOI21X1  g3276(.A0(new_n2438_), .A1(new_n2738_), .B0(new_n793_), .Y(new_n3326_));
  AND2X1   g3277(.A(new_n3326_), .B(new_n3325_), .Y(new_n3327_));
  NOR3X1   g3278(.A(new_n3327_), .B(new_n3324_), .C(new_n3321_), .Y(new_n3328_));
  OAI21X1  g3279(.A0(new_n3322_), .A1(new_n3312_), .B0(new_n3323_), .Y(new_n3329_));
  NAND3X1  g3280(.A(new_n3320_), .B(new_n3318_), .C(new_n3313_), .Y(new_n3330_));
  INVX1    g3281(.A(new_n3327_), .Y(new_n3331_));
  AOI21X1  g3282(.A0(new_n3330_), .A1(new_n3329_), .B0(new_n3331_), .Y(new_n3332_));
  NOR3X1   g3283(.A(new_n3332_), .B(new_n3328_), .C(new_n3311_), .Y(new_n3333_));
  NAND3X1  g3284(.A(new_n3331_), .B(new_n3330_), .C(new_n3329_), .Y(new_n3334_));
  OAI21X1  g3285(.A0(new_n3324_), .A1(new_n3321_), .B0(new_n3327_), .Y(new_n3335_));
  AOI21X1  g3286(.A0(new_n3335_), .A1(new_n3334_), .B0(new_n3310_), .Y(new_n3336_));
  OAI21X1  g3287(.A0(new_n3336_), .A1(new_n3333_), .B0(new_n3305_), .Y(new_n3337_));
  OR2X1    g3288(.A(new_n3289_), .B(new_n3292_), .Y(new_n3338_));
  AOI21X1  g3289(.A0(new_n3338_), .A1(new_n3270_), .B0(new_n3293_), .Y(new_n3339_));
  NAND3X1  g3290(.A(new_n3335_), .B(new_n3334_), .C(new_n3310_), .Y(new_n3340_));
  OAI21X1  g3291(.A0(new_n3332_), .A1(new_n3328_), .B0(new_n3311_), .Y(new_n3341_));
  NAND3X1  g3292(.A(new_n3341_), .B(new_n3340_), .C(new_n3339_), .Y(new_n3342_));
  AND2X1   g3293(.A(new_n3342_), .B(new_n3337_), .Y(new_n3343_));
  XOR2X1   g3294(.A(new_n3343_), .B(new_n3301_), .Y(new_n3344_));
  INVX1    g3295(.A(new_n3344_), .Y(new_n3345_));
  NAND2X1  g3296(.A(new_n3298_), .B(new_n3262_), .Y(new_n3346_));
  OAI21X1  g3297(.A0(new_n3346_), .A1(new_n3297_), .B0(new_n2504_), .Y(new_n3347_));
  XOR2X1   g3298(.A(new_n3347_), .B(new_n3345_), .Y(\sin[16] ));
  AOI21X1  g3299(.A0(new_n3342_), .A1(new_n3337_), .B0(new_n3301_), .Y(new_n3349_));
  AOI21X1  g3300(.A0(new_n3340_), .A1(new_n3305_), .B0(new_n3336_), .Y(new_n3350_));
  OR4X1    g3301(.A(new_n259_), .B(new_n256_), .C(new_n174_), .D(new_n127_), .Y(new_n3351_));
  NOR4X1   g3302(.A(new_n3351_), .B(new_n216_), .C(new_n212_), .D(new_n195_), .Y(new_n3352_));
  NOR4X1   g3303(.A(new_n442_), .B(new_n346_), .C(new_n280_), .D(new_n130_), .Y(new_n3353_));
  NAND2X1  g3304(.A(new_n3353_), .B(new_n3352_), .Y(new_n3354_));
  NOR4X1   g3305(.A(new_n3354_), .B(new_n2025_), .C(new_n570_), .D(new_n187_), .Y(new_n3355_));
  XOR2X1   g3306(.A(new_n3355_), .B(new_n3350_), .Y(new_n3356_));
  XOR2X1   g3307(.A(new_n3356_), .B(new_n3349_), .Y(new_n3357_));
  NOR3X1   g3308(.A(new_n3344_), .B(new_n3346_), .C(new_n3297_), .Y(new_n3358_));
  NOR2X1   g3309(.A(new_n3358_), .B(new_n2503_), .Y(new_n3359_));
  XOR2X1   g3310(.A(new_n3359_), .B(new_n3357_), .Y(\sin[17] ));
  AND2X1   g3311(.A(new_n3356_), .B(new_n3349_), .Y(new_n3361_));
  OAI21X1  g3312(.A0(new_n3333_), .A1(new_n3339_), .B0(new_n3341_), .Y(new_n3362_));
  INVX1    g3313(.A(new_n3355_), .Y(new_n3363_));
  NOR3X1   g3314(.A(new_n304_), .B(new_n141_), .C(new_n113_), .Y(new_n3364_));
  NAND3X1  g3315(.A(new_n3364_), .B(new_n215_), .C(new_n285_), .Y(new_n3365_));
  OR4X1    g3316(.A(new_n3365_), .B(new_n607_), .C(new_n1442_), .D(new_n385_), .Y(new_n3366_));
  OR4X1    g3317(.A(new_n3366_), .B(new_n1553_), .C(new_n718_), .D(new_n707_), .Y(new_n3367_));
  NOR4X1   g3318(.A(new_n3367_), .B(new_n2321_), .C(new_n558_), .D(new_n201_), .Y(new_n3368_));
  INVX1    g3319(.A(new_n3368_), .Y(new_n3369_));
  NAND3X1  g3320(.A(new_n3369_), .B(new_n3363_), .C(new_n3362_), .Y(new_n3370_));
  OAI21X1  g3321(.A0(new_n3355_), .A1(new_n3350_), .B0(new_n3368_), .Y(new_n3371_));
  AND2X1   g3322(.A(new_n3371_), .B(new_n3370_), .Y(new_n3372_));
  NAND3X1  g3323(.A(new_n3371_), .B(new_n3356_), .C(new_n3349_), .Y(new_n3373_));
  OAI21X1  g3324(.A0(new_n3372_), .A1(new_n3361_), .B0(new_n3373_), .Y(new_n3374_));
  NOR4X1   g3325(.A(new_n3357_), .B(new_n3344_), .C(new_n3346_), .D(new_n3297_), .Y(new_n3375_));
  OR2X1    g3326(.A(new_n3375_), .B(new_n2503_), .Y(new_n3376_));
  XOR2X1   g3327(.A(new_n3376_), .B(new_n3374_), .Y(\sin[18] ));
  NOR3X1   g3328(.A(new_n3368_), .B(new_n3355_), .C(new_n3350_), .Y(new_n3378_));
  OR4X1    g3329(.A(new_n214_), .B(new_n196_), .C(new_n193_), .D(new_n185_), .Y(new_n3379_));
  NOR3X1   g3330(.A(new_n292_), .B(new_n256_), .C(new_n213_), .Y(new_n3380_));
  NAND2X1  g3331(.A(new_n3380_), .B(new_n2719_), .Y(new_n3381_));
  OR4X1    g3332(.A(new_n3381_), .B(new_n3379_), .C(new_n1685_), .D(new_n296_), .Y(new_n3382_));
  NOR3X1   g3333(.A(new_n3382_), .B(new_n3271_), .C(new_n475_), .Y(new_n3383_));
  XOR2X1   g3334(.A(new_n3383_), .B(new_n3378_), .Y(new_n3384_));
  XOR2X1   g3335(.A(new_n3384_), .B(new_n3373_), .Y(new_n3385_));
  AOI21X1  g3336(.A0(new_n3375_), .A1(new_n3374_), .B0(new_n2503_), .Y(new_n3386_));
  XOR2X1   g3337(.A(new_n3386_), .B(new_n3385_), .Y(\sin[19] ));
  OR4X1    g3338(.A(new_n3383_), .B(new_n3368_), .C(new_n3355_), .D(new_n3350_), .Y(new_n3388_));
  OR4X1    g3339(.A(new_n346_), .B(new_n221_), .C(new_n173_), .D(new_n172_), .Y(new_n3389_));
  OR4X1    g3340(.A(new_n159_), .B(new_n149_), .C(new_n147_), .D(new_n134_), .Y(new_n3390_));
  OR4X1    g3341(.A(new_n3390_), .B(new_n294_), .C(new_n271_), .D(new_n113_), .Y(new_n3391_));
  OR4X1    g3342(.A(new_n3391_), .B(new_n3389_), .C(new_n365_), .D(new_n334_), .Y(new_n3392_));
  NOR4X1   g3343(.A(new_n3392_), .B(new_n2925_), .C(new_n496_), .D(new_n201_), .Y(new_n3393_));
  NOR2X1   g3344(.A(new_n3393_), .B(new_n3388_), .Y(new_n3394_));
  AND2X1   g3345(.A(new_n3393_), .B(new_n3388_), .Y(new_n3395_));
  OAI22X1  g3346(.A0(new_n3395_), .A1(new_n3394_), .B0(new_n3384_), .B1(new_n3373_), .Y(new_n3396_));
  XOR2X1   g3347(.A(new_n3383_), .B(new_n3370_), .Y(new_n3397_));
  NAND2X1  g3348(.A(new_n3393_), .B(new_n3388_), .Y(new_n3398_));
  NAND4X1  g3349(.A(new_n3398_), .B(new_n3397_), .C(new_n3371_), .D(new_n3361_), .Y(new_n3399_));
  AND2X1   g3350(.A(new_n3399_), .B(new_n3396_), .Y(new_n3400_));
  NAND2X1  g3351(.A(new_n3375_), .B(new_n3374_), .Y(new_n3401_));
  OR2X1    g3352(.A(new_n3401_), .B(new_n3385_), .Y(new_n3402_));
  AND2X1   g3353(.A(new_n3402_), .B(new_n2504_), .Y(new_n3403_));
  XOR2X1   g3354(.A(new_n3403_), .B(new_n3400_), .Y(\sin[20] ));
  OR4X1    g3355(.A(new_n326_), .B(new_n324_), .C(new_n329_), .D(new_n247_), .Y(new_n3405_));
  NOR4X1   g3356(.A(new_n3405_), .B(new_n2281_), .C(new_n400_), .D(new_n384_), .Y(new_n3406_));
  XOR2X1   g3357(.A(new_n3406_), .B(new_n3394_), .Y(new_n3407_));
  XOR2X1   g3358(.A(new_n3407_), .B(new_n3399_), .Y(new_n3408_));
  INVX1    g3359(.A(new_n3408_), .Y(new_n3409_));
  OAI21X1  g3360(.A0(new_n3402_), .A1(new_n3400_), .B0(new_n2504_), .Y(new_n3410_));
  XOR2X1   g3361(.A(new_n3410_), .B(new_n3409_), .Y(\sin[21] ));
  NOR2X1   g3362(.A(new_n3407_), .B(new_n3399_), .Y(new_n3412_));
  OR4X1    g3363(.A(new_n3406_), .B(new_n3393_), .C(new_n3383_), .D(new_n3370_), .Y(new_n3413_));
  NOR4X1   g3364(.A(new_n400_), .B(new_n384_), .C(new_n361_), .D(new_n345_), .Y(new_n3414_));
  AND2X1   g3365(.A(new_n3414_), .B(new_n3413_), .Y(new_n3415_));
  XOR2X1   g3366(.A(new_n3414_), .B(new_n3413_), .Y(new_n3416_));
  MX2X1    g3367(.A(new_n3416_), .B(new_n3415_), .S0(new_n3412_), .Y(new_n3417_));
  OR4X1    g3368(.A(new_n3408_), .B(new_n3400_), .C(new_n3401_), .D(new_n3385_), .Y(new_n3418_));
  AND2X1   g3369(.A(new_n3418_), .B(new_n2504_), .Y(new_n3419_));
  XOR2X1   g3370(.A(new_n3419_), .B(new_n3417_), .Y(\sin[22] ));
  NOR4X1   g3371(.A(new_n3414_), .B(new_n3406_), .C(new_n3393_), .D(new_n3388_), .Y(new_n3421_));
  NOR3X1   g3372(.A(new_n3415_), .B(new_n3407_), .C(new_n3399_), .Y(new_n3422_));
  XOR2X1   g3373(.A(new_n3422_), .B(new_n3421_), .Y(new_n3423_));
  OAI21X1  g3374(.A0(new_n3418_), .A1(new_n3417_), .B0(new_n2504_), .Y(new_n3424_));
  NOR3X1   g3375(.A(new_n75_), .B(\a[22] ), .C(\a[21] ), .Y(new_n3425_));
  AOI21X1  g3376(.A0(new_n3424_), .A1(new_n3423_), .B0(new_n3425_), .Y(new_n3426_));
  OAI21X1  g3377(.A0(new_n3424_), .A1(new_n3423_), .B0(new_n3426_), .Y(\sin[23] ));
  OR4X1    g3378(.A(new_n3414_), .B(new_n3407_), .C(new_n3413_), .D(new_n3399_), .Y(new_n3428_));
  OAI21X1  g3379(.A0(new_n3418_), .A1(new_n3417_), .B0(new_n3428_), .Y(new_n3429_));
  OR2X1    g3380(.A(new_n3422_), .B(new_n3421_), .Y(new_n3430_));
  NOR2X1   g3381(.A(new_n3418_), .B(new_n3417_), .Y(new_n3431_));
  AOI21X1  g3382(.A0(new_n3431_), .A1(new_n3430_), .B0(new_n3425_), .Y(new_n3432_));
  AOI21X1  g3383(.A0(new_n3432_), .A1(new_n3429_), .B0(new_n2503_), .Y(\sin[24] ));
endmodule


