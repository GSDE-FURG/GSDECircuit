//Converted to Combinational (Partial output: n676) , Module name: s9234_n676
module s9234_n676 ( g1, g2, g6, g24, g28, g693, g677, g683, g684, g41, g541, g682, g681, g676, g702, g699, g688, g536, g689, g685, g698, g516, g236, g465, g48, g230, g512, g520, g242, g524, g532, g278, g276, g277, g281, g279, g280, g212, g500, g224, g508, g528, g254, g504, g218, g248, g260, g206, g204, g205, g207, g208, g209, g1, g10, g18, g14, n676 );
input g1, g2, g6, g24, g28, g693, g677, g683, g684, g41, g541, g682, g681, g676, g702, g699, g688, g536, g689, g685, g698, g516, g236, g465, g48, g230, g512, g520, g242, g524, g532, g278, g276, g277, g281, g279, g280, g212, g500, g224, g508, g528, g254, g504, g218, g248, g260, g206, g204, g205, g207, g208, g209, g1, g10, g18, g14;
output n676;
wire n1011_1, n1497, n1010, n1007, n1009, n1349, n1496, n798, n826_1, n727, n1005, n1006_1, n1008, n1213, n991_1, n1495, n724, n726_1, n758, n789, n939, n990, n978, n981_1, n984, n1494, n1122, n870, n716_1, n723, n725, n989, n979, n980, n982, n983, n964, n869, n866_1, n867, n868, n719, n722, n988, n985, n986_1, n987, n793, n955, n963, n960, n961_1, n962, n717, n718, n720, n721_1;
MX2X1    g0788(.A(n1497), .B(g693), .S0(n1011_1), .Y(n676));
NOR4X1   g0302(.A(n1009), .B(n1007), .C(g677), .D(n1010), .Y(n1011_1));
NAND2X1  g0787(.A(n1496), .B(n1349), .Y(n1497));
NAND4X1  g0301(.A(n826_1), .B(g684), .C(n798), .D(g683), .Y(n1010));
OR4X1    g0298(.A(n1006_1), .B(g41), .C(n1005), .D(n727), .Y(n1007));
INVX1    g0300(.A(n1008), .Y(n1009));
INVX1    g0640(.A(g541), .Y(n1349));
NAND3X1  g0786(.A(n1495), .B(n991_1), .C(n1213), .Y(n1496));
INVX1    g0090(.A(g682), .Y(n798));
INVX1    g0118(.A(g681), .Y(n826_1));
OAI21X1  g0019(.A0(n726_1), .A1(n724), .B0(g676), .Y(n727));
INVX1    g0296(.A(g702), .Y(n1005));
INVX1    g0297(.A(g699), .Y(n1006_1));
NOR4X1   g0299(.A(n939), .B(n789), .C(n758), .D(g688), .Y(n1008));
INVX1    g0504(.A(g536), .Y(n1213));
NOR4X1   g0282(.A(n984), .B(n981_1), .C(n978), .D(n990), .Y(n991_1));
MX2X1    g0785(.A(n870), .B(n1122), .S0(n1494), .Y(n1495));
AND2X1   g0016(.A(n723), .B(n716_1), .Y(n724));
OAI21X1  g0018(.A0(n723), .A1(n716_1), .B0(n725), .Y(n726_1));
INVX1    g0050(.A(g689), .Y(n758));
INVX1    g0081(.A(g685), .Y(n789));
INVX1    g0230(.A(g698), .Y(n939));
INVX1    g0281(.A(n989), .Y(n990));
XOR2X1   g0269(.A(g236), .B(g516), .Y(n978));
OR2X1    g0272(.A(n980), .B(n979), .Y(n981_1));
NAND2X1  g0275(.A(n983), .B(n982), .Y(n984));
INVX1    g0784(.A(g465), .Y(n1494));
INVX1    g0413(.A(n964), .Y(n1122));
NOR4X1   g0162(.A(n868), .B(n867), .C(n866_1), .D(n869), .Y(n870));
INVX1    g0008(.A(g48), .Y(n716_1));
XOR2X1   g0015(.A(n722), .B(n719), .Y(n723));
INVX1    g0017(.A(g41), .Y(n725));
NOR4X1   g0280(.A(n987), .B(n986_1), .C(n985), .D(n988), .Y(n989));
XOR2X1   g0270(.A(g512), .B(g230), .Y(n979));
XOR2X1   g0271(.A(g242), .B(g520), .Y(n980));
XOR2X1   g0273(.A(g524), .B(n793), .Y(n982));
XOR2X1   g0274(.A(g532), .B(n955), .Y(n983));
OR4X1    g0255(.A(n962), .B(n961_1), .C(n960), .D(n963), .Y(n964));
NAND3X1  g0161(.A(g277), .B(g276), .C(g278), .Y(n869));
INVX1    g0158(.A(g281), .Y(n866_1));
INVX1    g0159(.A(g279), .Y(n867));
INVX1    g0160(.A(g280), .Y(n868));
XOR2X1   g0011(.A(n718), .B(n717), .Y(n719));
XOR2X1   g0014(.A(n721_1), .B(n720), .Y(n722));
XOR2X1   g0279(.A(g500), .B(g212), .Y(n988));
XOR2X1   g0276(.A(g508), .B(g224), .Y(n985));
XOR2X1   g0277(.A(g254), .B(g528), .Y(n986_1));
XOR2X1   g0278(.A(g218), .B(g504), .Y(n987));
INVX1    g0085(.A(g248), .Y(n793));
INVX1    g0246(.A(g260), .Y(n955));
NAND3X1  g0254(.A(g205), .B(g204), .C(g206), .Y(n963));
INVX1    g0251(.A(g207), .Y(n960));
INVX1    g0252(.A(g208), .Y(n961_1));
INVX1    g0253(.A(g209), .Y(n962));
XOR2X1   g0009(.A(g1), .B(g2), .Y(n717));
XOR2X1   g0010(.A(g10), .B(g6), .Y(n718));
XOR2X1   g0012(.A(g14), .B(g18), .Y(n720));
XOR2X1   g0013(.A(g28), .B(g24), .Y(n721_1));

endmodule
