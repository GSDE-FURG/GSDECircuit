//Converted to Combinational , Module name: s9234 , Timestamp: 2018-12-03T15:51:03.319453 
module s9234 ( g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23, g678, g332, g123, g207, g695, g461, g18, g292, g331, g689, g24, g465, g84, g291, g676, g622, g117, g278, g128, g598, g554, g496, g179, g48, g590, g551, g682, g606, g188, g646, g327, g361, g289, g398, g684, g619, g208, g248, g390, g625, g681, g437, g276, g323, g224, g685, g157, g282, g697, g206, g449, g118, g528, g284, g426, g634, g669, g520, g281, g175, g631, g693, g337, g457, g486, g471, g328, g285, g418, g402, g297, g212, g410, g430, g662, g453, g269, g574, g441, g664, g349, g211, g586, g571, g326, g698, g654, g293, g690, g445, g374, g687, g357, g386, g504, g665, g166, g541, g74, g338, g696, g516, g536, g683, g353, g545, g254, g341, g290, g287, g336, g345, g628, g679, g688, g283, g613, g14, g680, g143, g672, g667, g366, g279, g492, g170, g686, g288, g638, g602, g642, g280, g663, g610, g148, g209, g675, g478, g122, g594, g286, g489, g616, g79, g218, g242, g578, g184, g119, g668, g139, g422, g210, g394, g230, g204, g658, g650, g378, g508, g548, g370, g406, g236, g500, g205, g197, g666, g114, g524, g260, g111, g131, g677, g582, g485, g699, g193, g135, g382, g414, g434, g266, g152, g692, g277, g127, g161, g512, g532, g694, g691, g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102, g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098, n151, n156, n161, n166, n171, n176, n181, n186, n191, n196, n201, n206, n211, n216, n221, n226, n231, n236, n241, n246, n251, n256, n261, n266, n271, n276, n281, n286, n291, n296, n301, n306, n311, n316, n321, n326, n331, n336, n341, n346, n351, n356, n361, n366, n371, n376, n381, n386, n391, n396, n401, n406, n411, n416, n421, n426, n431, n436, n441, n446, n451, n456, n461, n466, n471, n476, n481, n486, n491, n496, n501, n506, n511, n516, n521, n526, n531, n536, n541, n546, n551, n556, n561, n566, n571, n576, n581, n586, n591, n596, n601, n606, n611, n616, n621, n626, n631, n636, n641, n646, n651, n656, n661, n666, n671, n676, n681, n686, n691, n696, n701, n706, n711, n716, n721, n726, n731, n736, n741, n746, n751, n756, n761, n766, n771, n776, n781, n786, n791, n796, n801, n806, n811, n816, n821, n826, n831, n836, n841, n846, n851, n856, n861, n866, n871, n876, n881, n886, n891, n896, n901, n906, n911, n916, n921, n926, n931, n936, n941, n946, n951, n956, n961, n966, n971, n976, n981, n986, n991, n996, n1001, n1006, n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201 );
input g43, g59, g54, g49, g64, g69, g3, g7, g11, g15, g25, g19, g33, g29, g28, g6, g10, g2, g1, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23, g678, g332, g123, g207, g695, g461, g18, g292, g331, g689, g24, g465, g84, g291, g676, g622, g117, g278, g128, g598, g554, g496, g179, g48, g590, g551, g682, g606, g188, g646, g327, g361, g289, g398, g684, g619, g208, g248, g390, g625, g681, g437, g276, g323, g224, g685, g157, g282, g697, g206, g449, g118, g528, g284, g426, g634, g669, g520, g281, g175, g631, g693, g337, g457, g486, g471, g328, g285, g418, g402, g297, g212, g410, g430, g662, g453, g269, g574, g441, g664, g349, g211, g586, g571, g326, g698, g654, g293, g690, g445, g374, g687, g357, g386, g504, g665, g166, g541, g74, g338, g696, g516, g536, g683, g353, g545, g254, g341, g290, g287, g336, g345, g628, g679, g688, g283, g613, g14, g680, g143, g672, g667, g366, g279, g492, g170, g686, g288, g638, g602, g642, g280, g663, g610, g148, g209, g675, g478, g122, g594, g286, g489, g616, g79, g218, g242, g578, g184, g119, g668, g139, g422, g210, g394, g230, g204, g658, g650, g378, g508, g548, g370, g406, g236, g500, g205, g197, g666, g114, g524, g260, g111, g131, g677, g582, g485, g699, g193, g135, g382, g414, g434, g266, g152, g692, g277, g127, g161, g512, g532, g694, g691;
output g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102, g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098, n151, n156, n161, n166, n171, n176, n181, n186, n191, n196, n201, n206, n211, n216, n221, n226, n231, n236, n241, n246, n251, n256, n261, n266, n271, n276, n281, n286, n291, n296, n301, n306, n311, n316, n321, n326, n331, n336, n341, n346, n351, n356, n361, n366, n371, n376, n381, n386, n391, n396, n401, n406, n411, n416, n421, n426, n431, n436, n441, n446, n451, n456, n461, n466, n471, n476, n481, n486, n491, n496, n501, n506, n511, n516, n521, n526, n531, n536, n541, n546, n551, n556, n561, n566, n571, n576, n581, n586, n591, n596, n601, n606, n611, n616, n621, n626, n631, n636, n641, n646, n651, n656, n661, n666, n671, n676, n681, n686, n691, n696, n701, n706, n711, n716, n721, n726, n731, n736, n741, n746, n751, n756, n761, n766, n771, n776, n781, n786, n791, n796, n801, n806, n811, n816, n821, n826, n831, n836, n841, n846, n851, n856, n861, n866, n871, n876, n881, n886, n891, n896, n901, n906, n911, n916, n921, n926, n931, n936, n941, n946, n951, n956, n961, n966, n971, n976, n981, n986, n991, n996, n1001, n1006, n1011, n1016, n1021, n1026, n1031, n1036, n1041, n1046, n1051, n1056, n1061, n1066, n1071, n1076, n1081, n1086, n1091, n1096, n1101, n1106, n1111, n1116, n1121, n1126, n1131, n1136, n1141, n1146, n1151, n1156, n1161, n1166, n1171, n1176, n1181, n1186, n1191, n1196, n1201;
wire n708, n710, n711_1, n714, n715, n716_1, n717, n718, n719, n720, n721_1, n722, n723, n724, n725, n726_1, n727, n729, n730, n731_1, n732, n733, n734, n735, n736_1, n748, n749, n750, n751_1, n752, n753, n754, n755, n756_1, n757, n758, n759, n760, n761_1, n762, n763, n764, n765, n766_1, n767, n768, n769, n770, n771_1, n772, n773, n774, n775, n776_1, n777, n778, n780, n781_1, n782, n783, n784, n785, n786_1, n787, n788, n789, n790, n791_1, n792, n793, n794, n795, n796_1, n797, n798, n799, n800, n801_1, n802, n803, n804, n805, n806_1, n807, n808, n809, n810, n811_1, n812, n813, n814, n815, n816_1, n817, n818, n819, n820, n821_1, n822, n823, n824, n825, n826_1, n827, n828, n829, n830, n831_1, n833, n834, n835, n836_1, n837, n838, n839, n841_1, n842, n843, n844, n845, n846_1, n847, n848, n849, n850, n851_1, n852, n853, n854, n855, n856_1, n857, n858, n859, n860, n861_1, n862, n863, n864, n865, n866_1, n867, n868, n869, n870, n871_1, n872, n873, n874, n875, n876_1, n877, n878, n879, n880, n881_1, n882, n883, n884, n885, n886_1, n887, n888, n889, n890, n891_1, n892, n893, n894, n895, n896_1, n897, n898, n899, n900, n901_1, n902, n903, n904, n905, n906_1, n907, n908, n909, n910, n911_1, n912, n913, n914, n915, n916_1, n917, n918, n919, n920, n921_1, n922, n923, n924, n926_1, n927, n928, n929, n930, n931_1, n932, n933, n934, n935, n936_1, n937, n938, n939, n940, n941_1, n942, n943, n944, n945, n946_1, n947, n948, n949, n950, n951_1, n952, n953, n954, n955, n956_1, n957, n958, n960, n961_1, n962, n963, n964, n965, n966_1, n967, n968, n969, n970, n971_1, n972, n973, n974, n975, n976_1, n978, n979, n980, n981_1, n982, n983, n984, n985, n986_1, n987, n988, n989, n990, n991_1, n992, n993, n995, n996_1, n997, n999, n1000, n1002, n1003, n1005, n1006_1, n1007, n1008, n1009, n1010, n1011_1, n1013, n1014, n1015, n1016_1, n1017, n1018, n1019, n1020, n1021_1, n1022, n1023, n1024, n1025, n1026_1, n1027, n1028, n1029, n1030, n1031_1, n1032, n1033, n1034, n1035, n1036_1, n1037, n1038, n1039, n1040, n1041_1, n1042, n1043, n1044, n1045, n1046_1, n1047, n1048, n1049, n1050, n1051_1, n1052, n1053, n1054, n1055, n1057, n1058, n1059, n1060, n1061_1, n1062, n1064, n1065, n1066_1, n1067, n1068, n1069, n1071_1, n1073, n1074, n1075, n1076_1, n1078, n1079, n1080, n1082, n1085, n1086_1, n1087, n1088, n1089, n1090, n1091_1, n1092, n1093, n1094, n1095, n1096_1, n1097, n1098, n1099, n1100, n1101_1, n1102, n1103, n1104, n1105, n1106_1, n1107, n1108, n1109, n1110, n1111_1, n1112, n1113, n1114, n1115, n1116_1, n1117, n1118, n1119, n1120, n1121_1, n1122, n1123, n1124, n1126_1, n1127, n1128, n1129, n1130, n1131_1, n1132, n1133, n1134, n1135, n1136_1, n1137, n1138, n1139, n1140, n1141_1, n1142, n1143, n1144, n1145, n1146_1, n1147, n1148, n1149, n1150, n1151_1, n1152, n1153, n1154, n1155, n1156_1, n1157, n1158, n1159, n1160, n1162, n1163, n1165, n1166_1, n1167, n1168, n1169, n1170, n1171_1, n1172, n1173, n1174, n1175, n1178, n1179, n1180, n1181_1, n1182, n1183, n1184, n1185, n1186_1, n1187, n1188, n1189, n1190, n1191_1, n1192, n1193, n1194, n1195, n1196_1, n1197, n1198, n1199, n1200, n1201_1, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1228, n1230, n1231, n1232, n1234, n1235, n1236, n1237, n1238, n1240, n1241, n1242, n1243, n1244, n1246, n1248, n1249, n1250, n1251, n1253, n1254, n1256, n1258, n1259, n1260, n1262, n1263, n1265, n1266, n1269, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1290, n1292, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1316, n1317, n1318, n1319, n1323, n1325, n1328, n1329, n1331, n1334, n1335, n1336, n1337, n1338, n1340, n1341, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1359, n1360, n1361, n1362, n1363, n1365, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1377, n1380, n1382, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1423, n1424, n1425, n1426, n1428, n1433, n1436, n1437, n1438, n1439, n1440, n1441, n1443, n1444, n1446, n1447, n1448, n1449, n1450, n1451, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1470, n1473, n1474, n1478, n1479, n1481, n1482, n1484, n1485, n1486, n1488, n1491, n1492, n1494, n1495, n1496, n1497, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1508, n1511, n1512, n1514, n1515, n1518, n1519, n1520, n1522, n1523, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1594, n1595, n1596, n1598, n1600, n1601, n1603, n1604, n1606, n1607, n1609, n1610, n1612, n1613, n1614, n1615, n1617, n1619, n1621, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1633, n1635, n1636, n1638, n1640, n1642, n1643, n1644, n1645, n1647, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1657, n1659, n1660, n1662, n1663, n1664, n1665, n1666, n1668, n1670, n1672, n1675, n1676, n1677, n1680, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1697, n1699, n1700, n1702, n1703, n1707, n1708, n1712, n1713, n1716, n1719, n1720, n1722, n1723, n1724, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1741, n1742, n1743, n1744, n1745, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1762, n1763, n1767, n1769, n1770, n1771, n1772, n1774, n1775, n1780, n1781, n1782, n1783, n1784, n1786, n1787, n1788, n1789, n1790, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1829, n1830, n1831, n1832, n1833, n1834, n1838, n1839, n1840, n1841, n1842, n1844, n1845, n1847, n1848, n1849, n1850, n1851;
INVX1    g0000(.A(g89), .Y(n708));
NOR2X1   g0001(.A(g102), .B(n708), .Y(g2584));
INVX1    g0002(.A(g486), .Y(n710));
INVX1    g0003(.A(g489), .Y(n711_1));
AOI22X1  g0004(.A0(g492), .A1(n711_1), .B0(n710), .B1(g496), .Y(g4809));
ZERO     g0005(.Y(g5692));
INVX1    g0006(.A(g675), .Y(n714));
OR2X1    g0007(.A(n714), .B(g22), .Y(n715));
INVX1    g0008(.A(g48), .Y(n716_1));
XOR2X1   g0009(.A(g1), .B(g2), .Y(n717));
XOR2X1   g0010(.A(g10), .B(g6), .Y(n718));
XOR2X1   g0011(.A(n718), .B(n717), .Y(n719));
XOR2X1   g0012(.A(g14), .B(g18), .Y(n720));
XOR2X1   g0013(.A(g28), .B(g24), .Y(n721_1));
XOR2X1   g0014(.A(n721_1), .B(n720), .Y(n722));
XOR2X1   g0015(.A(n722), .B(n719), .Y(n723));
AND2X1   g0016(.A(n723), .B(n716_1), .Y(n724));
INVX1    g0017(.A(g41), .Y(n725));
OAI21X1  g0018(.A0(n723), .A1(n716_1), .B0(n725), .Y(n726_1));
OAI21X1  g0019(.A0(n726_1), .A1(n724), .B0(g676), .Y(n727));
OR2X1    g0020(.A(n727), .B(n715), .Y(g6282));
NOR3X1   g0021(.A(n727), .B(n715), .C(n725), .Y(n729));
XOR2X1   g0022(.A(g29), .B(g33), .Y(n730));
XOR2X1   g0023(.A(g19), .B(g25), .Y(n731_1));
XOR2X1   g0024(.A(n731_1), .B(n730), .Y(n732));
XOR2X1   g0025(.A(g15), .B(g11), .Y(n733));
XOR2X1   g0026(.A(g7), .B(g3), .Y(n734));
XOR2X1   g0027(.A(n734), .B(n733), .Y(n735));
XOR2X1   g0028(.A(n735), .B(n732), .Y(n736_1));
NAND2X1  g0029(.A(n736_1), .B(n729), .Y(g6284));
OR4X1    g0030(.A(n715), .B(g25), .C(n725), .D(n727), .Y(g6360));
OR4X1    g0031(.A(n715), .B(g29), .C(n725), .D(n727), .Y(g6362));
OR4X1    g0032(.A(n715), .B(g3), .C(n725), .D(n727), .Y(g6364));
OR4X1    g0033(.A(n715), .B(g33), .C(n725), .D(n727), .Y(g6366));
OR4X1    g0034(.A(n715), .B(g7), .C(n725), .D(n727), .Y(g6368));
OR4X1    g0035(.A(n715), .B(g11), .C(n725), .D(n727), .Y(g6370));
OR4X1    g0036(.A(n715), .B(g15), .C(n725), .D(n727), .Y(g6372));
OR4X1    g0037(.A(n715), .B(g19), .C(n725), .D(n727), .Y(g6374));
ZERO     g0038(.Y(g6728));
NAND2X1  g0039(.A(g638), .B(g567), .Y(g4121));
INVX1    g0040(.A(g357), .Y(n748));
INVX1    g0041(.A(g353), .Y(n749));
NOR4X1   g0042(.A(g341), .B(g338), .C(g349), .D(g345), .Y(n750));
NAND4X1  g0043(.A(n749), .B(n748), .C(g323), .D(n750), .Y(n751_1));
NOR2X1   g0044(.A(g310), .B(g306), .Y(n752));
NOR2X1   g0045(.A(n752), .B(g332), .Y(n753));
MX2X1    g0046(.A(n753), .B(g332), .S0(n751_1), .Y(n754));
NOR4X1   g0047(.A(g310), .B(g306), .C(g301), .D(g314), .Y(n755));
INVX1    g0048(.A(g337), .Y(n756_1));
INVX1    g0049(.A(g687), .Y(n757));
INVX1    g0050(.A(g689), .Y(n758));
NOR2X1   g0051(.A(g698), .B(n758), .Y(n759));
INVX1    g0052(.A(g658), .Y(n760));
NAND2X1  g0053(.A(n760), .B(g662), .Y(n761_1));
NAND2X1  g0054(.A(g699), .B(g702), .Y(n762));
NOR4X1   g0055(.A(n761_1), .B(n727), .C(g41), .D(n762), .Y(n763));
NAND4X1  g0056(.A(n759), .B(g677), .C(n757), .D(n763), .Y(n764));
INVX1    g0057(.A(g677), .Y(n765));
NAND4X1  g0058(.A(n759), .B(n765), .C(n757), .D(n763), .Y(n766_1));
AND2X1   g0059(.A(g658), .B(g662), .Y(n767));
INVX1    g0060(.A(n767), .Y(n768));
OR4X1    g0061(.A(n761_1), .B(n727), .C(n725), .D(n762), .Y(n769));
NOR4X1   g0062(.A(g687), .B(g698), .C(n758), .D(n769), .Y(n770));
INVX1    g0063(.A(n770), .Y(n771_1));
NAND4X1  g0064(.A(n768), .B(n766_1), .C(n764), .D(n771_1), .Y(n772));
NAND4X1  g0065(.A(n759), .B(g677), .C(g687), .D(n763), .Y(n773));
NAND4X1  g0066(.A(n759), .B(n765), .C(g687), .D(n763), .Y(n774));
NOR4X1   g0067(.A(n757), .B(g698), .C(n758), .D(n769), .Y(n775));
INVX1    g0068(.A(n775), .Y(n776_1));
NAND4X1  g0069(.A(n774), .B(n773), .C(n768), .D(n776_1), .Y(n777));
NAND3X1  g0070(.A(n777), .B(n772), .C(n756_1), .Y(n778));
MX2X1    g0071(.A(n754), .B(n778), .S0(n755), .Y(n156));
INVX1    g0072(.A(g123), .Y(n780));
INVX1    g0073(.A(g139), .Y(n781_1));
NOR3X1   g0074(.A(g135), .B(g131), .C(g128), .Y(n782));
NAND3X1  g0075(.A(n782), .B(g114), .C(n781_1), .Y(n783));
INVX1    g0076(.A(n783), .Y(n784));
OR2X1    g0077(.A(g98), .B(g94), .Y(n785));
NAND3X1  g0078(.A(n784), .B(n785), .C(n780), .Y(n786_1));
OAI21X1  g0079(.A0(n784), .A1(n780), .B0(n786_1), .Y(n787));
NOR4X1   g0080(.A(g98), .B(g94), .C(g89), .D(g102), .Y(n788));
INVX1    g0081(.A(g685), .Y(n789));
INVX1    g0082(.A(g254), .Y(n790));
MX2X1    g0083(.A(n789), .B(n790), .S0(g658), .Y(n791_1));
INVX1    g0084(.A(g684), .Y(n792));
INVX1    g0085(.A(g248), .Y(n793));
MX2X1    g0086(.A(n792), .B(n793), .S0(g658), .Y(n794));
INVX1    g0087(.A(g683), .Y(n795));
INVX1    g0088(.A(g242), .Y(n796_1));
MX2X1    g0089(.A(n795), .B(n796_1), .S0(g658), .Y(n797));
INVX1    g0090(.A(g682), .Y(n798));
INVX1    g0091(.A(g236), .Y(n799));
MX2X1    g0092(.A(n798), .B(n799), .S0(g658), .Y(n800));
OAI22X1  g0093(.A0(n797), .A1(n800), .B0(n794), .B1(n791_1), .Y(n801_1));
INVX1    g0094(.A(g678), .Y(n802));
INVX1    g0095(.A(g212), .Y(n803));
MX2X1    g0096(.A(n802), .B(n803), .S0(g658), .Y(n804));
INVX1    g0097(.A(g679), .Y(n805));
INVX1    g0098(.A(g218), .Y(n806_1));
MX2X1    g0099(.A(n805), .B(n806_1), .S0(g658), .Y(n807));
INVX1    g0100(.A(g688), .Y(n808));
OR2X1    g0101(.A(g698), .B(g689), .Y(n809));
NOR3X1   g0102(.A(n809), .B(n808), .C(n757), .Y(n810));
AOI22X1  g0103(.A0(n767), .A1(g297), .B0(n763), .B1(n810), .Y(n811_1));
INVX1    g0104(.A(g224), .Y(n812));
INVX1    g0105(.A(g680), .Y(n813));
MX2X1    g0106(.A(n812), .B(n813), .S0(n760), .Y(n814));
NOR3X1   g0107(.A(n814), .B(n811_1), .C(n807), .Y(n815));
INVX1    g0108(.A(n807), .Y(n816_1));
INVX1    g0109(.A(n814), .Y(n817));
NOR3X1   g0110(.A(n817), .B(n811_1), .C(n816_1), .Y(n818));
OAI21X1  g0111(.A0(n818), .A1(n815), .B0(n804), .Y(n819));
INVX1    g0112(.A(n804), .Y(n820));
NOR3X1   g0113(.A(n814), .B(n811_1), .C(n816_1), .Y(n821_1));
OAI21X1  g0114(.A0(n821_1), .A1(n815), .B0(n820), .Y(n822));
NOR3X1   g0115(.A(n817), .B(n811_1), .C(n807), .Y(n823));
OAI21X1  g0116(.A0(n823), .A1(n821_1), .B0(n804), .Y(n824));
OAI21X1  g0117(.A0(n823), .A1(n818), .B0(n820), .Y(n825));
INVX1    g0118(.A(g681), .Y(n826_1));
INVX1    g0119(.A(g230), .Y(n827));
MX2X1    g0120(.A(n826_1), .B(n827), .S0(g658), .Y(n828));
NAND4X1  g0121(.A(n824), .B(n822), .C(n819), .D(n825), .Y(n829));
AND2X1   g0122(.A(n829), .B(n801_1), .Y(n830));
INVX1    g0123(.A(g567), .Y(n831_1));
INVX1    g0124(.A(g691), .Y(n916));
NOR4X1   g0125(.A(g634), .B(g598), .C(n831_1), .D(n916), .Y(n833));
INVX1    g0126(.A(g598), .Y(n834));
INVX1    g0127(.A(g697), .Y(n835));
INVX1    g0128(.A(g634), .Y(n836_1));
NOR4X1   g0129(.A(n835), .B(n834), .C(n831_1), .D(n836_1), .Y(n837));
INVX1    g0130(.A(g692), .Y(n838));
NOR4X1   g0131(.A(g634), .B(n834), .C(g567), .D(n838), .Y(n839));
INVX1    g0132(.A(g690), .Y(n496));
NOR4X1   g0133(.A(g634), .B(g598), .C(g567), .D(n496), .Y(n841_1));
NOR4X1   g0134(.A(n839), .B(n837), .C(n833), .D(n841_1), .Y(n842));
INVX1    g0135(.A(g693), .Y(n843));
NOR4X1   g0136(.A(g634), .B(n834), .C(n831_1), .D(n843), .Y(n844));
INVX1    g0137(.A(g695), .Y(n845));
NOR4X1   g0138(.A(g598), .B(n845), .C(n831_1), .D(n836_1), .Y(n846_1));
INVX1    g0139(.A(g696), .Y(n847));
NOR4X1   g0140(.A(n836_1), .B(n834), .C(g567), .D(n847), .Y(n848));
INVX1    g0141(.A(g694), .Y(n849));
NOR4X1   g0142(.A(n836_1), .B(g598), .C(g567), .D(n849), .Y(n850));
NOR4X1   g0143(.A(n848), .B(n846_1), .C(n844), .D(n850), .Y(n851_1));
XOR2X1   g0144(.A(g288), .B(g682), .Y(n852));
XOR2X1   g0145(.A(g683), .B(g289), .Y(n853));
XOR2X1   g0146(.A(g287), .B(g681), .Y(n854));
XOR2X1   g0147(.A(g286), .B(n813), .Y(n855));
XOR2X1   g0148(.A(g284), .B(n802), .Y(n856_1));
XOR2X1   g0149(.A(g290), .B(g684), .Y(n857));
XOR2X1   g0150(.A(g679), .B(g285), .Y(n858));
XOR2X1   g0151(.A(g685), .B(g291), .Y(n859));
XOR2X1   g0152(.A(g686), .B(g292), .Y(n860));
NOR4X1   g0153(.A(n859), .B(n858), .C(n857), .D(n860), .Y(n861_1));
NAND3X1  g0154(.A(n861_1), .B(n856_1), .C(n855), .Y(n862));
NOR4X1   g0155(.A(n854), .B(n853), .C(n852), .D(n862), .Y(n863));
AOI21X1  g0156(.A0(n851_1), .A1(n842), .B0(n863), .Y(n864));
INVX1    g0157(.A(n864), .Y(n865));
INVX1    g0158(.A(g281), .Y(n866_1));
INVX1    g0159(.A(g279), .Y(n867));
INVX1    g0160(.A(g280), .Y(n868));
NAND3X1  g0161(.A(g277), .B(g276), .C(g278), .Y(n869));
NOR4X1   g0162(.A(n868), .B(n867), .C(n866_1), .D(n869), .Y(n870));
INVX1    g0163(.A(n870), .Y(n871_1));
INVX1    g0164(.A(g478), .Y(n872));
AOI21X1  g0165(.A0(g696), .A1(g276), .B0(g277), .Y(n873));
OAI21X1  g0166(.A0(n835), .A1(g276), .B0(n873), .Y(n874));
INVX1    g0167(.A(g276), .Y(n875));
NAND2X1  g0168(.A(n875), .B(g695), .Y(n876_1));
INVX1    g0169(.A(g277), .Y(n877));
AOI21X1  g0170(.A0(g694), .A1(g276), .B0(n877), .Y(n878));
AOI21X1  g0171(.A0(n878), .A1(n876_1), .B0(g278), .Y(n879));
AOI21X1  g0172(.A0(g692), .A1(g276), .B0(g277), .Y(n880));
OAI21X1  g0173(.A0(n843), .A1(g276), .B0(n880), .Y(n881_1));
INVX1    g0174(.A(g278), .Y(n882));
NAND2X1  g0175(.A(g691), .B(n875), .Y(n883));
AOI21X1  g0176(.A0(g690), .A1(g276), .B0(n877), .Y(n884));
AOI21X1  g0177(.A0(n884), .A1(n883), .B0(n882), .Y(n885));
AOI22X1  g0178(.A0(n881_1), .A1(n885), .B0(n879), .B1(n874), .Y(n886_1));
NAND2X1  g0179(.A(n886_1), .B(n867), .Y(n887));
NAND2X1  g0180(.A(n886_1), .B(g279), .Y(n888));
AOI21X1  g0181(.A0(n888), .A1(n887), .B0(n872), .Y(n889));
NAND2X1  g0182(.A(g697), .B(n875), .Y(n890));
AND2X1   g0183(.A(n873), .B(n890), .Y(n891_1));
NOR2X1   g0184(.A(g276), .B(n845), .Y(n892));
OAI21X1  g0185(.A0(n849), .A1(n875), .B0(g277), .Y(n893));
OAI21X1  g0186(.A0(n893), .A1(n892), .B0(n882), .Y(n894));
NAND2X1  g0187(.A(g693), .B(n875), .Y(n895));
AND2X1   g0188(.A(n880), .B(n895), .Y(n896_1));
NOR2X1   g0189(.A(n916), .B(g276), .Y(n897));
OAI21X1  g0190(.A0(n496), .A1(n875), .B0(g277), .Y(n898));
OAI21X1  g0191(.A0(n898), .A1(n897), .B0(g278), .Y(n899));
OAI22X1  g0192(.A0(n896_1), .A1(n899), .B0(n894), .B1(n891_1), .Y(n900));
NOR2X1   g0193(.A(n900), .B(g279), .Y(n901_1));
NOR2X1   g0194(.A(n900), .B(n867), .Y(n902));
NOR3X1   g0195(.A(n902), .B(n901_1), .C(g478), .Y(n903));
INVX1    g0196(.A(g282), .Y(n904));
INVX1    g0197(.A(g283), .Y(n905));
XOR2X1   g0198(.A(g280), .B(n866_1), .Y(n906_1));
INVX1    g0199(.A(n906_1), .Y(n907));
NOR3X1   g0200(.A(n907), .B(n905), .C(n904), .Y(n908));
OAI21X1  g0201(.A0(n903), .A1(n889), .B0(n908), .Y(n909));
NOR4X1   g0202(.A(g280), .B(n867), .C(n866_1), .D(n869), .Y(n910));
NOR2X1   g0203(.A(n910), .B(n906_1), .Y(n911_1));
XOR2X1   g0204(.A(n911_1), .B(n872), .Y(n912));
NOR4X1   g0205(.A(n906_1), .B(n905), .C(n904), .D(n912), .Y(n913));
INVX1    g0206(.A(n913), .Y(n914));
AOI21X1  g0207(.A0(n914), .A1(n909), .B0(n871_1), .Y(n915));
NOR3X1   g0208(.A(n907), .B(g283), .C(n904), .Y(n916_1));
OAI21X1  g0209(.A0(n903), .A1(n889), .B0(n916_1), .Y(n917));
NOR2X1   g0210(.A(n917), .B(n871_1), .Y(n918));
NAND3X1  g0211(.A(n870), .B(g283), .C(n904), .Y(n919));
OR4X1    g0212(.A(g478), .B(g283), .C(g282), .D(n911_1), .Y(n920));
NAND2X1  g0213(.A(n920), .B(n919), .Y(n921_1));
NAND4X1  g0214(.A(n872), .B(n905), .C(n904), .D(n911_1), .Y(n922));
NAND3X1  g0215(.A(n907), .B(n905), .C(g282), .Y(n923));
OAI21X1  g0216(.A0(n923), .A1(n912), .B0(n922), .Y(n924));
OR4X1    g0217(.A(n921_1), .B(n918), .C(n915), .D(n905), .Y(n926_1));
AOI21X1  g0218(.A0(n914), .A1(n909), .B0(n870), .Y(n927));
NOR2X1   g0219(.A(n917), .B(n870), .Y(n928));
NOR3X1   g0220(.A(n871_1), .B(g283), .C(n904), .Y(n929));
AND2X1   g0221(.A(n929), .B(n917), .Y(n930));
NOR3X1   g0222(.A(n930), .B(n928), .C(n927), .Y(n931_1));
NAND2X1  g0223(.A(n931_1), .B(n926_1), .Y(n932));
OR4X1    g0224(.A(n927), .B(n924), .C(n904), .D(n928), .Y(n933));
NOR4X1   g0225(.A(n921_1), .B(n918), .C(n915), .D(n930), .Y(n934));
NAND2X1  g0226(.A(n934), .B(n933), .Y(n935));
NAND3X1  g0227(.A(n935), .B(n932), .C(n865), .Y(n936_1));
MX2X1    g0228(.A(g690), .B(n936_1), .S0(g658), .Y(n937));
OR4X1    g0229(.A(n761_1), .B(n727), .C(g41), .D(n762), .Y(n938));
INVX1    g0230(.A(g698), .Y(n939));
NOR3X1   g0231(.A(g688), .B(n939), .C(n758), .Y(n940));
INVX1    g0232(.A(n940), .Y(n941_1));
NOR4X1   g0233(.A(n938), .B(g685), .C(n792), .D(n941_1), .Y(n942));
NOR4X1   g0234(.A(n769), .B(g685), .C(n792), .D(n941_1), .Y(n943));
NOR3X1   g0235(.A(n943), .B(n942), .C(n767), .Y(n944));
MX2X1    g0236(.A(g683), .B(g571), .S0(g658), .Y(n945));
MX2X1    g0237(.A(g682), .B(g654), .S0(g658), .Y(n946_1));
AND2X1   g0238(.A(n946_1), .B(n945), .Y(n947));
NOR4X1   g0239(.A(n943), .B(n942), .C(n767), .D(n947), .Y(n948));
MX2X1    g0240(.A(g681), .B(g650), .S0(g658), .Y(n949));
MX2X1    g0241(.A(g680), .B(g646), .S0(g658), .Y(n950));
MX2X1    g0242(.A(g679), .B(g606), .S0(g658), .Y(n951_1));
MX2X1    g0243(.A(g678), .B(g642), .S0(g658), .Y(n952));
AOI22X1  g0244(.A0(n951_1), .A1(n952), .B0(n950), .B1(n949), .Y(n953));
INVX1    g0245(.A(g686), .Y(n954));
INVX1    g0246(.A(g260), .Y(n955));
MX2X1    g0247(.A(n954), .B(n955), .S0(g658), .Y(n956_1));
NOR4X1   g0248(.A(n953), .B(n948), .C(n944), .D(n956_1), .Y(n957));
OAI21X1  g0249(.A0(n937), .A1(n830), .B0(n957), .Y(n958));
MX2X1    g0250(.A(n787), .B(n958), .S0(n788), .Y(n161));
INVX1    g0251(.A(g207), .Y(n960));
INVX1    g0252(.A(g208), .Y(n961_1));
INVX1    g0253(.A(g209), .Y(n962));
NAND3X1  g0254(.A(g205), .B(g204), .C(g206), .Y(n963));
OR4X1    g0255(.A(n962), .B(n961_1), .C(n960), .D(n963), .Y(n964));
INVX1    g0256(.A(g471), .Y(n965));
INVX1    g0257(.A(g211), .Y(n966_1));
INVX1    g0258(.A(g210), .Y(n967));
NOR4X1   g0259(.A(n962), .B(g208), .C(n960), .D(n963), .Y(n968));
XOR2X1   g0260(.A(g209), .B(n961_1), .Y(n969));
NOR2X1   g0261(.A(n969), .B(n968), .Y(n970));
NAND4X1  g0262(.A(n967), .B(n966_1), .C(n965), .D(n970), .Y(n971_1));
AND2X1   g0263(.A(n971_1), .B(n964), .Y(n972));
XOR2X1   g0264(.A(n963), .B(g207), .Y(n973));
AND2X1   g0265(.A(n973), .B(n972), .Y(n974));
OR4X1    g0266(.A(g210), .B(g211), .C(g471), .D(n970), .Y(n975));
NAND2X1  g0267(.A(n975), .B(g197), .Y(n976_1));
OAI22X1  g0268(.A0(n974), .A1(n976_1), .B0(g197), .B1(n843), .Y(n166));
XOR2X1   g0269(.A(g236), .B(g516), .Y(n978));
XOR2X1   g0270(.A(g512), .B(g230), .Y(n979));
XOR2X1   g0271(.A(g242), .B(g520), .Y(n980));
OR2X1    g0272(.A(n980), .B(n979), .Y(n981_1));
XOR2X1   g0273(.A(g524), .B(n793), .Y(n982));
XOR2X1   g0274(.A(g532), .B(n955), .Y(n983));
NAND2X1  g0275(.A(n983), .B(n982), .Y(n984));
XOR2X1   g0276(.A(g508), .B(g224), .Y(n985));
XOR2X1   g0277(.A(g254), .B(g528), .Y(n986_1));
XOR2X1   g0278(.A(g218), .B(g504), .Y(n987));
XOR2X1   g0279(.A(g500), .B(g212), .Y(n988));
NOR4X1   g0280(.A(n987), .B(n986_1), .C(n985), .D(n988), .Y(n989));
INVX1    g0281(.A(n989), .Y(n990));
NOR4X1   g0282(.A(n984), .B(n981_1), .C(n978), .D(n990), .Y(n991_1));
INVX1    g0283(.A(n991_1), .Y(n992));
NOR3X1   g0284(.A(n992), .B(g536), .C(g541), .Y(n993));
MX2X1    g0285(.A(g461), .B(g430), .S0(n993), .Y(n176));
INVX1    g0286(.A(n729), .Y(n995));
NAND2X1  g0287(.A(n995), .B(g25), .Y(n996_1));
NAND2X1  g0288(.A(n729), .B(g25), .Y(n997));
NAND2X1  g0289(.A(n997), .B(n996_1), .Y(n181));
INVX1    g0290(.A(g328), .Y(n999));
NOR3X1   g0291(.A(g314), .B(g310), .C(g306), .Y(n1000));
NOR2X1   g0292(.A(n1000), .B(n999), .Y(n191));
NAND2X1  g0293(.A(n995), .B(g29), .Y(n1002));
NAND2X1  g0294(.A(n729), .B(g29), .Y(n1003));
NAND2X1  g0295(.A(n1003), .B(n1002), .Y(n201));
INVX1    g0296(.A(g702), .Y(n1005));
INVX1    g0297(.A(g699), .Y(n1006_1));
OR4X1    g0298(.A(n1006_1), .B(g41), .C(n1005), .D(n727), .Y(n1007));
NOR4X1   g0299(.A(n939), .B(n789), .C(n758), .D(g688), .Y(n1008));
INVX1    g0300(.A(n1008), .Y(n1009));
NAND4X1  g0301(.A(n826_1), .B(g684), .C(n798), .D(g683), .Y(n1010));
NOR4X1   g0302(.A(n1009), .B(n1007), .C(g677), .D(n1010), .Y(n1011_1));
MX2X1    g0303(.A(g465), .B(g691), .S0(n1011_1), .Y(n206));
INVX1    g0304(.A(g84), .Y(n1013));
INVX1    g0305(.A(n751_1), .Y(n1014));
INVX1    g0306(.A(g306), .Y(n1015));
INVX1    g0307(.A(g310), .Y(n1016_1));
INVX1    g0308(.A(g332), .Y(n1017));
AOI21X1  g0309(.A0(n1016_1), .A1(n1015), .B0(n1017), .Y(n1018));
INVX1    g0310(.A(g301), .Y(n1019));
INVX1    g0311(.A(g314), .Y(n1020));
NOR3X1   g0312(.A(g319), .B(n1020), .C(n1019), .Y(n1021_1));
OAI21X1  g0313(.A0(n1021_1), .A1(n1018), .B0(n1014), .Y(n1022));
OR2X1    g0314(.A(g310), .B(g301), .Y(n1023));
NOR4X1   g0315(.A(g319), .B(n1020), .C(g306), .D(n1023), .Y(n1024));
OAI21X1  g0316(.A0(n1024), .A1(g319), .B0(n1014), .Y(n1025));
NAND2X1  g0317(.A(n1025), .B(n1022), .Y(n1026_1));
INVX1    g0318(.A(g398), .Y(n1027));
INVX1    g0319(.A(g69), .Y(n1028));
INVX1    g0320(.A(g74), .Y(n1029));
INVX1    g0321(.A(g64), .Y(n1030));
NOR4X1   g0322(.A(g49), .B(g54), .C(g361), .D(g59), .Y(n1031_1));
NAND4X1  g0323(.A(n1030), .B(n1029), .C(n1028), .D(n1031_1), .Y(n1032));
OR2X1    g0324(.A(n1032), .B(g79), .Y(n1033));
NOR3X1   g0325(.A(g314), .B(n1016_1), .C(g306), .Y(n1034));
NOR2X1   g0326(.A(n1020), .B(g306), .Y(n1035));
NOR3X1   g0327(.A(g314), .B(g310), .C(n1015), .Y(n1036_1));
NOR3X1   g0328(.A(n1036_1), .B(n1035), .C(n1034), .Y(n1037));
NAND4X1  g0329(.A(g49), .B(g54), .C(g361), .D(g59), .Y(n1038));
NOR4X1   g0330(.A(n1030), .B(n1029), .C(n1028), .D(n1038), .Y(n1039));
NAND2X1  g0331(.A(n1039), .B(g79), .Y(n1040));
MX2X1    g0332(.A(n1040), .B(n1033), .S0(n1037), .Y(n1041_1));
MX2X1    g0333(.A(n1027), .B(n1041_1), .S0(n1025), .Y(n1042));
XOR2X1   g0334(.A(n1042), .B(g84), .Y(n1043));
MX2X1    g0335(.A(n1013), .B(n1043), .S0(n1026_1), .Y(n1044));
OR4X1    g0336(.A(n1035), .B(n1034), .C(g84), .D(n1036_1), .Y(n1045));
OR2X1    g0337(.A(n1045), .B(n1033), .Y(n1046_1));
INVX1    g0338(.A(g79), .Y(n1047));
INVX1    g0339(.A(n1039), .Y(n1048));
OR4X1    g0340(.A(n1037), .B(n1047), .C(n1013), .D(n1048), .Y(n1049));
AOI21X1  g0341(.A0(n1049), .A1(n1046_1), .B0(n1022), .Y(n1050));
OR2X1    g0342(.A(n1050), .B(n755), .Y(n1051_1));
AOI21X1  g0343(.A0(n1016_1), .A1(g306), .B0(n1021_1), .Y(n1052));
INVX1    g0344(.A(n1052), .Y(n1053));
NOR3X1   g0345(.A(n1053), .B(n755), .C(n1034), .Y(n1054));
OAI21X1  g0346(.A0(n1050), .A1(n755), .B0(n1054), .Y(n1055));
OAI21X1  g0347(.A0(n1051_1), .A1(n1044), .B0(n1055), .Y(n211));
XOR2X1   g0348(.A(g36), .B(g32), .Y(n1057));
XOR2X1   g0349(.A(g37), .B(g38), .Y(n1058));
XOR2X1   g0350(.A(n1058), .B(n1057), .Y(n1059));
XOR2X1   g0351(.A(g40), .B(g39), .Y(n1060));
XOR2X1   g0352(.A(n1060), .B(n1059), .Y(n1061_1));
XOR2X1   g0353(.A(n1061_1), .B(n723), .Y(n1062));
XOR2X1   g0354(.A(n1062), .B(g48), .Y(n221));
INVX1    g0355(.A(g639), .Y(n1064));
INVX1    g0356(.A(g622), .Y(n1065));
INVX1    g0357(.A(g619), .Y(n1066_1));
NAND4X1  g0358(.A(g610), .B(g602), .C(g613), .D(g616), .Y(n1067));
NOR2X1   g0359(.A(n1067), .B(n1066_1), .Y(n1068));
XOR2X1   g0360(.A(n1068), .B(n1065), .Y(n1069));
NOR2X1   g0361(.A(n1069), .B(n1064), .Y(n226));
NOR3X1   g0362(.A(g102), .B(g98), .C(g94), .Y(n1071_1));
OR2X1    g0363(.A(n1071_1), .B(g114), .Y(n231));
AND2X1   g0364(.A(n922), .B(n871_1), .Y(n1073));
AND2X1   g0365(.A(g277), .B(g276), .Y(n1074));
XOR2X1   g0366(.A(n1074), .B(g278), .Y(n1075));
NAND4X1  g0367(.A(n1073), .B(n920), .C(g269), .D(n1075), .Y(n1076_1));
OAI21X1  g0368(.A0(n838), .A1(g269), .B0(n1076_1), .Y(n236));
INVX1    g0369(.A(n788), .Y(n1078));
INVX1    g0370(.A(g128), .Y(n1079));
XOR2X1   g0371(.A(g114), .B(n1079), .Y(n1080));
NAND3X1  g0372(.A(n1080), .B(n1078), .C(n783), .Y(n241));
XOR2X1   g0373(.A(g598), .B(g567), .Y(n1082));
AND2X1   g0374(.A(n1082), .B(g638), .Y(n246));
MX2X1    g0375(.A(n932), .B(g554), .S0(n992), .Y(n251));
AOI21X1  g0376(.A0(g204), .A1(g696), .B0(g205), .Y(n1085));
OAI21X1  g0377(.A0(g204), .A1(n835), .B0(n1085), .Y(n1086_1));
INVX1    g0378(.A(g204), .Y(n1087));
NAND2X1  g0379(.A(n1087), .B(g695), .Y(n1088));
INVX1    g0380(.A(g205), .Y(n1089));
AOI21X1  g0381(.A0(g694), .A1(g204), .B0(n1089), .Y(n1090));
AOI21X1  g0382(.A0(n1090), .A1(n1088), .B0(g206), .Y(n1091_1));
AOI21X1  g0383(.A0(g692), .A1(g204), .B0(g205), .Y(n1092));
OAI21X1  g0384(.A0(g204), .A1(n843), .B0(n1092), .Y(n1093));
INVX1    g0385(.A(g206), .Y(n1094));
NAND2X1  g0386(.A(g691), .B(n1087), .Y(n1095));
AOI21X1  g0387(.A0(g204), .A1(g690), .B0(n1089), .Y(n1096_1));
AOI21X1  g0388(.A0(n1096_1), .A1(n1095), .B0(n1094), .Y(n1097));
AOI22X1  g0389(.A0(n1093), .A1(n1097), .B0(n1091_1), .B1(n1086_1), .Y(n1098));
NAND2X1  g0390(.A(n1098), .B(n960), .Y(n1099));
NAND2X1  g0391(.A(n1098), .B(g207), .Y(n1100));
AOI21X1  g0392(.A0(n1100), .A1(n1099), .B0(n965), .Y(n1101_1));
NAND2X1  g0393(.A(n1087), .B(g697), .Y(n1102));
AND2X1   g0394(.A(n1085), .B(n1102), .Y(n1103));
NOR2X1   g0395(.A(g204), .B(n845), .Y(n1104));
OAI21X1  g0396(.A0(n849), .A1(n1087), .B0(g205), .Y(n1105));
OAI21X1  g0397(.A0(n1105), .A1(n1104), .B0(n1094), .Y(n1106_1));
NAND2X1  g0398(.A(n1087), .B(g693), .Y(n1107));
AND2X1   g0399(.A(n1092), .B(n1107), .Y(n1108));
NOR2X1   g0400(.A(n916), .B(g204), .Y(n1109));
OAI21X1  g0401(.A0(n1087), .A1(n496), .B0(g205), .Y(n1110));
OAI21X1  g0402(.A0(n1110), .A1(n1109), .B0(g206), .Y(n1111_1));
OAI22X1  g0403(.A0(n1108), .A1(n1111_1), .B0(n1106_1), .B1(n1103), .Y(n1112));
NOR2X1   g0404(.A(n1112), .B(g207), .Y(n1113));
NOR2X1   g0405(.A(n1112), .B(n960), .Y(n1114));
NOR3X1   g0406(.A(n1114), .B(n1113), .C(g471), .Y(n1115));
INVX1    g0407(.A(n969), .Y(n1116_1));
NOR3X1   g0408(.A(n1116_1), .B(n967), .C(n966_1), .Y(n1117));
OAI21X1  g0409(.A0(n1115), .A1(n1101_1), .B0(n1117), .Y(n1118));
XOR2X1   g0410(.A(n970), .B(n965), .Y(n1119));
OR4X1    g0411(.A(n969), .B(n967), .C(n966_1), .D(n1119), .Y(n1120));
AOI21X1  g0412(.A0(n1120), .A1(n1118), .B0(n964), .Y(n1121_1));
INVX1    g0413(.A(n964), .Y(n1122));
AOI21X1  g0414(.A0(n1120), .A1(n1118), .B0(n1122), .Y(n1123));
OR2X1    g0415(.A(n1123), .B(g496), .Y(n1124));
OR2X1    g0416(.A(n1124), .B(n1121_1), .Y(n256));
INVX1    g0417(.A(g179), .Y(n1126_1));
INVX1    g0418(.A(g94), .Y(n1127));
INVX1    g0419(.A(g98), .Y(n1128));
AOI21X1  g0420(.A0(n1128), .A1(n1127), .B0(n780), .Y(n1129));
INVX1    g0421(.A(g102), .Y(n1130));
NOR3X1   g0422(.A(g107), .B(n1130), .C(n708), .Y(n1131_1));
OAI21X1  g0423(.A0(n1131_1), .A1(n1129), .B0(n784), .Y(n1132));
OR2X1    g0424(.A(g98), .B(g89), .Y(n1133));
NOR4X1   g0425(.A(g107), .B(n1130), .C(g94), .D(n1133), .Y(n1134));
OAI21X1  g0426(.A0(n1134), .A1(g107), .B0(n784), .Y(n1135));
NAND2X1  g0427(.A(n1135), .B(n1132), .Y(n1136_1));
INVX1    g0428(.A(g184), .Y(n1137));
NOR4X1   g0429(.A(g152), .B(g170), .C(g143), .D(g161), .Y(n1138));
INVX1    g0430(.A(n1138), .Y(n1139));
NOR3X1   g0431(.A(g102), .B(n1128), .C(g94), .Y(n1140));
NOR2X1   g0432(.A(n1130), .B(g94), .Y(n1141_1));
NOR3X1   g0433(.A(g102), .B(g98), .C(n1127), .Y(n1142));
NOR3X1   g0434(.A(n1142), .B(n1141_1), .C(n1140), .Y(n1143));
NAND4X1  g0435(.A(g152), .B(g170), .C(g143), .D(g161), .Y(n1144));
MX2X1    g0436(.A(n1144), .B(n1139), .S0(n1143), .Y(n1145));
MX2X1    g0437(.A(n1137), .B(n1145), .S0(n1135), .Y(n1146_1));
XOR2X1   g0438(.A(n1146_1), .B(g179), .Y(n1147));
MX2X1    g0439(.A(n1126_1), .B(n1147), .S0(n1136_1), .Y(n1148));
NAND2X1  g0440(.A(n1138), .B(n1126_1), .Y(n1149));
OR4X1    g0441(.A(n1141_1), .B(n1140), .C(g188), .D(n1142), .Y(n1150));
NOR2X1   g0442(.A(n1150), .B(n1149), .Y(n1151_1));
INVX1    g0443(.A(g188), .Y(n1152));
OR2X1    g0444(.A(n1144), .B(n1126_1), .Y(n1153));
NOR3X1   g0445(.A(n1153), .B(n1143), .C(n1152), .Y(n1154));
NOR2X1   g0446(.A(n1154), .B(n1151_1), .Y(n1155));
OAI21X1  g0447(.A0(n1155), .A1(n1132), .B0(n1078), .Y(n1156_1));
OR2X1    g0448(.A(n1155), .B(n1132), .Y(n1157));
AOI21X1  g0449(.A0(n1128), .A1(g94), .B0(n1131_1), .Y(n1158));
INVX1    g0450(.A(n1158), .Y(n1159));
OR4X1    g0451(.A(n1157), .B(n788), .C(n1140), .D(n1159), .Y(n1160));
OAI21X1  g0452(.A0(n1156_1), .A1(n1148), .B0(n1160), .Y(n261));
OR2X1    g0453(.A(n736_1), .B(n729), .Y(n1162));
OR4X1    g0454(.A(n727), .B(n715), .C(n725), .D(n736_1), .Y(n1163));
NAND2X1  g0455(.A(n1163), .B(n1162), .Y(n266));
INVX1    g0456(.A(g590), .Y(n1165));
INVX1    g0457(.A(g574), .Y(n1166_1));
INVX1    g0458(.A(g625), .Y(n1167));
NOR4X1   g0459(.A(n1167), .B(n1066_1), .C(n1065), .D(n1067), .Y(n1168));
AND2X1   g0460(.A(n1168), .B(g628), .Y(n1169));
AND2X1   g0461(.A(n1169), .B(g631), .Y(n1170));
NAND4X1  g0462(.A(g582), .B(g578), .C(g586), .D(n1170), .Y(n1171_1));
NOR3X1   g0463(.A(n1171_1), .B(n1166_1), .C(n1165), .Y(n1172));
AOI21X1  g0464(.A0(n1172), .A1(g594), .B0(n1064), .Y(n1173));
OR2X1    g0465(.A(n1171_1), .B(n1166_1), .Y(n1174));
XOR2X1   g0466(.A(n1174), .B(g590), .Y(n1175));
NAND2X1  g0467(.A(n1175), .B(n1173), .Y(n271));
MX2X1    g0468(.A(n935), .B(g551), .S0(n992), .Y(n276));
NOR4X1   g0469(.A(n769), .B(g685), .C(g684), .D(n941_1), .Y(n1178));
OAI21X1  g0470(.A0(g266), .A1(g662), .B0(n760), .Y(n1179));
OR4X1    g0471(.A(n1006_1), .B(n725), .C(n1005), .D(n1179), .Y(n1180));
NOR3X1   g0472(.A(n1180), .B(n795), .C(n792), .Y(n1181_1));
NAND4X1  g0473(.A(n1008), .B(n765), .C(g682), .D(n1181_1), .Y(n1182));
NAND4X1  g0474(.A(n1008), .B(g677), .C(g682), .D(n1181_1), .Y(n1183));
NAND2X1  g0475(.A(n1183), .B(n1182), .Y(n1184));
NOR3X1   g0476(.A(n1184), .B(n1178), .C(n943), .Y(n1185));
NOR4X1   g0477(.A(n769), .B(g688), .C(g687), .D(n809), .Y(n1186_1));
NOR4X1   g0478(.A(n769), .B(g688), .C(n757), .D(n809), .Y(n1187));
NOR4X1   g0479(.A(n1186_1), .B(n775), .C(n770), .D(n1187), .Y(n1188));
NAND3X1  g0480(.A(g688), .B(g698), .C(g689), .Y(n1189));
OR4X1    g0481(.A(g680), .B(n805), .C(n802), .D(n1189), .Y(n1190));
NOR4X1   g0482(.A(n1179), .B(n762), .C(n725), .D(n1190), .Y(n1191_1));
OR2X1    g0483(.A(g680), .B(g679), .Y(n1192));
NOR4X1   g0484(.A(n1189), .B(n1180), .C(n802), .D(n1192), .Y(n1193));
NOR4X1   g0485(.A(n1189), .B(n1180), .C(g678), .D(n1192), .Y(n1194));
OR4X1    g0486(.A(n813), .B(g679), .C(g678), .D(n1189), .Y(n1195));
NOR4X1   g0487(.A(n1179), .B(n762), .C(n725), .D(n1195), .Y(n1196_1));
OR4X1    g0488(.A(n1194), .B(n1193), .C(n1191_1), .D(n1196_1), .Y(n1197));
NOR4X1   g0489(.A(n1009), .B(g683), .C(n792), .D(n1180), .Y(n1198));
NOR4X1   g0490(.A(n826_1), .B(n792), .C(g682), .D(n795), .Y(n1199));
INVX1    g0491(.A(n1199), .Y(n1200));
NOR3X1   g0492(.A(n1200), .B(n1180), .C(n1009), .Y(n1201_1));
NAND4X1  g0493(.A(n1008), .B(n826_1), .C(n798), .D(n1181_1), .Y(n1202));
OR2X1    g0494(.A(n1202), .B(g677), .Y(n1203));
OR2X1    g0495(.A(n1202), .B(n765), .Y(n1204));
NAND2X1  g0496(.A(n1204), .B(n1203), .Y(n1205));
NOR4X1   g0497(.A(n1201_1), .B(n1198), .C(n1197), .D(n1205), .Y(n1206));
NAND3X1  g0498(.A(n1206), .B(n1188), .C(n1185), .Y(n1207));
INVX1    g0499(.A(n943), .Y(n1208));
NAND2X1  g0500(.A(n1198), .B(g293), .Y(n1209));
AOI22X1  g0501(.A0(n1191_1), .A1(g562), .B0(g551), .B1(n1201_1), .Y(n1210));
NAND2X1  g0502(.A(n1210), .B(n1209), .Y(n1211));
INVX1    g0503(.A(g453), .Y(n1212));
INVX1    g0504(.A(g536), .Y(n1213));
OAI22X1  g0505(.A0(n1182), .A1(n1212), .B0(n1213), .B1(n1203), .Y(n1214));
INVX1    g0506(.A(g410), .Y(n1215));
INVX1    g0507(.A(g508), .Y(n1216));
OAI22X1  g0508(.A0(n1183), .A1(n1215), .B0(n1216), .B1(n1204), .Y(n1217));
NOR3X1   g0509(.A(n1217), .B(n1214), .C(n1211), .Y(n1218));
OAI21X1  g0510(.A0(n1208), .A1(n838), .B0(n1218), .Y(n1219));
AOI21X1  g0511(.A0(n1178), .A1(g692), .B0(n1219), .Y(n1220));
NOR2X1   g0512(.A(n838), .B(g677), .Y(n1221));
AND2X1   g0513(.A(g692), .B(g677), .Y(n1222));
OAI22X1  g0514(.A0(n1221), .A1(n1222), .B0(n775), .B1(n770), .Y(n1223));
AND2X1   g0515(.A(g205), .B(g204), .Y(n1224));
XOR2X1   g0516(.A(n1224), .B(g206), .Y(n1225));
NAND4X1  g0517(.A(n975), .B(n972), .C(g197), .D(n1225), .Y(n1226));
OAI21X1  g0518(.A0(n838), .A1(g197), .B0(n1226), .Y(n411));
AOI22X1  g0519(.A0(n1187), .A1(n236), .B0(n1186_1), .B1(n411), .Y(n1228));
NAND4X1  g0520(.A(n1223), .B(n1220), .C(n1207), .D(n1228), .Y(n286));
INVX1    g0521(.A(g638), .Y(n1230));
NAND4X1  g0522(.A(g634), .B(g598), .C(g567), .D(g642), .Y(n1231));
XOR2X1   g0523(.A(n1231), .B(g606), .Y(n1232));
NOR2X1   g0524(.A(n1232), .B(n1230), .Y(n291));
INVX1    g0525(.A(g193), .Y(n1234));
MX2X1    g0526(.A(n1153), .B(n1149), .S0(n1143), .Y(n1235));
MX2X1    g0527(.A(n1234), .B(n1235), .S0(n1135), .Y(n1236));
XOR2X1   g0528(.A(n1236), .B(g188), .Y(n1237));
MX2X1    g0529(.A(n1152), .B(n1237), .S0(n1136_1), .Y(n1238));
OAI21X1  g0530(.A0(n1238), .A1(n1156_1), .B0(n1160), .Y(n296));
INVX1    g0531(.A(g606), .Y(n1240));
INVX1    g0532(.A(g642), .Y(n1241));
NAND3X1  g0533(.A(g634), .B(g598), .C(g567), .Y(n1242));
OR4X1    g0534(.A(n1241), .B(g646), .C(n1240), .D(n1242), .Y(n1243));
OAI21X1  g0535(.A0(n1231), .A1(n1240), .B0(g646), .Y(n1244));
AOI21X1  g0536(.A0(n1244), .A1(n1243), .B0(n1230), .Y(n301));
INVX1    g0537(.A(g326), .Y(n1246));
NOR2X1   g0538(.A(n1000), .B(n1246), .Y(n306));
INVX1    g0539(.A(g361), .Y(n1248));
NOR2X1   g0540(.A(n1025), .B(g366), .Y(n1249));
XOR2X1   g0541(.A(n1249), .B(g361), .Y(n1250));
MX2X1    g0542(.A(n1248), .B(n1250), .S0(n1026_1), .Y(n1251));
OAI21X1  g0543(.A0(n1251), .A1(n1051_1), .B0(n1055), .Y(n311));
NAND3X1  g0544(.A(n1014), .B(g319), .C(n1019), .Y(n1253));
NOR2X1   g0545(.A(n755), .B(n1027), .Y(n1254));
MX2X1    g0546(.A(g394), .B(n1254), .S0(n1253), .Y(n321));
XOR2X1   g0547(.A(n1067), .B(g619), .Y(n1256));
NOR2X1   g0548(.A(n1256), .B(n1064), .Y(n331));
NAND4X1  g0549(.A(g204), .B(g206), .C(g207), .D(g205), .Y(n1258));
XOR2X1   g0550(.A(n1258), .B(g208), .Y(n1259));
NAND4X1  g0551(.A(n975), .B(n971_1), .C(n964), .D(n1259), .Y(n1260));
MX2X1    g0552(.A(g694), .B(n1260), .S0(g197), .Y(n336));
INVX1    g0553(.A(g390), .Y(n1262));
NOR2X1   g0554(.A(n755), .B(n1262), .Y(n1263));
MX2X1    g0555(.A(g386), .B(n1263), .S0(n1253), .Y(n346));
NOR3X1   g0556(.A(n1067), .B(n1066_1), .C(n1065), .Y(n1265));
XOR2X1   g0557(.A(n1265), .B(n1167), .Y(n1266));
NOR2X1   g0558(.A(n1266), .B(n1064), .Y(n351));
MX2X1    g0559(.A(g437), .B(g441), .S0(n993), .Y(n361));
NAND4X1  g0560(.A(n920), .B(g269), .C(n875), .D(n1073), .Y(n1269));
OAI21X1  g0561(.A0(n496), .A1(g269), .B0(n1269), .Y(n366));
INVX1    g0562(.A(n1178), .Y(n1271));
AOI22X1  g0563(.A0(n1191_1), .A1(g564), .B0(g669), .B1(n1196_1), .Y(n1272));
AOI22X1  g0564(.A0(n1193), .A1(n710), .B0(g496), .B1(n1194), .Y(n1273));
AOI22X1  g0565(.A0(n1198), .A1(g197), .B0(g545), .B1(n1201_1), .Y(n1274));
NAND3X1  g0566(.A(n1274), .B(n1273), .C(n1272), .Y(n1275));
INVX1    g0567(.A(g461), .Y(n1276));
INVX1    g0568(.A(g532), .Y(n1277));
OAI22X1  g0569(.A0(n1182), .A1(n1276), .B0(n1277), .B1(n1203), .Y(n1278));
INVX1    g0570(.A(g402), .Y(n1279));
INVX1    g0571(.A(g500), .Y(n1280));
OAI22X1  g0572(.A0(n1183), .A1(n1279), .B0(n1280), .B1(n1204), .Y(n1281));
NOR3X1   g0573(.A(n1281), .B(n1278), .C(n1275), .Y(n1282));
OAI21X1  g0574(.A0(n1271), .A1(n496), .B0(n1282), .Y(n1283));
AOI21X1  g0575(.A0(n943), .A1(g690), .B0(n1283), .Y(n1284));
NOR2X1   g0576(.A(g677), .B(n496), .Y(n1285));
AND2X1   g0577(.A(g677), .B(g690), .Y(n1286));
OAI22X1  g0578(.A0(n1285), .A1(n1286), .B0(n775), .B1(n770), .Y(n1287));
NAND4X1  g0579(.A(n972), .B(g197), .C(n1087), .D(n975), .Y(n1288));
OAI21X1  g0580(.A0(g197), .A1(n496), .B0(n1288), .Y(n991));
AOI22X1  g0581(.A0(n366), .A1(n1187), .B0(n1186_1), .B1(n991), .Y(n1290));
NAND4X1  g0582(.A(n1287), .B(n1284), .C(n1207), .D(n1290), .Y(n371));
INVX1    g0583(.A(g331), .Y(n1292));
NOR2X1   g0584(.A(n1000), .B(n1292), .Y(n376));
INVX1    g0585(.A(g578), .Y(n1294));
INVX1    g0586(.A(g582), .Y(n1295));
OAI21X1  g0587(.A0(n1294), .A1(n847), .B0(n1295), .Y(n1296));
AOI21X1  g0588(.A0(n1294), .A1(g697), .B0(n1296), .Y(n1297));
INVX1    g0589(.A(g586), .Y(n1298));
NOR2X1   g0590(.A(g578), .B(n845), .Y(n1299));
OAI21X1  g0591(.A0(n849), .A1(n1294), .B0(g582), .Y(n1300));
OAI21X1  g0592(.A0(n1300), .A1(n1299), .B0(n1298), .Y(n1301));
OAI21X1  g0593(.A0(n838), .A1(n1294), .B0(n1295), .Y(n1302));
AOI21X1  g0594(.A0(n1294), .A1(g693), .B0(n1302), .Y(n1303));
NOR2X1   g0595(.A(n916), .B(g578), .Y(n1304));
OAI21X1  g0596(.A0(n1294), .A1(n496), .B0(g582), .Y(n1305));
OAI21X1  g0597(.A0(n1305), .A1(n1304), .B0(g586), .Y(n1306));
OAI22X1  g0598(.A0(n1303), .A1(n1306), .B0(n1301), .B1(n1297), .Y(n1307));
NOR2X1   g0599(.A(n1307), .B(n1166_1), .Y(n1308));
INVX1    g0600(.A(g594), .Y(n1309));
NOR4X1   g0601(.A(n1309), .B(n1298), .C(g590), .D(n1294), .Y(n1310));
NAND3X1  g0602(.A(n1310), .B(g582), .C(g574), .Y(n1311));
INVX1    g0603(.A(n1311), .Y(n1312));
OAI21X1  g0604(.A0(n1307), .A1(g574), .B0(n1311), .Y(n1313));
XOR2X1   g0605(.A(g594), .B(n1165), .Y(n1314));
OAI22X1  g0606(.A0(n1313), .A1(n1308), .B0(n1312), .B1(n1314), .Y(n391));
INVX1    g0607(.A(g107), .Y(n1316));
NOR3X1   g0608(.A(n783), .B(n1316), .C(g89), .Y(n1317));
INVX1    g0609(.A(g157), .Y(n1318));
NOR2X1   g0610(.A(n788), .B(n1318), .Y(n1319));
MX2X1    g0611(.A(n1319), .B(g148), .S0(n1317), .Y(n396));
MX2X1    g0612(.A(g696), .B(n935), .S0(g269), .Y(n401));
MX2X1    g0613(.A(g449), .B(g453), .S0(n993), .Y(n416));
INVX1    g0614(.A(g117), .Y(n1323));
NOR2X1   g0615(.A(n1071_1), .B(n1323), .Y(n421));
OR4X1    g0616(.A(n1009), .B(n1007), .C(n765), .D(n1010), .Y(n1325));
MX2X1    g0617(.A(g697), .B(g528), .S0(n1325), .Y(n426));
MX2X1    g0618(.A(g426), .B(g422), .S0(n993), .Y(n436));
AND2X1   g0619(.A(g598), .B(g567), .Y(n1328));
XOR2X1   g0620(.A(n1328), .B(n836_1), .Y(n1329));
NOR2X1   g0621(.A(n1329), .B(n1230), .Y(n441));
INVX1    g0622(.A(g669), .Y(n1331));
OAI21X1  g0623(.A0(n221), .A1(g22), .B0(n1331), .Y(n446));
MX2X1    g0624(.A(g695), .B(g520), .S0(n1325), .Y(n451));
NAND4X1  g0625(.A(g279), .B(g276), .C(g278), .D(g277), .Y(n1334));
NOR2X1   g0626(.A(n1334), .B(n868), .Y(n1335));
OAI21X1  g0627(.A0(n1335), .A1(n866_1), .B0(n920), .Y(n1336));
AOI21X1  g0628(.A0(n1335), .A1(n866_1), .B0(n1336), .Y(n1337));
NAND3X1  g0629(.A(n922), .B(n871_1), .C(g269), .Y(n1338));
OAI22X1  g0630(.A0(n1337), .A1(n1338), .B0(g269), .B1(n845), .Y(n456));
INVX1    g0631(.A(g175), .Y(n1340));
NOR2X1   g0632(.A(n788), .B(n1340), .Y(n1341));
MX2X1    g0633(.A(n1341), .B(g166), .S0(n1317), .Y(n461));
NAND2X1  g0634(.A(n1201_1), .B(g554), .Y(n1343));
AOI22X1  g0635(.A0(n1191_1), .A1(g561), .B0(g297), .B1(n1198), .Y(n1344));
NAND2X1  g0636(.A(n1344), .B(n1343), .Y(n1345));
INVX1    g0637(.A(g449), .Y(n1346));
INVX1    g0638(.A(g512), .Y(n1347));
OAI22X1  g0639(.A0(n1182), .A1(n1346), .B0(n1347), .B1(n1204), .Y(n1348));
INVX1    g0640(.A(g541), .Y(n1349));
INVX1    g0641(.A(g414), .Y(n1350));
OAI22X1  g0642(.A0(n1183), .A1(n1350), .B0(n1349), .B1(n1203), .Y(n1351));
NOR3X1   g0643(.A(n1351), .B(n1348), .C(n1345), .Y(n1352));
OAI21X1  g0644(.A0(n1208), .A1(n843), .B0(n1352), .Y(n1353));
AOI21X1  g0645(.A0(n1178), .A1(g693), .B0(n1353), .Y(n1354));
XOR2X1   g0646(.A(n869), .B(g279), .Y(n1355));
AND2X1   g0647(.A(n1355), .B(n1073), .Y(n1356));
NAND2X1  g0648(.A(n920), .B(g269), .Y(n1357));
OAI22X1  g0649(.A0(n1356), .A1(n1357), .B0(g269), .B1(n843), .Y(n821));
NAND2X1  g0650(.A(n765), .B(g693), .Y(n1359));
NAND2X1  g0651(.A(g677), .B(g693), .Y(n1360));
NAND2X1  g0652(.A(n1360), .B(n1359), .Y(n1361));
AOI22X1  g0653(.A0(n821), .A1(n1187), .B0(n770), .B1(n1361), .Y(n1362));
AOI22X1  g0654(.A0(n1186_1), .A1(n166), .B0(n775), .B1(n1361), .Y(n1363));
NAND4X1  g0655(.A(n1362), .B(n1354), .C(n1207), .D(n1363), .Y(n466));
XOR2X1   g0656(.A(n1169), .B(g631), .Y(n1365));
AND2X1   g0657(.A(n1365), .B(g639), .Y(n471));
INVX1    g0658(.A(g386), .Y(n1367));
NAND2X1  g0659(.A(n1031_1), .B(n1030), .Y(n1368));
OR2X1    g0660(.A(n1038), .B(n1030), .Y(n1369));
MX2X1    g0661(.A(n1369), .B(n1368), .S0(n1037), .Y(n1370));
MX2X1    g0662(.A(n1367), .B(n1370), .S0(n1025), .Y(n1371));
XOR2X1   g0663(.A(n1371), .B(g69), .Y(n1372));
MX2X1    g0664(.A(n1028), .B(n1372), .S0(n1026_1), .Y(n1373));
OAI21X1  g0665(.A0(n1373), .A1(n1051_1), .B0(n1055), .Y(n476));
NOR2X1   g0666(.A(g314), .B(n1019), .Y(n486));
MX2X1    g0667(.A(g457), .B(g461), .S0(n993), .Y(n491));
INVX1    g0668(.A(g327), .Y(n1377));
NOR2X1   g0669(.A(n1000), .B(n1377), .Y(n506));
MX2X1    g0670(.A(g418), .B(g414), .S0(n993), .Y(n516));
MX2X1    g0671(.A(g471), .B(g478), .S0(g465), .Y(n1380));
MX2X1    g0672(.A(g402), .B(n1380), .S0(n993), .Y(n521));
OR4X1    g0673(.A(n1007), .B(g683), .C(n792), .D(n1009), .Y(n1382));
MX2X1    g0674(.A(g693), .B(g297), .S0(n1382), .Y(n526));
MX2X1    g0675(.A(g410), .B(g406), .S0(n993), .Y(n536));
MX2X1    g0676(.A(g430), .B(g426), .S0(n993), .Y(n541));
AND2X1   g0677(.A(n943), .B(g697), .Y(n1386));
INVX1    g0678(.A(g528), .Y(n1387));
NOR3X1   g0679(.A(n1202), .B(n765), .C(n1387), .Y(n1388));
AND2X1   g0680(.A(n1191_1), .B(g557), .Y(n1389));
INVX1    g0681(.A(g430), .Y(n1390));
INVX1    g0682(.A(g434), .Y(n1391));
OAI22X1  g0683(.A0(n1182), .A1(n1391), .B0(n1390), .B1(n1183), .Y(n1392));
NOR3X1   g0684(.A(n1392), .B(n1389), .C(n1388), .Y(n1393));
OAI21X1  g0685(.A0(n1271), .A1(n835), .B0(n1393), .Y(n1394));
NAND2X1  g0686(.A(n765), .B(g697), .Y(n1395));
NAND2X1  g0687(.A(g677), .B(g697), .Y(n1396));
AOI22X1  g0688(.A0(n1395), .A1(n1396), .B0(n776_1), .B1(n771_1), .Y(n1397));
NOR3X1   g0689(.A(n1397), .B(n1394), .C(n1386), .Y(n1398));
NOR4X1   g0690(.A(n921_1), .B(n918), .C(n915), .D(n905), .Y(n1399));
OAI21X1  g0691(.A0(n902), .A1(n901_1), .B0(g478), .Y(n1400));
NAND3X1  g0692(.A(n888), .B(n887), .C(n872), .Y(n1401));
INVX1    g0693(.A(n908), .Y(n1402));
AOI21X1  g0694(.A0(n1401), .A1(n1400), .B0(n1402), .Y(n1403));
OAI21X1  g0695(.A0(n913), .A1(n1403), .B0(n871_1), .Y(n1404));
OR2X1    g0696(.A(n917), .B(n870), .Y(n1405));
NAND2X1  g0697(.A(n929), .B(n917), .Y(n1406));
NAND3X1  g0698(.A(n1406), .B(n1405), .C(n1404), .Y(n1407));
OAI21X1  g0699(.A0(n1407), .A1(n1399), .B0(g269), .Y(n1408));
NOR2X1   g0700(.A(g269), .B(n835), .Y(n1409));
INVX1    g0701(.A(n1409), .Y(n1410));
NAND2X1  g0702(.A(n1410), .B(n1408), .Y(n776));
OAI21X1  g0703(.A0(n1114), .A1(n1113), .B0(g471), .Y(n1412));
NAND3X1  g0704(.A(n1100), .B(n1099), .C(n965), .Y(n1413));
NAND3X1  g0705(.A(n969), .B(g210), .C(n966_1), .Y(n1414));
AOI21X1  g0706(.A0(n1413), .A1(n1412), .B0(n1414), .Y(n1415));
AND2X1   g0707(.A(n1415), .B(n1122), .Y(n1416));
NAND2X1  g0708(.A(n967), .B(g211), .Y(n1417));
OAI21X1  g0709(.A0(n1417), .A1(n964), .B0(n975), .Y(n1418));
NAND2X1  g0710(.A(g210), .B(n966_1), .Y(n1419));
OR2X1    g0711(.A(n1419), .B(n969), .Y(n1420));
OAI21X1  g0712(.A0(n1420), .A1(n1119), .B0(n971_1), .Y(n1421));
NOR4X1   g0713(.A(n1418), .B(n1416), .C(n1121_1), .D(n966_1), .Y(n1423));
AND2X1   g0714(.A(n1415), .B(n964), .Y(n1424));
NOR3X1   g0715(.A(n1415), .B(n1419), .C(n964), .Y(n1425));
OR4X1    g0716(.A(n1424), .B(n1423), .C(n1123), .D(n1425), .Y(n1426));
MX2X1    g0717(.A(g697), .B(n1426), .S0(g197), .Y(n586));
AOI22X1  g0718(.A0(n776), .A1(n1187), .B0(n1186_1), .B1(n586), .Y(n1428));
NAND3X1  g0719(.A(n1428), .B(n1398), .C(n1207), .Y(n546));
INVX1    g0720(.A(g266), .Y(n551));
MX2X1    g0721(.A(g453), .B(g457), .S0(n993), .Y(n556));
MX2X1    g0722(.A(g691), .B(g269), .S0(n1382), .Y(n561));
XOR2X1   g0723(.A(n1171_1), .B(g574), .Y(n1433));
NAND2X1  g0724(.A(n1433), .B(n1173), .Y(n566));
MX2X1    g0725(.A(g441), .B(g445), .S0(n993), .Y(n571));
INVX1    g0726(.A(n755), .Y(n1436));
AND2X1   g0727(.A(n1436), .B(n751_1), .Y(n1437));
INVX1    g0728(.A(n1437), .Y(n1438));
NOR3X1   g0729(.A(g345), .B(g341), .C(g338), .Y(n1439));
XOR2X1   g0730(.A(n1439), .B(g349), .Y(n1440));
MX2X1    g0731(.A(g349), .B(n1440), .S0(g323), .Y(n1441));
OR2X1    g0732(.A(n1441), .B(n1438), .Y(n581));
NAND4X1  g0733(.A(g582), .B(g578), .C(g631), .D(n1169), .Y(n1443));
XOR2X1   g0734(.A(n1443), .B(n1298), .Y(n1444));
AND2X1   g0735(.A(n1444), .B(n1173), .Y(n591));
INVX1    g0736(.A(g571), .Y(n1446));
INVX1    g0737(.A(g646), .Y(n1447));
INVX1    g0738(.A(g650), .Y(n1448));
NOR4X1   g0739(.A(n1448), .B(n1447), .C(n1240), .D(n1231), .Y(n1449));
AND2X1   g0740(.A(n1449), .B(g654), .Y(n1450));
XOR2X1   g0741(.A(n1450), .B(n1446), .Y(n1451));
NOR2X1   g0742(.A(n1451), .B(n1230), .Y(n596));
AND2X1   g0743(.A(n943), .B(g696), .Y(n1453));
INVX1    g0744(.A(g524), .Y(n1454));
NOR3X1   g0745(.A(n1202), .B(n765), .C(n1454), .Y(n1455));
AND2X1   g0746(.A(n1191_1), .B(g558), .Y(n1456));
INVX1    g0747(.A(g437), .Y(n1457));
INVX1    g0748(.A(g426), .Y(n1458));
OAI22X1  g0749(.A0(n1182), .A1(n1457), .B0(n1458), .B1(n1183), .Y(n1459));
NOR3X1   g0750(.A(n1459), .B(n1456), .C(n1455), .Y(n1460));
OAI21X1  g0751(.A0(n1271), .A1(n847), .B0(n1460), .Y(n1461));
NAND2X1  g0752(.A(n765), .B(g696), .Y(n1462));
NAND2X1  g0753(.A(g677), .B(g696), .Y(n1463));
AOI22X1  g0754(.A0(n1462), .A1(n1463), .B0(n776_1), .B1(n771_1), .Y(n1464));
NOR3X1   g0755(.A(n1464), .B(n1461), .C(n1453), .Y(n1465));
NOR4X1   g0756(.A(n1421), .B(n1123), .C(n967), .D(n1424), .Y(n1466));
OR4X1    g0757(.A(n1418), .B(n1416), .C(n1121_1), .D(n1425), .Y(n1467));
OR2X1    g0758(.A(n1467), .B(n1466), .Y(n1468));
MX2X1    g0759(.A(g696), .B(n1468), .S0(g197), .Y(n971));
AOI22X1  g0760(.A0(n401), .A1(n1187), .B0(n1186_1), .B1(n971), .Y(n1470));
NAND3X1  g0761(.A(n1470), .B(n1465), .C(n1207), .Y(n601));
OR2X1    g0762(.A(n1000), .B(g323), .Y(n606));
INVX1    g0763(.A(g654), .Y(n1473));
XOR2X1   g0764(.A(n1449), .B(n1473), .Y(n1474));
NOR2X1   g0765(.A(n1474), .B(n1230), .Y(n616));
MX2X1    g0766(.A(g692), .B(g293), .S0(n1382), .Y(n621));
MX2X1    g0767(.A(g445), .B(g449), .S0(n993), .Y(n631));
INVX1    g0768(.A(g374), .Y(n1478));
NOR2X1   g0769(.A(n755), .B(n1478), .Y(n1479));
MX2X1    g0770(.A(g370), .B(n1479), .S0(n1253), .Y(n636));
NAND2X1  g0771(.A(n995), .B(g11), .Y(n1481));
NAND2X1  g0772(.A(n729), .B(g11), .Y(n1482));
NAND2X1  g0773(.A(n1482), .B(n1481), .Y(n641));
AND2X1   g0774(.A(n750), .B(n749), .Y(n1484));
XOR2X1   g0775(.A(n1484), .B(n748), .Y(n1485));
MX2X1    g0776(.A(n748), .B(n1485), .S0(g323), .Y(n1486));
NAND2X1  g0777(.A(n1486), .B(n1437), .Y(n651));
NOR2X1   g0778(.A(n755), .B(n1367), .Y(n1488));
MX2X1    g0779(.A(g382), .B(n1488), .S0(n1253), .Y(n656));
MX2X1    g0780(.A(g691), .B(g504), .S0(n1325), .Y(n661));
INVX1    g0781(.A(g166), .Y(n1491));
NOR2X1   g0782(.A(n788), .B(n1491), .Y(n1492));
MX2X1    g0783(.A(n1492), .B(g157), .S0(n1317), .Y(n671));
INVX1    g0784(.A(g465), .Y(n1494));
MX2X1    g0785(.A(n870), .B(n1122), .S0(n1494), .Y(n1495));
NAND3X1  g0786(.A(n1495), .B(n991_1), .C(n1213), .Y(n1496));
NAND2X1  g0787(.A(n1496), .B(n1349), .Y(n1497));
MX2X1    g0788(.A(n1497), .B(g693), .S0(n1011_1), .Y(n676));
NAND3X1  g0789(.A(n1031_1), .B(n1030), .C(n1028), .Y(n1499));
INVX1    g0790(.A(g59), .Y(n1500));
NAND3X1  g0791(.A(g49), .B(g54), .C(g361), .Y(n1501));
OR4X1    g0792(.A(n1500), .B(n1030), .C(n1028), .D(n1501), .Y(n1502));
MX2X1    g0793(.A(n1502), .B(n1499), .S0(n1037), .Y(n1503));
MX2X1    g0794(.A(n1262), .B(n1503), .S0(n1025), .Y(n1504));
XOR2X1   g0795(.A(n1504), .B(g74), .Y(n1505));
MX2X1    g0796(.A(n1029), .B(n1505), .S0(n1026_1), .Y(n1506));
OAI21X1  g0797(.A0(n1506), .A1(n1051_1), .B0(n1055), .Y(n681));
XOR2X1   g0798(.A(g338), .B(g323), .Y(n1508));
OR2X1    g0799(.A(n1508), .B(n1438), .Y(n686));
MX2X1    g0800(.A(g694), .B(g516), .S0(n1325), .Y(n696));
MX2X1    g0801(.A(n910), .B(n968), .S0(n1494), .Y(n1511));
AOI21X1  g0802(.A0(n1511), .A1(n991_1), .B0(n1213), .Y(n1512));
MX2X1    g0803(.A(n1512), .B(g692), .S0(n1011_1), .Y(n701));
XOR2X1   g0804(.A(n750), .B(g353), .Y(n1514));
MX2X1    g0805(.A(g353), .B(n1514), .S0(g323), .Y(n1515));
AND2X1   g0806(.A(n1515), .B(n1437), .Y(n711));
MX2X1    g0807(.A(n1468), .B(g545), .S0(n992), .Y(n716));
INVX1    g0808(.A(g341), .Y(n1518));
XOR2X1   g0809(.A(g341), .B(g338), .Y(n1519));
MX2X1    g0810(.A(n1518), .B(n1519), .S0(g323), .Y(n1520));
NAND3X1  g0811(.A(n1520), .B(n1436), .C(n751_1), .Y(n726));
NAND2X1  g0812(.A(n995), .B(g7), .Y(n1522));
NAND2X1  g0813(.A(n729), .B(g7), .Y(n1523));
NAND2X1  g0814(.A(n1523), .B(n1522), .Y(n736));
AOI22X1  g0815(.A0(g314), .A1(g310), .B0(g301), .B1(g319), .Y(n1525));
INVX1    g0816(.A(n1525), .Y(n1526));
OAI21X1  g0817(.A0(n1526), .A1(n1021_1), .B0(n1017), .Y(n1527));
NAND3X1  g0818(.A(g332), .B(n1020), .C(g306), .Y(n1528));
AND2X1   g0819(.A(n1528), .B(n1527), .Y(n1529));
INVX1    g0820(.A(n1529), .Y(n1530));
AOI21X1  g0821(.A0(n1410), .A1(n1408), .B0(n1530), .Y(n1531));
INVX1    g0822(.A(g269), .Y(n1532));
AOI21X1  g0823(.A0(n931_1), .A1(n926_1), .B0(n1532), .Y(n1533));
NOR3X1   g0824(.A(n1529), .B(n1409), .C(n1533), .Y(n1534));
OAI21X1  g0825(.A0(g314), .A1(n1015), .B0(n1525), .Y(n1535));
NOR3X1   g0826(.A(n1535), .B(n1053), .C(n1024), .Y(n1536));
NOR4X1   g0827(.A(n486), .B(n1034), .C(n999), .D(n1536), .Y(n1537));
OAI21X1  g0828(.A0(n1534), .A1(n1531), .B0(n1537), .Y(n1538));
MX2X1    g0829(.A(n1034), .B(n1538), .S0(g336), .Y(n1539));
OR4X1    g0830(.A(g698), .B(g269), .C(g689), .D(g688), .Y(n1540));
NOR3X1   g0831(.A(n1540), .B(n938), .C(n757), .Y(n1541));
AND2X1   g0832(.A(g269), .B(g662), .Y(n1542));
NOR3X1   g0833(.A(n1542), .B(n1541), .C(n1187), .Y(n1543));
OR4X1    g0834(.A(g688), .B(g698), .C(g689), .D(g197), .Y(n1544));
NOR3X1   g0835(.A(n1544), .B(n938), .C(g687), .Y(n1545));
INVX1    g0836(.A(g197), .Y(n1546));
AOI21X1  g0837(.A0(n768), .A1(n761_1), .B0(n1546), .Y(n1547));
NOR3X1   g0838(.A(n1547), .B(n1545), .C(n1186_1), .Y(n1548));
MX2X1    g0839(.A(n1446), .B(n955), .S0(n760), .Y(n1549));
MX2X1    g0840(.A(n954), .B(n1549), .S0(g197), .Y(n1550));
OAI21X1  g0841(.A0(n1548), .A1(g337), .B0(n1550), .Y(n1551));
MX2X1    g0842(.A(n1241), .B(n827), .S0(n760), .Y(n1552));
NAND2X1  g0843(.A(n1546), .B(g681), .Y(n1553));
OAI21X1  g0844(.A0(n1552), .A1(n1546), .B0(n1553), .Y(n1554));
MX2X1    g0845(.A(n812), .B(n836_1), .S0(g658), .Y(n1555));
NAND2X1  g0846(.A(n1546), .B(g680), .Y(n1556));
OAI21X1  g0847(.A0(n1555), .A1(n1546), .B0(n1556), .Y(n1557));
MX2X1    g0848(.A(n834), .B(n806_1), .S0(n760), .Y(n1558));
NAND2X1  g0849(.A(n1546), .B(g679), .Y(n1559));
OAI21X1  g0850(.A0(n1558), .A1(n1546), .B0(n1559), .Y(n1560));
MX2X1    g0851(.A(n831_1), .B(n803), .S0(n760), .Y(n1561));
NAND2X1  g0852(.A(n1546), .B(g678), .Y(n1562));
OAI21X1  g0853(.A0(n1561), .A1(n1546), .B0(n1562), .Y(n1563));
AOI22X1  g0854(.A0(n1560), .A1(n1563), .B0(n1557), .B1(n1554), .Y(n1564));
MX2X1    g0855(.A(n1473), .B(n790), .S0(n760), .Y(n1565));
NAND2X1  g0856(.A(n1546), .B(g685), .Y(n1566));
OAI21X1  g0857(.A0(n1565), .A1(n1546), .B0(n1566), .Y(n1567));
MX2X1    g0858(.A(n793), .B(n1448), .S0(g658), .Y(n1568));
NAND2X1  g0859(.A(n1546), .B(g684), .Y(n1569));
OAI21X1  g0860(.A0(n1568), .A1(n1546), .B0(n1569), .Y(n1570));
MX2X1    g0861(.A(n1447), .B(n796_1), .S0(n760), .Y(n1571));
NAND2X1  g0862(.A(n1546), .B(g683), .Y(n1572));
OAI21X1  g0863(.A0(n1571), .A1(n1546), .B0(n1572), .Y(n1573));
MX2X1    g0864(.A(n1240), .B(n799), .S0(n760), .Y(n1574));
NAND2X1  g0865(.A(n1546), .B(g682), .Y(n1575));
OAI21X1  g0866(.A0(n1574), .A1(n1546), .B0(n1575), .Y(n1576));
AOI22X1  g0867(.A0(n1573), .A1(n1576), .B0(n1570), .B1(n1567), .Y(n1577));
NOR2X1   g0868(.A(n1577), .B(n1564), .Y(n1578));
AND2X1   g0869(.A(n1578), .B(n1551), .Y(n1579));
MX2X1    g0870(.A(n954), .B(n1549), .S0(g269), .Y(n1580));
OAI22X1  g0871(.A0(n1579), .A1(n1580), .B0(n1543), .B1(g337), .Y(n1581));
MX2X1    g0872(.A(n826_1), .B(n1552), .S0(g269), .Y(n1582));
MX2X1    g0873(.A(n813), .B(n1555), .S0(g269), .Y(n1583));
MX2X1    g0874(.A(n805), .B(n1558), .S0(g269), .Y(n1584));
MX2X1    g0875(.A(n802), .B(n1561), .S0(g269), .Y(n1585));
OAI22X1  g0876(.A0(n1584), .A1(n1585), .B0(n1583), .B1(n1582), .Y(n1586));
MX2X1    g0877(.A(n789), .B(n1565), .S0(g269), .Y(n1587));
MX2X1    g0878(.A(n792), .B(n1568), .S0(g269), .Y(n1588));
MX2X1    g0879(.A(n795), .B(n1571), .S0(g269), .Y(n1589));
MX2X1    g0880(.A(n798), .B(n1574), .S0(g269), .Y(n1590));
OAI22X1  g0881(.A0(n1589), .A1(n1590), .B0(n1588), .B1(n1587), .Y(n1591));
NAND3X1  g0882(.A(n1591), .B(n1586), .C(n1581), .Y(n1592));
MX2X1    g0883(.A(n1539), .B(n1592), .S0(n755), .Y(n746));
NOR2X1   g0884(.A(g341), .B(g338), .Y(n1594));
XOR2X1   g0885(.A(n1594), .B(g345), .Y(n1595));
MX2X1    g0886(.A(g345), .B(n1595), .S0(g323), .Y(n1596));
OR2X1    g0887(.A(n1596), .B(n1438), .Y(n751));
XOR2X1   g0888(.A(n1168), .B(g628), .Y(n1598));
AND2X1   g0889(.A(n1598), .B(g639), .Y(n756));
NAND2X1  g0890(.A(n995), .B(g33), .Y(n1600));
NAND2X1  g0891(.A(n729), .B(g33), .Y(n1601));
NAND2X1  g0892(.A(n1601), .B(n1600), .Y(n766));
NAND2X1  g0893(.A(g610), .B(g602), .Y(n1603));
XOR2X1   g0894(.A(n1603), .B(g613), .Y(n1604));
NAND2X1  g0895(.A(n1604), .B(g639), .Y(n781));
NAND2X1  g0896(.A(n995), .B(g15), .Y(n1606));
NAND2X1  g0897(.A(n729), .B(g15), .Y(n1607));
NAND2X1  g0898(.A(n1607), .B(n1606), .Y(n786));
NAND2X1  g0899(.A(n995), .B(g19), .Y(n1609));
NAND2X1  g0900(.A(n729), .B(g19), .Y(n1610));
NAND2X1  g0901(.A(n1610), .B(n1609), .Y(n791));
INVX1    g0902(.A(g143), .Y(n1612));
NOR2X1   g0903(.A(n1135), .B(g148), .Y(n1613));
XOR2X1   g0904(.A(n1613), .B(g143), .Y(n1614));
MX2X1    g0905(.A(n1612), .B(n1614), .S0(n1136_1), .Y(n1615));
OAI21X1  g0906(.A0(n1615), .A1(n1156_1), .B0(n1160), .Y(n801));
NOR3X1   g0907(.A(n726_1), .B(n724), .C(g22), .Y(n1617));
OR2X1    g0908(.A(n1617), .B(g672), .Y(n806));
MX2X1    g0909(.A(g398), .B(g366), .S0(n1253), .Y(n1619));
OR2X1    g0910(.A(n1619), .B(n755), .Y(n816));
NOR2X1   g0911(.A(n915), .B(g492), .Y(n1621));
NAND2X1  g0912(.A(n1621), .B(n1404), .Y(n826));
INVX1    g0913(.A(g170), .Y(n1623));
OR2X1    g0914(.A(g152), .B(g143), .Y(n1624));
OR2X1    g0915(.A(n1624), .B(g161), .Y(n1625));
NAND3X1  g0916(.A(g161), .B(g152), .C(g143), .Y(n1626));
MX2X1    g0917(.A(n1626), .B(n1625), .S0(n1143), .Y(n1627));
MX2X1    g0918(.A(n1340), .B(n1627), .S0(n1135), .Y(n1628));
XOR2X1   g0919(.A(n1628), .B(g170), .Y(n1629));
MX2X1    g0920(.A(n1623), .B(n1629), .S0(n1136_1), .Y(n1630));
OAI21X1  g0921(.A0(n1630), .A1(n1156_1), .B0(n1160), .Y(n831));
NOR2X1   g0922(.A(g602), .B(n1064), .Y(n851));
XOR2X1   g0923(.A(n1242), .B(g642), .Y(n1633));
NOR2X1   g0924(.A(n1633), .B(n1230), .Y(n856));
XOR2X1   g0925(.A(n1334), .B(g280), .Y(n1635));
NAND4X1  g0926(.A(n922), .B(n920), .C(n871_1), .D(n1635), .Y(n1636));
MX2X1    g0927(.A(g694), .B(n1636), .S0(g269), .Y(n861));
XOR2X1   g0928(.A(g610), .B(g602), .Y(n1638));
AND2X1   g0929(.A(n1638), .B(g639), .Y(n871));
MX2X1    g0930(.A(g148), .B(g193), .S0(n1317), .Y(n1640));
OR2X1    g0931(.A(n1640), .B(n788), .Y(n876));
NOR2X1   g0932(.A(n1258), .B(n961_1), .Y(n1642));
OAI21X1  g0933(.A0(n1642), .A1(n962), .B0(n975), .Y(n1643));
AOI21X1  g0934(.A0(n1642), .A1(n962), .B0(n1643), .Y(n1644));
NAND3X1  g0935(.A(n971_1), .B(n964), .C(g197), .Y(n1645));
OAI22X1  g0936(.A0(n1644), .A1(n1645), .B0(g197), .B1(n845), .Y(n881));
INVX1    g0937(.A(g119), .Y(n1647));
NOR2X1   g0938(.A(n1071_1), .B(n1647), .Y(n896));
INVX1    g0939(.A(g54), .Y(n1649));
OR2X1    g0940(.A(g49), .B(g361), .Y(n1650));
NAND2X1  g0941(.A(g49), .B(g361), .Y(n1651));
MX2X1    g0942(.A(n1651), .B(n1650), .S0(n1037), .Y(n1652));
MX2X1    g0943(.A(n1478), .B(n1652), .S0(n1025), .Y(n1653));
XOR2X1   g0944(.A(n1653), .B(g54), .Y(n1654));
MX2X1    g0945(.A(n1649), .B(n1654), .S0(n1026_1), .Y(n1655));
OAI21X1  g0946(.A0(n1655), .A1(n1051_1), .B0(n1055), .Y(n901));
XOR2X1   g0947(.A(n1172), .B(g594), .Y(n1657));
AND2X1   g0948(.A(n1657), .B(n1173), .Y(n906));
NAND3X1  g0949(.A(g610), .B(g602), .C(g613), .Y(n1659));
XOR2X1   g0950(.A(n1659), .B(g616), .Y(n1660));
NOR2X1   g0951(.A(n1660), .B(n1064), .Y(n921));
INVX1    g0952(.A(g394), .Y(n1662));
MX2X1    g0953(.A(n1048), .B(n1032), .S0(n1037), .Y(n1663));
MX2X1    g0954(.A(n1662), .B(n1663), .S0(n1025), .Y(n1664));
XOR2X1   g0955(.A(n1664), .B(g79), .Y(n1665));
MX2X1    g0956(.A(n1047), .B(n1665), .S0(n1026_1), .Y(n1666));
OAI21X1  g0957(.A0(n1666), .A1(n1051_1), .B0(n1055), .Y(n926));
XOR2X1   g0958(.A(n1170), .B(g578), .Y(n1668));
AND2X1   g0959(.A(n1668), .B(n1173), .Y(n941));
NOR2X1   g0960(.A(n788), .B(n1137), .Y(n1670));
MX2X1    g0961(.A(n1670), .B(g175), .S0(n1317), .Y(n946));
INVX1    g0962(.A(g118), .Y(n1672));
NOR2X1   g0963(.A(n1071_1), .B(n1672), .Y(n951));
NAND2X1  g0964(.A(n1468), .B(n1426), .Y(n956));
AND2X1   g0965(.A(n1078), .B(n783), .Y(n1675));
XOR2X1   g0966(.A(n782), .B(n781_1), .Y(n1676));
MX2X1    g0967(.A(n781_1), .B(n1676), .S0(g114), .Y(n1677));
NAND2X1  g0968(.A(n1677), .B(n1675), .Y(n961));
MX2X1    g0969(.A(g422), .B(g418), .S0(n993), .Y(n966));
NOR2X1   g0970(.A(n755), .B(n1662), .Y(n1680));
MX2X1    g0971(.A(g390), .B(n1680), .S0(n1253), .Y(n976));
AND2X1   g0972(.A(n943), .B(g695), .Y(n1682));
AND2X1   g0973(.A(n1178), .B(g695), .Y(n1683));
INVX1    g0974(.A(g520), .Y(n1684));
NAND2X1  g0975(.A(n1191_1), .B(g559), .Y(n1685));
OAI21X1  g0976(.A0(n1204), .A1(n1684), .B0(n1685), .Y(n1686));
INVX1    g0977(.A(g441), .Y(n1687));
INVX1    g0978(.A(g422), .Y(n1688));
OAI22X1  g0979(.A0(n1182), .A1(n1687), .B0(n1688), .B1(n1183), .Y(n1689));
NOR4X1   g0980(.A(n1686), .B(n1683), .C(n1682), .D(n1689), .Y(n1690));
NAND2X1  g0981(.A(n765), .B(g695), .Y(n1691));
NAND2X1  g0982(.A(g677), .B(g695), .Y(n1692));
NAND2X1  g0983(.A(n1692), .B(n1691), .Y(n1693));
AOI22X1  g0984(.A0(n456), .A1(n1187), .B0(n770), .B1(n1693), .Y(n1694));
AOI22X1  g0985(.A0(n881), .A1(n1186_1), .B0(n775), .B1(n1693), .Y(n1695));
NAND4X1  g0986(.A(n1694), .B(n1690), .C(n1207), .D(n1695), .Y(n986));
INVX1    g0987(.A(g45), .Y(n1697));
NOR2X1   g0988(.A(g658), .B(n1697), .Y(n996));
NOR3X1   g0989(.A(n1231), .B(n1447), .C(n1240), .Y(n1699));
XOR2X1   g0990(.A(n1699), .B(n1448), .Y(n1700));
NOR2X1   g0991(.A(n1700), .B(n1230), .Y(n1001));
INVX1    g0992(.A(g378), .Y(n1702));
NOR2X1   g0993(.A(n755), .B(n1702), .Y(n1703));
MX2X1    g0994(.A(g374), .B(n1703), .S0(n1253), .Y(n1006));
MX2X1    g0995(.A(g692), .B(g508), .S0(n1325), .Y(n1011));
MX2X1    g0996(.A(n1426), .B(g548), .S0(n992), .Y(n1016));
INVX1    g0997(.A(g370), .Y(n1707));
NOR2X1   g0998(.A(n755), .B(n1707), .Y(n1708));
MX2X1    g0999(.A(g366), .B(n1708), .S0(n1253), .Y(n1021));
MX2X1    g1000(.A(g406), .B(g402), .S0(n993), .Y(n1026));
MX2X1    g1001(.A(g690), .B(g500), .S0(n1325), .Y(n1036));
XOR2X1   g1002(.A(g205), .B(g204), .Y(n1712));
NAND4X1  g1003(.A(n975), .B(n972), .C(g197), .D(n1712), .Y(n1713));
OAI21X1  g1004(.A0(n916), .A1(g197), .B0(n1713), .Y(n1041));
MX2X1    g1005(.A(g690), .B(g197), .S0(n1382), .Y(n1046));
INVX1    g1006(.A(g122), .Y(n1716));
NOR2X1   g1007(.A(n1071_1), .B(n1716), .Y(n1056));
MX2X1    g1008(.A(g696), .B(g524), .S0(n1325), .Y(n1061));
OR4X1    g1009(.A(g107), .B(n1130), .C(n708), .D(n1157), .Y(n1719));
XOR2X1   g1010(.A(n1719), .B(g111), .Y(n1720));
NOR2X1   g1011(.A(n1720), .B(n788), .Y(n1071));
INVX1    g1012(.A(g131), .Y(n1722));
XOR2X1   g1013(.A(g131), .B(g128), .Y(n1723));
MX2X1    g1014(.A(n1722), .B(n1723), .S0(g114), .Y(n1724));
NAND3X1  g1015(.A(n1724), .B(n1078), .C(n783), .Y(n1076));
AOI22X1  g1016(.A0(n1191_1), .A1(g563), .B0(g492), .B1(n1194), .Y(n1726));
AOI22X1  g1017(.A0(n1193), .A1(n711_1), .B0(g672), .B1(n1196_1), .Y(n1727));
AOI22X1  g1018(.A0(n1198), .A1(g269), .B0(g548), .B1(n1201_1), .Y(n1728));
NAND3X1  g1019(.A(n1728), .B(n1727), .C(n1726), .Y(n1729));
INVX1    g1020(.A(g504), .Y(n1730));
OAI22X1  g1021(.A0(n1203), .A1(n1494), .B0(n1730), .B1(n1204), .Y(n1731));
INVX1    g1022(.A(g457), .Y(n1732));
INVX1    g1023(.A(g406), .Y(n1733));
OAI22X1  g1024(.A0(n1182), .A1(n1732), .B0(n1733), .B1(n1183), .Y(n1734));
NOR3X1   g1025(.A(n1734), .B(n1731), .C(n1729), .Y(n1735));
OAI21X1  g1026(.A0(n1208), .A1(n916), .B0(n1735), .Y(n1736));
AOI21X1  g1027(.A0(n1178), .A1(g691), .B0(n1736), .Y(n1737));
XOR2X1   g1028(.A(g277), .B(g276), .Y(n1738));
NAND4X1  g1029(.A(n1073), .B(n920), .C(g269), .D(n1738), .Y(n1739));
OAI21X1  g1030(.A0(n916), .A1(g269), .B0(n1739), .Y(n1156));
NAND2X1  g1031(.A(g691), .B(n765), .Y(n1741));
NAND2X1  g1032(.A(g691), .B(g677), .Y(n1742));
NAND2X1  g1033(.A(n1742), .B(n1741), .Y(n1743));
AOI22X1  g1034(.A0(n1156), .A1(n1187), .B0(n770), .B1(n1743), .Y(n1744));
AOI22X1  g1035(.A0(n1041), .A1(n1186_1), .B0(n775), .B1(n1743), .Y(n1745));
NAND4X1  g1036(.A(n1744), .B(n1737), .C(n1207), .D(n1745), .Y(n1081));
AND2X1   g1037(.A(n943), .B(g694), .Y(n1747));
AND2X1   g1038(.A(n1178), .B(g694), .Y(n1748));
INVX1    g1039(.A(g516), .Y(n1749));
NAND2X1  g1040(.A(n1191_1), .B(g560), .Y(n1750));
OAI21X1  g1041(.A0(n1204), .A1(n1749), .B0(n1750), .Y(n1751));
INVX1    g1042(.A(g418), .Y(n1752));
INVX1    g1043(.A(g445), .Y(n1753));
OAI22X1  g1044(.A0(n1182), .A1(n1753), .B0(n1752), .B1(n1183), .Y(n1754));
NOR4X1   g1045(.A(n1751), .B(n1748), .C(n1747), .D(n1754), .Y(n1755));
NAND2X1  g1046(.A(g694), .B(n765), .Y(n1756));
NAND2X1  g1047(.A(g694), .B(g677), .Y(n1757));
NAND2X1  g1048(.A(n1757), .B(n1756), .Y(n1758));
AOI22X1  g1049(.A0(n861), .A1(n1187), .B0(n770), .B1(n1758), .Y(n1759));
AOI22X1  g1050(.A0(n336), .A1(n1186_1), .B0(n775), .B1(n1758), .Y(n1760));
NAND4X1  g1051(.A(n1759), .B(n1755), .C(n1207), .D(n1760), .Y(n1086));
AND2X1   g1052(.A(n1170), .B(g578), .Y(n1762));
XOR2X1   g1053(.A(n1762), .B(g582), .Y(n1763));
AND2X1   g1054(.A(n1763), .B(n1173), .Y(n1096));
NAND2X1  g1055(.A(n935), .B(n932), .Y(n1101));
INVX1    g1056(.A(g47), .Y(n1106));
NOR2X1   g1057(.A(n788), .B(n1234), .Y(n1767));
MX2X1    g1058(.A(n1767), .B(g184), .S0(n1317), .Y(n1111));
INVX1    g1059(.A(g135), .Y(n1769));
NOR2X1   g1060(.A(g131), .B(g128), .Y(n1770));
XOR2X1   g1061(.A(n1770), .B(n1769), .Y(n1771));
MX2X1    g1062(.A(n1769), .B(n1771), .S0(g114), .Y(n1772));
NAND2X1  g1063(.A(n1772), .B(n1675), .Y(n1116));
INVX1    g1064(.A(g382), .Y(n1774));
NOR2X1   g1065(.A(n755), .B(n1774), .Y(n1775));
MX2X1    g1066(.A(g378), .B(n1775), .S0(n1253), .Y(n1121));
MX2X1    g1067(.A(g414), .B(g410), .S0(n993), .Y(n1126));
MX2X1    g1068(.A(g434), .B(g437), .S0(n993), .Y(n1131));
NOR2X1   g1069(.A(g266), .B(n1697), .Y(n1136));
INVX1    g1070(.A(g49), .Y(n1780));
XOR2X1   g1071(.A(n1037), .B(n1248), .Y(n1781));
MX2X1    g1072(.A(n1707), .B(n1781), .S0(n1025), .Y(n1782));
XOR2X1   g1073(.A(n1782), .B(g49), .Y(n1783));
MX2X1    g1074(.A(n1780), .B(n1783), .S0(n1026_1), .Y(n1784));
OAI21X1  g1075(.A0(n1784), .A1(n1051_1), .B0(n1055), .Y(n1141));
INVX1    g1076(.A(g152), .Y(n1786));
XOR2X1   g1077(.A(n1143), .B(n1612), .Y(n1787));
MX2X1    g1078(.A(n1318), .B(n1787), .S0(n1135), .Y(n1788));
XOR2X1   g1079(.A(n1788), .B(g152), .Y(n1789));
MX2X1    g1080(.A(n1786), .B(n1789), .S0(n1136_1), .Y(n1790));
OAI21X1  g1081(.A0(n1790), .A1(n1156_1), .B0(n1160), .Y(n1146));
INVX1    g1082(.A(g127), .Y(n1792));
NOR2X1   g1083(.A(g102), .B(n1127), .Y(n1793));
OAI22X1  g1084(.A0(n1130), .A1(n1128), .B0(n708), .B1(n1316), .Y(n1794));
OR2X1    g1085(.A(n1794), .B(n1131_1), .Y(n1795));
MX2X1    g1086(.A(n1793), .B(n1795), .S0(n780), .Y(n1796));
XOR2X1   g1087(.A(n1796), .B(g697), .Y(n1797));
NOR4X1   g1088(.A(n1159), .B(n1134), .C(n1793), .D(n1794), .Y(n1798));
NOR4X1   g1089(.A(g102), .B(n1128), .C(g94), .D(g111), .Y(n1799));
NOR4X1   g1090(.A(n1798), .B(g2584), .C(n1647), .D(n1799), .Y(n1800));
AOI21X1  g1091(.A0(n1800), .A1(n1797), .B0(n1792), .Y(n1801));
AND2X1   g1092(.A(n1799), .B(n1792), .Y(n1802));
OAI21X1  g1093(.A0(n1802), .A1(n1801), .B0(n1078), .Y(n1803));
NOR4X1   g1094(.A(n938), .B(n808), .C(g687), .D(n809), .Y(n1804));
AOI21X1  g1095(.A0(n767), .A1(g293), .B0(n1804), .Y(n1805));
NOR4X1   g1096(.A(n814), .B(n807), .C(n820), .D(n1805), .Y(n1806));
NOR4X1   g1097(.A(n817), .B(n816_1), .C(n820), .D(n1805), .Y(n1807));
NOR4X1   g1098(.A(n814), .B(n816_1), .C(n804), .D(n1805), .Y(n1808));
NOR4X1   g1099(.A(n814), .B(n807), .C(n804), .D(n1805), .Y(n1809));
NOR4X1   g1100(.A(n1808), .B(n1807), .C(n1806), .D(n1809), .Y(n1810));
NOR4X1   g1101(.A(n814), .B(n816_1), .C(n820), .D(n1805), .Y(n1811));
NOR4X1   g1102(.A(n817), .B(n807), .C(n820), .D(n1805), .Y(n1812));
NOR4X1   g1103(.A(n817), .B(n816_1), .C(n804), .D(n1805), .Y(n1813));
NOR4X1   g1104(.A(n817), .B(n807), .C(n804), .D(n1805), .Y(n1814));
NOR4X1   g1105(.A(n1813), .B(n1812), .C(n1811), .D(n1814), .Y(n1815));
NAND2X1  g1106(.A(n1815), .B(n1810), .Y(n1816));
AOI21X1  g1107(.A0(n1815), .A1(n1810), .B0(n828), .Y(n1817));
OAI21X1  g1108(.A0(n1817), .A1(n1816), .B0(n801_1), .Y(n1818));
NOR2X1   g1109(.A(g658), .B(n496), .Y(n1819));
NAND3X1  g1110(.A(n1468), .B(n1426), .C(n865), .Y(n1820));
AOI21X1  g1111(.A0(n1820), .A1(g658), .B0(n1819), .Y(n1821));
NOR2X1   g1112(.A(n956_1), .B(n953), .Y(n1822));
NAND4X1  g1113(.A(n763), .B(n789), .C(n792), .D(n940), .Y(n1823));
NAND3X1  g1114(.A(n1823), .B(n1271), .C(n768), .Y(n1824));
OR2X1    g1115(.A(n1824), .B(n947), .Y(n1825));
NAND3X1  g1116(.A(n1825), .B(n1824), .C(n1822), .Y(n1826));
AOI21X1  g1117(.A0(n1821), .A1(n1818), .B0(n1826), .Y(n1827));
OAI21X1  g1118(.A0(n1827), .A1(n1078), .B0(n1803), .Y(n1161));
INVX1    g1119(.A(g161), .Y(n1829));
NAND2X1  g1120(.A(g152), .B(g143), .Y(n1830));
MX2X1    g1121(.A(n1830), .B(n1624), .S0(n1143), .Y(n1831));
MX2X1    g1122(.A(n1491), .B(n1831), .S0(n1135), .Y(n1832));
XOR2X1   g1123(.A(n1832), .B(g161), .Y(n1833));
MX2X1    g1124(.A(n1829), .B(n1833), .S0(n1136_1), .Y(n1834));
OAI21X1  g1125(.A0(n1834), .A1(n1156_1), .B0(n1160), .Y(n1166));
MX2X1    g1126(.A(g693), .B(g512), .S0(n1325), .Y(n1171));
MX2X1    g1127(.A(g532), .B(g690), .S0(n1011_1), .Y(n1176));
INVX1    g1128(.A(n1031_1), .Y(n1838));
MX2X1    g1129(.A(n1038), .B(n1838), .S0(n1037), .Y(n1839));
MX2X1    g1130(.A(n1774), .B(n1839), .S0(n1025), .Y(n1840));
XOR2X1   g1131(.A(n1840), .B(g64), .Y(n1841));
MX2X1    g1132(.A(n1030), .B(n1841), .S0(n1026_1), .Y(n1842));
OAI21X1  g1133(.A0(n1842), .A1(n1051_1), .B0(n1055), .Y(n1181));
NAND2X1  g1134(.A(n995), .B(g3), .Y(n1844));
NAND2X1  g1135(.A(n729), .B(g3), .Y(n1845));
NAND2X1  g1136(.A(n1845), .B(n1844), .Y(n1196));
OR2X1    g1137(.A(n1650), .B(g54), .Y(n1847));
MX2X1    g1138(.A(n1501), .B(n1847), .S0(n1037), .Y(n1848));
MX2X1    g1139(.A(n1702), .B(n1848), .S0(n1025), .Y(n1849));
XOR2X1   g1140(.A(n1849), .B(g59), .Y(n1850));
MX2X1    g1141(.A(n1500), .B(n1850), .S0(n1026_1), .Y(n1851));
OAI21X1  g1142(.A0(n1851), .A1(n1051_1), .B0(n1055), .Y(n1201));
BUFX1    g1143(.A(g705), .Y(g3222));
BUFX1    g1144(.A(g43), .Y(g3600));
BUFX1    g1145(.A(g485), .Y(g4307));
BUFX1    g1146(.A(g668), .Y(g4321));
BUFX1    g1147(.A(g564), .Y(g4422));
BUFX1    g1148(.A(g43), .Y(g5137));
BUFX1    g1149(.A(g485), .Y(g5468));
BUFX1    g1150(.A(g668), .Y(g5469));
BUFX1    g1151(.A(g666), .Y(g1290));
BUFX1    g1152(.A(g45), .Y(g4108));
BUFX1    g1153(.A(g42), .Y(g4106));
BUFX1    g1154(.A(g39), .Y(g4103));
BUFX1    g1155(.A(g699), .Y(g1293));
BUFX1    g1156(.A(g32), .Y(g4099));
BUFX1    g1157(.A(g38), .Y(g4102));
BUFX1    g1158(.A(g46), .Y(g4109));
BUFX1    g1159(.A(g36), .Y(g4100));
BUFX1    g1160(.A(g47), .Y(g4112));
BUFX1    g1161(.A(g40), .Y(g4105));
BUFX1    g1162(.A(g37), .Y(g4101));
BUFX1    g1163(.A(g41), .Y(g4110));
BUFX1    g1164(.A(g22), .Y(g4104));
BUFX1    g1165(.A(g44), .Y(g4107));
BUFX1    g1166(.A(g23), .Y(g4098));
BUFX1    g1167(.A(g2), .Y(n151));
BUFX1    g1168(.A(g18), .Y(n171));
BUFX1    g1169(.A(g571), .Y(n186));
BUFX1    g1170(.A(g39), .Y(n196));
BUFX1    g1171(.A(g654), .Y(n216));
BUFX1    g1172(.A(g18), .Y(n281));
BUFX1    g1173(.A(g646), .Y(n316));
BUFX1    g1174(.A(g28), .Y(n326));
BUFX1    g1175(.A(g650), .Y(n341));
BUFX1    g1176(.A(g14), .Y(n356));
BUFX1    g1177(.A(g634), .Y(n381));
BUFX1    g1178(.A(g32), .Y(n386));
BUFX1    g1179(.A(g28), .Y(n406));
BUFX1    g1180(.A(g567), .Y(n431));
BUFX1    g1181(.A(g10), .Y(n481));
BUFX1    g1182(.A(g664), .Y(n501));
BUFX1    g1183(.A(g598), .Y(n511));
BUFX1    g1184(.A(g567), .Y(n531));
BUFX1    g1185(.A(g663), .Y(n576));
BUFX1    g1186(.A(g40), .Y(n611));
BUFX1    g1187(.A(g1), .Y(n626));
BUFX1    g1188(.A(g37), .Y(n646));
BUFX1    g1189(.A(g42), .Y(n666));
BUFX1    g1190(.A(g24), .Y(n691));
BUFX1    g1191(.A(g24), .Y(n706));
BUFX1    g1192(.A(g654), .Y(n721));
BUFX1    g1193(.A(g650), .Y(n731));
BUFX1    g1194(.A(g642), .Y(n741));
BUFX1    g1195(.A(g6), .Y(n761));
BUFX1    g1196(.A(g38), .Y(n771));
BUFX1    g1197(.A(g10), .Y(n796));
BUFX1    g1198(.A(g45), .Y(n811));
BUFX1    g1199(.A(g36), .Y(n836));
BUFX1    g1200(.A(g606), .Y(n841));
BUFX1    g1201(.A(g667), .Y(n846));
BUFX1    g1202(.A(g42), .Y(n866));
BUFX1    g1203(.A(g702), .Y(n886));
BUFX1    g1204(.A(g665), .Y(n891));
BUFX1    g1205(.A(g634), .Y(n911));
BUFX1    g1206(.A(g598), .Y(n931));
BUFX1    g1207(.A(g646), .Y(n936));
BUFX1    g1208(.A(g642), .Y(n981));
BUFX1    g1209(.A(g606), .Y(n1031));
BUFX1    g1210(.A(g46), .Y(n1051));
BUFX1    g1211(.A(g571), .Y(n1066));
BUFX1    g1212(.A(g1), .Y(n1091));
BUFX1    g1213(.A(g6), .Y(n1151));
BUFX1    g1214(.A(g14), .Y(n1186));
BUFX1    g1215(.A(g2), .Y(n1191));
endmodule
