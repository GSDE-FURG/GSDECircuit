//Converted to Combinational (Partial output: n104) , Module name: s953_n104
module s953_n104 ( Rdy2RtHS1, WantRtHS1, Rdy1RtHS1, WantBmHS1, State_0, Prog_0, FullOHS1, State_3, State_1, State_4, Rdy1BmHS1, Rdy2BmHS1, State_5, Prog_2, State_2, InDoneHS1, FullIHS1, n104 );
input Rdy2RtHS1, WantRtHS1, Rdy1RtHS1, WantBmHS1, State_0, Prog_0, FullOHS1, State_3, State_1, State_4, Rdy1BmHS1, Rdy2BmHS1, State_5, Prog_2, State_2, InDoneHS1, FullIHS1;
output n104;
wire n251, n242, n245, n248, n250, n209, n249, n241, n168, n235, n244, n246, n230, n247, n190, n132, n223, n206, n208, n178, n147, n148, n167, n131, n133_1, n205, n234, n243, n135, n139, n128, n229, n231, n189_1, n188, n136, n129_1, n127, n207, n162, n126, n153_1, n236, n187;
NAND4X1  g126(.A(n248), .B(n245), .C(n242), .D(n251), .Y(n104));
AOI21X1  g125(.A0(n249), .A1(n209), .B0(n250), .Y(n251));
NAND4X1  g116(.A(n168), .B(WantRtHS1), .C(Rdy2RtHS1), .D(n241), .Y(n242));
NAND2X1  g119(.A(n244), .B(n235), .Y(n245));
OAI21X1  g122(.A0(n247), .A1(n230), .B0(n246), .Y(n248));
OAI21X1  g124(.A0(n223), .A1(n132), .B0(n190), .Y(n250));
NOR3X1   g083(.A(n208), .B(n206), .C(n132), .Y(n209));
NOR2X1   g123(.A(n178), .B(Rdy1RtHS1), .Y(n249));
NAND3X1  g115(.A(WantBmHS1), .B(n148), .C(n147), .Y(n241));
NOR4X1   g042(.A(n133_1), .B(State_0), .C(n131), .D(n167), .Y(n168));
MX2X1    g109(.A(n234), .B(n205), .S0(Prog_0), .Y(n235));
NOR2X1   g118(.A(n243), .B(FullOHS1), .Y(n244));
NOR4X1   g120(.A(State_1), .B(State_3), .C(n139), .D(n135), .Y(n246));
OAI21X1  g104(.A0(n229), .A1(State_4), .B0(n128), .Y(n230));
AOI21X1  g121(.A0(Rdy2BmHS1), .A1(Rdy1BmHS1), .B0(n231), .Y(n247));
OAI21X1  g064(.A0(n188), .A1(State_3), .B0(n189_1), .Y(n190));
INVX1    g006(.A(State_1), .Y(n132));
OR4X1    g097(.A(n129_1), .B(n135), .C(State_4), .D(n136), .Y(n223));
NAND4X1  g080(.A(n128), .B(n127), .C(State_5), .D(n135), .Y(n206));
NOR2X1   g082(.A(n207), .B(State_4), .Y(n208));
INVX1    g052(.A(Rdy2RtHS1), .Y(n178));
INVX1    g021(.A(Rdy1BmHS1), .Y(n147));
INVX1    g022(.A(Rdy2BmHS1), .Y(n148));
NAND2X1  g041(.A(n136), .B(n162), .Y(n167));
INVX1    g005(.A(Prog_2), .Y(n131));
NAND4X1  g007(.A(n128), .B(n127), .C(State_5), .D(n132), .Y(n133_1));
NOR2X1   g079(.A(Rdy2RtHS1), .B(n126), .Y(n205));
NOR2X1   g108(.A(Rdy2BmHS1), .B(n147), .Y(n234));
NAND3X1  g117(.A(n236), .B(n153_1), .C(n131), .Y(n243));
INVX1    g009(.A(State_0), .Y(n135));
INVX1    g013(.A(State_5), .Y(n139));
INVX1    g002(.A(State_2), .Y(n128));
MX2X1    g103(.A(InDoneHS1), .B(n136), .S0(Prog_2), .Y(n229));
NOR2X1   g105(.A(State_4), .B(Prog_2), .Y(n231));
NOR4X1   g063(.A(State_2), .B(State_4), .C(State_5), .D(State_1), .Y(n189_1));
NOR4X1   g062(.A(State_0), .B(n148), .C(n147), .D(n187), .Y(n188));
NOR2X1   g010(.A(FullIHS1), .B(FullOHS1), .Y(n136));
NAND3X1  g003(.A(n128), .B(n127), .C(State_5), .Y(n129_1));
INVX1    g001(.A(State_3), .Y(n127));
NOR3X1   g081(.A(n131), .B(FullIHS1), .C(FullOHS1), .Y(n207));
INVX1    g036(.A(State_4), .Y(n162));
INVX1    g000(.A(Rdy1RtHS1), .Y(n126));
NOR4X1   g027(.A(State_2), .B(State_3), .C(n139), .D(State_0), .Y(n153_1));
NOR2X1   g110(.A(State_1), .B(State_4), .Y(n236));
OR2X1    g061(.A(FullIHS1), .B(FullOHS1), .Y(n187));

endmodule
