// Benchmark "i2c" written by ABC on Mon Sep 21 04:03:00 2020

module i2c ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire new_n291_, new_n292_, new_n293_, new_n294_, new_n295_, new_n296_,
    new_n297_, new_n298_, new_n299_, new_n300_, new_n301_, new_n302_,
    new_n303_, new_n304_, new_n305_, new_n306_, new_n307_, new_n308_,
    new_n309_, new_n310_, new_n311_, new_n312_, new_n313_, new_n314_,
    new_n315_, new_n316_, new_n317_, new_n318_, new_n319_, new_n320_,
    new_n321_, new_n322_, new_n323_, new_n324_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n375_, new_n376_, new_n377_,
    new_n378_, new_n379_, new_n380_, new_n381_, new_n382_, new_n383_,
    new_n384_, new_n386_, new_n387_, new_n388_, new_n389_, new_n390_,
    new_n392_, new_n393_, new_n394_, new_n395_, new_n396_, new_n397_,
    new_n398_, new_n399_, new_n400_, new_n401_, new_n402_, new_n404_,
    new_n405_, new_n406_, new_n407_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n426_, new_n427_, new_n428_, new_n429_, new_n431_, new_n432_,
    new_n433_, new_n434_, new_n435_, new_n436_, new_n438_, new_n439_,
    new_n440_, new_n441_, new_n442_, new_n444_, new_n445_, new_n446_,
    new_n447_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n455_, new_n456_, new_n457_, new_n459_, new_n460_, new_n461_,
    new_n462_, new_n463_, new_n464_, new_n465_, new_n466_, new_n467_,
    new_n468_, new_n469_, new_n470_, new_n471_, new_n472_, new_n473_,
    new_n474_, new_n475_, new_n476_, new_n477_, new_n478_, new_n479_,
    new_n481_, new_n482_, new_n483_, new_n485_, new_n486_, new_n487_,
    new_n488_, new_n489_, new_n490_, new_n492_, new_n493_, new_n495_,
    new_n496_, new_n497_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n520_, new_n521_,
    new_n522_, new_n523_, new_n524_, new_n526_, new_n527_, new_n528_,
    new_n529_, new_n531_, new_n532_, new_n534_, new_n535_, new_n536_,
    new_n537_, new_n538_, new_n539_, new_n540_, new_n541_, new_n542_,
    new_n543_, new_n544_, new_n545_, new_n546_, new_n547_, new_n548_,
    new_n549_, new_n550_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n591_, new_n592_, new_n593_,
    new_n594_, new_n595_, new_n596_, new_n598_, new_n599_, new_n600_,
    new_n601_, new_n602_, new_n603_, new_n604_, new_n605_, new_n606_,
    new_n607_, new_n608_, new_n609_, new_n610_, new_n611_, new_n612_,
    new_n613_, new_n614_, new_n615_, new_n616_, new_n617_, new_n619_,
    new_n620_, new_n621_, new_n622_, new_n623_, new_n624_, new_n625_,
    new_n626_, new_n627_, new_n628_, new_n629_, new_n630_, new_n631_,
    new_n632_, new_n633_, new_n634_, new_n635_, new_n637_, new_n638_,
    new_n640_, new_n641_, new_n643_, new_n644_, new_n646_, new_n647_,
    new_n649_, new_n650_, new_n652_, new_n653_, new_n655_, new_n656_,
    new_n658_, new_n659_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n677_,
    new_n678_, new_n679_, new_n680_, new_n681_, new_n682_, new_n684_,
    new_n685_, new_n686_, new_n687_, new_n688_, new_n689_, new_n690_,
    new_n691_, new_n692_, new_n693_, new_n694_, new_n695_, new_n697_,
    new_n698_, new_n699_, new_n700_, new_n701_, new_n702_, new_n703_,
    new_n704_, new_n705_, new_n707_, new_n708_, new_n709_, new_n710_,
    new_n711_, new_n712_, new_n713_, new_n714_, new_n715_, new_n716_,
    new_n717_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n735_, new_n736_, new_n737_,
    new_n738_, new_n739_, new_n740_, new_n741_, new_n742_, new_n743_,
    new_n744_, new_n745_, new_n746_, new_n747_, new_n749_, new_n750_,
    new_n751_, new_n752_, new_n753_, new_n754_, new_n755_, new_n756_,
    new_n757_, new_n758_, new_n759_, new_n761_, new_n762_, new_n763_,
    new_n764_, new_n765_, new_n766_, new_n767_, new_n768_, new_n769_,
    new_n771_, new_n772_, new_n773_, new_n774_, new_n775_, new_n776_,
    new_n777_, new_n778_, new_n779_, new_n780_, new_n781_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n807_, new_n808_, new_n810_,
    new_n811_, new_n813_, new_n814_, new_n815_, new_n816_, new_n817_,
    new_n818_, new_n819_, new_n820_, new_n822_, new_n824_, new_n827_,
    new_n828_, new_n829_, new_n830_, new_n831_, new_n832_, new_n833_,
    new_n834_, new_n835_, new_n836_, new_n837_, new_n838_, new_n839_,
    new_n841_, new_n842_, new_n843_, new_n844_, new_n845_, new_n846_,
    new_n847_, new_n848_, new_n849_, new_n850_, new_n852_, new_n853_,
    new_n854_, new_n856_, new_n857_, new_n858_, new_n859_, new_n860_,
    new_n861_, new_n862_, new_n863_, new_n864_, new_n865_, new_n866_,
    new_n867_, new_n869_, new_n872_, new_n873_, new_n874_, new_n875_,
    new_n876_, new_n877_, new_n879_, new_n880_, new_n882_, new_n883_,
    new_n885_, new_n886_, new_n888_, new_n889_, new_n891_, new_n892_,
    new_n894_, new_n895_, new_n897_, new_n898_, new_n900_, new_n901_,
    new_n903_, new_n904_, new_n906_, new_n908_, new_n910_, new_n912_,
    new_n914_, new_n916_, new_n918_, new_n919_, new_n920_, new_n922_,
    new_n924_, new_n926_, new_n928_, new_n930_, new_n931_, new_n932_,
    new_n933_, new_n934_, new_n935_, new_n936_, new_n937_, new_n939_,
    new_n941_, new_n942_, new_n944_, new_n946_, new_n948_, new_n949_,
    new_n951_, new_n953_, new_n955_, new_n957_, new_n959_, new_n961_,
    new_n962_, new_n963_, new_n965_, new_n966_, new_n967_, new_n968_,
    new_n969_, new_n970_, new_n972_, new_n973_, new_n975_, new_n976_,
    new_n978_, new_n980_, new_n982_, new_n983_, new_n985_, new_n986_,
    new_n987_, new_n988_, new_n989_, new_n990_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1006_, new_n1007_,
    new_n1008_, new_n1009_, new_n1010_, new_n1012_, new_n1013_, new_n1014_,
    new_n1015_, new_n1016_, new_n1017_, new_n1018_, new_n1019_, new_n1021_,
    new_n1023_, new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_,
    new_n1029_, new_n1030_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1040_, new_n1041_, new_n1042_,
    new_n1044_, new_n1046_, new_n1047_, new_n1048_, new_n1049_, new_n1051_,
    new_n1052_, new_n1053_, new_n1055_, new_n1056_, new_n1058_, new_n1059_,
    new_n1060_, new_n1062_, new_n1065_, new_n1066_, new_n1069_, new_n1071_,
    new_n1076_, new_n1078_, new_n1079_;
  INVX1    g000(.A(pi054), .Y(new_n291_));
  OR2X1    g001(.A(pi011), .B(pi009), .Y(new_n292_));
  OR4X1    g002(.A(pi022), .B(pi014), .C(pi013), .D(pi005), .Y(new_n293_));
  OR4X1    g003(.A(pi019), .B(pi018), .C(pi016), .D(pi004), .Y(new_n294_));
  INVX1    g004(.A(pi006), .Y(new_n295_));
  INVX1    g005(.A(pi007), .Y(new_n296_));
  INVX1    g006(.A(pi012), .Y(new_n297_));
  NOR3X1   g007(.A(pi021), .B(pi017), .C(pi008), .Y(new_n298_));
  NAND4X1  g008(.A(new_n298_), .B(new_n297_), .C(new_n296_), .D(new_n295_), .Y(new_n299_));
  NOR4X1   g009(.A(new_n299_), .B(new_n294_), .C(new_n293_), .D(new_n292_), .Y(new_n300_));
  NOR2X1   g010(.A(new_n300_), .B(new_n291_), .Y(new_n301_));
  OR2X1    g011(.A(pi022), .B(pi005), .Y(new_n302_));
  OR2X1    g012(.A(new_n302_), .B(pi056), .Y(new_n303_));
  INVX1    g013(.A(pi056), .Y(new_n304_));
  INVX1    g014(.A(pi014), .Y(new_n305_));
  INVX1    g015(.A(pi013), .Y(new_n306_));
  OR4X1    g016(.A(pi021), .B(new_n306_), .C(pi008), .D(pi007), .Y(new_n307_));
  OR2X1    g017(.A(pi021), .B(pi008), .Y(new_n308_));
  AND2X1   g018(.A(new_n308_), .B(pi007), .Y(new_n309_));
  AOI21X1  g019(.A0(pi021), .A1(pi008), .B0(pi013), .Y(new_n310_));
  OAI21X1  g020(.A0(new_n308_), .A1(pi007), .B0(new_n310_), .Y(new_n311_));
  OAI21X1  g021(.A0(new_n311_), .A1(new_n309_), .B0(new_n307_), .Y(new_n312_));
  NOR4X1   g022(.A(new_n308_), .B(new_n305_), .C(pi013), .D(pi007), .Y(new_n313_));
  AOI21X1  g023(.A0(new_n312_), .A1(new_n305_), .B0(new_n313_), .Y(new_n314_));
  INVX1    g024(.A(pi010), .Y(new_n315_));
  OR2X1    g025(.A(pi014), .B(pi013), .Y(new_n316_));
  OR4X1    g026(.A(new_n308_), .B(new_n316_), .C(new_n315_), .D(pi007), .Y(new_n317_));
  OAI21X1  g027(.A0(new_n314_), .A1(pi010), .B0(new_n317_), .Y(new_n318_));
  OR2X1    g028(.A(pi012), .B(pi006), .Y(new_n319_));
  NOR4X1   g029(.A(new_n319_), .B(new_n294_), .C(new_n302_), .D(pi017), .Y(new_n320_));
  AOI22X1  g030(.A0(new_n320_), .A1(new_n318_), .B0(new_n302_), .B1(new_n304_), .Y(new_n321_));
  MX2X1    g031(.A(new_n321_), .B(new_n303_), .S0(new_n292_), .Y(new_n322_));
  OAI22X1  g032(.A0(new_n322_), .A1(new_n291_), .B0(new_n301_), .B1(pi000), .Y(new_n323_));
  NOR2X1   g033(.A(pi129), .B(pi003), .Y(new_n324_));
  NAND2X1  g034(.A(new_n324_), .B(new_n323_), .Y(po015));
  OR2X1    g035(.A(pi012), .B(pi011), .Y(new_n326_));
  OR2X1    g036(.A(pi022), .B(pi010), .Y(new_n327_));
  OR4X1    g037(.A(new_n327_), .B(new_n326_), .C(new_n308_), .D(pi014), .Y(new_n328_));
  OR2X1    g038(.A(pi013), .B(pi007), .Y(new_n329_));
  OR4X1    g039(.A(new_n329_), .B(new_n294_), .C(pi006), .D(pi005), .Y(new_n330_));
  OR2X1    g040(.A(new_n330_), .B(new_n328_), .Y(new_n331_));
  INVX1    g041(.A(pi017), .Y(new_n332_));
  AND2X1   g042(.A(pi054), .B(new_n332_), .Y(new_n333_));
  AOI21X1  g043(.A0(new_n333_), .A1(new_n331_), .B0(pi001), .Y(new_n334_));
  INVX1    g044(.A(pi009), .Y(new_n335_));
  AND2X1   g045(.A(new_n319_), .B(pi005), .Y(new_n336_));
  NOR3X1   g046(.A(pi012), .B(pi006), .C(pi005), .Y(new_n337_));
  INVX1    g047(.A(new_n337_), .Y(new_n338_));
  AOI21X1  g048(.A0(pi012), .A1(pi006), .B0(pi007), .Y(new_n339_));
  OAI21X1  g049(.A0(new_n319_), .A1(pi005), .B0(new_n339_), .Y(new_n340_));
  OAI22X1  g050(.A0(new_n340_), .A1(new_n336_), .B0(new_n338_), .B1(new_n296_), .Y(new_n341_));
  NOR4X1   g051(.A(new_n319_), .B(new_n306_), .C(pi007), .D(pi005), .Y(new_n342_));
  AOI21X1  g052(.A0(new_n341_), .A1(new_n306_), .B0(new_n342_), .Y(new_n343_));
  NAND3X1  g053(.A(new_n337_), .B(new_n306_), .C(new_n296_), .Y(new_n344_));
  MX2X1    g054(.A(new_n344_), .B(new_n343_), .S0(new_n335_), .Y(new_n345_));
  NOR4X1   g055(.A(pi021), .B(pi017), .C(pi011), .D(pi008), .Y(new_n346_));
  INVX1    g056(.A(new_n346_), .Y(new_n347_));
  OR4X1    g057(.A(new_n291_), .B(pi022), .C(pi014), .D(pi010), .Y(new_n348_));
  NOR4X1   g058(.A(new_n348_), .B(new_n347_), .C(new_n345_), .D(new_n294_), .Y(new_n349_));
  OAI21X1  g059(.A0(new_n349_), .A1(new_n334_), .B0(new_n324_), .Y(po016));
  INVX1    g060(.A(pi065), .Y(new_n351_));
  OR2X1    g061(.A(pi047), .B(pi043), .Y(new_n352_));
  OR4X1    g062(.A(new_n352_), .B(pi048), .C(pi045), .D(pi002), .Y(new_n353_));
  OR2X1    g063(.A(pi044), .B(pi042), .Y(new_n354_));
  OR4X1    g064(.A(pi049), .B(pi024), .C(pi020), .D(pi015), .Y(new_n355_));
  OR4X1    g065(.A(pi050), .B(pi046), .C(pi041), .D(pi038), .Y(new_n356_));
  OR4X1    g066(.A(new_n356_), .B(new_n355_), .C(new_n354_), .D(pi040), .Y(new_n357_));
  OAI21X1  g067(.A0(new_n357_), .A1(new_n353_), .B0(pi082), .Y(new_n358_));
  AND2X1   g068(.A(pi127), .B(pi122), .Y(new_n359_));
  INVX1    g069(.A(new_n359_), .Y(new_n360_));
  NAND3X1  g070(.A(new_n360_), .B(new_n358_), .C(new_n351_), .Y(new_n361_));
  INVX1    g071(.A(pi082), .Y(new_n362_));
  INVX1    g072(.A(pi043), .Y(new_n363_));
  OR4X1    g073(.A(pi044), .B(pi042), .C(pi040), .D(pi038), .Y(new_n364_));
  NOR4X1   g074(.A(new_n364_), .B(pi050), .C(pi046), .D(pi041), .Y(new_n365_));
  AND2X1   g075(.A(new_n365_), .B(new_n363_), .Y(new_n366_));
  OR2X1    g076(.A(pi020), .B(pi015), .Y(new_n367_));
  OR2X1    g077(.A(pi045), .B(pi024), .Y(new_n368_));
  OR2X1    g078(.A(pi048), .B(pi047), .Y(new_n369_));
  NOR4X1   g079(.A(new_n369_), .B(new_n368_), .C(new_n367_), .D(pi049), .Y(new_n370_));
  AOI21X1  g080(.A0(new_n370_), .A1(new_n366_), .B0(new_n362_), .Y(new_n371_));
  AND2X1   g081(.A(new_n359_), .B(new_n362_), .Y(new_n372_));
  OAI21X1  g082(.A0(new_n372_), .A1(new_n371_), .B0(pi002), .Y(new_n373_));
  AOI21X1  g083(.A0(new_n373_), .A1(new_n361_), .B0(pi129), .Y(po017));
  NOR4X1   g084(.A(pi022), .B(pi014), .C(pi010), .D(pi009), .Y(new_n375_));
  INVX1    g085(.A(new_n375_), .Y(new_n376_));
  OR4X1    g086(.A(new_n376_), .B(new_n329_), .C(pi006), .D(pi005), .Y(new_n377_));
  OR2X1    g087(.A(pi017), .B(pi008), .Y(new_n378_));
  OR4X1    g088(.A(new_n378_), .B(new_n326_), .C(new_n294_), .D(pi021), .Y(new_n379_));
  NOR2X1   g089(.A(pi118), .B(pi061), .Y(new_n380_));
  OAI21X1  g090(.A0(new_n379_), .A1(new_n377_), .B0(new_n380_), .Y(new_n381_));
  INVX1    g091(.A(pi113), .Y(new_n382_));
  INVX1    g092(.A(pi123), .Y(new_n383_));
  NAND3X1  g093(.A(new_n383_), .B(new_n382_), .C(pi000), .Y(new_n384_));
  AOI21X1  g094(.A0(new_n384_), .A1(new_n381_), .B0(pi129), .Y(po018));
  INVX1    g095(.A(new_n324_), .Y(new_n386_));
  OR2X1    g096(.A(new_n294_), .B(new_n291_), .Y(new_n387_));
  OR4X1    g097(.A(pi022), .B(pi014), .C(new_n315_), .D(pi009), .Y(new_n388_));
  OR4X1    g098(.A(new_n388_), .B(new_n387_), .C(new_n347_), .D(new_n344_), .Y(new_n389_));
  NAND2X1  g099(.A(new_n291_), .B(pi004), .Y(new_n390_));
  AOI21X1  g100(.A0(new_n390_), .A1(new_n389_), .B0(new_n386_), .Y(po019));
  INVX1    g101(.A(pi005), .Y(new_n392_));
  OR2X1    g102(.A(pi054), .B(new_n392_), .Y(new_n393_));
  OR2X1    g103(.A(new_n291_), .B(pi016), .Y(new_n394_));
  OR4X1    g104(.A(pi012), .B(pi007), .C(pi006), .D(pi005), .Y(new_n395_));
  INVX1    g105(.A(pi025), .Y(new_n396_));
  INVX1    g106(.A(pi029), .Y(new_n397_));
  NOR3X1   g107(.A(pi019), .B(pi018), .C(pi004), .Y(new_n398_));
  NAND4X1  g108(.A(new_n398_), .B(new_n397_), .C(pi028), .D(new_n396_), .Y(new_n399_));
  INVX1    g109(.A(pi059), .Y(new_n400_));
  NAND4X1  g110(.A(new_n375_), .B(new_n346_), .C(new_n400_), .D(new_n306_), .Y(new_n401_));
  OR4X1    g111(.A(new_n401_), .B(new_n399_), .C(new_n395_), .D(new_n394_), .Y(new_n402_));
  AOI21X1  g112(.A0(new_n402_), .A1(new_n393_), .B0(new_n386_), .Y(po020));
  OR2X1    g113(.A(pi054), .B(new_n295_), .Y(new_n404_));
  INVX1    g114(.A(pi028), .Y(new_n405_));
  NAND4X1  g115(.A(new_n398_), .B(new_n397_), .C(new_n405_), .D(pi025), .Y(new_n406_));
  OR4X1    g116(.A(new_n406_), .B(new_n401_), .C(new_n395_), .D(new_n394_), .Y(new_n407_));
  AOI21X1  g117(.A0(new_n407_), .A1(new_n404_), .B0(new_n386_), .Y(po021));
  OR2X1    g118(.A(pi054), .B(new_n296_), .Y(new_n409_));
  NAND2X1  g119(.A(new_n375_), .B(new_n306_), .Y(new_n410_));
  OR2X1    g120(.A(pi021), .B(pi018), .Y(new_n411_));
  OR4X1    g121(.A(new_n291_), .B(pi019), .C(pi016), .D(pi004), .Y(new_n412_));
  NOR2X1   g122(.A(pi007), .B(pi005), .Y(new_n413_));
  NOR3X1   g123(.A(pi012), .B(pi011), .C(pi006), .Y(new_n414_));
  NAND4X1  g124(.A(new_n414_), .B(new_n413_), .C(new_n332_), .D(pi008), .Y(new_n415_));
  OR4X1    g125(.A(new_n415_), .B(new_n412_), .C(new_n411_), .D(new_n410_), .Y(new_n416_));
  AOI21X1  g126(.A0(new_n416_), .A1(new_n409_), .B0(new_n386_), .Y(po022));
  INVX1    g127(.A(pi008), .Y(new_n418_));
  OR2X1    g128(.A(pi054), .B(new_n418_), .Y(new_n419_));
  NAND4X1  g129(.A(new_n375_), .B(new_n337_), .C(new_n306_), .D(new_n296_), .Y(new_n420_));
  INVX1    g130(.A(pi011), .Y(new_n421_));
  NAND3X1  g131(.A(pi021), .B(new_n421_), .C(new_n418_), .Y(new_n422_));
  OR2X1    g132(.A(pi018), .B(pi017), .Y(new_n423_));
  OR4X1    g133(.A(new_n423_), .B(new_n422_), .C(new_n420_), .D(new_n412_), .Y(new_n424_));
  AOI21X1  g134(.A0(new_n424_), .A1(new_n419_), .B0(new_n386_), .Y(po023));
  OR2X1    g135(.A(pi054), .B(new_n335_), .Y(new_n426_));
  OR4X1    g136(.A(pi021), .B(pi018), .C(pi017), .D(pi008), .Y(new_n427_));
  OR4X1    g137(.A(new_n395_), .B(new_n316_), .C(new_n421_), .D(pi009), .Y(new_n428_));
  OR4X1    g138(.A(new_n428_), .B(new_n427_), .C(new_n412_), .D(new_n327_), .Y(new_n429_));
  AOI21X1  g139(.A0(new_n429_), .A1(new_n426_), .B0(new_n386_), .Y(po024));
  OR2X1    g140(.A(pi054), .B(new_n315_), .Y(new_n431_));
  OR2X1    g141(.A(pi019), .B(pi004), .Y(new_n432_));
  NAND2X1  g142(.A(new_n414_), .B(new_n413_), .Y(new_n433_));
  OR4X1    g143(.A(new_n291_), .B(pi016), .C(new_n305_), .D(pi013), .Y(new_n434_));
  OR4X1    g144(.A(new_n427_), .B(pi022), .C(pi010), .D(pi009), .Y(new_n435_));
  OR4X1    g145(.A(new_n435_), .B(new_n434_), .C(new_n433_), .D(new_n432_), .Y(new_n436_));
  AOI21X1  g146(.A0(new_n436_), .A1(new_n431_), .B0(new_n386_), .Y(po025));
  OR2X1    g147(.A(pi054), .B(new_n421_), .Y(new_n438_));
  OR4X1    g148(.A(new_n291_), .B(pi016), .C(pi014), .D(pi009), .Y(new_n439_));
  INVX1    g149(.A(pi022), .Y(new_n440_));
  OR4X1    g150(.A(new_n427_), .B(new_n440_), .C(pi011), .D(pi010), .Y(new_n441_));
  OR4X1    g151(.A(new_n441_), .B(new_n439_), .C(new_n432_), .D(new_n344_), .Y(new_n442_));
  AOI21X1  g152(.A0(new_n442_), .A1(new_n438_), .B0(new_n386_), .Y(po026));
  INVX1    g153(.A(pi018), .Y(new_n444_));
  INVX1    g154(.A(new_n298_), .Y(new_n445_));
  OR4X1    g155(.A(new_n412_), .B(new_n326_), .C(new_n445_), .D(new_n444_), .Y(new_n446_));
  OAI22X1  g156(.A0(new_n446_), .A1(new_n377_), .B0(pi054), .B1(new_n297_), .Y(new_n447_));
  AND2X1   g157(.A(new_n447_), .B(new_n324_), .Y(po027));
  OR2X1    g158(.A(pi054), .B(new_n306_), .Y(new_n449_));
  NOR3X1   g159(.A(new_n397_), .B(pi028), .C(pi025), .Y(new_n450_));
  NAND3X1  g160(.A(new_n450_), .B(new_n398_), .C(new_n375_), .Y(new_n451_));
  OR4X1    g161(.A(new_n394_), .B(new_n338_), .C(pi013), .D(pi007), .Y(new_n452_));
  OR4X1    g162(.A(new_n452_), .B(new_n451_), .C(new_n347_), .D(pi059), .Y(new_n453_));
  AOI21X1  g163(.A0(new_n453_), .A1(new_n449_), .B0(new_n386_), .Y(po028));
  OR2X1    g164(.A(pi054), .B(new_n305_), .Y(new_n455_));
  OR4X1    g165(.A(new_n427_), .B(pi016), .C(new_n306_), .D(pi009), .Y(new_n456_));
  OR4X1    g166(.A(new_n456_), .B(new_n433_), .C(new_n432_), .D(new_n348_), .Y(new_n457_));
  AOI21X1  g167(.A0(new_n457_), .A1(new_n455_), .B0(new_n386_), .Y(po029));
  INVX1    g168(.A(pi129), .Y(new_n459_));
  INVX1    g169(.A(pi015), .Y(new_n460_));
  NOR3X1   g170(.A(pi049), .B(pi045), .C(pi024), .Y(new_n461_));
  NOR3X1   g171(.A(pi048), .B(pi047), .C(pi043), .Y(new_n462_));
  AND2X1   g172(.A(new_n462_), .B(new_n461_), .Y(new_n463_));
  AOI21X1  g173(.A0(new_n463_), .A1(new_n365_), .B0(new_n460_), .Y(new_n464_));
  NOR3X1   g174(.A(pi049), .B(pi024), .C(pi015), .Y(new_n465_));
  OAI21X1  g175(.A0(pi020), .A1(pi002), .B0(new_n465_), .Y(new_n466_));
  NOR3X1   g176(.A(new_n466_), .B(new_n369_), .C(pi045), .Y(new_n467_));
  AOI21X1  g177(.A0(new_n467_), .A1(new_n366_), .B0(new_n464_), .Y(new_n468_));
  INVX1    g178(.A(pi046), .Y(new_n469_));
  NOR3X1   g179(.A(pi044), .B(pi042), .C(pi040), .Y(new_n470_));
  NOR2X1   g180(.A(pi050), .B(pi038), .Y(new_n471_));
  NAND3X1  g181(.A(new_n471_), .B(new_n470_), .C(new_n469_), .Y(new_n472_));
  NOR2X1   g182(.A(pi043), .B(pi041), .Y(new_n473_));
  NOR3X1   g183(.A(pi048), .B(pi047), .C(pi015), .Y(new_n474_));
  NAND3X1  g184(.A(new_n474_), .B(new_n473_), .C(new_n461_), .Y(new_n475_));
  OAI21X1  g185(.A0(new_n475_), .A1(new_n472_), .B0(pi082), .Y(new_n476_));
  AOI21X1  g186(.A0(pi127), .A1(pi122), .B0(pi070), .Y(new_n477_));
  AOI22X1  g187(.A0(new_n477_), .A1(new_n476_), .B0(new_n372_), .B1(pi015), .Y(new_n478_));
  OAI21X1  g188(.A0(new_n468_), .A1(new_n362_), .B0(new_n478_), .Y(new_n479_));
  AND2X1   g189(.A(new_n479_), .B(new_n459_), .Y(po030));
  NAND2X1  g190(.A(new_n291_), .B(pi016), .Y(new_n481_));
  OR4X1    g191(.A(new_n329_), .B(pi012), .C(new_n295_), .D(pi005), .Y(new_n482_));
  OR4X1    g192(.A(new_n482_), .B(new_n387_), .C(new_n376_), .D(new_n347_), .Y(new_n483_));
  AOI21X1  g193(.A0(new_n483_), .A1(new_n481_), .B0(new_n386_), .Y(po031));
  OR2X1    g194(.A(pi054), .B(new_n332_), .Y(new_n485_));
  OR2X1    g195(.A(new_n308_), .B(pi011), .Y(new_n486_));
  NAND4X1  g196(.A(new_n398_), .B(pi059), .C(new_n397_), .D(new_n405_), .Y(new_n487_));
  NOR4X1   g197(.A(pi025), .B(pi016), .C(pi012), .D(pi007), .Y(new_n488_));
  NAND4X1  g198(.A(new_n488_), .B(new_n333_), .C(new_n295_), .D(new_n392_), .Y(new_n489_));
  OR4X1    g199(.A(new_n489_), .B(new_n487_), .C(new_n486_), .D(new_n410_), .Y(new_n490_));
  AOI21X1  g200(.A0(new_n490_), .A1(new_n485_), .B0(new_n386_), .Y(po032));
  NAND4X1  g201(.A(new_n398_), .B(new_n346_), .C(pi054), .D(pi016), .Y(new_n492_));
  OAI22X1  g202(.A0(new_n492_), .A1(new_n420_), .B0(pi054), .B1(new_n444_), .Y(new_n493_));
  AND2X1   g203(.A(new_n493_), .B(new_n324_), .Y(po033));
  NAND2X1  g204(.A(new_n291_), .B(pi019), .Y(new_n495_));
  OR4X1    g205(.A(pi019), .B(pi018), .C(new_n332_), .D(pi004), .Y(new_n496_));
  OR4X1    g206(.A(new_n496_), .B(new_n486_), .C(new_n420_), .D(new_n394_), .Y(new_n497_));
  AOI21X1  g207(.A0(new_n497_), .A1(new_n495_), .B0(new_n386_), .Y(po034));
  INVX1    g208(.A(pi020), .Y(new_n499_));
  OR2X1    g209(.A(pi048), .B(pi045), .Y(new_n500_));
  OR4X1    g210(.A(pi047), .B(pi046), .C(pi043), .D(pi041), .Y(new_n501_));
  NOR3X1   g211(.A(new_n501_), .B(new_n500_), .C(pi024), .Y(new_n502_));
  INVX1    g212(.A(pi038), .Y(new_n503_));
  INVX1    g213(.A(pi040), .Y(new_n504_));
  INVX1    g214(.A(pi050), .Y(new_n505_));
  NAND3X1  g215(.A(new_n505_), .B(new_n504_), .C(new_n503_), .Y(new_n506_));
  NOR4X1   g216(.A(new_n506_), .B(new_n354_), .C(pi049), .D(pi015), .Y(new_n507_));
  AOI21X1  g217(.A0(new_n507_), .A1(new_n502_), .B0(new_n499_), .Y(new_n508_));
  INVX1    g218(.A(pi002), .Y(new_n509_));
  INVX1    g219(.A(pi044), .Y(new_n510_));
  NOR3X1   g220(.A(pi049), .B(pi020), .C(pi015), .Y(new_n511_));
  NOR4X1   g221(.A(pi050), .B(pi042), .C(pi040), .D(pi038), .Y(new_n512_));
  NAND4X1  g222(.A(new_n512_), .B(new_n502_), .C(new_n511_), .D(new_n510_), .Y(new_n513_));
  NOR2X1   g223(.A(new_n513_), .B(new_n509_), .Y(new_n514_));
  OAI21X1  g224(.A0(new_n514_), .A1(new_n508_), .B0(pi082), .Y(new_n515_));
  OR2X1    g225(.A(new_n359_), .B(pi071), .Y(new_n516_));
  AOI21X1  g226(.A0(new_n513_), .A1(pi082), .B0(new_n516_), .Y(new_n517_));
  AOI21X1  g227(.A0(new_n372_), .A1(pi020), .B0(new_n517_), .Y(new_n518_));
  AOI21X1  g228(.A0(new_n518_), .A1(new_n515_), .B0(pi129), .Y(po035));
  INVX1    g229(.A(pi021), .Y(new_n520_));
  OR2X1    g230(.A(pi054), .B(new_n520_), .Y(new_n521_));
  NAND3X1  g231(.A(pi054), .B(new_n520_), .C(pi019), .Y(new_n522_));
  OR4X1    g232(.A(pi016), .B(pi011), .C(pi008), .D(pi004), .Y(new_n523_));
  OR4X1    g233(.A(new_n523_), .B(new_n522_), .C(new_n423_), .D(new_n420_), .Y(new_n524_));
  AOI21X1  g234(.A0(new_n524_), .A1(new_n521_), .B0(new_n386_), .Y(po036));
  OR2X1    g235(.A(pi054), .B(new_n440_), .Y(new_n526_));
  INVX1    g236(.A(new_n414_), .Y(new_n527_));
  OR4X1    g237(.A(pi014), .B(pi013), .C(pi007), .D(new_n392_), .Y(new_n528_));
  OR4X1    g238(.A(new_n528_), .B(new_n435_), .C(new_n527_), .D(new_n412_), .Y(new_n529_));
  AOI21X1  g239(.A0(new_n529_), .A1(new_n526_), .B0(new_n386_), .Y(po037));
  INVX1    g240(.A(pi023), .Y(new_n531_));
  NAND2X1  g241(.A(new_n459_), .B(pi061), .Y(new_n532_));
  AOI21X1  g242(.A0(pi055), .A1(new_n531_), .B0(new_n532_), .Y(po038));
  INVX1    g243(.A(pi063), .Y(new_n534_));
  OR2X1    g244(.A(pi045), .B(pi002), .Y(new_n535_));
  NOR4X1   g245(.A(new_n535_), .B(new_n369_), .C(new_n367_), .D(pi049), .Y(new_n536_));
  AOI21X1  g246(.A0(new_n536_), .A1(new_n366_), .B0(new_n362_), .Y(new_n537_));
  NOR3X1   g247(.A(new_n537_), .B(new_n359_), .C(new_n534_), .Y(new_n538_));
  OR4X1    g248(.A(new_n500_), .B(pi047), .C(pi043), .D(pi041), .Y(new_n539_));
  OAI21X1  g249(.A0(new_n539_), .A1(new_n472_), .B0(pi082), .Y(new_n540_));
  OR4X1    g250(.A(pi049), .B(pi020), .C(pi015), .D(pi002), .Y(new_n541_));
  AND2X1   g251(.A(new_n541_), .B(pi082), .Y(new_n542_));
  OR2X1    g252(.A(new_n542_), .B(new_n360_), .Y(new_n543_));
  AOI21X1  g253(.A0(new_n543_), .A1(new_n540_), .B0(pi024), .Y(new_n544_));
  INVX1    g254(.A(pi041), .Y(new_n545_));
  NAND3X1  g255(.A(new_n469_), .B(new_n363_), .C(new_n545_), .Y(new_n546_));
  OR4X1    g256(.A(new_n546_), .B(pi048), .C(pi047), .D(pi045), .Y(new_n547_));
  INVX1    g257(.A(pi042), .Y(new_n548_));
  NAND4X1  g258(.A(pi082), .B(new_n510_), .C(new_n548_), .D(pi024), .Y(new_n549_));
  NOR3X1   g259(.A(new_n549_), .B(new_n547_), .C(new_n506_), .Y(new_n550_));
  NOR4X1   g260(.A(new_n550_), .B(new_n544_), .C(new_n538_), .D(pi129), .Y(po039));
  INVX1    g261(.A(pi026), .Y(new_n552_));
  INVX1    g262(.A(pi116), .Y(new_n553_));
  NAND3X1  g263(.A(new_n553_), .B(new_n552_), .C(pi025), .Y(new_n554_));
  INVX1    g264(.A(pi053), .Y(new_n555_));
  INVX1    g265(.A(pi085), .Y(new_n556_));
  INVX1    g266(.A(pi100), .Y(new_n557_));
  NOR3X1   g267(.A(pi110), .B(pi096), .C(pi085), .Y(new_n558_));
  AOI21X1  g268(.A0(pi116), .A1(pi085), .B0(new_n558_), .Y(new_n559_));
  OR2X1    g269(.A(pi116), .B(new_n396_), .Y(new_n560_));
  OAI22X1  g270(.A0(new_n560_), .A1(new_n556_), .B0(new_n559_), .B1(new_n557_), .Y(new_n561_));
  NOR3X1   g271(.A(pi052), .B(pi051), .C(pi039), .Y(new_n562_));
  NOR3X1   g272(.A(pi100), .B(pi097), .C(pi095), .Y(new_n563_));
  OR2X1    g273(.A(new_n563_), .B(pi110), .Y(new_n564_));
  AND2X1   g274(.A(pi116), .B(pi026), .Y(new_n565_));
  AOI21X1  g275(.A0(new_n564_), .A1(pi025), .B0(new_n565_), .Y(new_n566_));
  OAI22X1  g276(.A0(new_n566_), .A1(new_n562_), .B0(new_n560_), .B1(new_n552_), .Y(new_n567_));
  AOI22X1  g277(.A0(new_n567_), .A1(new_n556_), .B0(new_n561_), .B1(new_n552_), .Y(new_n568_));
  AND2X1   g278(.A(new_n564_), .B(pi025), .Y(new_n569_));
  NOR3X1   g279(.A(pi052), .B(pi051), .C(pi039), .Y(new_n570_));
  MX2X1    g280(.A(new_n570_), .B(pi025), .S0(new_n553_), .Y(new_n571_));
  AOI22X1  g281(.A0(new_n571_), .A1(pi027), .B0(new_n569_), .B1(new_n562_), .Y(new_n572_));
  OR2X1    g282(.A(pi085), .B(pi026), .Y(new_n573_));
  OAI22X1  g283(.A0(new_n573_), .A1(new_n572_), .B0(new_n568_), .B1(pi027), .Y(new_n574_));
  NOR4X1   g284(.A(new_n554_), .B(pi085), .C(new_n555_), .D(pi027), .Y(new_n575_));
  AOI21X1  g285(.A0(new_n574_), .A1(new_n555_), .B0(new_n575_), .Y(new_n576_));
  INVX1    g286(.A(pi058), .Y(new_n577_));
  OR4X1    g287(.A(pi085), .B(new_n577_), .C(pi053), .D(pi027), .Y(new_n578_));
  OAI22X1  g288(.A0(new_n578_), .A1(new_n554_), .B0(new_n576_), .B1(pi058), .Y(new_n579_));
  AND2X1   g289(.A(new_n579_), .B(new_n324_), .Y(po040));
  NAND2X1  g290(.A(pi116), .B(pi085), .Y(new_n581_));
  INVX1    g291(.A(pi110), .Y(new_n582_));
  OAI21X1  g292(.A0(pi116), .A1(new_n556_), .B0(new_n582_), .Y(new_n583_));
  OR2X1    g293(.A(new_n565_), .B(pi096), .Y(new_n584_));
  OAI22X1  g294(.A0(new_n584_), .A1(new_n583_), .B0(new_n581_), .B1(pi026), .Y(new_n585_));
  AOI21X1  g295(.A0(new_n570_), .A1(pi116), .B0(pi085), .Y(new_n586_));
  AOI22X1  g296(.A0(new_n586_), .A1(pi026), .B0(new_n585_), .B1(pi100), .Y(new_n587_));
  INVX1    g297(.A(pi027), .Y(new_n588_));
  NAND3X1  g298(.A(new_n577_), .B(new_n555_), .C(new_n588_), .Y(new_n589_));
  NOR3X1   g299(.A(new_n589_), .B(new_n587_), .C(new_n386_), .Y(po041));
  INVX1    g300(.A(pi096), .Y(new_n591_));
  NAND2X1  g301(.A(pi116), .B(pi027), .Y(new_n592_));
  NAND3X1  g302(.A(new_n592_), .B(new_n591_), .C(pi095), .Y(new_n593_));
  OAI22X1  g303(.A0(new_n593_), .A1(new_n583_), .B0(new_n581_), .B1(pi027), .Y(new_n594_));
  AOI22X1  g304(.A0(new_n594_), .A1(new_n557_), .B0(new_n586_), .B1(pi027), .Y(new_n595_));
  OR2X1    g305(.A(pi058), .B(pi053), .Y(new_n596_));
  NOR4X1   g306(.A(new_n596_), .B(new_n595_), .C(new_n386_), .D(pi026), .Y(po042));
  INVX1    g307(.A(pi051), .Y(new_n598_));
  NOR2X1   g308(.A(pi052), .B(pi039), .Y(new_n599_));
  NAND2X1  g309(.A(new_n599_), .B(new_n598_), .Y(new_n600_));
  OR2X1    g310(.A(new_n562_), .B(pi026), .Y(new_n601_));
  OAI21X1  g311(.A0(new_n600_), .A1(pi027), .B0(new_n601_), .Y(new_n602_));
  XOR2X1   g312(.A(pi027), .B(pi026), .Y(new_n603_));
  AOI22X1  g313(.A0(new_n603_), .A1(new_n553_), .B0(new_n602_), .B1(new_n564_), .Y(new_n604_));
  NOR2X1   g314(.A(new_n604_), .B(new_n405_), .Y(new_n605_));
  AND2X1   g315(.A(new_n591_), .B(pi095), .Y(new_n606_));
  NOR3X1   g316(.A(pi110), .B(pi100), .C(pi026), .Y(new_n607_));
  AOI22X1  g317(.A0(new_n607_), .A1(new_n606_), .B0(new_n570_), .B1(new_n565_), .Y(new_n608_));
  OAI22X1  g318(.A0(new_n608_), .A1(pi027), .B0(new_n601_), .B1(new_n592_), .Y(new_n609_));
  OAI21X1  g319(.A0(new_n609_), .A1(new_n605_), .B0(new_n556_), .Y(new_n610_));
  MX2X1    g320(.A(pi100), .B(new_n405_), .S0(new_n553_), .Y(new_n611_));
  OR4X1    g321(.A(new_n611_), .B(new_n556_), .C(pi027), .D(pi026), .Y(new_n612_));
  AOI21X1  g322(.A0(new_n612_), .A1(new_n610_), .B0(pi053), .Y(new_n613_));
  NAND3X1  g323(.A(new_n553_), .B(pi028), .C(new_n588_), .Y(new_n614_));
  NOR4X1   g324(.A(new_n614_), .B(pi085), .C(new_n555_), .D(pi026), .Y(new_n615_));
  OAI21X1  g325(.A0(new_n615_), .A1(new_n613_), .B0(new_n577_), .Y(new_n616_));
  OR4X1    g326(.A(new_n614_), .B(new_n573_), .C(new_n577_), .D(pi053), .Y(new_n617_));
  AOI21X1  g327(.A0(new_n617_), .A1(new_n616_), .B0(new_n386_), .Y(po043));
  AND2X1   g328(.A(pi110), .B(pi029), .Y(new_n619_));
  OR2X1    g329(.A(pi100), .B(pi095), .Y(new_n620_));
  NAND3X1  g330(.A(new_n582_), .B(pi097), .C(new_n591_), .Y(new_n621_));
  OR2X1    g331(.A(pi097), .B(new_n397_), .Y(new_n622_));
  AOI21X1  g332(.A0(new_n622_), .A1(new_n621_), .B0(new_n620_), .Y(new_n623_));
  OAI21X1  g333(.A0(new_n623_), .A1(new_n619_), .B0(new_n577_), .Y(new_n624_));
  MX2X1    g334(.A(pi029), .B(pi097), .S0(pi116), .Y(new_n625_));
  NAND2X1  g335(.A(new_n625_), .B(pi058), .Y(new_n626_));
  AOI21X1  g336(.A0(new_n626_), .A1(new_n624_), .B0(pi053), .Y(new_n627_));
  NOR4X1   g337(.A(pi116), .B(pi058), .C(new_n555_), .D(new_n397_), .Y(new_n628_));
  OAI21X1  g338(.A0(new_n628_), .A1(new_n627_), .B0(new_n588_), .Y(new_n629_));
  OR4X1    g339(.A(new_n596_), .B(pi116), .C(new_n397_), .D(new_n588_), .Y(new_n630_));
  AOI21X1  g340(.A0(new_n630_), .A1(new_n629_), .B0(pi085), .Y(new_n631_));
  NOR4X1   g341(.A(new_n589_), .B(pi116), .C(new_n556_), .D(new_n397_), .Y(new_n632_));
  OAI21X1  g342(.A0(new_n632_), .A1(new_n631_), .B0(new_n552_), .Y(new_n633_));
  NOR4X1   g343(.A(new_n596_), .B(pi085), .C(pi027), .D(new_n552_), .Y(new_n634_));
  NAND3X1  g344(.A(new_n634_), .B(new_n553_), .C(pi029), .Y(new_n635_));
  AOI21X1  g345(.A0(new_n635_), .A1(new_n633_), .B0(new_n386_), .Y(po044));
  MX2X1    g346(.A(pi030), .B(pi060), .S0(pi109), .Y(new_n637_));
  MX2X1    g347(.A(new_n637_), .B(pi088), .S0(pi106), .Y(new_n638_));
  AND2X1   g348(.A(new_n638_), .B(new_n459_), .Y(po045));
  MX2X1    g349(.A(pi031), .B(pi030), .S0(pi109), .Y(new_n640_));
  MX2X1    g350(.A(new_n640_), .B(pi089), .S0(pi106), .Y(new_n641_));
  AND2X1   g351(.A(new_n641_), .B(new_n459_), .Y(po046));
  MX2X1    g352(.A(pi032), .B(pi031), .S0(pi109), .Y(new_n643_));
  MX2X1    g353(.A(new_n643_), .B(pi099), .S0(pi106), .Y(new_n644_));
  AND2X1   g354(.A(new_n644_), .B(new_n459_), .Y(po047));
  MX2X1    g355(.A(pi033), .B(pi032), .S0(pi109), .Y(new_n646_));
  MX2X1    g356(.A(new_n646_), .B(pi090), .S0(pi106), .Y(new_n647_));
  AND2X1   g357(.A(new_n647_), .B(new_n459_), .Y(po048));
  MX2X1    g358(.A(pi034), .B(pi033), .S0(pi109), .Y(new_n649_));
  MX2X1    g359(.A(new_n649_), .B(pi091), .S0(pi106), .Y(new_n650_));
  AND2X1   g360(.A(new_n650_), .B(new_n459_), .Y(po049));
  MX2X1    g361(.A(pi035), .B(pi034), .S0(pi109), .Y(new_n652_));
  MX2X1    g362(.A(new_n652_), .B(pi092), .S0(pi106), .Y(new_n653_));
  AND2X1   g363(.A(new_n653_), .B(new_n459_), .Y(po050));
  MX2X1    g364(.A(pi036), .B(pi035), .S0(pi109), .Y(new_n655_));
  MX2X1    g365(.A(new_n655_), .B(pi098), .S0(pi106), .Y(new_n656_));
  AND2X1   g366(.A(new_n656_), .B(new_n459_), .Y(po051));
  MX2X1    g367(.A(pi037), .B(pi036), .S0(pi109), .Y(new_n658_));
  MX2X1    g368(.A(new_n658_), .B(pi093), .S0(pi106), .Y(new_n659_));
  AND2X1   g369(.A(new_n659_), .B(new_n459_), .Y(po052));
  NOR3X1   g370(.A(pi050), .B(pi046), .C(pi041), .Y(new_n661_));
  AND2X1   g371(.A(new_n462_), .B(new_n661_), .Y(new_n662_));
  NOR2X1   g372(.A(new_n535_), .B(new_n355_), .Y(new_n663_));
  AOI21X1  g373(.A0(new_n663_), .A1(new_n662_), .B0(new_n362_), .Y(new_n664_));
  OAI22X1  g374(.A0(new_n664_), .A1(new_n360_), .B0(new_n470_), .B1(new_n362_), .Y(new_n665_));
  INVX1    g375(.A(new_n511_), .Y(new_n666_));
  NOR4X1   g376(.A(new_n368_), .B(new_n666_), .C(pi048), .D(pi002), .Y(new_n667_));
  NOR4X1   g377(.A(new_n501_), .B(new_n354_), .C(pi050), .D(pi040), .Y(new_n668_));
  AOI21X1  g378(.A0(new_n668_), .A1(new_n667_), .B0(new_n362_), .Y(new_n669_));
  INVX1    g379(.A(pi074), .Y(new_n670_));
  OR2X1    g380(.A(new_n359_), .B(new_n670_), .Y(new_n671_));
  OR2X1    g381(.A(pi042), .B(pi040), .Y(new_n672_));
  OR4X1    g382(.A(new_n672_), .B(new_n362_), .C(pi044), .D(new_n503_), .Y(new_n673_));
  AND2X1   g383(.A(new_n673_), .B(new_n459_), .Y(new_n674_));
  OAI21X1  g384(.A0(new_n671_), .A1(new_n669_), .B0(new_n674_), .Y(new_n675_));
  AOI21X1  g385(.A0(new_n665_), .A1(new_n503_), .B0(new_n675_), .Y(po053));
  NOR2X1   g386(.A(pi052), .B(pi051), .Y(new_n677_));
  NAND2X1  g387(.A(new_n677_), .B(pi109), .Y(new_n678_));
  NAND2X1  g388(.A(new_n678_), .B(pi039), .Y(new_n679_));
  INVX1    g389(.A(pi109), .Y(new_n680_));
  NOR4X1   g390(.A(new_n680_), .B(pi052), .C(pi051), .D(pi039), .Y(new_n681_));
  NOR2X1   g391(.A(new_n681_), .B(pi106), .Y(new_n682_));
  AOI21X1  g392(.A0(new_n682_), .A1(new_n679_), .B0(pi129), .Y(po054));
  OAI21X1  g393(.A0(pi044), .A1(pi042), .B0(pi082), .Y(new_n684_));
  INVX1    g394(.A(new_n356_), .Y(new_n685_));
  NOR4X1   g395(.A(new_n535_), .B(new_n355_), .C(new_n352_), .D(pi048), .Y(new_n686_));
  AOI21X1  g396(.A0(new_n686_), .A1(new_n685_), .B0(new_n362_), .Y(new_n687_));
  OAI21X1  g397(.A0(new_n687_), .A1(new_n360_), .B0(new_n684_), .Y(new_n688_));
  NOR4X1   g398(.A(new_n501_), .B(new_n354_), .C(pi050), .D(pi038), .Y(new_n689_));
  AOI21X1  g399(.A0(new_n689_), .A1(new_n667_), .B0(new_n362_), .Y(new_n690_));
  INVX1    g400(.A(pi073), .Y(new_n691_));
  OR2X1    g401(.A(new_n359_), .B(new_n691_), .Y(new_n692_));
  NOR3X1   g402(.A(new_n354_), .B(new_n362_), .C(new_n504_), .Y(new_n693_));
  NOR2X1   g403(.A(new_n693_), .B(pi129), .Y(new_n694_));
  OAI21X1  g404(.A0(new_n692_), .A1(new_n690_), .B0(new_n694_), .Y(new_n695_));
  AOI21X1  g405(.A0(new_n688_), .A1(new_n504_), .B0(new_n695_), .Y(po055));
  NAND2X1  g406(.A(new_n472_), .B(pi082), .Y(new_n697_));
  OAI21X1  g407(.A0(new_n686_), .A1(new_n362_), .B0(new_n359_), .Y(new_n698_));
  AOI21X1  g408(.A0(new_n698_), .A1(new_n697_), .B0(pi041), .Y(new_n699_));
  INVX1    g409(.A(pi076), .Y(new_n700_));
  NOR4X1   g410(.A(new_n364_), .B(new_n352_), .C(pi050), .D(pi046), .Y(new_n701_));
  AOI21X1  g411(.A0(new_n701_), .A1(new_n667_), .B0(new_n362_), .Y(new_n702_));
  NOR3X1   g412(.A(new_n702_), .B(new_n359_), .C(new_n700_), .Y(new_n703_));
  OR4X1    g413(.A(pi050), .B(pi046), .C(pi040), .D(pi038), .Y(new_n704_));
  NOR4X1   g414(.A(new_n704_), .B(new_n354_), .C(new_n362_), .D(new_n545_), .Y(new_n705_));
  NOR4X1   g415(.A(new_n705_), .B(new_n703_), .C(new_n699_), .D(pi129), .Y(po056));
  NOR4X1   g416(.A(new_n704_), .B(pi047), .C(pi043), .D(pi041), .Y(new_n707_));
  AOI21X1  g417(.A0(new_n707_), .A1(new_n667_), .B0(new_n362_), .Y(new_n708_));
  OAI22X1  g418(.A0(new_n708_), .A1(new_n360_), .B0(new_n362_), .B1(new_n510_), .Y(new_n709_));
  AND2X1   g419(.A(new_n709_), .B(new_n548_), .Y(new_n710_));
  INVX1    g420(.A(new_n667_), .Y(new_n711_));
  OR4X1    g421(.A(new_n711_), .B(new_n506_), .C(new_n501_), .D(pi044), .Y(new_n712_));
  INVX1    g422(.A(pi072), .Y(new_n713_));
  OR2X1    g423(.A(new_n359_), .B(new_n713_), .Y(new_n714_));
  AOI21X1  g424(.A0(new_n712_), .A1(pi082), .B0(new_n714_), .Y(new_n715_));
  OR2X1    g425(.A(new_n362_), .B(pi044), .Y(new_n716_));
  OAI21X1  g426(.A0(new_n716_), .A1(new_n548_), .B0(new_n459_), .Y(new_n717_));
  NOR3X1   g427(.A(new_n717_), .B(new_n715_), .C(new_n710_), .Y(po057));
  INVX1    g428(.A(pi047), .Y(new_n719_));
  NAND3X1  g429(.A(new_n667_), .B(new_n365_), .C(new_n719_), .Y(new_n720_));
  INVX1    g430(.A(pi077), .Y(new_n721_));
  OR2X1    g431(.A(new_n359_), .B(new_n721_), .Y(new_n722_));
  AOI21X1  g432(.A0(new_n720_), .A1(pi082), .B0(new_n722_), .Y(new_n723_));
  OR2X1    g433(.A(new_n365_), .B(new_n362_), .Y(new_n724_));
  NOR3X1   g434(.A(new_n535_), .B(new_n369_), .C(new_n355_), .Y(new_n725_));
  OAI21X1  g435(.A0(new_n725_), .A1(new_n362_), .B0(new_n359_), .Y(new_n726_));
  AOI21X1  g436(.A0(new_n726_), .A1(new_n724_), .B0(pi043), .Y(new_n727_));
  NOR4X1   g437(.A(new_n716_), .B(new_n672_), .C(new_n356_), .D(new_n363_), .Y(new_n728_));
  NOR4X1   g438(.A(new_n728_), .B(new_n727_), .C(new_n723_), .D(pi129), .Y(po058));
  OR4X1    g439(.A(new_n672_), .B(new_n501_), .C(pi050), .D(pi038), .Y(new_n730_));
  OAI21X1  g440(.A0(new_n730_), .A1(new_n711_), .B0(pi082), .Y(new_n731_));
  MX2X1    g441(.A(pi067), .B(new_n510_), .S0(new_n359_), .Y(new_n732_));
  OAI21X1  g442(.A0(new_n362_), .A1(new_n510_), .B0(new_n459_), .Y(new_n733_));
  AOI21X1  g443(.A0(new_n732_), .A1(new_n731_), .B0(new_n733_), .Y(po059));
  INVX1    g444(.A(pi068), .Y(new_n735_));
  NOR3X1   g445(.A(new_n369_), .B(new_n355_), .C(pi002), .Y(new_n736_));
  AOI21X1  g446(.A0(new_n736_), .A1(new_n366_), .B0(new_n362_), .Y(new_n737_));
  NOR3X1   g447(.A(new_n737_), .B(new_n359_), .C(new_n735_), .Y(new_n738_));
  NAND2X1  g448(.A(new_n471_), .B(new_n470_), .Y(new_n739_));
  OR4X1    g449(.A(new_n739_), .B(new_n546_), .C(pi048), .D(pi047), .Y(new_n740_));
  OAI21X1  g450(.A0(new_n541_), .A1(pi024), .B0(pi082), .Y(new_n741_));
  AOI22X1  g451(.A0(new_n741_), .A1(new_n359_), .B0(new_n740_), .B1(pi082), .Y(new_n742_));
  NOR2X1   g452(.A(new_n742_), .B(pi045), .Y(new_n743_));
  INVX1    g453(.A(new_n661_), .Y(new_n744_));
  NOR3X1   g454(.A(pi042), .B(pi040), .C(pi038), .Y(new_n745_));
  NAND4X1  g455(.A(new_n745_), .B(pi082), .C(pi045), .D(new_n510_), .Y(new_n746_));
  NOR4X1   g456(.A(new_n746_), .B(new_n744_), .C(new_n352_), .D(pi048), .Y(new_n747_));
  NOR4X1   g457(.A(new_n747_), .B(new_n743_), .C(new_n738_), .D(pi129), .Y(po060));
  AOI21X1  g458(.A0(new_n471_), .A1(new_n470_), .B0(new_n362_), .Y(new_n749_));
  NAND3X1  g459(.A(new_n667_), .B(new_n473_), .C(new_n719_), .Y(new_n750_));
  AOI21X1  g460(.A0(new_n750_), .A1(pi082), .B0(new_n360_), .Y(new_n751_));
  OAI21X1  g461(.A0(new_n751_), .A1(new_n749_), .B0(new_n469_), .Y(new_n752_));
  OR2X1    g462(.A(new_n364_), .B(pi050), .Y(new_n753_));
  OAI21X1  g463(.A0(new_n753_), .A1(new_n750_), .B0(pi082), .Y(new_n754_));
  INVX1    g464(.A(pi075), .Y(new_n755_));
  NOR2X1   g465(.A(new_n359_), .B(new_n755_), .Y(new_n756_));
  NOR4X1   g466(.A(new_n364_), .B(new_n362_), .C(pi050), .D(new_n469_), .Y(new_n757_));
  OR2X1    g467(.A(new_n757_), .B(pi129), .Y(new_n758_));
  AOI21X1  g468(.A0(new_n756_), .A1(new_n754_), .B0(new_n758_), .Y(new_n759_));
  AND2X1   g469(.A(new_n759_), .B(new_n752_), .Y(po061));
  INVX1    g470(.A(pi064), .Y(new_n761_));
  AOI21X1  g471(.A0(new_n667_), .A1(new_n366_), .B0(new_n362_), .Y(new_n762_));
  NOR3X1   g472(.A(new_n762_), .B(new_n359_), .C(new_n761_), .Y(new_n763_));
  OR2X1    g473(.A(new_n366_), .B(new_n362_), .Y(new_n764_));
  OAI21X1  g474(.A0(new_n667_), .A1(new_n362_), .B0(new_n359_), .Y(new_n765_));
  AOI21X1  g475(.A0(new_n765_), .A1(new_n764_), .B0(pi047), .Y(new_n766_));
  NAND2X1  g476(.A(new_n471_), .B(new_n469_), .Y(new_n767_));
  NAND2X1  g477(.A(new_n473_), .B(pi047), .Y(new_n768_));
  NOR4X1   g478(.A(new_n768_), .B(new_n716_), .C(new_n672_), .D(new_n767_), .Y(new_n769_));
  NOR4X1   g479(.A(new_n769_), .B(new_n766_), .C(new_n763_), .D(pi129), .Y(po062));
  NOR3X1   g480(.A(new_n368_), .B(new_n367_), .C(pi049), .Y(new_n771_));
  NAND4X1  g481(.A(new_n771_), .B(new_n366_), .C(new_n719_), .D(new_n509_), .Y(new_n772_));
  INVX1    g482(.A(pi062), .Y(new_n773_));
  OR2X1    g483(.A(new_n359_), .B(new_n773_), .Y(new_n774_));
  AOI21X1  g484(.A0(new_n772_), .A1(pi082), .B0(new_n774_), .Y(new_n775_));
  OAI21X1  g485(.A0(new_n739_), .A1(new_n501_), .B0(pi082), .Y(new_n776_));
  OAI21X1  g486(.A0(new_n663_), .A1(new_n362_), .B0(new_n359_), .Y(new_n777_));
  AOI21X1  g487(.A0(new_n777_), .A1(new_n776_), .B0(pi048), .Y(new_n778_));
  INVX1    g488(.A(pi048), .Y(new_n779_));
  NAND2X1  g489(.A(new_n745_), .B(new_n661_), .Y(new_n780_));
  NOR4X1   g490(.A(new_n780_), .B(new_n716_), .C(new_n352_), .D(new_n779_), .Y(new_n781_));
  NOR4X1   g491(.A(new_n781_), .B(new_n778_), .C(new_n775_), .D(pi129), .Y(po063));
  OR4X1    g492(.A(pi050), .B(pi044), .C(pi040), .D(pi038), .Y(new_n783_));
  OR4X1    g493(.A(new_n783_), .B(new_n547_), .C(pi042), .D(pi024), .Y(new_n784_));
  NOR4X1   g494(.A(new_n364_), .B(pi050), .C(pi049), .D(pi024), .Y(new_n785_));
  NOR3X1   g495(.A(pi020), .B(pi015), .C(pi002), .Y(new_n786_));
  NOR3X1   g496(.A(new_n786_), .B(new_n501_), .C(new_n500_), .Y(new_n787_));
  AOI22X1  g497(.A0(new_n787_), .A1(new_n785_), .B0(new_n784_), .B1(pi049), .Y(new_n788_));
  INVX1    g498(.A(new_n785_), .Y(new_n789_));
  OAI21X1  g499(.A0(new_n789_), .A1(new_n547_), .B0(pi082), .Y(new_n790_));
  AOI21X1  g500(.A0(pi127), .A1(pi122), .B0(pi069), .Y(new_n791_));
  AOI22X1  g501(.A0(new_n791_), .A1(new_n790_), .B0(new_n372_), .B1(pi049), .Y(new_n792_));
  OAI21X1  g502(.A0(new_n788_), .A1(new_n362_), .B0(new_n792_), .Y(new_n793_));
  AND2X1   g503(.A(new_n793_), .B(new_n459_), .Y(po064));
  NAND2X1  g504(.A(new_n364_), .B(pi082), .Y(new_n795_));
  NOR3X1   g505(.A(new_n546_), .B(new_n369_), .C(pi002), .Y(new_n796_));
  AOI21X1  g506(.A0(new_n796_), .A1(new_n771_), .B0(new_n362_), .Y(new_n797_));
  OAI21X1  g507(.A0(new_n797_), .A1(new_n360_), .B0(new_n795_), .Y(new_n798_));
  NOR2X1   g508(.A(new_n501_), .B(new_n364_), .Y(new_n799_));
  AOI21X1  g509(.A0(new_n799_), .A1(new_n667_), .B0(new_n362_), .Y(new_n800_));
  INVX1    g510(.A(pi066), .Y(new_n801_));
  OR2X1    g511(.A(new_n359_), .B(new_n801_), .Y(new_n802_));
  NAND4X1  g512(.A(new_n745_), .B(pi082), .C(pi050), .D(new_n510_), .Y(new_n803_));
  AND2X1   g513(.A(new_n803_), .B(new_n459_), .Y(new_n804_));
  OAI21X1  g514(.A0(new_n802_), .A1(new_n800_), .B0(new_n804_), .Y(new_n805_));
  AOI21X1  g515(.A0(new_n798_), .A1(new_n505_), .B0(new_n805_), .Y(po065));
  OR2X1    g516(.A(pi109), .B(new_n598_), .Y(new_n807_));
  AOI21X1  g517(.A0(pi109), .A1(new_n598_), .B0(pi106), .Y(new_n808_));
  AOI21X1  g518(.A0(new_n808_), .A1(new_n807_), .B0(pi129), .Y(po066));
  OAI21X1  g519(.A0(new_n680_), .A1(pi051), .B0(pi052), .Y(new_n810_));
  AOI21X1  g520(.A0(new_n677_), .A1(pi109), .B0(pi106), .Y(new_n811_));
  AOI21X1  g521(.A0(new_n811_), .A1(new_n810_), .B0(pi129), .Y(po067));
  AND2X1   g522(.A(new_n577_), .B(pi053), .Y(new_n813_));
  INVX1    g523(.A(new_n813_), .Y(new_n814_));
  NOR4X1   g524(.A(new_n620_), .B(pi110), .C(pi096), .D(pi058), .Y(new_n815_));
  AOI21X1  g525(.A0(pi116), .A1(pi058), .B0(new_n815_), .Y(new_n816_));
  INVX1    g526(.A(pi097), .Y(new_n817_));
  OR2X1    g527(.A(new_n817_), .B(pi053), .Y(new_n818_));
  OAI22X1  g528(.A0(new_n818_), .A1(new_n816_), .B0(new_n814_), .B1(pi116), .Y(new_n819_));
  NOR4X1   g529(.A(new_n386_), .B(pi085), .C(pi027), .D(pi026), .Y(new_n820_));
  AND2X1   g530(.A(new_n820_), .B(new_n819_), .Y(po068));
  AOI21X1  g531(.A0(new_n725_), .A1(new_n366_), .B0(new_n362_), .Y(new_n822_));
  OAI21X1  g532(.A0(new_n822_), .A1(new_n359_), .B0(new_n459_), .Y(po069));
  INVX1    g533(.A(pi114), .Y(new_n824_));
  OR2X1    g534(.A(pi129), .B(pi123), .Y(po129));
  NOR3X1   g535(.A(po129), .B(pi122), .C(new_n824_), .Y(po070));
  INVX1    g536(.A(pi094), .Y(new_n827_));
  INVX1    g537(.A(new_n565_), .Y(new_n828_));
  MX2X1    g538(.A(new_n828_), .B(pi026), .S0(pi058), .Y(new_n829_));
  AND2X1   g539(.A(new_n553_), .B(pi058), .Y(new_n830_));
  AOI22X1  g540(.A0(new_n553_), .A1(pi037), .B0(pi058), .B1(new_n552_), .Y(new_n831_));
  OAI22X1  g541(.A0(new_n831_), .A1(new_n830_), .B0(new_n829_), .B1(new_n827_), .Y(new_n832_));
  INVX1    g542(.A(pi037), .Y(new_n833_));
  NOR3X1   g543(.A(pi058), .B(new_n833_), .C(pi026), .Y(new_n834_));
  AOI21X1  g544(.A0(new_n832_), .A1(new_n555_), .B0(new_n834_), .Y(new_n835_));
  OR4X1    g545(.A(pi058), .B(pi053), .C(new_n833_), .D(pi026), .Y(new_n836_));
  OAI21X1  g546(.A0(new_n835_), .A1(pi085), .B0(new_n836_), .Y(new_n837_));
  NOR4X1   g547(.A(new_n596_), .B(pi085), .C(new_n833_), .D(pi026), .Y(new_n838_));
  AOI21X1  g548(.A0(new_n837_), .A1(new_n588_), .B0(new_n838_), .Y(new_n839_));
  NOR2X1   g549(.A(new_n839_), .B(new_n386_), .Y(po071));
  INVX1    g550(.A(pi057), .Y(new_n841_));
  NOR2X1   g551(.A(pi053), .B(pi026), .Y(new_n842_));
  AOI21X1  g552(.A0(pi053), .A1(pi026), .B0(pi085), .Y(new_n843_));
  OAI21X1  g553(.A0(new_n843_), .A1(new_n842_), .B0(new_n577_), .Y(new_n844_));
  OR4X1    g554(.A(pi116), .B(pi085), .C(pi053), .D(pi026), .Y(new_n845_));
  AOI21X1  g555(.A0(new_n845_), .A1(new_n844_), .B0(new_n841_), .Y(new_n846_));
  NAND3X1  g556(.A(pi116), .B(pi060), .C(pi058), .Y(new_n847_));
  NOR4X1   g557(.A(new_n847_), .B(pi085), .C(pi053), .D(pi026), .Y(new_n848_));
  OAI21X1  g558(.A0(new_n848_), .A1(new_n846_), .B0(new_n588_), .Y(new_n849_));
  NAND4X1  g559(.A(new_n842_), .B(new_n556_), .C(new_n577_), .D(pi057), .Y(new_n850_));
  AOI21X1  g560(.A0(new_n850_), .A1(new_n849_), .B0(new_n386_), .Y(po072));
  OR4X1    g561(.A(pi116), .B(new_n577_), .C(pi027), .D(pi026), .Y(new_n852_));
  NAND4X1  g562(.A(new_n603_), .B(new_n570_), .C(pi116), .D(new_n577_), .Y(new_n853_));
  OR4X1    g563(.A(pi129), .B(pi085), .C(pi053), .D(pi003), .Y(new_n854_));
  AOI21X1  g564(.A0(new_n853_), .A1(new_n852_), .B0(new_n854_), .Y(po073));
  INVX1    g565(.A(new_n596_), .Y(new_n856_));
  XOR2X1   g566(.A(pi058), .B(pi053), .Y(new_n857_));
  AOI22X1  g567(.A0(new_n857_), .A1(new_n553_), .B0(new_n856_), .B1(new_n564_), .Y(new_n858_));
  NOR2X1   g568(.A(new_n858_), .B(new_n400_), .Y(new_n859_));
  NOR4X1   g569(.A(new_n596_), .B(new_n563_), .C(pi110), .D(new_n591_), .Y(new_n860_));
  OAI21X1  g570(.A0(new_n860_), .A1(new_n859_), .B0(new_n556_), .Y(new_n861_));
  OR4X1    g571(.A(new_n596_), .B(pi116), .C(new_n556_), .D(new_n400_), .Y(new_n862_));
  AOI21X1  g572(.A0(new_n862_), .A1(new_n861_), .B0(pi027), .Y(new_n863_));
  NAND3X1  g573(.A(new_n553_), .B(pi059), .C(pi027), .Y(new_n864_));
  NOR3X1   g574(.A(new_n864_), .B(new_n596_), .C(pi085), .Y(new_n865_));
  OAI21X1  g575(.A0(new_n865_), .A1(new_n863_), .B0(new_n552_), .Y(new_n866_));
  NAND3X1  g576(.A(new_n634_), .B(new_n553_), .C(pi059), .Y(new_n867_));
  AOI21X1  g577(.A0(new_n867_), .A1(new_n866_), .B0(new_n386_), .Y(po074));
  OR2X1    g578(.A(pi122), .B(pi117), .Y(new_n869_));
  MX2X1    g579(.A(pi123), .B(pi060), .S0(new_n869_), .Y(po075));
  NOR4X1   g580(.A(pi129), .B(new_n383_), .C(pi122), .D(pi114), .Y(po076));
  INVX1    g581(.A(pi136), .Y(new_n872_));
  NAND3X1  g582(.A(pi133), .B(pi132), .C(pi131), .Y(new_n873_));
  OR4X1    g583(.A(new_n873_), .B(pi138), .C(pi137), .D(new_n872_), .Y(new_n874_));
  NOR2X1   g584(.A(new_n873_), .B(pi138), .Y(new_n875_));
  NOR3X1   g585(.A(pi140), .B(pi137), .C(new_n872_), .Y(new_n876_));
  AOI22X1  g586(.A0(new_n876_), .A1(new_n875_), .B0(new_n874_), .B1(pi062), .Y(new_n877_));
  OR2X1    g587(.A(new_n877_), .B(pi129), .Y(po077));
  NOR3X1   g588(.A(pi142), .B(pi137), .C(new_n872_), .Y(new_n879_));
  AOI22X1  g589(.A0(new_n879_), .A1(new_n875_), .B0(new_n874_), .B1(pi063), .Y(new_n880_));
  OR2X1    g590(.A(new_n880_), .B(pi129), .Y(po078));
  NOR3X1   g591(.A(pi139), .B(pi137), .C(new_n872_), .Y(new_n882_));
  AOI22X1  g592(.A0(new_n882_), .A1(new_n875_), .B0(new_n874_), .B1(pi064), .Y(new_n883_));
  OR2X1    g593(.A(new_n883_), .B(pi129), .Y(po079));
  NOR3X1   g594(.A(pi146), .B(pi137), .C(new_n872_), .Y(new_n885_));
  AOI22X1  g595(.A0(new_n885_), .A1(new_n875_), .B0(new_n874_), .B1(pi065), .Y(new_n886_));
  OR2X1    g596(.A(new_n886_), .B(pi129), .Y(po080));
  OR4X1    g597(.A(new_n873_), .B(pi138), .C(pi137), .D(pi136), .Y(new_n888_));
  MX2X1    g598(.A(pi143), .B(new_n801_), .S0(new_n888_), .Y(new_n889_));
  OR2X1    g599(.A(new_n889_), .B(pi129), .Y(po081));
  INVX1    g600(.A(pi067), .Y(new_n891_));
  MX2X1    g601(.A(pi139), .B(new_n891_), .S0(new_n888_), .Y(new_n892_));
  OR2X1    g602(.A(new_n892_), .B(pi129), .Y(po082));
  NOR3X1   g603(.A(pi141), .B(pi137), .C(new_n872_), .Y(new_n894_));
  AOI22X1  g604(.A0(new_n894_), .A1(new_n875_), .B0(new_n874_), .B1(pi068), .Y(new_n895_));
  OR2X1    g605(.A(new_n895_), .B(pi129), .Y(po083));
  NOR3X1   g606(.A(pi143), .B(pi137), .C(new_n872_), .Y(new_n897_));
  AOI22X1  g607(.A0(new_n897_), .A1(new_n875_), .B0(new_n874_), .B1(pi069), .Y(new_n898_));
  OR2X1    g608(.A(new_n898_), .B(pi129), .Y(po084));
  NOR3X1   g609(.A(pi144), .B(pi137), .C(new_n872_), .Y(new_n900_));
  AOI22X1  g610(.A0(new_n900_), .A1(new_n875_), .B0(new_n874_), .B1(pi070), .Y(new_n901_));
  OR2X1    g611(.A(new_n901_), .B(pi129), .Y(po085));
  NOR3X1   g612(.A(pi145), .B(pi137), .C(new_n872_), .Y(new_n903_));
  AOI22X1  g613(.A0(new_n903_), .A1(new_n875_), .B0(new_n874_), .B1(pi071), .Y(new_n904_));
  OR2X1    g614(.A(new_n904_), .B(pi129), .Y(po086));
  MX2X1    g615(.A(pi140), .B(new_n713_), .S0(new_n888_), .Y(new_n906_));
  OR2X1    g616(.A(new_n906_), .B(pi129), .Y(po087));
  MX2X1    g617(.A(pi141), .B(new_n691_), .S0(new_n888_), .Y(new_n908_));
  OR2X1    g618(.A(new_n908_), .B(pi129), .Y(po088));
  MX2X1    g619(.A(pi142), .B(new_n670_), .S0(new_n888_), .Y(new_n910_));
  OR2X1    g620(.A(new_n910_), .B(pi129), .Y(po089));
  MX2X1    g621(.A(pi144), .B(new_n755_), .S0(new_n888_), .Y(new_n912_));
  OR2X1    g622(.A(new_n912_), .B(pi129), .Y(po090));
  MX2X1    g623(.A(pi145), .B(new_n700_), .S0(new_n888_), .Y(new_n914_));
  OR2X1    g624(.A(new_n914_), .B(pi129), .Y(po091));
  MX2X1    g625(.A(pi146), .B(new_n721_), .S0(new_n888_), .Y(new_n916_));
  OR2X1    g626(.A(new_n916_), .B(pi129), .Y(po092));
  INVX1    g627(.A(pi137), .Y(new_n918_));
  OR4X1    g628(.A(new_n873_), .B(pi138), .C(new_n918_), .D(pi136), .Y(new_n919_));
  MX2X1    g629(.A(pi142), .B(pi078), .S0(new_n919_), .Y(new_n920_));
  AND2X1   g630(.A(new_n920_), .B(new_n459_), .Y(po093));
  MX2X1    g631(.A(pi143), .B(pi079), .S0(new_n919_), .Y(new_n922_));
  AND2X1   g632(.A(new_n922_), .B(new_n459_), .Y(po094));
  MX2X1    g633(.A(pi144), .B(pi080), .S0(new_n919_), .Y(new_n924_));
  AND2X1   g634(.A(new_n924_), .B(new_n459_), .Y(po095));
  MX2X1    g635(.A(pi145), .B(pi081), .S0(new_n919_), .Y(new_n926_));
  AND2X1   g636(.A(new_n926_), .B(new_n459_), .Y(po096));
  MX2X1    g637(.A(pi146), .B(pi082), .S0(new_n919_), .Y(new_n928_));
  AND2X1   g638(.A(new_n928_), .B(new_n459_), .Y(po097));
  INVX1    g639(.A(pi138), .Y(new_n930_));
  MX2X1    g640(.A(pi089), .B(new_n773_), .S0(new_n930_), .Y(new_n931_));
  MX2X1    g641(.A(pi119), .B(new_n713_), .S0(new_n930_), .Y(new_n932_));
  MX2X1    g642(.A(new_n932_), .B(new_n931_), .S0(pi136), .Y(new_n933_));
  INVX1    g643(.A(pi087), .Y(new_n934_));
  MX2X1    g644(.A(pi115), .B(new_n934_), .S0(new_n930_), .Y(new_n935_));
  NAND3X1  g645(.A(new_n930_), .B(pi136), .C(pi031), .Y(new_n936_));
  OAI21X1  g646(.A0(new_n935_), .A1(pi136), .B0(new_n936_), .Y(new_n937_));
  MX2X1    g647(.A(new_n937_), .B(new_n933_), .S0(new_n918_), .Y(po098));
  MX2X1    g648(.A(pi141), .B(pi084), .S0(new_n919_), .Y(new_n939_));
  AND2X1   g649(.A(new_n939_), .B(new_n459_), .Y(po099));
  NOR3X1   g650(.A(new_n563_), .B(pi110), .C(pi085), .Y(new_n941_));
  AOI22X1  g651(.A0(new_n941_), .A1(pi096), .B0(new_n553_), .B1(pi085), .Y(new_n942_));
  NOR4X1   g652(.A(new_n942_), .B(new_n589_), .C(new_n386_), .D(pi026), .Y(po100));
  MX2X1    g653(.A(pi139), .B(pi086), .S0(new_n919_), .Y(new_n944_));
  AND2X1   g654(.A(new_n944_), .B(new_n459_), .Y(po101));
  MX2X1    g655(.A(pi140), .B(pi087), .S0(new_n919_), .Y(new_n946_));
  AND2X1   g656(.A(new_n946_), .B(new_n459_), .Y(po102));
  OR4X1    g657(.A(new_n873_), .B(pi138), .C(new_n918_), .D(new_n872_), .Y(new_n948_));
  MX2X1    g658(.A(pi139), .B(pi088), .S0(new_n948_), .Y(new_n949_));
  AND2X1   g659(.A(new_n949_), .B(new_n459_), .Y(po103));
  MX2X1    g660(.A(pi140), .B(pi089), .S0(new_n948_), .Y(new_n951_));
  AND2X1   g661(.A(new_n951_), .B(new_n459_), .Y(po104));
  MX2X1    g662(.A(pi142), .B(pi090), .S0(new_n948_), .Y(new_n953_));
  AND2X1   g663(.A(new_n953_), .B(new_n459_), .Y(po105));
  MX2X1    g664(.A(pi143), .B(pi091), .S0(new_n948_), .Y(new_n955_));
  AND2X1   g665(.A(new_n955_), .B(new_n459_), .Y(po106));
  MX2X1    g666(.A(pi144), .B(pi092), .S0(new_n948_), .Y(new_n957_));
  AND2X1   g667(.A(new_n957_), .B(new_n459_), .Y(po107));
  MX2X1    g668(.A(pi146), .B(pi093), .S0(new_n948_), .Y(new_n959_));
  AND2X1   g669(.A(new_n959_), .B(new_n459_), .Y(po108));
  NAND4X1  g670(.A(pi138), .B(pi133), .C(pi132), .D(pi131), .Y(new_n961_));
  OR4X1    g671(.A(new_n961_), .B(pi137), .C(pi136), .D(new_n362_), .Y(new_n962_));
  MX2X1    g672(.A(pi142), .B(pi094), .S0(new_n962_), .Y(new_n963_));
  AND2X1   g673(.A(new_n963_), .B(new_n459_), .Y(po109));
  INVX1    g674(.A(pi095), .Y(new_n965_));
  INVX1    g675(.A(pi143), .Y(new_n966_));
  OR2X1    g676(.A(pi110), .B(pi003), .Y(new_n967_));
  NOR4X1   g677(.A(new_n930_), .B(pi137), .C(pi136), .D(new_n362_), .Y(new_n968_));
  MX2X1    g678(.A(new_n968_), .B(new_n967_), .S0(new_n873_), .Y(new_n969_));
  OAI22X1  g679(.A0(new_n969_), .A1(new_n965_), .B0(new_n962_), .B1(new_n966_), .Y(new_n970_));
  AND2X1   g680(.A(new_n970_), .B(new_n459_), .Y(po110));
  INVX1    g681(.A(pi146), .Y(new_n972_));
  OAI22X1  g682(.A0(new_n969_), .A1(new_n591_), .B0(new_n962_), .B1(new_n972_), .Y(new_n973_));
  AND2X1   g683(.A(new_n973_), .B(new_n459_), .Y(po111));
  INVX1    g684(.A(pi145), .Y(new_n975_));
  OAI22X1  g685(.A0(new_n969_), .A1(new_n817_), .B0(new_n962_), .B1(new_n975_), .Y(new_n976_));
  AND2X1   g686(.A(new_n976_), .B(new_n459_), .Y(po112));
  MX2X1    g687(.A(pi145), .B(pi098), .S0(new_n948_), .Y(new_n978_));
  AND2X1   g688(.A(new_n978_), .B(new_n459_), .Y(po113));
  MX2X1    g689(.A(pi141), .B(pi099), .S0(new_n948_), .Y(new_n980_));
  AND2X1   g690(.A(new_n980_), .B(new_n459_), .Y(po114));
  INVX1    g691(.A(pi144), .Y(new_n982_));
  OAI22X1  g692(.A0(new_n969_), .A1(new_n557_), .B0(new_n962_), .B1(new_n982_), .Y(new_n983_));
  AND2X1   g693(.A(new_n983_), .B(new_n459_), .Y(po115));
  MX2X1    g694(.A(pi124), .B(new_n721_), .S0(new_n930_), .Y(new_n985_));
  MX2X1    g695(.A(pi093), .B(new_n351_), .S0(new_n930_), .Y(new_n986_));
  MX2X1    g696(.A(new_n986_), .B(new_n985_), .S0(new_n872_), .Y(new_n987_));
  NAND3X1  g697(.A(new_n930_), .B(pi136), .C(pi037), .Y(new_n988_));
  MX2X1    g698(.A(new_n591_), .B(new_n362_), .S0(new_n930_), .Y(new_n989_));
  OAI21X1  g699(.A0(new_n989_), .A1(pi136), .B0(new_n988_), .Y(new_n990_));
  MX2X1    g700(.A(new_n990_), .B(new_n987_), .S0(new_n918_), .Y(po116));
  OR2X1    g701(.A(new_n918_), .B(pi136), .Y(new_n992_));
  NAND3X1  g702(.A(new_n918_), .B(pi136), .C(pi091), .Y(new_n993_));
  OAI21X1  g703(.A0(new_n992_), .A1(new_n965_), .B0(new_n993_), .Y(new_n994_));
  MX2X1    g704(.A(pi079), .B(pi034), .S0(pi136), .Y(new_n995_));
  INVX1    g705(.A(pi069), .Y(new_n996_));
  MX2X1    g706(.A(new_n996_), .B(new_n801_), .S0(new_n872_), .Y(new_n997_));
  MX2X1    g707(.A(new_n997_), .B(new_n995_), .S0(pi137), .Y(new_n998_));
  MX2X1    g708(.A(new_n998_), .B(new_n994_), .S0(pi138), .Y(po117));
  NAND3X1  g709(.A(new_n918_), .B(pi136), .C(pi090), .Y(new_n1000_));
  OAI21X1  g710(.A0(new_n992_), .A1(new_n827_), .B0(new_n1000_), .Y(new_n1001_));
  MX2X1    g711(.A(pi078), .B(pi033), .S0(pi136), .Y(new_n1002_));
  MX2X1    g712(.A(new_n670_), .B(new_n534_), .S0(pi136), .Y(new_n1003_));
  MX2X1    g713(.A(new_n1003_), .B(new_n1002_), .S0(pi137), .Y(new_n1004_));
  MX2X1    g714(.A(new_n1004_), .B(new_n1001_), .S0(pi138), .Y(po118));
  NAND3X1  g715(.A(new_n918_), .B(pi136), .C(pi099), .Y(new_n1006_));
  OAI21X1  g716(.A0(new_n992_), .A1(pi112), .B0(new_n1006_), .Y(new_n1007_));
  MX2X1    g717(.A(new_n691_), .B(new_n735_), .S0(pi136), .Y(new_n1008_));
  MX2X1    g718(.A(pi084), .B(pi032), .S0(pi136), .Y(new_n1009_));
  MX2X1    g719(.A(new_n1009_), .B(new_n1008_), .S0(new_n918_), .Y(new_n1010_));
  MX2X1    g720(.A(new_n1010_), .B(new_n1007_), .S0(pi138), .Y(po119));
  INVX1    g721(.A(pi070), .Y(new_n1012_));
  MX2X1    g722(.A(pi092), .B(new_n1012_), .S0(new_n930_), .Y(new_n1013_));
  MX2X1    g723(.A(pi125), .B(new_n755_), .S0(new_n930_), .Y(new_n1014_));
  MX2X1    g724(.A(new_n1014_), .B(new_n1013_), .S0(pi136), .Y(new_n1015_));
  INVX1    g725(.A(pi080), .Y(new_n1016_));
  MX2X1    g726(.A(new_n557_), .B(new_n1016_), .S0(new_n930_), .Y(new_n1017_));
  NAND3X1  g727(.A(new_n930_), .B(pi136), .C(pi035), .Y(new_n1018_));
  OAI21X1  g728(.A0(new_n1017_), .A1(pi136), .B0(new_n1018_), .Y(new_n1019_));
  MX2X1    g729(.A(new_n1019_), .B(new_n1015_), .S0(new_n918_), .Y(po120));
  NAND4X1  g730(.A(new_n941_), .B(new_n856_), .C(new_n588_), .D(new_n552_), .Y(new_n1021_));
  AOI21X1  g731(.A0(new_n1021_), .A1(new_n581_), .B0(new_n386_), .Y(po121));
  INVX1    g732(.A(pi071), .Y(new_n1023_));
  MX2X1    g733(.A(pi098), .B(new_n1023_), .S0(new_n930_), .Y(new_n1024_));
  MX2X1    g734(.A(new_n700_), .B(pi023), .S0(pi138), .Y(new_n1025_));
  MX2X1    g735(.A(new_n1025_), .B(new_n1024_), .S0(pi136), .Y(new_n1026_));
  NAND3X1  g736(.A(new_n930_), .B(pi136), .C(pi036), .Y(new_n1027_));
  INVX1    g737(.A(pi081), .Y(new_n1028_));
  MX2X1    g738(.A(new_n817_), .B(new_n1028_), .S0(new_n930_), .Y(new_n1029_));
  OAI21X1  g739(.A0(new_n1029_), .A1(pi136), .B0(new_n1027_), .Y(new_n1030_));
  MX2X1    g740(.A(new_n1030_), .B(new_n1026_), .S0(new_n918_), .Y(po122));
  MX2X1    g741(.A(pi088), .B(new_n761_), .S0(new_n930_), .Y(new_n1032_));
  MX2X1    g742(.A(pi120), .B(new_n891_), .S0(new_n930_), .Y(new_n1033_));
  MX2X1    g743(.A(new_n1033_), .B(new_n1032_), .S0(pi136), .Y(new_n1034_));
  AND2X1   g744(.A(pi138), .B(pi111), .Y(new_n1035_));
  AOI21X1  g745(.A0(new_n930_), .A1(pi086), .B0(new_n1035_), .Y(new_n1036_));
  NAND3X1  g746(.A(new_n930_), .B(pi136), .C(pi030), .Y(new_n1037_));
  OAI21X1  g747(.A0(new_n1036_), .A1(pi136), .B0(new_n1037_), .Y(new_n1038_));
  MX2X1    g748(.A(new_n1038_), .B(new_n1034_), .S0(new_n918_), .Y(po123));
  OR2X1    g749(.A(pi027), .B(new_n552_), .Y(new_n1040_));
  NAND3X1  g750(.A(new_n600_), .B(pi027), .C(new_n552_), .Y(new_n1041_));
  NAND2X1  g751(.A(new_n324_), .B(pi116), .Y(new_n1042_));
  AOI21X1  g752(.A0(new_n1041_), .A1(new_n1040_), .B0(new_n1042_), .Y(po124));
  NAND3X1  g753(.A(new_n817_), .B(pi058), .C(new_n555_), .Y(new_n1044_));
  AOI21X1  g754(.A0(new_n1044_), .A1(new_n814_), .B0(new_n1042_), .Y(po125));
  INVX1    g755(.A(new_n968_), .Y(new_n1046_));
  NOR3X1   g756(.A(new_n930_), .B(pi137), .C(new_n362_), .Y(new_n1047_));
  AND2X1   g757(.A(pi139), .B(new_n872_), .Y(new_n1048_));
  AOI22X1  g758(.A0(new_n1048_), .A1(new_n1047_), .B0(new_n1046_), .B1(pi111), .Y(new_n1049_));
  NOR3X1   g759(.A(new_n1049_), .B(new_n873_), .C(pi129), .Y(po126));
  AND2X1   g760(.A(pi141), .B(new_n872_), .Y(new_n1051_));
  NOR2X1   g761(.A(new_n968_), .B(pi112), .Y(new_n1052_));
  AOI21X1  g762(.A0(new_n1051_), .A1(new_n1047_), .B0(new_n1052_), .Y(new_n1053_));
  NOR3X1   g763(.A(new_n1053_), .B(new_n873_), .C(pi129), .Y(po127));
  OR2X1    g764(.A(pi113), .B(pi054), .Y(new_n1055_));
  OAI21X1  g765(.A0(pi022), .A1(pi011), .B0(pi054), .Y(new_n1056_));
  AOI21X1  g766(.A0(new_n1056_), .A1(new_n1055_), .B0(new_n386_), .Y(po128));
  AND2X1   g767(.A(pi140), .B(new_n872_), .Y(new_n1058_));
  NOR2X1   g768(.A(new_n968_), .B(pi115), .Y(new_n1059_));
  AOI21X1  g769(.A0(new_n1058_), .A1(new_n1047_), .B0(new_n1059_), .Y(new_n1060_));
  NOR3X1   g770(.A(new_n1060_), .B(new_n873_), .C(pi129), .Y(po130));
  NOR4X1   g771(.A(pi012), .B(pi009), .C(pi007), .D(pi004), .Y(new_n1062_));
  NOR4X1   g772(.A(new_n1062_), .B(pi129), .C(new_n291_), .D(pi003), .Y(po131));
  NAND2X1  g773(.A(new_n459_), .B(pi122), .Y(po132));
  NAND2X1  g774(.A(pi118), .B(new_n291_), .Y(new_n1065_));
  NAND3X1  g775(.A(new_n450_), .B(new_n400_), .C(pi054), .Y(new_n1066_));
  AOI21X1  g776(.A0(new_n1066_), .A1(new_n1065_), .B0(pi129), .Y(po133));
  AND2X1   g777(.A(new_n620_), .B(new_n459_), .Y(po134));
  NOR3X1   g778(.A(pi120), .B(pi110), .C(pi003), .Y(new_n1069_));
  NOR3X1   g779(.A(new_n1069_), .B(pi129), .C(pi111), .Y(po135));
  AND2X1   g780(.A(pi120), .B(pi081), .Y(new_n1071_));
  AND2X1   g781(.A(new_n1071_), .B(new_n459_), .Y(po136));
  OR2X1    g782(.A(pi134), .B(pi129), .Y(po137));
  OR2X1    g783(.A(pi135), .B(pi129), .Y(po138));
  AND2X1   g784(.A(new_n459_), .B(pi057), .Y(po139));
  AOI21X1  g785(.A0(pi125), .A1(new_n591_), .B0(pi003), .Y(new_n1076_));
  NOR2X1   g786(.A(new_n1076_), .B(pi129), .Y(po140));
  INVX1    g787(.A(pi132), .Y(new_n1078_));
  INVX1    g788(.A(pi133), .Y(new_n1079_));
  NOR3X1   g789(.A(new_n1079_), .B(new_n1078_), .C(pi126), .Y(po141));
  ONE      g790(.Y(po012));
  BUFX1    g791(.A(pi108), .Y(po000));
  BUFX1    g792(.A(pi083), .Y(po001));
  BUFX1    g793(.A(pi104), .Y(po002));
  BUFX1    g794(.A(pi103), .Y(po003));
  BUFX1    g795(.A(pi102), .Y(po004));
  BUFX1    g796(.A(pi105), .Y(po005));
  BUFX1    g797(.A(pi107), .Y(po006));
  BUFX1    g798(.A(pi101), .Y(po007));
  BUFX1    g799(.A(pi126), .Y(po008));
  BUFX1    g800(.A(pi121), .Y(po009));
  BUFX1    g801(.A(pi001), .Y(po010));
  BUFX1    g802(.A(pi000), .Y(po011));
  BUFX1    g803(.A(pi130), .Y(po013));
  BUFX1    g804(.A(pi128), .Y(po014));
endmodule


