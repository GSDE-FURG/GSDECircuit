// Benchmark "top" written by ABC on Mon Sep 21 03:40:29 2020

module top ( 
    \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] ,
    \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] ,
    \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] ,
    \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31]   );
  input  \a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] ,
    \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] ,
    \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] ,
    \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] ;
  wire new_n65_, new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_,
    new_n72_, new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_,
    new_n79_, new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_,
    new_n86_, new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_,
    new_n93_, new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_,
    new_n100_, new_n101_, new_n102_, new_n103_, new_n104_, new_n105_,
    new_n106_, new_n107_, new_n108_, new_n109_, new_n110_, new_n111_,
    new_n112_, new_n113_, new_n114_, new_n115_, new_n116_, new_n117_,
    new_n118_, new_n119_, new_n120_, new_n121_, new_n122_, new_n123_,
    new_n124_, new_n125_, new_n126_, new_n127_, new_n128_, new_n129_,
    new_n130_, new_n131_, new_n132_, new_n133_, new_n134_, new_n135_,
    new_n136_, new_n137_, new_n138_, new_n139_, new_n140_, new_n141_,
    new_n142_, new_n143_, new_n144_, new_n145_, new_n146_, new_n147_,
    new_n148_, new_n149_, new_n150_, new_n151_, new_n152_, new_n153_,
    new_n154_, new_n155_, new_n156_, new_n157_, new_n158_, new_n159_,
    new_n160_, new_n161_, new_n162_, new_n163_, new_n164_, new_n165_,
    new_n166_, new_n167_, new_n168_, new_n169_, new_n170_, new_n171_,
    new_n172_, new_n173_, new_n174_, new_n175_, new_n176_, new_n177_,
    new_n178_, new_n179_, new_n180_, new_n181_, new_n182_, new_n183_,
    new_n184_, new_n185_, new_n186_, new_n187_, new_n188_, new_n189_,
    new_n190_, new_n191_, new_n192_, new_n193_, new_n194_, new_n195_,
    new_n196_, new_n197_, new_n198_, new_n199_, new_n200_, new_n201_,
    new_n202_, new_n203_, new_n204_, new_n205_, new_n206_, new_n207_,
    new_n208_, new_n209_, new_n210_, new_n211_, new_n212_, new_n213_,
    new_n214_, new_n215_, new_n216_, new_n217_, new_n218_, new_n219_,
    new_n220_, new_n221_, new_n222_, new_n223_, new_n224_, new_n225_,
    new_n226_, new_n227_, new_n228_, new_n229_, new_n230_, new_n231_,
    new_n232_, new_n233_, new_n234_, new_n235_, new_n236_, new_n237_,
    new_n238_, new_n239_, new_n240_, new_n241_, new_n242_, new_n243_,
    new_n244_, new_n245_, new_n246_, new_n247_, new_n248_, new_n249_,
    new_n250_, new_n251_, new_n252_, new_n253_, new_n254_, new_n255_,
    new_n256_, new_n257_, new_n258_, new_n259_, new_n260_, new_n261_,
    new_n262_, new_n263_, new_n264_, new_n265_, new_n266_, new_n267_,
    new_n268_, new_n269_, new_n270_, new_n271_, new_n272_, new_n273_,
    new_n274_, new_n275_, new_n276_, new_n277_, new_n278_, new_n279_,
    new_n280_, new_n281_, new_n282_, new_n283_, new_n284_, new_n285_,
    new_n286_, new_n287_, new_n288_, new_n289_, new_n290_, new_n291_,
    new_n292_, new_n293_, new_n294_, new_n295_, new_n296_, new_n297_,
    new_n298_, new_n299_, new_n300_, new_n301_, new_n302_, new_n303_,
    new_n304_, new_n305_, new_n306_, new_n307_, new_n308_, new_n309_,
    new_n310_, new_n311_, new_n312_, new_n313_, new_n314_, new_n315_,
    new_n316_, new_n317_, new_n318_, new_n319_, new_n320_, new_n321_,
    new_n322_, new_n323_, new_n324_, new_n325_, new_n326_, new_n327_,
    new_n328_, new_n329_, new_n330_, new_n331_, new_n332_, new_n333_,
    new_n334_, new_n335_, new_n336_, new_n337_, new_n338_, new_n339_,
    new_n340_, new_n341_, new_n342_, new_n343_, new_n344_, new_n345_,
    new_n346_, new_n347_, new_n348_, new_n349_, new_n350_, new_n351_,
    new_n352_, new_n353_, new_n354_, new_n355_, new_n356_, new_n357_,
    new_n358_, new_n359_, new_n360_, new_n361_, new_n362_, new_n363_,
    new_n364_, new_n365_, new_n366_, new_n367_, new_n368_, new_n369_,
    new_n370_, new_n371_, new_n372_, new_n373_, new_n374_, new_n375_,
    new_n376_, new_n377_, new_n378_, new_n379_, new_n380_, new_n381_,
    new_n382_, new_n383_, new_n384_, new_n385_, new_n386_, new_n387_,
    new_n388_, new_n389_, new_n390_, new_n391_, new_n392_, new_n393_,
    new_n394_, new_n395_, new_n396_, new_n397_, new_n398_, new_n399_,
    new_n400_, new_n401_, new_n402_, new_n403_, new_n404_, new_n405_,
    new_n406_, new_n407_, new_n408_, new_n409_, new_n410_, new_n411_,
    new_n412_, new_n413_, new_n414_, new_n415_, new_n416_, new_n417_,
    new_n418_, new_n419_, new_n420_, new_n421_, new_n422_, new_n423_,
    new_n424_, new_n425_, new_n426_, new_n427_, new_n428_, new_n429_,
    new_n430_, new_n431_, new_n432_, new_n433_, new_n434_, new_n435_,
    new_n436_, new_n437_, new_n438_, new_n439_, new_n440_, new_n441_,
    new_n442_, new_n443_, new_n444_, new_n445_, new_n446_, new_n447_,
    new_n448_, new_n449_, new_n450_, new_n451_, new_n452_, new_n453_,
    new_n454_, new_n455_, new_n456_, new_n457_, new_n458_, new_n459_,
    new_n460_, new_n461_, new_n462_, new_n463_, new_n464_, new_n465_,
    new_n466_, new_n467_, new_n468_, new_n469_, new_n470_, new_n471_,
    new_n472_, new_n473_, new_n474_, new_n475_, new_n476_, new_n477_,
    new_n478_, new_n479_, new_n480_, new_n481_, new_n482_, new_n483_,
    new_n484_, new_n485_, new_n486_, new_n487_, new_n488_, new_n489_,
    new_n490_, new_n491_, new_n492_, new_n493_, new_n494_, new_n495_,
    new_n496_, new_n497_, new_n498_, new_n499_, new_n500_, new_n501_,
    new_n502_, new_n503_, new_n504_, new_n505_, new_n506_, new_n507_,
    new_n508_, new_n509_, new_n510_, new_n511_, new_n512_, new_n513_,
    new_n514_, new_n515_, new_n516_, new_n517_, new_n518_, new_n519_,
    new_n520_, new_n521_, new_n522_, new_n523_, new_n524_, new_n525_,
    new_n526_, new_n527_, new_n528_, new_n529_, new_n530_, new_n531_,
    new_n532_, new_n533_, new_n534_, new_n535_, new_n536_, new_n537_,
    new_n538_, new_n539_, new_n540_, new_n541_, new_n542_, new_n543_,
    new_n544_, new_n545_, new_n546_, new_n547_, new_n548_, new_n549_,
    new_n550_, new_n551_, new_n552_, new_n553_, new_n554_, new_n555_,
    new_n556_, new_n557_, new_n558_, new_n559_, new_n560_, new_n561_,
    new_n562_, new_n563_, new_n564_, new_n565_, new_n566_, new_n567_,
    new_n568_, new_n569_, new_n570_, new_n571_, new_n572_, new_n573_,
    new_n574_, new_n575_, new_n576_, new_n577_, new_n578_, new_n579_,
    new_n580_, new_n581_, new_n582_, new_n583_, new_n584_, new_n585_,
    new_n586_, new_n587_, new_n588_, new_n589_, new_n590_, new_n591_,
    new_n592_, new_n593_, new_n594_, new_n595_, new_n596_, new_n597_,
    new_n598_, new_n599_, new_n600_, new_n601_, new_n602_, new_n603_,
    new_n604_, new_n605_, new_n606_, new_n607_, new_n608_, new_n609_,
    new_n610_, new_n611_, new_n612_, new_n613_, new_n614_, new_n615_,
    new_n616_, new_n617_, new_n618_, new_n619_, new_n620_, new_n621_,
    new_n622_, new_n623_, new_n624_, new_n625_, new_n626_, new_n627_,
    new_n628_, new_n629_, new_n630_, new_n631_, new_n632_, new_n633_,
    new_n634_, new_n635_, new_n636_, new_n637_, new_n638_, new_n639_,
    new_n640_, new_n641_, new_n642_, new_n643_, new_n644_, new_n645_,
    new_n646_, new_n647_, new_n648_, new_n649_, new_n650_, new_n651_,
    new_n652_, new_n653_, new_n654_, new_n655_, new_n656_, new_n657_,
    new_n658_, new_n659_, new_n660_, new_n661_, new_n662_, new_n663_,
    new_n664_, new_n665_, new_n666_, new_n667_, new_n668_, new_n669_,
    new_n670_, new_n671_, new_n672_, new_n673_, new_n674_, new_n675_,
    new_n676_, new_n677_, new_n678_, new_n679_, new_n680_, new_n681_,
    new_n682_, new_n683_, new_n684_, new_n685_, new_n686_, new_n687_,
    new_n688_, new_n689_, new_n690_, new_n691_, new_n692_, new_n693_,
    new_n694_, new_n695_, new_n696_, new_n697_, new_n698_, new_n699_,
    new_n700_, new_n701_, new_n702_, new_n703_, new_n704_, new_n705_,
    new_n706_, new_n707_, new_n708_, new_n709_, new_n710_, new_n711_,
    new_n712_, new_n713_, new_n714_, new_n715_, new_n716_, new_n717_,
    new_n718_, new_n719_, new_n720_, new_n721_, new_n722_, new_n723_,
    new_n724_, new_n725_, new_n726_, new_n727_, new_n728_, new_n729_,
    new_n730_, new_n731_, new_n732_, new_n733_, new_n734_, new_n735_,
    new_n736_, new_n737_, new_n738_, new_n739_, new_n740_, new_n741_,
    new_n742_, new_n743_, new_n744_, new_n745_, new_n746_, new_n747_,
    new_n748_, new_n749_, new_n750_, new_n751_, new_n752_, new_n753_,
    new_n754_, new_n755_, new_n756_, new_n757_, new_n758_, new_n759_,
    new_n760_, new_n761_, new_n762_, new_n763_, new_n764_, new_n765_,
    new_n766_, new_n767_, new_n768_, new_n769_, new_n770_, new_n771_,
    new_n772_, new_n773_, new_n774_, new_n775_, new_n776_, new_n777_,
    new_n778_, new_n779_, new_n780_, new_n781_, new_n782_, new_n783_,
    new_n784_, new_n785_, new_n786_, new_n787_, new_n788_, new_n789_,
    new_n790_, new_n791_, new_n792_, new_n793_, new_n794_, new_n795_,
    new_n796_, new_n797_, new_n798_, new_n799_, new_n800_, new_n801_,
    new_n802_, new_n803_, new_n804_, new_n805_, new_n806_, new_n807_,
    new_n808_, new_n809_, new_n810_, new_n811_, new_n812_, new_n813_,
    new_n814_, new_n815_, new_n816_, new_n817_, new_n818_, new_n819_,
    new_n820_, new_n821_, new_n822_, new_n823_, new_n824_, new_n825_,
    new_n826_, new_n827_, new_n828_, new_n829_, new_n830_, new_n831_,
    new_n832_, new_n833_, new_n834_, new_n835_, new_n836_, new_n837_,
    new_n838_, new_n839_, new_n840_, new_n841_, new_n842_, new_n843_,
    new_n844_, new_n845_, new_n846_, new_n847_, new_n848_, new_n849_,
    new_n850_, new_n851_, new_n852_, new_n853_, new_n854_, new_n855_,
    new_n856_, new_n857_, new_n858_, new_n859_, new_n860_, new_n861_,
    new_n862_, new_n863_, new_n864_, new_n865_, new_n866_, new_n867_,
    new_n868_, new_n869_, new_n870_, new_n871_, new_n872_, new_n873_,
    new_n874_, new_n875_, new_n876_, new_n877_, new_n878_, new_n879_,
    new_n880_, new_n881_, new_n882_, new_n883_, new_n884_, new_n885_,
    new_n886_, new_n887_, new_n888_, new_n889_, new_n890_, new_n891_,
    new_n892_, new_n893_, new_n894_, new_n895_, new_n896_, new_n897_,
    new_n898_, new_n899_, new_n900_, new_n901_, new_n902_, new_n903_,
    new_n904_, new_n905_, new_n906_, new_n907_, new_n908_, new_n909_,
    new_n910_, new_n911_, new_n912_, new_n913_, new_n914_, new_n915_,
    new_n916_, new_n917_, new_n918_, new_n919_, new_n920_, new_n921_,
    new_n922_, new_n923_, new_n924_, new_n925_, new_n926_, new_n927_,
    new_n928_, new_n929_, new_n930_, new_n931_, new_n932_, new_n933_,
    new_n934_, new_n935_, new_n936_, new_n937_, new_n938_, new_n939_,
    new_n940_, new_n941_, new_n942_, new_n943_, new_n944_, new_n945_,
    new_n946_, new_n947_, new_n948_, new_n949_, new_n950_, new_n951_,
    new_n952_, new_n953_, new_n954_, new_n955_, new_n956_, new_n957_,
    new_n958_, new_n959_, new_n960_, new_n961_, new_n962_, new_n963_,
    new_n964_, new_n965_, new_n966_, new_n967_, new_n968_, new_n969_,
    new_n970_, new_n971_, new_n972_, new_n973_, new_n974_, new_n975_,
    new_n976_, new_n977_, new_n978_, new_n979_, new_n980_, new_n981_,
    new_n982_, new_n983_, new_n984_, new_n985_, new_n986_, new_n987_,
    new_n988_, new_n989_, new_n990_, new_n991_, new_n992_, new_n993_,
    new_n994_, new_n995_, new_n996_, new_n997_, new_n998_, new_n999_,
    new_n1000_, new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_,
    new_n1006_, new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_,
    new_n1012_, new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_,
    new_n1018_, new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_,
    new_n1024_, new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_,
    new_n1030_, new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_,
    new_n1036_, new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_,
    new_n1042_, new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_,
    new_n1048_, new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_,
    new_n1054_, new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_,
    new_n1060_, new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_,
    new_n1066_, new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_,
    new_n1072_, new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_,
    new_n1078_, new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_,
    new_n1084_, new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_,
    new_n1090_, new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_,
    new_n1096_, new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_,
    new_n1102_, new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_,
    new_n1108_, new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_,
    new_n1114_, new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_,
    new_n1120_, new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_,
    new_n1126_, new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_,
    new_n1132_, new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_,
    new_n1138_, new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_,
    new_n1144_, new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_,
    new_n1150_, new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_,
    new_n1156_, new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_,
    new_n1162_, new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_,
    new_n1168_, new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_,
    new_n1174_, new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_,
    new_n1180_, new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_,
    new_n1186_, new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_,
    new_n1192_, new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_,
    new_n1198_, new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_,
    new_n1204_, new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_,
    new_n1210_, new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_,
    new_n1216_, new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_,
    new_n1222_, new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_,
    new_n1228_, new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_,
    new_n1234_, new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_,
    new_n1240_, new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_,
    new_n1246_, new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_,
    new_n1252_, new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_,
    new_n1258_, new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_,
    new_n1264_, new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_,
    new_n1270_, new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_,
    new_n1276_, new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_,
    new_n1282_, new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_,
    new_n1288_, new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_,
    new_n1294_, new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_,
    new_n1300_, new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_,
    new_n1306_, new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_,
    new_n1312_, new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_,
    new_n1318_, new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_,
    new_n1324_, new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_,
    new_n1330_, new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_,
    new_n1336_, new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_,
    new_n1342_, new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_,
    new_n1348_, new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_,
    new_n1354_, new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_,
    new_n1360_, new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_,
    new_n1366_, new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_,
    new_n1372_, new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_,
    new_n1378_, new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_,
    new_n1384_, new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_,
    new_n1390_, new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_,
    new_n1396_, new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_,
    new_n1402_, new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_,
    new_n1408_, new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_,
    new_n1414_, new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_,
    new_n1420_, new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_,
    new_n1426_, new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_,
    new_n1432_, new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_,
    new_n1438_, new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_,
    new_n1444_, new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_,
    new_n1450_, new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_,
    new_n1456_, new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_,
    new_n1462_, new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_,
    new_n1468_, new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_,
    new_n1474_, new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_,
    new_n1480_, new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_,
    new_n1486_, new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_,
    new_n1492_, new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_,
    new_n1498_, new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_,
    new_n1504_, new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_,
    new_n1510_, new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_,
    new_n1516_, new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_,
    new_n1522_, new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_,
    new_n1528_, new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_,
    new_n1534_, new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_,
    new_n1540_, new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_,
    new_n1546_, new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_,
    new_n1552_, new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_,
    new_n1558_, new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_,
    new_n1564_, new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_,
    new_n1570_, new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_,
    new_n1576_, new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_,
    new_n1582_, new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_,
    new_n1588_, new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_,
    new_n1594_, new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_,
    new_n1600_, new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_,
    new_n1606_, new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_,
    new_n1612_, new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_,
    new_n1618_, new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_,
    new_n1624_, new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_,
    new_n1630_, new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_,
    new_n1636_, new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_,
    new_n1642_, new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_,
    new_n1648_, new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_,
    new_n1654_, new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_,
    new_n1660_, new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_,
    new_n1666_, new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_,
    new_n1672_, new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_,
    new_n1678_, new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_,
    new_n1684_, new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_,
    new_n1690_, new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_,
    new_n1696_, new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_,
    new_n1702_, new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_,
    new_n1708_, new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_,
    new_n1714_, new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_,
    new_n1720_, new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_,
    new_n1726_, new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_,
    new_n1732_, new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_,
    new_n1738_, new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_,
    new_n1744_, new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_,
    new_n1750_, new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_,
    new_n1756_, new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_,
    new_n1762_, new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_,
    new_n1768_, new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_,
    new_n1774_, new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_,
    new_n1780_, new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_,
    new_n1786_, new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_,
    new_n1792_, new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_,
    new_n1798_, new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_,
    new_n1804_, new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_,
    new_n1810_, new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_,
    new_n1816_, new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_,
    new_n1822_, new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_,
    new_n1828_, new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_,
    new_n1834_, new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_,
    new_n1840_, new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_,
    new_n1846_, new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_,
    new_n1852_, new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_,
    new_n1858_, new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_,
    new_n1864_, new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_,
    new_n1870_, new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_,
    new_n1876_, new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_,
    new_n1882_, new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_,
    new_n1888_, new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_,
    new_n1894_, new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_,
    new_n1900_, new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_,
    new_n1906_, new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_,
    new_n1912_, new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_,
    new_n1918_, new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_,
    new_n1924_, new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_,
    new_n1930_, new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_,
    new_n1936_, new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_,
    new_n1942_, new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_,
    new_n1948_, new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_,
    new_n1954_, new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_,
    new_n1960_, new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_,
    new_n1966_, new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_,
    new_n1972_, new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_,
    new_n1978_, new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_,
    new_n1984_, new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_,
    new_n1990_, new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_,
    new_n1996_, new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_,
    new_n2002_, new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_,
    new_n2008_, new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_,
    new_n2014_, new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_,
    new_n2020_, new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_,
    new_n2026_, new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_,
    new_n2032_, new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_,
    new_n2038_, new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_,
    new_n2044_, new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_,
    new_n2050_, new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_,
    new_n2056_, new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_,
    new_n2062_, new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_,
    new_n2068_, new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_,
    new_n2074_, new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_,
    new_n2080_, new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_,
    new_n2086_, new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_,
    new_n2092_, new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_,
    new_n2098_, new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_,
    new_n2104_, new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_,
    new_n2110_, new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_,
    new_n2116_, new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_,
    new_n2122_, new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_,
    new_n2128_, new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_,
    new_n2134_, new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_,
    new_n2140_, new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_,
    new_n2146_, new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_,
    new_n2152_, new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_,
    new_n2158_, new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_,
    new_n2164_, new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_,
    new_n2170_, new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_,
    new_n2176_, new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_,
    new_n2182_, new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_,
    new_n2188_, new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_,
    new_n2194_, new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_,
    new_n2200_, new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_,
    new_n2206_, new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_,
    new_n2212_, new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_,
    new_n2218_, new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_,
    new_n2224_, new_n2225_, new_n2226_, new_n2227_, new_n2228_, new_n2229_,
    new_n2230_, new_n2231_, new_n2232_, new_n2233_, new_n2234_, new_n2235_,
    new_n2236_, new_n2237_, new_n2238_, new_n2239_, new_n2240_, new_n2241_,
    new_n2242_, new_n2243_, new_n2244_, new_n2245_, new_n2246_, new_n2247_,
    new_n2248_, new_n2249_, new_n2250_, new_n2251_, new_n2252_, new_n2253_,
    new_n2254_, new_n2255_, new_n2256_, new_n2257_, new_n2258_, new_n2259_,
    new_n2260_, new_n2261_, new_n2262_, new_n2263_, new_n2264_, new_n2265_,
    new_n2266_, new_n2267_, new_n2268_, new_n2269_, new_n2270_, new_n2271_,
    new_n2272_, new_n2273_, new_n2274_, new_n2275_, new_n2276_, new_n2277_,
    new_n2278_, new_n2279_, new_n2280_, new_n2281_, new_n2282_, new_n2283_,
    new_n2284_, new_n2285_, new_n2286_, new_n2287_, new_n2288_, new_n2289_,
    new_n2290_, new_n2291_, new_n2292_, new_n2293_, new_n2294_, new_n2295_,
    new_n2296_, new_n2297_, new_n2298_, new_n2299_, new_n2300_, new_n2301_,
    new_n2302_, new_n2303_, new_n2304_, new_n2305_, new_n2306_, new_n2307_,
    new_n2308_, new_n2309_, new_n2310_, new_n2311_, new_n2312_, new_n2313_,
    new_n2314_, new_n2315_, new_n2316_, new_n2317_, new_n2318_, new_n2319_,
    new_n2320_, new_n2321_, new_n2322_, new_n2323_, new_n2324_, new_n2325_,
    new_n2326_, new_n2327_, new_n2328_, new_n2329_, new_n2330_, new_n2331_,
    new_n2332_, new_n2333_, new_n2334_, new_n2335_, new_n2336_, new_n2337_,
    new_n2338_, new_n2339_, new_n2340_, new_n2341_, new_n2342_, new_n2343_,
    new_n2344_, new_n2345_, new_n2346_, new_n2347_, new_n2348_, new_n2349_,
    new_n2350_, new_n2351_, new_n2352_, new_n2353_, new_n2354_, new_n2355_,
    new_n2356_, new_n2357_, new_n2358_, new_n2359_, new_n2360_, new_n2361_,
    new_n2362_, new_n2363_, new_n2364_, new_n2365_, new_n2366_, new_n2367_,
    new_n2368_, new_n2369_, new_n2370_, new_n2371_, new_n2372_, new_n2373_,
    new_n2374_, new_n2375_, new_n2376_, new_n2377_, new_n2378_, new_n2379_,
    new_n2380_, new_n2381_, new_n2382_, new_n2383_, new_n2384_, new_n2385_,
    new_n2386_, new_n2387_, new_n2388_, new_n2389_, new_n2390_, new_n2391_,
    new_n2392_, new_n2393_, new_n2394_, new_n2395_, new_n2396_, new_n2397_,
    new_n2398_, new_n2399_, new_n2400_, new_n2401_, new_n2402_, new_n2403_,
    new_n2404_, new_n2405_, new_n2406_, new_n2407_, new_n2408_, new_n2409_,
    new_n2410_, new_n2411_, new_n2412_, new_n2413_, new_n2414_, new_n2415_,
    new_n2416_, new_n2417_, new_n2418_, new_n2419_, new_n2420_, new_n2421_,
    new_n2422_, new_n2423_, new_n2424_, new_n2425_, new_n2426_, new_n2427_,
    new_n2428_, new_n2429_, new_n2430_, new_n2431_, new_n2432_, new_n2433_,
    new_n2434_, new_n2435_, new_n2436_, new_n2437_, new_n2438_, new_n2439_,
    new_n2440_, new_n2441_, new_n2442_, new_n2443_, new_n2444_, new_n2445_,
    new_n2446_, new_n2447_, new_n2448_, new_n2449_, new_n2450_, new_n2451_,
    new_n2452_, new_n2453_, new_n2454_, new_n2455_, new_n2456_, new_n2457_,
    new_n2458_, new_n2459_, new_n2460_, new_n2461_, new_n2462_, new_n2463_,
    new_n2464_, new_n2465_, new_n2466_, new_n2467_, new_n2468_, new_n2469_,
    new_n2470_, new_n2471_, new_n2472_, new_n2473_, new_n2474_, new_n2475_,
    new_n2476_, new_n2477_, new_n2478_, new_n2479_, new_n2480_, new_n2481_,
    new_n2482_, new_n2483_, new_n2484_, new_n2485_, new_n2486_, new_n2487_,
    new_n2488_, new_n2489_, new_n2490_, new_n2491_, new_n2492_, new_n2493_,
    new_n2494_, new_n2495_, new_n2496_, new_n2497_, new_n2498_, new_n2499_,
    new_n2500_, new_n2501_, new_n2502_, new_n2503_, new_n2504_, new_n2505_,
    new_n2506_, new_n2507_, new_n2508_, new_n2509_, new_n2510_, new_n2511_,
    new_n2512_, new_n2513_, new_n2514_, new_n2515_, new_n2516_, new_n2517_,
    new_n2518_, new_n2519_, new_n2520_, new_n2521_, new_n2522_, new_n2523_,
    new_n2524_, new_n2525_, new_n2526_, new_n2527_, new_n2528_, new_n2529_,
    new_n2530_, new_n2531_, new_n2532_, new_n2533_, new_n2534_, new_n2535_,
    new_n2536_, new_n2537_, new_n2538_, new_n2539_, new_n2540_, new_n2541_,
    new_n2542_, new_n2543_, new_n2544_, new_n2545_, new_n2546_, new_n2547_,
    new_n2548_, new_n2549_, new_n2550_, new_n2551_, new_n2552_, new_n2553_,
    new_n2554_, new_n2555_, new_n2556_, new_n2557_, new_n2558_, new_n2559_,
    new_n2560_, new_n2561_, new_n2562_, new_n2563_, new_n2564_, new_n2565_,
    new_n2566_, new_n2567_, new_n2568_, new_n2569_, new_n2570_, new_n2571_,
    new_n2572_, new_n2573_, new_n2574_, new_n2575_, new_n2576_, new_n2577_,
    new_n2578_, new_n2579_, new_n2580_, new_n2581_, new_n2582_, new_n2583_,
    new_n2584_, new_n2585_, new_n2586_, new_n2587_, new_n2588_, new_n2589_,
    new_n2590_, new_n2591_, new_n2592_, new_n2593_, new_n2594_, new_n2595_,
    new_n2596_, new_n2597_, new_n2598_, new_n2599_, new_n2600_, new_n2601_,
    new_n2602_, new_n2603_, new_n2604_, new_n2605_, new_n2606_, new_n2607_,
    new_n2608_, new_n2609_, new_n2610_, new_n2611_, new_n2612_, new_n2613_,
    new_n2614_, new_n2615_, new_n2616_, new_n2617_, new_n2618_, new_n2619_,
    new_n2620_, new_n2621_, new_n2622_, new_n2623_, new_n2624_, new_n2625_,
    new_n2626_, new_n2627_, new_n2628_, new_n2629_, new_n2630_, new_n2631_,
    new_n2632_, new_n2633_, new_n2634_, new_n2635_, new_n2636_, new_n2637_,
    new_n2638_, new_n2639_, new_n2640_, new_n2641_, new_n2642_, new_n2643_,
    new_n2644_, new_n2645_, new_n2646_, new_n2647_, new_n2648_, new_n2649_,
    new_n2650_, new_n2651_, new_n2652_, new_n2653_, new_n2654_, new_n2655_,
    new_n2656_, new_n2657_, new_n2658_, new_n2659_, new_n2660_, new_n2661_,
    new_n2662_, new_n2663_, new_n2664_, new_n2665_, new_n2666_, new_n2667_,
    new_n2668_, new_n2669_, new_n2670_, new_n2671_, new_n2672_, new_n2673_,
    new_n2674_, new_n2675_, new_n2676_, new_n2677_, new_n2678_, new_n2679_,
    new_n2680_, new_n2681_, new_n2682_, new_n2683_, new_n2684_, new_n2685_,
    new_n2686_, new_n2687_, new_n2688_, new_n2689_, new_n2690_, new_n2691_,
    new_n2692_, new_n2693_, new_n2694_, new_n2695_, new_n2696_, new_n2697_,
    new_n2698_, new_n2699_, new_n2700_, new_n2701_, new_n2702_, new_n2703_,
    new_n2704_, new_n2705_, new_n2706_, new_n2707_, new_n2708_, new_n2709_,
    new_n2710_, new_n2711_, new_n2712_, new_n2713_, new_n2714_, new_n2715_,
    new_n2716_, new_n2717_, new_n2718_, new_n2719_, new_n2720_, new_n2721_,
    new_n2722_, new_n2723_, new_n2724_, new_n2725_, new_n2726_, new_n2727_,
    new_n2728_, new_n2729_, new_n2730_, new_n2731_, new_n2732_, new_n2733_,
    new_n2734_, new_n2735_, new_n2736_, new_n2737_, new_n2738_, new_n2739_,
    new_n2740_, new_n2741_, new_n2742_, new_n2743_, new_n2744_, new_n2745_,
    new_n2746_, new_n2747_, new_n2748_, new_n2749_, new_n2750_, new_n2751_,
    new_n2752_, new_n2753_, new_n2754_, new_n2755_, new_n2756_, new_n2757_,
    new_n2758_, new_n2759_, new_n2760_, new_n2761_, new_n2762_, new_n2763_,
    new_n2764_, new_n2765_, new_n2766_, new_n2767_, new_n2768_, new_n2769_,
    new_n2770_, new_n2771_, new_n2772_, new_n2773_, new_n2774_, new_n2775_,
    new_n2776_, new_n2777_, new_n2778_, new_n2779_, new_n2780_, new_n2781_,
    new_n2782_, new_n2783_, new_n2784_, new_n2785_, new_n2786_, new_n2787_,
    new_n2788_, new_n2789_, new_n2790_, new_n2791_, new_n2792_, new_n2793_,
    new_n2794_, new_n2795_, new_n2796_, new_n2797_, new_n2798_, new_n2799_,
    new_n2800_, new_n2801_, new_n2802_, new_n2803_, new_n2804_, new_n2805_,
    new_n2806_, new_n2807_, new_n2808_, new_n2809_, new_n2810_, new_n2811_,
    new_n2812_, new_n2813_, new_n2814_, new_n2815_, new_n2816_, new_n2817_,
    new_n2818_, new_n2819_, new_n2820_, new_n2821_, new_n2822_, new_n2823_,
    new_n2824_, new_n2825_, new_n2826_, new_n2827_, new_n2828_, new_n2829_,
    new_n2830_, new_n2831_, new_n2832_, new_n2833_, new_n2834_, new_n2835_,
    new_n2836_, new_n2837_, new_n2838_, new_n2839_, new_n2840_, new_n2841_,
    new_n2842_, new_n2843_, new_n2844_, new_n2845_, new_n2846_, new_n2847_,
    new_n2848_, new_n2849_, new_n2850_, new_n2851_, new_n2852_, new_n2853_,
    new_n2854_, new_n2855_, new_n2856_, new_n2857_, new_n2858_, new_n2859_,
    new_n2860_, new_n2861_, new_n2862_, new_n2863_, new_n2864_, new_n2865_,
    new_n2866_, new_n2867_, new_n2868_, new_n2869_, new_n2870_, new_n2871_,
    new_n2872_, new_n2873_, new_n2874_, new_n2875_, new_n2876_, new_n2877_,
    new_n2878_, new_n2879_, new_n2880_, new_n2881_, new_n2882_, new_n2883_,
    new_n2884_, new_n2885_, new_n2886_, new_n2887_, new_n2888_, new_n2889_,
    new_n2890_, new_n2891_, new_n2892_, new_n2893_, new_n2894_, new_n2895_,
    new_n2896_, new_n2897_, new_n2898_, new_n2899_, new_n2900_, new_n2901_,
    new_n2902_, new_n2903_, new_n2904_, new_n2905_, new_n2906_, new_n2907_,
    new_n2908_, new_n2909_, new_n2910_, new_n2911_, new_n2912_, new_n2913_,
    new_n2914_, new_n2915_, new_n2916_, new_n2917_, new_n2918_, new_n2919_,
    new_n2920_, new_n2921_, new_n2922_, new_n2923_, new_n2924_, new_n2925_,
    new_n2926_, new_n2927_, new_n2928_, new_n2929_, new_n2930_, new_n2931_,
    new_n2932_, new_n2933_, new_n2934_, new_n2935_, new_n2936_, new_n2937_,
    new_n2938_, new_n2939_, new_n2940_, new_n2941_, new_n2942_, new_n2943_,
    new_n2944_, new_n2945_, new_n2946_, new_n2947_, new_n2948_, new_n2949_,
    new_n2950_, new_n2951_, new_n2952_, new_n2953_, new_n2954_, new_n2955_,
    new_n2956_, new_n2957_, new_n2958_, new_n2959_, new_n2960_, new_n2961_,
    new_n2962_, new_n2963_, new_n2964_, new_n2965_, new_n2966_, new_n2967_,
    new_n2968_, new_n2969_, new_n2970_, new_n2971_, new_n2972_, new_n2973_,
    new_n2974_, new_n2975_, new_n2976_, new_n2977_, new_n2978_, new_n2979_,
    new_n2980_, new_n2981_, new_n2982_, new_n2983_, new_n2984_, new_n2985_,
    new_n2986_, new_n2987_, new_n2988_, new_n2989_, new_n2990_, new_n2991_,
    new_n2992_, new_n2993_, new_n2994_, new_n2995_, new_n2996_, new_n2997_,
    new_n2998_, new_n2999_, new_n3000_, new_n3001_, new_n3002_, new_n3003_,
    new_n3004_, new_n3005_, new_n3006_, new_n3007_, new_n3008_, new_n3009_,
    new_n3010_, new_n3011_, new_n3012_, new_n3013_, new_n3014_, new_n3015_,
    new_n3016_, new_n3017_, new_n3018_, new_n3019_, new_n3020_, new_n3021_,
    new_n3022_, new_n3023_, new_n3024_, new_n3025_, new_n3026_, new_n3027_,
    new_n3028_, new_n3029_, new_n3030_, new_n3031_, new_n3032_, new_n3033_,
    new_n3034_, new_n3035_, new_n3036_, new_n3037_, new_n3038_, new_n3039_,
    new_n3040_, new_n3041_, new_n3042_, new_n3043_, new_n3044_, new_n3045_,
    new_n3046_, new_n3047_, new_n3048_, new_n3049_, new_n3050_, new_n3051_,
    new_n3052_, new_n3053_, new_n3054_, new_n3055_, new_n3056_, new_n3057_,
    new_n3058_, new_n3059_, new_n3060_, new_n3061_, new_n3062_, new_n3063_,
    new_n3064_, new_n3065_, new_n3066_, new_n3067_, new_n3068_, new_n3069_,
    new_n3070_, new_n3071_, new_n3072_, new_n3073_, new_n3074_, new_n3075_,
    new_n3076_, new_n3077_, new_n3078_, new_n3079_, new_n3080_, new_n3081_,
    new_n3082_, new_n3083_, new_n3084_, new_n3085_, new_n3086_, new_n3087_,
    new_n3088_, new_n3089_, new_n3090_, new_n3091_, new_n3092_, new_n3093_,
    new_n3094_, new_n3095_, new_n3096_, new_n3097_, new_n3098_, new_n3099_,
    new_n3100_, new_n3101_, new_n3102_, new_n3103_, new_n3104_, new_n3105_,
    new_n3106_, new_n3107_, new_n3108_, new_n3109_, new_n3110_, new_n3111_,
    new_n3112_, new_n3113_, new_n3114_, new_n3115_, new_n3116_, new_n3117_,
    new_n3118_, new_n3119_, new_n3120_, new_n3121_, new_n3122_, new_n3123_,
    new_n3124_, new_n3125_, new_n3126_, new_n3127_, new_n3128_, new_n3129_,
    new_n3130_, new_n3131_, new_n3132_, new_n3133_, new_n3134_, new_n3135_,
    new_n3136_, new_n3137_, new_n3138_, new_n3139_, new_n3140_, new_n3141_,
    new_n3142_, new_n3143_, new_n3144_, new_n3145_, new_n3146_, new_n3147_,
    new_n3148_, new_n3149_, new_n3150_, new_n3151_, new_n3152_, new_n3153_,
    new_n3154_, new_n3155_, new_n3156_, new_n3157_, new_n3158_, new_n3159_,
    new_n3160_, new_n3161_, new_n3162_, new_n3163_, new_n3164_, new_n3165_,
    new_n3166_, new_n3167_, new_n3168_, new_n3169_, new_n3170_, new_n3171_,
    new_n3172_, new_n3173_, new_n3174_, new_n3175_, new_n3176_, new_n3177_,
    new_n3178_, new_n3179_, new_n3180_, new_n3181_, new_n3182_, new_n3183_,
    new_n3184_, new_n3185_, new_n3186_, new_n3187_, new_n3188_, new_n3189_,
    new_n3190_, new_n3191_, new_n3192_, new_n3193_, new_n3194_, new_n3195_,
    new_n3196_, new_n3197_, new_n3198_, new_n3199_, new_n3200_, new_n3201_,
    new_n3202_, new_n3203_, new_n3204_, new_n3205_, new_n3206_, new_n3207_,
    new_n3208_, new_n3209_, new_n3210_, new_n3211_, new_n3212_, new_n3213_,
    new_n3214_, new_n3215_, new_n3216_, new_n3217_, new_n3218_, new_n3219_,
    new_n3220_, new_n3221_, new_n3222_, new_n3223_, new_n3224_, new_n3225_,
    new_n3226_, new_n3227_, new_n3228_, new_n3229_, new_n3230_, new_n3231_,
    new_n3232_, new_n3233_, new_n3234_, new_n3235_, new_n3236_, new_n3237_,
    new_n3238_, new_n3239_, new_n3240_, new_n3241_, new_n3242_, new_n3243_,
    new_n3244_, new_n3245_, new_n3246_, new_n3247_, new_n3248_, new_n3249_,
    new_n3250_, new_n3251_, new_n3252_, new_n3253_, new_n3254_, new_n3255_,
    new_n3256_, new_n3257_, new_n3258_, new_n3259_, new_n3260_, new_n3261_,
    new_n3262_, new_n3263_, new_n3264_, new_n3265_, new_n3266_, new_n3267_,
    new_n3268_, new_n3269_, new_n3270_, new_n3271_, new_n3272_, new_n3273_,
    new_n3274_, new_n3275_, new_n3276_, new_n3277_, new_n3278_, new_n3279_,
    new_n3280_, new_n3281_, new_n3282_, new_n3283_, new_n3284_, new_n3285_,
    new_n3286_, new_n3287_, new_n3288_, new_n3289_, new_n3290_, new_n3291_,
    new_n3292_, new_n3293_, new_n3294_, new_n3295_, new_n3296_, new_n3297_,
    new_n3298_, new_n3299_, new_n3300_, new_n3301_, new_n3302_, new_n3303_,
    new_n3304_, new_n3305_, new_n3306_, new_n3307_, new_n3308_, new_n3309_,
    new_n3310_, new_n3311_, new_n3312_, new_n3313_, new_n3314_, new_n3315_,
    new_n3316_, new_n3317_, new_n3318_, new_n3319_, new_n3320_, new_n3321_,
    new_n3322_, new_n3323_, new_n3324_, new_n3325_, new_n3326_, new_n3327_,
    new_n3328_, new_n3329_, new_n3330_, new_n3331_, new_n3332_, new_n3333_,
    new_n3334_, new_n3335_, new_n3336_, new_n3337_, new_n3338_, new_n3339_,
    new_n3340_, new_n3341_, new_n3342_, new_n3343_, new_n3344_, new_n3345_,
    new_n3346_, new_n3347_, new_n3348_, new_n3349_, new_n3350_, new_n3351_,
    new_n3352_, new_n3353_, new_n3354_, new_n3355_, new_n3356_, new_n3357_,
    new_n3358_, new_n3359_, new_n3360_, new_n3361_, new_n3362_, new_n3363_,
    new_n3364_, new_n3365_, new_n3366_, new_n3367_, new_n3368_, new_n3369_,
    new_n3370_, new_n3371_, new_n3372_, new_n3373_, new_n3374_, new_n3375_,
    new_n3376_, new_n3377_, new_n3378_, new_n3379_, new_n3380_, new_n3381_,
    new_n3382_, new_n3383_, new_n3384_, new_n3385_, new_n3386_, new_n3387_,
    new_n3388_, new_n3389_, new_n3390_, new_n3391_, new_n3392_, new_n3393_,
    new_n3394_, new_n3395_, new_n3396_, new_n3397_, new_n3398_, new_n3399_,
    new_n3400_, new_n3401_, new_n3402_, new_n3403_, new_n3404_, new_n3405_,
    new_n3406_, new_n3407_, new_n3408_, new_n3409_, new_n3410_, new_n3411_,
    new_n3412_, new_n3413_, new_n3414_, new_n3415_, new_n3416_, new_n3417_,
    new_n3418_, new_n3419_, new_n3420_, new_n3421_, new_n3422_, new_n3423_,
    new_n3424_, new_n3425_, new_n3426_, new_n3427_, new_n3428_, new_n3429_,
    new_n3430_, new_n3431_, new_n3432_, new_n3433_, new_n3434_, new_n3435_,
    new_n3436_, new_n3437_, new_n3438_, new_n3439_, new_n3440_, new_n3441_,
    new_n3442_, new_n3443_, new_n3444_, new_n3445_, new_n3446_, new_n3447_,
    new_n3448_, new_n3449_, new_n3450_, new_n3451_, new_n3452_, new_n3453_,
    new_n3454_, new_n3455_, new_n3456_, new_n3457_, new_n3458_, new_n3459_,
    new_n3460_, new_n3461_, new_n3462_, new_n3463_, new_n3464_, new_n3465_,
    new_n3466_, new_n3467_, new_n3468_, new_n3469_, new_n3470_, new_n3471_,
    new_n3472_, new_n3473_, new_n3474_, new_n3475_, new_n3476_, new_n3477_,
    new_n3478_, new_n3479_, new_n3480_, new_n3481_, new_n3482_, new_n3483_,
    new_n3484_, new_n3485_, new_n3486_, new_n3487_, new_n3488_, new_n3489_,
    new_n3490_, new_n3491_, new_n3492_, new_n3493_, new_n3494_, new_n3495_,
    new_n3496_, new_n3497_, new_n3498_, new_n3499_, new_n3500_, new_n3501_,
    new_n3502_, new_n3503_, new_n3504_, new_n3505_, new_n3506_, new_n3507_,
    new_n3508_, new_n3509_, new_n3510_, new_n3511_, new_n3512_, new_n3513_,
    new_n3514_, new_n3515_, new_n3516_, new_n3517_, new_n3518_, new_n3519_,
    new_n3520_, new_n3521_, new_n3522_, new_n3523_, new_n3524_, new_n3525_,
    new_n3526_, new_n3527_, new_n3528_, new_n3529_, new_n3530_, new_n3531_,
    new_n3532_, new_n3533_, new_n3534_, new_n3535_, new_n3536_, new_n3537_,
    new_n3538_, new_n3539_, new_n3540_, new_n3541_, new_n3542_, new_n3543_,
    new_n3544_, new_n3545_, new_n3546_, new_n3547_, new_n3548_, new_n3549_,
    new_n3550_, new_n3551_, new_n3552_, new_n3553_, new_n3554_, new_n3555_,
    new_n3556_, new_n3557_, new_n3558_, new_n3559_, new_n3560_, new_n3561_,
    new_n3562_, new_n3563_, new_n3564_, new_n3565_, new_n3566_, new_n3567_,
    new_n3568_, new_n3569_, new_n3570_, new_n3571_, new_n3572_, new_n3573_,
    new_n3574_, new_n3575_, new_n3576_, new_n3577_, new_n3578_, new_n3579_,
    new_n3580_, new_n3581_, new_n3582_, new_n3583_, new_n3584_, new_n3585_,
    new_n3586_, new_n3587_, new_n3588_, new_n3589_, new_n3590_, new_n3591_,
    new_n3592_, new_n3593_, new_n3594_, new_n3595_, new_n3596_, new_n3597_,
    new_n3598_, new_n3599_, new_n3600_, new_n3601_, new_n3602_, new_n3603_,
    new_n3604_, new_n3605_, new_n3606_, new_n3607_, new_n3608_, new_n3609_,
    new_n3610_, new_n3611_, new_n3612_, new_n3613_, new_n3614_, new_n3615_,
    new_n3616_, new_n3617_, new_n3618_, new_n3619_, new_n3620_, new_n3621_,
    new_n3622_, new_n3623_, new_n3624_, new_n3625_, new_n3626_, new_n3627_,
    new_n3628_, new_n3629_, new_n3630_, new_n3631_, new_n3632_, new_n3633_,
    new_n3634_, new_n3635_, new_n3636_, new_n3637_, new_n3638_, new_n3639_,
    new_n3640_, new_n3641_, new_n3642_, new_n3643_, new_n3644_, new_n3645_,
    new_n3646_, new_n3647_, new_n3648_, new_n3649_, new_n3650_, new_n3651_,
    new_n3652_, new_n3653_, new_n3654_, new_n3655_, new_n3656_, new_n3657_,
    new_n3658_, new_n3659_, new_n3660_, new_n3661_, new_n3662_, new_n3663_,
    new_n3664_, new_n3665_, new_n3666_, new_n3667_, new_n3668_, new_n3669_,
    new_n3670_, new_n3671_, new_n3672_, new_n3673_, new_n3674_, new_n3675_,
    new_n3676_, new_n3677_, new_n3678_, new_n3679_, new_n3680_, new_n3681_,
    new_n3682_, new_n3683_, new_n3684_, new_n3685_, new_n3686_, new_n3687_,
    new_n3688_, new_n3689_, new_n3690_, new_n3691_, new_n3692_, new_n3693_,
    new_n3694_, new_n3695_, new_n3696_, new_n3697_, new_n3698_, new_n3699_,
    new_n3700_, new_n3701_, new_n3702_, new_n3703_, new_n3704_, new_n3705_,
    new_n3706_, new_n3707_, new_n3708_, new_n3709_, new_n3710_, new_n3711_,
    new_n3712_, new_n3713_, new_n3714_, new_n3715_, new_n3716_, new_n3717_,
    new_n3718_, new_n3719_, new_n3720_, new_n3721_, new_n3722_, new_n3723_,
    new_n3724_, new_n3725_, new_n3726_, new_n3727_, new_n3728_, new_n3729_,
    new_n3730_, new_n3731_, new_n3732_, new_n3733_, new_n3734_, new_n3735_,
    new_n3736_, new_n3737_, new_n3738_, new_n3739_, new_n3740_, new_n3741_,
    new_n3742_, new_n3743_, new_n3744_, new_n3745_, new_n3746_, new_n3747_,
    new_n3748_, new_n3749_, new_n3750_, new_n3751_, new_n3752_, new_n3753_,
    new_n3754_, new_n3755_, new_n3756_, new_n3757_, new_n3758_, new_n3759_,
    new_n3760_, new_n3761_, new_n3762_, new_n3763_, new_n3764_, new_n3765_,
    new_n3766_, new_n3767_, new_n3768_, new_n3769_, new_n3770_, new_n3771_,
    new_n3772_, new_n3773_, new_n3774_, new_n3775_, new_n3776_, new_n3777_,
    new_n3778_, new_n3779_, new_n3780_, new_n3781_, new_n3782_, new_n3783_,
    new_n3784_, new_n3785_, new_n3786_, new_n3787_, new_n3788_, new_n3789_,
    new_n3790_, new_n3791_, new_n3792_, new_n3793_, new_n3794_, new_n3795_,
    new_n3796_, new_n3797_, new_n3798_, new_n3799_, new_n3800_, new_n3801_,
    new_n3802_, new_n3803_, new_n3804_, new_n3805_, new_n3806_, new_n3807_,
    new_n3808_, new_n3809_, new_n3810_, new_n3811_, new_n3812_, new_n3813_,
    new_n3814_, new_n3815_, new_n3816_, new_n3817_, new_n3818_, new_n3819_,
    new_n3820_, new_n3821_, new_n3822_, new_n3823_, new_n3824_, new_n3825_,
    new_n3826_, new_n3827_, new_n3828_, new_n3829_, new_n3830_, new_n3831_,
    new_n3832_, new_n3833_, new_n3834_, new_n3835_, new_n3836_, new_n3837_,
    new_n3838_, new_n3839_, new_n3840_, new_n3841_, new_n3842_, new_n3843_,
    new_n3844_, new_n3845_, new_n3846_, new_n3847_, new_n3848_, new_n3849_,
    new_n3850_, new_n3851_, new_n3852_, new_n3853_, new_n3854_, new_n3855_,
    new_n3856_, new_n3857_, new_n3858_, new_n3859_, new_n3860_, new_n3861_,
    new_n3862_, new_n3863_, new_n3864_, new_n3865_, new_n3866_, new_n3867_,
    new_n3868_, new_n3869_, new_n3870_, new_n3871_, new_n3872_, new_n3873_,
    new_n3874_, new_n3875_, new_n3876_, new_n3877_, new_n3878_, new_n3879_,
    new_n3880_, new_n3881_, new_n3882_, new_n3883_, new_n3884_, new_n3885_,
    new_n3886_, new_n3887_, new_n3888_, new_n3889_, new_n3890_, new_n3891_,
    new_n3892_, new_n3893_, new_n3894_, new_n3895_, new_n3896_, new_n3897_,
    new_n3898_, new_n3899_, new_n3900_, new_n3901_, new_n3902_, new_n3903_,
    new_n3904_, new_n3905_, new_n3906_, new_n3907_, new_n3908_, new_n3909_,
    new_n3910_, new_n3911_, new_n3912_, new_n3913_, new_n3914_, new_n3915_,
    new_n3916_, new_n3917_, new_n3918_, new_n3919_, new_n3920_, new_n3921_,
    new_n3922_, new_n3923_, new_n3924_, new_n3925_, new_n3926_, new_n3927_,
    new_n3928_, new_n3929_, new_n3930_, new_n3931_, new_n3932_, new_n3933_,
    new_n3934_, new_n3935_, new_n3936_, new_n3937_, new_n3938_, new_n3939_,
    new_n3940_, new_n3941_, new_n3942_, new_n3943_, new_n3944_, new_n3945_,
    new_n3946_, new_n3947_, new_n3948_, new_n3949_, new_n3950_, new_n3951_,
    new_n3952_, new_n3953_, new_n3954_, new_n3955_, new_n3956_, new_n3957_,
    new_n3958_, new_n3959_, new_n3960_, new_n3961_, new_n3962_, new_n3963_,
    new_n3964_, new_n3965_, new_n3966_, new_n3967_, new_n3968_, new_n3969_,
    new_n3970_, new_n3971_, new_n3972_, new_n3973_, new_n3974_, new_n3975_,
    new_n3976_, new_n3977_, new_n3978_, new_n3979_, new_n3980_, new_n3981_,
    new_n3982_, new_n3983_, new_n3984_, new_n3985_, new_n3986_, new_n3987_,
    new_n3988_, new_n3989_, new_n3990_, new_n3991_, new_n3992_, new_n3993_,
    new_n3994_, new_n3995_, new_n3996_, new_n3997_, new_n3998_, new_n3999_,
    new_n4000_, new_n4001_, new_n4002_, new_n4003_, new_n4004_, new_n4005_,
    new_n4006_, new_n4007_, new_n4008_, new_n4009_, new_n4010_, new_n4011_,
    new_n4012_, new_n4013_, new_n4014_, new_n4015_, new_n4016_, new_n4017_,
    new_n4018_, new_n4019_, new_n4020_, new_n4021_, new_n4022_, new_n4023_,
    new_n4024_, new_n4025_, new_n4026_, new_n4027_, new_n4028_, new_n4029_,
    new_n4030_, new_n4031_, new_n4032_, new_n4033_, new_n4034_, new_n4035_,
    new_n4036_, new_n4037_, new_n4038_, new_n4039_, new_n4040_, new_n4041_,
    new_n4042_, new_n4043_, new_n4044_, new_n4045_, new_n4046_, new_n4047_,
    new_n4048_, new_n4049_, new_n4050_, new_n4051_, new_n4052_, new_n4053_,
    new_n4054_, new_n4055_, new_n4056_, new_n4057_, new_n4058_, new_n4059_,
    new_n4060_, new_n4061_, new_n4062_, new_n4063_, new_n4064_, new_n4065_,
    new_n4066_, new_n4067_, new_n4068_, new_n4069_, new_n4070_, new_n4071_,
    new_n4072_, new_n4073_, new_n4074_, new_n4075_, new_n4076_, new_n4077_,
    new_n4078_, new_n4079_, new_n4080_, new_n4081_, new_n4082_, new_n4083_,
    new_n4084_, new_n4085_, new_n4086_, new_n4087_, new_n4088_, new_n4089_,
    new_n4090_, new_n4091_, new_n4092_, new_n4093_, new_n4094_, new_n4095_,
    new_n4096_, new_n4097_, new_n4098_, new_n4099_, new_n4100_, new_n4101_,
    new_n4102_, new_n4103_, new_n4104_, new_n4105_, new_n4106_, new_n4107_,
    new_n4108_, new_n4109_, new_n4110_, new_n4111_, new_n4112_, new_n4113_,
    new_n4114_, new_n4115_, new_n4116_, new_n4117_, new_n4118_, new_n4119_,
    new_n4120_, new_n4121_, new_n4122_, new_n4123_, new_n4124_, new_n4125_,
    new_n4126_, new_n4127_, new_n4128_, new_n4129_, new_n4130_, new_n4131_,
    new_n4132_, new_n4133_, new_n4134_, new_n4135_, new_n4136_, new_n4137_,
    new_n4138_, new_n4139_, new_n4140_, new_n4141_, new_n4142_, new_n4143_,
    new_n4144_, new_n4145_, new_n4146_, new_n4147_, new_n4148_, new_n4149_,
    new_n4150_, new_n4151_, new_n4152_, new_n4153_, new_n4154_, new_n4155_,
    new_n4156_, new_n4157_, new_n4158_, new_n4159_, new_n4160_, new_n4161_,
    new_n4162_, new_n4163_, new_n4164_, new_n4165_, new_n4166_, new_n4167_,
    new_n4168_, new_n4169_, new_n4170_, new_n4171_, new_n4172_, new_n4173_,
    new_n4174_, new_n4175_, new_n4176_, new_n4177_, new_n4178_, new_n4179_,
    new_n4180_, new_n4181_, new_n4182_, new_n4183_, new_n4184_, new_n4185_,
    new_n4186_, new_n4187_, new_n4188_, new_n4189_, new_n4190_, new_n4191_,
    new_n4192_, new_n4193_, new_n4194_, new_n4195_, new_n4196_, new_n4197_,
    new_n4198_, new_n4199_, new_n4200_, new_n4201_, new_n4202_, new_n4203_,
    new_n4204_, new_n4205_, new_n4206_, new_n4207_, new_n4208_, new_n4209_,
    new_n4210_, new_n4211_, new_n4212_, new_n4213_, new_n4214_, new_n4215_,
    new_n4216_, new_n4217_, new_n4218_, new_n4219_, new_n4220_, new_n4221_,
    new_n4222_, new_n4223_, new_n4224_, new_n4225_, new_n4226_, new_n4227_,
    new_n4228_, new_n4229_, new_n4230_, new_n4231_, new_n4232_, new_n4233_,
    new_n4234_, new_n4235_, new_n4236_, new_n4237_, new_n4238_, new_n4239_,
    new_n4240_, new_n4241_, new_n4242_, new_n4243_, new_n4244_, new_n4245_,
    new_n4246_, new_n4247_, new_n4248_, new_n4249_, new_n4250_, new_n4251_,
    new_n4252_, new_n4253_, new_n4254_, new_n4255_, new_n4256_, new_n4257_,
    new_n4258_, new_n4259_, new_n4260_, new_n4261_, new_n4262_, new_n4263_,
    new_n4264_, new_n4265_, new_n4266_, new_n4267_, new_n4268_, new_n4269_,
    new_n4270_, new_n4271_, new_n4272_, new_n4273_, new_n4274_, new_n4275_,
    new_n4276_, new_n4277_, new_n4278_, new_n4279_, new_n4280_, new_n4281_,
    new_n4282_, new_n4283_, new_n4284_, new_n4285_, new_n4286_, new_n4287_,
    new_n4288_, new_n4289_, new_n4290_, new_n4291_, new_n4292_, new_n4293_,
    new_n4294_, new_n4295_, new_n4296_, new_n4297_, new_n4298_, new_n4299_,
    new_n4300_, new_n4301_, new_n4302_, new_n4303_, new_n4304_, new_n4305_,
    new_n4306_, new_n4307_, new_n4308_, new_n4309_, new_n4310_, new_n4311_,
    new_n4312_, new_n4313_, new_n4314_, new_n4315_, new_n4316_, new_n4317_,
    new_n4318_, new_n4319_, new_n4320_, new_n4321_, new_n4322_, new_n4323_,
    new_n4324_, new_n4325_, new_n4326_, new_n4327_, new_n4328_, new_n4329_,
    new_n4330_, new_n4331_, new_n4332_, new_n4333_, new_n4334_, new_n4335_,
    new_n4336_, new_n4337_, new_n4338_, new_n4339_, new_n4340_, new_n4341_,
    new_n4342_, new_n4343_, new_n4344_, new_n4345_, new_n4346_, new_n4347_,
    new_n4348_, new_n4349_, new_n4350_, new_n4351_, new_n4352_, new_n4353_,
    new_n4354_, new_n4355_, new_n4356_, new_n4357_, new_n4358_, new_n4359_,
    new_n4360_, new_n4361_, new_n4362_, new_n4363_, new_n4364_, new_n4365_,
    new_n4366_, new_n4367_, new_n4368_, new_n4369_, new_n4370_, new_n4371_,
    new_n4372_, new_n4373_, new_n4374_, new_n4375_, new_n4376_, new_n4377_,
    new_n4378_, new_n4379_, new_n4380_, new_n4381_, new_n4382_, new_n4383_,
    new_n4384_, new_n4385_, new_n4386_, new_n4387_, new_n4388_, new_n4389_,
    new_n4390_, new_n4391_, new_n4392_, new_n4393_, new_n4394_, new_n4395_,
    new_n4396_, new_n4397_, new_n4398_, new_n4399_, new_n4400_, new_n4401_,
    new_n4402_, new_n4403_, new_n4404_, new_n4405_, new_n4406_, new_n4407_,
    new_n4408_, new_n4409_, new_n4410_, new_n4411_, new_n4412_, new_n4413_,
    new_n4414_, new_n4415_, new_n4416_, new_n4417_, new_n4418_, new_n4419_,
    new_n4420_, new_n4421_, new_n4422_, new_n4423_, new_n4424_, new_n4425_,
    new_n4426_, new_n4427_, new_n4428_, new_n4429_, new_n4430_, new_n4431_,
    new_n4432_, new_n4433_, new_n4434_, new_n4435_, new_n4436_, new_n4437_,
    new_n4438_, new_n4439_, new_n4440_, new_n4441_, new_n4442_, new_n4443_,
    new_n4444_, new_n4445_, new_n4446_, new_n4447_, new_n4448_, new_n4449_,
    new_n4450_, new_n4451_, new_n4452_, new_n4453_, new_n4454_, new_n4455_,
    new_n4456_, new_n4457_, new_n4458_, new_n4459_, new_n4460_, new_n4461_,
    new_n4462_, new_n4463_, new_n4464_, new_n4465_, new_n4466_, new_n4467_,
    new_n4468_, new_n4469_, new_n4470_, new_n4471_, new_n4472_, new_n4473_,
    new_n4474_, new_n4475_, new_n4476_, new_n4477_, new_n4478_, new_n4479_,
    new_n4480_, new_n4481_, new_n4482_, new_n4483_, new_n4484_, new_n4485_,
    new_n4486_, new_n4487_, new_n4488_, new_n4489_, new_n4490_, new_n4491_,
    new_n4492_, new_n4493_, new_n4494_, new_n4495_, new_n4496_, new_n4497_,
    new_n4498_, new_n4499_, new_n4500_, new_n4501_, new_n4502_, new_n4503_,
    new_n4504_, new_n4505_, new_n4506_, new_n4507_, new_n4508_, new_n4509_,
    new_n4510_, new_n4511_, new_n4512_, new_n4513_, new_n4514_, new_n4515_,
    new_n4516_, new_n4517_, new_n4518_, new_n4519_, new_n4520_, new_n4521_,
    new_n4522_, new_n4523_, new_n4524_, new_n4525_, new_n4526_, new_n4527_,
    new_n4528_, new_n4529_, new_n4530_, new_n4531_, new_n4532_, new_n4533_,
    new_n4534_, new_n4535_, new_n4536_, new_n4537_, new_n4538_, new_n4539_,
    new_n4540_, new_n4541_, new_n4542_, new_n4543_, new_n4544_, new_n4545_,
    new_n4546_, new_n4547_, new_n4548_, new_n4549_, new_n4550_, new_n4551_,
    new_n4552_, new_n4553_, new_n4554_, new_n4555_, new_n4556_, new_n4557_,
    new_n4558_, new_n4559_, new_n4560_, new_n4561_, new_n4562_, new_n4563_,
    new_n4564_, new_n4565_, new_n4566_, new_n4567_, new_n4568_, new_n4569_,
    new_n4570_, new_n4571_, new_n4572_, new_n4573_, new_n4574_, new_n4575_,
    new_n4576_, new_n4577_, new_n4578_, new_n4579_, new_n4580_, new_n4581_,
    new_n4582_, new_n4583_, new_n4584_, new_n4585_, new_n4586_, new_n4587_,
    new_n4588_, new_n4589_, new_n4590_, new_n4591_, new_n4592_, new_n4593_,
    new_n4594_, new_n4595_, new_n4596_, new_n4597_, new_n4598_, new_n4599_,
    new_n4600_, new_n4601_, new_n4602_, new_n4603_, new_n4604_, new_n4605_,
    new_n4606_, new_n4607_, new_n4608_, new_n4609_, new_n4610_, new_n4611_,
    new_n4612_, new_n4613_, new_n4614_, new_n4615_, new_n4616_, new_n4617_,
    new_n4618_, new_n4619_, new_n4620_, new_n4621_, new_n4622_, new_n4623_,
    new_n4624_, new_n4625_, new_n4626_, new_n4627_, new_n4628_, new_n4629_,
    new_n4630_, new_n4631_, new_n4632_, new_n4633_, new_n4634_, new_n4635_,
    new_n4636_, new_n4637_, new_n4638_, new_n4639_, new_n4640_, new_n4641_,
    new_n4642_, new_n4643_, new_n4644_, new_n4645_, new_n4646_, new_n4647_,
    new_n4648_, new_n4649_, new_n4650_, new_n4651_, new_n4652_, new_n4653_,
    new_n4654_, new_n4655_, new_n4656_, new_n4657_, new_n4658_, new_n4659_,
    new_n4660_, new_n4661_, new_n4662_, new_n4663_, new_n4664_, new_n4665_,
    new_n4666_, new_n4667_, new_n4668_, new_n4669_, new_n4670_, new_n4671_,
    new_n4672_, new_n4673_, new_n4674_, new_n4675_, new_n4676_, new_n4677_,
    new_n4678_, new_n4679_, new_n4680_, new_n4681_, new_n4682_, new_n4683_,
    new_n4684_, new_n4685_, new_n4686_, new_n4687_, new_n4688_, new_n4689_,
    new_n4690_, new_n4691_, new_n4692_, new_n4693_, new_n4694_, new_n4695_,
    new_n4696_, new_n4697_, new_n4698_, new_n4699_, new_n4700_, new_n4701_,
    new_n4702_, new_n4703_, new_n4704_, new_n4705_, new_n4706_, new_n4707_,
    new_n4708_, new_n4709_, new_n4710_, new_n4711_, new_n4712_, new_n4713_,
    new_n4714_, new_n4715_, new_n4716_, new_n4717_, new_n4718_, new_n4719_,
    new_n4720_, new_n4721_, new_n4722_, new_n4723_, new_n4724_, new_n4725_,
    new_n4726_, new_n4727_, new_n4728_, new_n4729_, new_n4730_, new_n4731_,
    new_n4732_, new_n4733_, new_n4734_, new_n4735_, new_n4736_, new_n4737_,
    new_n4738_, new_n4739_, new_n4740_, new_n4741_, new_n4742_, new_n4743_,
    new_n4744_, new_n4745_, new_n4746_, new_n4747_, new_n4748_, new_n4749_,
    new_n4750_, new_n4751_, new_n4752_, new_n4753_, new_n4754_, new_n4755_,
    new_n4756_, new_n4757_, new_n4758_, new_n4759_, new_n4760_, new_n4761_,
    new_n4762_, new_n4763_, new_n4764_, new_n4765_, new_n4766_, new_n4767_,
    new_n4768_, new_n4769_, new_n4770_, new_n4771_, new_n4772_, new_n4773_,
    new_n4774_, new_n4775_, new_n4776_, new_n4777_, new_n4778_, new_n4779_,
    new_n4780_, new_n4781_, new_n4782_, new_n4783_, new_n4784_, new_n4785_,
    new_n4786_, new_n4787_, new_n4788_, new_n4789_, new_n4790_, new_n4791_,
    new_n4792_, new_n4793_, new_n4794_, new_n4795_, new_n4796_, new_n4797_,
    new_n4798_, new_n4799_, new_n4800_, new_n4801_, new_n4802_, new_n4803_,
    new_n4804_, new_n4805_, new_n4806_, new_n4807_, new_n4808_, new_n4809_,
    new_n4810_, new_n4811_, new_n4812_, new_n4813_, new_n4814_, new_n4815_,
    new_n4816_, new_n4817_, new_n4818_, new_n4819_, new_n4820_, new_n4821_,
    new_n4822_, new_n4823_, new_n4824_, new_n4825_, new_n4826_, new_n4827_,
    new_n4828_, new_n4829_, new_n4830_, new_n4831_, new_n4832_, new_n4833_,
    new_n4834_, new_n4835_, new_n4836_, new_n4837_, new_n4838_, new_n4839_,
    new_n4840_, new_n4841_, new_n4842_, new_n4843_, new_n4844_, new_n4845_,
    new_n4846_, new_n4847_, new_n4848_, new_n4849_, new_n4850_, new_n4851_,
    new_n4852_, new_n4853_, new_n4854_, new_n4855_, new_n4856_, new_n4857_,
    new_n4858_, new_n4859_, new_n4860_, new_n4861_, new_n4862_, new_n4863_,
    new_n4864_, new_n4865_, new_n4866_, new_n4867_, new_n4868_, new_n4869_,
    new_n4870_, new_n4871_, new_n4872_, new_n4873_, new_n4874_, new_n4875_,
    new_n4876_, new_n4877_, new_n4878_, new_n4879_, new_n4880_, new_n4881_,
    new_n4882_, new_n4883_, new_n4884_, new_n4885_, new_n4886_, new_n4887_,
    new_n4888_, new_n4889_, new_n4890_, new_n4891_, new_n4892_, new_n4893_,
    new_n4894_, new_n4895_, new_n4896_, new_n4897_, new_n4898_, new_n4899_,
    new_n4900_, new_n4901_, new_n4902_, new_n4903_, new_n4904_, new_n4905_,
    new_n4906_, new_n4907_, new_n4908_, new_n4909_, new_n4910_, new_n4911_,
    new_n4912_, new_n4913_, new_n4914_, new_n4915_, new_n4916_, new_n4917_,
    new_n4918_, new_n4919_, new_n4920_, new_n4921_, new_n4922_, new_n4923_,
    new_n4924_, new_n4925_, new_n4926_, new_n4927_, new_n4928_, new_n4929_,
    new_n4930_, new_n4931_, new_n4932_, new_n4933_, new_n4934_, new_n4935_,
    new_n4936_, new_n4937_, new_n4938_, new_n4939_, new_n4940_, new_n4941_,
    new_n4942_, new_n4943_, new_n4944_, new_n4945_, new_n4946_, new_n4947_,
    new_n4948_, new_n4949_, new_n4950_, new_n4951_, new_n4952_, new_n4953_,
    new_n4954_, new_n4955_, new_n4956_, new_n4957_, new_n4958_, new_n4959_,
    new_n4960_, new_n4961_, new_n4962_, new_n4963_, new_n4964_, new_n4965_,
    new_n4966_, new_n4967_, new_n4968_, new_n4969_, new_n4970_, new_n4971_,
    new_n4972_, new_n4973_, new_n4974_, new_n4975_, new_n4976_, new_n4977_,
    new_n4978_, new_n4979_, new_n4980_, new_n4981_, new_n4982_, new_n4983_,
    new_n4984_, new_n4985_, new_n4986_, new_n4987_, new_n4988_, new_n4989_,
    new_n4990_, new_n4991_, new_n4992_, new_n4993_, new_n4994_, new_n4995_,
    new_n4996_, new_n4997_, new_n4998_, new_n4999_, new_n5000_, new_n5001_,
    new_n5002_, new_n5003_, new_n5004_, new_n5005_, new_n5006_, new_n5007_,
    new_n5008_, new_n5009_, new_n5010_, new_n5011_, new_n5012_, new_n5013_,
    new_n5014_, new_n5015_, new_n5016_, new_n5017_, new_n5018_, new_n5019_,
    new_n5020_, new_n5021_, new_n5022_, new_n5023_, new_n5024_, new_n5025_,
    new_n5026_, new_n5027_, new_n5028_, new_n5029_, new_n5030_, new_n5031_,
    new_n5032_, new_n5033_, new_n5034_, new_n5035_, new_n5036_, new_n5037_,
    new_n5038_, new_n5039_, new_n5040_, new_n5041_, new_n5042_, new_n5043_,
    new_n5044_, new_n5045_, new_n5046_, new_n5047_, new_n5048_, new_n5049_,
    new_n5050_, new_n5051_, new_n5052_, new_n5053_, new_n5054_, new_n5055_,
    new_n5056_, new_n5057_, new_n5058_, new_n5059_, new_n5060_, new_n5061_,
    new_n5062_, new_n5063_, new_n5064_, new_n5065_, new_n5066_, new_n5067_,
    new_n5068_, new_n5069_, new_n5070_, new_n5071_, new_n5072_, new_n5073_,
    new_n5074_, new_n5075_, new_n5076_, new_n5077_, new_n5078_, new_n5079_,
    new_n5080_, new_n5081_, new_n5082_, new_n5083_, new_n5084_, new_n5085_,
    new_n5086_, new_n5087_, new_n5088_, new_n5089_, new_n5090_, new_n5091_,
    new_n5092_, new_n5093_, new_n5094_, new_n5095_, new_n5096_, new_n5097_,
    new_n5098_, new_n5099_, new_n5100_, new_n5101_, new_n5102_, new_n5103_,
    new_n5104_, new_n5105_, new_n5106_, new_n5107_, new_n5108_, new_n5109_,
    new_n5110_, new_n5111_, new_n5112_, new_n5113_, new_n5114_, new_n5115_,
    new_n5116_, new_n5117_, new_n5118_, new_n5119_, new_n5120_, new_n5121_,
    new_n5122_, new_n5123_, new_n5124_, new_n5125_, new_n5126_, new_n5127_,
    new_n5128_, new_n5129_, new_n5130_, new_n5131_, new_n5132_, new_n5133_,
    new_n5134_, new_n5135_, new_n5136_, new_n5137_, new_n5138_, new_n5139_,
    new_n5140_, new_n5141_, new_n5142_, new_n5143_, new_n5144_, new_n5145_,
    new_n5146_, new_n5147_, new_n5148_, new_n5149_, new_n5150_, new_n5151_,
    new_n5152_, new_n5153_, new_n5154_, new_n5155_, new_n5156_, new_n5157_,
    new_n5158_, new_n5159_, new_n5160_, new_n5161_, new_n5162_, new_n5163_,
    new_n5164_, new_n5165_, new_n5166_, new_n5167_, new_n5168_, new_n5169_,
    new_n5170_, new_n5171_, new_n5172_, new_n5173_, new_n5174_, new_n5175_,
    new_n5176_, new_n5177_, new_n5178_, new_n5179_, new_n5180_, new_n5181_,
    new_n5182_, new_n5183_, new_n5184_, new_n5185_, new_n5186_, new_n5187_,
    new_n5188_, new_n5189_, new_n5190_, new_n5191_, new_n5192_, new_n5193_,
    new_n5194_, new_n5195_, new_n5196_, new_n5197_, new_n5198_, new_n5199_,
    new_n5200_, new_n5201_, new_n5202_, new_n5203_, new_n5204_, new_n5205_,
    new_n5206_, new_n5207_, new_n5208_, new_n5209_, new_n5210_, new_n5211_,
    new_n5212_, new_n5213_, new_n5214_, new_n5215_, new_n5216_, new_n5217_,
    new_n5218_, new_n5219_, new_n5220_, new_n5221_, new_n5222_, new_n5223_,
    new_n5224_, new_n5225_, new_n5226_, new_n5227_, new_n5228_, new_n5229_,
    new_n5230_, new_n5231_, new_n5232_, new_n5233_, new_n5234_, new_n5235_,
    new_n5236_, new_n5237_, new_n5238_, new_n5239_, new_n5240_, new_n5241_,
    new_n5242_, new_n5243_, new_n5244_, new_n5245_, new_n5246_, new_n5247_,
    new_n5248_, new_n5249_, new_n5250_, new_n5251_, new_n5252_, new_n5253_,
    new_n5254_, new_n5255_, new_n5256_, new_n5257_, new_n5258_, new_n5259_,
    new_n5260_, new_n5261_, new_n5262_, new_n5263_, new_n5264_, new_n5265_,
    new_n5266_, new_n5267_, new_n5268_, new_n5269_, new_n5270_, new_n5271_,
    new_n5272_, new_n5273_, new_n5274_, new_n5275_, new_n5276_, new_n5277_,
    new_n5278_, new_n5279_, new_n5280_, new_n5281_, new_n5282_, new_n5283_,
    new_n5284_, new_n5285_, new_n5286_, new_n5287_, new_n5288_, new_n5289_,
    new_n5290_, new_n5291_, new_n5292_, new_n5293_, new_n5294_, new_n5295_,
    new_n5296_, new_n5297_, new_n5298_, new_n5299_, new_n5300_, new_n5301_,
    new_n5302_, new_n5303_, new_n5304_, new_n5305_, new_n5306_, new_n5307_,
    new_n5308_, new_n5309_, new_n5310_, new_n5311_, new_n5312_, new_n5313_,
    new_n5314_, new_n5315_, new_n5316_, new_n5317_, new_n5318_, new_n5319_,
    new_n5320_, new_n5321_, new_n5322_, new_n5323_, new_n5324_, new_n5325_,
    new_n5326_, new_n5327_, new_n5328_, new_n5329_, new_n5330_, new_n5331_,
    new_n5332_, new_n5333_, new_n5334_, new_n5335_, new_n5336_, new_n5337_,
    new_n5338_, new_n5339_, new_n5340_, new_n5341_, new_n5342_, new_n5343_,
    new_n5344_, new_n5345_, new_n5346_, new_n5347_, new_n5348_, new_n5349_,
    new_n5350_, new_n5351_, new_n5352_, new_n5353_, new_n5354_, new_n5355_,
    new_n5356_, new_n5357_, new_n5358_, new_n5359_, new_n5360_, new_n5361_,
    new_n5362_, new_n5363_, new_n5364_, new_n5365_, new_n5366_, new_n5367_,
    new_n5368_, new_n5369_, new_n5370_, new_n5371_, new_n5372_, new_n5373_,
    new_n5374_, new_n5375_, new_n5376_, new_n5377_, new_n5378_, new_n5379_,
    new_n5380_, new_n5381_, new_n5382_, new_n5383_, new_n5384_, new_n5385_,
    new_n5386_, new_n5387_, new_n5388_, new_n5389_, new_n5390_, new_n5391_,
    new_n5392_, new_n5393_, new_n5394_, new_n5395_, new_n5396_, new_n5397_,
    new_n5398_, new_n5399_, new_n5400_, new_n5401_, new_n5402_, new_n5403_,
    new_n5404_, new_n5405_, new_n5406_, new_n5407_, new_n5408_, new_n5409_,
    new_n5410_, new_n5411_, new_n5412_, new_n5413_, new_n5414_, new_n5415_,
    new_n5416_, new_n5417_, new_n5418_, new_n5419_, new_n5420_, new_n5421_,
    new_n5422_, new_n5423_, new_n5424_, new_n5425_, new_n5426_, new_n5427_,
    new_n5428_, new_n5429_, new_n5430_, new_n5431_, new_n5432_, new_n5433_,
    new_n5434_, new_n5435_, new_n5436_, new_n5437_, new_n5438_, new_n5439_,
    new_n5440_, new_n5441_, new_n5442_, new_n5443_, new_n5444_, new_n5445_,
    new_n5446_, new_n5447_, new_n5448_, new_n5449_, new_n5450_, new_n5451_,
    new_n5452_, new_n5453_, new_n5454_, new_n5455_, new_n5456_, new_n5457_,
    new_n5458_, new_n5459_, new_n5460_, new_n5461_, new_n5462_, new_n5463_,
    new_n5464_, new_n5465_, new_n5466_, new_n5467_, new_n5468_, new_n5469_,
    new_n5470_, new_n5471_, new_n5472_, new_n5473_, new_n5474_, new_n5475_,
    new_n5476_, new_n5477_, new_n5478_, new_n5479_, new_n5480_, new_n5481_,
    new_n5482_, new_n5483_, new_n5484_, new_n5485_, new_n5486_, new_n5487_,
    new_n5488_, new_n5489_, new_n5490_, new_n5491_, new_n5492_, new_n5493_,
    new_n5494_, new_n5495_, new_n5496_, new_n5497_, new_n5498_, new_n5499_,
    new_n5500_, new_n5501_, new_n5502_, new_n5503_, new_n5504_, new_n5505_,
    new_n5506_, new_n5507_, new_n5508_, new_n5509_, new_n5510_, new_n5511_,
    new_n5512_, new_n5513_, new_n5514_, new_n5515_, new_n5516_, new_n5517_,
    new_n5518_, new_n5519_, new_n5520_, new_n5521_, new_n5522_, new_n5523_,
    new_n5524_, new_n5525_, new_n5526_, new_n5527_, new_n5528_, new_n5529_,
    new_n5530_, new_n5531_, new_n5532_, new_n5533_, new_n5534_, new_n5535_,
    new_n5536_, new_n5537_, new_n5538_, new_n5539_, new_n5540_, new_n5541_,
    new_n5542_, new_n5543_, new_n5544_, new_n5545_, new_n5546_, new_n5547_,
    new_n5548_, new_n5549_, new_n5550_, new_n5551_, new_n5552_, new_n5553_,
    new_n5554_, new_n5555_, new_n5556_, new_n5557_, new_n5558_, new_n5559_,
    new_n5560_, new_n5561_, new_n5562_, new_n5563_, new_n5564_, new_n5565_,
    new_n5566_, new_n5567_, new_n5568_, new_n5569_, new_n5570_, new_n5571_,
    new_n5572_, new_n5573_, new_n5574_, new_n5575_, new_n5576_, new_n5577_,
    new_n5578_, new_n5579_, new_n5580_, new_n5581_, new_n5582_, new_n5583_,
    new_n5584_, new_n5585_, new_n5586_, new_n5587_, new_n5588_, new_n5589_,
    new_n5590_, new_n5591_, new_n5592_, new_n5593_, new_n5594_, new_n5595_,
    new_n5596_, new_n5597_, new_n5598_, new_n5599_, new_n5600_, new_n5601_,
    new_n5602_, new_n5603_, new_n5604_, new_n5605_, new_n5606_, new_n5607_,
    new_n5608_, new_n5609_, new_n5610_, new_n5611_, new_n5612_, new_n5613_,
    new_n5614_, new_n5615_, new_n5616_, new_n5617_, new_n5618_, new_n5619_,
    new_n5620_, new_n5621_, new_n5622_, new_n5623_, new_n5624_, new_n5625_,
    new_n5626_, new_n5627_, new_n5628_, new_n5629_, new_n5630_, new_n5631_,
    new_n5632_, new_n5633_, new_n5634_, new_n5635_, new_n5636_, new_n5637_,
    new_n5638_, new_n5639_, new_n5640_, new_n5641_, new_n5642_, new_n5643_,
    new_n5644_, new_n5645_, new_n5646_, new_n5647_, new_n5648_, new_n5649_,
    new_n5650_, new_n5651_, new_n5652_, new_n5653_, new_n5654_, new_n5655_,
    new_n5656_, new_n5657_, new_n5658_, new_n5659_, new_n5660_, new_n5661_,
    new_n5662_, new_n5663_, new_n5664_, new_n5665_, new_n5666_, new_n5667_,
    new_n5668_, new_n5669_, new_n5670_, new_n5671_, new_n5672_, new_n5673_,
    new_n5674_, new_n5675_, new_n5676_, new_n5677_, new_n5678_, new_n5679_,
    new_n5680_, new_n5681_, new_n5682_, new_n5683_, new_n5684_, new_n5685_,
    new_n5686_, new_n5687_, new_n5688_, new_n5689_, new_n5690_, new_n5691_,
    new_n5692_, new_n5693_, new_n5694_, new_n5695_, new_n5696_, new_n5697_,
    new_n5698_, new_n5699_, new_n5700_, new_n5701_, new_n5702_, new_n5703_,
    new_n5704_, new_n5705_, new_n5706_, new_n5707_, new_n5708_, new_n5709_,
    new_n5710_, new_n5711_, new_n5712_, new_n5713_, new_n5714_, new_n5715_,
    new_n5716_, new_n5717_, new_n5718_, new_n5719_, new_n5720_, new_n5721_,
    new_n5722_, new_n5723_, new_n5724_, new_n5725_, new_n5726_, new_n5727_,
    new_n5728_, new_n5729_, new_n5730_, new_n5731_, new_n5732_, new_n5733_,
    new_n5734_, new_n5735_, new_n5736_, new_n5737_, new_n5738_, new_n5739_,
    new_n5740_, new_n5741_, new_n5742_, new_n5743_, new_n5744_, new_n5745_,
    new_n5746_, new_n5747_, new_n5748_, new_n5749_, new_n5750_, new_n5751_,
    new_n5752_, new_n5753_, new_n5754_, new_n5755_, new_n5756_, new_n5757_,
    new_n5758_, new_n5759_, new_n5760_, new_n5761_, new_n5762_, new_n5763_,
    new_n5764_, new_n5765_, new_n5766_, new_n5767_, new_n5768_, new_n5769_,
    new_n5770_, new_n5771_, new_n5772_, new_n5773_, new_n5774_, new_n5775_,
    new_n5776_, new_n5777_, new_n5778_, new_n5779_, new_n5780_, new_n5781_,
    new_n5782_, new_n5783_, new_n5784_, new_n5785_, new_n5786_, new_n5787_,
    new_n5788_, new_n5789_, new_n5790_, new_n5791_, new_n5792_, new_n5793_,
    new_n5794_, new_n5795_, new_n5796_, new_n5797_, new_n5798_, new_n5799_,
    new_n5800_, new_n5801_, new_n5802_, new_n5803_, new_n5804_, new_n5805_,
    new_n5806_, new_n5807_, new_n5808_, new_n5809_, new_n5810_, new_n5811_,
    new_n5812_, new_n5813_, new_n5814_, new_n5815_, new_n5816_, new_n5817_,
    new_n5818_, new_n5819_, new_n5820_, new_n5821_, new_n5822_, new_n5823_,
    new_n5824_, new_n5825_, new_n5826_, new_n5827_, new_n5828_, new_n5829_,
    new_n5830_, new_n5831_, new_n5832_, new_n5833_, new_n5834_, new_n5835_,
    new_n5836_, new_n5837_, new_n5838_, new_n5839_, new_n5840_, new_n5841_,
    new_n5842_, new_n5843_, new_n5844_, new_n5845_, new_n5846_, new_n5847_,
    new_n5848_, new_n5849_, new_n5850_, new_n5851_, new_n5852_, new_n5853_,
    new_n5854_, new_n5855_, new_n5856_, new_n5857_, new_n5858_, new_n5859_,
    new_n5860_, new_n5861_, new_n5862_, new_n5863_, new_n5864_, new_n5865_,
    new_n5866_, new_n5867_, new_n5868_, new_n5869_, new_n5870_, new_n5871_,
    new_n5872_, new_n5873_, new_n5874_, new_n5875_, new_n5876_, new_n5877_,
    new_n5878_, new_n5879_, new_n5880_, new_n5881_, new_n5882_, new_n5883_,
    new_n5884_, new_n5885_, new_n5886_, new_n5887_, new_n5888_, new_n5889_,
    new_n5890_, new_n5891_, new_n5892_, new_n5893_, new_n5894_, new_n5895_,
    new_n5896_, new_n5897_, new_n5898_, new_n5899_, new_n5900_, new_n5901_,
    new_n5902_, new_n5903_, new_n5904_, new_n5905_, new_n5906_, new_n5907_,
    new_n5908_, new_n5909_, new_n5910_, new_n5911_, new_n5912_, new_n5913_,
    new_n5914_, new_n5915_, new_n5916_, new_n5917_, new_n5918_, new_n5919_,
    new_n5920_, new_n5921_, new_n5922_, new_n5923_, new_n5924_, new_n5925_,
    new_n5926_, new_n5927_, new_n5928_, new_n5929_, new_n5930_, new_n5931_,
    new_n5932_, new_n5933_, new_n5934_, new_n5935_, new_n5936_, new_n5937_,
    new_n5938_, new_n5939_, new_n5940_, new_n5941_, new_n5942_, new_n5943_,
    new_n5944_, new_n5945_, new_n5946_, new_n5947_, new_n5948_, new_n5949_,
    new_n5950_, new_n5951_, new_n5952_, new_n5953_, new_n5954_, new_n5955_,
    new_n5956_, new_n5957_, new_n5958_, new_n5959_, new_n5960_, new_n5961_,
    new_n5962_, new_n5963_, new_n5964_, new_n5965_, new_n5966_, new_n5967_,
    new_n5968_, new_n5969_, new_n5970_, new_n5971_, new_n5972_, new_n5973_,
    new_n5974_, new_n5975_, new_n5976_, new_n5977_, new_n5978_, new_n5979_,
    new_n5980_, new_n5981_, new_n5982_, new_n5983_, new_n5984_, new_n5985_,
    new_n5986_, new_n5987_, new_n5988_, new_n5989_, new_n5990_, new_n5991_,
    new_n5992_, new_n5993_, new_n5994_, new_n5995_, new_n5996_, new_n5997_,
    new_n5998_, new_n5999_, new_n6000_, new_n6001_, new_n6002_, new_n6003_,
    new_n6004_, new_n6005_, new_n6006_, new_n6007_, new_n6008_, new_n6009_,
    new_n6010_, new_n6011_, new_n6012_, new_n6013_, new_n6014_, new_n6015_,
    new_n6016_, new_n6017_, new_n6018_, new_n6019_, new_n6020_, new_n6021_,
    new_n6022_, new_n6023_, new_n6024_, new_n6025_, new_n6026_, new_n6027_,
    new_n6028_, new_n6029_, new_n6030_, new_n6031_, new_n6032_, new_n6033_,
    new_n6034_, new_n6035_, new_n6036_, new_n6037_, new_n6038_, new_n6039_,
    new_n6040_, new_n6041_, new_n6042_, new_n6043_, new_n6044_, new_n6045_,
    new_n6046_, new_n6047_, new_n6048_, new_n6049_, new_n6050_, new_n6051_,
    new_n6052_, new_n6053_, new_n6054_, new_n6055_, new_n6056_, new_n6057_,
    new_n6058_, new_n6059_, new_n6060_, new_n6061_, new_n6062_, new_n6063_,
    new_n6064_, new_n6065_, new_n6066_, new_n6067_, new_n6068_, new_n6069_,
    new_n6070_, new_n6071_, new_n6072_, new_n6073_, new_n6074_, new_n6075_,
    new_n6076_, new_n6077_, new_n6078_, new_n6079_, new_n6080_, new_n6081_,
    new_n6082_, new_n6083_, new_n6084_, new_n6085_, new_n6086_, new_n6087_,
    new_n6088_, new_n6089_, new_n6090_, new_n6091_, new_n6092_, new_n6093_,
    new_n6094_, new_n6095_, new_n6096_, new_n6097_, new_n6098_, new_n6099_,
    new_n6100_, new_n6101_, new_n6102_, new_n6103_, new_n6104_, new_n6105_,
    new_n6106_, new_n6107_, new_n6108_, new_n6109_, new_n6110_, new_n6111_,
    new_n6112_, new_n6113_, new_n6114_, new_n6115_, new_n6116_, new_n6117_,
    new_n6118_, new_n6119_, new_n6120_, new_n6121_, new_n6122_, new_n6123_,
    new_n6124_, new_n6125_, new_n6126_, new_n6127_, new_n6128_, new_n6129_,
    new_n6130_, new_n6131_, new_n6132_, new_n6133_, new_n6134_, new_n6135_,
    new_n6136_, new_n6137_, new_n6138_, new_n6139_, new_n6140_, new_n6141_,
    new_n6142_, new_n6143_, new_n6144_, new_n6145_, new_n6146_, new_n6147_,
    new_n6148_, new_n6149_, new_n6150_, new_n6151_, new_n6152_, new_n6153_,
    new_n6154_, new_n6155_, new_n6156_, new_n6157_, new_n6158_, new_n6159_,
    new_n6160_, new_n6161_, new_n6162_, new_n6163_, new_n6164_, new_n6165_,
    new_n6166_, new_n6167_, new_n6168_, new_n6169_, new_n6170_, new_n6171_,
    new_n6172_, new_n6173_, new_n6174_, new_n6175_, new_n6176_, new_n6177_,
    new_n6178_, new_n6179_, new_n6180_, new_n6181_, new_n6182_, new_n6183_,
    new_n6184_, new_n6185_, new_n6186_, new_n6187_, new_n6188_, new_n6189_,
    new_n6190_, new_n6191_, new_n6192_, new_n6193_, new_n6194_, new_n6195_,
    new_n6196_, new_n6197_, new_n6198_, new_n6199_, new_n6200_, new_n6201_,
    new_n6202_, new_n6203_, new_n6204_, new_n6205_, new_n6206_, new_n6207_,
    new_n6208_, new_n6209_, new_n6210_, new_n6211_, new_n6212_, new_n6213_,
    new_n6214_, new_n6215_, new_n6216_, new_n6217_, new_n6218_, new_n6219_,
    new_n6220_, new_n6221_, new_n6222_, new_n6223_, new_n6224_, new_n6225_,
    new_n6226_, new_n6227_, new_n6228_, new_n6229_, new_n6230_, new_n6231_,
    new_n6232_, new_n6233_, new_n6234_, new_n6235_, new_n6236_, new_n6237_,
    new_n6238_, new_n6239_, new_n6240_, new_n6241_, new_n6242_, new_n6243_,
    new_n6244_, new_n6245_, new_n6246_, new_n6247_, new_n6248_, new_n6249_,
    new_n6250_, new_n6251_, new_n6252_, new_n6253_, new_n6254_, new_n6255_,
    new_n6256_, new_n6257_, new_n6258_, new_n6259_, new_n6260_, new_n6261_,
    new_n6262_, new_n6263_, new_n6264_, new_n6265_, new_n6266_, new_n6267_,
    new_n6268_, new_n6269_, new_n6270_, new_n6271_, new_n6272_, new_n6273_,
    new_n6274_, new_n6275_, new_n6276_, new_n6277_, new_n6278_, new_n6279_,
    new_n6280_, new_n6281_, new_n6282_, new_n6283_, new_n6284_, new_n6285_,
    new_n6286_, new_n6287_, new_n6288_, new_n6289_, new_n6290_, new_n6291_,
    new_n6292_, new_n6293_, new_n6294_, new_n6295_, new_n6296_, new_n6297_,
    new_n6298_, new_n6299_, new_n6300_, new_n6301_, new_n6302_, new_n6303_,
    new_n6304_, new_n6305_, new_n6306_, new_n6307_, new_n6308_, new_n6309_,
    new_n6310_, new_n6311_, new_n6312_, new_n6313_, new_n6314_, new_n6315_,
    new_n6316_, new_n6317_, new_n6318_, new_n6319_, new_n6320_, new_n6321_,
    new_n6322_, new_n6323_, new_n6324_, new_n6325_, new_n6326_, new_n6327_,
    new_n6328_, new_n6329_, new_n6330_, new_n6331_, new_n6332_, new_n6333_,
    new_n6334_, new_n6335_, new_n6336_, new_n6337_, new_n6338_, new_n6339_,
    new_n6340_, new_n6341_, new_n6342_, new_n6343_, new_n6344_, new_n6345_,
    new_n6346_, new_n6347_, new_n6348_, new_n6349_, new_n6350_, new_n6351_,
    new_n6352_, new_n6353_, new_n6354_, new_n6355_, new_n6356_, new_n6357_,
    new_n6358_, new_n6359_, new_n6360_, new_n6361_, new_n6362_, new_n6363_,
    new_n6364_, new_n6365_, new_n6366_, new_n6367_, new_n6368_, new_n6369_,
    new_n6370_, new_n6371_, new_n6372_, new_n6373_, new_n6374_, new_n6375_,
    new_n6376_, new_n6377_, new_n6378_, new_n6379_, new_n6380_, new_n6381_,
    new_n6382_, new_n6383_, new_n6384_, new_n6385_, new_n6386_, new_n6387_,
    new_n6388_, new_n6389_, new_n6390_, new_n6391_, new_n6392_, new_n6393_,
    new_n6394_, new_n6395_, new_n6396_, new_n6397_, new_n6398_, new_n6399_,
    new_n6400_, new_n6401_, new_n6402_, new_n6403_, new_n6404_, new_n6405_,
    new_n6406_, new_n6407_, new_n6408_, new_n6409_, new_n6410_, new_n6411_,
    new_n6412_, new_n6413_, new_n6414_, new_n6415_, new_n6416_, new_n6417_,
    new_n6418_, new_n6419_, new_n6420_, new_n6421_, new_n6422_, new_n6423_,
    new_n6424_, new_n6425_, new_n6426_, new_n6427_, new_n6428_, new_n6429_,
    new_n6430_, new_n6431_, new_n6432_, new_n6433_, new_n6434_, new_n6435_,
    new_n6436_, new_n6437_, new_n6438_, new_n6439_, new_n6440_, new_n6441_,
    new_n6442_, new_n6443_, new_n6444_, new_n6445_, new_n6446_, new_n6447_,
    new_n6448_, new_n6449_, new_n6450_, new_n6451_, new_n6452_, new_n6453_,
    new_n6454_, new_n6455_, new_n6456_, new_n6457_, new_n6458_, new_n6459_,
    new_n6460_, new_n6461_, new_n6462_, new_n6463_, new_n6464_, new_n6465_,
    new_n6466_, new_n6467_, new_n6468_, new_n6469_, new_n6470_, new_n6471_,
    new_n6472_, new_n6473_, new_n6474_, new_n6475_, new_n6476_, new_n6477_,
    new_n6478_, new_n6479_, new_n6480_, new_n6481_, new_n6482_, new_n6483_,
    new_n6484_, new_n6485_, new_n6486_, new_n6487_, new_n6488_, new_n6489_,
    new_n6490_, new_n6491_, new_n6492_, new_n6493_, new_n6494_, new_n6495_,
    new_n6496_, new_n6497_, new_n6498_, new_n6499_, new_n6500_, new_n6501_,
    new_n6502_, new_n6503_, new_n6504_, new_n6505_, new_n6506_, new_n6507_,
    new_n6508_, new_n6509_, new_n6510_, new_n6511_, new_n6512_, new_n6513_,
    new_n6514_, new_n6515_, new_n6516_, new_n6517_, new_n6518_, new_n6519_,
    new_n6520_, new_n6521_, new_n6522_, new_n6523_, new_n6524_, new_n6525_,
    new_n6526_, new_n6527_, new_n6528_, new_n6529_, new_n6530_, new_n6531_,
    new_n6532_, new_n6533_, new_n6534_, new_n6535_, new_n6536_, new_n6537_,
    new_n6538_, new_n6539_, new_n6540_, new_n6541_, new_n6542_, new_n6543_,
    new_n6544_, new_n6545_, new_n6546_, new_n6547_, new_n6548_, new_n6549_,
    new_n6550_, new_n6551_, new_n6552_, new_n6553_, new_n6554_, new_n6555_,
    new_n6556_, new_n6557_, new_n6558_, new_n6559_, new_n6560_, new_n6561_,
    new_n6562_, new_n6563_, new_n6564_, new_n6565_, new_n6566_, new_n6567_,
    new_n6568_, new_n6569_, new_n6570_, new_n6571_, new_n6572_, new_n6573_,
    new_n6574_, new_n6575_, new_n6576_, new_n6577_, new_n6578_, new_n6579_,
    new_n6580_, new_n6581_, new_n6582_, new_n6583_, new_n6584_, new_n6585_,
    new_n6586_, new_n6587_, new_n6588_, new_n6589_, new_n6590_, new_n6591_,
    new_n6592_, new_n6593_, new_n6594_, new_n6595_, new_n6596_, new_n6597_,
    new_n6598_, new_n6599_, new_n6600_, new_n6601_, new_n6602_, new_n6603_,
    new_n6604_, new_n6605_, new_n6606_, new_n6607_, new_n6608_, new_n6609_,
    new_n6610_, new_n6611_, new_n6612_, new_n6613_, new_n6614_, new_n6615_,
    new_n6616_, new_n6617_, new_n6618_, new_n6619_, new_n6620_, new_n6621_,
    new_n6622_, new_n6623_, new_n6624_, new_n6625_, new_n6626_, new_n6627_,
    new_n6628_, new_n6629_, new_n6630_, new_n6631_, new_n6632_, new_n6633_,
    new_n6634_, new_n6635_, new_n6636_, new_n6637_, new_n6638_, new_n6639_,
    new_n6640_, new_n6641_, new_n6642_, new_n6643_, new_n6644_, new_n6645_,
    new_n6646_, new_n6647_, new_n6648_, new_n6649_, new_n6650_, new_n6651_,
    new_n6652_, new_n6653_, new_n6654_, new_n6655_, new_n6656_, new_n6657_,
    new_n6658_, new_n6659_, new_n6660_, new_n6661_, new_n6662_, new_n6663_,
    new_n6664_, new_n6665_, new_n6666_, new_n6667_, new_n6668_, new_n6669_,
    new_n6670_, new_n6671_, new_n6672_, new_n6673_, new_n6674_, new_n6675_,
    new_n6676_, new_n6677_, new_n6678_, new_n6679_, new_n6680_, new_n6681_,
    new_n6682_, new_n6683_, new_n6684_, new_n6685_, new_n6686_, new_n6687_,
    new_n6688_, new_n6689_, new_n6690_, new_n6691_, new_n6692_, new_n6693_,
    new_n6694_, new_n6695_, new_n6696_, new_n6697_, new_n6698_, new_n6699_,
    new_n6700_, new_n6701_, new_n6702_, new_n6703_, new_n6704_, new_n6705_,
    new_n6706_, new_n6707_, new_n6708_, new_n6709_, new_n6710_, new_n6711_,
    new_n6712_, new_n6713_, new_n6714_, new_n6715_, new_n6716_, new_n6717_,
    new_n6718_, new_n6719_, new_n6720_, new_n6721_, new_n6722_, new_n6723_,
    new_n6724_, new_n6725_, new_n6726_, new_n6727_, new_n6728_, new_n6729_,
    new_n6730_, new_n6731_, new_n6732_, new_n6733_, new_n6734_, new_n6735_,
    new_n6736_, new_n6737_, new_n6738_, new_n6739_, new_n6740_, new_n6741_,
    new_n6742_, new_n6743_, new_n6744_, new_n6745_, new_n6746_, new_n6747_,
    new_n6748_, new_n6749_, new_n6750_, new_n6751_, new_n6752_, new_n6753_,
    new_n6754_, new_n6755_, new_n6756_, new_n6757_, new_n6758_, new_n6759_,
    new_n6760_, new_n6761_, new_n6762_, new_n6763_, new_n6764_, new_n6765_,
    new_n6766_, new_n6767_, new_n6768_, new_n6769_, new_n6770_, new_n6771_,
    new_n6772_, new_n6773_, new_n6774_, new_n6775_, new_n6776_, new_n6777_,
    new_n6778_, new_n6779_, new_n6780_, new_n6781_, new_n6782_, new_n6783_,
    new_n6784_, new_n6785_, new_n6786_, new_n6787_, new_n6788_, new_n6789_,
    new_n6790_, new_n6791_, new_n6792_, new_n6793_, new_n6794_, new_n6795_,
    new_n6796_, new_n6797_, new_n6798_, new_n6799_, new_n6800_, new_n6801_,
    new_n6802_, new_n6803_, new_n6804_, new_n6805_, new_n6806_, new_n6807_,
    new_n6808_, new_n6809_, new_n6810_, new_n6811_, new_n6812_, new_n6813_,
    new_n6814_, new_n6815_, new_n6816_, new_n6817_, new_n6818_, new_n6819_,
    new_n6820_, new_n6821_, new_n6822_, new_n6823_, new_n6824_, new_n6825_,
    new_n6826_, new_n6827_, new_n6828_, new_n6829_, new_n6830_, new_n6831_,
    new_n6832_, new_n6833_, new_n6834_, new_n6835_, new_n6836_, new_n6837_,
    new_n6838_, new_n6839_, new_n6840_, new_n6841_, new_n6842_, new_n6843_,
    new_n6844_, new_n6845_, new_n6846_, new_n6847_, new_n6848_, new_n6849_,
    new_n6850_, new_n6851_, new_n6852_, new_n6853_, new_n6854_, new_n6855_,
    new_n6856_, new_n6857_, new_n6858_, new_n6859_, new_n6860_, new_n6861_,
    new_n6862_, new_n6863_, new_n6864_, new_n6865_, new_n6866_, new_n6867_,
    new_n6868_, new_n6869_, new_n6870_, new_n6871_, new_n6872_, new_n6873_,
    new_n6874_, new_n6875_, new_n6876_, new_n6877_, new_n6878_, new_n6879_,
    new_n6880_, new_n6881_, new_n6882_, new_n6883_, new_n6884_, new_n6885_,
    new_n6886_, new_n6887_, new_n6888_, new_n6889_, new_n6890_, new_n6891_,
    new_n6892_, new_n6893_, new_n6894_, new_n6895_, new_n6896_, new_n6897_,
    new_n6898_, new_n6899_, new_n6900_, new_n6901_, new_n6902_, new_n6903_,
    new_n6904_, new_n6905_, new_n6906_, new_n6907_, new_n6908_, new_n6909_,
    new_n6910_, new_n6911_, new_n6912_, new_n6913_, new_n6914_, new_n6915_,
    new_n6916_, new_n6917_, new_n6918_, new_n6919_, new_n6920_, new_n6921_,
    new_n6922_, new_n6923_, new_n6924_, new_n6925_, new_n6926_, new_n6927_,
    new_n6928_, new_n6929_, new_n6930_, new_n6931_, new_n6932_, new_n6933_,
    new_n6934_, new_n6935_, new_n6936_, new_n6937_, new_n6938_, new_n6939_,
    new_n6940_, new_n6941_, new_n6942_, new_n6943_, new_n6944_, new_n6945_,
    new_n6946_, new_n6947_, new_n6948_, new_n6949_, new_n6950_, new_n6951_,
    new_n6952_, new_n6953_, new_n6954_, new_n6955_, new_n6956_, new_n6957_,
    new_n6958_, new_n6959_, new_n6960_, new_n6961_, new_n6962_, new_n6963_,
    new_n6964_, new_n6965_, new_n6966_, new_n6967_, new_n6968_, new_n6969_,
    new_n6970_, new_n6971_, new_n6972_, new_n6973_, new_n6974_, new_n6975_,
    new_n6976_, new_n6977_, new_n6978_, new_n6979_, new_n6980_, new_n6981_,
    new_n6982_, new_n6983_, new_n6984_, new_n6985_, new_n6986_, new_n6987_,
    new_n6988_, new_n6989_, new_n6990_, new_n6991_, new_n6992_, new_n6993_,
    new_n6994_, new_n6995_, new_n6996_, new_n6997_, new_n6998_, new_n6999_,
    new_n7000_, new_n7001_, new_n7002_, new_n7003_, new_n7004_, new_n7005_,
    new_n7006_, new_n7007_, new_n7008_, new_n7009_, new_n7010_, new_n7011_,
    new_n7012_, new_n7013_, new_n7014_, new_n7015_, new_n7016_, new_n7017_,
    new_n7018_, new_n7019_, new_n7020_, new_n7021_, new_n7022_, new_n7023_,
    new_n7024_, new_n7025_, new_n7026_, new_n7027_, new_n7028_, new_n7029_,
    new_n7030_, new_n7031_, new_n7032_, new_n7033_, new_n7034_, new_n7035_,
    new_n7036_, new_n7037_, new_n7038_, new_n7039_, new_n7040_, new_n7041_,
    new_n7042_, new_n7043_, new_n7044_, new_n7045_, new_n7046_, new_n7047_,
    new_n7048_, new_n7049_, new_n7050_, new_n7051_, new_n7052_, new_n7053_,
    new_n7054_, new_n7055_, new_n7056_, new_n7057_, new_n7058_, new_n7059_,
    new_n7060_, new_n7061_, new_n7062_, new_n7063_, new_n7064_, new_n7065_,
    new_n7066_, new_n7067_, new_n7068_, new_n7069_, new_n7070_, new_n7071_,
    new_n7072_, new_n7073_, new_n7074_, new_n7075_, new_n7076_, new_n7077_,
    new_n7078_, new_n7079_, new_n7080_, new_n7081_, new_n7082_, new_n7083_,
    new_n7084_, new_n7085_, new_n7086_, new_n7087_, new_n7088_, new_n7089_,
    new_n7090_, new_n7091_, new_n7092_, new_n7093_, new_n7094_, new_n7095_,
    new_n7096_, new_n7097_, new_n7098_, new_n7099_, new_n7100_, new_n7101_,
    new_n7102_, new_n7103_, new_n7104_, new_n7105_, new_n7106_, new_n7107_,
    new_n7108_, new_n7109_, new_n7110_, new_n7111_, new_n7112_, new_n7113_,
    new_n7114_, new_n7115_, new_n7116_, new_n7117_, new_n7118_, new_n7119_,
    new_n7120_, new_n7121_, new_n7122_, new_n7123_, new_n7124_, new_n7125_,
    new_n7126_, new_n7127_, new_n7128_, new_n7129_, new_n7130_, new_n7131_,
    new_n7132_, new_n7133_, new_n7134_, new_n7135_, new_n7136_, new_n7137_,
    new_n7138_, new_n7139_, new_n7140_, new_n7141_, new_n7142_, new_n7143_,
    new_n7144_, new_n7145_, new_n7146_, new_n7147_, new_n7148_, new_n7149_,
    new_n7150_, new_n7151_, new_n7152_, new_n7153_, new_n7154_, new_n7155_,
    new_n7156_, new_n7157_, new_n7158_, new_n7159_, new_n7160_, new_n7161_,
    new_n7162_, new_n7163_, new_n7164_, new_n7165_, new_n7166_, new_n7167_,
    new_n7168_, new_n7169_, new_n7170_, new_n7171_, new_n7172_, new_n7173_,
    new_n7174_, new_n7175_, new_n7176_, new_n7177_, new_n7178_, new_n7179_,
    new_n7180_, new_n7181_, new_n7182_, new_n7183_, new_n7184_, new_n7185_,
    new_n7186_, new_n7187_, new_n7188_, new_n7189_, new_n7190_, new_n7191_,
    new_n7192_, new_n7193_, new_n7194_, new_n7195_, new_n7196_, new_n7197_,
    new_n7198_, new_n7199_, new_n7200_, new_n7201_, new_n7202_, new_n7203_,
    new_n7204_, new_n7205_, new_n7206_, new_n7207_, new_n7208_, new_n7209_,
    new_n7210_, new_n7211_, new_n7212_, new_n7213_, new_n7214_, new_n7215_,
    new_n7216_, new_n7217_, new_n7218_, new_n7219_, new_n7220_, new_n7221_,
    new_n7222_, new_n7223_, new_n7224_, new_n7225_, new_n7226_, new_n7227_,
    new_n7228_, new_n7229_, new_n7230_, new_n7231_, new_n7232_, new_n7233_,
    new_n7234_, new_n7235_, new_n7236_, new_n7237_, new_n7238_, new_n7239_,
    new_n7240_, new_n7241_, new_n7242_, new_n7243_, new_n7244_, new_n7245_,
    new_n7246_, new_n7247_, new_n7248_, new_n7249_, new_n7250_, new_n7251_,
    new_n7252_, new_n7253_, new_n7254_, new_n7255_, new_n7256_, new_n7257_,
    new_n7258_, new_n7259_, new_n7260_, new_n7261_, new_n7262_, new_n7263_,
    new_n7264_, new_n7265_, new_n7266_, new_n7267_, new_n7268_, new_n7269_,
    new_n7270_, new_n7271_, new_n7272_, new_n7273_, new_n7274_, new_n7275_,
    new_n7276_, new_n7277_, new_n7278_, new_n7279_, new_n7280_, new_n7281_,
    new_n7282_, new_n7283_, new_n7284_, new_n7285_, new_n7286_, new_n7287_,
    new_n7288_, new_n7289_, new_n7290_, new_n7291_, new_n7292_, new_n7293_,
    new_n7294_, new_n7295_, new_n7296_, new_n7297_, new_n7298_, new_n7299_,
    new_n7300_, new_n7301_, new_n7302_, new_n7303_, new_n7304_, new_n7305_,
    new_n7306_, new_n7307_, new_n7308_, new_n7309_, new_n7310_, new_n7311_,
    new_n7312_, new_n7313_, new_n7314_, new_n7315_, new_n7316_, new_n7317_,
    new_n7318_, new_n7319_, new_n7320_, new_n7321_, new_n7322_, new_n7323_,
    new_n7324_, new_n7325_, new_n7326_, new_n7327_, new_n7328_, new_n7329_,
    new_n7330_, new_n7331_, new_n7332_, new_n7333_, new_n7334_, new_n7335_,
    new_n7336_, new_n7337_, new_n7338_, new_n7339_, new_n7340_, new_n7341_,
    new_n7342_, new_n7343_, new_n7344_, new_n7345_, new_n7346_, new_n7347_,
    new_n7348_, new_n7349_, new_n7350_, new_n7351_, new_n7352_, new_n7353_,
    new_n7354_, new_n7355_, new_n7356_, new_n7357_, new_n7358_, new_n7359_,
    new_n7360_, new_n7361_, new_n7362_, new_n7363_, new_n7364_, new_n7365_,
    new_n7366_, new_n7367_, new_n7368_, new_n7369_, new_n7370_, new_n7371_,
    new_n7372_, new_n7373_, new_n7374_, new_n7375_, new_n7376_, new_n7377_,
    new_n7378_, new_n7379_, new_n7380_, new_n7381_, new_n7382_, new_n7383_,
    new_n7384_, new_n7385_, new_n7386_, new_n7387_, new_n7388_, new_n7389_,
    new_n7390_, new_n7391_, new_n7392_, new_n7393_, new_n7394_, new_n7395_,
    new_n7396_, new_n7397_, new_n7398_, new_n7399_, new_n7400_, new_n7401_,
    new_n7402_, new_n7403_, new_n7404_, new_n7405_, new_n7406_, new_n7407_,
    new_n7408_, new_n7409_, new_n7410_, new_n7411_, new_n7412_, new_n7413_,
    new_n7414_, new_n7415_, new_n7416_, new_n7417_, new_n7418_, new_n7419_,
    new_n7420_, new_n7421_, new_n7422_, new_n7423_, new_n7424_, new_n7425_,
    new_n7426_, new_n7427_, new_n7428_, new_n7429_, new_n7430_, new_n7431_,
    new_n7432_, new_n7433_, new_n7434_, new_n7435_, new_n7436_, new_n7437_,
    new_n7438_, new_n7439_, new_n7440_, new_n7441_, new_n7442_, new_n7443_,
    new_n7444_, new_n7445_, new_n7446_, new_n7447_, new_n7448_, new_n7449_,
    new_n7450_, new_n7451_, new_n7452_, new_n7453_, new_n7454_, new_n7455_,
    new_n7456_, new_n7457_, new_n7458_, new_n7459_, new_n7460_, new_n7461_,
    new_n7462_, new_n7463_, new_n7464_, new_n7465_, new_n7466_, new_n7467_,
    new_n7468_, new_n7469_, new_n7470_, new_n7471_, new_n7472_, new_n7473_,
    new_n7474_, new_n7475_, new_n7476_, new_n7477_, new_n7478_, new_n7479_,
    new_n7480_, new_n7481_, new_n7482_, new_n7483_, new_n7484_, new_n7485_,
    new_n7486_, new_n7487_, new_n7488_, new_n7489_, new_n7490_, new_n7491_,
    new_n7492_, new_n7493_, new_n7494_, new_n7495_, new_n7496_, new_n7497_,
    new_n7498_, new_n7499_, new_n7500_, new_n7501_, new_n7502_, new_n7503_,
    new_n7504_, new_n7505_, new_n7506_, new_n7507_, new_n7508_, new_n7509_,
    new_n7510_, new_n7511_, new_n7512_, new_n7513_, new_n7514_, new_n7515_,
    new_n7516_, new_n7517_, new_n7518_, new_n7519_, new_n7520_, new_n7521_,
    new_n7522_, new_n7523_, new_n7524_, new_n7525_, new_n7526_, new_n7527_,
    new_n7528_, new_n7529_, new_n7530_, new_n7531_, new_n7532_, new_n7533_,
    new_n7534_, new_n7535_, new_n7536_, new_n7537_, new_n7538_, new_n7539_,
    new_n7540_, new_n7541_, new_n7542_, new_n7543_, new_n7544_, new_n7545_,
    new_n7546_, new_n7547_, new_n7548_, new_n7549_, new_n7550_, new_n7551_,
    new_n7552_, new_n7553_, new_n7554_, new_n7555_, new_n7556_, new_n7557_,
    new_n7558_, new_n7559_, new_n7560_, new_n7561_, new_n7562_, new_n7563_,
    new_n7564_, new_n7565_, new_n7566_, new_n7567_, new_n7568_, new_n7569_,
    new_n7570_, new_n7571_, new_n7572_, new_n7573_, new_n7574_, new_n7575_,
    new_n7576_, new_n7577_, new_n7578_, new_n7579_, new_n7580_, new_n7581_,
    new_n7582_, new_n7583_, new_n7584_, new_n7585_, new_n7586_, new_n7587_,
    new_n7588_, new_n7589_, new_n7590_, new_n7591_, new_n7592_, new_n7593_,
    new_n7594_, new_n7595_, new_n7596_, new_n7597_, new_n7598_, new_n7599_,
    new_n7600_, new_n7601_, new_n7602_, new_n7603_, new_n7604_, new_n7605_,
    new_n7606_, new_n7607_, new_n7608_, new_n7609_, new_n7610_, new_n7611_,
    new_n7612_, new_n7613_, new_n7614_, new_n7615_, new_n7616_, new_n7617_,
    new_n7618_, new_n7619_, new_n7620_, new_n7621_, new_n7622_, new_n7623_,
    new_n7624_, new_n7625_, new_n7626_, new_n7627_, new_n7628_, new_n7629_,
    new_n7630_, new_n7631_, new_n7632_, new_n7633_, new_n7634_, new_n7635_,
    new_n7636_, new_n7637_, new_n7638_, new_n7639_, new_n7640_, new_n7641_,
    new_n7642_, new_n7643_, new_n7644_, new_n7645_, new_n7646_, new_n7647_,
    new_n7648_, new_n7649_, new_n7650_, new_n7651_, new_n7652_, new_n7653_,
    new_n7654_, new_n7655_, new_n7656_, new_n7657_, new_n7658_, new_n7659_,
    new_n7660_, new_n7661_, new_n7662_, new_n7663_, new_n7664_, new_n7665_,
    new_n7666_, new_n7667_, new_n7668_, new_n7669_, new_n7670_, new_n7671_,
    new_n7672_, new_n7673_, new_n7674_, new_n7675_, new_n7676_, new_n7677_,
    new_n7678_, new_n7679_, new_n7680_, new_n7681_, new_n7682_, new_n7683_,
    new_n7684_, new_n7685_, new_n7686_, new_n7687_, new_n7688_, new_n7689_,
    new_n7690_, new_n7691_, new_n7692_, new_n7693_, new_n7694_, new_n7695_,
    new_n7696_, new_n7697_, new_n7698_, new_n7699_, new_n7700_, new_n7701_,
    new_n7702_, new_n7703_, new_n7704_, new_n7705_, new_n7706_, new_n7707_,
    new_n7708_, new_n7709_, new_n7710_, new_n7711_, new_n7712_, new_n7713_,
    new_n7714_, new_n7715_, new_n7716_, new_n7717_, new_n7718_, new_n7719_,
    new_n7720_, new_n7721_, new_n7722_, new_n7723_, new_n7724_, new_n7725_,
    new_n7726_, new_n7727_, new_n7728_, new_n7729_, new_n7730_, new_n7731_,
    new_n7732_, new_n7733_, new_n7734_, new_n7735_, new_n7736_, new_n7737_,
    new_n7738_, new_n7739_, new_n7740_, new_n7741_, new_n7742_, new_n7743_,
    new_n7744_, new_n7745_, new_n7746_, new_n7747_, new_n7748_, new_n7749_,
    new_n7750_, new_n7751_, new_n7752_, new_n7753_, new_n7754_, new_n7755_,
    new_n7756_, new_n7757_, new_n7758_, new_n7759_, new_n7760_, new_n7761_,
    new_n7762_, new_n7763_, new_n7764_, new_n7765_, new_n7766_, new_n7767_,
    new_n7768_, new_n7769_, new_n7770_, new_n7771_, new_n7772_, new_n7773_,
    new_n7774_, new_n7775_, new_n7776_, new_n7777_, new_n7778_, new_n7779_,
    new_n7780_, new_n7781_, new_n7782_, new_n7783_, new_n7784_, new_n7785_,
    new_n7786_, new_n7787_, new_n7788_, new_n7789_, new_n7790_, new_n7791_,
    new_n7792_, new_n7793_, new_n7794_, new_n7795_, new_n7796_, new_n7797_,
    new_n7798_, new_n7799_, new_n7800_, new_n7801_, new_n7802_, new_n7803_,
    new_n7804_, new_n7805_, new_n7806_, new_n7807_, new_n7808_, new_n7809_,
    new_n7810_, new_n7811_, new_n7812_, new_n7813_, new_n7814_, new_n7815_,
    new_n7816_, new_n7817_, new_n7818_, new_n7819_, new_n7820_, new_n7821_,
    new_n7822_, new_n7823_, new_n7824_, new_n7825_, new_n7826_, new_n7827_,
    new_n7828_, new_n7829_, new_n7830_, new_n7831_, new_n7832_, new_n7833_,
    new_n7834_, new_n7835_, new_n7836_, new_n7837_, new_n7838_, new_n7839_,
    new_n7840_, new_n7841_, new_n7842_, new_n7843_, new_n7844_, new_n7845_,
    new_n7846_, new_n7847_, new_n7848_, new_n7849_, new_n7850_, new_n7851_,
    new_n7852_, new_n7853_, new_n7854_, new_n7855_, new_n7856_, new_n7857_,
    new_n7858_, new_n7859_, new_n7860_, new_n7861_, new_n7862_, new_n7863_,
    new_n7864_, new_n7865_, new_n7866_, new_n7867_, new_n7868_, new_n7869_,
    new_n7870_, new_n7871_, new_n7872_, new_n7873_, new_n7874_, new_n7875_,
    new_n7876_, new_n7877_, new_n7878_, new_n7879_, new_n7880_, new_n7881_,
    new_n7882_, new_n7883_, new_n7884_, new_n7885_, new_n7886_, new_n7887_,
    new_n7888_, new_n7889_, new_n7890_, new_n7891_, new_n7892_, new_n7893_,
    new_n7894_, new_n7895_, new_n7896_, new_n7897_, new_n7898_, new_n7899_,
    new_n7900_, new_n7901_, new_n7902_, new_n7903_, new_n7904_, new_n7905_,
    new_n7906_, new_n7907_, new_n7908_, new_n7909_, new_n7910_, new_n7911_,
    new_n7912_, new_n7913_, new_n7914_, new_n7915_, new_n7916_, new_n7917_,
    new_n7918_, new_n7919_, new_n7920_, new_n7921_, new_n7922_, new_n7923_,
    new_n7924_, new_n7925_, new_n7926_, new_n7927_, new_n7928_, new_n7929_,
    new_n7930_, new_n7931_, new_n7932_, new_n7933_, new_n7934_, new_n7935_,
    new_n7936_, new_n7937_, new_n7938_, new_n7939_, new_n7940_, new_n7941_,
    new_n7942_, new_n7943_, new_n7944_, new_n7945_, new_n7946_, new_n7947_,
    new_n7948_, new_n7949_, new_n7950_, new_n7951_, new_n7952_, new_n7953_,
    new_n7954_, new_n7955_, new_n7956_, new_n7957_, new_n7958_, new_n7959_,
    new_n7960_, new_n7961_, new_n7962_, new_n7963_, new_n7964_, new_n7965_,
    new_n7966_, new_n7967_, new_n7968_, new_n7969_, new_n7970_, new_n7971_,
    new_n7972_, new_n7973_, new_n7974_, new_n7975_, new_n7976_, new_n7977_,
    new_n7978_, new_n7979_, new_n7980_, new_n7981_, new_n7982_, new_n7983_,
    new_n7984_, new_n7985_, new_n7986_, new_n7987_, new_n7988_, new_n7989_,
    new_n7990_, new_n7991_, new_n7992_, new_n7993_, new_n7994_, new_n7995_,
    new_n7996_, new_n7997_, new_n7998_, new_n7999_, new_n8000_, new_n8001_,
    new_n8002_, new_n8003_, new_n8004_, new_n8005_, new_n8006_, new_n8007_,
    new_n8008_, new_n8009_, new_n8010_, new_n8011_, new_n8012_, new_n8013_,
    new_n8014_, new_n8015_, new_n8016_, new_n8017_, new_n8018_, new_n8019_,
    new_n8020_, new_n8021_, new_n8022_, new_n8023_, new_n8024_, new_n8025_,
    new_n8026_, new_n8027_, new_n8028_, new_n8029_, new_n8030_, new_n8031_,
    new_n8032_, new_n8033_, new_n8034_, new_n8035_, new_n8036_, new_n8037_,
    new_n8038_, new_n8039_, new_n8040_, new_n8041_, new_n8042_, new_n8043_,
    new_n8044_, new_n8045_, new_n8046_, new_n8047_, new_n8048_, new_n8049_,
    new_n8050_, new_n8051_, new_n8052_, new_n8053_, new_n8054_, new_n8055_,
    new_n8056_, new_n8057_, new_n8058_, new_n8059_, new_n8060_, new_n8061_,
    new_n8062_, new_n8063_, new_n8064_, new_n8065_, new_n8066_, new_n8067_,
    new_n8068_, new_n8069_, new_n8070_, new_n8071_, new_n8072_, new_n8073_,
    new_n8074_, new_n8075_, new_n8076_, new_n8077_, new_n8078_, new_n8079_,
    new_n8080_, new_n8081_, new_n8082_, new_n8083_, new_n8084_, new_n8085_,
    new_n8086_, new_n8087_, new_n8088_, new_n8089_, new_n8090_, new_n8091_,
    new_n8092_, new_n8093_, new_n8094_, new_n8095_, new_n8096_, new_n8097_,
    new_n8098_, new_n8099_, new_n8100_, new_n8101_, new_n8102_, new_n8103_,
    new_n8104_, new_n8105_, new_n8106_, new_n8107_, new_n8108_, new_n8109_,
    new_n8110_, new_n8111_, new_n8112_, new_n8113_, new_n8114_, new_n8115_,
    new_n8116_, new_n8117_, new_n8118_, new_n8119_, new_n8120_, new_n8121_,
    new_n8122_, new_n8123_, new_n8124_, new_n8125_, new_n8126_, new_n8127_,
    new_n8128_, new_n8129_, new_n8130_, new_n8131_, new_n8132_, new_n8133_,
    new_n8134_, new_n8135_, new_n8136_, new_n8137_, new_n8138_, new_n8139_,
    new_n8140_, new_n8141_, new_n8142_, new_n8143_, new_n8144_, new_n8145_,
    new_n8146_, new_n8147_, new_n8148_, new_n8149_, new_n8150_, new_n8151_,
    new_n8152_, new_n8153_, new_n8154_, new_n8155_, new_n8156_, new_n8157_,
    new_n8158_, new_n8159_, new_n8160_, new_n8161_, new_n8162_, new_n8163_,
    new_n8164_, new_n8165_, new_n8166_, new_n8167_, new_n8168_, new_n8169_,
    new_n8170_, new_n8171_, new_n8172_, new_n8173_, new_n8174_, new_n8175_,
    new_n8176_, new_n8177_, new_n8178_, new_n8179_, new_n8180_, new_n8181_,
    new_n8182_, new_n8183_, new_n8184_, new_n8185_, new_n8186_, new_n8187_,
    new_n8188_, new_n8189_, new_n8190_, new_n8191_, new_n8192_, new_n8193_,
    new_n8194_, new_n8195_, new_n8196_, new_n8197_, new_n8198_, new_n8199_,
    new_n8200_, new_n8201_, new_n8202_, new_n8203_, new_n8204_, new_n8205_,
    new_n8206_, new_n8207_, new_n8208_, new_n8209_, new_n8210_, new_n8211_,
    new_n8212_, new_n8213_, new_n8214_, new_n8215_, new_n8216_, new_n8217_,
    new_n8218_, new_n8219_, new_n8220_, new_n8221_, new_n8222_, new_n8223_,
    new_n8224_, new_n8225_, new_n8226_, new_n8227_, new_n8228_, new_n8229_,
    new_n8230_, new_n8231_, new_n8232_, new_n8233_, new_n8234_, new_n8235_,
    new_n8236_, new_n8237_, new_n8238_, new_n8239_, new_n8240_, new_n8241_,
    new_n8242_, new_n8243_, new_n8244_, new_n8245_, new_n8246_, new_n8247_,
    new_n8248_, new_n8249_, new_n8250_, new_n8251_, new_n8252_, new_n8253_,
    new_n8254_, new_n8255_, new_n8256_, new_n8257_, new_n8258_, new_n8259_,
    new_n8260_, new_n8261_, new_n8262_, new_n8263_, new_n8264_, new_n8265_,
    new_n8266_, new_n8267_, new_n8268_, new_n8269_, new_n8270_, new_n8271_,
    new_n8272_, new_n8273_, new_n8274_, new_n8275_, new_n8276_, new_n8277_,
    new_n8278_, new_n8279_, new_n8280_, new_n8281_, new_n8282_, new_n8283_,
    new_n8284_, new_n8285_, new_n8286_, new_n8287_, new_n8288_, new_n8289_,
    new_n8290_, new_n8291_, new_n8292_, new_n8293_, new_n8294_, new_n8295_,
    new_n8296_, new_n8297_, new_n8298_, new_n8299_, new_n8300_, new_n8301_,
    new_n8302_, new_n8303_, new_n8304_, new_n8305_, new_n8306_, new_n8307_,
    new_n8308_, new_n8309_, new_n8310_, new_n8311_, new_n8312_, new_n8313_,
    new_n8314_, new_n8315_, new_n8316_, new_n8317_, new_n8318_, new_n8319_,
    new_n8320_, new_n8321_, new_n8322_, new_n8323_, new_n8324_, new_n8325_,
    new_n8326_, new_n8327_, new_n8328_, new_n8329_, new_n8330_, new_n8331_,
    new_n8332_, new_n8333_, new_n8334_, new_n8335_, new_n8336_, new_n8337_,
    new_n8338_, new_n8339_, new_n8340_, new_n8341_, new_n8342_, new_n8343_,
    new_n8344_, new_n8345_, new_n8346_, new_n8347_, new_n8348_, new_n8349_,
    new_n8350_, new_n8351_, new_n8352_, new_n8353_, new_n8354_, new_n8355_,
    new_n8356_, new_n8357_, new_n8358_, new_n8359_, new_n8360_, new_n8361_,
    new_n8362_, new_n8363_, new_n8364_, new_n8365_, new_n8366_, new_n8367_,
    new_n8368_, new_n8369_, new_n8370_, new_n8371_, new_n8372_, new_n8373_,
    new_n8374_, new_n8375_, new_n8376_, new_n8377_, new_n8378_, new_n8379_,
    new_n8380_, new_n8381_, new_n8382_, new_n8383_, new_n8384_, new_n8385_,
    new_n8386_, new_n8387_, new_n8388_, new_n8389_, new_n8390_, new_n8391_,
    new_n8392_, new_n8393_, new_n8394_, new_n8395_, new_n8396_, new_n8397_,
    new_n8398_, new_n8399_, new_n8400_, new_n8401_, new_n8402_, new_n8403_,
    new_n8404_, new_n8405_, new_n8406_, new_n8407_, new_n8408_, new_n8409_,
    new_n8410_, new_n8411_, new_n8412_, new_n8413_, new_n8414_, new_n8415_,
    new_n8416_, new_n8417_, new_n8418_, new_n8419_, new_n8420_, new_n8421_,
    new_n8422_, new_n8423_, new_n8424_, new_n8425_, new_n8426_, new_n8427_,
    new_n8428_, new_n8429_, new_n8430_, new_n8431_, new_n8432_, new_n8433_,
    new_n8434_, new_n8435_, new_n8436_, new_n8437_, new_n8438_, new_n8439_,
    new_n8440_, new_n8441_, new_n8442_, new_n8443_, new_n8444_, new_n8445_,
    new_n8446_, new_n8447_, new_n8448_, new_n8449_, new_n8450_, new_n8451_,
    new_n8452_, new_n8453_, new_n8454_, new_n8455_, new_n8456_, new_n8457_,
    new_n8458_, new_n8459_, new_n8460_, new_n8461_, new_n8462_, new_n8463_,
    new_n8464_, new_n8465_, new_n8466_, new_n8467_, new_n8468_, new_n8469_,
    new_n8470_, new_n8471_, new_n8472_, new_n8473_, new_n8474_, new_n8475_,
    new_n8476_, new_n8477_, new_n8478_, new_n8479_, new_n8480_, new_n8481_,
    new_n8482_, new_n8483_, new_n8484_, new_n8485_, new_n8486_, new_n8487_,
    new_n8488_, new_n8489_, new_n8490_, new_n8491_, new_n8492_, new_n8493_,
    new_n8494_, new_n8495_, new_n8496_, new_n8497_, new_n8498_, new_n8499_,
    new_n8500_, new_n8501_, new_n8502_, new_n8503_, new_n8504_, new_n8505_,
    new_n8506_, new_n8507_, new_n8508_, new_n8509_, new_n8510_, new_n8511_,
    new_n8512_, new_n8513_, new_n8514_, new_n8515_, new_n8516_, new_n8517_,
    new_n8518_, new_n8519_, new_n8520_, new_n8521_, new_n8522_, new_n8523_,
    new_n8524_, new_n8525_, new_n8526_, new_n8527_, new_n8528_, new_n8529_,
    new_n8530_, new_n8531_, new_n8532_, new_n8533_, new_n8534_, new_n8535_,
    new_n8536_, new_n8537_, new_n8538_, new_n8539_, new_n8540_, new_n8541_,
    new_n8542_, new_n8543_, new_n8544_, new_n8545_, new_n8546_, new_n8547_,
    new_n8548_, new_n8549_, new_n8550_, new_n8551_, new_n8552_, new_n8553_,
    new_n8554_, new_n8555_, new_n8556_, new_n8557_, new_n8558_, new_n8559_,
    new_n8560_, new_n8561_, new_n8562_, new_n8563_, new_n8564_, new_n8565_,
    new_n8566_, new_n8567_, new_n8568_, new_n8569_, new_n8570_, new_n8571_,
    new_n8572_, new_n8573_, new_n8574_, new_n8575_, new_n8576_, new_n8577_,
    new_n8578_, new_n8579_, new_n8580_, new_n8581_, new_n8582_, new_n8583_,
    new_n8584_, new_n8585_, new_n8586_, new_n8587_, new_n8588_, new_n8589_,
    new_n8590_, new_n8591_, new_n8592_, new_n8593_, new_n8594_, new_n8595_,
    new_n8596_, new_n8597_, new_n8598_, new_n8599_, new_n8600_, new_n8601_,
    new_n8602_, new_n8603_, new_n8604_, new_n8605_, new_n8606_, new_n8607_,
    new_n8608_, new_n8609_, new_n8610_, new_n8611_, new_n8612_, new_n8613_,
    new_n8614_, new_n8615_, new_n8616_, new_n8617_, new_n8618_, new_n8619_,
    new_n8620_, new_n8621_, new_n8622_, new_n8623_, new_n8624_, new_n8625_,
    new_n8626_, new_n8627_, new_n8628_, new_n8629_, new_n8630_, new_n8631_,
    new_n8632_, new_n8633_, new_n8634_, new_n8635_, new_n8636_, new_n8637_,
    new_n8638_, new_n8639_, new_n8640_, new_n8641_, new_n8642_, new_n8643_,
    new_n8644_, new_n8645_, new_n8646_, new_n8647_, new_n8648_, new_n8649_,
    new_n8650_, new_n8651_, new_n8652_, new_n8653_, new_n8654_, new_n8655_,
    new_n8656_, new_n8657_, new_n8658_, new_n8659_, new_n8660_, new_n8661_,
    new_n8662_, new_n8663_, new_n8664_, new_n8665_, new_n8666_, new_n8667_,
    new_n8668_, new_n8669_, new_n8670_, new_n8671_, new_n8672_, new_n8673_,
    new_n8674_, new_n8675_, new_n8676_, new_n8677_, new_n8678_, new_n8679_,
    new_n8680_, new_n8681_, new_n8682_, new_n8683_, new_n8684_, new_n8685_,
    new_n8686_, new_n8687_, new_n8688_, new_n8689_, new_n8690_, new_n8691_,
    new_n8692_, new_n8693_, new_n8694_, new_n8695_, new_n8696_, new_n8697_,
    new_n8698_, new_n8699_, new_n8700_, new_n8701_, new_n8702_, new_n8703_,
    new_n8704_, new_n8705_, new_n8706_, new_n8707_, new_n8708_, new_n8709_,
    new_n8710_, new_n8711_, new_n8712_, new_n8713_, new_n8714_, new_n8715_,
    new_n8716_, new_n8717_, new_n8718_, new_n8719_, new_n8720_, new_n8721_,
    new_n8722_, new_n8723_, new_n8724_, new_n8725_, new_n8726_, new_n8727_,
    new_n8728_, new_n8729_, new_n8730_, new_n8731_, new_n8732_, new_n8733_,
    new_n8734_, new_n8735_, new_n8736_, new_n8737_, new_n8738_, new_n8739_,
    new_n8740_, new_n8741_, new_n8742_, new_n8743_, new_n8744_, new_n8745_,
    new_n8746_, new_n8747_, new_n8748_, new_n8749_, new_n8750_, new_n8751_,
    new_n8752_, new_n8753_, new_n8754_, new_n8755_, new_n8756_, new_n8757_,
    new_n8758_, new_n8759_, new_n8760_, new_n8761_, new_n8762_, new_n8763_,
    new_n8764_, new_n8765_, new_n8766_, new_n8767_, new_n8768_, new_n8769_,
    new_n8770_, new_n8771_, new_n8772_, new_n8773_, new_n8774_, new_n8775_,
    new_n8776_, new_n8777_, new_n8778_, new_n8779_, new_n8780_, new_n8781_,
    new_n8782_, new_n8783_, new_n8784_, new_n8785_, new_n8786_, new_n8787_,
    new_n8788_, new_n8789_, new_n8790_, new_n8791_, new_n8792_, new_n8793_,
    new_n8794_, new_n8795_, new_n8796_, new_n8797_, new_n8798_, new_n8799_,
    new_n8800_, new_n8801_, new_n8802_, new_n8803_, new_n8804_, new_n8805_,
    new_n8806_, new_n8807_, new_n8808_, new_n8809_, new_n8810_, new_n8811_,
    new_n8812_, new_n8813_, new_n8814_, new_n8815_, new_n8816_, new_n8817_,
    new_n8818_, new_n8819_, new_n8820_, new_n8821_, new_n8822_, new_n8823_,
    new_n8824_, new_n8825_, new_n8826_, new_n8827_, new_n8828_, new_n8829_,
    new_n8830_, new_n8831_, new_n8832_, new_n8833_, new_n8834_, new_n8835_,
    new_n8836_, new_n8837_, new_n8838_, new_n8839_, new_n8840_, new_n8841_,
    new_n8842_, new_n8843_, new_n8844_, new_n8845_, new_n8846_, new_n8847_,
    new_n8848_, new_n8849_, new_n8850_, new_n8851_, new_n8852_, new_n8853_,
    new_n8854_, new_n8855_, new_n8856_, new_n8857_, new_n8858_, new_n8859_,
    new_n8860_, new_n8861_, new_n8862_, new_n8863_, new_n8864_, new_n8865_,
    new_n8866_, new_n8867_, new_n8868_, new_n8869_, new_n8870_, new_n8871_,
    new_n8872_, new_n8873_, new_n8874_, new_n8875_, new_n8876_, new_n8877_,
    new_n8878_, new_n8879_, new_n8880_, new_n8881_, new_n8882_, new_n8883_,
    new_n8884_, new_n8885_, new_n8886_, new_n8887_, new_n8888_, new_n8889_,
    new_n8890_, new_n8891_, new_n8892_, new_n8893_, new_n8894_, new_n8895_,
    new_n8896_, new_n8897_, new_n8898_, new_n8899_, new_n8900_, new_n8901_,
    new_n8902_, new_n8903_, new_n8904_, new_n8905_, new_n8906_, new_n8907_,
    new_n8908_, new_n8909_, new_n8910_, new_n8911_, new_n8912_, new_n8913_,
    new_n8914_, new_n8915_, new_n8916_, new_n8917_, new_n8918_, new_n8919_,
    new_n8920_, new_n8921_, new_n8922_, new_n8923_, new_n8924_, new_n8925_,
    new_n8926_, new_n8927_, new_n8928_, new_n8929_, new_n8930_, new_n8931_,
    new_n8932_, new_n8933_, new_n8934_, new_n8935_, new_n8936_, new_n8937_,
    new_n8938_, new_n8939_, new_n8940_, new_n8941_, new_n8942_, new_n8943_,
    new_n8944_, new_n8945_, new_n8946_, new_n8947_, new_n8948_, new_n8949_,
    new_n8950_, new_n8951_, new_n8952_, new_n8953_, new_n8954_, new_n8955_,
    new_n8956_, new_n8957_, new_n8958_, new_n8959_, new_n8960_, new_n8961_,
    new_n8962_, new_n8963_, new_n8964_, new_n8965_, new_n8966_, new_n8967_,
    new_n8968_, new_n8969_, new_n8970_, new_n8971_, new_n8972_, new_n8973_,
    new_n8974_, new_n8975_, new_n8976_, new_n8977_, new_n8978_, new_n8979_,
    new_n8980_, new_n8981_, new_n8982_, new_n8983_, new_n8984_, new_n8985_,
    new_n8986_, new_n8987_, new_n8988_, new_n8989_, new_n8990_, new_n8991_,
    new_n8992_, new_n8993_, new_n8994_, new_n8995_, new_n8996_, new_n8997_,
    new_n8998_, new_n8999_, new_n9000_, new_n9001_, new_n9002_, new_n9003_,
    new_n9004_, new_n9005_, new_n9006_, new_n9007_, new_n9008_, new_n9009_,
    new_n9010_, new_n9011_, new_n9012_, new_n9013_, new_n9014_, new_n9015_,
    new_n9016_, new_n9017_, new_n9018_, new_n9019_, new_n9020_, new_n9021_,
    new_n9022_, new_n9023_, new_n9024_, new_n9025_, new_n9026_, new_n9027_,
    new_n9028_, new_n9029_, new_n9030_, new_n9031_, new_n9032_, new_n9033_,
    new_n9034_, new_n9035_, new_n9036_, new_n9037_, new_n9038_, new_n9039_,
    new_n9040_, new_n9041_, new_n9042_, new_n9043_, new_n9044_, new_n9045_,
    new_n9046_, new_n9047_, new_n9048_, new_n9049_, new_n9050_, new_n9051_,
    new_n9052_, new_n9053_, new_n9054_, new_n9055_, new_n9056_, new_n9057_,
    new_n9058_, new_n9059_, new_n9060_, new_n9061_, new_n9062_, new_n9063_,
    new_n9064_, new_n9065_, new_n9066_, new_n9067_, new_n9068_, new_n9069_,
    new_n9070_, new_n9071_, new_n9072_, new_n9073_, new_n9074_, new_n9075_,
    new_n9076_, new_n9077_, new_n9078_, new_n9079_, new_n9080_, new_n9081_,
    new_n9082_, new_n9083_, new_n9084_, new_n9085_, new_n9086_, new_n9087_,
    new_n9088_, new_n9089_, new_n9090_, new_n9091_, new_n9092_, new_n9093_,
    new_n9094_, new_n9095_, new_n9096_, new_n9097_, new_n9098_, new_n9099_,
    new_n9100_, new_n9101_, new_n9102_, new_n9103_, new_n9104_, new_n9105_,
    new_n9106_, new_n9107_, new_n9108_, new_n9109_, new_n9110_, new_n9111_,
    new_n9112_, new_n9113_, new_n9114_, new_n9115_, new_n9116_, new_n9117_,
    new_n9118_, new_n9119_, new_n9120_, new_n9121_, new_n9122_, new_n9123_,
    new_n9124_, new_n9125_, new_n9126_, new_n9127_, new_n9128_, new_n9129_,
    new_n9130_, new_n9131_, new_n9132_, new_n9133_, new_n9134_, new_n9135_,
    new_n9136_, new_n9137_, new_n9138_, new_n9139_, new_n9140_, new_n9141_,
    new_n9142_, new_n9143_, new_n9144_, new_n9145_, new_n9146_, new_n9147_,
    new_n9148_, new_n9149_, new_n9150_, new_n9151_, new_n9152_, new_n9153_,
    new_n9154_, new_n9155_, new_n9156_, new_n9157_, new_n9158_, new_n9159_,
    new_n9160_, new_n9161_, new_n9162_, new_n9163_, new_n9164_, new_n9165_,
    new_n9166_, new_n9167_, new_n9168_, new_n9169_, new_n9170_, new_n9171_,
    new_n9172_, new_n9173_, new_n9174_, new_n9175_, new_n9176_, new_n9177_,
    new_n9178_, new_n9179_, new_n9180_, new_n9181_, new_n9182_, new_n9183_,
    new_n9184_, new_n9185_, new_n9186_, new_n9187_, new_n9188_, new_n9189_,
    new_n9190_, new_n9191_, new_n9192_, new_n9193_, new_n9194_, new_n9195_,
    new_n9196_, new_n9197_, new_n9198_, new_n9199_, new_n9200_, new_n9201_,
    new_n9202_, new_n9203_, new_n9204_, new_n9205_, new_n9206_, new_n9207_,
    new_n9208_, new_n9209_, new_n9210_, new_n9211_, new_n9212_, new_n9213_,
    new_n9214_, new_n9215_, new_n9216_, new_n9217_, new_n9218_, new_n9219_,
    new_n9220_, new_n9221_, new_n9222_, new_n9223_, new_n9224_, new_n9225_,
    new_n9226_, new_n9227_, new_n9228_, new_n9229_, new_n9230_, new_n9231_,
    new_n9232_, new_n9233_, new_n9234_, new_n9235_, new_n9236_, new_n9237_,
    new_n9238_, new_n9239_, new_n9240_, new_n9241_, new_n9242_, new_n9243_,
    new_n9244_, new_n9245_, new_n9246_, new_n9247_, new_n9248_, new_n9249_,
    new_n9250_, new_n9251_, new_n9252_, new_n9253_, new_n9254_, new_n9255_,
    new_n9256_, new_n9257_, new_n9258_, new_n9259_, new_n9260_, new_n9261_,
    new_n9262_, new_n9263_, new_n9264_, new_n9265_, new_n9266_, new_n9267_,
    new_n9268_, new_n9269_, new_n9270_, new_n9271_, new_n9272_, new_n9273_,
    new_n9274_, new_n9275_, new_n9276_, new_n9277_, new_n9278_, new_n9279_,
    new_n9280_, new_n9281_, new_n9282_, new_n9283_, new_n9284_, new_n9285_,
    new_n9286_, new_n9287_, new_n9288_, new_n9289_, new_n9290_, new_n9291_,
    new_n9292_, new_n9293_, new_n9294_, new_n9295_, new_n9296_, new_n9297_,
    new_n9298_, new_n9299_, new_n9300_, new_n9301_, new_n9302_, new_n9303_,
    new_n9304_, new_n9305_, new_n9306_, new_n9307_, new_n9308_, new_n9309_,
    new_n9310_, new_n9311_, new_n9312_, new_n9313_, new_n9314_, new_n9315_,
    new_n9316_, new_n9317_, new_n9318_, new_n9319_, new_n9320_, new_n9321_,
    new_n9322_, new_n9323_, new_n9324_, new_n9325_, new_n9326_, new_n9327_,
    new_n9328_, new_n9329_, new_n9330_, new_n9331_, new_n9332_, new_n9333_,
    new_n9334_, new_n9335_, new_n9336_, new_n9337_, new_n9338_, new_n9339_,
    new_n9340_, new_n9341_, new_n9342_, new_n9343_, new_n9344_, new_n9345_,
    new_n9346_, new_n9347_, new_n9348_, new_n9349_, new_n9350_, new_n9351_,
    new_n9352_, new_n9353_, new_n9354_, new_n9355_, new_n9356_, new_n9357_,
    new_n9358_, new_n9359_, new_n9360_, new_n9361_, new_n9362_, new_n9363_,
    new_n9364_, new_n9365_, new_n9366_, new_n9367_, new_n9368_, new_n9369_,
    new_n9370_, new_n9371_, new_n9372_, new_n9373_, new_n9374_, new_n9375_,
    new_n9376_, new_n9377_, new_n9378_, new_n9379_, new_n9380_, new_n9381_,
    new_n9382_, new_n9383_, new_n9384_, new_n9385_, new_n9386_, new_n9387_,
    new_n9388_, new_n9389_, new_n9390_, new_n9391_, new_n9392_, new_n9393_,
    new_n9394_, new_n9395_, new_n9396_, new_n9397_, new_n9398_, new_n9399_,
    new_n9400_, new_n9401_, new_n9402_, new_n9403_, new_n9404_, new_n9405_,
    new_n9406_, new_n9407_, new_n9408_, new_n9409_, new_n9410_, new_n9411_,
    new_n9412_, new_n9413_, new_n9414_, new_n9415_, new_n9416_, new_n9417_,
    new_n9418_, new_n9419_, new_n9420_, new_n9421_, new_n9422_, new_n9423_,
    new_n9424_, new_n9425_, new_n9426_, new_n9427_, new_n9428_, new_n9429_,
    new_n9430_, new_n9431_, new_n9432_, new_n9433_, new_n9434_, new_n9435_,
    new_n9436_, new_n9437_, new_n9438_, new_n9439_, new_n9440_, new_n9441_,
    new_n9442_, new_n9443_, new_n9444_, new_n9445_, new_n9446_, new_n9447_,
    new_n9448_, new_n9449_, new_n9450_, new_n9451_, new_n9452_, new_n9453_,
    new_n9454_, new_n9455_, new_n9456_, new_n9457_, new_n9458_, new_n9459_,
    new_n9460_, new_n9461_, new_n9462_, new_n9463_, new_n9464_, new_n9465_,
    new_n9466_, new_n9467_, new_n9468_, new_n9469_, new_n9470_, new_n9471_,
    new_n9472_, new_n9473_, new_n9474_, new_n9475_, new_n9476_, new_n9477_,
    new_n9478_, new_n9479_, new_n9480_, new_n9481_, new_n9482_, new_n9483_,
    new_n9484_, new_n9485_, new_n9486_, new_n9487_, new_n9488_, new_n9489_,
    new_n9490_, new_n9491_, new_n9492_, new_n9493_, new_n9494_, new_n9495_,
    new_n9496_, new_n9497_, new_n9498_, new_n9499_, new_n9500_, new_n9501_,
    new_n9502_, new_n9503_, new_n9504_, new_n9505_, new_n9506_, new_n9507_,
    new_n9508_, new_n9509_, new_n9510_, new_n9511_, new_n9512_, new_n9513_,
    new_n9514_, new_n9515_, new_n9516_, new_n9517_, new_n9518_, new_n9519_,
    new_n9520_, new_n9521_, new_n9522_, new_n9523_, new_n9524_, new_n9525_,
    new_n9526_, new_n9527_, new_n9528_, new_n9529_, new_n9530_, new_n9531_,
    new_n9532_, new_n9533_, new_n9534_, new_n9535_, new_n9536_, new_n9537_,
    new_n9538_, new_n9539_, new_n9540_, new_n9541_, new_n9542_, new_n9543_,
    new_n9544_, new_n9545_, new_n9546_, new_n9547_, new_n9548_, new_n9549_,
    new_n9550_, new_n9551_, new_n9552_, new_n9553_, new_n9554_, new_n9555_,
    new_n9556_, new_n9557_, new_n9558_, new_n9559_, new_n9560_, new_n9561_,
    new_n9562_, new_n9563_, new_n9564_, new_n9565_, new_n9566_, new_n9567_,
    new_n9568_, new_n9569_, new_n9570_, new_n9571_, new_n9572_, new_n9573_,
    new_n9574_, new_n9575_, new_n9576_, new_n9577_, new_n9578_, new_n9579_,
    new_n9580_, new_n9581_, new_n9582_, new_n9583_, new_n9584_, new_n9585_,
    new_n9586_, new_n9587_, new_n9588_, new_n9589_, new_n9590_, new_n9591_,
    new_n9592_, new_n9593_, new_n9594_, new_n9595_, new_n9596_, new_n9597_,
    new_n9598_, new_n9599_, new_n9600_, new_n9601_, new_n9602_, new_n9603_,
    new_n9604_, new_n9605_, new_n9606_, new_n9607_, new_n9608_, new_n9609_,
    new_n9610_, new_n9611_, new_n9612_, new_n9613_, new_n9614_, new_n9615_,
    new_n9616_, new_n9617_, new_n9618_, new_n9619_, new_n9620_, new_n9621_,
    new_n9622_, new_n9623_, new_n9624_, new_n9625_, new_n9626_, new_n9627_,
    new_n9628_, new_n9629_, new_n9630_, new_n9631_, new_n9632_, new_n9633_,
    new_n9634_, new_n9635_, new_n9636_, new_n9637_, new_n9638_, new_n9639_,
    new_n9640_, new_n9641_, new_n9642_, new_n9643_, new_n9644_, new_n9645_,
    new_n9646_, new_n9647_, new_n9648_, new_n9649_, new_n9650_, new_n9651_,
    new_n9652_, new_n9653_, new_n9654_, new_n9655_, new_n9656_, new_n9657_,
    new_n9658_, new_n9659_, new_n9660_, new_n9661_, new_n9662_, new_n9663_,
    new_n9664_, new_n9665_, new_n9666_, new_n9667_, new_n9668_, new_n9669_,
    new_n9670_, new_n9671_, new_n9672_, new_n9673_, new_n9674_, new_n9675_,
    new_n9676_, new_n9677_, new_n9678_, new_n9679_, new_n9680_, new_n9681_,
    new_n9682_, new_n9683_, new_n9684_, new_n9685_, new_n9686_, new_n9687_,
    new_n9688_, new_n9689_, new_n9690_, new_n9691_, new_n9692_, new_n9693_,
    new_n9694_, new_n9695_, new_n9696_, new_n9697_, new_n9698_, new_n9699_,
    new_n9700_, new_n9701_, new_n9702_, new_n9703_, new_n9704_, new_n9705_,
    new_n9706_, new_n9707_, new_n9708_, new_n9709_, new_n9710_, new_n9711_,
    new_n9712_, new_n9713_, new_n9714_, new_n9715_, new_n9716_, new_n9717_,
    new_n9718_, new_n9719_, new_n9720_, new_n9721_, new_n9722_, new_n9723_,
    new_n9724_, new_n9725_, new_n9726_, new_n9727_, new_n9728_, new_n9729_,
    new_n9730_, new_n9731_, new_n9732_, new_n9733_, new_n9734_, new_n9735_,
    new_n9736_, new_n9737_, new_n9738_, new_n9739_, new_n9740_, new_n9741_,
    new_n9742_, new_n9743_, new_n9744_, new_n9745_, new_n9746_, new_n9747_,
    new_n9748_, new_n9749_, new_n9750_, new_n9751_, new_n9752_, new_n9753_,
    new_n9754_, new_n9755_, new_n9756_, new_n9757_, new_n9758_, new_n9759_,
    new_n9760_, new_n9761_, new_n9762_, new_n9763_, new_n9764_, new_n9765_,
    new_n9766_, new_n9767_, new_n9768_, new_n9769_, new_n9770_, new_n9771_,
    new_n9772_, new_n9773_, new_n9774_, new_n9775_, new_n9776_, new_n9777_,
    new_n9778_, new_n9779_, new_n9780_, new_n9781_, new_n9782_, new_n9783_,
    new_n9784_, new_n9785_, new_n9786_, new_n9787_, new_n9788_, new_n9789_,
    new_n9790_, new_n9791_, new_n9792_, new_n9793_, new_n9794_, new_n9795_,
    new_n9796_, new_n9797_, new_n9798_, new_n9799_, new_n9800_, new_n9801_,
    new_n9802_, new_n9803_, new_n9804_, new_n9805_, new_n9806_, new_n9807_,
    new_n9808_, new_n9809_, new_n9810_, new_n9811_, new_n9812_, new_n9813_,
    new_n9814_, new_n9815_, new_n9816_, new_n9817_, new_n9818_, new_n9819_,
    new_n9820_, new_n9821_, new_n9822_, new_n9823_, new_n9824_, new_n9825_,
    new_n9826_, new_n9827_, new_n9828_, new_n9829_, new_n9830_, new_n9831_,
    new_n9832_, new_n9833_, new_n9834_, new_n9835_, new_n9836_, new_n9837_,
    new_n9838_, new_n9839_, new_n9840_, new_n9841_, new_n9842_, new_n9843_,
    new_n9844_, new_n9845_, new_n9846_, new_n9847_, new_n9848_, new_n9849_,
    new_n9850_, new_n9851_, new_n9852_, new_n9853_, new_n9854_, new_n9855_,
    new_n9856_, new_n9857_, new_n9858_, new_n9859_, new_n9860_, new_n9861_,
    new_n9862_, new_n9863_, new_n9864_, new_n9865_, new_n9866_, new_n9867_,
    new_n9868_, new_n9869_, new_n9870_, new_n9871_, new_n9872_, new_n9873_,
    new_n9874_, new_n9875_, new_n9876_, new_n9877_, new_n9878_, new_n9879_,
    new_n9880_, new_n9881_, new_n9882_, new_n9883_, new_n9884_, new_n9885_,
    new_n9886_, new_n9887_, new_n9888_, new_n9889_, new_n9890_, new_n9891_,
    new_n9892_, new_n9893_, new_n9894_, new_n9895_, new_n9896_, new_n9897_,
    new_n9898_, new_n9899_, new_n9900_, new_n9901_, new_n9902_, new_n9903_,
    new_n9904_, new_n9905_, new_n9906_, new_n9907_, new_n9908_, new_n9909_,
    new_n9910_, new_n9911_, new_n9912_, new_n9913_, new_n9914_, new_n9915_,
    new_n9916_, new_n9917_, new_n9918_, new_n9919_, new_n9920_, new_n9921_,
    new_n9922_, new_n9923_, new_n9924_, new_n9925_, new_n9926_, new_n9927_,
    new_n9928_, new_n9929_, new_n9930_, new_n9931_, new_n9932_, new_n9933_,
    new_n9934_, new_n9935_, new_n9936_, new_n9937_, new_n9938_, new_n9939_,
    new_n9940_, new_n9941_, new_n9942_, new_n9943_, new_n9944_, new_n9945_,
    new_n9946_, new_n9947_, new_n9948_, new_n9949_, new_n9950_, new_n9951_,
    new_n9952_, new_n9953_, new_n9954_, new_n9955_, new_n9956_, new_n9957_,
    new_n9958_, new_n9959_, new_n9960_, new_n9961_, new_n9962_, new_n9963_,
    new_n9964_, new_n9965_, new_n9966_, new_n9967_, new_n9968_, new_n9969_,
    new_n9970_, new_n9971_, new_n9972_, new_n9973_, new_n9974_, new_n9975_,
    new_n9976_, new_n9977_, new_n9978_, new_n9979_, new_n9980_, new_n9981_,
    new_n9982_, new_n9983_, new_n9984_, new_n9985_, new_n9986_, new_n9987_,
    new_n9988_, new_n9989_, new_n9990_, new_n9991_, new_n9992_, new_n9993_,
    new_n9994_, new_n9995_, new_n9996_, new_n9997_, new_n9998_, new_n9999_,
    new_n10000_, new_n10001_, new_n10002_, new_n10003_, new_n10004_,
    new_n10005_, new_n10006_, new_n10007_, new_n10008_, new_n10009_,
    new_n10010_, new_n10011_, new_n10012_, new_n10013_, new_n10014_,
    new_n10015_, new_n10016_, new_n10017_, new_n10018_, new_n10019_,
    new_n10020_, new_n10021_, new_n10022_, new_n10023_, new_n10024_,
    new_n10025_, new_n10026_, new_n10027_, new_n10028_, new_n10029_,
    new_n10030_, new_n10031_, new_n10032_, new_n10033_, new_n10034_,
    new_n10035_, new_n10036_, new_n10037_, new_n10038_, new_n10039_,
    new_n10040_, new_n10041_, new_n10042_, new_n10043_, new_n10044_,
    new_n10045_, new_n10046_, new_n10047_, new_n10048_, new_n10049_,
    new_n10050_, new_n10051_, new_n10052_, new_n10053_, new_n10054_,
    new_n10055_, new_n10056_, new_n10057_, new_n10058_, new_n10059_,
    new_n10060_, new_n10061_, new_n10062_, new_n10063_, new_n10064_,
    new_n10065_, new_n10066_, new_n10067_, new_n10068_, new_n10069_,
    new_n10070_, new_n10071_, new_n10072_, new_n10073_, new_n10074_,
    new_n10075_, new_n10076_, new_n10077_, new_n10078_, new_n10079_,
    new_n10080_, new_n10081_, new_n10082_, new_n10083_, new_n10084_,
    new_n10085_, new_n10086_, new_n10087_, new_n10088_, new_n10089_,
    new_n10090_, new_n10091_, new_n10092_, new_n10093_, new_n10094_,
    new_n10095_, new_n10096_, new_n10097_, new_n10098_, new_n10099_,
    new_n10100_, new_n10101_, new_n10102_, new_n10103_, new_n10104_,
    new_n10105_, new_n10106_, new_n10107_, new_n10108_, new_n10109_,
    new_n10110_, new_n10111_, new_n10112_, new_n10113_, new_n10114_,
    new_n10115_, new_n10116_, new_n10117_, new_n10118_, new_n10119_,
    new_n10120_, new_n10121_, new_n10122_, new_n10123_, new_n10124_,
    new_n10125_, new_n10126_, new_n10127_, new_n10128_, new_n10129_,
    new_n10130_, new_n10131_, new_n10132_, new_n10133_, new_n10134_,
    new_n10135_, new_n10136_, new_n10137_, new_n10138_, new_n10139_,
    new_n10140_, new_n10141_, new_n10142_, new_n10143_, new_n10144_,
    new_n10145_, new_n10146_, new_n10147_, new_n10148_, new_n10149_,
    new_n10150_, new_n10151_, new_n10152_, new_n10153_, new_n10154_,
    new_n10155_, new_n10156_, new_n10157_, new_n10158_, new_n10159_,
    new_n10160_, new_n10161_, new_n10162_, new_n10163_, new_n10164_,
    new_n10165_, new_n10166_, new_n10167_, new_n10168_, new_n10169_,
    new_n10170_, new_n10171_, new_n10172_, new_n10173_, new_n10174_,
    new_n10175_, new_n10176_, new_n10177_, new_n10178_, new_n10179_,
    new_n10180_, new_n10181_, new_n10182_, new_n10183_, new_n10184_,
    new_n10185_, new_n10186_, new_n10187_, new_n10188_, new_n10189_,
    new_n10190_, new_n10191_, new_n10192_, new_n10193_, new_n10194_,
    new_n10195_, new_n10196_, new_n10197_, new_n10198_, new_n10199_,
    new_n10200_, new_n10201_, new_n10202_, new_n10203_, new_n10204_,
    new_n10205_, new_n10206_, new_n10207_, new_n10208_, new_n10209_,
    new_n10210_, new_n10211_, new_n10212_, new_n10213_, new_n10214_,
    new_n10215_, new_n10216_, new_n10217_, new_n10218_, new_n10219_,
    new_n10220_, new_n10221_, new_n10222_, new_n10223_, new_n10224_,
    new_n10225_, new_n10226_, new_n10227_, new_n10228_, new_n10229_,
    new_n10230_, new_n10231_, new_n10232_, new_n10233_, new_n10234_,
    new_n10235_, new_n10236_, new_n10237_, new_n10238_, new_n10239_,
    new_n10240_, new_n10241_, new_n10242_, new_n10243_, new_n10244_,
    new_n10245_, new_n10246_, new_n10247_, new_n10248_, new_n10249_,
    new_n10250_, new_n10251_, new_n10252_, new_n10253_, new_n10254_,
    new_n10255_, new_n10256_, new_n10257_, new_n10258_, new_n10259_,
    new_n10260_, new_n10261_, new_n10262_, new_n10263_, new_n10264_,
    new_n10265_, new_n10266_, new_n10267_, new_n10268_, new_n10269_,
    new_n10270_, new_n10271_, new_n10272_, new_n10273_, new_n10274_,
    new_n10275_, new_n10276_, new_n10277_, new_n10278_, new_n10279_,
    new_n10280_, new_n10281_, new_n10282_, new_n10283_, new_n10284_,
    new_n10285_, new_n10286_, new_n10287_, new_n10288_, new_n10289_,
    new_n10290_, new_n10291_, new_n10292_, new_n10293_, new_n10294_,
    new_n10295_, new_n10296_, new_n10297_, new_n10298_, new_n10299_,
    new_n10300_, new_n10301_, new_n10302_, new_n10303_, new_n10304_,
    new_n10305_, new_n10306_, new_n10307_, new_n10308_, new_n10309_,
    new_n10310_, new_n10311_, new_n10312_, new_n10313_, new_n10314_,
    new_n10315_, new_n10316_, new_n10317_, new_n10318_, new_n10319_,
    new_n10320_, new_n10321_, new_n10322_, new_n10323_, new_n10324_,
    new_n10325_, new_n10326_, new_n10327_, new_n10328_, new_n10329_,
    new_n10330_, new_n10331_, new_n10332_, new_n10333_, new_n10334_,
    new_n10335_, new_n10336_, new_n10337_, new_n10338_, new_n10339_,
    new_n10340_, new_n10341_, new_n10342_, new_n10343_, new_n10344_,
    new_n10345_, new_n10346_, new_n10347_, new_n10348_, new_n10349_,
    new_n10350_, new_n10351_, new_n10352_, new_n10353_, new_n10354_,
    new_n10355_, new_n10356_, new_n10357_, new_n10358_, new_n10359_,
    new_n10360_, new_n10361_, new_n10362_, new_n10363_, new_n10364_,
    new_n10365_, new_n10366_, new_n10367_, new_n10368_, new_n10369_,
    new_n10370_, new_n10371_, new_n10372_, new_n10373_, new_n10374_,
    new_n10375_, new_n10376_, new_n10377_, new_n10378_, new_n10379_,
    new_n10380_, new_n10381_, new_n10382_, new_n10383_, new_n10384_,
    new_n10385_, new_n10386_, new_n10387_, new_n10388_, new_n10389_,
    new_n10390_, new_n10391_, new_n10392_, new_n10393_, new_n10394_,
    new_n10395_, new_n10396_, new_n10397_, new_n10398_, new_n10399_,
    new_n10400_, new_n10401_, new_n10402_, new_n10403_, new_n10404_,
    new_n10405_, new_n10406_, new_n10407_, new_n10408_, new_n10409_,
    new_n10410_, new_n10411_, new_n10412_, new_n10413_, new_n10414_,
    new_n10415_, new_n10416_, new_n10417_, new_n10418_, new_n10419_,
    new_n10420_, new_n10421_, new_n10422_, new_n10423_, new_n10424_,
    new_n10425_, new_n10426_, new_n10427_, new_n10428_, new_n10429_,
    new_n10430_, new_n10431_, new_n10432_, new_n10433_, new_n10434_,
    new_n10435_, new_n10436_, new_n10437_, new_n10438_, new_n10439_,
    new_n10440_, new_n10441_, new_n10442_, new_n10443_, new_n10444_,
    new_n10445_, new_n10446_, new_n10447_, new_n10448_, new_n10449_,
    new_n10450_, new_n10451_, new_n10452_, new_n10453_, new_n10454_,
    new_n10455_, new_n10456_, new_n10457_, new_n10458_, new_n10459_,
    new_n10460_, new_n10461_, new_n10462_, new_n10463_, new_n10464_,
    new_n10465_, new_n10466_, new_n10467_, new_n10468_, new_n10469_,
    new_n10470_, new_n10471_, new_n10472_, new_n10473_, new_n10474_,
    new_n10475_, new_n10476_, new_n10477_, new_n10478_, new_n10479_,
    new_n10480_, new_n10481_, new_n10482_, new_n10483_, new_n10484_,
    new_n10485_, new_n10486_, new_n10487_, new_n10488_, new_n10489_,
    new_n10490_, new_n10491_, new_n10492_, new_n10493_, new_n10494_,
    new_n10495_, new_n10496_, new_n10497_, new_n10498_, new_n10499_,
    new_n10500_, new_n10501_, new_n10502_, new_n10503_, new_n10504_,
    new_n10505_, new_n10506_, new_n10507_, new_n10508_, new_n10509_,
    new_n10510_, new_n10511_, new_n10512_, new_n10513_, new_n10514_,
    new_n10515_, new_n10516_, new_n10517_, new_n10518_, new_n10519_,
    new_n10520_, new_n10521_, new_n10522_, new_n10523_, new_n10524_,
    new_n10525_, new_n10526_, new_n10527_, new_n10528_, new_n10529_,
    new_n10530_, new_n10531_, new_n10532_, new_n10533_, new_n10534_,
    new_n10535_, new_n10536_, new_n10537_, new_n10538_, new_n10539_,
    new_n10540_, new_n10541_, new_n10542_, new_n10543_, new_n10544_,
    new_n10545_, new_n10546_, new_n10547_, new_n10548_, new_n10549_,
    new_n10550_, new_n10551_, new_n10552_, new_n10553_, new_n10554_,
    new_n10555_, new_n10556_, new_n10557_, new_n10558_, new_n10559_,
    new_n10560_, new_n10561_, new_n10562_, new_n10563_, new_n10564_,
    new_n10565_, new_n10566_, new_n10567_, new_n10568_, new_n10569_,
    new_n10570_, new_n10571_, new_n10572_, new_n10573_, new_n10574_,
    new_n10575_, new_n10576_, new_n10577_, new_n10578_, new_n10579_,
    new_n10580_, new_n10581_, new_n10582_, new_n10583_, new_n10584_,
    new_n10585_, new_n10586_, new_n10587_, new_n10588_, new_n10589_,
    new_n10590_, new_n10591_, new_n10592_, new_n10593_, new_n10594_,
    new_n10595_, new_n10596_, new_n10597_, new_n10598_, new_n10599_,
    new_n10600_, new_n10601_, new_n10602_, new_n10603_, new_n10604_,
    new_n10605_, new_n10606_, new_n10607_, new_n10608_, new_n10609_,
    new_n10610_, new_n10611_, new_n10612_, new_n10613_, new_n10614_,
    new_n10615_, new_n10616_, new_n10617_, new_n10618_, new_n10619_,
    new_n10620_, new_n10621_, new_n10622_, new_n10623_, new_n10624_,
    new_n10625_, new_n10626_, new_n10627_, new_n10628_, new_n10629_,
    new_n10630_, new_n10631_, new_n10632_, new_n10633_, new_n10634_,
    new_n10635_, new_n10636_, new_n10637_, new_n10638_, new_n10639_,
    new_n10640_, new_n10641_, new_n10642_, new_n10643_, new_n10644_,
    new_n10645_, new_n10646_, new_n10647_, new_n10648_, new_n10649_,
    new_n10650_, new_n10651_, new_n10652_, new_n10653_, new_n10654_,
    new_n10655_, new_n10656_, new_n10657_, new_n10658_, new_n10659_,
    new_n10660_, new_n10661_, new_n10662_, new_n10663_, new_n10664_,
    new_n10665_, new_n10666_, new_n10667_, new_n10668_, new_n10669_,
    new_n10670_, new_n10671_, new_n10672_, new_n10673_, new_n10674_,
    new_n10675_, new_n10676_, new_n10677_, new_n10678_, new_n10679_,
    new_n10680_, new_n10681_, new_n10682_, new_n10683_, new_n10684_,
    new_n10685_, new_n10686_, new_n10687_, new_n10688_, new_n10689_,
    new_n10690_, new_n10691_, new_n10692_, new_n10693_, new_n10694_,
    new_n10695_, new_n10696_, new_n10697_, new_n10698_, new_n10699_,
    new_n10700_, new_n10701_, new_n10702_, new_n10703_, new_n10704_,
    new_n10705_, new_n10706_, new_n10707_, new_n10708_, new_n10709_,
    new_n10710_, new_n10711_, new_n10712_, new_n10713_, new_n10714_,
    new_n10715_, new_n10716_, new_n10717_, new_n10718_, new_n10719_,
    new_n10720_, new_n10721_, new_n10722_, new_n10723_, new_n10724_,
    new_n10725_, new_n10726_, new_n10727_, new_n10728_, new_n10729_,
    new_n10730_, new_n10731_, new_n10732_, new_n10733_, new_n10734_,
    new_n10735_, new_n10736_, new_n10737_, new_n10738_, new_n10739_,
    new_n10740_, new_n10741_, new_n10742_, new_n10743_, new_n10744_,
    new_n10745_, new_n10746_, new_n10747_, new_n10748_, new_n10749_,
    new_n10750_, new_n10751_, new_n10752_, new_n10753_, new_n10754_,
    new_n10755_, new_n10756_, new_n10757_, new_n10758_, new_n10759_,
    new_n10760_, new_n10761_, new_n10762_, new_n10763_, new_n10764_,
    new_n10765_, new_n10766_, new_n10767_, new_n10768_, new_n10769_,
    new_n10770_, new_n10771_, new_n10772_, new_n10773_, new_n10774_,
    new_n10775_, new_n10776_, new_n10777_, new_n10778_, new_n10779_,
    new_n10780_, new_n10781_, new_n10782_, new_n10783_, new_n10784_,
    new_n10785_, new_n10786_, new_n10787_, new_n10788_, new_n10789_,
    new_n10790_, new_n10791_, new_n10792_, new_n10793_, new_n10794_,
    new_n10795_, new_n10796_, new_n10797_, new_n10798_, new_n10799_,
    new_n10800_, new_n10801_, new_n10802_, new_n10803_, new_n10804_,
    new_n10805_, new_n10806_, new_n10807_, new_n10808_, new_n10809_,
    new_n10810_, new_n10811_, new_n10812_, new_n10813_, new_n10814_,
    new_n10815_, new_n10816_, new_n10817_, new_n10818_, new_n10819_,
    new_n10820_, new_n10821_, new_n10822_, new_n10823_, new_n10824_,
    new_n10825_, new_n10826_, new_n10827_, new_n10828_, new_n10829_,
    new_n10830_, new_n10831_, new_n10832_, new_n10833_, new_n10834_,
    new_n10835_, new_n10836_, new_n10837_, new_n10838_, new_n10839_,
    new_n10840_, new_n10841_, new_n10842_, new_n10843_, new_n10844_,
    new_n10845_, new_n10846_, new_n10847_, new_n10848_, new_n10849_,
    new_n10850_, new_n10851_, new_n10852_, new_n10853_, new_n10854_,
    new_n10855_, new_n10856_, new_n10857_, new_n10858_, new_n10859_,
    new_n10860_, new_n10861_, new_n10862_, new_n10863_, new_n10864_,
    new_n10865_, new_n10866_, new_n10867_, new_n10868_, new_n10869_,
    new_n10870_, new_n10871_, new_n10872_, new_n10873_, new_n10874_,
    new_n10875_, new_n10876_, new_n10877_, new_n10878_, new_n10879_,
    new_n10880_, new_n10881_, new_n10882_, new_n10883_, new_n10884_,
    new_n10885_, new_n10886_, new_n10887_, new_n10888_, new_n10889_,
    new_n10890_, new_n10891_, new_n10892_, new_n10893_, new_n10894_,
    new_n10895_, new_n10896_, new_n10897_, new_n10898_, new_n10899_,
    new_n10900_, new_n10901_, new_n10902_, new_n10903_, new_n10904_,
    new_n10905_, new_n10906_, new_n10907_, new_n10908_, new_n10909_,
    new_n10910_, new_n10911_, new_n10912_, new_n10913_, new_n10914_,
    new_n10915_, new_n10916_, new_n10917_, new_n10918_, new_n10919_,
    new_n10920_, new_n10921_, new_n10922_, new_n10923_, new_n10924_,
    new_n10925_, new_n10926_, new_n10927_, new_n10928_, new_n10929_,
    new_n10930_, new_n10931_, new_n10932_, new_n10933_, new_n10934_,
    new_n10935_, new_n10936_, new_n10937_, new_n10938_, new_n10939_,
    new_n10940_, new_n10941_, new_n10942_, new_n10943_, new_n10944_,
    new_n10945_, new_n10946_, new_n10947_, new_n10948_, new_n10949_,
    new_n10950_, new_n10951_, new_n10952_, new_n10953_, new_n10954_,
    new_n10955_, new_n10956_, new_n10957_, new_n10958_, new_n10959_,
    new_n10960_, new_n10961_, new_n10962_, new_n10963_, new_n10964_,
    new_n10965_, new_n10966_, new_n10967_, new_n10968_, new_n10969_,
    new_n10970_, new_n10971_, new_n10972_, new_n10973_, new_n10974_,
    new_n10975_, new_n10976_, new_n10977_, new_n10978_, new_n10979_,
    new_n10980_, new_n10981_, new_n10982_, new_n10983_, new_n10984_,
    new_n10985_, new_n10986_, new_n10987_, new_n10988_, new_n10989_,
    new_n10990_, new_n10991_, new_n10992_, new_n10993_, new_n10994_,
    new_n10995_, new_n10996_, new_n10997_, new_n10998_, new_n10999_,
    new_n11000_, new_n11001_, new_n11002_, new_n11003_, new_n11004_,
    new_n11005_, new_n11006_, new_n11007_, new_n11008_, new_n11009_,
    new_n11010_, new_n11011_, new_n11012_, new_n11013_, new_n11014_,
    new_n11015_, new_n11016_, new_n11017_, new_n11018_, new_n11019_,
    new_n11020_, new_n11021_, new_n11022_, new_n11023_, new_n11024_,
    new_n11025_, new_n11026_, new_n11027_, new_n11028_, new_n11029_,
    new_n11030_, new_n11031_, new_n11032_, new_n11033_, new_n11034_,
    new_n11035_, new_n11036_, new_n11037_, new_n11038_, new_n11039_,
    new_n11040_, new_n11041_, new_n11042_, new_n11043_, new_n11044_,
    new_n11045_, new_n11046_, new_n11047_, new_n11048_, new_n11049_,
    new_n11050_, new_n11051_, new_n11052_, new_n11053_, new_n11054_,
    new_n11055_, new_n11056_, new_n11057_, new_n11058_, new_n11059_,
    new_n11060_, new_n11061_, new_n11062_, new_n11063_, new_n11064_,
    new_n11065_, new_n11066_, new_n11067_, new_n11068_, new_n11069_,
    new_n11070_, new_n11071_, new_n11072_, new_n11073_, new_n11074_,
    new_n11075_, new_n11076_, new_n11077_, new_n11078_, new_n11079_,
    new_n11080_, new_n11081_, new_n11082_, new_n11083_, new_n11084_,
    new_n11085_, new_n11086_, new_n11087_, new_n11088_, new_n11089_,
    new_n11090_, new_n11091_, new_n11092_, new_n11093_, new_n11094_,
    new_n11095_, new_n11096_, new_n11097_, new_n11098_, new_n11099_,
    new_n11100_, new_n11101_, new_n11102_, new_n11103_, new_n11104_,
    new_n11105_, new_n11106_, new_n11107_, new_n11108_, new_n11109_,
    new_n11110_, new_n11111_, new_n11112_, new_n11113_, new_n11114_,
    new_n11115_, new_n11116_, new_n11117_, new_n11118_, new_n11119_,
    new_n11120_, new_n11121_, new_n11122_, new_n11123_, new_n11124_,
    new_n11125_, new_n11126_, new_n11127_, new_n11128_, new_n11129_,
    new_n11130_, new_n11131_, new_n11132_, new_n11133_, new_n11134_,
    new_n11135_, new_n11136_, new_n11137_, new_n11138_, new_n11139_,
    new_n11140_, new_n11141_, new_n11142_, new_n11143_, new_n11144_,
    new_n11145_, new_n11146_, new_n11147_, new_n11148_, new_n11149_,
    new_n11150_, new_n11151_, new_n11152_, new_n11153_, new_n11154_,
    new_n11155_, new_n11156_, new_n11157_, new_n11158_, new_n11159_,
    new_n11160_, new_n11161_, new_n11162_, new_n11163_, new_n11164_,
    new_n11165_, new_n11166_, new_n11167_, new_n11168_, new_n11169_,
    new_n11170_, new_n11171_, new_n11172_, new_n11173_, new_n11174_,
    new_n11175_, new_n11176_, new_n11177_, new_n11178_, new_n11179_,
    new_n11180_, new_n11181_, new_n11182_, new_n11183_, new_n11184_,
    new_n11185_, new_n11186_, new_n11187_, new_n11188_, new_n11189_,
    new_n11190_, new_n11191_, new_n11192_, new_n11193_, new_n11194_,
    new_n11195_, new_n11196_, new_n11197_, new_n11198_, new_n11199_,
    new_n11200_, new_n11201_, new_n11202_, new_n11203_, new_n11204_,
    new_n11205_, new_n11206_, new_n11207_, new_n11208_, new_n11209_,
    new_n11210_, new_n11211_, new_n11212_, new_n11213_, new_n11214_,
    new_n11215_, new_n11216_, new_n11217_, new_n11218_, new_n11219_,
    new_n11220_, new_n11221_, new_n11222_, new_n11223_, new_n11224_,
    new_n11225_, new_n11226_, new_n11227_, new_n11228_, new_n11229_,
    new_n11230_, new_n11231_, new_n11232_, new_n11233_, new_n11234_,
    new_n11235_, new_n11236_, new_n11237_, new_n11238_, new_n11239_,
    new_n11240_, new_n11241_, new_n11242_, new_n11243_, new_n11244_,
    new_n11245_, new_n11246_, new_n11247_, new_n11248_, new_n11249_,
    new_n11250_, new_n11251_, new_n11252_, new_n11253_, new_n11254_,
    new_n11255_, new_n11256_, new_n11257_, new_n11258_, new_n11259_,
    new_n11260_, new_n11261_, new_n11262_, new_n11263_, new_n11264_,
    new_n11265_, new_n11266_, new_n11267_, new_n11268_, new_n11269_,
    new_n11270_, new_n11271_, new_n11272_, new_n11273_, new_n11274_,
    new_n11275_, new_n11276_, new_n11277_, new_n11278_, new_n11279_,
    new_n11280_, new_n11281_, new_n11282_, new_n11283_, new_n11284_,
    new_n11285_, new_n11286_, new_n11287_, new_n11288_, new_n11289_,
    new_n11290_, new_n11291_, new_n11292_, new_n11293_, new_n11294_,
    new_n11295_, new_n11296_, new_n11297_, new_n11298_, new_n11299_,
    new_n11300_, new_n11301_, new_n11302_, new_n11303_, new_n11304_,
    new_n11305_, new_n11306_, new_n11307_, new_n11308_, new_n11309_,
    new_n11310_, new_n11311_, new_n11312_, new_n11313_, new_n11314_,
    new_n11315_, new_n11316_, new_n11317_, new_n11318_, new_n11319_,
    new_n11320_, new_n11321_, new_n11322_, new_n11323_, new_n11324_,
    new_n11325_, new_n11326_, new_n11327_, new_n11328_, new_n11329_,
    new_n11330_, new_n11331_, new_n11332_, new_n11333_, new_n11334_,
    new_n11335_, new_n11336_, new_n11337_, new_n11338_, new_n11339_,
    new_n11340_, new_n11341_, new_n11342_, new_n11343_, new_n11344_,
    new_n11345_, new_n11346_, new_n11347_, new_n11348_, new_n11349_,
    new_n11350_, new_n11351_, new_n11352_, new_n11353_, new_n11354_,
    new_n11355_, new_n11356_, new_n11357_, new_n11358_, new_n11359_,
    new_n11360_, new_n11361_, new_n11362_, new_n11363_, new_n11364_,
    new_n11365_, new_n11366_, new_n11367_, new_n11368_, new_n11369_,
    new_n11370_, new_n11371_, new_n11372_, new_n11373_, new_n11374_,
    new_n11375_, new_n11376_, new_n11377_, new_n11378_, new_n11379_,
    new_n11380_, new_n11381_, new_n11382_, new_n11383_, new_n11384_,
    new_n11385_, new_n11386_, new_n11387_, new_n11388_, new_n11389_,
    new_n11390_, new_n11391_, new_n11392_, new_n11393_, new_n11394_,
    new_n11395_, new_n11396_, new_n11397_, new_n11398_, new_n11399_,
    new_n11400_, new_n11401_, new_n11402_, new_n11403_, new_n11404_,
    new_n11405_, new_n11406_, new_n11407_, new_n11408_, new_n11409_,
    new_n11410_, new_n11411_, new_n11412_, new_n11413_, new_n11414_,
    new_n11415_, new_n11416_, new_n11417_, new_n11418_, new_n11419_,
    new_n11420_, new_n11421_, new_n11422_, new_n11423_, new_n11424_,
    new_n11425_, new_n11426_, new_n11427_, new_n11428_, new_n11429_,
    new_n11430_, new_n11431_, new_n11432_, new_n11433_, new_n11434_,
    new_n11435_, new_n11436_, new_n11437_, new_n11438_, new_n11439_,
    new_n11440_, new_n11441_, new_n11442_, new_n11443_, new_n11444_,
    new_n11445_, new_n11446_, new_n11447_, new_n11448_, new_n11449_,
    new_n11450_, new_n11451_, new_n11452_, new_n11453_, new_n11454_,
    new_n11455_, new_n11456_, new_n11457_, new_n11458_, new_n11459_,
    new_n11460_, new_n11461_, new_n11462_, new_n11463_, new_n11464_,
    new_n11465_, new_n11466_, new_n11467_, new_n11468_, new_n11469_,
    new_n11470_, new_n11471_, new_n11472_, new_n11473_, new_n11474_,
    new_n11475_, new_n11476_, new_n11477_, new_n11478_, new_n11479_,
    new_n11480_, new_n11481_, new_n11482_, new_n11483_, new_n11484_,
    new_n11485_, new_n11486_, new_n11487_, new_n11488_, new_n11489_,
    new_n11490_, new_n11491_, new_n11492_, new_n11493_, new_n11494_,
    new_n11495_, new_n11496_, new_n11497_, new_n11498_, new_n11499_,
    new_n11500_, new_n11501_, new_n11502_, new_n11503_, new_n11504_,
    new_n11505_, new_n11506_, new_n11507_, new_n11508_, new_n11509_,
    new_n11510_, new_n11511_, new_n11512_, new_n11513_, new_n11514_,
    new_n11515_, new_n11516_, new_n11517_, new_n11518_, new_n11519_,
    new_n11520_, new_n11521_, new_n11522_, new_n11523_, new_n11524_,
    new_n11525_, new_n11526_, new_n11527_, new_n11528_, new_n11529_,
    new_n11530_, new_n11531_, new_n11532_, new_n11533_, new_n11534_,
    new_n11535_, new_n11536_, new_n11537_, new_n11538_, new_n11539_,
    new_n11540_, new_n11541_, new_n11542_, new_n11543_, new_n11544_,
    new_n11545_, new_n11546_, new_n11547_, new_n11548_, new_n11549_,
    new_n11550_, new_n11551_, new_n11552_, new_n11553_, new_n11554_,
    new_n11555_, new_n11556_, new_n11557_, new_n11558_, new_n11559_,
    new_n11560_, new_n11561_, new_n11562_, new_n11563_, new_n11564_,
    new_n11565_, new_n11566_, new_n11567_, new_n11568_, new_n11569_,
    new_n11570_, new_n11571_, new_n11572_, new_n11573_, new_n11574_,
    new_n11575_, new_n11576_, new_n11577_, new_n11578_, new_n11579_,
    new_n11580_, new_n11581_, new_n11582_, new_n11583_, new_n11584_,
    new_n11585_, new_n11586_, new_n11587_, new_n11588_, new_n11589_,
    new_n11590_, new_n11591_, new_n11592_, new_n11593_, new_n11594_,
    new_n11595_, new_n11596_, new_n11597_, new_n11598_, new_n11599_,
    new_n11600_, new_n11601_, new_n11602_, new_n11603_, new_n11604_,
    new_n11605_, new_n11606_, new_n11607_, new_n11608_, new_n11609_,
    new_n11610_, new_n11611_, new_n11612_, new_n11613_, new_n11614_,
    new_n11615_, new_n11616_, new_n11617_, new_n11618_, new_n11619_,
    new_n11620_, new_n11621_, new_n11622_, new_n11623_, new_n11624_,
    new_n11625_, new_n11626_, new_n11627_, new_n11628_, new_n11629_,
    new_n11630_, new_n11631_, new_n11632_, new_n11633_, new_n11634_,
    new_n11635_, new_n11636_, new_n11637_, new_n11638_, new_n11639_,
    new_n11640_, new_n11641_, new_n11642_, new_n11643_, new_n11644_,
    new_n11645_, new_n11646_, new_n11647_, new_n11648_, new_n11649_,
    new_n11650_, new_n11651_, new_n11652_, new_n11653_, new_n11654_,
    new_n11655_, new_n11656_, new_n11657_, new_n11658_, new_n11659_,
    new_n11660_, new_n11661_, new_n11662_, new_n11663_, new_n11664_,
    new_n11665_, new_n11666_, new_n11667_, new_n11668_, new_n11669_,
    new_n11670_, new_n11671_, new_n11672_, new_n11673_, new_n11674_,
    new_n11675_, new_n11676_, new_n11677_, new_n11678_, new_n11679_,
    new_n11680_, new_n11681_, new_n11682_, new_n11683_, new_n11684_,
    new_n11685_, new_n11686_, new_n11687_, new_n11688_, new_n11689_,
    new_n11690_, new_n11691_, new_n11692_, new_n11693_, new_n11694_,
    new_n11695_, new_n11696_, new_n11697_, new_n11698_, new_n11699_,
    new_n11700_, new_n11701_, new_n11702_, new_n11703_, new_n11704_,
    new_n11705_, new_n11706_, new_n11707_, new_n11708_, new_n11709_,
    new_n11710_, new_n11711_, new_n11712_, new_n11713_, new_n11714_,
    new_n11715_, new_n11716_, new_n11717_, new_n11718_, new_n11719_,
    new_n11720_, new_n11721_, new_n11722_, new_n11723_, new_n11724_,
    new_n11725_, new_n11726_, new_n11727_, new_n11728_, new_n11729_,
    new_n11730_, new_n11731_, new_n11732_, new_n11733_, new_n11734_,
    new_n11735_, new_n11736_, new_n11737_, new_n11738_, new_n11739_,
    new_n11740_, new_n11741_, new_n11742_, new_n11743_, new_n11744_,
    new_n11745_, new_n11746_, new_n11747_, new_n11748_, new_n11749_,
    new_n11750_, new_n11751_, new_n11752_, new_n11753_, new_n11754_,
    new_n11755_, new_n11756_, new_n11757_, new_n11758_, new_n11759_,
    new_n11760_, new_n11761_, new_n11762_, new_n11763_, new_n11764_,
    new_n11765_, new_n11766_, new_n11767_, new_n11768_, new_n11769_,
    new_n11770_, new_n11771_, new_n11772_, new_n11773_, new_n11774_,
    new_n11775_, new_n11776_, new_n11777_, new_n11778_, new_n11779_,
    new_n11780_, new_n11781_, new_n11782_, new_n11783_, new_n11784_,
    new_n11785_, new_n11786_, new_n11787_, new_n11788_, new_n11789_,
    new_n11790_, new_n11791_, new_n11792_, new_n11793_, new_n11794_,
    new_n11795_, new_n11796_, new_n11797_, new_n11798_, new_n11799_,
    new_n11800_, new_n11801_, new_n11802_, new_n11803_, new_n11804_,
    new_n11805_, new_n11806_, new_n11807_, new_n11808_, new_n11809_,
    new_n11810_, new_n11811_, new_n11812_, new_n11813_, new_n11814_,
    new_n11815_, new_n11816_, new_n11817_, new_n11818_, new_n11819_,
    new_n11820_, new_n11821_, new_n11822_, new_n11823_, new_n11824_,
    new_n11825_, new_n11826_, new_n11827_, new_n11828_, new_n11829_,
    new_n11830_, new_n11831_, new_n11832_, new_n11833_, new_n11834_,
    new_n11835_, new_n11836_, new_n11837_, new_n11838_, new_n11839_,
    new_n11840_, new_n11841_, new_n11842_, new_n11843_, new_n11844_,
    new_n11845_, new_n11846_, new_n11847_, new_n11848_, new_n11849_,
    new_n11850_, new_n11851_, new_n11852_, new_n11853_, new_n11854_,
    new_n11855_, new_n11856_, new_n11857_, new_n11858_, new_n11859_,
    new_n11860_, new_n11861_, new_n11862_, new_n11863_, new_n11864_,
    new_n11865_, new_n11866_, new_n11867_, new_n11868_, new_n11869_,
    new_n11870_, new_n11871_, new_n11872_, new_n11873_, new_n11874_,
    new_n11875_, new_n11876_, new_n11877_, new_n11878_, new_n11879_,
    new_n11880_, new_n11881_, new_n11882_, new_n11883_, new_n11884_,
    new_n11885_, new_n11886_, new_n11887_, new_n11888_, new_n11889_,
    new_n11890_, new_n11891_, new_n11892_, new_n11893_, new_n11894_,
    new_n11895_, new_n11896_, new_n11897_, new_n11898_, new_n11899_,
    new_n11900_, new_n11901_, new_n11902_, new_n11903_, new_n11904_,
    new_n11905_, new_n11906_, new_n11907_, new_n11908_, new_n11909_,
    new_n11910_, new_n11911_, new_n11912_, new_n11913_, new_n11914_,
    new_n11915_, new_n11916_, new_n11917_, new_n11918_, new_n11919_,
    new_n11920_, new_n11921_, new_n11922_, new_n11923_, new_n11924_,
    new_n11925_, new_n11926_, new_n11927_, new_n11928_, new_n11929_,
    new_n11930_, new_n11931_, new_n11932_, new_n11933_, new_n11934_,
    new_n11935_, new_n11936_, new_n11937_, new_n11938_, new_n11939_,
    new_n11940_, new_n11941_, new_n11942_, new_n11943_, new_n11944_,
    new_n11945_, new_n11946_, new_n11947_, new_n11948_, new_n11949_,
    new_n11950_, new_n11951_, new_n11952_, new_n11953_, new_n11954_,
    new_n11955_, new_n11956_, new_n11957_, new_n11958_, new_n11959_,
    new_n11960_, new_n11961_, new_n11962_, new_n11963_, new_n11964_,
    new_n11965_, new_n11966_, new_n11967_, new_n11968_, new_n11969_,
    new_n11970_, new_n11971_, new_n11972_, new_n11973_, new_n11974_,
    new_n11975_, new_n11976_, new_n11977_, new_n11978_, new_n11979_,
    new_n11980_, new_n11981_, new_n11982_, new_n11983_, new_n11984_,
    new_n11985_, new_n11986_, new_n11987_, new_n11988_, new_n11989_,
    new_n11990_, new_n11991_, new_n11992_, new_n11993_, new_n11994_,
    new_n11995_, new_n11996_, new_n11997_, new_n11998_, new_n11999_,
    new_n12000_, new_n12001_, new_n12002_, new_n12003_, new_n12004_,
    new_n12005_, new_n12006_, new_n12007_, new_n12008_, new_n12009_,
    new_n12010_, new_n12011_, new_n12012_, new_n12013_, new_n12014_,
    new_n12015_, new_n12016_, new_n12017_, new_n12018_, new_n12019_,
    new_n12020_, new_n12021_, new_n12022_, new_n12023_, new_n12024_,
    new_n12025_, new_n12026_, new_n12027_, new_n12028_, new_n12029_,
    new_n12030_, new_n12031_, new_n12032_, new_n12033_, new_n12034_,
    new_n12035_, new_n12036_, new_n12037_, new_n12038_, new_n12039_,
    new_n12040_, new_n12041_, new_n12042_, new_n12043_, new_n12044_,
    new_n12045_, new_n12046_, new_n12047_, new_n12048_, new_n12049_,
    new_n12050_, new_n12051_, new_n12052_, new_n12053_, new_n12054_,
    new_n12055_, new_n12056_, new_n12057_, new_n12058_, new_n12059_,
    new_n12060_, new_n12061_, new_n12062_, new_n12063_, new_n12064_,
    new_n12065_, new_n12066_, new_n12067_, new_n12068_, new_n12069_,
    new_n12070_, new_n12071_, new_n12072_, new_n12073_, new_n12074_,
    new_n12075_, new_n12076_, new_n12077_, new_n12078_, new_n12079_,
    new_n12080_, new_n12081_, new_n12082_, new_n12083_, new_n12084_,
    new_n12085_, new_n12086_, new_n12087_, new_n12088_, new_n12089_,
    new_n12090_, new_n12091_, new_n12092_, new_n12093_, new_n12094_,
    new_n12095_, new_n12096_, new_n12097_, new_n12098_, new_n12099_,
    new_n12100_, new_n12101_, new_n12102_, new_n12103_, new_n12104_,
    new_n12105_, new_n12106_, new_n12107_, new_n12108_, new_n12109_,
    new_n12110_, new_n12111_, new_n12112_, new_n12113_, new_n12114_,
    new_n12115_, new_n12116_, new_n12117_, new_n12118_, new_n12119_,
    new_n12120_, new_n12121_, new_n12122_, new_n12123_, new_n12124_,
    new_n12125_, new_n12126_, new_n12127_, new_n12128_, new_n12129_,
    new_n12130_, new_n12131_, new_n12132_, new_n12133_, new_n12134_,
    new_n12135_, new_n12136_, new_n12137_, new_n12138_, new_n12139_,
    new_n12140_, new_n12141_, new_n12142_, new_n12143_, new_n12144_,
    new_n12145_, new_n12146_, new_n12147_, new_n12148_, new_n12149_,
    new_n12150_, new_n12151_, new_n12152_, new_n12153_, new_n12154_,
    new_n12155_, new_n12156_, new_n12157_, new_n12158_, new_n12159_,
    new_n12160_, new_n12161_, new_n12162_, new_n12163_, new_n12164_,
    new_n12165_, new_n12166_, new_n12167_, new_n12168_, new_n12169_,
    new_n12170_, new_n12171_, new_n12172_, new_n12173_, new_n12174_,
    new_n12175_, new_n12176_, new_n12177_, new_n12178_, new_n12179_,
    new_n12180_, new_n12181_, new_n12182_, new_n12183_, new_n12184_,
    new_n12185_, new_n12186_, new_n12187_, new_n12188_, new_n12189_,
    new_n12190_, new_n12191_, new_n12192_, new_n12193_, new_n12194_,
    new_n12195_, new_n12196_, new_n12197_, new_n12198_, new_n12199_,
    new_n12200_, new_n12201_, new_n12202_, new_n12203_, new_n12204_,
    new_n12205_, new_n12206_, new_n12207_, new_n12208_, new_n12209_,
    new_n12210_, new_n12211_, new_n12212_, new_n12213_, new_n12214_,
    new_n12215_, new_n12216_, new_n12217_, new_n12218_, new_n12219_,
    new_n12220_, new_n12221_, new_n12222_, new_n12223_, new_n12224_,
    new_n12225_, new_n12226_, new_n12227_, new_n12228_, new_n12229_,
    new_n12230_, new_n12231_, new_n12232_, new_n12233_, new_n12234_,
    new_n12235_, new_n12236_, new_n12237_, new_n12238_, new_n12239_,
    new_n12240_, new_n12241_, new_n12242_, new_n12243_, new_n12244_,
    new_n12245_, new_n12246_, new_n12247_, new_n12248_, new_n12249_,
    new_n12250_, new_n12251_, new_n12252_, new_n12253_, new_n12254_,
    new_n12255_, new_n12256_, new_n12257_, new_n12258_, new_n12259_,
    new_n12260_, new_n12261_, new_n12262_, new_n12263_, new_n12264_,
    new_n12265_, new_n12266_, new_n12267_, new_n12268_, new_n12269_,
    new_n12270_, new_n12271_, new_n12272_, new_n12273_, new_n12274_,
    new_n12275_, new_n12276_, new_n12277_, new_n12278_, new_n12279_,
    new_n12280_, new_n12281_, new_n12282_, new_n12283_, new_n12284_,
    new_n12285_, new_n12286_, new_n12287_, new_n12288_, new_n12289_,
    new_n12290_, new_n12291_, new_n12292_, new_n12293_, new_n12294_,
    new_n12295_, new_n12296_, new_n12297_, new_n12298_, new_n12299_,
    new_n12300_, new_n12301_, new_n12302_, new_n12303_, new_n12304_,
    new_n12305_, new_n12306_, new_n12307_, new_n12308_, new_n12309_,
    new_n12310_, new_n12311_, new_n12312_, new_n12313_, new_n12314_,
    new_n12315_, new_n12316_, new_n12317_, new_n12318_, new_n12319_,
    new_n12320_, new_n12321_, new_n12322_, new_n12323_, new_n12324_,
    new_n12325_, new_n12326_, new_n12327_, new_n12328_, new_n12329_,
    new_n12330_, new_n12331_, new_n12332_, new_n12333_, new_n12334_,
    new_n12335_, new_n12336_, new_n12337_, new_n12338_, new_n12339_,
    new_n12340_, new_n12341_, new_n12342_, new_n12343_, new_n12344_,
    new_n12345_, new_n12346_, new_n12347_, new_n12348_, new_n12349_,
    new_n12350_, new_n12351_, new_n12352_, new_n12353_, new_n12354_,
    new_n12355_, new_n12356_, new_n12357_, new_n12358_, new_n12359_,
    new_n12360_, new_n12361_, new_n12362_, new_n12363_, new_n12364_,
    new_n12365_, new_n12366_, new_n12367_, new_n12368_, new_n12369_,
    new_n12370_, new_n12371_, new_n12372_, new_n12373_, new_n12374_,
    new_n12375_, new_n12376_, new_n12377_, new_n12378_, new_n12379_,
    new_n12380_, new_n12381_, new_n12382_, new_n12383_, new_n12384_,
    new_n12385_, new_n12386_, new_n12387_, new_n12388_, new_n12389_,
    new_n12390_, new_n12391_, new_n12392_, new_n12393_, new_n12394_,
    new_n12395_, new_n12396_, new_n12397_, new_n12398_, new_n12399_,
    new_n12400_, new_n12401_, new_n12402_, new_n12403_, new_n12404_,
    new_n12405_, new_n12406_, new_n12407_, new_n12408_, new_n12409_,
    new_n12410_, new_n12411_, new_n12412_, new_n12413_, new_n12414_,
    new_n12415_, new_n12416_, new_n12417_, new_n12418_, new_n12419_,
    new_n12420_, new_n12421_, new_n12422_, new_n12423_, new_n12424_,
    new_n12425_, new_n12426_, new_n12427_, new_n12428_, new_n12429_,
    new_n12430_, new_n12431_, new_n12432_, new_n12433_, new_n12434_,
    new_n12435_, new_n12436_, new_n12437_, new_n12438_, new_n12439_,
    new_n12440_, new_n12441_, new_n12442_, new_n12443_, new_n12444_,
    new_n12445_, new_n12446_, new_n12447_, new_n12448_, new_n12449_,
    new_n12450_, new_n12451_, new_n12452_, new_n12453_, new_n12454_,
    new_n12455_, new_n12456_, new_n12457_, new_n12458_, new_n12459_,
    new_n12460_, new_n12461_, new_n12462_, new_n12463_, new_n12464_,
    new_n12465_, new_n12466_, new_n12467_, new_n12468_, new_n12469_,
    new_n12470_, new_n12471_, new_n12472_, new_n12473_, new_n12474_,
    new_n12475_, new_n12476_, new_n12477_, new_n12478_, new_n12479_,
    new_n12480_, new_n12481_, new_n12482_, new_n12483_, new_n12484_,
    new_n12485_, new_n12486_, new_n12487_, new_n12488_, new_n12489_,
    new_n12490_, new_n12491_, new_n12492_, new_n12493_, new_n12494_,
    new_n12495_, new_n12496_, new_n12497_, new_n12498_, new_n12499_,
    new_n12500_, new_n12501_, new_n12502_, new_n12503_, new_n12504_,
    new_n12505_, new_n12506_, new_n12507_, new_n12508_, new_n12509_,
    new_n12510_, new_n12511_, new_n12512_, new_n12513_, new_n12514_,
    new_n12515_, new_n12516_, new_n12517_, new_n12518_, new_n12519_,
    new_n12520_, new_n12521_, new_n12522_, new_n12523_, new_n12524_,
    new_n12525_, new_n12526_, new_n12527_, new_n12528_, new_n12529_,
    new_n12530_, new_n12531_, new_n12532_, new_n12533_, new_n12534_,
    new_n12535_, new_n12536_, new_n12537_, new_n12538_, new_n12539_,
    new_n12540_, new_n12541_, new_n12542_, new_n12543_, new_n12544_,
    new_n12545_, new_n12546_, new_n12547_, new_n12548_, new_n12549_,
    new_n12550_, new_n12551_, new_n12552_, new_n12553_, new_n12554_,
    new_n12555_, new_n12556_, new_n12557_, new_n12558_, new_n12559_,
    new_n12560_, new_n12561_, new_n12562_, new_n12563_, new_n12564_,
    new_n12565_, new_n12566_, new_n12567_, new_n12568_, new_n12569_,
    new_n12570_, new_n12571_, new_n12572_, new_n12573_, new_n12574_,
    new_n12575_, new_n12576_, new_n12577_, new_n12578_, new_n12579_,
    new_n12580_, new_n12581_, new_n12582_, new_n12583_, new_n12584_,
    new_n12585_, new_n12586_, new_n12587_, new_n12588_, new_n12589_,
    new_n12590_, new_n12591_, new_n12592_, new_n12593_, new_n12594_,
    new_n12595_, new_n12596_, new_n12597_, new_n12598_, new_n12599_,
    new_n12600_, new_n12601_, new_n12602_, new_n12603_, new_n12604_,
    new_n12605_, new_n12606_, new_n12607_, new_n12608_, new_n12609_,
    new_n12610_, new_n12611_, new_n12612_, new_n12613_, new_n12614_,
    new_n12615_, new_n12616_, new_n12617_, new_n12618_, new_n12619_,
    new_n12620_, new_n12621_, new_n12622_, new_n12623_, new_n12624_,
    new_n12625_, new_n12626_, new_n12627_, new_n12628_, new_n12629_,
    new_n12630_, new_n12631_, new_n12632_, new_n12633_, new_n12634_,
    new_n12635_, new_n12636_, new_n12637_, new_n12638_, new_n12639_,
    new_n12640_, new_n12641_, new_n12642_, new_n12643_, new_n12644_,
    new_n12645_, new_n12646_, new_n12647_, new_n12648_, new_n12649_,
    new_n12650_, new_n12651_, new_n12652_, new_n12653_, new_n12654_,
    new_n12655_, new_n12656_, new_n12657_, new_n12658_, new_n12659_,
    new_n12660_, new_n12661_, new_n12662_, new_n12663_, new_n12664_,
    new_n12665_, new_n12666_, new_n12667_, new_n12668_, new_n12669_,
    new_n12670_, new_n12671_, new_n12672_, new_n12673_, new_n12674_,
    new_n12675_, new_n12676_, new_n12677_, new_n12678_, new_n12679_,
    new_n12680_, new_n12681_, new_n12682_, new_n12683_, new_n12684_,
    new_n12685_, new_n12686_, new_n12687_, new_n12688_, new_n12689_,
    new_n12690_, new_n12691_, new_n12692_, new_n12693_, new_n12694_,
    new_n12695_, new_n12696_, new_n12697_, new_n12698_, new_n12699_,
    new_n12700_, new_n12701_, new_n12702_, new_n12703_, new_n12704_,
    new_n12705_, new_n12706_, new_n12707_, new_n12708_, new_n12709_,
    new_n12710_, new_n12711_, new_n12712_, new_n12713_, new_n12714_,
    new_n12715_, new_n12716_, new_n12717_, new_n12718_, new_n12719_,
    new_n12720_, new_n12721_, new_n12722_, new_n12723_, new_n12724_,
    new_n12725_, new_n12726_, new_n12727_, new_n12728_, new_n12729_,
    new_n12730_, new_n12731_, new_n12732_, new_n12733_, new_n12734_,
    new_n12735_, new_n12736_, new_n12737_, new_n12738_, new_n12739_,
    new_n12740_, new_n12741_, new_n12742_, new_n12743_, new_n12744_,
    new_n12745_, new_n12746_, new_n12747_, new_n12748_, new_n12749_,
    new_n12750_, new_n12751_, new_n12752_, new_n12753_, new_n12754_,
    new_n12755_, new_n12756_, new_n12757_, new_n12758_, new_n12759_,
    new_n12760_, new_n12761_, new_n12762_, new_n12763_, new_n12764_,
    new_n12765_, new_n12766_, new_n12767_, new_n12768_, new_n12769_,
    new_n12770_, new_n12771_, new_n12772_, new_n12773_, new_n12774_,
    new_n12775_, new_n12776_, new_n12777_, new_n12778_, new_n12779_,
    new_n12780_, new_n12781_, new_n12782_, new_n12783_, new_n12784_,
    new_n12785_, new_n12786_, new_n12787_, new_n12788_, new_n12789_,
    new_n12790_, new_n12791_, new_n12792_, new_n12793_, new_n12794_,
    new_n12795_, new_n12796_, new_n12797_, new_n12798_, new_n12799_,
    new_n12800_, new_n12801_, new_n12802_, new_n12803_, new_n12804_,
    new_n12805_, new_n12806_, new_n12807_, new_n12808_, new_n12809_,
    new_n12810_, new_n12811_, new_n12812_, new_n12813_, new_n12814_,
    new_n12815_, new_n12816_, new_n12817_, new_n12818_, new_n12819_,
    new_n12820_, new_n12821_, new_n12822_, new_n12823_, new_n12824_,
    new_n12825_, new_n12826_, new_n12827_, new_n12828_, new_n12829_,
    new_n12830_, new_n12831_, new_n12832_, new_n12833_, new_n12834_,
    new_n12835_, new_n12836_, new_n12837_, new_n12838_, new_n12839_,
    new_n12840_, new_n12841_, new_n12842_, new_n12843_, new_n12844_,
    new_n12845_, new_n12846_, new_n12847_, new_n12848_, new_n12849_,
    new_n12850_, new_n12851_, new_n12852_, new_n12853_, new_n12854_,
    new_n12855_, new_n12856_, new_n12857_, new_n12858_, new_n12859_,
    new_n12860_, new_n12861_, new_n12862_, new_n12863_, new_n12864_,
    new_n12865_, new_n12866_, new_n12867_, new_n12868_, new_n12869_,
    new_n12870_, new_n12871_, new_n12872_, new_n12873_, new_n12874_,
    new_n12875_, new_n12876_, new_n12877_, new_n12878_, new_n12879_,
    new_n12880_, new_n12881_, new_n12882_, new_n12883_, new_n12884_,
    new_n12885_, new_n12886_, new_n12887_, new_n12888_, new_n12889_,
    new_n12890_, new_n12891_, new_n12892_, new_n12893_, new_n12894_,
    new_n12895_, new_n12896_, new_n12897_, new_n12898_, new_n12899_,
    new_n12900_, new_n12901_, new_n12902_, new_n12903_, new_n12904_,
    new_n12905_, new_n12906_, new_n12907_, new_n12908_, new_n12909_,
    new_n12910_, new_n12911_, new_n12912_, new_n12913_, new_n12914_,
    new_n12915_, new_n12916_, new_n12917_, new_n12918_, new_n12919_,
    new_n12920_, new_n12921_, new_n12922_, new_n12923_, new_n12924_,
    new_n12925_, new_n12926_, new_n12927_, new_n12928_, new_n12929_,
    new_n12930_, new_n12931_, new_n12932_, new_n12933_, new_n12934_,
    new_n12935_, new_n12936_, new_n12937_, new_n12938_, new_n12939_,
    new_n12940_, new_n12941_, new_n12942_, new_n12943_, new_n12944_,
    new_n12945_, new_n12946_, new_n12947_, new_n12948_, new_n12949_,
    new_n12950_, new_n12951_, new_n12952_, new_n12953_, new_n12954_,
    new_n12955_, new_n12956_, new_n12957_, new_n12958_, new_n12959_,
    new_n12960_, new_n12961_, new_n12962_, new_n12963_, new_n12964_,
    new_n12965_, new_n12966_, new_n12967_, new_n12968_, new_n12969_,
    new_n12970_, new_n12971_, new_n12972_, new_n12973_, new_n12974_,
    new_n12975_, new_n12976_, new_n12977_, new_n12978_, new_n12979_,
    new_n12980_, new_n12981_, new_n12982_, new_n12983_, new_n12984_,
    new_n12985_, new_n12986_, new_n12987_, new_n12988_, new_n12989_,
    new_n12990_, new_n12991_, new_n12992_, new_n12993_, new_n12994_,
    new_n12995_, new_n12996_, new_n12997_, new_n12998_, new_n12999_,
    new_n13000_, new_n13001_, new_n13002_, new_n13003_, new_n13004_,
    new_n13005_, new_n13006_, new_n13007_, new_n13008_, new_n13009_,
    new_n13010_, new_n13011_, new_n13012_, new_n13013_, new_n13014_,
    new_n13015_, new_n13016_, new_n13017_, new_n13018_, new_n13019_,
    new_n13020_, new_n13021_, new_n13022_, new_n13023_, new_n13024_,
    new_n13025_, new_n13026_, new_n13027_, new_n13028_, new_n13029_,
    new_n13030_, new_n13031_, new_n13032_, new_n13033_, new_n13034_,
    new_n13035_, new_n13036_, new_n13037_, new_n13038_, new_n13039_,
    new_n13040_, new_n13041_, new_n13042_, new_n13043_, new_n13044_,
    new_n13045_, new_n13046_, new_n13047_, new_n13048_, new_n13049_,
    new_n13050_, new_n13051_, new_n13052_, new_n13053_, new_n13054_,
    new_n13055_, new_n13056_, new_n13057_, new_n13058_, new_n13059_,
    new_n13060_, new_n13061_, new_n13062_, new_n13063_, new_n13064_,
    new_n13065_, new_n13066_, new_n13067_, new_n13068_, new_n13069_,
    new_n13070_, new_n13071_, new_n13072_, new_n13073_, new_n13074_,
    new_n13075_, new_n13076_, new_n13077_, new_n13078_, new_n13079_,
    new_n13080_, new_n13081_, new_n13082_, new_n13083_, new_n13084_,
    new_n13085_, new_n13086_, new_n13087_, new_n13088_, new_n13089_,
    new_n13090_, new_n13091_, new_n13092_, new_n13093_, new_n13094_,
    new_n13095_, new_n13096_, new_n13097_, new_n13098_, new_n13099_,
    new_n13100_, new_n13101_, new_n13102_, new_n13103_, new_n13104_,
    new_n13105_, new_n13106_, new_n13107_, new_n13108_, new_n13109_,
    new_n13110_, new_n13111_, new_n13112_, new_n13113_, new_n13114_,
    new_n13115_, new_n13116_, new_n13117_, new_n13118_, new_n13119_,
    new_n13120_, new_n13121_, new_n13122_, new_n13123_, new_n13124_,
    new_n13125_, new_n13126_, new_n13127_, new_n13128_, new_n13129_,
    new_n13130_, new_n13131_, new_n13132_, new_n13133_, new_n13134_,
    new_n13135_, new_n13136_, new_n13137_, new_n13138_, new_n13139_,
    new_n13140_, new_n13141_, new_n13142_, new_n13143_, new_n13144_,
    new_n13145_, new_n13146_, new_n13147_, new_n13148_, new_n13149_,
    new_n13150_, new_n13151_, new_n13152_, new_n13153_, new_n13154_,
    new_n13155_, new_n13156_, new_n13157_, new_n13158_, new_n13159_,
    new_n13160_, new_n13161_, new_n13162_, new_n13163_, new_n13164_,
    new_n13165_, new_n13166_, new_n13167_, new_n13168_, new_n13169_,
    new_n13170_, new_n13171_, new_n13172_, new_n13173_, new_n13174_,
    new_n13175_, new_n13176_, new_n13177_, new_n13178_, new_n13179_,
    new_n13180_, new_n13181_, new_n13182_, new_n13183_, new_n13184_,
    new_n13185_, new_n13186_, new_n13187_, new_n13188_, new_n13189_,
    new_n13190_, new_n13191_, new_n13192_, new_n13193_, new_n13194_,
    new_n13195_, new_n13196_, new_n13197_, new_n13198_, new_n13199_,
    new_n13200_, new_n13201_, new_n13202_, new_n13203_, new_n13204_,
    new_n13205_, new_n13206_, new_n13207_, new_n13208_, new_n13209_,
    new_n13210_, new_n13211_, new_n13212_, new_n13213_, new_n13214_,
    new_n13215_, new_n13216_, new_n13217_, new_n13218_, new_n13219_,
    new_n13220_, new_n13221_, new_n13222_, new_n13223_, new_n13224_,
    new_n13225_, new_n13226_, new_n13227_, new_n13228_, new_n13229_,
    new_n13230_, new_n13231_, new_n13232_, new_n13233_, new_n13234_,
    new_n13235_, new_n13236_, new_n13237_, new_n13238_, new_n13239_,
    new_n13240_, new_n13241_, new_n13242_, new_n13243_, new_n13244_,
    new_n13245_, new_n13246_, new_n13247_, new_n13248_, new_n13249_,
    new_n13250_, new_n13251_, new_n13252_, new_n13253_, new_n13254_,
    new_n13255_, new_n13256_, new_n13257_, new_n13258_, new_n13259_,
    new_n13260_, new_n13261_, new_n13262_, new_n13263_, new_n13264_,
    new_n13265_, new_n13266_, new_n13267_, new_n13268_, new_n13269_,
    new_n13270_, new_n13271_, new_n13272_, new_n13273_, new_n13274_,
    new_n13275_, new_n13276_, new_n13277_, new_n13278_, new_n13279_,
    new_n13280_, new_n13281_, new_n13282_, new_n13283_, new_n13284_,
    new_n13285_, new_n13286_, new_n13287_, new_n13288_, new_n13289_,
    new_n13290_, new_n13291_, new_n13292_, new_n13293_, new_n13294_,
    new_n13295_, new_n13296_, new_n13297_, new_n13298_, new_n13299_,
    new_n13300_, new_n13301_, new_n13302_, new_n13303_, new_n13304_,
    new_n13305_, new_n13306_, new_n13307_, new_n13308_, new_n13309_,
    new_n13310_, new_n13311_, new_n13312_, new_n13313_, new_n13314_,
    new_n13315_, new_n13316_, new_n13317_, new_n13318_, new_n13319_,
    new_n13320_, new_n13321_, new_n13322_, new_n13323_, new_n13324_,
    new_n13325_, new_n13326_, new_n13327_, new_n13328_, new_n13329_,
    new_n13330_, new_n13331_, new_n13332_, new_n13333_, new_n13334_,
    new_n13335_, new_n13336_, new_n13337_, new_n13338_, new_n13339_,
    new_n13340_, new_n13341_, new_n13342_, new_n13343_, new_n13344_,
    new_n13345_, new_n13346_, new_n13347_, new_n13348_, new_n13349_,
    new_n13350_, new_n13351_, new_n13352_, new_n13353_, new_n13354_,
    new_n13355_, new_n13356_, new_n13357_, new_n13358_, new_n13359_,
    new_n13360_, new_n13361_, new_n13362_, new_n13363_, new_n13364_,
    new_n13365_, new_n13366_, new_n13367_, new_n13368_, new_n13369_,
    new_n13370_, new_n13371_, new_n13372_, new_n13373_, new_n13374_,
    new_n13375_, new_n13376_, new_n13377_, new_n13378_, new_n13379_,
    new_n13380_, new_n13381_, new_n13382_, new_n13383_, new_n13384_,
    new_n13385_, new_n13386_, new_n13387_, new_n13388_, new_n13389_,
    new_n13390_, new_n13391_, new_n13392_, new_n13393_, new_n13394_,
    new_n13395_, new_n13396_, new_n13397_, new_n13398_, new_n13399_,
    new_n13400_, new_n13401_, new_n13402_, new_n13403_, new_n13404_,
    new_n13405_, new_n13406_, new_n13407_, new_n13408_, new_n13409_,
    new_n13410_, new_n13411_, new_n13412_, new_n13413_, new_n13414_,
    new_n13415_, new_n13416_, new_n13417_, new_n13418_, new_n13419_,
    new_n13420_, new_n13421_, new_n13422_, new_n13423_, new_n13424_,
    new_n13425_, new_n13426_, new_n13427_, new_n13428_, new_n13429_,
    new_n13430_, new_n13431_, new_n13432_, new_n13433_, new_n13434_,
    new_n13435_, new_n13436_, new_n13437_, new_n13438_, new_n13439_,
    new_n13440_, new_n13441_, new_n13442_, new_n13443_, new_n13444_,
    new_n13445_, new_n13446_, new_n13447_, new_n13448_, new_n13449_,
    new_n13450_, new_n13451_, new_n13452_, new_n13453_, new_n13454_,
    new_n13455_, new_n13456_, new_n13457_, new_n13458_, new_n13459_,
    new_n13460_, new_n13461_, new_n13462_, new_n13463_, new_n13464_,
    new_n13465_, new_n13466_, new_n13467_, new_n13468_, new_n13469_,
    new_n13470_, new_n13471_, new_n13472_, new_n13473_, new_n13474_,
    new_n13475_, new_n13476_, new_n13477_, new_n13478_, new_n13479_,
    new_n13480_, new_n13481_, new_n13482_, new_n13483_, new_n13484_,
    new_n13485_, new_n13486_, new_n13487_, new_n13488_, new_n13489_,
    new_n13490_, new_n13491_, new_n13492_, new_n13493_, new_n13494_,
    new_n13495_, new_n13496_, new_n13497_, new_n13498_, new_n13499_,
    new_n13500_, new_n13501_, new_n13502_, new_n13503_, new_n13504_,
    new_n13505_, new_n13506_, new_n13507_, new_n13508_, new_n13509_,
    new_n13510_, new_n13511_, new_n13512_, new_n13513_, new_n13514_,
    new_n13515_, new_n13516_, new_n13517_, new_n13518_, new_n13519_,
    new_n13520_, new_n13521_, new_n13522_, new_n13523_, new_n13524_,
    new_n13525_, new_n13526_, new_n13527_, new_n13528_, new_n13529_,
    new_n13530_, new_n13531_, new_n13532_, new_n13533_, new_n13534_,
    new_n13535_, new_n13536_, new_n13537_, new_n13538_, new_n13539_,
    new_n13540_, new_n13541_, new_n13542_, new_n13543_, new_n13544_,
    new_n13545_, new_n13546_, new_n13547_, new_n13548_, new_n13549_,
    new_n13550_, new_n13551_, new_n13552_, new_n13553_, new_n13554_,
    new_n13555_, new_n13556_, new_n13557_, new_n13558_, new_n13559_,
    new_n13560_, new_n13561_, new_n13562_, new_n13563_, new_n13564_,
    new_n13565_, new_n13566_, new_n13567_, new_n13568_, new_n13569_,
    new_n13570_, new_n13571_, new_n13572_, new_n13573_, new_n13574_,
    new_n13575_, new_n13576_, new_n13577_, new_n13578_, new_n13579_,
    new_n13580_, new_n13581_, new_n13582_, new_n13583_, new_n13584_,
    new_n13585_, new_n13586_, new_n13587_, new_n13588_, new_n13589_,
    new_n13590_, new_n13591_, new_n13592_, new_n13593_, new_n13594_,
    new_n13595_, new_n13596_, new_n13597_, new_n13598_, new_n13599_,
    new_n13600_, new_n13601_, new_n13602_, new_n13603_, new_n13604_,
    new_n13605_, new_n13606_, new_n13607_, new_n13608_, new_n13609_,
    new_n13610_, new_n13611_, new_n13612_, new_n13613_, new_n13614_,
    new_n13615_, new_n13616_, new_n13617_, new_n13618_, new_n13619_,
    new_n13620_, new_n13621_, new_n13622_, new_n13623_, new_n13624_,
    new_n13625_, new_n13626_, new_n13627_, new_n13628_, new_n13629_,
    new_n13630_, new_n13631_, new_n13632_, new_n13633_, new_n13634_,
    new_n13635_, new_n13636_, new_n13637_, new_n13638_, new_n13639_,
    new_n13640_, new_n13641_, new_n13642_, new_n13643_, new_n13644_,
    new_n13645_, new_n13646_, new_n13647_, new_n13648_, new_n13649_,
    new_n13650_, new_n13651_, new_n13652_, new_n13653_, new_n13654_,
    new_n13655_, new_n13656_, new_n13657_, new_n13658_, new_n13659_,
    new_n13660_, new_n13661_, new_n13662_, new_n13663_, new_n13664_,
    new_n13665_, new_n13666_, new_n13667_, new_n13668_, new_n13669_,
    new_n13670_, new_n13671_, new_n13672_, new_n13673_, new_n13674_,
    new_n13675_, new_n13676_, new_n13677_, new_n13678_, new_n13679_,
    new_n13680_, new_n13681_, new_n13682_, new_n13683_, new_n13684_,
    new_n13685_, new_n13686_, new_n13687_, new_n13688_, new_n13689_,
    new_n13690_, new_n13691_, new_n13692_, new_n13693_, new_n13694_,
    new_n13695_, new_n13696_, new_n13697_, new_n13698_, new_n13699_,
    new_n13700_, new_n13701_, new_n13702_, new_n13703_, new_n13704_,
    new_n13705_, new_n13706_, new_n13707_, new_n13708_, new_n13709_,
    new_n13710_, new_n13711_, new_n13712_, new_n13713_, new_n13714_,
    new_n13715_, new_n13716_, new_n13717_, new_n13718_, new_n13719_,
    new_n13720_, new_n13721_, new_n13722_, new_n13723_, new_n13724_,
    new_n13725_, new_n13726_, new_n13727_, new_n13728_, new_n13729_,
    new_n13730_, new_n13731_, new_n13732_, new_n13733_, new_n13734_,
    new_n13735_, new_n13736_, new_n13737_, new_n13738_, new_n13739_,
    new_n13740_, new_n13741_, new_n13742_, new_n13743_, new_n13744_,
    new_n13745_, new_n13746_, new_n13747_, new_n13748_, new_n13749_,
    new_n13750_, new_n13751_, new_n13752_, new_n13753_, new_n13754_,
    new_n13755_, new_n13756_, new_n13757_, new_n13758_, new_n13759_,
    new_n13760_, new_n13761_, new_n13762_, new_n13763_, new_n13764_,
    new_n13765_, new_n13766_, new_n13767_, new_n13768_, new_n13769_,
    new_n13770_, new_n13771_, new_n13772_, new_n13773_, new_n13774_,
    new_n13775_, new_n13776_, new_n13777_, new_n13778_, new_n13779_,
    new_n13780_, new_n13781_, new_n13782_, new_n13783_, new_n13784_,
    new_n13785_, new_n13786_, new_n13787_, new_n13788_, new_n13789_,
    new_n13790_, new_n13791_, new_n13792_, new_n13793_, new_n13794_,
    new_n13795_, new_n13796_, new_n13797_, new_n13798_, new_n13799_,
    new_n13800_, new_n13801_, new_n13802_, new_n13803_, new_n13804_,
    new_n13805_, new_n13806_, new_n13807_, new_n13808_, new_n13809_,
    new_n13810_, new_n13811_, new_n13812_, new_n13813_, new_n13814_,
    new_n13815_, new_n13816_, new_n13817_, new_n13818_, new_n13819_,
    new_n13820_, new_n13821_, new_n13822_, new_n13823_, new_n13824_,
    new_n13825_, new_n13826_, new_n13827_, new_n13828_, new_n13829_,
    new_n13830_, new_n13831_, new_n13832_, new_n13833_, new_n13834_,
    new_n13835_, new_n13836_, new_n13837_, new_n13838_, new_n13839_,
    new_n13840_, new_n13841_, new_n13842_, new_n13843_, new_n13844_,
    new_n13845_, new_n13846_, new_n13847_, new_n13848_, new_n13849_,
    new_n13850_, new_n13851_, new_n13852_, new_n13853_, new_n13854_,
    new_n13855_, new_n13856_, new_n13857_, new_n13858_, new_n13859_,
    new_n13860_, new_n13861_, new_n13862_, new_n13863_, new_n13864_,
    new_n13865_, new_n13866_, new_n13867_, new_n13868_, new_n13869_,
    new_n13870_, new_n13871_, new_n13872_, new_n13873_, new_n13874_,
    new_n13875_, new_n13876_, new_n13877_, new_n13878_, new_n13879_,
    new_n13880_, new_n13881_, new_n13882_, new_n13883_, new_n13884_,
    new_n13885_, new_n13886_, new_n13887_, new_n13888_, new_n13889_,
    new_n13890_, new_n13891_, new_n13892_, new_n13893_, new_n13894_,
    new_n13895_, new_n13896_, new_n13897_, new_n13898_, new_n13899_,
    new_n13900_, new_n13901_, new_n13902_, new_n13903_, new_n13904_,
    new_n13905_, new_n13906_, new_n13907_, new_n13908_, new_n13909_,
    new_n13910_, new_n13911_, new_n13912_, new_n13913_, new_n13914_,
    new_n13915_, new_n13916_, new_n13917_, new_n13918_, new_n13919_,
    new_n13920_, new_n13921_, new_n13922_, new_n13923_, new_n13924_,
    new_n13925_, new_n13926_, new_n13927_, new_n13928_, new_n13929_,
    new_n13930_, new_n13931_, new_n13932_, new_n13933_, new_n13934_,
    new_n13935_, new_n13936_, new_n13937_, new_n13938_, new_n13939_,
    new_n13940_, new_n13941_, new_n13942_, new_n13943_, new_n13944_,
    new_n13945_, new_n13946_, new_n13947_, new_n13948_, new_n13949_,
    new_n13950_, new_n13951_, new_n13952_, new_n13953_, new_n13954_,
    new_n13955_, new_n13956_, new_n13957_, new_n13958_, new_n13959_,
    new_n13960_, new_n13961_, new_n13962_, new_n13963_, new_n13964_,
    new_n13965_, new_n13966_, new_n13967_, new_n13968_, new_n13969_,
    new_n13970_, new_n13971_, new_n13972_, new_n13973_, new_n13974_,
    new_n13975_, new_n13976_, new_n13977_, new_n13978_, new_n13979_,
    new_n13980_, new_n13981_, new_n13982_, new_n13983_, new_n13984_,
    new_n13985_, new_n13986_, new_n13987_, new_n13988_, new_n13989_,
    new_n13990_, new_n13991_, new_n13992_, new_n13993_, new_n13994_,
    new_n13995_, new_n13996_, new_n13997_, new_n13998_, new_n13999_,
    new_n14000_, new_n14001_, new_n14002_, new_n14003_, new_n14004_,
    new_n14005_, new_n14006_, new_n14007_, new_n14008_, new_n14009_,
    new_n14010_, new_n14011_, new_n14012_, new_n14013_, new_n14014_,
    new_n14015_, new_n14016_, new_n14017_, new_n14018_, new_n14019_,
    new_n14020_, new_n14021_, new_n14022_, new_n14023_, new_n14024_,
    new_n14025_, new_n14026_, new_n14027_, new_n14028_, new_n14029_,
    new_n14030_, new_n14031_, new_n14032_, new_n14033_, new_n14034_,
    new_n14035_, new_n14036_, new_n14037_, new_n14038_, new_n14039_,
    new_n14040_, new_n14041_, new_n14042_, new_n14043_, new_n14044_,
    new_n14045_, new_n14046_, new_n14047_, new_n14048_, new_n14049_,
    new_n14050_, new_n14051_, new_n14052_, new_n14053_, new_n14054_,
    new_n14055_, new_n14056_, new_n14057_, new_n14058_, new_n14059_,
    new_n14060_, new_n14061_, new_n14062_, new_n14063_, new_n14064_,
    new_n14065_, new_n14066_, new_n14067_, new_n14068_, new_n14069_,
    new_n14070_, new_n14071_, new_n14072_, new_n14073_, new_n14074_,
    new_n14075_, new_n14076_, new_n14077_, new_n14078_, new_n14079_,
    new_n14080_, new_n14081_, new_n14082_, new_n14083_, new_n14084_,
    new_n14085_, new_n14086_, new_n14087_, new_n14088_, new_n14089_,
    new_n14090_, new_n14091_, new_n14092_, new_n14093_, new_n14094_,
    new_n14095_, new_n14096_, new_n14097_, new_n14098_, new_n14099_,
    new_n14100_, new_n14101_, new_n14102_, new_n14103_, new_n14104_,
    new_n14105_, new_n14106_, new_n14107_, new_n14108_, new_n14109_,
    new_n14110_, new_n14111_, new_n14112_, new_n14113_, new_n14114_,
    new_n14115_, new_n14116_, new_n14117_, new_n14118_, new_n14119_,
    new_n14120_, new_n14121_, new_n14122_, new_n14123_, new_n14124_,
    new_n14125_, new_n14126_, new_n14127_, new_n14128_, new_n14129_,
    new_n14130_, new_n14131_, new_n14132_, new_n14133_, new_n14134_,
    new_n14135_, new_n14136_, new_n14137_, new_n14138_, new_n14139_,
    new_n14140_, new_n14141_, new_n14142_, new_n14143_, new_n14144_,
    new_n14145_, new_n14146_, new_n14147_, new_n14148_, new_n14149_,
    new_n14150_, new_n14151_, new_n14152_, new_n14153_, new_n14154_,
    new_n14155_, new_n14156_, new_n14157_, new_n14158_, new_n14159_,
    new_n14160_, new_n14161_, new_n14162_, new_n14163_, new_n14164_,
    new_n14165_, new_n14166_, new_n14167_, new_n14168_, new_n14169_,
    new_n14170_, new_n14171_, new_n14172_, new_n14173_, new_n14174_,
    new_n14175_, new_n14176_, new_n14177_, new_n14178_, new_n14179_,
    new_n14180_, new_n14181_, new_n14182_, new_n14183_, new_n14184_,
    new_n14185_, new_n14186_, new_n14187_, new_n14188_, new_n14189_,
    new_n14190_, new_n14191_, new_n14192_, new_n14193_, new_n14194_,
    new_n14195_, new_n14196_, new_n14197_, new_n14198_, new_n14199_,
    new_n14200_, new_n14201_, new_n14202_, new_n14203_, new_n14204_,
    new_n14205_, new_n14206_, new_n14207_, new_n14208_, new_n14209_,
    new_n14210_, new_n14211_, new_n14212_, new_n14213_, new_n14214_,
    new_n14215_, new_n14216_, new_n14217_, new_n14218_, new_n14219_,
    new_n14220_, new_n14221_, new_n14222_, new_n14223_, new_n14224_,
    new_n14225_, new_n14226_, new_n14227_, new_n14228_, new_n14229_,
    new_n14230_, new_n14231_, new_n14232_, new_n14233_, new_n14234_,
    new_n14235_, new_n14236_, new_n14237_, new_n14238_, new_n14239_,
    new_n14240_, new_n14241_, new_n14242_, new_n14243_, new_n14244_,
    new_n14245_, new_n14246_, new_n14247_, new_n14248_, new_n14249_,
    new_n14250_, new_n14251_, new_n14252_, new_n14253_, new_n14254_,
    new_n14255_, new_n14256_, new_n14257_, new_n14258_, new_n14259_,
    new_n14260_, new_n14261_, new_n14262_, new_n14263_, new_n14264_,
    new_n14265_, new_n14266_, new_n14267_, new_n14268_, new_n14269_,
    new_n14270_, new_n14271_, new_n14272_, new_n14273_, new_n14274_,
    new_n14275_, new_n14276_, new_n14277_, new_n14278_, new_n14279_,
    new_n14280_, new_n14281_, new_n14282_, new_n14283_, new_n14284_,
    new_n14285_, new_n14286_, new_n14287_, new_n14288_, new_n14289_,
    new_n14290_, new_n14291_, new_n14292_, new_n14293_, new_n14294_,
    new_n14295_, new_n14296_, new_n14297_, new_n14298_, new_n14299_,
    new_n14300_, new_n14301_, new_n14302_, new_n14303_, new_n14304_,
    new_n14305_, new_n14306_, new_n14307_, new_n14308_, new_n14309_,
    new_n14310_, new_n14311_, new_n14312_, new_n14313_, new_n14314_,
    new_n14315_, new_n14316_, new_n14317_, new_n14318_, new_n14319_,
    new_n14320_, new_n14321_, new_n14322_, new_n14323_, new_n14324_,
    new_n14325_, new_n14326_, new_n14327_, new_n14328_, new_n14329_,
    new_n14330_, new_n14331_, new_n14332_, new_n14333_, new_n14334_,
    new_n14335_, new_n14336_, new_n14337_, new_n14338_, new_n14339_,
    new_n14340_, new_n14341_, new_n14342_, new_n14343_, new_n14344_,
    new_n14345_, new_n14346_, new_n14347_, new_n14348_, new_n14349_,
    new_n14350_, new_n14351_, new_n14352_, new_n14353_, new_n14354_,
    new_n14355_, new_n14356_, new_n14357_, new_n14358_, new_n14359_,
    new_n14360_, new_n14361_, new_n14362_, new_n14363_, new_n14364_,
    new_n14365_, new_n14366_, new_n14367_, new_n14368_, new_n14369_,
    new_n14370_, new_n14371_, new_n14372_, new_n14373_, new_n14374_,
    new_n14375_, new_n14376_, new_n14377_, new_n14378_, new_n14379_,
    new_n14380_, new_n14381_, new_n14382_, new_n14383_, new_n14384_,
    new_n14385_, new_n14386_, new_n14387_, new_n14388_, new_n14389_,
    new_n14390_, new_n14391_, new_n14392_, new_n14393_, new_n14394_,
    new_n14395_, new_n14396_, new_n14397_, new_n14398_, new_n14399_,
    new_n14400_, new_n14401_, new_n14402_, new_n14403_, new_n14404_,
    new_n14405_, new_n14406_, new_n14407_, new_n14408_, new_n14409_,
    new_n14410_, new_n14411_, new_n14412_, new_n14413_, new_n14414_,
    new_n14415_, new_n14416_, new_n14417_, new_n14418_, new_n14419_,
    new_n14420_, new_n14421_, new_n14422_, new_n14423_, new_n14424_,
    new_n14425_, new_n14426_, new_n14427_, new_n14428_, new_n14429_,
    new_n14430_, new_n14431_, new_n14432_, new_n14433_, new_n14434_,
    new_n14435_, new_n14436_, new_n14437_, new_n14438_, new_n14439_,
    new_n14440_, new_n14441_, new_n14442_, new_n14443_, new_n14444_,
    new_n14445_, new_n14446_, new_n14447_, new_n14448_, new_n14449_,
    new_n14450_, new_n14451_, new_n14452_, new_n14453_, new_n14454_,
    new_n14455_, new_n14456_, new_n14457_, new_n14458_, new_n14459_,
    new_n14460_, new_n14461_, new_n14462_, new_n14463_, new_n14464_,
    new_n14465_, new_n14466_, new_n14467_, new_n14468_, new_n14469_,
    new_n14470_, new_n14471_, new_n14472_, new_n14473_, new_n14474_,
    new_n14475_, new_n14476_, new_n14477_, new_n14478_, new_n14479_,
    new_n14480_, new_n14481_, new_n14482_, new_n14483_, new_n14484_,
    new_n14485_, new_n14486_, new_n14487_, new_n14488_, new_n14489_,
    new_n14490_, new_n14491_, new_n14492_, new_n14493_, new_n14494_,
    new_n14495_, new_n14496_, new_n14497_, new_n14498_, new_n14499_,
    new_n14500_, new_n14501_, new_n14502_, new_n14503_, new_n14504_,
    new_n14505_, new_n14506_, new_n14507_, new_n14508_, new_n14509_,
    new_n14510_, new_n14511_, new_n14512_, new_n14513_, new_n14514_,
    new_n14515_, new_n14516_, new_n14517_, new_n14518_, new_n14519_,
    new_n14520_, new_n14521_, new_n14522_, new_n14523_, new_n14524_,
    new_n14525_, new_n14526_, new_n14527_, new_n14528_, new_n14529_,
    new_n14530_, new_n14531_, new_n14532_, new_n14533_, new_n14534_,
    new_n14535_, new_n14536_, new_n14537_, new_n14538_, new_n14539_,
    new_n14540_, new_n14541_, new_n14542_, new_n14543_, new_n14544_,
    new_n14545_, new_n14546_, new_n14547_, new_n14548_, new_n14549_,
    new_n14550_, new_n14551_, new_n14552_, new_n14553_, new_n14554_,
    new_n14555_, new_n14556_, new_n14557_, new_n14558_, new_n14559_,
    new_n14560_, new_n14561_, new_n14562_, new_n14563_, new_n14564_,
    new_n14565_, new_n14566_, new_n14567_, new_n14568_, new_n14569_,
    new_n14570_, new_n14571_, new_n14572_, new_n14573_, new_n14574_,
    new_n14575_, new_n14576_, new_n14577_, new_n14578_, new_n14579_,
    new_n14580_, new_n14581_, new_n14582_, new_n14583_, new_n14584_,
    new_n14585_, new_n14586_, new_n14587_, new_n14588_, new_n14589_,
    new_n14590_, new_n14591_, new_n14592_, new_n14593_, new_n14594_,
    new_n14595_, new_n14596_, new_n14597_, new_n14598_, new_n14599_,
    new_n14600_, new_n14601_, new_n14602_, new_n14603_, new_n14604_,
    new_n14605_, new_n14606_, new_n14607_, new_n14608_, new_n14609_,
    new_n14610_, new_n14611_, new_n14612_, new_n14613_, new_n14614_,
    new_n14615_, new_n14616_, new_n14617_, new_n14618_, new_n14619_,
    new_n14620_, new_n14621_, new_n14622_, new_n14623_, new_n14624_,
    new_n14625_, new_n14626_, new_n14627_, new_n14628_, new_n14629_,
    new_n14630_, new_n14631_, new_n14632_, new_n14633_, new_n14634_,
    new_n14635_, new_n14636_, new_n14637_, new_n14638_, new_n14639_,
    new_n14640_, new_n14641_, new_n14642_, new_n14643_, new_n14644_,
    new_n14645_, new_n14646_, new_n14647_, new_n14648_, new_n14649_,
    new_n14650_, new_n14651_, new_n14652_, new_n14653_, new_n14654_,
    new_n14655_, new_n14656_, new_n14657_, new_n14658_, new_n14660_,
    new_n14661_, new_n14662_, new_n14663_, new_n14664_, new_n14665_,
    new_n14666_, new_n14667_, new_n14668_, new_n14669_, new_n14670_,
    new_n14671_, new_n14672_, new_n14673_, new_n14674_, new_n14675_,
    new_n14676_, new_n14677_, new_n14678_, new_n14679_, new_n14680_,
    new_n14681_, new_n14682_, new_n14683_, new_n14684_, new_n14685_,
    new_n14686_, new_n14687_, new_n14688_, new_n14689_, new_n14690_,
    new_n14691_, new_n14692_, new_n14693_, new_n14694_, new_n14695_,
    new_n14696_, new_n14697_, new_n14698_, new_n14699_, new_n14700_,
    new_n14701_, new_n14702_, new_n14703_, new_n14704_, new_n14705_,
    new_n14706_, new_n14707_, new_n14708_, new_n14709_, new_n14710_,
    new_n14711_, new_n14712_, new_n14713_, new_n14714_, new_n14715_,
    new_n14716_, new_n14717_, new_n14718_, new_n14719_, new_n14720_,
    new_n14721_, new_n14722_, new_n14723_, new_n14724_, new_n14725_,
    new_n14726_, new_n14727_, new_n14728_, new_n14729_, new_n14730_,
    new_n14731_, new_n14732_, new_n14733_, new_n14734_, new_n14735_,
    new_n14736_, new_n14737_, new_n14738_, new_n14739_, new_n14740_,
    new_n14741_, new_n14742_, new_n14743_, new_n14744_, new_n14745_,
    new_n14746_, new_n14747_, new_n14748_, new_n14749_, new_n14750_,
    new_n14751_, new_n14752_, new_n14753_, new_n14754_, new_n14755_,
    new_n14756_, new_n14757_, new_n14758_, new_n14759_, new_n14760_,
    new_n14761_, new_n14762_, new_n14763_, new_n14764_, new_n14765_,
    new_n14766_, new_n14767_, new_n14768_, new_n14769_, new_n14770_,
    new_n14771_, new_n14772_, new_n14773_, new_n14774_, new_n14775_,
    new_n14776_, new_n14777_, new_n14778_, new_n14779_, new_n14780_,
    new_n14781_, new_n14782_, new_n14783_, new_n14784_, new_n14785_,
    new_n14786_, new_n14787_, new_n14788_, new_n14789_, new_n14790_,
    new_n14791_, new_n14792_, new_n14793_, new_n14794_, new_n14795_,
    new_n14796_, new_n14797_, new_n14798_, new_n14799_, new_n14800_,
    new_n14801_, new_n14802_, new_n14803_, new_n14804_, new_n14805_,
    new_n14806_, new_n14807_, new_n14808_, new_n14809_, new_n14810_,
    new_n14811_, new_n14812_, new_n14813_, new_n14815_, new_n14816_,
    new_n14817_, new_n14818_, new_n14819_, new_n14820_, new_n14821_,
    new_n14822_, new_n14823_, new_n14824_, new_n14825_, new_n14826_,
    new_n14827_, new_n14828_, new_n14829_, new_n14830_, new_n14831_,
    new_n14832_, new_n14833_, new_n14834_, new_n14835_, new_n14836_,
    new_n14837_, new_n14838_, new_n14839_, new_n14840_, new_n14841_,
    new_n14842_, new_n14843_, new_n14844_, new_n14845_, new_n14846_,
    new_n14847_, new_n14848_, new_n14849_, new_n14850_, new_n14851_,
    new_n14852_, new_n14853_, new_n14854_, new_n14855_, new_n14856_,
    new_n14857_, new_n14858_, new_n14859_, new_n14860_, new_n14861_,
    new_n14862_, new_n14863_, new_n14864_, new_n14865_, new_n14866_,
    new_n14867_, new_n14868_, new_n14869_, new_n14870_, new_n14871_,
    new_n14872_, new_n14873_, new_n14874_, new_n14875_, new_n14876_,
    new_n14877_, new_n14878_, new_n14879_, new_n14880_, new_n14881_,
    new_n14882_, new_n14883_, new_n14884_, new_n14885_, new_n14886_,
    new_n14887_, new_n14888_, new_n14889_, new_n14890_, new_n14891_,
    new_n14892_, new_n14893_, new_n14894_, new_n14895_, new_n14896_,
    new_n14897_, new_n14898_, new_n14899_, new_n14900_, new_n14901_,
    new_n14902_, new_n14903_, new_n14904_, new_n14905_, new_n14906_,
    new_n14907_, new_n14908_, new_n14909_, new_n14910_, new_n14911_,
    new_n14912_, new_n14913_, new_n14914_, new_n14915_, new_n14916_,
    new_n14917_, new_n14918_, new_n14919_, new_n14920_, new_n14921_,
    new_n14922_, new_n14923_, new_n14924_, new_n14925_, new_n14926_,
    new_n14927_, new_n14928_, new_n14929_, new_n14930_, new_n14931_,
    new_n14932_, new_n14933_, new_n14934_, new_n14935_, new_n14936_,
    new_n14937_, new_n14938_, new_n14939_, new_n14940_, new_n14941_,
    new_n14942_, new_n14943_, new_n14944_, new_n14945_, new_n14946_,
    new_n14947_, new_n14948_, new_n14949_, new_n14950_, new_n14951_,
    new_n14952_, new_n14953_, new_n14954_, new_n14955_, new_n14956_,
    new_n14957_, new_n14959_, new_n14960_, new_n14961_, new_n14962_,
    new_n14963_, new_n14964_, new_n14965_, new_n14966_, new_n14967_,
    new_n14968_, new_n14969_, new_n14970_, new_n14971_, new_n14972_,
    new_n14973_, new_n14974_, new_n14975_, new_n14976_, new_n14977_,
    new_n14978_, new_n14979_, new_n14980_, new_n14981_, new_n14982_,
    new_n14983_, new_n14984_, new_n14985_, new_n14986_, new_n14987_,
    new_n14988_, new_n14989_, new_n14990_, new_n14991_, new_n14992_,
    new_n14993_, new_n14994_, new_n14995_, new_n14996_, new_n14997_,
    new_n14998_, new_n14999_, new_n15000_, new_n15001_, new_n15002_,
    new_n15003_, new_n15004_, new_n15005_, new_n15006_, new_n15007_,
    new_n15008_, new_n15009_, new_n15010_, new_n15011_, new_n15012_,
    new_n15013_, new_n15014_, new_n15015_, new_n15016_, new_n15017_,
    new_n15018_, new_n15019_, new_n15020_, new_n15021_, new_n15022_,
    new_n15023_, new_n15024_, new_n15025_, new_n15026_, new_n15027_,
    new_n15028_, new_n15029_, new_n15030_, new_n15031_, new_n15032_,
    new_n15033_, new_n15034_, new_n15035_, new_n15036_, new_n15037_,
    new_n15038_, new_n15039_, new_n15040_, new_n15041_, new_n15042_,
    new_n15043_, new_n15044_, new_n15045_, new_n15046_, new_n15047_,
    new_n15048_, new_n15049_, new_n15050_, new_n15051_, new_n15052_,
    new_n15053_, new_n15054_, new_n15055_, new_n15056_, new_n15057_,
    new_n15058_, new_n15059_, new_n15060_, new_n15061_, new_n15062_,
    new_n15063_, new_n15064_, new_n15065_, new_n15066_, new_n15067_,
    new_n15068_, new_n15069_, new_n15070_, new_n15071_, new_n15072_,
    new_n15073_, new_n15074_, new_n15075_, new_n15076_, new_n15077_,
    new_n15078_, new_n15079_, new_n15080_, new_n15081_, new_n15082_,
    new_n15083_, new_n15084_, new_n15085_, new_n15086_, new_n15087_,
    new_n15088_, new_n15089_, new_n15090_, new_n15091_, new_n15092_,
    new_n15093_, new_n15094_, new_n15095_, new_n15096_, new_n15097_,
    new_n15098_, new_n15099_, new_n15100_, new_n15101_, new_n15102_,
    new_n15103_, new_n15105_, new_n15106_, new_n15107_, new_n15108_,
    new_n15109_, new_n15110_, new_n15111_, new_n15112_, new_n15113_,
    new_n15114_, new_n15115_, new_n15116_, new_n15117_, new_n15118_,
    new_n15119_, new_n15120_, new_n15121_, new_n15122_, new_n15123_,
    new_n15124_, new_n15125_, new_n15126_, new_n15127_, new_n15128_,
    new_n15129_, new_n15130_, new_n15131_, new_n15132_, new_n15133_,
    new_n15134_, new_n15135_, new_n15136_, new_n15137_, new_n15138_,
    new_n15139_, new_n15140_, new_n15141_, new_n15142_, new_n15143_,
    new_n15144_, new_n15145_, new_n15146_, new_n15147_, new_n15148_,
    new_n15149_, new_n15150_, new_n15151_, new_n15152_, new_n15153_,
    new_n15154_, new_n15155_, new_n15156_, new_n15157_, new_n15158_,
    new_n15159_, new_n15160_, new_n15161_, new_n15162_, new_n15163_,
    new_n15164_, new_n15165_, new_n15166_, new_n15167_, new_n15168_,
    new_n15169_, new_n15170_, new_n15171_, new_n15172_, new_n15173_,
    new_n15174_, new_n15175_, new_n15176_, new_n15177_, new_n15178_,
    new_n15179_, new_n15180_, new_n15181_, new_n15182_, new_n15183_,
    new_n15184_, new_n15185_, new_n15186_, new_n15187_, new_n15188_,
    new_n15189_, new_n15190_, new_n15191_, new_n15192_, new_n15193_,
    new_n15194_, new_n15195_, new_n15196_, new_n15197_, new_n15198_,
    new_n15199_, new_n15200_, new_n15201_, new_n15202_, new_n15203_,
    new_n15204_, new_n15205_, new_n15206_, new_n15207_, new_n15208_,
    new_n15209_, new_n15210_, new_n15211_, new_n15212_, new_n15213_,
    new_n15214_, new_n15215_, new_n15216_, new_n15217_, new_n15218_,
    new_n15219_, new_n15220_, new_n15221_, new_n15222_, new_n15223_,
    new_n15224_, new_n15225_, new_n15226_, new_n15227_, new_n15228_,
    new_n15229_, new_n15230_, new_n15231_, new_n15232_, new_n15233_,
    new_n15234_, new_n15235_, new_n15236_, new_n15237_, new_n15238_,
    new_n15239_, new_n15240_, new_n15241_, new_n15242_, new_n15243_,
    new_n15244_, new_n15245_, new_n15247_, new_n15248_, new_n15249_,
    new_n15250_, new_n15251_, new_n15252_, new_n15253_, new_n15254_,
    new_n15255_, new_n15256_, new_n15257_, new_n15258_, new_n15259_,
    new_n15260_, new_n15261_, new_n15262_, new_n15263_, new_n15264_,
    new_n15265_, new_n15266_, new_n15267_, new_n15268_, new_n15269_,
    new_n15270_, new_n15271_, new_n15272_, new_n15273_, new_n15274_,
    new_n15275_, new_n15276_, new_n15277_, new_n15278_, new_n15279_,
    new_n15280_, new_n15281_, new_n15282_, new_n15283_, new_n15284_,
    new_n15285_, new_n15286_, new_n15287_, new_n15288_, new_n15289_,
    new_n15290_, new_n15291_, new_n15292_, new_n15293_, new_n15294_,
    new_n15295_, new_n15296_, new_n15297_, new_n15298_, new_n15299_,
    new_n15300_, new_n15301_, new_n15302_, new_n15303_, new_n15304_,
    new_n15305_, new_n15306_, new_n15307_, new_n15308_, new_n15309_,
    new_n15310_, new_n15311_, new_n15312_, new_n15313_, new_n15314_,
    new_n15315_, new_n15316_, new_n15317_, new_n15318_, new_n15319_,
    new_n15320_, new_n15321_, new_n15322_, new_n15323_, new_n15324_,
    new_n15325_, new_n15326_, new_n15327_, new_n15328_, new_n15329_,
    new_n15330_, new_n15331_, new_n15332_, new_n15333_, new_n15334_,
    new_n15335_, new_n15336_, new_n15337_, new_n15338_, new_n15339_,
    new_n15340_, new_n15341_, new_n15342_, new_n15343_, new_n15344_,
    new_n15345_, new_n15346_, new_n15347_, new_n15348_, new_n15349_,
    new_n15350_, new_n15351_, new_n15352_, new_n15353_, new_n15354_,
    new_n15355_, new_n15356_, new_n15357_, new_n15358_, new_n15359_,
    new_n15360_, new_n15361_, new_n15362_, new_n15363_, new_n15364_,
    new_n15365_, new_n15366_, new_n15367_, new_n15368_, new_n15369_,
    new_n15370_, new_n15371_, new_n15372_, new_n15373_, new_n15374_,
    new_n15375_, new_n15376_, new_n15377_, new_n15378_, new_n15380_,
    new_n15381_, new_n15382_, new_n15383_, new_n15384_, new_n15385_,
    new_n15386_, new_n15387_, new_n15388_, new_n15389_, new_n15390_,
    new_n15391_, new_n15392_, new_n15393_, new_n15394_, new_n15395_,
    new_n15396_, new_n15397_, new_n15398_, new_n15399_, new_n15400_,
    new_n15401_, new_n15402_, new_n15403_, new_n15404_, new_n15405_,
    new_n15406_, new_n15407_, new_n15408_, new_n15409_, new_n15410_,
    new_n15411_, new_n15412_, new_n15413_, new_n15414_, new_n15415_,
    new_n15416_, new_n15417_, new_n15418_, new_n15419_, new_n15420_,
    new_n15421_, new_n15422_, new_n15423_, new_n15424_, new_n15425_,
    new_n15426_, new_n15427_, new_n15428_, new_n15429_, new_n15430_,
    new_n15431_, new_n15432_, new_n15433_, new_n15434_, new_n15435_,
    new_n15436_, new_n15437_, new_n15438_, new_n15439_, new_n15440_,
    new_n15441_, new_n15442_, new_n15443_, new_n15444_, new_n15445_,
    new_n15446_, new_n15447_, new_n15448_, new_n15449_, new_n15450_,
    new_n15451_, new_n15452_, new_n15453_, new_n15454_, new_n15455_,
    new_n15456_, new_n15457_, new_n15458_, new_n15459_, new_n15460_,
    new_n15461_, new_n15462_, new_n15463_, new_n15464_, new_n15465_,
    new_n15466_, new_n15467_, new_n15468_, new_n15469_, new_n15470_,
    new_n15471_, new_n15472_, new_n15473_, new_n15474_, new_n15475_,
    new_n15476_, new_n15477_, new_n15478_, new_n15479_, new_n15480_,
    new_n15481_, new_n15482_, new_n15483_, new_n15484_, new_n15485_,
    new_n15486_, new_n15487_, new_n15488_, new_n15489_, new_n15490_,
    new_n15491_, new_n15492_, new_n15493_, new_n15494_, new_n15495_,
    new_n15496_, new_n15497_, new_n15498_, new_n15500_, new_n15501_,
    new_n15502_, new_n15503_, new_n15504_, new_n15505_, new_n15506_,
    new_n15507_, new_n15508_, new_n15509_, new_n15510_, new_n15511_,
    new_n15512_, new_n15513_, new_n15514_, new_n15515_, new_n15516_,
    new_n15517_, new_n15518_, new_n15519_, new_n15520_, new_n15521_,
    new_n15522_, new_n15523_, new_n15524_, new_n15525_, new_n15526_,
    new_n15527_, new_n15528_, new_n15529_, new_n15530_, new_n15531_,
    new_n15532_, new_n15533_, new_n15534_, new_n15535_, new_n15536_,
    new_n15537_, new_n15538_, new_n15539_, new_n15540_, new_n15541_,
    new_n15542_, new_n15543_, new_n15544_, new_n15545_, new_n15546_,
    new_n15547_, new_n15548_, new_n15549_, new_n15550_, new_n15551_,
    new_n15552_, new_n15553_, new_n15554_, new_n15555_, new_n15556_,
    new_n15557_, new_n15558_, new_n15559_, new_n15560_, new_n15561_,
    new_n15562_, new_n15563_, new_n15564_, new_n15565_, new_n15566_,
    new_n15567_, new_n15568_, new_n15569_, new_n15570_, new_n15571_,
    new_n15572_, new_n15573_, new_n15574_, new_n15575_, new_n15576_,
    new_n15577_, new_n15578_, new_n15579_, new_n15580_, new_n15581_,
    new_n15582_, new_n15583_, new_n15584_, new_n15585_, new_n15586_,
    new_n15587_, new_n15588_, new_n15589_, new_n15590_, new_n15591_,
    new_n15592_, new_n15593_, new_n15594_, new_n15595_, new_n15596_,
    new_n15597_, new_n15598_, new_n15599_, new_n15600_, new_n15601_,
    new_n15602_, new_n15603_, new_n15604_, new_n15605_, new_n15606_,
    new_n15607_, new_n15608_, new_n15609_, new_n15610_, new_n15611_,
    new_n15612_, new_n15613_, new_n15614_, new_n15615_, new_n15616_,
    new_n15617_, new_n15618_, new_n15619_, new_n15620_, new_n15621_,
    new_n15622_, new_n15623_, new_n15624_, new_n15625_, new_n15626_,
    new_n15627_, new_n15628_, new_n15629_, new_n15630_, new_n15631_,
    new_n15632_, new_n15633_, new_n15634_, new_n15635_, new_n15636_,
    new_n15637_, new_n15638_, new_n15639_, new_n15640_, new_n15641_,
    new_n15642_, new_n15643_, new_n15644_, new_n15645_, new_n15646_,
    new_n15647_, new_n15648_, new_n15649_, new_n15650_, new_n15651_,
    new_n15652_, new_n15653_, new_n15654_, new_n15655_, new_n15656_,
    new_n15657_, new_n15658_, new_n15659_, new_n15660_, new_n15661_,
    new_n15662_, new_n15663_, new_n15664_, new_n15665_, new_n15666_,
    new_n15667_, new_n15668_, new_n15669_, new_n15670_, new_n15671_,
    new_n15672_, new_n15673_, new_n15674_, new_n15675_, new_n15676_,
    new_n15677_, new_n15678_, new_n15679_, new_n15680_, new_n15681_,
    new_n15682_, new_n15683_, new_n15684_, new_n15685_, new_n15686_,
    new_n15687_, new_n15688_, new_n15689_, new_n15690_, new_n15692_,
    new_n15693_, new_n15694_, new_n15695_, new_n15696_, new_n15697_,
    new_n15698_, new_n15699_, new_n15700_, new_n15701_, new_n15702_,
    new_n15703_, new_n15704_, new_n15705_, new_n15706_, new_n15707_,
    new_n15708_, new_n15709_, new_n15710_, new_n15711_, new_n15712_,
    new_n15713_, new_n15714_, new_n15715_, new_n15716_, new_n15717_,
    new_n15718_, new_n15719_, new_n15720_, new_n15721_, new_n15722_,
    new_n15723_, new_n15724_, new_n15725_, new_n15726_, new_n15727_,
    new_n15728_, new_n15729_, new_n15730_, new_n15731_, new_n15732_,
    new_n15733_, new_n15734_, new_n15735_, new_n15736_, new_n15737_,
    new_n15738_, new_n15739_, new_n15740_, new_n15741_, new_n15742_,
    new_n15743_, new_n15744_, new_n15745_, new_n15746_, new_n15747_,
    new_n15748_, new_n15749_, new_n15750_, new_n15751_, new_n15752_,
    new_n15753_, new_n15754_, new_n15755_, new_n15756_, new_n15757_,
    new_n15758_, new_n15759_, new_n15760_, new_n15761_, new_n15762_,
    new_n15763_, new_n15764_, new_n15765_, new_n15766_, new_n15767_,
    new_n15768_, new_n15769_, new_n15770_, new_n15771_, new_n15772_,
    new_n15773_, new_n15774_, new_n15775_, new_n15776_, new_n15777_,
    new_n15778_, new_n15779_, new_n15780_, new_n15781_, new_n15782_,
    new_n15783_, new_n15784_, new_n15785_, new_n15786_, new_n15787_,
    new_n15788_, new_n15789_, new_n15790_, new_n15791_, new_n15792_,
    new_n15793_, new_n15794_, new_n15795_, new_n15796_, new_n15797_,
    new_n15798_, new_n15799_, new_n15800_, new_n15801_, new_n15802_,
    new_n15803_, new_n15804_, new_n15805_, new_n15806_, new_n15807_,
    new_n15808_, new_n15809_, new_n15810_, new_n15811_, new_n15812_,
    new_n15813_, new_n15814_, new_n15815_, new_n15816_, new_n15817_,
    new_n15818_, new_n15819_, new_n15820_, new_n15821_, new_n15822_,
    new_n15823_, new_n15824_, new_n15825_, new_n15826_, new_n15827_,
    new_n15828_, new_n15829_, new_n15830_, new_n15831_, new_n15832_,
    new_n15833_, new_n15834_, new_n15835_, new_n15836_, new_n15837_,
    new_n15838_, new_n15839_, new_n15840_, new_n15841_, new_n15842_,
    new_n15843_, new_n15844_, new_n15845_, new_n15846_, new_n15847_,
    new_n15848_, new_n15849_, new_n15850_, new_n15851_, new_n15852_,
    new_n15853_, new_n15854_, new_n15855_, new_n15856_, new_n15857_,
    new_n15858_, new_n15859_, new_n15860_, new_n15861_, new_n15863_,
    new_n15864_, new_n15865_, new_n15866_, new_n15867_, new_n15868_,
    new_n15869_, new_n15870_, new_n15871_, new_n15872_, new_n15873_,
    new_n15874_, new_n15875_, new_n15876_, new_n15877_, new_n15878_,
    new_n15879_, new_n15880_, new_n15881_, new_n15882_, new_n15883_,
    new_n15884_, new_n15885_, new_n15886_, new_n15887_, new_n15888_,
    new_n15889_, new_n15890_, new_n15891_, new_n15892_, new_n15893_,
    new_n15894_, new_n15895_, new_n15896_, new_n15897_, new_n15898_,
    new_n15899_, new_n15900_, new_n15901_, new_n15902_, new_n15903_,
    new_n15904_, new_n15905_, new_n15906_, new_n15907_, new_n15908_,
    new_n15909_, new_n15910_, new_n15911_, new_n15912_, new_n15913_,
    new_n15914_, new_n15915_, new_n15916_, new_n15917_, new_n15918_,
    new_n15919_, new_n15920_, new_n15921_, new_n15922_, new_n15923_,
    new_n15924_, new_n15925_, new_n15926_, new_n15927_, new_n15928_,
    new_n15929_, new_n15930_, new_n15931_, new_n15932_, new_n15933_,
    new_n15934_, new_n15935_, new_n15936_, new_n15937_, new_n15938_,
    new_n15939_, new_n15940_, new_n15941_, new_n15942_, new_n15943_,
    new_n15944_, new_n15945_, new_n15946_, new_n15947_, new_n15948_,
    new_n15949_, new_n15950_, new_n15951_, new_n15952_, new_n15953_,
    new_n15955_, new_n15956_, new_n15957_, new_n15958_, new_n15959_,
    new_n15960_, new_n15961_, new_n15962_, new_n15963_, new_n15964_,
    new_n15965_, new_n15966_, new_n15967_, new_n15968_, new_n15969_,
    new_n15970_, new_n15971_, new_n15972_, new_n15973_, new_n15974_,
    new_n15975_, new_n15976_, new_n15977_, new_n15978_, new_n15979_,
    new_n15980_, new_n15981_, new_n15982_, new_n15983_, new_n15984_,
    new_n15985_, new_n15986_, new_n15987_, new_n15988_, new_n15989_,
    new_n15990_, new_n15991_, new_n15992_, new_n15993_, new_n15994_,
    new_n15995_, new_n15996_, new_n15997_, new_n15998_, new_n15999_,
    new_n16000_, new_n16001_, new_n16002_, new_n16003_, new_n16004_,
    new_n16005_, new_n16006_, new_n16007_, new_n16008_, new_n16009_,
    new_n16010_, new_n16011_, new_n16012_, new_n16013_, new_n16014_,
    new_n16015_, new_n16016_, new_n16017_, new_n16018_, new_n16019_,
    new_n16020_, new_n16021_, new_n16022_, new_n16023_, new_n16024_,
    new_n16025_, new_n16026_, new_n16027_, new_n16028_, new_n16029_,
    new_n16030_, new_n16031_, new_n16032_, new_n16033_, new_n16034_,
    new_n16035_, new_n16036_, new_n16037_, new_n16038_, new_n16039_,
    new_n16040_, new_n16041_, new_n16042_, new_n16043_, new_n16044_,
    new_n16045_, new_n16046_, new_n16047_, new_n16048_, new_n16049_,
    new_n16050_, new_n16051_, new_n16052_, new_n16053_, new_n16054_,
    new_n16055_, new_n16056_, new_n16057_, new_n16058_, new_n16059_,
    new_n16060_, new_n16061_, new_n16062_, new_n16063_, new_n16064_,
    new_n16065_, new_n16066_, new_n16068_, new_n16069_, new_n16070_,
    new_n16071_, new_n16072_, new_n16073_, new_n16074_, new_n16075_,
    new_n16076_, new_n16077_, new_n16078_, new_n16079_, new_n16080_,
    new_n16081_, new_n16082_, new_n16083_, new_n16084_, new_n16085_,
    new_n16086_, new_n16087_, new_n16088_, new_n16089_, new_n16090_,
    new_n16091_, new_n16092_, new_n16093_, new_n16094_, new_n16095_,
    new_n16096_, new_n16097_, new_n16098_, new_n16099_, new_n16100_,
    new_n16101_, new_n16102_, new_n16103_, new_n16104_, new_n16105_,
    new_n16106_, new_n16107_, new_n16108_, new_n16109_, new_n16110_,
    new_n16111_, new_n16112_, new_n16113_, new_n16114_, new_n16115_,
    new_n16116_, new_n16117_, new_n16118_, new_n16119_, new_n16120_,
    new_n16121_, new_n16122_, new_n16123_, new_n16124_, new_n16125_,
    new_n16126_, new_n16127_, new_n16128_, new_n16129_, new_n16130_,
    new_n16131_, new_n16132_, new_n16133_, new_n16134_, new_n16135_,
    new_n16136_, new_n16137_, new_n16138_, new_n16139_, new_n16140_,
    new_n16141_, new_n16142_, new_n16143_, new_n16144_, new_n16145_,
    new_n16146_, new_n16147_, new_n16148_, new_n16149_, new_n16150_,
    new_n16151_, new_n16152_, new_n16153_, new_n16154_, new_n16155_,
    new_n16156_, new_n16157_, new_n16158_, new_n16159_, new_n16160_,
    new_n16161_, new_n16162_, new_n16163_, new_n16164_, new_n16165_,
    new_n16167_, new_n16168_, new_n16169_, new_n16170_, new_n16171_,
    new_n16172_, new_n16173_, new_n16174_, new_n16175_, new_n16176_,
    new_n16177_, new_n16178_, new_n16179_, new_n16180_, new_n16181_,
    new_n16182_, new_n16183_, new_n16184_, new_n16185_, new_n16186_,
    new_n16187_, new_n16188_, new_n16189_, new_n16190_, new_n16191_,
    new_n16192_, new_n16193_, new_n16194_, new_n16195_, new_n16196_,
    new_n16197_, new_n16198_, new_n16199_, new_n16200_, new_n16201_,
    new_n16202_, new_n16203_, new_n16204_, new_n16205_, new_n16206_,
    new_n16207_, new_n16208_, new_n16209_, new_n16210_, new_n16211_,
    new_n16212_, new_n16213_, new_n16214_, new_n16215_, new_n16216_,
    new_n16217_, new_n16218_, new_n16219_, new_n16220_, new_n16221_,
    new_n16222_, new_n16223_, new_n16224_, new_n16225_, new_n16226_,
    new_n16227_, new_n16228_, new_n16229_, new_n16230_, new_n16231_,
    new_n16232_, new_n16233_, new_n16234_, new_n16235_, new_n16236_,
    new_n16237_, new_n16238_, new_n16239_, new_n16240_, new_n16241_,
    new_n16242_, new_n16243_, new_n16244_, new_n16245_, new_n16246_,
    new_n16247_, new_n16248_, new_n16249_, new_n16250_, new_n16251_,
    new_n16252_, new_n16253_, new_n16254_, new_n16255_, new_n16256_,
    new_n16257_, new_n16258_, new_n16259_, new_n16260_, new_n16261_,
    new_n16262_, new_n16263_, new_n16264_, new_n16265_, new_n16266_,
    new_n16267_, new_n16268_, new_n16269_, new_n16270_, new_n16271_,
    new_n16272_, new_n16273_, new_n16275_, new_n16276_, new_n16277_,
    new_n16278_, new_n16279_, new_n16280_, new_n16281_, new_n16282_,
    new_n16283_, new_n16284_, new_n16285_, new_n16286_, new_n16287_,
    new_n16288_, new_n16289_, new_n16290_, new_n16291_, new_n16292_,
    new_n16293_, new_n16294_, new_n16295_, new_n16296_, new_n16297_,
    new_n16298_, new_n16299_, new_n16300_, new_n16301_, new_n16302_,
    new_n16303_, new_n16304_, new_n16305_, new_n16306_, new_n16307_,
    new_n16308_, new_n16309_, new_n16310_, new_n16311_, new_n16312_,
    new_n16313_, new_n16314_, new_n16315_, new_n16316_, new_n16317_,
    new_n16318_, new_n16319_, new_n16320_, new_n16321_, new_n16322_,
    new_n16323_, new_n16324_, new_n16325_, new_n16326_, new_n16327_,
    new_n16328_, new_n16329_, new_n16330_, new_n16331_, new_n16332_,
    new_n16333_, new_n16334_, new_n16335_, new_n16336_, new_n16337_,
    new_n16338_, new_n16339_, new_n16340_, new_n16341_, new_n16342_,
    new_n16343_, new_n16344_, new_n16345_, new_n16346_, new_n16347_,
    new_n16348_, new_n16349_, new_n16350_, new_n16351_, new_n16352_,
    new_n16353_, new_n16354_, new_n16355_, new_n16356_, new_n16357_,
    new_n16358_, new_n16359_, new_n16360_, new_n16361_, new_n16362_,
    new_n16363_, new_n16364_, new_n16366_, new_n16367_, new_n16368_,
    new_n16369_, new_n16370_, new_n16371_, new_n16372_, new_n16373_,
    new_n16374_, new_n16375_, new_n16376_, new_n16377_, new_n16378_,
    new_n16379_, new_n16380_, new_n16381_, new_n16382_, new_n16383_,
    new_n16384_, new_n16385_, new_n16386_, new_n16387_, new_n16388_,
    new_n16389_, new_n16390_, new_n16391_, new_n16392_, new_n16393_,
    new_n16394_, new_n16395_, new_n16396_, new_n16397_, new_n16398_,
    new_n16399_, new_n16400_, new_n16401_, new_n16402_, new_n16403_,
    new_n16404_, new_n16405_, new_n16406_, new_n16407_, new_n16408_,
    new_n16409_, new_n16410_, new_n16411_, new_n16412_, new_n16413_,
    new_n16414_, new_n16415_, new_n16416_, new_n16417_, new_n16418_,
    new_n16419_, new_n16420_, new_n16421_, new_n16422_, new_n16423_,
    new_n16424_, new_n16425_, new_n16426_, new_n16427_, new_n16428_,
    new_n16429_, new_n16430_, new_n16431_, new_n16432_, new_n16433_,
    new_n16434_, new_n16435_, new_n16436_, new_n16437_, new_n16438_,
    new_n16439_, new_n16440_, new_n16441_, new_n16442_, new_n16443_,
    new_n16444_, new_n16445_, new_n16446_, new_n16447_, new_n16448_,
    new_n16449_, new_n16450_, new_n16451_, new_n16452_, new_n16453_,
    new_n16454_, new_n16455_, new_n16456_, new_n16457_, new_n16458_,
    new_n16459_, new_n16460_, new_n16461_, new_n16462_, new_n16463_,
    new_n16464_, new_n16465_, new_n16466_, new_n16467_, new_n16469_,
    new_n16470_, new_n16471_, new_n16472_, new_n16473_, new_n16474_,
    new_n16475_, new_n16476_, new_n16477_, new_n16478_, new_n16479_,
    new_n16480_, new_n16481_, new_n16482_, new_n16483_, new_n16484_,
    new_n16485_, new_n16486_, new_n16487_, new_n16488_, new_n16489_,
    new_n16490_, new_n16491_, new_n16492_, new_n16493_, new_n16494_,
    new_n16495_, new_n16496_, new_n16497_, new_n16498_, new_n16499_,
    new_n16500_, new_n16501_, new_n16502_, new_n16503_, new_n16504_,
    new_n16505_, new_n16506_, new_n16507_, new_n16508_, new_n16509_,
    new_n16510_, new_n16511_, new_n16512_, new_n16513_, new_n16514_,
    new_n16515_, new_n16516_, new_n16517_, new_n16518_, new_n16519_,
    new_n16520_, new_n16521_, new_n16522_, new_n16523_, new_n16524_,
    new_n16525_, new_n16526_, new_n16527_, new_n16528_, new_n16529_,
    new_n16530_, new_n16531_, new_n16532_, new_n16533_, new_n16534_,
    new_n16535_, new_n16536_, new_n16537_, new_n16538_, new_n16539_,
    new_n16540_, new_n16541_, new_n16542_, new_n16543_, new_n16544_,
    new_n16545_, new_n16546_, new_n16547_, new_n16548_, new_n16549_,
    new_n16550_, new_n16551_, new_n16552_, new_n16553_, new_n16554_,
    new_n16555_, new_n16556_, new_n16557_, new_n16558_, new_n16559_,
    new_n16560_, new_n16561_, new_n16562_, new_n16564_, new_n16565_,
    new_n16566_, new_n16567_, new_n16568_, new_n16569_, new_n16570_,
    new_n16571_, new_n16572_, new_n16573_, new_n16574_, new_n16575_,
    new_n16576_, new_n16577_, new_n16578_, new_n16579_, new_n16580_,
    new_n16581_, new_n16582_, new_n16583_, new_n16584_, new_n16585_,
    new_n16586_, new_n16587_, new_n16588_, new_n16589_, new_n16590_,
    new_n16591_, new_n16592_, new_n16593_, new_n16594_, new_n16595_,
    new_n16596_, new_n16597_, new_n16598_, new_n16599_, new_n16600_,
    new_n16601_, new_n16602_, new_n16603_, new_n16604_, new_n16605_,
    new_n16606_, new_n16607_, new_n16608_, new_n16609_, new_n16610_,
    new_n16611_, new_n16612_, new_n16613_, new_n16614_, new_n16615_,
    new_n16616_, new_n16617_, new_n16618_, new_n16619_, new_n16620_,
    new_n16621_, new_n16622_, new_n16623_, new_n16624_, new_n16625_,
    new_n16626_, new_n16627_, new_n16628_, new_n16629_, new_n16630_,
    new_n16631_, new_n16632_, new_n16633_, new_n16634_, new_n16635_,
    new_n16636_, new_n16637_, new_n16638_, new_n16639_, new_n16640_,
    new_n16641_, new_n16642_, new_n16643_, new_n16644_, new_n16645_,
    new_n16646_, new_n16647_, new_n16648_, new_n16650_, new_n16651_,
    new_n16652_, new_n16653_, new_n16654_, new_n16655_, new_n16656_,
    new_n16657_, new_n16658_, new_n16659_, new_n16660_, new_n16661_,
    new_n16662_, new_n16663_, new_n16664_, new_n16665_, new_n16666_,
    new_n16667_, new_n16668_, new_n16669_, new_n16670_, new_n16671_,
    new_n16672_, new_n16673_, new_n16674_, new_n16675_, new_n16676_,
    new_n16677_, new_n16678_, new_n16679_, new_n16680_, new_n16681_,
    new_n16682_, new_n16683_, new_n16684_, new_n16685_, new_n16686_,
    new_n16687_, new_n16688_, new_n16689_, new_n16690_, new_n16691_,
    new_n16692_, new_n16693_, new_n16694_, new_n16695_, new_n16696_,
    new_n16697_, new_n16698_, new_n16699_, new_n16700_, new_n16701_,
    new_n16702_, new_n16703_, new_n16704_, new_n16705_, new_n16706_,
    new_n16707_, new_n16708_, new_n16709_, new_n16710_, new_n16711_,
    new_n16712_, new_n16713_, new_n16714_, new_n16715_, new_n16716_,
    new_n16717_, new_n16718_, new_n16719_, new_n16720_, new_n16721_,
    new_n16722_, new_n16723_, new_n16724_, new_n16725_, new_n16726_,
    new_n16728_, new_n16729_, new_n16730_, new_n16731_, new_n16732_,
    new_n16733_, new_n16734_, new_n16735_, new_n16736_, new_n16737_,
    new_n16738_, new_n16739_, new_n16740_, new_n16741_, new_n16742_,
    new_n16743_, new_n16744_, new_n16745_, new_n16746_, new_n16747_,
    new_n16748_, new_n16749_, new_n16750_, new_n16751_, new_n16752_,
    new_n16753_, new_n16754_, new_n16755_, new_n16756_, new_n16757_,
    new_n16758_, new_n16759_, new_n16760_, new_n16761_, new_n16762_,
    new_n16763_, new_n16764_, new_n16765_, new_n16766_, new_n16767_,
    new_n16768_, new_n16769_, new_n16770_, new_n16771_, new_n16772_,
    new_n16773_, new_n16774_, new_n16775_, new_n16776_, new_n16777_,
    new_n16778_, new_n16779_, new_n16780_, new_n16781_, new_n16782_,
    new_n16783_, new_n16784_, new_n16785_, new_n16786_, new_n16787_,
    new_n16788_, new_n16789_, new_n16790_, new_n16791_, new_n16792_,
    new_n16793_, new_n16794_, new_n16795_, new_n16796_, new_n16797_,
    new_n16798_, new_n16799_, new_n16800_, new_n16801_, new_n16802_,
    new_n16803_, new_n16804_, new_n16805_, new_n16806_, new_n16807_,
    new_n16809_, new_n16810_, new_n16811_, new_n16812_, new_n16813_,
    new_n16814_, new_n16815_, new_n16816_, new_n16817_, new_n16818_,
    new_n16819_, new_n16820_, new_n16821_, new_n16822_, new_n16823_,
    new_n16824_, new_n16825_, new_n16826_, new_n16827_, new_n16828_,
    new_n16829_, new_n16830_, new_n16831_, new_n16832_, new_n16833_,
    new_n16834_, new_n16835_, new_n16836_, new_n16837_, new_n16838_,
    new_n16839_, new_n16840_, new_n16841_, new_n16842_, new_n16843_,
    new_n16844_, new_n16845_, new_n16846_, new_n16847_, new_n16848_,
    new_n16849_, new_n16850_, new_n16851_, new_n16852_, new_n16853_,
    new_n16854_, new_n16855_, new_n16856_, new_n16857_, new_n16858_,
    new_n16859_, new_n16860_, new_n16861_, new_n16862_, new_n16863_,
    new_n16864_, new_n16865_, new_n16866_, new_n16867_, new_n16868_,
    new_n16869_, new_n16870_, new_n16871_, new_n16872_, new_n16873_,
    new_n16874_, new_n16875_, new_n16876_, new_n16877_, new_n16878_,
    new_n16879_, new_n16880_, new_n16881_, new_n16883_, new_n16884_,
    new_n16885_, new_n16886_, new_n16887_, new_n16888_, new_n16889_,
    new_n16890_, new_n16891_, new_n16892_, new_n16893_, new_n16894_,
    new_n16895_, new_n16896_, new_n16897_, new_n16898_, new_n16899_,
    new_n16900_, new_n16901_, new_n16902_, new_n16903_, new_n16904_,
    new_n16905_, new_n16906_, new_n16907_, new_n16908_, new_n16909_,
    new_n16910_, new_n16911_, new_n16912_, new_n16913_, new_n16914_,
    new_n16915_, new_n16916_, new_n16917_, new_n16918_, new_n16919_,
    new_n16920_, new_n16921_, new_n16922_, new_n16923_, new_n16924_,
    new_n16925_, new_n16926_, new_n16927_, new_n16928_, new_n16929_,
    new_n16930_, new_n16931_, new_n16932_, new_n16933_, new_n16934_,
    new_n16935_, new_n16936_, new_n16937_, new_n16938_, new_n16939_,
    new_n16940_, new_n16941_, new_n16942_, new_n16943_, new_n16944_,
    new_n16945_, new_n16946_, new_n16947_, new_n16948_, new_n16949_,
    new_n16950_, new_n16951_, new_n16952_, new_n16953_, new_n16954_,
    new_n16955_, new_n16956_, new_n16957_, new_n16958_, new_n16959_,
    new_n16960_, new_n16961_, new_n16962_, new_n16963_, new_n16965_,
    new_n16966_, new_n16967_, new_n16968_, new_n16969_, new_n16970_,
    new_n16971_, new_n16972_, new_n16973_, new_n16974_, new_n16975_,
    new_n16976_, new_n16977_, new_n16978_, new_n16979_, new_n16980_,
    new_n16981_, new_n16982_, new_n16983_, new_n16984_, new_n16985_,
    new_n16986_, new_n16987_, new_n16988_, new_n16989_, new_n16990_,
    new_n16991_, new_n16992_, new_n16993_, new_n16994_, new_n16995_,
    new_n16996_, new_n16997_, new_n16998_, new_n16999_, new_n17000_,
    new_n17001_, new_n17002_, new_n17003_, new_n17004_, new_n17005_,
    new_n17006_, new_n17007_, new_n17008_, new_n17009_, new_n17010_,
    new_n17011_, new_n17012_, new_n17013_, new_n17014_, new_n17015_,
    new_n17016_, new_n17017_, new_n17018_, new_n17019_, new_n17020_,
    new_n17021_, new_n17022_, new_n17023_, new_n17024_, new_n17025_,
    new_n17026_, new_n17027_, new_n17028_, new_n17029_, new_n17030_,
    new_n17031_, new_n17032_, new_n17033_, new_n17034_, new_n17035_,
    new_n17036_, new_n17037_, new_n17038_, new_n17039_, new_n17040_,
    new_n17042_, new_n17043_, new_n17044_, new_n17045_, new_n17046_,
    new_n17047_, new_n17048_, new_n17049_, new_n17050_, new_n17051_,
    new_n17052_, new_n17053_, new_n17054_, new_n17055_, new_n17056_,
    new_n17057_, new_n17058_, new_n17059_, new_n17060_, new_n17061_,
    new_n17062_, new_n17063_, new_n17064_, new_n17065_, new_n17066_,
    new_n17067_, new_n17068_, new_n17069_, new_n17070_, new_n17071_,
    new_n17072_, new_n17073_, new_n17074_, new_n17075_, new_n17076_,
    new_n17077_, new_n17078_, new_n17079_, new_n17080_, new_n17081_,
    new_n17082_, new_n17083_, new_n17084_, new_n17085_, new_n17086_,
    new_n17087_, new_n17088_, new_n17089_, new_n17090_, new_n17091_,
    new_n17092_, new_n17093_, new_n17094_, new_n17095_, new_n17096_,
    new_n17097_, new_n17098_, new_n17099_, new_n17100_, new_n17101_,
    new_n17102_, new_n17103_, new_n17104_, new_n17105_, new_n17107_,
    new_n17108_, new_n17109_, new_n17110_, new_n17111_, new_n17112_,
    new_n17113_, new_n17114_, new_n17115_, new_n17116_, new_n17117_,
    new_n17118_, new_n17119_, new_n17120_, new_n17121_, new_n17122_,
    new_n17123_, new_n17124_, new_n17125_, new_n17126_, new_n17127_,
    new_n17128_, new_n17129_, new_n17130_, new_n17131_, new_n17132_,
    new_n17133_, new_n17134_, new_n17135_, new_n17136_, new_n17137_,
    new_n17138_, new_n17139_, new_n17140_, new_n17141_, new_n17142_,
    new_n17143_, new_n17144_, new_n17145_, new_n17146_, new_n17147_,
    new_n17148_, new_n17149_, new_n17150_, new_n17151_, new_n17152_,
    new_n17153_, new_n17154_, new_n17155_, new_n17156_, new_n17157_,
    new_n17158_, new_n17159_, new_n17160_, new_n17161_, new_n17162_,
    new_n17163_, new_n17164_, new_n17165_, new_n17166_, new_n17167_,
    new_n17169_, new_n17170_, new_n17171_, new_n17172_, new_n17173_,
    new_n17174_, new_n17175_, new_n17176_, new_n17177_, new_n17178_,
    new_n17179_, new_n17180_, new_n17181_, new_n17182_, new_n17183_,
    new_n17184_, new_n17185_, new_n17186_, new_n17187_, new_n17188_,
    new_n17189_, new_n17190_, new_n17191_, new_n17192_, new_n17193_,
    new_n17194_, new_n17195_, new_n17196_, new_n17197_, new_n17198_,
    new_n17199_, new_n17200_, new_n17201_, new_n17202_, new_n17203_,
    new_n17204_, new_n17205_, new_n17206_, new_n17207_, new_n17208_,
    new_n17209_, new_n17210_, new_n17211_, new_n17212_, new_n17213_,
    new_n17214_, new_n17215_, new_n17216_, new_n17217_, new_n17218_,
    new_n17219_, new_n17220_, new_n17221_, new_n17222_, new_n17223_,
    new_n17224_, new_n17225_, new_n17226_, new_n17227_, new_n17228_,
    new_n17230_, new_n17231_, new_n17232_, new_n17233_, new_n17234_,
    new_n17235_, new_n17236_, new_n17237_, new_n17238_, new_n17239_,
    new_n17240_, new_n17241_, new_n17242_, new_n17243_, new_n17244_,
    new_n17245_, new_n17246_, new_n17247_, new_n17248_, new_n17249_,
    new_n17250_, new_n17251_, new_n17252_, new_n17253_, new_n17254_,
    new_n17255_, new_n17256_, new_n17257_, new_n17258_, new_n17259_,
    new_n17260_, new_n17261_, new_n17262_, new_n17263_, new_n17264_,
    new_n17265_, new_n17266_, new_n17267_, new_n17268_, new_n17269_,
    new_n17270_, new_n17271_, new_n17272_, new_n17273_, new_n17274_,
    new_n17275_, new_n17276_, new_n17277_, new_n17278_, new_n17279_,
    new_n17280_, new_n17281_, new_n17282_, new_n17283_, new_n17284_,
    new_n17285_, new_n17286_, new_n17287_, new_n17288_, new_n17289_,
    new_n17291_, new_n17292_, new_n17293_, new_n17294_, new_n17295_,
    new_n17296_, new_n17297_, new_n17298_, new_n17299_, new_n17300_,
    new_n17301_, new_n17302_, new_n17303_, new_n17304_, new_n17305_,
    new_n17306_, new_n17307_, new_n17308_, new_n17309_, new_n17310_,
    new_n17311_, new_n17312_, new_n17313_, new_n17314_, new_n17315_,
    new_n17316_, new_n17317_, new_n17318_, new_n17319_, new_n17320_,
    new_n17321_, new_n17322_, new_n17323_, new_n17324_, new_n17325_,
    new_n17326_, new_n17327_, new_n17328_, new_n17329_, new_n17330_,
    new_n17331_, new_n17332_, new_n17333_, new_n17334_, new_n17335_,
    new_n17336_, new_n17337_, new_n17338_, new_n17339_, new_n17340_,
    new_n17341_, new_n17342_, new_n17343_, new_n17344_, new_n17346_,
    new_n17347_, new_n17348_, new_n17349_, new_n17350_, new_n17351_,
    new_n17352_, new_n17353_, new_n17354_, new_n17355_, new_n17356_,
    new_n17357_, new_n17358_, new_n17359_, new_n17360_, new_n17361_,
    new_n17362_, new_n17363_, new_n17364_, new_n17365_, new_n17366_,
    new_n17367_, new_n17368_, new_n17369_, new_n17370_, new_n17371_,
    new_n17372_, new_n17373_, new_n17374_, new_n17375_, new_n17376_,
    new_n17377_, new_n17378_, new_n17379_, new_n17380_, new_n17381_,
    new_n17382_, new_n17383_, new_n17384_, new_n17385_, new_n17386_,
    new_n17387_, new_n17388_, new_n17389_, new_n17390_, new_n17391_,
    new_n17392_, new_n17393_, new_n17394_, new_n17395_, new_n17396_,
    new_n17397_, new_n17399_, new_n17400_, new_n17401_, new_n17402_,
    new_n17403_, new_n17404_, new_n17405_, new_n17406_, new_n17407_,
    new_n17408_, new_n17409_, new_n17410_, new_n17411_, new_n17412_,
    new_n17413_, new_n17414_, new_n17415_, new_n17416_, new_n17417_,
    new_n17418_, new_n17419_, new_n17420_, new_n17421_, new_n17422_,
    new_n17423_, new_n17424_, new_n17425_, new_n17426_, new_n17427_,
    new_n17428_, new_n17429_, new_n17430_, new_n17431_, new_n17432_,
    new_n17433_, new_n17434_, new_n17435_, new_n17436_, new_n17437_,
    new_n17438_, new_n17439_, new_n17440_, new_n17442_, new_n17443_,
    new_n17444_, new_n17445_, new_n17446_, new_n17447_, new_n17448_,
    new_n17449_, new_n17450_, new_n17451_, new_n17452_, new_n17453_,
    new_n17454_, new_n17455_, new_n17456_, new_n17457_, new_n17458_,
    new_n17459_, new_n17460_, new_n17461_, new_n17462_, new_n17463_,
    new_n17464_, new_n17465_, new_n17466_, new_n17467_, new_n17468_,
    new_n17469_, new_n17470_, new_n17471_, new_n17472_, new_n17473_,
    new_n17474_, new_n17475_, new_n17476_, new_n17477_, new_n17478_,
    new_n17479_, new_n17480_, new_n17481_, new_n17482_, new_n17483_,
    new_n17485_, new_n17486_, new_n17487_, new_n17488_, new_n17489_,
    new_n17490_, new_n17491_, new_n17492_, new_n17493_, new_n17494_,
    new_n17495_, new_n17496_, new_n17497_, new_n17498_, new_n17499_,
    new_n17500_, new_n17501_, new_n17502_, new_n17503_, new_n17504_,
    new_n17505_, new_n17506_, new_n17507_, new_n17508_, new_n17509_,
    new_n17510_, new_n17511_, new_n17512_, new_n17513_, new_n17514_,
    new_n17515_, new_n17516_, new_n17517_, new_n17518_, new_n17519_,
    new_n17520_, new_n17521_, new_n17522_, new_n17523_, new_n17524_,
    new_n17525_, new_n17526_, new_n17528_, new_n17529_, new_n17530_,
    new_n17531_, new_n17532_, new_n17533_, new_n17534_, new_n17535_,
    new_n17536_, new_n17537_, new_n17538_, new_n17539_, new_n17540_,
    new_n17541_, new_n17542_, new_n17543_, new_n17544_, new_n17545_,
    new_n17546_, new_n17547_, new_n17548_, new_n17549_, new_n17550_,
    new_n17551_, new_n17552_;
  XOR2X1   g00000(.A(\a[5] ), .B(\a[4] ), .Y(new_n65_));
  XOR2X1   g00001(.A(\a[3] ), .B(\a[2] ), .Y(new_n66_));
  AND2X1   g00002(.A(new_n66_), .B(new_n65_), .Y(new_n67_));
  INVX1    g00003(.A(\a[30] ), .Y(new_n68_));
  OR4X1    g00004(.A(new_n68_), .B(\a[29] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n69_));
  INVX1    g00005(.A(\a[23] ), .Y(new_n70_));
  INVX1    g00006(.A(\a[24] ), .Y(new_n71_));
  OR4X1    g00007(.A(\a[26] ), .B(\a[25] ), .C(new_n71_), .D(new_n70_), .Y(new_n72_));
  INVX1    g00008(.A(\a[27] ), .Y(new_n73_));
  INVX1    g00009(.A(\a[29] ), .Y(new_n74_));
  OR4X1    g00010(.A(\a[30] ), .B(new_n74_), .C(\a[28] ), .D(new_n73_), .Y(new_n75_));
  AOI21X1  g00011(.A0(new_n75_), .A1(new_n69_), .B0(new_n72_), .Y(new_n76_));
  INVX1    g00012(.A(\a[25] ), .Y(new_n77_));
  OR4X1    g00013(.A(\a[26] ), .B(new_n77_), .C(\a[24] ), .D(new_n70_), .Y(new_n78_));
  OR4X1    g00014(.A(\a[30] ), .B(new_n74_), .C(\a[28] ), .D(\a[27] ), .Y(new_n79_));
  NOR2X1   g00015(.A(new_n79_), .B(new_n78_), .Y(new_n80_));
  OR4X1    g00016(.A(\a[26] ), .B(\a[25] ), .C(new_n71_), .D(\a[23] ), .Y(new_n81_));
  AND2X1   g00017(.A(\a[28] ), .B(\a[27] ), .Y(new_n82_));
  NOR2X1   g00018(.A(\a[30] ), .B(\a[29] ), .Y(new_n83_));
  NAND2X1  g00019(.A(new_n83_), .B(new_n82_), .Y(new_n84_));
  NOR2X1   g00020(.A(new_n84_), .B(new_n81_), .Y(new_n85_));
  NOR2X1   g00021(.A(new_n81_), .B(new_n69_), .Y(new_n86_));
  OR4X1    g00022(.A(new_n86_), .B(new_n85_), .C(new_n80_), .D(new_n76_), .Y(new_n87_));
  NAND3X1  g00023(.A(new_n83_), .B(\a[28] ), .C(new_n73_), .Y(new_n88_));
  INVX1    g00024(.A(\a[26] ), .Y(new_n89_));
  OR4X1    g00025(.A(new_n89_), .B(new_n77_), .C(\a[24] ), .D(\a[23] ), .Y(new_n90_));
  NAND3X1  g00026(.A(new_n82_), .B(new_n68_), .C(\a[29] ), .Y(new_n91_));
  OR4X1    g00027(.A(new_n89_), .B(\a[25] ), .C(new_n71_), .D(\a[23] ), .Y(new_n92_));
  OAI22X1  g00028(.A0(new_n92_), .A1(new_n91_), .B0(new_n90_), .B1(new_n88_), .Y(new_n93_));
  OR4X1    g00029(.A(new_n89_), .B(\a[25] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n94_));
  INVX1    g00030(.A(\a[28] ), .Y(new_n95_));
  OR4X1    g00031(.A(\a[30] ), .B(new_n74_), .C(new_n95_), .D(\a[27] ), .Y(new_n96_));
  OAI22X1  g00032(.A0(new_n96_), .A1(new_n92_), .B0(new_n94_), .B1(new_n91_), .Y(new_n97_));
  OR2X1    g00033(.A(\a[28] ), .B(\a[27] ), .Y(new_n98_));
  OR4X1    g00034(.A(\a[26] ), .B(\a[25] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n99_));
  NOR4X1   g00035(.A(new_n99_), .B(new_n98_), .C(new_n68_), .D(new_n74_), .Y(new_n100_));
  OR2X1    g00036(.A(\a[25] ), .B(\a[24] ), .Y(new_n101_));
  OR4X1    g00037(.A(\a[30] ), .B(\a[29] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n102_));
  NOR4X1   g00038(.A(new_n102_), .B(new_n101_), .C(new_n89_), .D(\a[23] ), .Y(new_n103_));
  OR2X1    g00039(.A(new_n103_), .B(new_n100_), .Y(new_n104_));
  OR4X1    g00040(.A(\a[26] ), .B(new_n77_), .C(new_n71_), .D(new_n70_), .Y(new_n105_));
  NAND3X1  g00041(.A(new_n82_), .B(\a[30] ), .C(new_n74_), .Y(new_n106_));
  NAND2X1  g00042(.A(\a[26] ), .B(\a[23] ), .Y(new_n107_));
  OR2X1    g00043(.A(new_n107_), .B(new_n101_), .Y(new_n108_));
  OAI22X1  g00044(.A0(new_n108_), .A1(new_n106_), .B0(new_n105_), .B1(new_n88_), .Y(new_n109_));
  OR4X1    g00045(.A(new_n109_), .B(new_n104_), .C(new_n97_), .D(new_n93_), .Y(new_n110_));
  NOR2X1   g00046(.A(new_n102_), .B(new_n90_), .Y(new_n111_));
  OAI22X1  g00047(.A0(new_n92_), .A1(new_n84_), .B0(new_n88_), .B1(new_n81_), .Y(new_n112_));
  OR2X1    g00048(.A(new_n112_), .B(new_n111_), .Y(new_n113_));
  NOR2X1   g00049(.A(new_n99_), .B(new_n75_), .Y(new_n114_));
  OR4X1    g00050(.A(new_n68_), .B(new_n74_), .C(\a[28] ), .D(\a[27] ), .Y(new_n115_));
  NOR2X1   g00051(.A(new_n108_), .B(new_n115_), .Y(new_n116_));
  OR4X1    g00052(.A(new_n68_), .B(new_n74_), .C(new_n95_), .D(\a[27] ), .Y(new_n117_));
  NOR2X1   g00053(.A(new_n117_), .B(new_n108_), .Y(new_n118_));
  OR4X1    g00054(.A(new_n68_), .B(\a[29] ), .C(\a[28] ), .D(new_n73_), .Y(new_n119_));
  NOR2X1   g00055(.A(new_n119_), .B(new_n72_), .Y(new_n120_));
  OR4X1    g00056(.A(new_n120_), .B(new_n118_), .C(new_n116_), .D(new_n114_), .Y(new_n121_));
  OR4X1    g00057(.A(new_n121_), .B(new_n113_), .C(new_n110_), .D(new_n87_), .Y(new_n122_));
  NAND3X1  g00058(.A(new_n83_), .B(new_n95_), .C(\a[27] ), .Y(new_n123_));
  NOR2X1   g00059(.A(new_n123_), .B(new_n81_), .Y(new_n124_));
  NAND4X1  g00060(.A(\a[26] ), .B(\a[25] ), .C(\a[24] ), .D(\a[23] ), .Y(new_n125_));
  NOR4X1   g00061(.A(new_n125_), .B(new_n98_), .C(new_n68_), .D(new_n74_), .Y(new_n126_));
  OR4X1    g00062(.A(new_n89_), .B(new_n77_), .C(\a[24] ), .D(new_n70_), .Y(new_n127_));
  OAI22X1  g00063(.A0(new_n127_), .A1(new_n117_), .B0(new_n106_), .B1(new_n99_), .Y(new_n128_));
  OR4X1    g00064(.A(\a[26] ), .B(\a[25] ), .C(\a[24] ), .D(new_n70_), .Y(new_n129_));
  OAI22X1  g00065(.A0(new_n129_), .A1(new_n106_), .B0(new_n127_), .B1(new_n88_), .Y(new_n130_));
  OR4X1    g00066(.A(new_n89_), .B(\a[25] ), .C(new_n71_), .D(new_n70_), .Y(new_n131_));
  OAI22X1  g00067(.A0(new_n131_), .A1(new_n102_), .B0(new_n119_), .B1(new_n94_), .Y(new_n132_));
  NOR2X1   g00068(.A(new_n131_), .B(new_n96_), .Y(new_n133_));
  NOR2X1   g00069(.A(new_n96_), .B(new_n72_), .Y(new_n134_));
  OR4X1    g00070(.A(new_n134_), .B(new_n133_), .C(new_n132_), .D(new_n130_), .Y(new_n135_));
  OR4X1    g00071(.A(new_n135_), .B(new_n128_), .C(new_n126_), .D(new_n124_), .Y(new_n136_));
  NOR2X1   g00072(.A(new_n117_), .B(new_n90_), .Y(new_n137_));
  NOR2X1   g00073(.A(new_n123_), .B(new_n99_), .Y(new_n138_));
  NOR2X1   g00074(.A(new_n119_), .B(new_n78_), .Y(new_n139_));
  NOR3X1   g00075(.A(new_n139_), .B(new_n138_), .C(new_n137_), .Y(new_n140_));
  NOR2X1   g00076(.A(new_n102_), .B(new_n81_), .Y(new_n141_));
  NOR2X1   g00077(.A(new_n125_), .B(new_n96_), .Y(new_n142_));
  OR4X1    g00078(.A(new_n89_), .B(new_n77_), .C(new_n71_), .D(\a[23] ), .Y(new_n143_));
  NOR2X1   g00079(.A(new_n143_), .B(new_n106_), .Y(new_n144_));
  NOR3X1   g00080(.A(new_n144_), .B(new_n142_), .C(new_n141_), .Y(new_n145_));
  OAI22X1  g00081(.A0(new_n117_), .A1(new_n81_), .B0(new_n115_), .B1(new_n78_), .Y(new_n146_));
  NOR2X1   g00082(.A(new_n131_), .B(new_n119_), .Y(new_n147_));
  OR4X1    g00083(.A(new_n68_), .B(\a[29] ), .C(new_n95_), .D(\a[27] ), .Y(new_n148_));
  NOR2X1   g00084(.A(new_n148_), .B(new_n125_), .Y(new_n149_));
  NOR3X1   g00085(.A(new_n149_), .B(new_n147_), .C(new_n146_), .Y(new_n150_));
  NAND3X1  g00086(.A(new_n150_), .B(new_n145_), .C(new_n140_), .Y(new_n151_));
  OR4X1    g00087(.A(new_n68_), .B(new_n74_), .C(\a[28] ), .D(new_n73_), .Y(new_n152_));
  OAI22X1  g00088(.A0(new_n152_), .A1(new_n143_), .B0(new_n125_), .B1(new_n84_), .Y(new_n153_));
  AOI21X1  g00089(.A0(new_n92_), .A1(new_n90_), .B0(new_n152_), .Y(new_n154_));
  NOR2X1   g00090(.A(new_n84_), .B(new_n78_), .Y(new_n155_));
  NOR2X1   g00091(.A(new_n131_), .B(new_n115_), .Y(new_n156_));
  OR4X1    g00092(.A(new_n156_), .B(new_n155_), .C(new_n154_), .D(new_n153_), .Y(new_n157_));
  NOR2X1   g00093(.A(new_n91_), .B(new_n78_), .Y(new_n158_));
  NOR2X1   g00094(.A(new_n105_), .B(new_n91_), .Y(new_n159_));
  NOR2X1   g00095(.A(new_n108_), .B(new_n84_), .Y(new_n160_));
  OR4X1    g00096(.A(\a[26] ), .B(new_n77_), .C(\a[24] ), .D(\a[23] ), .Y(new_n161_));
  NOR2X1   g00097(.A(new_n161_), .B(new_n84_), .Y(new_n162_));
  OR4X1    g00098(.A(new_n162_), .B(new_n160_), .C(new_n159_), .D(new_n158_), .Y(new_n163_));
  OAI22X1  g00099(.A0(new_n161_), .A1(new_n106_), .B0(new_n125_), .B1(new_n75_), .Y(new_n164_));
  OAI22X1  g00100(.A0(new_n96_), .A1(new_n78_), .B0(new_n90_), .B1(new_n69_), .Y(new_n165_));
  OR4X1    g00101(.A(new_n165_), .B(new_n164_), .C(new_n163_), .D(new_n157_), .Y(new_n166_));
  OR4X1    g00102(.A(new_n166_), .B(new_n151_), .C(new_n136_), .D(new_n122_), .Y(new_n167_));
  NAND4X1  g00103(.A(\a[30] ), .B(\a[29] ), .C(\a[28] ), .D(\a[27] ), .Y(new_n168_));
  OAI22X1  g00104(.A0(new_n168_), .A1(new_n90_), .B0(new_n143_), .B1(new_n119_), .Y(new_n169_));
  OAI22X1  g00105(.A0(new_n127_), .A1(new_n119_), .B0(new_n90_), .B1(new_n75_), .Y(new_n170_));
  OR2X1    g00106(.A(new_n143_), .B(new_n79_), .Y(new_n171_));
  INVX1    g00107(.A(new_n171_), .Y(new_n172_));
  NOR2X1   g00108(.A(new_n168_), .B(new_n72_), .Y(new_n173_));
  NOR4X1   g00109(.A(new_n173_), .B(new_n172_), .C(new_n170_), .D(new_n169_), .Y(new_n174_));
  NOR2X1   g00110(.A(new_n108_), .B(new_n91_), .Y(new_n175_));
  NOR2X1   g00111(.A(new_n88_), .B(new_n78_), .Y(new_n176_));
  NOR2X1   g00112(.A(new_n148_), .B(new_n81_), .Y(new_n177_));
  NOR2X1   g00113(.A(new_n106_), .B(new_n105_), .Y(new_n178_));
  NOR4X1   g00114(.A(new_n178_), .B(new_n177_), .C(new_n176_), .D(new_n175_), .Y(new_n179_));
  NOR2X1   g00115(.A(new_n115_), .B(new_n94_), .Y(new_n180_));
  NOR2X1   g00116(.A(new_n125_), .B(new_n117_), .Y(new_n181_));
  OR4X1    g00117(.A(\a[26] ), .B(new_n77_), .C(new_n71_), .D(\a[23] ), .Y(new_n182_));
  NOR2X1   g00118(.A(new_n182_), .B(new_n106_), .Y(new_n183_));
  NOR2X1   g00119(.A(new_n148_), .B(new_n105_), .Y(new_n184_));
  NOR4X1   g00120(.A(new_n184_), .B(new_n183_), .C(new_n181_), .D(new_n180_), .Y(new_n185_));
  NAND3X1  g00121(.A(new_n185_), .B(new_n179_), .C(new_n174_), .Y(new_n186_));
  NOR4X1   g00122(.A(new_n107_), .B(new_n102_), .C(new_n77_), .D(\a[24] ), .Y(new_n187_));
  OAI22X1  g00123(.A0(new_n182_), .A1(new_n148_), .B0(new_n94_), .B1(new_n75_), .Y(new_n188_));
  OR2X1    g00124(.A(new_n188_), .B(new_n187_), .Y(new_n189_));
  OAI22X1  g00125(.A0(new_n168_), .A1(new_n131_), .B0(new_n123_), .B1(new_n105_), .Y(new_n190_));
  NOR2X1   g00126(.A(new_n148_), .B(new_n131_), .Y(new_n191_));
  OR2X1    g00127(.A(new_n108_), .B(new_n79_), .Y(new_n192_));
  INVX1    g00128(.A(new_n192_), .Y(new_n193_));
  NOR2X1   g00129(.A(new_n79_), .B(new_n72_), .Y(new_n194_));
  OR4X1    g00130(.A(new_n194_), .B(new_n193_), .C(new_n191_), .D(new_n190_), .Y(new_n195_));
  NOR2X1   g00131(.A(new_n143_), .B(new_n115_), .Y(new_n196_));
  NOR2X1   g00132(.A(new_n127_), .B(new_n84_), .Y(new_n197_));
  NAND2X1  g00133(.A(\a[25] ), .B(\a[24] ), .Y(new_n198_));
  NOR4X1   g00134(.A(new_n168_), .B(new_n198_), .C(\a[26] ), .D(\a[23] ), .Y(new_n199_));
  NOR2X1   g00135(.A(new_n123_), .B(new_n90_), .Y(new_n200_));
  NOR2X1   g00136(.A(new_n117_), .B(new_n105_), .Y(new_n201_));
  NOR4X1   g00137(.A(new_n125_), .B(new_n98_), .C(\a[30] ), .D(new_n74_), .Y(new_n202_));
  NOR3X1   g00138(.A(new_n107_), .B(new_n102_), .C(new_n101_), .Y(new_n203_));
  OR4X1    g00139(.A(new_n203_), .B(new_n202_), .C(new_n201_), .D(new_n200_), .Y(new_n204_));
  OR4X1    g00140(.A(new_n204_), .B(new_n199_), .C(new_n197_), .D(new_n196_), .Y(new_n205_));
  NOR4X1   g00141(.A(new_n198_), .B(new_n102_), .C(\a[26] ), .D(new_n70_), .Y(new_n206_));
  NOR2X1   g00142(.A(new_n108_), .B(new_n75_), .Y(new_n207_));
  NOR2X1   g00143(.A(new_n148_), .B(new_n90_), .Y(new_n208_));
  AOI21X1  g00144(.A0(new_n182_), .A1(new_n129_), .B0(new_n69_), .Y(new_n209_));
  OR4X1    g00145(.A(new_n209_), .B(new_n208_), .C(new_n207_), .D(new_n206_), .Y(new_n210_));
  OR4X1    g00146(.A(new_n210_), .B(new_n205_), .C(new_n195_), .D(new_n189_), .Y(new_n211_));
  OR2X1    g00147(.A(new_n211_), .B(new_n186_), .Y(new_n212_));
  NOR2X1   g00148(.A(new_n143_), .B(new_n75_), .Y(new_n213_));
  OR4X1    g00149(.A(new_n168_), .B(new_n198_), .C(\a[26] ), .D(new_n70_), .Y(new_n214_));
  OAI21X1  g00150(.A0(new_n161_), .A1(new_n117_), .B0(new_n214_), .Y(new_n215_));
  OR2X1    g00151(.A(new_n215_), .B(new_n213_), .Y(new_n216_));
  NOR2X1   g00152(.A(new_n168_), .B(new_n99_), .Y(new_n217_));
  NOR2X1   g00153(.A(new_n152_), .B(new_n129_), .Y(new_n218_));
  NOR2X1   g00154(.A(new_n182_), .B(new_n119_), .Y(new_n219_));
  NOR2X1   g00155(.A(new_n106_), .B(new_n78_), .Y(new_n220_));
  OR4X1    g00156(.A(new_n220_), .B(new_n219_), .C(new_n218_), .D(new_n217_), .Y(new_n221_));
  OAI22X1  g00157(.A0(new_n182_), .A1(new_n91_), .B0(new_n148_), .B1(new_n78_), .Y(new_n222_));
  NOR2X1   g00158(.A(new_n105_), .B(new_n75_), .Y(new_n223_));
  NOR2X1   g00159(.A(new_n84_), .B(new_n72_), .Y(new_n224_));
  OR4X1    g00160(.A(new_n224_), .B(new_n223_), .C(new_n222_), .D(new_n221_), .Y(new_n225_));
  NOR2X1   g00161(.A(new_n117_), .B(new_n92_), .Y(new_n226_));
  NOR2X1   g00162(.A(new_n106_), .B(new_n81_), .Y(new_n227_));
  NOR2X1   g00163(.A(new_n148_), .B(new_n129_), .Y(new_n228_));
  NOR2X1   g00164(.A(new_n125_), .B(new_n106_), .Y(new_n229_));
  OR4X1    g00165(.A(new_n229_), .B(new_n228_), .C(new_n227_), .D(new_n226_), .Y(new_n230_));
  NOR2X1   g00166(.A(new_n129_), .B(new_n88_), .Y(new_n231_));
  NOR2X1   g00167(.A(new_n102_), .B(new_n92_), .Y(new_n232_));
  NOR2X1   g00168(.A(new_n161_), .B(new_n102_), .Y(new_n233_));
  NOR2X1   g00169(.A(new_n152_), .B(new_n94_), .Y(new_n234_));
  OR4X1    g00170(.A(new_n234_), .B(new_n233_), .C(new_n232_), .D(new_n231_), .Y(new_n235_));
  OR2X1    g00171(.A(new_n235_), .B(new_n230_), .Y(new_n236_));
  OAI22X1  g00172(.A0(new_n182_), .A1(new_n152_), .B0(new_n148_), .B1(new_n143_), .Y(new_n237_));
  OAI22X1  g00173(.A0(new_n161_), .A1(new_n123_), .B0(new_n129_), .B1(new_n79_), .Y(new_n238_));
  NOR2X1   g00174(.A(new_n117_), .B(new_n99_), .Y(new_n239_));
  NOR2X1   g00175(.A(new_n161_), .B(new_n115_), .Y(new_n240_));
  OR4X1    g00176(.A(new_n240_), .B(new_n239_), .C(new_n238_), .D(new_n237_), .Y(new_n241_));
  OR4X1    g00177(.A(new_n241_), .B(new_n236_), .C(new_n225_), .D(new_n216_), .Y(new_n242_));
  NOR2X1   g00178(.A(new_n94_), .B(new_n79_), .Y(new_n243_));
  OR2X1    g00179(.A(new_n81_), .B(new_n75_), .Y(new_n244_));
  INVX1    g00180(.A(new_n244_), .Y(new_n245_));
  NOR2X1   g00181(.A(new_n161_), .B(new_n152_), .Y(new_n246_));
  NOR2X1   g00182(.A(new_n115_), .B(new_n90_), .Y(new_n247_));
  NOR4X1   g00183(.A(new_n247_), .B(new_n246_), .C(new_n245_), .D(new_n243_), .Y(new_n248_));
  OAI22X1  g00184(.A0(new_n182_), .A1(new_n123_), .B0(new_n129_), .B1(new_n96_), .Y(new_n249_));
  OR2X1    g00185(.A(new_n91_), .B(new_n90_), .Y(new_n250_));
  INVX1    g00186(.A(new_n250_), .Y(new_n251_));
  NOR2X1   g00187(.A(new_n161_), .B(new_n91_), .Y(new_n252_));
  NOR3X1   g00188(.A(new_n252_), .B(new_n251_), .C(new_n249_), .Y(new_n253_));
  OAI22X1  g00189(.A0(new_n168_), .A1(new_n81_), .B0(new_n106_), .B1(new_n94_), .Y(new_n254_));
  OAI22X1  g00190(.A0(new_n129_), .A1(new_n75_), .B0(new_n108_), .B1(new_n88_), .Y(new_n255_));
  NOR2X1   g00191(.A(new_n119_), .B(new_n92_), .Y(new_n256_));
  OAI22X1  g00192(.A0(new_n131_), .A1(new_n91_), .B0(new_n129_), .B1(new_n84_), .Y(new_n257_));
  NOR4X1   g00193(.A(new_n257_), .B(new_n256_), .C(new_n255_), .D(new_n254_), .Y(new_n258_));
  NOR2X1   g00194(.A(new_n106_), .B(new_n72_), .Y(new_n259_));
  NOR2X1   g00195(.A(new_n129_), .B(new_n119_), .Y(new_n260_));
  NOR2X1   g00196(.A(new_n108_), .B(new_n69_), .Y(new_n261_));
  OAI22X1  g00197(.A0(new_n143_), .A1(new_n96_), .B0(new_n102_), .B1(new_n99_), .Y(new_n262_));
  NOR2X1   g00198(.A(new_n96_), .B(new_n94_), .Y(new_n263_));
  NOR2X1   g00199(.A(new_n143_), .B(new_n69_), .Y(new_n264_));
  NOR2X1   g00200(.A(new_n148_), .B(new_n127_), .Y(new_n265_));
  OR4X1    g00201(.A(new_n265_), .B(new_n264_), .C(new_n263_), .D(new_n262_), .Y(new_n266_));
  NOR4X1   g00202(.A(new_n266_), .B(new_n261_), .C(new_n260_), .D(new_n259_), .Y(new_n267_));
  NAND4X1  g00203(.A(new_n267_), .B(new_n258_), .C(new_n253_), .D(new_n248_), .Y(new_n268_));
  NOR4X1   g00204(.A(new_n268_), .B(new_n242_), .C(new_n212_), .D(new_n167_), .Y(new_n269_));
  INVX1    g00205(.A(new_n269_), .Y(new_n270_));
  OAI22X1  g00206(.A0(new_n108_), .A1(new_n75_), .B0(new_n99_), .B1(new_n91_), .Y(new_n271_));
  AOI21X1  g00207(.A0(new_n108_), .A1(new_n105_), .B0(new_n115_), .Y(new_n272_));
  NOR2X1   g00208(.A(new_n152_), .B(new_n125_), .Y(new_n273_));
  NOR2X1   g00209(.A(new_n119_), .B(new_n108_), .Y(new_n274_));
  OR4X1    g00210(.A(new_n274_), .B(new_n273_), .C(new_n272_), .D(new_n271_), .Y(new_n275_));
  NOR2X1   g00211(.A(new_n127_), .B(new_n79_), .Y(new_n276_));
  OAI22X1  g00212(.A0(new_n168_), .A1(new_n131_), .B0(new_n148_), .B1(new_n78_), .Y(new_n277_));
  OR2X1    g00213(.A(new_n277_), .B(new_n276_), .Y(new_n278_));
  INVX1    g00214(.A(new_n173_), .Y(new_n279_));
  NOR2X1   g00215(.A(new_n148_), .B(new_n108_), .Y(new_n280_));
  INVX1    g00216(.A(new_n280_), .Y(new_n281_));
  NOR2X1   g00217(.A(new_n152_), .B(new_n72_), .Y(new_n282_));
  INVX1    g00218(.A(new_n282_), .Y(new_n283_));
  NAND3X1  g00219(.A(new_n283_), .B(new_n281_), .C(new_n279_), .Y(new_n284_));
  NOR2X1   g00220(.A(new_n123_), .B(new_n108_), .Y(new_n285_));
  NOR2X1   g00221(.A(new_n182_), .B(new_n79_), .Y(new_n286_));
  OR4X1    g00222(.A(new_n286_), .B(new_n285_), .C(new_n193_), .D(new_n142_), .Y(new_n287_));
  OR4X1    g00223(.A(new_n287_), .B(new_n284_), .C(new_n278_), .D(new_n275_), .Y(new_n288_));
  OAI22X1  g00224(.A0(new_n108_), .A1(new_n69_), .B0(new_n92_), .B1(new_n75_), .Y(new_n289_));
  NOR3X1   g00225(.A(new_n289_), .B(new_n263_), .C(new_n183_), .Y(new_n290_));
  NOR2X1   g00226(.A(new_n125_), .B(new_n84_), .Y(new_n291_));
  NOR2X1   g00227(.A(new_n143_), .B(new_n96_), .Y(new_n292_));
  NOR2X1   g00228(.A(new_n94_), .B(new_n84_), .Y(new_n293_));
  NOR2X1   g00229(.A(new_n143_), .B(new_n84_), .Y(new_n294_));
  NOR4X1   g00230(.A(new_n294_), .B(new_n293_), .C(new_n292_), .D(new_n291_), .Y(new_n295_));
  NOR2X1   g00231(.A(new_n161_), .B(new_n123_), .Y(new_n296_));
  OAI22X1  g00232(.A0(new_n161_), .A1(new_n106_), .B0(new_n96_), .B1(new_n72_), .Y(new_n297_));
  OR2X1    g00233(.A(new_n297_), .B(new_n296_), .Y(new_n298_));
  NOR2X1   g00234(.A(new_n143_), .B(new_n117_), .Y(new_n299_));
  NOR2X1   g00235(.A(new_n94_), .B(new_n88_), .Y(new_n300_));
  NOR2X1   g00236(.A(new_n131_), .B(new_n123_), .Y(new_n301_));
  NOR4X1   g00237(.A(new_n301_), .B(new_n300_), .C(new_n299_), .D(new_n298_), .Y(new_n302_));
  NOR2X1   g00238(.A(new_n152_), .B(new_n143_), .Y(new_n303_));
  NOR2X1   g00239(.A(new_n105_), .B(new_n69_), .Y(new_n304_));
  AOI21X1  g00240(.A0(new_n119_), .A1(new_n91_), .B0(new_n127_), .Y(new_n305_));
  OR4X1    g00241(.A(new_n305_), .B(new_n304_), .C(new_n256_), .D(new_n303_), .Y(new_n306_));
  NOR2X1   g00242(.A(new_n105_), .B(new_n88_), .Y(new_n307_));
  OAI22X1  g00243(.A0(new_n168_), .A1(new_n161_), .B0(new_n125_), .B1(new_n123_), .Y(new_n308_));
  OAI22X1  g00244(.A0(new_n152_), .A1(new_n99_), .B0(new_n131_), .B1(new_n106_), .Y(new_n309_));
  OR4X1    g00245(.A(new_n309_), .B(new_n308_), .C(new_n219_), .D(new_n307_), .Y(new_n310_));
  OAI22X1  g00246(.A0(new_n152_), .A1(new_n92_), .B0(new_n125_), .B1(new_n119_), .Y(new_n311_));
  OAI22X1  g00247(.A0(new_n148_), .A1(new_n81_), .B0(new_n143_), .B1(new_n88_), .Y(new_n312_));
  OAI22X1  g00248(.A0(new_n182_), .A1(new_n102_), .B0(new_n115_), .B1(new_n92_), .Y(new_n313_));
  OAI22X1  g00249(.A0(new_n152_), .A1(new_n105_), .B0(new_n127_), .B1(new_n115_), .Y(new_n314_));
  OR4X1    g00250(.A(new_n314_), .B(new_n313_), .C(new_n312_), .D(new_n311_), .Y(new_n315_));
  NOR3X1   g00251(.A(new_n315_), .B(new_n310_), .C(new_n306_), .Y(new_n316_));
  NAND4X1  g00252(.A(new_n316_), .B(new_n302_), .C(new_n295_), .D(new_n290_), .Y(new_n317_));
  OR2X1    g00253(.A(new_n317_), .B(new_n288_), .Y(new_n318_));
  NOR2X1   g00254(.A(new_n94_), .B(new_n69_), .Y(new_n319_));
  INVX1    g00255(.A(new_n319_), .Y(new_n320_));
  NOR2X1   g00256(.A(new_n123_), .B(new_n72_), .Y(new_n321_));
  INVX1    g00257(.A(new_n321_), .Y(new_n322_));
  NOR2X1   g00258(.A(new_n117_), .B(new_n72_), .Y(new_n323_));
  INVX1    g00259(.A(new_n323_), .Y(new_n324_));
  NAND3X1  g00260(.A(new_n324_), .B(new_n322_), .C(new_n320_), .Y(new_n325_));
  OR2X1    g00261(.A(new_n168_), .B(new_n90_), .Y(new_n326_));
  INVX1    g00262(.A(new_n326_), .Y(new_n327_));
  NOR2X1   g00263(.A(new_n99_), .B(new_n96_), .Y(new_n328_));
  NOR2X1   g00264(.A(new_n127_), .B(new_n75_), .Y(new_n329_));
  OR4X1    g00265(.A(new_n329_), .B(new_n328_), .C(new_n208_), .D(new_n327_), .Y(new_n330_));
  NOR4X1   g00266(.A(new_n330_), .B(new_n325_), .C(new_n231_), .D(new_n86_), .Y(new_n331_));
  OAI22X1  g00267(.A0(new_n127_), .A1(new_n69_), .B0(new_n125_), .B1(new_n91_), .Y(new_n332_));
  OAI22X1  g00268(.A0(new_n125_), .A1(new_n106_), .B0(new_n78_), .B1(new_n75_), .Y(new_n333_));
  OAI22X1  g00269(.A0(new_n131_), .A1(new_n79_), .B0(new_n125_), .B1(new_n115_), .Y(new_n334_));
  OAI22X1  g00270(.A0(new_n143_), .A1(new_n79_), .B0(new_n92_), .B1(new_n84_), .Y(new_n335_));
  NOR4X1   g00271(.A(new_n335_), .B(new_n334_), .C(new_n333_), .D(new_n332_), .Y(new_n336_));
  NOR2X1   g00272(.A(new_n90_), .B(new_n88_), .Y(new_n337_));
  NOR2X1   g00273(.A(new_n106_), .B(new_n99_), .Y(new_n338_));
  OR4X1    g00274(.A(new_n247_), .B(new_n338_), .C(new_n114_), .D(new_n337_), .Y(new_n339_));
  OAI22X1  g00275(.A0(new_n127_), .A1(new_n88_), .B0(new_n125_), .B1(new_n102_), .Y(new_n340_));
  OR4X1    g00276(.A(new_n168_), .B(new_n198_), .C(new_n89_), .D(\a[23] ), .Y(new_n341_));
  OAI21X1  g00277(.A0(new_n105_), .A1(new_n84_), .B0(new_n341_), .Y(new_n342_));
  OR2X1    g00278(.A(new_n342_), .B(new_n340_), .Y(new_n343_));
  OR2X1    g00279(.A(new_n119_), .B(new_n72_), .Y(new_n344_));
  OR2X1    g00280(.A(new_n143_), .B(new_n91_), .Y(new_n345_));
  OR2X1    g00281(.A(new_n168_), .B(new_n78_), .Y(new_n346_));
  NAND3X1  g00282(.A(new_n346_), .B(new_n345_), .C(new_n344_), .Y(new_n347_));
  NOR2X1   g00283(.A(new_n108_), .B(new_n96_), .Y(new_n348_));
  OR2X1    g00284(.A(new_n127_), .B(new_n123_), .Y(new_n349_));
  INVX1    g00285(.A(new_n349_), .Y(new_n350_));
  OR4X1    g00286(.A(new_n350_), .B(new_n348_), .C(new_n240_), .D(new_n137_), .Y(new_n351_));
  NOR4X1   g00287(.A(new_n351_), .B(new_n347_), .C(new_n343_), .D(new_n339_), .Y(new_n352_));
  NAND3X1  g00288(.A(new_n352_), .B(new_n336_), .C(new_n331_), .Y(new_n353_));
  NOR2X1   g00289(.A(new_n115_), .B(new_n81_), .Y(new_n354_));
  NOR2X1   g00290(.A(new_n161_), .B(new_n96_), .Y(new_n355_));
  NOR2X1   g00291(.A(new_n99_), .B(new_n84_), .Y(new_n356_));
  NOR2X1   g00292(.A(new_n129_), .B(new_n69_), .Y(new_n357_));
  NOR2X1   g00293(.A(new_n81_), .B(new_n79_), .Y(new_n358_));
  OR4X1    g00294(.A(new_n358_), .B(new_n357_), .C(new_n200_), .D(new_n184_), .Y(new_n359_));
  OR4X1    g00295(.A(new_n359_), .B(new_n356_), .C(new_n355_), .D(new_n354_), .Y(new_n360_));
  NOR4X1   g00296(.A(new_n99_), .B(new_n98_), .C(new_n68_), .D(\a[29] ), .Y(new_n361_));
  OAI22X1  g00297(.A0(new_n119_), .A1(new_n81_), .B0(new_n117_), .B1(new_n105_), .Y(new_n362_));
  OR2X1    g00298(.A(new_n362_), .B(new_n361_), .Y(new_n363_));
  OR4X1    g00299(.A(new_n198_), .B(new_n102_), .C(new_n89_), .D(\a[23] ), .Y(new_n364_));
  INVX1    g00300(.A(new_n364_), .Y(new_n365_));
  OR4X1    g00301(.A(new_n102_), .B(new_n101_), .C(\a[26] ), .D(new_n70_), .Y(new_n366_));
  OAI21X1  g00302(.A0(new_n72_), .A1(new_n69_), .B0(new_n366_), .Y(new_n367_));
  OR2X1    g00303(.A(new_n367_), .B(new_n365_), .Y(new_n368_));
  OAI22X1  g00304(.A0(new_n143_), .A1(new_n69_), .B0(new_n106_), .B1(new_n81_), .Y(new_n369_));
  NOR2X1   g00305(.A(new_n117_), .B(new_n94_), .Y(new_n370_));
  NOR2X1   g00306(.A(new_n129_), .B(new_n91_), .Y(new_n371_));
  NOR4X1   g00307(.A(new_n168_), .B(new_n107_), .C(new_n77_), .D(\a[24] ), .Y(new_n372_));
  OR4X1    g00308(.A(new_n372_), .B(new_n371_), .C(new_n370_), .D(new_n369_), .Y(new_n373_));
  AOI21X1  g00309(.A0(new_n182_), .A1(new_n131_), .B0(new_n152_), .Y(new_n374_));
  OAI22X1  g00310(.A0(new_n168_), .A1(new_n81_), .B0(new_n90_), .B1(new_n75_), .Y(new_n375_));
  AOI21X1  g00311(.A0(new_n125_), .A1(new_n81_), .B0(new_n75_), .Y(new_n376_));
  OR4X1    g00312(.A(new_n376_), .B(new_n375_), .C(new_n374_), .D(new_n373_), .Y(new_n377_));
  OR4X1    g00313(.A(new_n377_), .B(new_n368_), .C(new_n363_), .D(new_n360_), .Y(new_n378_));
  NOR2X1   g00314(.A(new_n117_), .B(new_n81_), .Y(new_n379_));
  OR2X1    g00315(.A(new_n123_), .B(new_n105_), .Y(new_n380_));
  INVX1    g00316(.A(new_n380_), .Y(new_n381_));
  NOR2X1   g00317(.A(new_n125_), .B(new_n88_), .Y(new_n382_));
  NOR2X1   g00318(.A(new_n127_), .B(new_n106_), .Y(new_n383_));
  OR4X1    g00319(.A(new_n383_), .B(new_n382_), .C(new_n381_), .D(new_n379_), .Y(new_n384_));
  NOR2X1   g00320(.A(new_n161_), .B(new_n88_), .Y(new_n385_));
  NOR2X1   g00321(.A(new_n102_), .B(new_n78_), .Y(new_n386_));
  NOR2X1   g00322(.A(new_n168_), .B(new_n125_), .Y(new_n387_));
  OR4X1    g00323(.A(new_n387_), .B(new_n386_), .C(new_n385_), .D(new_n223_), .Y(new_n388_));
  OR4X1    g00324(.A(new_n388_), .B(new_n384_), .C(new_n194_), .D(new_n160_), .Y(new_n389_));
  NOR2X1   g00325(.A(new_n127_), .B(new_n117_), .Y(new_n390_));
  NOR2X1   g00326(.A(new_n91_), .B(new_n81_), .Y(new_n391_));
  NOR3X1   g00327(.A(new_n391_), .B(new_n233_), .C(new_n390_), .Y(new_n392_));
  NOR2X1   g00328(.A(new_n91_), .B(new_n72_), .Y(new_n393_));
  NOR2X1   g00329(.A(new_n182_), .B(new_n84_), .Y(new_n394_));
  NOR2X1   g00330(.A(new_n119_), .B(new_n90_), .Y(new_n395_));
  NOR2X1   g00331(.A(new_n161_), .B(new_n148_), .Y(new_n396_));
  NOR4X1   g00332(.A(new_n396_), .B(new_n395_), .C(new_n394_), .D(new_n393_), .Y(new_n397_));
  NOR2X1   g00333(.A(new_n148_), .B(new_n143_), .Y(new_n398_));
  NOR2X1   g00334(.A(new_n106_), .B(new_n94_), .Y(new_n399_));
  NOR2X1   g00335(.A(new_n102_), .B(new_n99_), .Y(new_n400_));
  NOR4X1   g00336(.A(new_n400_), .B(new_n399_), .C(new_n398_), .D(new_n138_), .Y(new_n401_));
  NAND3X1  g00337(.A(new_n401_), .B(new_n397_), .C(new_n392_), .Y(new_n402_));
  OR2X1    g00338(.A(new_n402_), .B(new_n389_), .Y(new_n403_));
  NOR4X1   g00339(.A(new_n403_), .B(new_n378_), .C(new_n353_), .D(new_n318_), .Y(new_n404_));
  NOR2X1   g00340(.A(new_n404_), .B(new_n270_), .Y(new_n405_));
  XOR2X1   g00341(.A(\a[30] ), .B(\a[29] ), .Y(new_n406_));
  AND2X1   g00342(.A(new_n406_), .B(\a[31] ), .Y(new_n407_));
  NOR2X1   g00343(.A(new_n92_), .B(new_n88_), .Y(new_n408_));
  NOR2X1   g00344(.A(new_n408_), .B(new_n260_), .Y(new_n409_));
  NOR2X1   g00345(.A(new_n96_), .B(new_n78_), .Y(new_n410_));
  NOR4X1   g00346(.A(new_n200_), .B(new_n410_), .C(new_n147_), .D(new_n144_), .Y(new_n411_));
  NOR2X1   g00347(.A(new_n182_), .B(new_n115_), .Y(new_n412_));
  NOR3X1   g00348(.A(new_n412_), .B(new_n356_), .C(new_n390_), .Y(new_n413_));
  NOR2X1   g00349(.A(new_n90_), .B(new_n84_), .Y(new_n414_));
  NOR3X1   g00350(.A(new_n414_), .B(new_n382_), .C(new_n294_), .Y(new_n415_));
  NAND4X1  g00351(.A(new_n415_), .B(new_n413_), .C(new_n411_), .D(new_n409_), .Y(new_n416_));
  AOI21X1  g00352(.A0(new_n182_), .A1(new_n131_), .B0(new_n75_), .Y(new_n417_));
  NOR2X1   g00353(.A(new_n131_), .B(new_n117_), .Y(new_n418_));
  OR2X1    g00354(.A(new_n418_), .B(new_n417_), .Y(new_n419_));
  NOR2X1   g00355(.A(new_n119_), .B(new_n81_), .Y(new_n420_));
  NOR2X1   g00356(.A(new_n152_), .B(new_n131_), .Y(new_n421_));
  NOR2X1   g00357(.A(new_n161_), .B(new_n69_), .Y(new_n422_));
  NOR2X1   g00358(.A(new_n115_), .B(new_n92_), .Y(new_n423_));
  OR4X1    g00359(.A(new_n395_), .B(new_n423_), .C(new_n293_), .D(new_n180_), .Y(new_n424_));
  OR4X1    g00360(.A(new_n424_), .B(new_n422_), .C(new_n421_), .D(new_n420_), .Y(new_n425_));
  NOR2X1   g00361(.A(new_n127_), .B(new_n119_), .Y(new_n426_));
  OAI22X1  g00362(.A0(new_n161_), .A1(new_n123_), .B0(new_n125_), .B1(new_n102_), .Y(new_n427_));
  OAI22X1  g00363(.A0(new_n106_), .A1(new_n81_), .B0(new_n91_), .B1(new_n90_), .Y(new_n428_));
  NOR2X1   g00364(.A(new_n148_), .B(new_n72_), .Y(new_n429_));
  OR4X1    g00365(.A(new_n429_), .B(new_n428_), .C(new_n427_), .D(new_n426_), .Y(new_n430_));
  NOR4X1   g00366(.A(new_n107_), .B(new_n102_), .C(\a[25] ), .D(new_n71_), .Y(new_n431_));
  OAI22X1  g00367(.A0(new_n131_), .A1(new_n106_), .B0(new_n115_), .B1(new_n90_), .Y(new_n432_));
  OAI22X1  g00368(.A0(new_n92_), .A1(new_n79_), .B0(new_n88_), .B1(new_n78_), .Y(new_n433_));
  OAI22X1  g00369(.A0(new_n168_), .A1(new_n92_), .B0(new_n84_), .B1(new_n78_), .Y(new_n434_));
  OR2X1    g00370(.A(new_n434_), .B(new_n433_), .Y(new_n435_));
  OR4X1    g00371(.A(new_n435_), .B(new_n432_), .C(new_n431_), .D(new_n85_), .Y(new_n436_));
  OR4X1    g00372(.A(new_n436_), .B(new_n430_), .C(new_n425_), .D(new_n419_), .Y(new_n437_));
  OR2X1    g00373(.A(new_n437_), .B(new_n416_), .Y(new_n438_));
  NOR2X1   g00374(.A(new_n182_), .B(new_n69_), .Y(new_n439_));
  AOI21X1  g00375(.A0(new_n168_), .A1(new_n79_), .B0(new_n108_), .Y(new_n440_));
  AOI21X1  g00376(.A0(new_n108_), .A1(new_n90_), .B0(new_n69_), .Y(new_n441_));
  OR4X1    g00377(.A(new_n441_), .B(new_n440_), .C(new_n439_), .D(new_n379_), .Y(new_n442_));
  INVX1    g00378(.A(new_n442_), .Y(new_n443_));
  AOI21X1  g00379(.A0(new_n131_), .A1(new_n90_), .B0(new_n79_), .Y(new_n444_));
  OAI22X1  g00380(.A0(new_n148_), .A1(new_n81_), .B0(new_n115_), .B1(new_n99_), .Y(new_n445_));
  AOI21X1  g00381(.A0(new_n129_), .A1(new_n72_), .B0(new_n88_), .Y(new_n446_));
  OAI22X1  g00382(.A0(new_n148_), .A1(new_n131_), .B0(new_n72_), .B1(new_n69_), .Y(new_n447_));
  NOR4X1   g00383(.A(new_n447_), .B(new_n446_), .C(new_n445_), .D(new_n444_), .Y(new_n448_));
  NOR2X1   g00384(.A(new_n115_), .B(new_n78_), .Y(new_n449_));
  OAI21X1  g00385(.A0(new_n94_), .A1(new_n88_), .B0(new_n214_), .Y(new_n450_));
  OAI22X1  g00386(.A0(new_n148_), .A1(new_n125_), .B0(new_n91_), .B1(new_n78_), .Y(new_n451_));
  NOR4X1   g00387(.A(new_n451_), .B(new_n450_), .C(new_n276_), .D(new_n449_), .Y(new_n452_));
  NAND3X1  g00388(.A(new_n452_), .B(new_n448_), .C(new_n443_), .Y(new_n453_));
  OAI22X1  g00389(.A0(new_n182_), .A1(new_n117_), .B0(new_n119_), .B1(new_n78_), .Y(new_n454_));
  NOR2X1   g00390(.A(new_n125_), .B(new_n123_), .Y(new_n455_));
  OR4X1    g00391(.A(new_n348_), .B(new_n455_), .C(new_n220_), .D(new_n181_), .Y(new_n456_));
  NOR2X1   g00392(.A(new_n161_), .B(new_n117_), .Y(new_n457_));
  OR4X1    g00393(.A(new_n252_), .B(new_n457_), .C(new_n213_), .D(new_n134_), .Y(new_n458_));
  NOR2X1   g00394(.A(new_n161_), .B(new_n79_), .Y(new_n459_));
  NOR2X1   g00395(.A(new_n119_), .B(new_n99_), .Y(new_n460_));
  OR4X1    g00396(.A(new_n460_), .B(new_n459_), .C(new_n387_), .D(new_n319_), .Y(new_n461_));
  OR4X1    g00397(.A(new_n461_), .B(new_n458_), .C(new_n456_), .D(new_n454_), .Y(new_n462_));
  OAI22X1  g00398(.A0(new_n105_), .A1(new_n102_), .B0(new_n79_), .B1(new_n78_), .Y(new_n463_));
  OAI22X1  g00399(.A0(new_n168_), .A1(new_n161_), .B0(new_n152_), .B1(new_n127_), .Y(new_n464_));
  OAI22X1  g00400(.A0(new_n148_), .A1(new_n105_), .B0(new_n119_), .B1(new_n72_), .Y(new_n465_));
  OR4X1    g00401(.A(new_n465_), .B(new_n464_), .C(new_n463_), .D(new_n262_), .Y(new_n466_));
  INVX1    g00402(.A(new_n223_), .Y(new_n467_));
  NOR2X1   g00403(.A(new_n102_), .B(new_n72_), .Y(new_n468_));
  INVX1    g00404(.A(new_n468_), .Y(new_n469_));
  NAND3X1  g00405(.A(new_n469_), .B(new_n283_), .C(new_n467_), .Y(new_n470_));
  OAI22X1  g00406(.A0(new_n168_), .A1(new_n99_), .B0(new_n94_), .B1(new_n91_), .Y(new_n471_));
  OR2X1    g00407(.A(new_n471_), .B(new_n172_), .Y(new_n472_));
  OR4X1    g00408(.A(new_n472_), .B(new_n470_), .C(new_n466_), .D(new_n462_), .Y(new_n473_));
  NOR2X1   g00409(.A(new_n127_), .B(new_n91_), .Y(new_n474_));
  NOR2X1   g00410(.A(new_n131_), .B(new_n69_), .Y(new_n475_));
  NOR3X1   g00411(.A(new_n475_), .B(new_n370_), .C(new_n474_), .Y(new_n476_));
  INVX1    g00412(.A(new_n476_), .Y(new_n477_));
  INVX1    g00413(.A(new_n345_), .Y(new_n478_));
  NOR2X1   g00414(.A(new_n168_), .B(new_n81_), .Y(new_n479_));
  NOR2X1   g00415(.A(new_n152_), .B(new_n78_), .Y(new_n480_));
  OR4X1    g00416(.A(new_n480_), .B(new_n399_), .C(new_n479_), .D(new_n114_), .Y(new_n481_));
  OR4X1    g00417(.A(new_n481_), .B(new_n478_), .C(new_n264_), .D(new_n126_), .Y(new_n482_));
  NOR2X1   g00418(.A(new_n127_), .B(new_n69_), .Y(new_n483_));
  OAI22X1  g00419(.A0(new_n152_), .A1(new_n125_), .B0(new_n129_), .B1(new_n91_), .Y(new_n484_));
  OAI22X1  g00420(.A0(new_n129_), .A1(new_n79_), .B0(new_n127_), .B1(new_n75_), .Y(new_n485_));
  OR4X1    g00421(.A(new_n485_), .B(new_n484_), .C(new_n483_), .D(new_n219_), .Y(new_n486_));
  OAI22X1  g00422(.A0(new_n148_), .A1(new_n143_), .B0(new_n92_), .B1(new_n75_), .Y(new_n487_));
  OAI22X1  g00423(.A0(new_n143_), .A1(new_n115_), .B0(new_n92_), .B1(new_n84_), .Y(new_n488_));
  AOI21X1  g00424(.A0(new_n106_), .A1(new_n84_), .B0(new_n182_), .Y(new_n489_));
  OAI22X1  g00425(.A0(new_n131_), .A1(new_n123_), .B0(new_n102_), .B1(new_n90_), .Y(new_n490_));
  OR4X1    g00426(.A(new_n490_), .B(new_n489_), .C(new_n488_), .D(new_n487_), .Y(new_n491_));
  OR4X1    g00427(.A(new_n491_), .B(new_n486_), .C(new_n482_), .D(new_n477_), .Y(new_n492_));
  NOR2X1   g00428(.A(new_n129_), .B(new_n75_), .Y(new_n493_));
  NOR2X1   g00429(.A(new_n129_), .B(new_n84_), .Y(new_n494_));
  OR4X1    g00430(.A(new_n494_), .B(new_n493_), .C(new_n228_), .D(new_n175_), .Y(new_n495_));
  NOR2X1   g00431(.A(new_n105_), .B(new_n96_), .Y(new_n496_));
  NOR4X1   g00432(.A(new_n125_), .B(new_n98_), .C(new_n68_), .D(\a[29] ), .Y(new_n497_));
  OAI22X1  g00433(.A0(new_n161_), .A1(new_n119_), .B0(new_n105_), .B1(new_n69_), .Y(new_n498_));
  OR4X1    g00434(.A(new_n498_), .B(new_n497_), .C(new_n496_), .D(new_n495_), .Y(new_n499_));
  NOR2X1   g00435(.A(new_n152_), .B(new_n108_), .Y(new_n500_));
  OAI22X1  g00436(.A0(new_n108_), .A1(new_n88_), .B0(new_n99_), .B1(new_n96_), .Y(new_n501_));
  OR2X1    g00437(.A(new_n501_), .B(new_n500_), .Y(new_n502_));
  OR2X1    g00438(.A(new_n115_), .B(new_n72_), .Y(new_n503_));
  INVX1    g00439(.A(new_n503_), .Y(new_n504_));
  NOR4X1   g00440(.A(new_n99_), .B(new_n98_), .C(\a[30] ), .D(new_n74_), .Y(new_n505_));
  NOR2X1   g00441(.A(new_n131_), .B(new_n88_), .Y(new_n506_));
  OR4X1    g00442(.A(new_n506_), .B(new_n505_), .C(new_n504_), .D(new_n502_), .Y(new_n507_));
  OAI22X1  g00443(.A0(new_n182_), .A1(new_n148_), .B0(new_n168_), .B1(new_n90_), .Y(new_n508_));
  NOR2X1   g00444(.A(new_n96_), .B(new_n90_), .Y(new_n509_));
  NOR2X1   g00445(.A(new_n123_), .B(new_n78_), .Y(new_n510_));
  OAI22X1  g00446(.A0(new_n182_), .A1(new_n102_), .B0(new_n129_), .B1(new_n115_), .Y(new_n511_));
  OR4X1    g00447(.A(new_n511_), .B(new_n510_), .C(new_n509_), .D(new_n508_), .Y(new_n512_));
  OAI21X1  g00448(.A0(new_n92_), .A1(new_n69_), .B0(new_n366_), .Y(new_n513_));
  OAI22X1  g00449(.A0(new_n168_), .A1(new_n78_), .B0(new_n129_), .B1(new_n123_), .Y(new_n514_));
  OAI22X1  g00450(.A0(new_n152_), .A1(new_n105_), .B0(new_n78_), .B1(new_n69_), .Y(new_n515_));
  OAI22X1  g00451(.A0(new_n152_), .A1(new_n129_), .B0(new_n125_), .B1(new_n79_), .Y(new_n516_));
  OR4X1    g00452(.A(new_n516_), .B(new_n515_), .C(new_n514_), .D(new_n513_), .Y(new_n517_));
  OR4X1    g00453(.A(new_n517_), .B(new_n512_), .C(new_n507_), .D(new_n499_), .Y(new_n518_));
  OR4X1    g00454(.A(new_n518_), .B(new_n492_), .C(new_n473_), .D(new_n453_), .Y(new_n519_));
  NOR2X1   g00455(.A(new_n519_), .B(new_n438_), .Y(new_n520_));
  NOR2X1   g00456(.A(new_n92_), .B(new_n91_), .Y(new_n521_));
  NOR2X1   g00457(.A(new_n182_), .B(new_n91_), .Y(new_n522_));
  NOR2X1   g00458(.A(new_n131_), .B(new_n75_), .Y(new_n523_));
  OAI22X1  g00459(.A0(new_n123_), .A1(new_n92_), .B0(new_n84_), .B1(new_n81_), .Y(new_n524_));
  OR4X1    g00460(.A(new_n524_), .B(new_n523_), .C(new_n522_), .D(new_n521_), .Y(new_n525_));
  OR2X1    g00461(.A(new_n148_), .B(new_n92_), .Y(new_n526_));
  INVX1    g00462(.A(new_n526_), .Y(new_n527_));
  OAI22X1  g00463(.A0(new_n161_), .A1(new_n119_), .B0(new_n148_), .B1(new_n72_), .Y(new_n528_));
  OR4X1    g00464(.A(new_n285_), .B(new_n282_), .C(new_n256_), .D(new_n162_), .Y(new_n529_));
  OAI22X1  g00465(.A0(new_n182_), .A1(new_n96_), .B0(new_n108_), .B1(new_n115_), .Y(new_n530_));
  OAI22X1  g00466(.A0(new_n143_), .A1(new_n96_), .B0(new_n123_), .B1(new_n99_), .Y(new_n531_));
  OR2X1    g00467(.A(new_n531_), .B(new_n530_), .Y(new_n532_));
  OR4X1    g00468(.A(new_n532_), .B(new_n529_), .C(new_n528_), .D(new_n527_), .Y(new_n533_));
  OR2X1    g00469(.A(new_n533_), .B(new_n525_), .Y(new_n534_));
  NOR2X1   g00470(.A(new_n127_), .B(new_n88_), .Y(new_n535_));
  NOR2X1   g00471(.A(new_n148_), .B(new_n78_), .Y(new_n536_));
  AOI21X1  g00472(.A0(new_n105_), .A1(new_n78_), .B0(new_n75_), .Y(new_n537_));
  NOR3X1   g00473(.A(new_n537_), .B(new_n536_), .C(new_n535_), .Y(new_n538_));
  NOR2X1   g00474(.A(new_n182_), .B(new_n152_), .Y(new_n539_));
  INVX1    g00475(.A(new_n366_), .Y(new_n540_));
  NOR2X1   g00476(.A(new_n106_), .B(new_n92_), .Y(new_n541_));
  NOR4X1   g00477(.A(new_n541_), .B(new_n540_), .C(new_n539_), .D(new_n303_), .Y(new_n542_));
  NOR4X1   g00478(.A(new_n168_), .B(new_n101_), .C(new_n89_), .D(\a[23] ), .Y(new_n543_));
  NOR3X1   g00479(.A(new_n543_), .B(new_n252_), .C(new_n219_), .Y(new_n544_));
  NAND3X1  g00480(.A(new_n544_), .B(new_n542_), .C(new_n538_), .Y(new_n545_));
  NOR2X1   g00481(.A(new_n129_), .B(new_n123_), .Y(new_n546_));
  NOR2X1   g00482(.A(new_n78_), .B(new_n69_), .Y(new_n547_));
  OR4X1    g00483(.A(new_n365_), .B(new_n233_), .C(new_n218_), .D(new_n114_), .Y(new_n548_));
  OR4X1    g00484(.A(new_n548_), .B(new_n547_), .C(new_n546_), .D(new_n207_), .Y(new_n549_));
  OAI22X1  g00485(.A0(new_n161_), .A1(new_n96_), .B0(new_n91_), .B1(new_n90_), .Y(new_n550_));
  OR4X1    g00486(.A(new_n99_), .B(new_n98_), .C(\a[30] ), .D(new_n74_), .Y(new_n551_));
  OAI21X1  g00487(.A0(new_n91_), .A1(new_n81_), .B0(new_n551_), .Y(new_n552_));
  OAI22X1  g00488(.A0(new_n117_), .A1(new_n94_), .B0(new_n105_), .B1(new_n84_), .Y(new_n553_));
  NOR4X1   g00489(.A(\a[26] ), .B(\a[25] ), .C(new_n71_), .D(\a[23] ), .Y(new_n554_));
  NOR3X1   g00490(.A(new_n98_), .B(new_n68_), .C(new_n74_), .Y(new_n555_));
  NOR2X1   g00491(.A(new_n107_), .B(new_n198_), .Y(new_n556_));
  NOR4X1   g00492(.A(new_n68_), .B(\a[29] ), .C(new_n95_), .D(\a[27] ), .Y(new_n557_));
  AOI22X1  g00493(.A0(new_n557_), .A1(new_n556_), .B0(new_n555_), .B1(new_n554_), .Y(new_n558_));
  INVX1    g00494(.A(new_n558_), .Y(new_n559_));
  OAI22X1  g00495(.A0(new_n127_), .A1(new_n106_), .B0(new_n105_), .B1(new_n115_), .Y(new_n560_));
  OAI22X1  g00496(.A0(new_n152_), .A1(new_n131_), .B0(new_n102_), .B1(new_n92_), .Y(new_n561_));
  OR4X1    g00497(.A(new_n561_), .B(new_n560_), .C(new_n559_), .D(new_n433_), .Y(new_n562_));
  OR4X1    g00498(.A(new_n562_), .B(new_n553_), .C(new_n552_), .D(new_n550_), .Y(new_n563_));
  OR4X1    g00499(.A(new_n563_), .B(new_n549_), .C(new_n545_), .D(new_n534_), .Y(new_n564_));
  NOR4X1   g00500(.A(new_n198_), .B(new_n102_), .C(\a[26] ), .D(\a[23] ), .Y(new_n565_));
  AOI21X1  g00501(.A0(new_n81_), .A1(new_n72_), .B0(new_n102_), .Y(new_n566_));
  OR4X1    g00502(.A(new_n566_), .B(new_n565_), .C(new_n193_), .D(new_n103_), .Y(new_n567_));
  OAI22X1  g00503(.A0(new_n152_), .A1(new_n125_), .B0(new_n119_), .B1(new_n108_), .Y(new_n568_));
  OAI22X1  g00504(.A0(new_n117_), .A1(new_n105_), .B0(new_n94_), .B1(new_n91_), .Y(new_n569_));
  OAI22X1  g00505(.A0(new_n182_), .A1(new_n117_), .B0(new_n115_), .B1(new_n72_), .Y(new_n570_));
  OAI22X1  g00506(.A0(new_n161_), .A1(new_n106_), .B0(new_n72_), .B1(new_n69_), .Y(new_n571_));
  OAI22X1  g00507(.A0(new_n129_), .A1(new_n75_), .B0(new_n125_), .B1(new_n96_), .Y(new_n572_));
  OR4X1    g00508(.A(new_n572_), .B(new_n571_), .C(new_n570_), .D(new_n569_), .Y(new_n573_));
  NOR2X1   g00509(.A(new_n131_), .B(new_n79_), .Y(new_n574_));
  OR4X1    g00510(.A(new_n574_), .B(new_n144_), .C(new_n126_), .D(new_n111_), .Y(new_n575_));
  OR4X1    g00511(.A(new_n575_), .B(new_n573_), .C(new_n464_), .D(new_n568_), .Y(new_n576_));
  OR2X1    g00512(.A(new_n576_), .B(new_n567_), .Y(new_n577_));
  NOR2X1   g00513(.A(new_n108_), .B(new_n88_), .Y(new_n578_));
  NOR3X1   g00514(.A(new_n168_), .B(new_n107_), .C(new_n101_), .Y(new_n579_));
  OR4X1    g00515(.A(new_n579_), .B(new_n348_), .C(new_n578_), .D(new_n410_), .Y(new_n580_));
  NOR2X1   g00516(.A(new_n152_), .B(new_n90_), .Y(new_n581_));
  OAI22X1  g00517(.A0(new_n106_), .A1(new_n105_), .B0(new_n96_), .B1(new_n81_), .Y(new_n582_));
  OR4X1    g00518(.A(new_n582_), .B(new_n494_), .C(new_n581_), .D(new_n118_), .Y(new_n583_));
  OR2X1    g00519(.A(new_n583_), .B(new_n580_), .Y(new_n584_));
  NOR2X1   g00520(.A(new_n96_), .B(new_n92_), .Y(new_n585_));
  NOR2X1   g00521(.A(new_n161_), .B(new_n75_), .Y(new_n586_));
  OR4X1    g00522(.A(new_n586_), .B(new_n213_), .C(new_n134_), .D(new_n585_), .Y(new_n587_));
  INVX1    g00523(.A(new_n500_), .Y(new_n588_));
  NOR2X1   g00524(.A(new_n152_), .B(new_n81_), .Y(new_n589_));
  INVX1    g00525(.A(new_n589_), .Y(new_n590_));
  NAND3X1  g00526(.A(new_n590_), .B(new_n588_), .C(new_n344_), .Y(new_n591_));
  OR4X1    g00527(.A(new_n591_), .B(new_n381_), .C(new_n180_), .D(new_n291_), .Y(new_n592_));
  NOR4X1   g00528(.A(new_n592_), .B(new_n587_), .C(new_n584_), .D(new_n577_), .Y(new_n593_));
  NOR2X1   g00529(.A(new_n143_), .B(new_n123_), .Y(new_n594_));
  OAI22X1  g00530(.A0(new_n125_), .A1(new_n91_), .B0(new_n96_), .B1(new_n94_), .Y(new_n595_));
  NOR2X1   g00531(.A(new_n148_), .B(new_n99_), .Y(new_n596_));
  OR4X1    g00532(.A(new_n596_), .B(new_n496_), .C(new_n480_), .D(new_n361_), .Y(new_n597_));
  NOR2X1   g00533(.A(new_n143_), .B(new_n88_), .Y(new_n598_));
  OR4X1    g00534(.A(new_n422_), .B(new_n394_), .C(new_n371_), .D(new_n598_), .Y(new_n599_));
  OR4X1    g00535(.A(new_n599_), .B(new_n597_), .C(new_n595_), .D(new_n594_), .Y(new_n600_));
  OR4X1    g00536(.A(new_n358_), .B(new_n239_), .C(new_n203_), .D(new_n124_), .Y(new_n601_));
  OAI22X1  g00537(.A0(new_n182_), .A1(new_n79_), .B0(new_n168_), .B1(new_n127_), .Y(new_n602_));
  NOR2X1   g00538(.A(new_n125_), .B(new_n102_), .Y(new_n603_));
  OR4X1    g00539(.A(new_n603_), .B(new_n296_), .C(new_n327_), .D(new_n337_), .Y(new_n604_));
  OR4X1    g00540(.A(new_n604_), .B(new_n602_), .C(new_n601_), .D(new_n600_), .Y(new_n605_));
  NOR4X1   g00541(.A(new_n234_), .B(new_n202_), .C(new_n184_), .D(new_n173_), .Y(new_n606_));
  OAI22X1  g00542(.A0(new_n129_), .A1(new_n106_), .B0(new_n125_), .B1(new_n117_), .Y(new_n607_));
  OAI22X1  g00543(.A0(new_n152_), .A1(new_n99_), .B0(new_n119_), .B1(new_n78_), .Y(new_n608_));
  NOR2X1   g00544(.A(new_n608_), .B(new_n607_), .Y(new_n609_));
  NOR2X1   g00545(.A(new_n152_), .B(new_n92_), .Y(new_n610_));
  NOR3X1   g00546(.A(new_n300_), .B(new_n246_), .C(new_n610_), .Y(new_n611_));
  NOR2X1   g00547(.A(new_n129_), .B(new_n115_), .Y(new_n612_));
  NOR4X1   g00548(.A(new_n612_), .B(new_n459_), .C(new_n412_), .D(new_n265_), .Y(new_n613_));
  NAND4X1  g00549(.A(new_n613_), .B(new_n611_), .C(new_n609_), .D(new_n606_), .Y(new_n614_));
  NOR2X1   g00550(.A(new_n152_), .B(new_n105_), .Y(new_n615_));
  NOR2X1   g00551(.A(new_n182_), .B(new_n123_), .Y(new_n616_));
  OAI22X1  g00552(.A0(new_n143_), .A1(new_n117_), .B0(new_n123_), .B1(new_n94_), .Y(new_n617_));
  OAI22X1  g00553(.A0(new_n182_), .A1(new_n88_), .B0(new_n123_), .B1(new_n90_), .Y(new_n618_));
  OR4X1    g00554(.A(new_n618_), .B(new_n617_), .C(new_n616_), .D(new_n183_), .Y(new_n619_));
  OR4X1    g00555(.A(new_n619_), .B(new_n615_), .C(new_n474_), .D(new_n426_), .Y(new_n620_));
  NOR3X1   g00556(.A(new_n620_), .B(new_n614_), .C(new_n605_), .Y(new_n621_));
  NAND2X1  g00557(.A(new_n621_), .B(new_n593_), .Y(new_n622_));
  NOR2X1   g00558(.A(new_n622_), .B(new_n564_), .Y(new_n623_));
  NOR2X1   g00559(.A(new_n623_), .B(new_n520_), .Y(new_n624_));
  OAI22X1  g00560(.A0(new_n105_), .A1(new_n115_), .B0(new_n92_), .B1(new_n88_), .Y(new_n625_));
  OR2X1    g00561(.A(new_n625_), .B(new_n589_), .Y(new_n626_));
  NOR2X1   g00562(.A(new_n125_), .B(new_n91_), .Y(new_n627_));
  OR4X1    g00563(.A(new_n627_), .B(new_n232_), .C(new_n220_), .D(new_n303_), .Y(new_n628_));
  OAI22X1  g00564(.A0(new_n148_), .A1(new_n81_), .B0(new_n90_), .B1(new_n79_), .Y(new_n629_));
  OR4X1    g00565(.A(new_n629_), .B(new_n628_), .C(new_n626_), .D(new_n552_), .Y(new_n630_));
  NOR2X1   g00566(.A(new_n123_), .B(new_n92_), .Y(new_n631_));
  NOR2X1   g00567(.A(new_n96_), .B(new_n81_), .Y(new_n632_));
  OAI22X1  g00568(.A0(new_n125_), .A1(new_n106_), .B0(new_n105_), .B1(new_n69_), .Y(new_n633_));
  NOR2X1   g00569(.A(new_n105_), .B(new_n79_), .Y(new_n634_));
  OR4X1    g00570(.A(new_n634_), .B(new_n633_), .C(new_n632_), .D(new_n631_), .Y(new_n635_));
  NOR2X1   g00571(.A(new_n117_), .B(new_n78_), .Y(new_n636_));
  OR4X1    g00572(.A(new_n636_), .B(new_n527_), .C(new_n393_), .D(new_n439_), .Y(new_n637_));
  OAI21X1  g00573(.A0(new_n75_), .A1(new_n72_), .B0(new_n364_), .Y(new_n638_));
  OR4X1    g00574(.A(new_n638_), .B(new_n637_), .C(new_n256_), .D(new_n218_), .Y(new_n639_));
  AOI21X1  g00575(.A0(new_n123_), .A1(new_n84_), .B0(new_n81_), .Y(new_n640_));
  AOI21X1  g00576(.A0(new_n129_), .A1(new_n108_), .B0(new_n102_), .Y(new_n641_));
  NOR2X1   g00577(.A(new_n127_), .B(new_n96_), .Y(new_n642_));
  OR4X1    g00578(.A(new_n642_), .B(new_n641_), .C(new_n640_), .D(new_n160_), .Y(new_n643_));
  NOR4X1   g00579(.A(new_n643_), .B(new_n639_), .C(new_n635_), .D(new_n630_), .Y(new_n644_));
  INVX1    g00580(.A(new_n644_), .Y(new_n645_));
  OAI22X1  g00581(.A0(new_n152_), .A1(new_n125_), .B0(new_n143_), .B1(new_n84_), .Y(new_n646_));
  AOI21X1  g00582(.A0(new_n161_), .A1(new_n72_), .B0(new_n69_), .Y(new_n647_));
  NOR2X1   g00583(.A(new_n125_), .B(new_n75_), .Y(new_n648_));
  OR4X1    g00584(.A(new_n172_), .B(new_n648_), .C(new_n139_), .D(new_n585_), .Y(new_n649_));
  OR4X1    g00585(.A(new_n649_), .B(new_n647_), .C(new_n646_), .D(new_n395_), .Y(new_n650_));
  NOR2X1   g00586(.A(new_n119_), .B(new_n94_), .Y(new_n651_));
  OAI22X1  g00587(.A0(new_n127_), .A1(new_n117_), .B0(new_n125_), .B1(new_n96_), .Y(new_n652_));
  OAI22X1  g00588(.A0(new_n182_), .A1(new_n106_), .B0(new_n168_), .B1(new_n161_), .Y(new_n653_));
  OR4X1    g00589(.A(new_n653_), .B(new_n652_), .C(new_n616_), .D(new_n651_), .Y(new_n654_));
  OAI22X1  g00590(.A0(new_n161_), .A1(new_n115_), .B0(new_n117_), .B1(new_n99_), .Y(new_n655_));
  OAI22X1  g00591(.A0(new_n148_), .A1(new_n108_), .B0(new_n129_), .B1(new_n119_), .Y(new_n656_));
  OAI22X1  g00592(.A0(new_n129_), .A1(new_n69_), .B0(new_n117_), .B1(new_n90_), .Y(new_n657_));
  OR4X1    g00593(.A(new_n657_), .B(new_n656_), .C(new_n655_), .D(new_n190_), .Y(new_n658_));
  OAI22X1  g00594(.A0(new_n161_), .A1(new_n84_), .B0(new_n131_), .B1(new_n91_), .Y(new_n659_));
  OAI22X1  g00595(.A0(new_n129_), .A1(new_n106_), .B0(new_n125_), .B1(new_n115_), .Y(new_n660_));
  OR4X1    g00596(.A(new_n660_), .B(new_n659_), .C(new_n423_), .D(new_n309_), .Y(new_n661_));
  OR4X1    g00597(.A(new_n661_), .B(new_n658_), .C(new_n654_), .D(new_n650_), .Y(new_n662_));
  OR4X1    g00598(.A(new_n412_), .B(new_n276_), .C(new_n191_), .D(new_n337_), .Y(new_n663_));
  NOR2X1   g00599(.A(new_n90_), .B(new_n75_), .Y(new_n664_));
  OR4X1    g00600(.A(new_n479_), .B(new_n664_), .C(new_n156_), .D(new_n155_), .Y(new_n665_));
  OAI22X1  g00601(.A0(new_n125_), .A1(new_n117_), .B0(new_n119_), .B1(new_n81_), .Y(new_n666_));
  OAI22X1  g00602(.A0(new_n106_), .A1(new_n81_), .B0(new_n84_), .B1(new_n72_), .Y(new_n667_));
  OAI22X1  g00603(.A0(new_n161_), .A1(new_n117_), .B0(new_n94_), .B1(new_n69_), .Y(new_n668_));
  OAI22X1  g00604(.A0(new_n182_), .A1(new_n119_), .B0(new_n94_), .B1(new_n84_), .Y(new_n669_));
  OR4X1    g00605(.A(new_n669_), .B(new_n668_), .C(new_n667_), .D(new_n666_), .Y(new_n670_));
  OAI22X1  g00606(.A0(new_n125_), .A1(new_n123_), .B0(new_n108_), .B1(new_n96_), .Y(new_n671_));
  OR2X1    g00607(.A(new_n671_), .B(new_n417_), .Y(new_n672_));
  OAI22X1  g00608(.A0(new_n168_), .A1(new_n127_), .B0(new_n148_), .B1(new_n72_), .Y(new_n673_));
  OR4X1    g00609(.A(new_n673_), .B(new_n672_), .C(new_n478_), .D(new_n251_), .Y(new_n674_));
  OR4X1    g00610(.A(new_n674_), .B(new_n670_), .C(new_n665_), .D(new_n663_), .Y(new_n675_));
  AOI21X1  g00611(.A0(new_n182_), .A1(new_n161_), .B0(new_n88_), .Y(new_n676_));
  NOR4X1   g00612(.A(new_n676_), .B(new_n440_), .C(new_n493_), .D(new_n134_), .Y(new_n677_));
  NOR2X1   g00613(.A(new_n78_), .B(new_n75_), .Y(new_n678_));
  NOR2X1   g00614(.A(new_n152_), .B(new_n127_), .Y(new_n679_));
  NOR3X1   g00615(.A(new_n612_), .B(new_n679_), .C(new_n678_), .Y(new_n680_));
  NOR2X1   g00616(.A(new_n125_), .B(new_n119_), .Y(new_n681_));
  NOR4X1   g00617(.A(new_n394_), .B(new_n598_), .C(new_n681_), .D(new_n197_), .Y(new_n682_));
  NAND3X1  g00618(.A(new_n682_), .B(new_n680_), .C(new_n677_), .Y(new_n683_));
  OAI22X1  g00619(.A0(new_n127_), .A1(new_n88_), .B0(new_n102_), .B1(new_n94_), .Y(new_n684_));
  OR2X1    g00620(.A(new_n684_), .B(new_n383_), .Y(new_n685_));
  OR2X1    g00621(.A(new_n450_), .B(new_n399_), .Y(new_n686_));
  OR4X1    g00622(.A(new_n686_), .B(new_n387_), .C(new_n118_), .D(new_n307_), .Y(new_n687_));
  OR4X1    g00623(.A(new_n687_), .B(new_n685_), .C(new_n683_), .D(new_n675_), .Y(new_n688_));
  OR2X1    g00624(.A(new_n688_), .B(new_n662_), .Y(new_n689_));
  NOR2X1   g00625(.A(new_n689_), .B(new_n645_), .Y(new_n690_));
  NOR2X1   g00626(.A(new_n92_), .B(new_n75_), .Y(new_n691_));
  NOR4X1   g00627(.A(new_n427_), .B(new_n372_), .C(new_n328_), .D(new_n691_), .Y(new_n692_));
  NOR4X1   g00628(.A(new_n541_), .B(new_n447_), .C(new_n321_), .D(new_n282_), .Y(new_n693_));
  AOI21X1  g00629(.A0(new_n92_), .A1(new_n90_), .B0(new_n168_), .Y(new_n694_));
  OAI22X1  g00630(.A0(new_n105_), .A1(new_n102_), .B0(new_n90_), .B1(new_n75_), .Y(new_n695_));
  OR4X1    g00631(.A(new_n695_), .B(new_n694_), .C(new_n396_), .D(new_n285_), .Y(new_n696_));
  INVX1    g00632(.A(new_n696_), .Y(new_n697_));
  NAND3X1  g00633(.A(new_n697_), .B(new_n693_), .C(new_n692_), .Y(new_n698_));
  OR4X1    g00634(.A(new_n233_), .B(new_n158_), .C(new_n337_), .D(new_n80_), .Y(new_n699_));
  AOI21X1  g00635(.A0(new_n161_), .A1(new_n143_), .B0(new_n96_), .Y(new_n700_));
  OAI22X1  g00636(.A0(new_n117_), .A1(new_n78_), .B0(new_n102_), .B1(new_n94_), .Y(new_n701_));
  NOR2X1   g00637(.A(new_n92_), .B(new_n79_), .Y(new_n702_));
  OR4X1    g00638(.A(new_n547_), .B(new_n500_), .C(new_n273_), .D(new_n183_), .Y(new_n703_));
  OR4X1    g00639(.A(new_n703_), .B(new_n632_), .C(new_n702_), .D(new_n356_), .Y(new_n704_));
  OR4X1    g00640(.A(new_n704_), .B(new_n701_), .C(new_n700_), .D(new_n699_), .Y(new_n705_));
  OR2X1    g00641(.A(new_n148_), .B(new_n78_), .Y(new_n706_));
  INVX1    g00642(.A(new_n247_), .Y(new_n707_));
  NAND3X1  g00643(.A(new_n707_), .B(new_n706_), .C(new_n214_), .Y(new_n708_));
  OR4X1    g00644(.A(new_n546_), .B(new_n421_), .C(new_n598_), .D(new_n261_), .Y(new_n709_));
  OAI22X1  g00645(.A0(new_n182_), .A1(new_n152_), .B0(new_n115_), .B1(new_n94_), .Y(new_n710_));
  OAI22X1  g00646(.A0(new_n143_), .A1(new_n75_), .B0(new_n108_), .B1(new_n102_), .Y(new_n711_));
  OR4X1    g00647(.A(new_n711_), .B(new_n710_), .C(new_n709_), .D(new_n708_), .Y(new_n712_));
  OR4X1    g00648(.A(new_n480_), .B(new_n414_), .C(new_n114_), .D(new_n521_), .Y(new_n713_));
  OAI22X1  g00649(.A0(new_n143_), .A1(new_n84_), .B0(new_n129_), .B1(new_n79_), .Y(new_n714_));
  NOR2X1   g00650(.A(new_n293_), .B(new_n239_), .Y(new_n715_));
  INVX1    g00651(.A(new_n715_), .Y(new_n716_));
  NOR2X1   g00652(.A(new_n131_), .B(new_n106_), .Y(new_n717_));
  INVX1    g00653(.A(new_n717_), .Y(new_n718_));
  OR2X1    g00654(.A(new_n143_), .B(new_n123_), .Y(new_n719_));
  NOR2X1   g00655(.A(new_n106_), .B(new_n90_), .Y(new_n720_));
  INVX1    g00656(.A(new_n720_), .Y(new_n721_));
  NAND3X1  g00657(.A(new_n721_), .B(new_n719_), .C(new_n718_), .Y(new_n722_));
  NOR4X1   g00658(.A(new_n168_), .B(new_n101_), .C(\a[26] ), .D(new_n70_), .Y(new_n723_));
  NOR2X1   g00659(.A(new_n131_), .B(new_n84_), .Y(new_n724_));
  OR4X1    g00660(.A(new_n724_), .B(new_n723_), .C(new_n722_), .D(new_n418_), .Y(new_n725_));
  OR4X1    g00661(.A(new_n725_), .B(new_n716_), .C(new_n714_), .D(new_n713_), .Y(new_n726_));
  OR4X1    g00662(.A(new_n726_), .B(new_n712_), .C(new_n705_), .D(new_n698_), .Y(new_n727_));
  OAI22X1  g00663(.A0(new_n123_), .A1(new_n92_), .B0(new_n117_), .B1(new_n72_), .Y(new_n728_));
  OAI22X1  g00664(.A0(new_n119_), .A1(new_n90_), .B0(new_n92_), .B1(new_n69_), .Y(new_n729_));
  OR4X1    g00665(.A(new_n729_), .B(new_n728_), .C(new_n354_), .D(new_n423_), .Y(new_n730_));
  OAI22X1  g00666(.A0(new_n143_), .A1(new_n106_), .B0(new_n129_), .B1(new_n69_), .Y(new_n731_));
  OR2X1    g00667(.A(new_n731_), .B(new_n642_), .Y(new_n732_));
  OAI22X1  g00668(.A0(new_n125_), .A1(new_n75_), .B0(new_n119_), .B1(new_n94_), .Y(new_n733_));
  OR2X1    g00669(.A(new_n733_), .B(new_n634_), .Y(new_n734_));
  OR4X1    g00670(.A(new_n394_), .B(new_n627_), .C(new_n479_), .D(new_n223_), .Y(new_n735_));
  OR4X1    g00671(.A(new_n735_), .B(new_n734_), .C(new_n732_), .D(new_n730_), .Y(new_n736_));
  OAI22X1  g00672(.A0(new_n125_), .A1(new_n84_), .B0(new_n108_), .B1(new_n91_), .Y(new_n737_));
  OR2X1    g00673(.A(new_n737_), .B(new_n178_), .Y(new_n738_));
  OR4X1    g00674(.A(new_n510_), .B(new_n300_), .C(new_n616_), .D(new_n232_), .Y(new_n739_));
  NOR2X1   g00675(.A(new_n161_), .B(new_n119_), .Y(new_n740_));
  NOR2X1   g00676(.A(new_n119_), .B(new_n105_), .Y(new_n741_));
  OR4X1    g00677(.A(new_n741_), .B(new_n740_), .C(new_n361_), .D(new_n585_), .Y(new_n742_));
  AOI21X1  g00678(.A0(new_n94_), .A1(new_n90_), .B0(new_n96_), .Y(new_n743_));
  OAI22X1  g00679(.A0(new_n131_), .A1(new_n123_), .B0(new_n127_), .B1(new_n106_), .Y(new_n744_));
  OR4X1    g00680(.A(new_n744_), .B(new_n743_), .C(new_n199_), .D(new_n100_), .Y(new_n745_));
  NOR2X1   g00681(.A(new_n161_), .B(new_n106_), .Y(new_n746_));
  NOR2X1   g00682(.A(new_n105_), .B(new_n84_), .Y(new_n747_));
  OR4X1    g00683(.A(new_n370_), .B(new_n747_), .C(new_n219_), .D(new_n746_), .Y(new_n748_));
  OR2X1    g00684(.A(new_n168_), .B(new_n125_), .Y(new_n749_));
  OAI21X1  g00685(.A0(new_n119_), .A1(new_n108_), .B0(new_n749_), .Y(new_n750_));
  AOI21X1  g00686(.A0(new_n143_), .A1(new_n108_), .B0(new_n117_), .Y(new_n751_));
  OR4X1    g00687(.A(new_n751_), .B(new_n750_), .C(new_n748_), .D(new_n745_), .Y(new_n752_));
  OR4X1    g00688(.A(new_n752_), .B(new_n742_), .C(new_n739_), .D(new_n738_), .Y(new_n753_));
  OR2X1    g00689(.A(new_n753_), .B(new_n736_), .Y(new_n754_));
  NOR2X1   g00690(.A(new_n123_), .B(new_n94_), .Y(new_n755_));
  OR4X1    g00691(.A(new_n755_), .B(new_n612_), .C(new_n420_), .D(new_n286_), .Y(new_n756_));
  NOR2X1   g00692(.A(new_n94_), .B(new_n75_), .Y(new_n757_));
  NOR4X1   g00693(.A(new_n168_), .B(new_n107_), .C(\a[25] ), .D(new_n71_), .Y(new_n758_));
  OR4X1    g00694(.A(new_n758_), .B(new_n757_), .C(new_n535_), .D(new_n86_), .Y(new_n759_));
  OR4X1    g00695(.A(new_n759_), .B(new_n271_), .C(new_n251_), .D(new_n431_), .Y(new_n760_));
  OR4X1    g00696(.A(new_n629_), .B(new_n276_), .C(new_n426_), .D(new_n449_), .Y(new_n761_));
  INVX1    g00697(.A(new_n439_), .Y(new_n762_));
  NOR3X1   g00698(.A(new_n596_), .B(new_n338_), .C(new_n126_), .Y(new_n763_));
  NAND3X1  g00699(.A(new_n763_), .B(new_n281_), .C(new_n762_), .Y(new_n764_));
  OR4X1    g00700(.A(new_n764_), .B(new_n761_), .C(new_n760_), .D(new_n756_), .Y(new_n765_));
  OAI22X1  g00701(.A0(new_n161_), .A1(new_n152_), .B0(new_n108_), .B1(new_n79_), .Y(new_n766_));
  AOI21X1  g00702(.A0(new_n125_), .A1(new_n92_), .B0(new_n148_), .Y(new_n767_));
  OAI22X1  g00703(.A0(new_n125_), .A1(new_n69_), .B0(new_n119_), .B1(new_n99_), .Y(new_n768_));
  OAI21X1  g00704(.A0(new_n161_), .A1(new_n91_), .B0(new_n341_), .Y(new_n769_));
  NOR4X1   g00705(.A(new_n769_), .B(new_n768_), .C(new_n767_), .D(new_n766_), .Y(new_n770_));
  NOR3X1   g00706(.A(new_n543_), .B(new_n505_), .C(new_n579_), .Y(new_n771_));
  OAI22X1  g00707(.A0(new_n106_), .A1(new_n81_), .B0(new_n92_), .B1(new_n84_), .Y(new_n772_));
  NOR3X1   g00708(.A(new_n772_), .B(new_n615_), .C(new_n400_), .Y(new_n773_));
  NAND3X1  g00709(.A(new_n773_), .B(new_n771_), .C(new_n770_), .Y(new_n774_));
  OAI22X1  g00710(.A0(new_n182_), .A1(new_n88_), .B0(new_n143_), .B1(new_n79_), .Y(new_n775_));
  OR4X1    g00711(.A(new_n107_), .B(new_n102_), .C(new_n77_), .D(\a[24] ), .Y(new_n776_));
  OAI21X1  g00712(.A0(new_n131_), .A1(new_n119_), .B0(new_n776_), .Y(new_n777_));
  OAI22X1  g00713(.A0(new_n102_), .A1(new_n90_), .B0(new_n96_), .B1(new_n78_), .Y(new_n778_));
  OR4X1    g00714(.A(new_n778_), .B(new_n777_), .C(new_n775_), .D(new_n652_), .Y(new_n779_));
  OR4X1    g00715(.A(new_n496_), .B(new_n412_), .C(new_n391_), .D(new_n234_), .Y(new_n780_));
  OR4X1    g00716(.A(new_n780_), .B(new_n779_), .C(new_n333_), .D(new_n154_), .Y(new_n781_));
  OR4X1    g00717(.A(new_n781_), .B(new_n774_), .C(new_n765_), .D(new_n754_), .Y(new_n782_));
  NOR2X1   g00718(.A(new_n782_), .B(new_n727_), .Y(new_n783_));
  NOR2X1   g00719(.A(new_n783_), .B(new_n690_), .Y(new_n784_));
  OAI22X1  g00720(.A0(new_n182_), .A1(new_n79_), .B0(new_n123_), .B1(new_n108_), .Y(new_n785_));
  OAI22X1  g00721(.A0(new_n143_), .A1(new_n79_), .B0(new_n123_), .B1(new_n78_), .Y(new_n786_));
  OAI22X1  g00722(.A0(new_n148_), .A1(new_n92_), .B0(new_n143_), .B1(new_n75_), .Y(new_n787_));
  OR4X1    g00723(.A(new_n787_), .B(new_n786_), .C(new_n607_), .D(new_n569_), .Y(new_n788_));
  OR4X1    g00724(.A(new_n399_), .B(new_n243_), .C(new_n522_), .D(new_n137_), .Y(new_n789_));
  OR4X1    g00725(.A(new_n789_), .B(new_n788_), .C(new_n444_), .D(new_n785_), .Y(new_n790_));
  OR2X1    g00726(.A(new_n790_), .B(new_n764_), .Y(new_n791_));
  NOR2X1   g00727(.A(new_n90_), .B(new_n69_), .Y(new_n792_));
  NOR2X1   g00728(.A(new_n598_), .B(new_n792_), .Y(new_n793_));
  NAND2X1  g00729(.A(new_n793_), .B(new_n693_), .Y(new_n794_));
  OAI21X1  g00730(.A0(new_n161_), .A1(new_n115_), .B0(new_n749_), .Y(new_n795_));
  NOR2X1   g00731(.A(new_n795_), .B(new_n755_), .Y(new_n796_));
  NOR2X1   g00732(.A(new_n105_), .B(new_n115_), .Y(new_n797_));
  NOR3X1   g00733(.A(new_n354_), .B(new_n797_), .C(new_n194_), .Y(new_n798_));
  OAI22X1  g00734(.A0(new_n125_), .A1(new_n91_), .B0(new_n119_), .B1(new_n92_), .Y(new_n799_));
  NOR3X1   g00735(.A(new_n799_), .B(new_n156_), .C(new_n521_), .Y(new_n800_));
  NAND3X1  g00736(.A(new_n800_), .B(new_n798_), .C(new_n796_), .Y(new_n801_));
  OR2X1    g00737(.A(new_n566_), .B(new_n103_), .Y(new_n802_));
  AOI21X1  g00738(.A0(new_n123_), .A1(new_n79_), .B0(new_n81_), .Y(new_n803_));
  INVX1    g00739(.A(new_n199_), .Y(new_n804_));
  INVX1    g00740(.A(new_n455_), .Y(new_n805_));
  NOR2X1   g00741(.A(new_n127_), .B(new_n115_), .Y(new_n806_));
  INVX1    g00742(.A(new_n806_), .Y(new_n807_));
  NAND3X1  g00743(.A(new_n807_), .B(new_n805_), .C(new_n804_), .Y(new_n808_));
  OR4X1    g00744(.A(new_n808_), .B(new_n803_), .C(new_n802_), .D(new_n239_), .Y(new_n809_));
  OR4X1    g00745(.A(new_n809_), .B(new_n801_), .C(new_n794_), .D(new_n791_), .Y(new_n810_));
  OR4X1    g00746(.A(new_n460_), .B(new_n483_), .C(new_n323_), .D(new_n293_), .Y(new_n811_));
  NOR2X1   g00747(.A(new_n129_), .B(new_n79_), .Y(new_n812_));
  OR4X1    g00748(.A(new_n812_), .B(new_n173_), .C(new_n426_), .D(new_n303_), .Y(new_n813_));
  NOR2X1   g00749(.A(new_n131_), .B(new_n91_), .Y(new_n814_));
  NOR2X1   g00750(.A(new_n88_), .B(new_n72_), .Y(new_n815_));
  OR4X1    g00751(.A(new_n815_), .B(new_n429_), .C(new_n814_), .D(new_n307_), .Y(new_n816_));
  INVX1    g00752(.A(new_n139_), .Y(new_n817_));
  OR2X1    g00753(.A(new_n182_), .B(new_n106_), .Y(new_n818_));
  NOR2X1   g00754(.A(new_n99_), .B(new_n91_), .Y(new_n819_));
  INVX1    g00755(.A(new_n819_), .Y(new_n820_));
  NAND4X1  g00756(.A(new_n413_), .B(new_n820_), .C(new_n818_), .D(new_n817_), .Y(new_n821_));
  OR4X1    g00757(.A(new_n821_), .B(new_n816_), .C(new_n813_), .D(new_n811_), .Y(new_n822_));
  OAI22X1  g00758(.A0(new_n127_), .A1(new_n79_), .B0(new_n123_), .B1(new_n99_), .Y(new_n823_));
  OR4X1    g00759(.A(new_n823_), .B(new_n304_), .C(new_n648_), .D(new_n379_), .Y(new_n824_));
  NOR2X1   g00760(.A(new_n182_), .B(new_n148_), .Y(new_n825_));
  OR4X1    g00761(.A(new_n459_), .B(new_n681_), .C(new_n159_), .D(new_n155_), .Y(new_n826_));
  OAI22X1  g00762(.A0(new_n168_), .A1(new_n129_), .B0(new_n106_), .B1(new_n78_), .Y(new_n827_));
  OR4X1    g00763(.A(new_n827_), .B(new_n826_), .C(new_n825_), .D(new_n581_), .Y(new_n828_));
  OAI22X1  g00764(.A0(new_n115_), .A1(new_n94_), .B0(new_n96_), .B1(new_n90_), .Y(new_n829_));
  OAI22X1  g00765(.A0(new_n182_), .A1(new_n84_), .B0(new_n143_), .B1(new_n69_), .Y(new_n830_));
  OAI22X1  g00766(.A0(new_n148_), .A1(new_n143_), .B0(new_n129_), .B1(new_n75_), .Y(new_n831_));
  OR4X1    g00767(.A(new_n831_), .B(new_n830_), .C(new_n829_), .D(new_n828_), .Y(new_n832_));
  NOR2X1   g00768(.A(new_n365_), .B(new_n233_), .Y(new_n833_));
  INVX1    g00769(.A(new_n833_), .Y(new_n834_));
  OAI22X1  g00770(.A0(new_n182_), .A1(new_n96_), .B0(new_n99_), .B1(new_n88_), .Y(new_n835_));
  OR4X1    g00771(.A(new_n835_), .B(new_n834_), .C(new_n477_), .D(new_n431_), .Y(new_n836_));
  AOI21X1  g00772(.A0(new_n84_), .A1(new_n69_), .B0(new_n81_), .Y(new_n837_));
  OAI21X1  g00773(.A0(new_n182_), .A1(new_n123_), .B0(new_n214_), .Y(new_n838_));
  OR4X1    g00774(.A(new_n838_), .B(new_n561_), .C(new_n550_), .D(new_n837_), .Y(new_n839_));
  NOR4X1   g00775(.A(new_n168_), .B(new_n198_), .C(new_n89_), .D(\a[23] ), .Y(new_n840_));
  NOR4X1   g00776(.A(new_n840_), .B(new_n328_), .C(new_n247_), .D(new_n219_), .Y(new_n841_));
  INVX1    g00777(.A(new_n841_), .Y(new_n842_));
  NOR2X1   g00778(.A(new_n152_), .B(new_n99_), .Y(new_n843_));
  OR4X1    g00779(.A(new_n702_), .B(new_n396_), .C(new_n843_), .D(new_n261_), .Y(new_n844_));
  OR4X1    g00780(.A(new_n844_), .B(new_n842_), .C(new_n839_), .D(new_n836_), .Y(new_n845_));
  OR4X1    g00781(.A(new_n845_), .B(new_n832_), .C(new_n824_), .D(new_n822_), .Y(new_n846_));
  NOR2X1   g00782(.A(new_n846_), .B(new_n810_), .Y(new_n847_));
  NOR2X1   g00783(.A(new_n99_), .B(new_n88_), .Y(new_n848_));
  OR4X1    g00784(.A(new_n848_), .B(new_n527_), .C(new_n815_), .D(new_n259_), .Y(new_n849_));
  NOR2X1   g00785(.A(new_n129_), .B(new_n96_), .Y(new_n850_));
  OR4X1    g00786(.A(new_n263_), .B(new_n850_), .C(new_n648_), .D(new_n116_), .Y(new_n851_));
  OR4X1    g00787(.A(new_n851_), .B(new_n849_), .C(new_n642_), .D(new_n843_), .Y(new_n852_));
  NOR4X1   g00788(.A(new_n543_), .B(new_n812_), .C(new_n177_), .D(new_n431_), .Y(new_n853_));
  NOR3X1   g00789(.A(new_n489_), .B(new_n256_), .C(new_n232_), .Y(new_n854_));
  NOR2X1   g00790(.A(new_n741_), .B(new_n524_), .Y(new_n855_));
  NAND4X1  g00791(.A(new_n855_), .B(new_n854_), .C(new_n853_), .D(new_n611_), .Y(new_n856_));
  OAI22X1  g00792(.A0(new_n127_), .A1(new_n75_), .B0(new_n119_), .B1(new_n90_), .Y(new_n857_));
  OR4X1    g00793(.A(new_n857_), .B(new_n694_), .C(new_n506_), .D(new_n717_), .Y(new_n858_));
  NOR4X1   g00794(.A(new_n858_), .B(new_n856_), .C(new_n852_), .D(new_n373_), .Y(new_n859_));
  INVX1    g00795(.A(new_n859_), .Y(new_n860_));
  INVX1    g00796(.A(new_n418_), .Y(new_n861_));
  INVX1    g00797(.A(new_n546_), .Y(new_n862_));
  NAND3X1  g00798(.A(new_n862_), .B(new_n861_), .C(new_n467_), .Y(new_n863_));
  OR4X1    g00799(.A(new_n579_), .B(new_n578_), .C(new_n457_), .D(new_n449_), .Y(new_n864_));
  OR4X1    g00800(.A(new_n864_), .B(new_n356_), .C(new_n350_), .D(new_n296_), .Y(new_n865_));
  OR2X1    g00801(.A(new_n865_), .B(new_n863_), .Y(new_n866_));
  OAI22X1  g00802(.A0(new_n182_), .A1(new_n168_), .B0(new_n115_), .B1(new_n92_), .Y(new_n867_));
  OR2X1    g00803(.A(new_n867_), .B(new_n280_), .Y(new_n868_));
  NOR2X1   g00804(.A(new_n90_), .B(new_n79_), .Y(new_n869_));
  OR4X1    g00805(.A(new_n869_), .B(new_n412_), .C(new_n396_), .D(new_n294_), .Y(new_n870_));
  OR4X1    g00806(.A(new_n870_), .B(new_n224_), .C(new_n213_), .D(new_n209_), .Y(new_n871_));
  OR2X1    g00807(.A(new_n871_), .B(new_n868_), .Y(new_n872_));
  OR2X1    g00808(.A(new_n387_), .B(new_n758_), .Y(new_n873_));
  OAI22X1  g00809(.A0(new_n182_), .A1(new_n96_), .B0(new_n105_), .B1(new_n88_), .Y(new_n874_));
  OAI22X1  g00810(.A0(new_n182_), .A1(new_n88_), .B0(new_n105_), .B1(new_n84_), .Y(new_n875_));
  OR4X1    g00811(.A(new_n875_), .B(new_n874_), .C(new_n873_), .D(new_n571_), .Y(new_n876_));
  NOR2X1   g00812(.A(new_n480_), .B(new_n114_), .Y(new_n877_));
  INVX1    g00813(.A(new_n877_), .Y(new_n878_));
  OR4X1    g00814(.A(new_n559_), .B(new_n516_), .C(new_n487_), .D(new_n878_), .Y(new_n879_));
  OR4X1    g00815(.A(new_n879_), .B(new_n876_), .C(new_n872_), .D(new_n866_), .Y(new_n880_));
  OAI22X1  g00816(.A0(new_n129_), .A1(new_n119_), .B0(new_n106_), .B1(new_n99_), .Y(new_n881_));
  AOI21X1  g00817(.A0(new_n96_), .A1(new_n69_), .B0(new_n99_), .Y(new_n882_));
  OR4X1    g00818(.A(new_n882_), .B(new_n881_), .C(new_n803_), .D(new_n422_), .Y(new_n883_));
  NOR2X1   g00819(.A(new_n92_), .B(new_n84_), .Y(new_n884_));
  NOR2X1   g00820(.A(new_n168_), .B(new_n161_), .Y(new_n885_));
  OR4X1    g00821(.A(new_n806_), .B(new_n885_), .C(new_n379_), .D(new_n884_), .Y(new_n886_));
  OAI22X1  g00822(.A0(new_n148_), .A1(new_n127_), .B0(new_n102_), .B1(new_n78_), .Y(new_n887_));
  OR4X1    g00823(.A(new_n887_), .B(new_n886_), .C(new_n219_), .D(new_n184_), .Y(new_n888_));
  OR4X1    g00824(.A(new_n888_), .B(new_n786_), .C(new_n652_), .D(new_n93_), .Y(new_n889_));
  OR4X1    g00825(.A(new_n586_), .B(new_n612_), .C(new_n414_), .D(new_n286_), .Y(new_n890_));
  AOI21X1  g00826(.A0(new_n161_), .A1(new_n94_), .B0(new_n91_), .Y(new_n891_));
  OAI22X1  g00827(.A0(new_n148_), .A1(new_n129_), .B0(new_n94_), .B1(new_n79_), .Y(new_n892_));
  OR4X1    g00828(.A(new_n892_), .B(new_n891_), .C(new_n187_), .D(new_n581_), .Y(new_n893_));
  OR2X1    g00829(.A(new_n893_), .B(new_n890_), .Y(new_n894_));
  NOR2X1   g00830(.A(new_n301_), .B(new_n200_), .Y(new_n895_));
  INVX1    g00831(.A(new_n895_), .Y(new_n896_));
  OR2X1    g00832(.A(new_n498_), .B(new_n191_), .Y(new_n897_));
  OR4X1    g00833(.A(new_n681_), .B(new_n285_), .C(new_n201_), .D(new_n176_), .Y(new_n898_));
  OR4X1    g00834(.A(new_n898_), .B(new_n897_), .C(new_n896_), .D(new_n382_), .Y(new_n899_));
  OR4X1    g00835(.A(new_n899_), .B(new_n894_), .C(new_n889_), .D(new_n883_), .Y(new_n900_));
  OR2X1    g00836(.A(new_n900_), .B(new_n880_), .Y(new_n901_));
  OAI22X1  g00837(.A0(new_n901_), .A1(new_n860_), .B0(new_n846_), .B1(new_n810_), .Y(new_n902_));
  NOR2X1   g00838(.A(new_n901_), .B(new_n860_), .Y(new_n903_));
  OAI22X1  g00839(.A0(new_n143_), .A1(new_n119_), .B0(new_n105_), .B1(new_n84_), .Y(new_n904_));
  OAI22X1  g00840(.A0(new_n148_), .A1(new_n131_), .B0(new_n108_), .B1(new_n115_), .Y(new_n905_));
  OR4X1    g00841(.A(new_n905_), .B(new_n904_), .C(new_n226_), .D(new_n338_), .Y(new_n906_));
  OAI22X1  g00842(.A0(new_n129_), .A1(new_n119_), .B0(new_n106_), .B1(new_n90_), .Y(new_n907_));
  OR2X1    g00843(.A(new_n907_), .B(new_n757_), .Y(new_n908_));
  OR4X1    g00844(.A(new_n632_), .B(new_n385_), .C(new_n819_), .D(new_n245_), .Y(new_n909_));
  OR4X1    g00845(.A(new_n541_), .B(new_n574_), .C(new_n265_), .D(new_n173_), .Y(new_n910_));
  OR4X1    g00846(.A(new_n910_), .B(new_n909_), .C(new_n908_), .D(new_n906_), .Y(new_n911_));
  OAI22X1  g00847(.A0(new_n123_), .A1(new_n72_), .B0(new_n108_), .B1(new_n96_), .Y(new_n912_));
  OR4X1    g00848(.A(new_n912_), .B(new_n523_), .C(new_n246_), .D(new_n85_), .Y(new_n913_));
  NOR4X1   g00849(.A(new_n913_), .B(new_n506_), .C(new_n301_), .D(new_n196_), .Y(new_n914_));
  INVX1    g00850(.A(new_n914_), .Y(new_n915_));
  OR4X1    g00851(.A(new_n627_), .B(new_n299_), .C(new_n280_), .D(new_n539_), .Y(new_n916_));
  OR4X1    g00852(.A(new_n724_), .B(new_n603_), .C(new_n304_), .D(new_n535_), .Y(new_n917_));
  OR4X1    g00853(.A(new_n917_), .B(new_n500_), .C(new_n206_), .D(new_n202_), .Y(new_n918_));
  OR4X1    g00854(.A(new_n918_), .B(new_n916_), .C(new_n641_), .D(new_n785_), .Y(new_n919_));
  OR4X1    g00855(.A(new_n772_), .B(new_n393_), .C(new_n231_), .D(new_n209_), .Y(new_n920_));
  AOI21X1  g00856(.A0(new_n129_), .A1(new_n99_), .B0(new_n96_), .Y(new_n921_));
  OR4X1    g00857(.A(new_n921_), .B(new_n920_), .C(new_n823_), .D(new_n768_), .Y(new_n922_));
  NOR4X1   g00858(.A(new_n922_), .B(new_n919_), .C(new_n915_), .D(new_n911_), .Y(new_n923_));
  AOI21X1  g00859(.A0(new_n92_), .A1(new_n81_), .B0(new_n102_), .Y(new_n924_));
  OR4X1    g00860(.A(new_n924_), .B(new_n510_), .C(new_n207_), .D(new_n426_), .Y(new_n925_));
  OAI22X1  g00861(.A0(new_n161_), .A1(new_n91_), .B0(new_n106_), .B1(new_n72_), .Y(new_n926_));
  OR2X1    g00862(.A(new_n926_), .B(new_n797_), .Y(new_n927_));
  NOR2X1   g00863(.A(new_n129_), .B(new_n106_), .Y(new_n928_));
  OR4X1    g00864(.A(new_n843_), .B(new_n200_), .C(new_n159_), .D(new_n928_), .Y(new_n929_));
  OR4X1    g00865(.A(new_n168_), .B(new_n101_), .C(new_n89_), .D(\a[23] ), .Y(new_n930_));
  OAI21X1  g00866(.A0(new_n182_), .A1(new_n115_), .B0(new_n930_), .Y(new_n931_));
  OR4X1    g00867(.A(new_n931_), .B(new_n803_), .C(new_n586_), .D(new_n494_), .Y(new_n932_));
  OR4X1    g00868(.A(new_n932_), .B(new_n929_), .C(new_n927_), .D(new_n925_), .Y(new_n933_));
  OR4X1    g00869(.A(new_n329_), .B(new_n825_), .C(new_n746_), .D(new_n651_), .Y(new_n934_));
  AOI21X1  g00870(.A0(new_n148_), .A1(new_n115_), .B0(new_n90_), .Y(new_n935_));
  OR4X1    g00871(.A(new_n935_), .B(new_n934_), .C(new_n414_), .D(new_n691_), .Y(new_n936_));
  OR4X1    g00872(.A(new_n936_), .B(new_n679_), .C(new_n356_), .D(new_n423_), .Y(new_n937_));
  NOR2X1   g00873(.A(new_n129_), .B(new_n117_), .Y(new_n938_));
  OR4X1    g00874(.A(new_n938_), .B(new_n505_), .C(new_n565_), .D(new_n223_), .Y(new_n939_));
  OR4X1    g00875(.A(new_n292_), .B(new_n134_), .C(new_n120_), .D(new_n307_), .Y(new_n940_));
  OR4X1    g00876(.A(new_n940_), .B(new_n433_), .C(new_n483_), .D(new_n219_), .Y(new_n941_));
  OR4X1    g00877(.A(new_n941_), .B(new_n939_), .C(new_n937_), .D(new_n933_), .Y(new_n942_));
  OR4X1    g00878(.A(new_n634_), .B(new_n372_), .C(new_n228_), .D(new_n100_), .Y(new_n943_));
  OR4X1    g00879(.A(new_n612_), .B(new_n256_), .C(new_n160_), .D(new_n337_), .Y(new_n944_));
  OAI22X1  g00880(.A0(new_n152_), .A1(new_n129_), .B0(new_n84_), .B1(new_n78_), .Y(new_n945_));
  OR2X1    g00881(.A(new_n945_), .B(new_n263_), .Y(new_n946_));
  OAI22X1  g00882(.A0(new_n143_), .A1(new_n75_), .B0(new_n108_), .B1(new_n91_), .Y(new_n947_));
  NOR3X1   g00883(.A(new_n947_), .B(new_n504_), .C(new_n382_), .Y(new_n948_));
  INVX1    g00884(.A(new_n948_), .Y(new_n949_));
  OR4X1    g00885(.A(new_n949_), .B(new_n946_), .C(new_n944_), .D(new_n943_), .Y(new_n950_));
  OAI22X1  g00886(.A0(new_n161_), .A1(new_n84_), .B0(new_n119_), .B1(new_n105_), .Y(new_n951_));
  OR4X1    g00887(.A(new_n951_), .B(new_n629_), .C(new_n243_), .D(new_n133_), .Y(new_n952_));
  OR4X1    g00888(.A(new_n363_), .B(new_n282_), .C(new_n240_), .D(new_n222_), .Y(new_n953_));
  OR4X1    g00889(.A(new_n953_), .B(new_n952_), .C(new_n950_), .D(new_n836_), .Y(new_n954_));
  NOR2X1   g00890(.A(new_n954_), .B(new_n942_), .Y(new_n955_));
  AOI21X1  g00891(.A0(new_n955_), .A1(new_n923_), .B0(new_n903_), .Y(new_n956_));
  AND2X1   g00892(.A(new_n955_), .B(new_n923_), .Y(new_n957_));
  OR4X1    g00893(.A(new_n823_), .B(new_n429_), .C(new_n691_), .D(new_n398_), .Y(new_n958_));
  AOI21X1  g00894(.A0(new_n91_), .A1(new_n69_), .B0(new_n94_), .Y(new_n959_));
  OR4X1    g00895(.A(new_n959_), .B(new_n921_), .C(new_n640_), .D(new_n272_), .Y(new_n960_));
  OR2X1    g00896(.A(new_n960_), .B(new_n696_), .Y(new_n961_));
  NOR3X1   g00897(.A(new_n393_), .B(new_n385_), .C(new_n806_), .Y(new_n962_));
  NOR4X1   g00898(.A(new_n356_), .B(new_n294_), .C(new_n264_), .D(new_n184_), .Y(new_n963_));
  NOR4X1   g00899(.A(new_n191_), .B(new_n825_), .C(new_n792_), .D(new_n103_), .Y(new_n964_));
  NAND3X1  g00900(.A(new_n964_), .B(new_n963_), .C(new_n962_), .Y(new_n965_));
  OR4X1    g00901(.A(new_n965_), .B(new_n961_), .C(new_n958_), .D(new_n774_), .Y(new_n966_));
  INVX1    g00902(.A(new_n966_), .Y(new_n967_));
  NOR2X1   g00903(.A(new_n182_), .B(new_n75_), .Y(new_n968_));
  OR4X1    g00904(.A(new_n863_), .B(new_n509_), .C(new_n968_), .D(new_n178_), .Y(new_n969_));
  OR4X1    g00905(.A(new_n594_), .B(new_n578_), .C(new_n812_), .D(new_n200_), .Y(new_n970_));
  INVX1    g00906(.A(new_n232_), .Y(new_n971_));
  INVX1    g00907(.A(new_n636_), .Y(new_n972_));
  NAND3X1  g00908(.A(new_n972_), .B(new_n345_), .C(new_n971_), .Y(new_n973_));
  INVX1    g00909(.A(new_n214_), .Y(new_n974_));
  OAI22X1  g00910(.A0(new_n161_), .A1(new_n69_), .B0(new_n123_), .B1(new_n105_), .Y(new_n975_));
  OR4X1    g00911(.A(new_n975_), .B(new_n974_), .C(new_n197_), .D(new_n76_), .Y(new_n976_));
  OR2X1    g00912(.A(new_n976_), .B(new_n310_), .Y(new_n977_));
  OR4X1    g00913(.A(new_n977_), .B(new_n973_), .C(new_n970_), .D(new_n969_), .Y(new_n978_));
  OAI22X1  g00914(.A0(new_n105_), .A1(new_n91_), .B0(new_n96_), .B1(new_n72_), .Y(new_n979_));
  OR2X1    g00915(.A(new_n979_), .B(new_n589_), .Y(new_n980_));
  NOR2X1   g00916(.A(new_n88_), .B(new_n81_), .Y(new_n981_));
  OR4X1    g00917(.A(new_n459_), .B(new_n479_), .C(new_n181_), .D(new_n981_), .Y(new_n982_));
  OR4X1    g00918(.A(new_n982_), .B(new_n980_), .C(new_n358_), .D(new_n350_), .Y(new_n983_));
  NOR4X1   g00919(.A(new_n983_), .B(new_n978_), .C(new_n954_), .D(new_n781_), .Y(new_n984_));
  AND2X1   g00920(.A(new_n984_), .B(new_n967_), .Y(new_n985_));
  OR2X1    g00921(.A(new_n985_), .B(new_n957_), .Y(new_n986_));
  INVX1    g00922(.A(new_n356_), .Y(new_n987_));
  INVX1    g00923(.A(new_n702_), .Y(new_n988_));
  INVX1    g00924(.A(new_n632_), .Y(new_n989_));
  NAND3X1  g00925(.A(new_n989_), .B(new_n988_), .C(new_n987_), .Y(new_n990_));
  NOR2X1   g00926(.A(new_n292_), .B(new_n291_), .Y(new_n991_));
  INVX1    g00927(.A(new_n991_), .Y(new_n992_));
  OAI22X1  g00928(.A0(new_n102_), .A1(new_n72_), .B0(new_n99_), .B1(new_n91_), .Y(new_n993_));
  OAI22X1  g00929(.A0(new_n129_), .A1(new_n91_), .B0(new_n105_), .B1(new_n102_), .Y(new_n994_));
  OR4X1    g00930(.A(new_n994_), .B(new_n993_), .C(new_n332_), .D(new_n992_), .Y(new_n995_));
  OR4X1    g00931(.A(new_n510_), .B(new_n386_), .C(new_n299_), .D(new_n203_), .Y(new_n996_));
  OR4X1    g00932(.A(new_n996_), .B(new_n995_), .C(new_n734_), .D(new_n990_), .Y(new_n997_));
  NOR2X1   g00933(.A(new_n168_), .B(new_n78_), .Y(new_n998_));
  NOR3X1   g00934(.A(new_n848_), .B(new_n358_), .C(new_n998_), .Y(new_n999_));
  OAI22X1  g00935(.A0(new_n148_), .A1(new_n92_), .B0(new_n91_), .B1(new_n81_), .Y(new_n1000_));
  NOR3X1   g00936(.A(new_n1000_), .B(new_n319_), .C(new_n806_), .Y(new_n1001_));
  AOI21X1  g00937(.A0(new_n92_), .A1(new_n72_), .B0(new_n96_), .Y(new_n1002_));
  NOR3X1   g00938(.A(new_n1002_), .B(new_n280_), .C(new_n928_), .Y(new_n1003_));
  NAND4X1  g00939(.A(new_n1003_), .B(new_n1001_), .C(new_n999_), .D(new_n476_), .Y(new_n1004_));
  OAI22X1  g00940(.A0(new_n148_), .A1(new_n78_), .B0(new_n129_), .B1(new_n84_), .Y(new_n1005_));
  AOI21X1  g00941(.A0(new_n92_), .A1(new_n81_), .B0(new_n117_), .Y(new_n1006_));
  OR4X1    g00942(.A(new_n1006_), .B(new_n1005_), .C(new_n717_), .D(new_n118_), .Y(new_n1007_));
  NOR2X1   g00943(.A(new_n108_), .B(new_n106_), .Y(new_n1008_));
  OR4X1    g00944(.A(new_n256_), .B(new_n539_), .C(new_n426_), .D(new_n1008_), .Y(new_n1009_));
  OR4X1    g00945(.A(new_n1009_), .B(new_n1007_), .C(new_n904_), .D(new_n513_), .Y(new_n1010_));
  OR4X1    g00946(.A(new_n508_), .B(new_n812_), .C(new_n296_), .D(new_n160_), .Y(new_n1011_));
  OAI22X1  g00947(.A0(new_n143_), .A1(new_n79_), .B0(new_n102_), .B1(new_n81_), .Y(new_n1012_));
  OR4X1    g00948(.A(new_n1012_), .B(new_n489_), .C(new_n408_), .D(new_n350_), .Y(new_n1013_));
  OR4X1    g00949(.A(new_n1013_), .B(new_n1011_), .C(new_n1010_), .D(new_n1004_), .Y(new_n1014_));
  OR2X1    g00950(.A(new_n1014_), .B(new_n997_), .Y(new_n1015_));
  OAI22X1  g00951(.A0(new_n182_), .A1(new_n75_), .B0(new_n96_), .B1(new_n78_), .Y(new_n1016_));
  OR2X1    g00952(.A(new_n1016_), .B(new_n612_), .Y(new_n1017_));
  OAI22X1  g00953(.A0(new_n106_), .A1(new_n99_), .B0(new_n79_), .B1(new_n72_), .Y(new_n1018_));
  OR4X1    g00954(.A(new_n480_), .B(new_n396_), .C(new_n304_), .D(new_n196_), .Y(new_n1019_));
  OR4X1    g00955(.A(new_n1019_), .B(new_n1018_), .C(new_n1017_), .D(new_n691_), .Y(new_n1020_));
  OAI22X1  g00956(.A0(new_n123_), .A1(new_n81_), .B0(new_n106_), .B1(new_n105_), .Y(new_n1021_));
  OAI22X1  g00957(.A0(new_n182_), .A1(new_n91_), .B0(new_n75_), .B1(new_n72_), .Y(new_n1022_));
  OR4X1    g00958(.A(new_n1022_), .B(new_n1021_), .C(new_n678_), .D(new_n176_), .Y(new_n1023_));
  OR4X1    g00959(.A(new_n293_), .B(new_n239_), .C(new_n139_), .D(new_n120_), .Y(new_n1024_));
  OR4X1    g00960(.A(new_n1024_), .B(new_n1023_), .C(new_n423_), .D(new_n681_), .Y(new_n1025_));
  OAI22X1  g00961(.A0(new_n168_), .A1(new_n72_), .B0(new_n161_), .B1(new_n102_), .Y(new_n1026_));
  OR2X1    g00962(.A(new_n1026_), .B(new_n224_), .Y(new_n1027_));
  NOR2X1   g00963(.A(new_n148_), .B(new_n94_), .Y(new_n1028_));
  OAI22X1  g00964(.A0(new_n152_), .A1(new_n105_), .B0(new_n125_), .B1(new_n123_), .Y(new_n1029_));
  OR4X1    g00965(.A(new_n1029_), .B(new_n1028_), .C(new_n175_), .D(new_n137_), .Y(new_n1030_));
  OR2X1    g00966(.A(new_n1030_), .B(new_n1027_), .Y(new_n1031_));
  OR4X1    g00967(.A(new_n252_), .B(new_n616_), .C(new_n220_), .D(new_n457_), .Y(new_n1032_));
  INVX1    g00968(.A(new_n337_), .Y(new_n1033_));
  INVX1    g00969(.A(new_n207_), .Y(new_n1034_));
  INVX1    g00970(.A(new_n234_), .Y(new_n1035_));
  NAND3X1  g00971(.A(new_n1035_), .B(new_n1034_), .C(new_n1033_), .Y(new_n1036_));
  OAI22X1  g00972(.A0(new_n152_), .A1(new_n131_), .B0(new_n99_), .B1(new_n96_), .Y(new_n1037_));
  OR2X1    g00973(.A(new_n1037_), .B(new_n724_), .Y(new_n1038_));
  OR4X1    g00974(.A(new_n1038_), .B(new_n1036_), .C(new_n1032_), .D(new_n945_), .Y(new_n1039_));
  NOR4X1   g00975(.A(new_n1039_), .B(new_n1031_), .C(new_n1025_), .D(new_n1020_), .Y(new_n1040_));
  INVX1    g00976(.A(new_n1040_), .Y(new_n1041_));
  NOR4X1   g00977(.A(new_n701_), .B(new_n440_), .C(new_n814_), .D(new_n227_), .Y(new_n1042_));
  NOR3X1   g00978(.A(new_n506_), .B(new_n300_), .C(new_n758_), .Y(new_n1043_));
  NOR2X1   g00979(.A(new_n182_), .B(new_n96_), .Y(new_n1044_));
  NOR3X1   g00980(.A(new_n1044_), .B(new_n869_), .C(new_n603_), .Y(new_n1045_));
  NOR2X1   g00981(.A(new_n94_), .B(new_n91_), .Y(new_n1046_));
  NOR4X1   g00982(.A(new_n197_), .B(new_n746_), .C(new_n303_), .D(new_n1046_), .Y(new_n1047_));
  NAND4X1  g00983(.A(new_n1047_), .B(new_n1045_), .C(new_n1043_), .D(new_n1042_), .Y(new_n1048_));
  AND2X1   g00984(.A(new_n345_), .B(new_n250_), .Y(new_n1049_));
  NOR4X1   g00985(.A(new_n500_), .B(new_n395_), .C(new_n354_), .D(new_n974_), .Y(new_n1050_));
  NOR4X1   g00986(.A(new_n755_), .B(new_n496_), .C(new_n246_), .D(new_n162_), .Y(new_n1051_));
  NAND3X1  g00987(.A(new_n1051_), .B(new_n1050_), .C(new_n1049_), .Y(new_n1052_));
  NOR3X1   g00988(.A(new_n98_), .B(new_n68_), .C(\a[29] ), .Y(new_n1053_));
  NOR3X1   g00989(.A(new_n107_), .B(new_n77_), .C(\a[24] ), .Y(new_n1054_));
  NOR3X1   g00990(.A(new_n198_), .B(new_n89_), .C(\a[23] ), .Y(new_n1055_));
  AOI22X1  g00991(.A0(new_n557_), .A1(new_n1054_), .B0(new_n1055_), .B1(new_n1053_), .Y(new_n1056_));
  INVX1    g00992(.A(new_n1056_), .Y(new_n1057_));
  OR4X1    g00993(.A(new_n586_), .B(new_n460_), .C(new_n429_), .D(new_n240_), .Y(new_n1058_));
  OR4X1    g00994(.A(new_n232_), .B(new_n223_), .C(new_n535_), .D(new_n390_), .Y(new_n1059_));
  OR4X1    g00995(.A(new_n1059_), .B(new_n1058_), .C(new_n823_), .D(new_n1057_), .Y(new_n1060_));
  OAI22X1  g00996(.A0(new_n148_), .A1(new_n99_), .B0(new_n119_), .B1(new_n105_), .Y(new_n1061_));
  OAI22X1  g00997(.A0(new_n115_), .A1(new_n78_), .B0(new_n90_), .B1(new_n69_), .Y(new_n1062_));
  OR4X1    g00998(.A(new_n1062_), .B(new_n1061_), .C(new_n843_), .D(new_n282_), .Y(new_n1063_));
  OR4X1    g00999(.A(new_n1063_), .B(new_n1060_), .C(new_n1052_), .D(new_n745_), .Y(new_n1064_));
  NOR4X1   g01000(.A(new_n1064_), .B(new_n1048_), .C(new_n1041_), .D(new_n1015_), .Y(new_n1065_));
  AOI21X1  g01001(.A0(new_n984_), .A1(new_n967_), .B0(new_n1065_), .Y(new_n1066_));
  OAI22X1  g01002(.A0(new_n143_), .A1(new_n117_), .B0(new_n90_), .B1(new_n84_), .Y(new_n1067_));
  OR4X1    g01003(.A(new_n1067_), .B(new_n931_), .C(new_n819_), .D(new_n137_), .Y(new_n1068_));
  OR4X1    g01004(.A(new_n228_), .B(new_n224_), .C(new_n664_), .D(new_n521_), .Y(new_n1069_));
  OR2X1    g01005(.A(new_n127_), .B(new_n91_), .Y(new_n1070_));
  OR2X1    g01006(.A(new_n168_), .B(new_n161_), .Y(new_n1071_));
  NAND3X1  g01007(.A(new_n590_), .B(new_n1071_), .C(new_n1070_), .Y(new_n1072_));
  OR4X1    g01008(.A(new_n1072_), .B(new_n1069_), .C(new_n1068_), .D(new_n970_), .Y(new_n1073_));
  OAI22X1  g01009(.A0(new_n99_), .A1(new_n84_), .B0(new_n79_), .B1(new_n78_), .Y(new_n1074_));
  OR2X1    g01010(.A(new_n1074_), .B(new_n354_), .Y(new_n1075_));
  NOR3X1   g01011(.A(new_n239_), .B(new_n199_), .C(new_n173_), .Y(new_n1076_));
  INVX1    g01012(.A(new_n1076_), .Y(new_n1077_));
  AOI21X1  g01013(.A0(new_n125_), .A1(new_n94_), .B0(new_n119_), .Y(new_n1078_));
  OR2X1    g01014(.A(new_n1078_), .B(new_n395_), .Y(new_n1079_));
  OR4X1    g01015(.A(new_n1079_), .B(new_n1077_), .C(new_n1075_), .D(new_n927_), .Y(new_n1080_));
  OR4X1    g01016(.A(new_n945_), .B(new_n938_), .C(new_n743_), .D(new_n547_), .Y(new_n1081_));
  NOR2X1   g01017(.A(new_n182_), .B(new_n88_), .Y(new_n1082_));
  OR4X1    g01018(.A(new_n265_), .B(new_n264_), .C(new_n479_), .D(new_n338_), .Y(new_n1083_));
  OR4X1    g01019(.A(new_n1083_), .B(new_n1082_), .C(new_n385_), .D(new_n785_), .Y(new_n1084_));
  OR4X1    g01020(.A(new_n1084_), .B(new_n1081_), .C(new_n1080_), .D(new_n1073_), .Y(new_n1085_));
  NOR3X1   g01021(.A(new_n1085_), .B(new_n834_), .C(new_n758_), .Y(new_n1086_));
  NOR2X1   g01022(.A(new_n143_), .B(new_n119_), .Y(new_n1087_));
  NOR3X1   g01023(.A(new_n968_), .B(new_n1087_), .C(new_n610_), .Y(new_n1088_));
  OR4X1    g01024(.A(new_n741_), .B(new_n400_), .C(new_n220_), .D(new_n187_), .Y(new_n1089_));
  OAI22X1  g01025(.A0(new_n152_), .A1(new_n143_), .B0(new_n131_), .B1(new_n117_), .Y(new_n1090_));
  NOR4X1   g01026(.A(new_n1090_), .B(new_n1089_), .C(new_n632_), .D(new_n357_), .Y(new_n1091_));
  NAND2X1  g01027(.A(new_n1091_), .B(new_n1088_), .Y(new_n1092_));
  NOR2X1   g01028(.A(new_n243_), .B(new_n133_), .Y(new_n1093_));
  INVX1    g01029(.A(new_n1093_), .Y(new_n1094_));
  OAI22X1  g01030(.A0(new_n161_), .A1(new_n75_), .B0(new_n148_), .B1(new_n94_), .Y(new_n1095_));
  OAI22X1  g01031(.A0(new_n125_), .A1(new_n123_), .B0(new_n99_), .B1(new_n88_), .Y(new_n1096_));
  OR4X1    g01032(.A(new_n1096_), .B(new_n1095_), .C(new_n504_), .D(new_n300_), .Y(new_n1097_));
  OR4X1    g01033(.A(new_n541_), .B(new_n475_), .C(new_n648_), .D(new_n126_), .Y(new_n1098_));
  OR4X1    g01034(.A(new_n1098_), .B(new_n1097_), .C(new_n1094_), .D(new_n76_), .Y(new_n1099_));
  OAI22X1  g01035(.A0(new_n161_), .A1(new_n96_), .B0(new_n94_), .B1(new_n69_), .Y(new_n1100_));
  OAI22X1  g01036(.A0(new_n106_), .A1(new_n94_), .B0(new_n90_), .B1(new_n69_), .Y(new_n1101_));
  OR4X1    g01037(.A(new_n1101_), .B(new_n1100_), .C(new_n510_), .D(new_n307_), .Y(new_n1102_));
  NOR4X1   g01038(.A(new_n1102_), .B(new_n1099_), .C(new_n1092_), .D(new_n761_), .Y(new_n1103_));
  OAI22X1  g01039(.A0(new_n161_), .A1(new_n152_), .B0(new_n129_), .B1(new_n88_), .Y(new_n1104_));
  OAI22X1  g01040(.A0(new_n127_), .A1(new_n84_), .B0(new_n99_), .B1(new_n75_), .Y(new_n1105_));
  OAI22X1  g01041(.A0(new_n168_), .A1(new_n99_), .B0(new_n143_), .B1(new_n84_), .Y(new_n1106_));
  OR4X1    g01042(.A(new_n1106_), .B(new_n1105_), .C(new_n1104_), .D(new_n1000_), .Y(new_n1107_));
  OAI22X1  g01043(.A0(new_n108_), .A1(new_n102_), .B0(new_n96_), .B1(new_n78_), .Y(new_n1108_));
  OR2X1    g01044(.A(new_n1108_), .B(new_n422_), .Y(new_n1109_));
  NOR4X1   g01045(.A(new_n755_), .B(new_n282_), .C(new_n172_), .D(new_n160_), .Y(new_n1110_));
  INVX1    g01046(.A(new_n1110_), .Y(new_n1111_));
  OR4X1    g01047(.A(new_n596_), .B(new_n840_), .C(new_n423_), .D(new_n746_), .Y(new_n1112_));
  NOR4X1   g01048(.A(new_n1112_), .B(new_n1111_), .C(new_n1109_), .D(new_n1107_), .Y(new_n1113_));
  AOI21X1  g01049(.A0(new_n131_), .A1(new_n92_), .B0(new_n88_), .Y(new_n1114_));
  OR4X1    g01050(.A(new_n806_), .B(new_n184_), .C(new_n180_), .D(new_n327_), .Y(new_n1115_));
  OR4X1    g01051(.A(new_n500_), .B(new_n301_), .C(new_n201_), .D(new_n757_), .Y(new_n1116_));
  OR4X1    g01052(.A(new_n1116_), .B(new_n603_), .C(new_n493_), .D(new_n379_), .Y(new_n1117_));
  OAI22X1  g01053(.A0(new_n131_), .A1(new_n91_), .B0(new_n102_), .B1(new_n78_), .Y(new_n1118_));
  OAI22X1  g01054(.A0(new_n168_), .A1(new_n129_), .B0(new_n152_), .B1(new_n127_), .Y(new_n1119_));
  NOR3X1   g01055(.A(new_n1119_), .B(new_n1118_), .C(new_n333_), .Y(new_n1120_));
  NOR4X1   g01056(.A(new_n720_), .B(new_n642_), .C(new_n505_), .D(new_n497_), .Y(new_n1121_));
  NOR4X1   g01057(.A(new_n387_), .B(new_n372_), .C(new_n293_), .D(new_n206_), .Y(new_n1122_));
  NAND3X1  g01058(.A(new_n1122_), .B(new_n1121_), .C(new_n1120_), .Y(new_n1123_));
  NOR4X1   g01059(.A(new_n1123_), .B(new_n1117_), .C(new_n1115_), .D(new_n1114_), .Y(new_n1124_));
  AND2X1   g01060(.A(new_n1124_), .B(new_n1113_), .Y(new_n1125_));
  NAND3X1  g01061(.A(new_n1125_), .B(new_n1103_), .C(new_n1086_), .Y(new_n1126_));
  INVX1    g01062(.A(new_n1126_), .Y(new_n1127_));
  OR4X1    g01063(.A(new_n391_), .B(new_n387_), .C(new_n234_), .D(new_n439_), .Y(new_n1128_));
  INVX1    g01064(.A(new_n142_), .Y(new_n1129_));
  INVX1    g01065(.A(new_n328_), .Y(new_n1130_));
  NAND3X1  g01066(.A(new_n1130_), .B(new_n380_), .C(new_n1129_), .Y(new_n1131_));
  OR4X1    g01067(.A(new_n1131_), .B(new_n1128_), .C(new_n1018_), .D(new_n691_), .Y(new_n1132_));
  INVX1    g01068(.A(new_n1049_), .Y(new_n1133_));
  AOI21X1  g01069(.A0(new_n96_), .A1(new_n75_), .B0(new_n81_), .Y(new_n1134_));
  OAI22X1  g01070(.A0(new_n148_), .A1(new_n129_), .B0(new_n90_), .B1(new_n75_), .Y(new_n1135_));
  AOI21X1  g01071(.A0(new_n115_), .A1(new_n91_), .B0(new_n125_), .Y(new_n1136_));
  OR4X1    g01072(.A(new_n1136_), .B(new_n1135_), .C(new_n1134_), .D(new_n710_), .Y(new_n1137_));
  OR4X1    g01073(.A(new_n565_), .B(new_n423_), .C(new_n578_), .D(new_n457_), .Y(new_n1138_));
  OR4X1    g01074(.A(new_n1138_), .B(new_n1137_), .C(new_n1133_), .D(new_n531_), .Y(new_n1139_));
  OAI22X1  g01075(.A0(new_n152_), .A1(new_n131_), .B0(new_n143_), .B1(new_n117_), .Y(new_n1140_));
  OR4X1    g01076(.A(new_n1140_), .B(new_n385_), .C(new_n286_), .D(new_n200_), .Y(new_n1141_));
  AOI21X1  g01077(.A0(new_n125_), .A1(new_n105_), .B0(new_n79_), .Y(new_n1142_));
  OR4X1    g01078(.A(new_n1142_), .B(new_n321_), .C(new_n536_), .D(new_n522_), .Y(new_n1143_));
  OR2X1    g01079(.A(new_n1143_), .B(new_n1141_), .Y(new_n1144_));
  NOR4X1   g01080(.A(new_n1144_), .B(new_n1139_), .C(new_n1132_), .D(new_n1048_), .Y(new_n1145_));
  AOI21X1  g01081(.A0(new_n79_), .A1(new_n69_), .B0(new_n92_), .Y(new_n1146_));
  OR2X1    g01082(.A(new_n1146_), .B(new_n723_), .Y(new_n1147_));
  OR4X1    g01083(.A(new_n678_), .B(new_n850_), .C(new_n231_), .D(new_n337_), .Y(new_n1148_));
  NOR4X1   g01084(.A(new_n1148_), .B(new_n1147_), .C(new_n1102_), .D(new_n485_), .Y(new_n1149_));
  INVX1    g01085(.A(new_n259_), .Y(new_n1150_));
  INVX1    g01086(.A(new_n408_), .Y(new_n1151_));
  INVX1    g01087(.A(new_n679_), .Y(new_n1152_));
  NAND3X1  g01088(.A(new_n1152_), .B(new_n1151_), .C(new_n1150_), .Y(new_n1153_));
  OR4X1    g01089(.A(new_n509_), .B(new_n574_), .C(new_n806_), .D(new_n455_), .Y(new_n1154_));
  NOR4X1   g01090(.A(new_n1154_), .B(new_n1153_), .C(new_n176_), .D(new_n116_), .Y(new_n1155_));
  OAI22X1  g01091(.A0(new_n161_), .A1(new_n148_), .B0(new_n123_), .B1(new_n94_), .Y(new_n1156_));
  OAI22X1  g01092(.A0(new_n108_), .A1(new_n91_), .B0(new_n75_), .B1(new_n72_), .Y(new_n1157_));
  AOI21X1  g01093(.A0(new_n129_), .A1(new_n72_), .B0(new_n91_), .Y(new_n1158_));
  OAI22X1  g01094(.A0(new_n117_), .A1(new_n72_), .B0(new_n115_), .B1(new_n90_), .Y(new_n1159_));
  OR4X1    g01095(.A(new_n1159_), .B(new_n1158_), .C(new_n1157_), .D(new_n1156_), .Y(new_n1160_));
  INVX1    g01096(.A(new_n581_), .Y(new_n1161_));
  INVX1    g01097(.A(new_n285_), .Y(new_n1162_));
  NAND3X1  g01098(.A(new_n721_), .B(new_n1162_), .C(new_n1161_), .Y(new_n1163_));
  NOR3X1   g01099(.A(new_n543_), .B(new_n974_), .C(new_n173_), .Y(new_n1164_));
  INVX1    g01100(.A(new_n1164_), .Y(new_n1165_));
  NOR2X1   g01101(.A(new_n182_), .B(new_n117_), .Y(new_n1166_));
  OR4X1    g01102(.A(new_n1166_), .B(new_n358_), .C(new_n356_), .D(new_n681_), .Y(new_n1167_));
  NOR4X1   g01103(.A(new_n1167_), .B(new_n1165_), .C(new_n1163_), .D(new_n1160_), .Y(new_n1168_));
  NAND3X1  g01104(.A(new_n1168_), .B(new_n1155_), .C(new_n1149_), .Y(new_n1169_));
  INVX1    g01105(.A(new_n1169_), .Y(new_n1170_));
  OAI22X1  g01106(.A0(new_n131_), .A1(new_n69_), .B0(new_n108_), .B1(new_n96_), .Y(new_n1171_));
  OAI22X1  g01107(.A0(new_n105_), .A1(new_n75_), .B0(new_n88_), .B1(new_n72_), .Y(new_n1172_));
  OAI21X1  g01108(.A0(new_n106_), .A1(new_n92_), .B0(new_n551_), .Y(new_n1173_));
  NOR4X1   g01109(.A(new_n1173_), .B(new_n1172_), .C(new_n1171_), .D(new_n1095_), .Y(new_n1174_));
  NOR3X1   g01110(.A(new_n527_), .B(new_n540_), .C(new_n124_), .Y(new_n1175_));
  NOR3X1   g01111(.A(new_n155_), .B(new_n141_), .C(new_n521_), .Y(new_n1176_));
  NOR3X1   g01112(.A(new_n514_), .B(new_n410_), .C(new_n162_), .Y(new_n1177_));
  NAND4X1  g01113(.A(new_n1177_), .B(new_n1176_), .C(new_n1175_), .D(new_n1174_), .Y(new_n1178_));
  OR4X1    g01114(.A(new_n596_), .B(new_n498_), .C(new_n417_), .D(new_n494_), .Y(new_n1179_));
  OR4X1    g01115(.A(new_n1179_), .B(new_n496_), .C(new_n350_), .D(new_n233_), .Y(new_n1180_));
  NOR4X1   g01116(.A(new_n504_), .B(new_n412_), .C(new_n819_), .D(new_n177_), .Y(new_n1181_));
  NOR4X1   g01117(.A(new_n199_), .B(new_n181_), .C(new_n884_), .D(new_n86_), .Y(new_n1182_));
  OAI22X1  g01118(.A0(new_n182_), .A1(new_n119_), .B0(new_n148_), .B1(new_n105_), .Y(new_n1183_));
  NOR3X1   g01119(.A(new_n1183_), .B(new_n493_), .C(new_n149_), .Y(new_n1184_));
  NAND3X1  g01120(.A(new_n1184_), .B(new_n1182_), .C(new_n1181_), .Y(new_n1185_));
  NOR4X1   g01121(.A(new_n1185_), .B(new_n1180_), .C(new_n1178_), .D(new_n650_), .Y(new_n1186_));
  NAND3X1  g01122(.A(new_n1186_), .B(new_n1170_), .C(new_n1145_), .Y(new_n1187_));
  AND2X1   g01123(.A(new_n1187_), .B(new_n1126_), .Y(new_n1188_));
  INVX1    g01124(.A(new_n1187_), .Y(new_n1189_));
  OR4X1    g01125(.A(new_n755_), .B(new_n843_), .C(new_n885_), .D(new_n301_), .Y(new_n1190_));
  OAI22X1  g01126(.A0(new_n161_), .A1(new_n88_), .B0(new_n106_), .B1(new_n72_), .Y(new_n1191_));
  OR4X1    g01127(.A(new_n1191_), .B(new_n516_), .C(new_n740_), .D(new_n227_), .Y(new_n1192_));
  OR2X1    g01128(.A(new_n1192_), .B(new_n1190_), .Y(new_n1193_));
  NOR4X1   g01129(.A(new_n286_), .B(new_n825_), .C(new_n303_), .D(new_n535_), .Y(new_n1194_));
  NOR3X1   g01130(.A(new_n217_), .B(new_n165_), .C(new_n648_), .Y(new_n1195_));
  NOR3X1   g01131(.A(new_n642_), .B(new_n197_), .C(new_n184_), .Y(new_n1196_));
  OAI21X1  g01132(.A0(new_n102_), .A1(new_n72_), .B0(new_n930_), .Y(new_n1197_));
  NOR3X1   g01133(.A(new_n1197_), .B(new_n596_), .C(new_n496_), .Y(new_n1198_));
  NAND4X1  g01134(.A(new_n1198_), .B(new_n1196_), .C(new_n1195_), .D(new_n1194_), .Y(new_n1199_));
  OAI22X1  g01135(.A0(new_n161_), .A1(new_n115_), .B0(new_n125_), .B1(new_n117_), .Y(new_n1200_));
  OR4X1    g01136(.A(new_n1200_), .B(new_n249_), .C(new_n138_), .D(new_n1008_), .Y(new_n1201_));
  OAI22X1  g01137(.A0(new_n127_), .A1(new_n123_), .B0(new_n94_), .B1(new_n69_), .Y(new_n1202_));
  OR4X1    g01138(.A(new_n1202_), .B(new_n391_), .C(new_n252_), .D(new_n357_), .Y(new_n1203_));
  OR4X1    g01139(.A(new_n1203_), .B(new_n1201_), .C(new_n1199_), .D(new_n1193_), .Y(new_n1204_));
  OAI22X1  g01140(.A0(new_n129_), .A1(new_n75_), .B0(new_n88_), .B1(new_n81_), .Y(new_n1205_));
  OR4X1    g01141(.A(new_n1205_), .B(new_n975_), .C(new_n86_), .D(new_n85_), .Y(new_n1206_));
  OR2X1    g01142(.A(new_n365_), .B(new_n271_), .Y(new_n1207_));
  NAND3X1  g01143(.A(new_n503_), .B(new_n281_), .C(new_n171_), .Y(new_n1208_));
  OR4X1    g01144(.A(new_n1208_), .B(new_n1207_), .C(new_n1206_), .D(new_n477_), .Y(new_n1209_));
  AOI21X1  g01145(.A0(new_n102_), .A1(new_n84_), .B0(new_n131_), .Y(new_n1210_));
  OAI22X1  g01146(.A0(new_n168_), .A1(new_n131_), .B0(new_n75_), .B1(new_n72_), .Y(new_n1211_));
  OR4X1    g01147(.A(new_n1211_), .B(new_n1210_), .C(new_n1158_), .D(new_n716_), .Y(new_n1212_));
  OR4X1    g01148(.A(new_n998_), .B(new_n260_), .C(new_n219_), .D(new_n651_), .Y(new_n1213_));
  OR4X1    g01149(.A(new_n1213_), .B(new_n432_), .C(new_n276_), .D(new_n449_), .Y(new_n1214_));
  AOI21X1  g01150(.A0(new_n129_), .A1(new_n125_), .B0(new_n84_), .Y(new_n1215_));
  OR2X1    g01151(.A(new_n1215_), .B(new_n523_), .Y(new_n1216_));
  OR4X1    g01152(.A(new_n1216_), .B(new_n1214_), .C(new_n1212_), .D(new_n1069_), .Y(new_n1217_));
  NOR2X1   g01153(.A(new_n1217_), .B(new_n1209_), .Y(new_n1218_));
  INVX1    g01154(.A(new_n1218_), .Y(new_n1219_));
  OAI22X1  g01155(.A0(new_n161_), .A1(new_n84_), .B0(new_n148_), .B1(new_n94_), .Y(new_n1220_));
  OAI22X1  g01156(.A0(new_n129_), .A1(new_n79_), .B0(new_n125_), .B1(new_n69_), .Y(new_n1221_));
  OR4X1    g01157(.A(new_n1221_), .B(new_n1220_), .C(new_n974_), .D(new_n137_), .Y(new_n1222_));
  AOI21X1  g01158(.A0(new_n143_), .A1(new_n81_), .B0(new_n168_), .Y(new_n1223_));
  OAI22X1  g01159(.A0(new_n119_), .A1(new_n99_), .B0(new_n92_), .B1(new_n88_), .Y(new_n1224_));
  OAI22X1  g01160(.A0(new_n182_), .A1(new_n115_), .B0(new_n148_), .B1(new_n143_), .Y(new_n1225_));
  OR2X1    g01161(.A(new_n1225_), .B(new_n1224_), .Y(new_n1226_));
  AOI21X1  g01162(.A0(new_n96_), .A1(new_n69_), .B0(new_n92_), .Y(new_n1227_));
  OR4X1    g01163(.A(new_n1227_), .B(new_n1006_), .C(new_n561_), .D(new_n440_), .Y(new_n1228_));
  OR4X1    g01164(.A(new_n1228_), .B(new_n1226_), .C(new_n1223_), .D(new_n1222_), .Y(new_n1229_));
  OR4X1    g01165(.A(new_n387_), .B(new_n245_), .C(new_n203_), .D(new_n124_), .Y(new_n1230_));
  OR4X1    g01166(.A(new_n1230_), .B(new_n546_), .C(new_n505_), .D(new_n420_), .Y(new_n1231_));
  NOR4X1   g01167(.A(new_n527_), .B(new_n506_), .C(new_n457_), .D(new_n757_), .Y(new_n1232_));
  INVX1    g01168(.A(new_n1232_), .Y(new_n1233_));
  OR4X1    g01169(.A(new_n627_), .B(new_n483_), .C(new_n455_), .D(new_n126_), .Y(new_n1234_));
  OR4X1    g01170(.A(new_n1234_), .B(new_n1233_), .C(new_n1231_), .D(new_n705_), .Y(new_n1235_));
  NOR4X1   g01171(.A(new_n1235_), .B(new_n1229_), .C(new_n1219_), .D(new_n1204_), .Y(new_n1236_));
  OR2X1    g01172(.A(new_n1236_), .B(new_n1189_), .Y(new_n1237_));
  OAI22X1  g01173(.A0(new_n168_), .A1(new_n99_), .B0(new_n106_), .B1(new_n92_), .Y(new_n1238_));
  NOR4X1   g01174(.A(new_n1238_), .B(new_n835_), .C(new_n184_), .D(new_n307_), .Y(new_n1239_));
  NOR4X1   g01175(.A(new_n586_), .B(new_n321_), .C(new_n474_), .D(new_n285_), .Y(new_n1240_));
  OR2X1    g01176(.A(new_n775_), .B(new_n522_), .Y(new_n1241_));
  NOR4X1   g01177(.A(new_n1241_), .B(new_n527_), .C(new_n540_), .D(new_n124_), .Y(new_n1242_));
  NAND4X1  g01178(.A(new_n1242_), .B(new_n1240_), .C(new_n1239_), .D(new_n763_), .Y(new_n1243_));
  OAI22X1  g01179(.A0(new_n131_), .A1(new_n84_), .B0(new_n81_), .B1(new_n75_), .Y(new_n1244_));
  OR2X1    g01180(.A(new_n1244_), .B(new_n814_), .Y(new_n1245_));
  OR4X1    g01181(.A(new_n615_), .B(new_n156_), .C(new_n149_), .D(new_n116_), .Y(new_n1246_));
  OR4X1    g01182(.A(new_n1246_), .B(new_n1245_), .C(new_n508_), .D(new_n154_), .Y(new_n1247_));
  NOR3X1   g01183(.A(new_n468_), .B(new_n247_), .C(new_n158_), .Y(new_n1248_));
  OAI22X1  g01184(.A0(new_n148_), .A1(new_n131_), .B0(new_n129_), .B1(new_n115_), .Y(new_n1249_));
  NOR3X1   g01185(.A(new_n1249_), .B(new_n355_), .C(new_n273_), .Y(new_n1250_));
  NOR4X1   g01186(.A(new_n998_), .B(new_n400_), .C(new_n147_), .D(new_n134_), .Y(new_n1251_));
  NAND3X1  g01187(.A(new_n1251_), .B(new_n1250_), .C(new_n1248_), .Y(new_n1252_));
  OAI22X1  g01188(.A0(new_n168_), .A1(new_n72_), .B0(new_n127_), .B1(new_n119_), .Y(new_n1253_));
  OR4X1    g01189(.A(new_n1253_), .B(new_n598_), .C(new_n197_), .D(new_n144_), .Y(new_n1254_));
  OAI22X1  g01190(.A0(new_n106_), .A1(new_n105_), .B0(new_n92_), .B1(new_n91_), .Y(new_n1255_));
  AOI21X1  g01191(.A0(new_n91_), .A1(new_n88_), .B0(new_n129_), .Y(new_n1256_));
  OR4X1    g01192(.A(new_n1256_), .B(new_n1255_), .C(new_n1254_), .D(new_n769_), .Y(new_n1257_));
  OR4X1    g01193(.A(new_n1257_), .B(new_n1252_), .C(new_n1247_), .D(new_n1243_), .Y(new_n1258_));
  OAI22X1  g01194(.A0(new_n105_), .A1(new_n84_), .B0(new_n102_), .B1(new_n94_), .Y(new_n1259_));
  OR4X1    g01195(.A(new_n603_), .B(new_n423_), .C(new_n681_), .D(new_n535_), .Y(new_n1260_));
  NOR2X1   g01196(.A(new_n168_), .B(new_n92_), .Y(new_n1261_));
  OR4X1    g01197(.A(new_n702_), .B(new_n422_), .C(new_n421_), .D(new_n111_), .Y(new_n1262_));
  OR4X1    g01198(.A(new_n1262_), .B(new_n723_), .C(new_n547_), .D(new_n1261_), .Y(new_n1263_));
  OR4X1    g01199(.A(new_n1263_), .B(new_n1260_), .C(new_n1259_), .D(new_n1258_), .Y(new_n1264_));
  OR4X1    g01200(.A(new_n412_), .B(new_n260_), .C(new_n256_), .D(new_n203_), .Y(new_n1265_));
  OR4X1    g01201(.A(new_n480_), .B(new_n226_), .C(new_n220_), .D(new_n114_), .Y(new_n1266_));
  OR4X1    g01202(.A(new_n740_), .B(new_n372_), .C(new_n812_), .D(new_n227_), .Y(new_n1267_));
  OR4X1    g01203(.A(new_n1267_), .B(new_n1266_), .C(new_n1265_), .D(new_n1116_), .Y(new_n1268_));
  OAI22X1  g01204(.A0(new_n182_), .A1(new_n69_), .B0(new_n148_), .B1(new_n90_), .Y(new_n1269_));
  OR4X1    g01205(.A(new_n1269_), .B(new_n391_), .C(new_n382_), .D(new_n265_), .Y(new_n1270_));
  AOI21X1  g01206(.A0(new_n105_), .A1(new_n78_), .B0(new_n79_), .Y(new_n1271_));
  OAI22X1  g01207(.A0(new_n148_), .A1(new_n72_), .B0(new_n123_), .B1(new_n92_), .Y(new_n1272_));
  OR4X1    g01208(.A(new_n1272_), .B(new_n1271_), .C(new_n286_), .D(new_n494_), .Y(new_n1273_));
  OAI22X1  g01209(.A0(new_n168_), .A1(new_n81_), .B0(new_n127_), .B1(new_n117_), .Y(new_n1274_));
  OAI22X1  g01210(.A0(new_n182_), .A1(new_n84_), .B0(new_n161_), .B1(new_n115_), .Y(new_n1275_));
  OAI22X1  g01211(.A0(new_n152_), .A1(new_n127_), .B0(new_n94_), .B1(new_n79_), .Y(new_n1276_));
  OAI22X1  g01212(.A0(new_n143_), .A1(new_n117_), .B0(new_n127_), .B1(new_n79_), .Y(new_n1277_));
  OR4X1    g01213(.A(new_n1277_), .B(new_n1276_), .C(new_n1275_), .D(new_n1274_), .Y(new_n1278_));
  NOR4X1   g01214(.A(new_n1278_), .B(new_n1273_), .C(new_n1270_), .D(new_n1268_), .Y(new_n1279_));
  INVX1    g01215(.A(new_n1279_), .Y(new_n1280_));
  NOR3X1   g01216(.A(new_n632_), .B(new_n968_), .C(new_n365_), .Y(new_n1281_));
  NOR3X1   g01217(.A(new_n261_), .B(new_n177_), .C(new_n1008_), .Y(new_n1282_));
  NAND3X1  g01218(.A(new_n1282_), .B(new_n1281_), .C(new_n1043_), .Y(new_n1283_));
  NOR2X1   g01219(.A(new_n72_), .B(new_n69_), .Y(new_n1284_));
  OR4X1    g01220(.A(new_n294_), .B(new_n159_), .C(new_n291_), .D(new_n1284_), .Y(new_n1285_));
  OR4X1    g01221(.A(new_n1285_), .B(new_n669_), .C(new_n478_), .D(new_n251_), .Y(new_n1286_));
  OR4X1    g01222(.A(new_n264_), .B(new_n224_), .C(new_n536_), .D(new_n162_), .Y(new_n1287_));
  OR4X1    g01223(.A(new_n1287_), .B(new_n594_), .C(new_n459_), .D(new_n843_), .Y(new_n1288_));
  OAI22X1  g01224(.A0(new_n117_), .A1(new_n94_), .B0(new_n106_), .B1(new_n90_), .Y(new_n1289_));
  OAI22X1  g01225(.A0(new_n127_), .A1(new_n96_), .B0(new_n91_), .B1(new_n72_), .Y(new_n1290_));
  OR4X1    g01226(.A(new_n1290_), .B(new_n1289_), .C(new_n187_), .D(new_n85_), .Y(new_n1291_));
  OR4X1    g01227(.A(new_n959_), .B(new_n766_), .C(new_n497_), .D(new_n475_), .Y(new_n1292_));
  OR4X1    g01228(.A(new_n1292_), .B(new_n1291_), .C(new_n1288_), .D(new_n1286_), .Y(new_n1293_));
  NOR4X1   g01229(.A(new_n1293_), .B(new_n1283_), .C(new_n1280_), .D(new_n1264_), .Y(new_n1294_));
  NOR2X1   g01230(.A(new_n1294_), .B(new_n1236_), .Y(new_n1295_));
  OAI22X1  g01231(.A0(new_n152_), .A1(new_n78_), .B0(new_n117_), .B1(new_n92_), .Y(new_n1296_));
  NOR4X1   g01232(.A(new_n1296_), .B(new_n1256_), .C(new_n673_), .D(new_n342_), .Y(new_n1297_));
  NOR3X1   g01233(.A(new_n938_), .B(new_n586_), .C(new_n615_), .Y(new_n1298_));
  NOR4X1   g01234(.A(new_n358_), .B(new_n292_), .C(new_n252_), .D(new_n381_), .Y(new_n1299_));
  NAND3X1  g01235(.A(new_n1299_), .B(new_n1298_), .C(new_n1297_), .Y(new_n1300_));
  OR4X1    g01236(.A(new_n741_), .B(new_n968_), .C(new_n319_), .D(new_n299_), .Y(new_n1301_));
  OR4X1    g01237(.A(new_n681_), .B(new_n239_), .C(new_n610_), .D(new_n338_), .Y(new_n1302_));
  OR4X1    g01238(.A(new_n1302_), .B(new_n1301_), .C(new_n744_), .D(new_n582_), .Y(new_n1303_));
  OR4X1    g01239(.A(new_n395_), .B(new_n385_), .C(new_n797_), .D(new_n261_), .Y(new_n1304_));
  OR4X1    g01240(.A(new_n1304_), .B(new_n887_), .C(new_n103_), .D(new_n100_), .Y(new_n1305_));
  AOI21X1  g01241(.A0(new_n92_), .A1(new_n90_), .B0(new_n79_), .Y(new_n1306_));
  OR4X1    g01242(.A(new_n1306_), .B(new_n1210_), .C(new_n474_), .D(new_n291_), .Y(new_n1307_));
  NOR4X1   g01243(.A(new_n1307_), .B(new_n1305_), .C(new_n1303_), .D(new_n1300_), .Y(new_n1308_));
  NOR2X1   g01244(.A(new_n616_), .B(new_n758_), .Y(new_n1309_));
  NAND2X1  g01245(.A(new_n1309_), .B(new_n1308_), .Y(new_n1310_));
  NOR4X1   g01246(.A(new_n510_), .B(new_n354_), .C(new_n400_), .D(new_n260_), .Y(new_n1311_));
  NOR4X1   g01247(.A(new_n494_), .B(new_n251_), .C(new_n194_), .D(new_n191_), .Y(new_n1312_));
  NAND3X1  g01248(.A(new_n1312_), .B(new_n1311_), .C(new_n140_), .Y(new_n1313_));
  AOI21X1  g01249(.A0(new_n108_), .A1(new_n81_), .B0(new_n117_), .Y(new_n1314_));
  OR4X1    g01250(.A(new_n1314_), .B(new_n158_), .C(new_n581_), .D(new_n126_), .Y(new_n1315_));
  AOI21X1  g01251(.A0(new_n168_), .A1(new_n88_), .B0(new_n108_), .Y(new_n1316_));
  OR4X1    g01252(.A(new_n1119_), .B(new_n618_), .C(new_n1316_), .D(new_n427_), .Y(new_n1317_));
  OR4X1    g01253(.A(new_n1317_), .B(new_n1315_), .C(new_n1313_), .D(new_n852_), .Y(new_n1318_));
  AOI21X1  g01254(.A0(new_n125_), .A1(new_n81_), .B0(new_n88_), .Y(new_n1319_));
  OAI22X1  g01255(.A0(new_n131_), .A1(new_n106_), .B0(new_n129_), .B1(new_n115_), .Y(new_n1320_));
  OAI22X1  g01256(.A0(new_n182_), .A1(new_n152_), .B0(new_n125_), .B1(new_n123_), .Y(new_n1321_));
  OR2X1    g01257(.A(new_n1321_), .B(new_n589_), .Y(new_n1322_));
  OR4X1    g01258(.A(new_n224_), .B(new_n201_), .C(new_n664_), .D(new_n426_), .Y(new_n1323_));
  OR4X1    g01259(.A(new_n1323_), .B(new_n1322_), .C(new_n1320_), .D(new_n1087_), .Y(new_n1324_));
  OR4X1    g01260(.A(new_n1324_), .B(new_n1319_), .C(new_n1289_), .D(new_n785_), .Y(new_n1325_));
  NOR4X1   g01261(.A(new_n768_), .B(new_n607_), .C(new_n1002_), .D(new_n498_), .Y(new_n1326_));
  NOR3X1   g01262(.A(new_n355_), .B(new_n282_), .C(new_n399_), .Y(new_n1327_));
  NOR4X1   g01263(.A(new_n422_), .B(new_n998_), .C(new_n812_), .D(new_n196_), .Y(new_n1328_));
  NAND3X1  g01264(.A(new_n1328_), .B(new_n1327_), .C(new_n1326_), .Y(new_n1329_));
  OR2X1    g01265(.A(new_n79_), .B(new_n78_), .Y(new_n1330_));
  NOR3X1   g01266(.A(new_n570_), .B(new_n365_), .C(new_n233_), .Y(new_n1331_));
  NAND4X1  g01267(.A(new_n1331_), .B(new_n719_), .C(new_n244_), .D(new_n1330_), .Y(new_n1332_));
  OAI22X1  g01268(.A0(new_n148_), .A1(new_n78_), .B0(new_n105_), .B1(new_n91_), .Y(new_n1333_));
  OAI21X1  g01269(.A0(new_n152_), .A1(new_n108_), .B0(new_n551_), .Y(new_n1334_));
  OR4X1    g01270(.A(new_n1334_), .B(new_n1333_), .C(new_n418_), .D(new_n651_), .Y(new_n1335_));
  OAI22X1  g01271(.A0(new_n182_), .A1(new_n168_), .B0(new_n91_), .B1(new_n72_), .Y(new_n1336_));
  OR4X1    g01272(.A(new_n1336_), .B(new_n1142_), .C(new_n361_), .D(new_n328_), .Y(new_n1337_));
  OR4X1    g01273(.A(new_n1337_), .B(new_n1335_), .C(new_n1332_), .D(new_n1329_), .Y(new_n1338_));
  NOR4X1   g01274(.A(new_n1338_), .B(new_n1325_), .C(new_n1318_), .D(new_n1310_), .Y(new_n1339_));
  OR2X1    g01275(.A(new_n1339_), .B(new_n1294_), .Y(new_n1340_));
  OR4X1    g01276(.A(new_n656_), .B(new_n740_), .C(new_n229_), .D(new_n180_), .Y(new_n1341_));
  OR4X1    g01277(.A(new_n497_), .B(new_n323_), .C(new_n806_), .D(new_n111_), .Y(new_n1342_));
  INVX1    g01278(.A(new_n574_), .Y(new_n1343_));
  NAND3X1  g01279(.A(new_n366_), .B(new_n341_), .C(new_n1343_), .Y(new_n1344_));
  OR4X1    g01280(.A(new_n1225_), .B(new_n1171_), .C(new_n664_), .D(new_n156_), .Y(new_n1345_));
  OR4X1    g01281(.A(new_n1345_), .B(new_n1344_), .C(new_n1342_), .D(new_n1341_), .Y(new_n1346_));
  OAI21X1  g01282(.A0(new_n90_), .A1(new_n84_), .B0(new_n364_), .Y(new_n1347_));
  OR4X1    g01283(.A(new_n1347_), .B(new_n1005_), .C(new_n938_), .D(new_n547_), .Y(new_n1348_));
  OR4X1    g01284(.A(new_n1348_), .B(new_n206_), .C(new_n757_), .D(new_n928_), .Y(new_n1349_));
  NOR3X1   g01285(.A(new_n723_), .B(new_n797_), .C(new_n1087_), .Y(new_n1350_));
  OR4X1    g01286(.A(new_n523_), .B(new_n998_), .C(new_n565_), .D(new_n191_), .Y(new_n1351_));
  OAI22X1  g01287(.A0(new_n125_), .A1(new_n79_), .B0(new_n119_), .B1(new_n108_), .Y(new_n1352_));
  OR2X1    g01288(.A(new_n1352_), .B(new_n702_), .Y(new_n1353_));
  NOR2X1   g01289(.A(new_n1353_), .B(new_n1351_), .Y(new_n1354_));
  NAND3X1  g01290(.A(new_n1354_), .B(new_n1350_), .C(new_n1248_), .Y(new_n1355_));
  NOR4X1   g01291(.A(new_n1355_), .B(new_n1349_), .C(new_n1346_), .D(new_n983_), .Y(new_n1356_));
  NAND3X1  g01292(.A(new_n1356_), .B(new_n1040_), .C(new_n859_), .Y(new_n1357_));
  INVX1    g01293(.A(new_n1357_), .Y(new_n1358_));
  NOR2X1   g01294(.A(new_n1358_), .B(new_n1339_), .Y(new_n1359_));
  OAI22X1  g01295(.A0(new_n182_), .A1(new_n88_), .B0(new_n115_), .B1(new_n99_), .Y(new_n1360_));
  OR4X1    g01296(.A(new_n489_), .B(new_n400_), .C(new_n256_), .D(new_n303_), .Y(new_n1361_));
  OR4X1    g01297(.A(new_n506_), .B(new_n496_), .C(new_n459_), .D(new_n118_), .Y(new_n1362_));
  OR4X1    g01298(.A(new_n493_), .B(new_n398_), .C(new_n457_), .D(new_n651_), .Y(new_n1363_));
  OR2X1    g01299(.A(new_n1173_), .B(new_n1135_), .Y(new_n1364_));
  NOR4X1   g01300(.A(new_n1364_), .B(new_n1363_), .C(new_n1362_), .D(new_n1361_), .Y(new_n1365_));
  OAI22X1  g01301(.A0(new_n88_), .A1(new_n72_), .B0(new_n81_), .B1(new_n75_), .Y(new_n1366_));
  OR2X1    g01302(.A(new_n1366_), .B(new_n612_), .Y(new_n1367_));
  NOR4X1   g01303(.A(new_n720_), .B(new_n475_), .C(new_n1087_), .D(new_n160_), .Y(new_n1368_));
  INVX1    g01304(.A(new_n1368_), .Y(new_n1369_));
  OAI21X1  g01305(.A0(new_n182_), .A1(new_n148_), .B0(new_n214_), .Y(new_n1370_));
  OR2X1    g01306(.A(new_n1370_), .B(new_n806_), .Y(new_n1371_));
  NOR3X1   g01307(.A(new_n1371_), .B(new_n1369_), .C(new_n1367_), .Y(new_n1372_));
  OR4X1    g01308(.A(new_n874_), .B(new_n566_), .C(new_n521_), .D(new_n337_), .Y(new_n1373_));
  OR4X1    g01309(.A(new_n540_), .B(new_n478_), .C(new_n187_), .D(new_n884_), .Y(new_n1374_));
  OR4X1    g01310(.A(new_n850_), .B(new_n449_), .C(new_n981_), .D(new_n1046_), .Y(new_n1375_));
  NOR3X1   g01311(.A(new_n1375_), .B(new_n1374_), .C(new_n1373_), .Y(new_n1376_));
  NAND3X1  g01312(.A(new_n1376_), .B(new_n1372_), .C(new_n1365_), .Y(new_n1377_));
  INVX1    g01313(.A(new_n331_), .Y(new_n1378_));
  NOR4X1   g01314(.A(new_n1227_), .B(new_n827_), .C(new_n638_), .D(new_n1316_), .Y(new_n1379_));
  NOR4X1   g01315(.A(new_n596_), .B(new_n543_), .C(new_n510_), .D(new_n740_), .Y(new_n1380_));
  NOR4X1   g01316(.A(new_n202_), .B(new_n381_), .C(new_n175_), .D(new_n162_), .Y(new_n1381_));
  NAND3X1  g01317(.A(new_n1381_), .B(new_n1380_), .C(new_n1379_), .Y(new_n1382_));
  OR4X1    g01318(.A(new_n1006_), .B(new_n354_), .C(new_n149_), .D(new_n80_), .Y(new_n1383_));
  OAI22X1  g01319(.A0(new_n125_), .A1(new_n75_), .B0(new_n117_), .B1(new_n99_), .Y(new_n1384_));
  OAI22X1  g01320(.A0(new_n161_), .A1(new_n75_), .B0(new_n143_), .B1(new_n69_), .Y(new_n1385_));
  OAI22X1  g01321(.A0(new_n152_), .A1(new_n81_), .B0(new_n143_), .B1(new_n115_), .Y(new_n1386_));
  OR4X1    g01322(.A(new_n1386_), .B(new_n1385_), .C(new_n1384_), .D(new_n1383_), .Y(new_n1387_));
  OR4X1    g01323(.A(new_n1387_), .B(new_n1382_), .C(new_n1378_), .D(new_n288_), .Y(new_n1388_));
  NOR4X1   g01324(.A(new_n1388_), .B(new_n1377_), .C(new_n1360_), .D(new_n438_), .Y(new_n1389_));
  OAI22X1  g01325(.A0(new_n123_), .A1(new_n78_), .B0(new_n96_), .B1(new_n90_), .Y(new_n1390_));
  OAI22X1  g01326(.A0(new_n117_), .A1(new_n92_), .B0(new_n105_), .B1(new_n91_), .Y(new_n1391_));
  OR4X1    g01327(.A(new_n1391_), .B(new_n778_), .C(new_n1390_), .D(new_n169_), .Y(new_n1392_));
  OAI22X1  g01328(.A0(new_n131_), .A1(new_n119_), .B0(new_n105_), .B1(new_n88_), .Y(new_n1393_));
  OR2X1    g01329(.A(new_n1393_), .B(new_n265_), .Y(new_n1394_));
  OR4X1    g01330(.A(new_n603_), .B(new_n286_), .C(new_n155_), .D(new_n133_), .Y(new_n1395_));
  OR4X1    g01331(.A(new_n1395_), .B(new_n1394_), .C(new_n1392_), .D(new_n1353_), .Y(new_n1396_));
  NOR4X1   g01332(.A(new_n292_), .B(new_n261_), .C(new_n180_), .D(new_n746_), .Y(new_n1397_));
  NOR2X1   g01333(.A(new_n92_), .B(new_n69_), .Y(new_n1398_));
  NOR4X1   g01334(.A(new_n596_), .B(new_n1398_), .C(new_n418_), .D(new_n615_), .Y(new_n1399_));
  NOR4X1   g01335(.A(new_n678_), .B(new_n627_), .C(new_n885_), .D(new_n162_), .Y(new_n1400_));
  NAND3X1  g01336(.A(new_n1400_), .B(new_n1399_), .C(new_n1397_), .Y(new_n1401_));
  OAI22X1  g01337(.A0(new_n182_), .A1(new_n123_), .B0(new_n102_), .B1(new_n81_), .Y(new_n1402_));
  OR4X1    g01338(.A(new_n1402_), .B(new_n815_), .C(new_n539_), .D(new_n229_), .Y(new_n1403_));
  OR4X1    g01339(.A(new_n714_), .B(new_n272_), .C(new_n379_), .D(new_n118_), .Y(new_n1404_));
  NOR3X1   g01340(.A(new_n454_), .B(new_n400_), .C(new_n209_), .Y(new_n1405_));
  INVX1    g01341(.A(new_n1405_), .Y(new_n1406_));
  AOI21X1  g01342(.A0(new_n106_), .A1(new_n96_), .B0(new_n72_), .Y(new_n1407_));
  AOI21X1  g01343(.A0(new_n92_), .A1(new_n90_), .B0(new_n84_), .Y(new_n1408_));
  OR4X1    g01344(.A(new_n1408_), .B(new_n1407_), .C(new_n1134_), .D(new_n233_), .Y(new_n1409_));
  OR4X1    g01345(.A(new_n1409_), .B(new_n1406_), .C(new_n1404_), .D(new_n1403_), .Y(new_n1410_));
  NOR3X1   g01346(.A(new_n1410_), .B(new_n1401_), .C(new_n1396_), .Y(new_n1411_));
  OR4X1    g01347(.A(new_n1261_), .B(new_n232_), .C(new_n223_), .D(new_n149_), .Y(new_n1412_));
  OR4X1    g01348(.A(new_n591_), .B(new_n1044_), .C(new_n358_), .D(new_n296_), .Y(new_n1413_));
  OAI22X1  g01349(.A0(new_n125_), .A1(new_n119_), .B0(new_n115_), .B1(new_n92_), .Y(new_n1414_));
  OAI22X1  g01350(.A0(new_n125_), .A1(new_n88_), .B0(new_n123_), .B1(new_n72_), .Y(new_n1415_));
  OAI22X1  g01351(.A0(new_n161_), .A1(new_n148_), .B0(new_n79_), .B1(new_n78_), .Y(new_n1416_));
  OAI22X1  g01352(.A0(new_n143_), .A1(new_n91_), .B0(new_n123_), .B1(new_n99_), .Y(new_n1417_));
  OR4X1    g01353(.A(new_n1417_), .B(new_n1416_), .C(new_n1415_), .D(new_n1238_), .Y(new_n1418_));
  OR4X1    g01354(.A(new_n395_), .B(new_n329_), .C(new_n137_), .D(new_n535_), .Y(new_n1419_));
  OR4X1    g01355(.A(new_n1419_), .B(new_n1418_), .C(new_n1414_), .D(new_n1018_), .Y(new_n1420_));
  OR4X1    g01356(.A(new_n1420_), .B(new_n1413_), .C(new_n1412_), .D(new_n1254_), .Y(new_n1421_));
  NOR3X1   g01357(.A(new_n1421_), .B(new_n1217_), .C(new_n1209_), .Y(new_n1422_));
  AND2X1   g01358(.A(new_n1422_), .B(new_n1411_), .Y(new_n1423_));
  NOR2X1   g01359(.A(new_n1423_), .B(new_n1389_), .Y(new_n1424_));
  OAI22X1  g01360(.A0(new_n123_), .A1(new_n90_), .B0(new_n117_), .B1(new_n105_), .Y(new_n1425_));
  OAI22X1  g01361(.A0(new_n148_), .A1(new_n99_), .B0(new_n91_), .B1(new_n78_), .Y(new_n1426_));
  OR2X1    g01362(.A(new_n206_), .B(new_n126_), .Y(new_n1427_));
  OR4X1    g01363(.A(new_n1427_), .B(new_n1426_), .C(new_n1425_), .D(new_n132_), .Y(new_n1428_));
  OR4X1    g01364(.A(new_n598_), .B(new_n294_), .C(new_n400_), .D(new_n142_), .Y(new_n1429_));
  OR4X1    g01365(.A(new_n1429_), .B(new_n395_), .C(new_n319_), .D(new_n806_), .Y(new_n1430_));
  OR4X1    g01366(.A(new_n1430_), .B(new_n1428_), .C(new_n222_), .D(new_n149_), .Y(new_n1431_));
  NOR4X1   g01367(.A(new_n468_), .B(new_n815_), .C(new_n393_), .D(new_n420_), .Y(new_n1432_));
  NOR4X1   g01368(.A(new_n387_), .B(new_n358_), .C(new_n178_), .D(new_n303_), .Y(new_n1433_));
  NOR4X1   g01369(.A(new_n276_), .B(new_n247_), .C(new_n449_), .D(new_n116_), .Y(new_n1434_));
  NAND3X1  g01370(.A(new_n1434_), .B(new_n1433_), .C(new_n1432_), .Y(new_n1435_));
  OAI22X1  g01371(.A0(new_n125_), .A1(new_n75_), .B0(new_n102_), .B1(new_n90_), .Y(new_n1436_));
  OR4X1    g01372(.A(new_n1436_), .B(new_n711_), .C(new_n589_), .D(new_n265_), .Y(new_n1437_));
  OAI22X1  g01373(.A0(new_n152_), .A1(new_n90_), .B0(new_n129_), .B1(new_n117_), .Y(new_n1438_));
  OR4X1    g01374(.A(new_n1438_), .B(new_n1407_), .C(new_n550_), .D(new_n441_), .Y(new_n1439_));
  OR4X1    g01375(.A(new_n1439_), .B(new_n1437_), .C(new_n1435_), .D(new_n1011_), .Y(new_n1440_));
  OR4X1    g01376(.A(new_n292_), .B(new_n226_), .C(new_n291_), .D(new_n379_), .Y(new_n1441_));
  OR4X1    g01377(.A(new_n1441_), .B(new_n547_), .C(new_n483_), .D(new_n286_), .Y(new_n1442_));
  AOI21X1  g01378(.A0(new_n92_), .A1(new_n81_), .B0(new_n115_), .Y(new_n1443_));
  OR4X1    g01379(.A(new_n951_), .B(new_n1443_), .C(new_n586_), .D(new_n494_), .Y(new_n1444_));
  OR4X1    g01380(.A(new_n361_), .B(new_n797_), .C(new_n234_), .D(new_n197_), .Y(new_n1445_));
  OR4X1    g01381(.A(new_n1445_), .B(new_n1444_), .C(new_n1316_), .D(new_n434_), .Y(new_n1446_));
  OAI22X1  g01382(.A0(new_n161_), .A1(new_n69_), .B0(new_n106_), .B1(new_n81_), .Y(new_n1447_));
  OR4X1    g01383(.A(new_n565_), .B(new_n814_), .C(new_n252_), .D(new_n85_), .Y(new_n1448_));
  OR4X1    g01384(.A(new_n1448_), .B(new_n755_), .C(new_n475_), .D(new_n323_), .Y(new_n1449_));
  OR4X1    g01385(.A(new_n1449_), .B(new_n1447_), .C(new_n701_), .D(new_n673_), .Y(new_n1450_));
  NAND3X1  g01386(.A(new_n820_), .B(new_n818_), .C(new_n817_), .Y(new_n1451_));
  OR4X1    g01387(.A(new_n273_), .B(new_n245_), .C(new_n240_), .D(new_n144_), .Y(new_n1452_));
  OR4X1    g01388(.A(new_n1452_), .B(new_n1320_), .C(new_n1451_), .D(new_n1087_), .Y(new_n1453_));
  OR4X1    g01389(.A(new_n1453_), .B(new_n1450_), .C(new_n1446_), .D(new_n1442_), .Y(new_n1454_));
  NOR4X1   g01390(.A(new_n421_), .B(new_n243_), .C(new_n208_), .D(new_n133_), .Y(new_n1455_));
  NOR3X1   g01391(.A(new_n418_), .B(new_n998_), .C(new_n156_), .Y(new_n1456_));
  OR4X1    g01392(.A(new_n1166_), .B(new_n408_), .C(new_n681_), .D(new_n301_), .Y(new_n1457_));
  OR4X1    g01393(.A(new_n256_), .B(new_n399_), .C(new_n229_), .D(new_n120_), .Y(new_n1458_));
  OAI22X1  g01394(.A0(new_n161_), .A1(new_n106_), .B0(new_n152_), .B1(new_n78_), .Y(new_n1459_));
  OR4X1    g01395(.A(new_n1459_), .B(new_n1415_), .C(new_n118_), .D(new_n86_), .Y(new_n1460_));
  OAI22X1  g01396(.A0(new_n152_), .A1(new_n99_), .B0(new_n127_), .B1(new_n96_), .Y(new_n1461_));
  OR4X1    g01397(.A(new_n1347_), .B(new_n931_), .C(new_n1461_), .D(new_n464_), .Y(new_n1462_));
  NOR4X1   g01398(.A(new_n1462_), .B(new_n1460_), .C(new_n1458_), .D(new_n1457_), .Y(new_n1463_));
  NAND4X1  g01399(.A(new_n1463_), .B(new_n1456_), .C(new_n1455_), .D(new_n1232_), .Y(new_n1464_));
  NOR4X1   g01400(.A(new_n1464_), .B(new_n1454_), .C(new_n1440_), .D(new_n1431_), .Y(new_n1465_));
  OR2X1    g01401(.A(new_n1465_), .B(new_n1423_), .Y(new_n1466_));
  OAI22X1  g01402(.A0(new_n161_), .A1(new_n117_), .B0(new_n96_), .B1(new_n72_), .Y(new_n1467_));
  INVX1    g01403(.A(new_n579_), .Y(new_n1468_));
  OR2X1    g01404(.A(new_n119_), .B(new_n105_), .Y(new_n1469_));
  NAND3X1  g01405(.A(new_n1469_), .B(new_n551_), .C(new_n1468_), .Y(new_n1470_));
  OR4X1    g01406(.A(new_n429_), .B(new_n431_), .C(new_n116_), .D(new_n1008_), .Y(new_n1471_));
  OR4X1    g01407(.A(new_n1471_), .B(new_n1470_), .C(new_n1094_), .D(new_n1467_), .Y(new_n1472_));
  OAI22X1  g01408(.A0(new_n161_), .A1(new_n115_), .B0(new_n143_), .B1(new_n106_), .Y(new_n1473_));
  OAI22X1  g01409(.A0(new_n148_), .A1(new_n90_), .B0(new_n115_), .B1(new_n78_), .Y(new_n1474_));
  OR4X1    g01410(.A(new_n1474_), .B(new_n1473_), .C(new_n1095_), .D(new_n1023_), .Y(new_n1475_));
  OR4X1    g01411(.A(new_n1475_), .B(new_n1472_), .C(new_n1344_), .D(new_n1342_), .Y(new_n1476_));
  NOR3X1   g01412(.A(new_n947_), .B(new_n772_), .C(new_n694_), .Y(new_n1477_));
  OAI22X1  g01413(.A0(new_n143_), .A1(new_n88_), .B0(new_n127_), .B1(new_n123_), .Y(new_n1478_));
  NOR3X1   g01414(.A(new_n1478_), .B(new_n441_), .C(new_n539_), .Y(new_n1479_));
  NOR3X1   g01415(.A(new_n1351_), .B(new_n432_), .C(new_n390_), .Y(new_n1480_));
  NAND3X1  g01416(.A(new_n1480_), .B(new_n1479_), .C(new_n1477_), .Y(new_n1481_));
  INVX1    g01417(.A(new_n692_), .Y(new_n1482_));
  OR4X1    g01418(.A(new_n1005_), .B(new_n570_), .C(new_n541_), .D(new_n217_), .Y(new_n1483_));
  OAI22X1  g01419(.A0(new_n182_), .A1(new_n123_), .B0(new_n117_), .B1(new_n108_), .Y(new_n1484_));
  OR2X1    g01420(.A(new_n1484_), .B(new_n142_), .Y(new_n1485_));
  OR4X1    g01421(.A(new_n1485_), .B(new_n561_), .C(new_n394_), .D(new_n86_), .Y(new_n1486_));
  OR4X1    g01422(.A(new_n1486_), .B(new_n1483_), .C(new_n1482_), .D(new_n635_), .Y(new_n1487_));
  NOR3X1   g01423(.A(new_n1487_), .B(new_n1481_), .C(new_n1476_), .Y(new_n1488_));
  AOI21X1  g01424(.A0(new_n1488_), .A1(new_n1086_), .B0(new_n1465_), .Y(new_n1489_));
  NAND2X1  g01425(.A(new_n1488_), .B(new_n1086_), .Y(new_n1490_));
  OR4X1    g01426(.A(new_n741_), .B(new_n546_), .C(new_n421_), .D(new_n282_), .Y(new_n1491_));
  OR4X1    g01427(.A(new_n792_), .B(new_n156_), .C(new_n155_), .D(new_n111_), .Y(new_n1492_));
  OAI22X1  g01428(.A0(new_n131_), .A1(new_n88_), .B0(new_n117_), .B1(new_n105_), .Y(new_n1493_));
  OR4X1    g01429(.A(new_n1493_), .B(new_n1492_), .C(new_n1491_), .D(new_n1427_), .Y(new_n1494_));
  OR4X1    g01430(.A(new_n1494_), .B(new_n929_), .C(new_n926_), .D(new_n797_), .Y(new_n1495_));
  OR4X1    g01431(.A(new_n446_), .B(new_n237_), .C(new_n233_), .D(new_n337_), .Y(new_n1496_));
  OAI22X1  g01432(.A0(new_n127_), .A1(new_n119_), .B0(new_n115_), .B1(new_n81_), .Y(new_n1497_));
  OR4X1    g01433(.A(new_n1497_), .B(new_n1496_), .C(new_n1371_), .D(new_n720_), .Y(new_n1498_));
  OAI22X1  g01434(.A0(new_n182_), .A1(new_n168_), .B0(new_n117_), .B1(new_n90_), .Y(new_n1499_));
  OR2X1    g01435(.A(new_n1499_), .B(new_n429_), .Y(new_n1500_));
  OR4X1    g01436(.A(new_n1500_), .B(new_n1287_), .C(new_n739_), .D(new_n384_), .Y(new_n1501_));
  OAI22X1  g01437(.A0(new_n152_), .A1(new_n127_), .B0(new_n143_), .B1(new_n123_), .Y(new_n1502_));
  NOR4X1   g01438(.A(new_n1502_), .B(new_n1090_), .C(new_n465_), .D(new_n169_), .Y(new_n1503_));
  NOR4X1   g01439(.A(new_n615_), .B(new_n273_), .C(new_n203_), .D(new_n191_), .Y(new_n1504_));
  NOR4X1   g01440(.A(new_n234_), .B(new_n218_), .C(new_n651_), .D(new_n86_), .Y(new_n1505_));
  NAND3X1  g01441(.A(new_n1505_), .B(new_n1504_), .C(new_n1503_), .Y(new_n1506_));
  NOR4X1   g01442(.A(new_n1506_), .B(new_n1501_), .C(new_n1498_), .D(new_n1495_), .Y(new_n1507_));
  OR4X1    g01443(.A(new_n700_), .B(new_n691_), .C(new_n493_), .D(new_n142_), .Y(new_n1508_));
  OR4X1    g01444(.A(new_n921_), .B(new_n1044_), .C(new_n757_), .D(new_n648_), .Y(new_n1509_));
  OR4X1    g01445(.A(new_n642_), .B(new_n523_), .C(new_n968_), .D(new_n410_), .Y(new_n1510_));
  NOR4X1   g01446(.A(new_n1510_), .B(new_n1509_), .C(new_n1508_), .D(new_n587_), .Y(new_n1511_));
  NOR2X1   g01447(.A(new_n702_), .B(new_n114_), .Y(new_n1512_));
  NAND2X1  g01448(.A(new_n1512_), .B(new_n1511_), .Y(new_n1513_));
  OAI22X1  g01449(.A0(new_n117_), .A1(new_n92_), .B0(new_n84_), .B1(new_n81_), .Y(new_n1514_));
  OAI22X1  g01450(.A0(new_n148_), .A1(new_n129_), .B0(new_n88_), .B1(new_n78_), .Y(new_n1515_));
  OAI22X1  g01451(.A0(new_n148_), .A1(new_n99_), .B0(new_n129_), .B1(new_n84_), .Y(new_n1516_));
  OAI22X1  g01452(.A0(new_n106_), .A1(new_n81_), .B0(new_n115_), .B1(new_n99_), .Y(new_n1517_));
  OR4X1    g01453(.A(new_n1517_), .B(new_n1473_), .C(new_n1516_), .D(new_n311_), .Y(new_n1518_));
  OR4X1    g01454(.A(new_n1518_), .B(new_n504_), .C(new_n497_), .D(new_n356_), .Y(new_n1519_));
  OR4X1    g01455(.A(new_n1519_), .B(new_n1515_), .C(new_n1514_), .D(new_n1474_), .Y(new_n1520_));
  OR4X1    g01456(.A(new_n571_), .B(new_n451_), .C(new_n396_), .D(new_n323_), .Y(new_n1521_));
  OR4X1    g01457(.A(new_n755_), .B(new_n579_), .C(new_n422_), .D(new_n197_), .Y(new_n1522_));
  OR4X1    g01458(.A(new_n1522_), .B(new_n483_), .C(new_n261_), .D(new_n357_), .Y(new_n1523_));
  OAI22X1  g01459(.A0(new_n152_), .A1(new_n90_), .B0(new_n92_), .B1(new_n91_), .Y(new_n1524_));
  OR4X1    g01460(.A(new_n1524_), .B(new_n656_), .C(new_n342_), .D(new_n196_), .Y(new_n1525_));
  OR4X1    g01461(.A(new_n1525_), .B(new_n1523_), .C(new_n1521_), .D(new_n1013_), .Y(new_n1526_));
  OR4X1    g01462(.A(new_n1142_), .B(new_n714_), .C(new_n291_), .D(new_n80_), .Y(new_n1527_));
  OR4X1    g01463(.A(new_n1527_), .B(new_n505_), .C(new_n194_), .D(new_n193_), .Y(new_n1528_));
  OAI22X1  g01464(.A0(new_n168_), .A1(new_n81_), .B0(new_n117_), .B1(new_n99_), .Y(new_n1529_));
  OAI22X1  g01465(.A0(new_n131_), .A1(new_n84_), .B0(new_n102_), .B1(new_n78_), .Y(new_n1530_));
  OAI22X1  g01466(.A0(new_n161_), .A1(new_n123_), .B0(new_n115_), .B1(new_n94_), .Y(new_n1531_));
  OR4X1    g01467(.A(new_n1531_), .B(new_n1530_), .C(new_n1529_), .D(new_n799_), .Y(new_n1532_));
  OR4X1    g01468(.A(new_n1532_), .B(new_n361_), .C(new_n321_), .D(new_n304_), .Y(new_n1533_));
  OR2X1    g01469(.A(new_n1533_), .B(new_n1528_), .Y(new_n1534_));
  NOR4X1   g01470(.A(new_n1534_), .B(new_n1526_), .C(new_n1520_), .D(new_n1513_), .Y(new_n1535_));
  NAND2X1  g01471(.A(new_n1535_), .B(new_n1507_), .Y(new_n1536_));
  NAND2X1  g01472(.A(new_n1536_), .B(new_n1490_), .Y(new_n1537_));
  OAI22X1  g01473(.A0(new_n127_), .A1(new_n88_), .B0(new_n102_), .B1(new_n78_), .Y(new_n1538_));
  OR4X1    g01474(.A(new_n1538_), .B(new_n1276_), .C(new_n1220_), .D(new_n488_), .Y(new_n1539_));
  OAI22X1  g01475(.A0(new_n143_), .A1(new_n123_), .B0(new_n108_), .B1(new_n84_), .Y(new_n1540_));
  OR2X1    g01476(.A(new_n1540_), .B(new_n390_), .Y(new_n1541_));
  OR4X1    g01477(.A(new_n631_), .B(new_n355_), .C(new_n181_), .D(new_n1087_), .Y(new_n1542_));
  OR4X1    g01478(.A(new_n156_), .B(new_n981_), .C(new_n1008_), .D(new_n307_), .Y(new_n1543_));
  OR4X1    g01479(.A(new_n1543_), .B(new_n1542_), .C(new_n1541_), .D(new_n1539_), .Y(new_n1544_));
  NOR3X1   g01480(.A(new_n217_), .B(new_n178_), .C(new_n431_), .Y(new_n1545_));
  NOR4X1   g01481(.A(new_n1082_), .B(new_n304_), .C(new_n187_), .D(new_n180_), .Y(new_n1546_));
  OAI22X1  g01482(.A0(new_n168_), .A1(new_n90_), .B0(new_n96_), .B1(new_n92_), .Y(new_n1547_));
  NOR3X1   g01483(.A(new_n1547_), .B(new_n193_), .C(new_n159_), .Y(new_n1548_));
  NAND3X1  g01484(.A(new_n1548_), .B(new_n1546_), .C(new_n1545_), .Y(new_n1549_));
  OAI22X1  g01485(.A0(new_n119_), .A1(new_n99_), .B0(new_n81_), .B1(new_n79_), .Y(new_n1550_));
  OR4X1    g01486(.A(new_n1550_), .B(new_n1256_), .C(new_n823_), .D(new_n778_), .Y(new_n1551_));
  OR4X1    g01487(.A(new_n194_), .B(new_n176_), .C(new_n103_), .D(new_n100_), .Y(new_n1552_));
  OR4X1    g01488(.A(new_n264_), .B(new_n292_), .C(new_n227_), .D(new_n291_), .Y(new_n1553_));
  OR4X1    g01489(.A(new_n723_), .B(new_n541_), .C(new_n459_), .D(new_n474_), .Y(new_n1554_));
  OR4X1    g01490(.A(new_n1554_), .B(new_n1553_), .C(new_n1552_), .D(new_n502_), .Y(new_n1555_));
  NOR4X1   g01491(.A(new_n1555_), .B(new_n1551_), .C(new_n1549_), .D(new_n1544_), .Y(new_n1556_));
  OR4X1    g01492(.A(new_n1171_), .B(new_n396_), .C(new_n362_), .D(new_n361_), .Y(new_n1557_));
  OAI22X1  g01493(.A0(new_n182_), .A1(new_n84_), .B0(new_n152_), .B1(new_n72_), .Y(new_n1558_));
  NOR4X1   g01494(.A(new_n1558_), .B(new_n678_), .C(new_n479_), .D(new_n141_), .Y(new_n1559_));
  OAI22X1  g01495(.A0(new_n119_), .A1(new_n90_), .B0(new_n106_), .B1(new_n99_), .Y(new_n1560_));
  NOR4X1   g01496(.A(new_n1560_), .B(new_n743_), .C(new_n374_), .D(new_n615_), .Y(new_n1561_));
  NAND2X1  g01497(.A(new_n1561_), .B(new_n1559_), .Y(new_n1562_));
  OR2X1    g01498(.A(new_n1562_), .B(new_n1557_), .Y(new_n1563_));
  INVX1    g01499(.A(new_n385_), .Y(new_n1564_));
  NAND3X1  g01500(.A(new_n1564_), .B(new_n346_), .C(new_n341_), .Y(new_n1565_));
  OR4X1    g01501(.A(new_n681_), .B(new_n399_), .C(new_n245_), .D(new_n610_), .Y(new_n1566_));
  OR4X1    g01502(.A(new_n1566_), .B(new_n1565_), .C(new_n1485_), .D(new_n732_), .Y(new_n1567_));
  OR4X1    g01503(.A(new_n1426_), .B(new_n506_), .C(new_n434_), .D(new_n717_), .Y(new_n1568_));
  OR4X1    g01504(.A(new_n1568_), .B(new_n1567_), .C(new_n1563_), .D(new_n1143_), .Y(new_n1569_));
  OR2X1    g01505(.A(new_n161_), .B(new_n119_), .Y(new_n1570_));
  NAND3X1  g01506(.A(new_n930_), .B(new_n503_), .C(new_n1570_), .Y(new_n1571_));
  OR4X1    g01507(.A(new_n294_), .B(new_n260_), .C(new_n296_), .D(new_n203_), .Y(new_n1572_));
  OR4X1    g01508(.A(new_n1572_), .B(new_n1571_), .C(new_n218_), .D(new_n792_), .Y(new_n1573_));
  OAI22X1  g01509(.A0(new_n127_), .A1(new_n75_), .B0(new_n123_), .B1(new_n90_), .Y(new_n1574_));
  OR2X1    g01510(.A(new_n1574_), .B(new_n455_), .Y(new_n1575_));
  OAI22X1  g01511(.A0(new_n161_), .A1(new_n91_), .B0(new_n125_), .B1(new_n106_), .Y(new_n1576_));
  OR4X1    g01512(.A(new_n383_), .B(new_n247_), .C(new_n439_), .D(new_n133_), .Y(new_n1577_));
  OR4X1    g01513(.A(new_n1577_), .B(new_n1576_), .C(new_n1575_), .D(new_n197_), .Y(new_n1578_));
  NOR2X1   g01514(.A(new_n75_), .B(new_n72_), .Y(new_n1579_));
  OR4X1    g01515(.A(new_n1044_), .B(new_n251_), .C(new_n457_), .D(new_n116_), .Y(new_n1580_));
  OR4X1    g01516(.A(new_n1580_), .B(new_n579_), .C(new_n825_), .D(new_n1579_), .Y(new_n1581_));
  OR4X1    g01517(.A(new_n799_), .B(new_n653_), .C(new_n487_), .D(new_n785_), .Y(new_n1582_));
  OR4X1    g01518(.A(new_n1582_), .B(new_n1581_), .C(new_n1578_), .D(new_n1573_), .Y(new_n1583_));
  NOR2X1   g01519(.A(new_n1583_), .B(new_n1569_), .Y(new_n1584_));
  AOI22X1  g01520(.A0(new_n1584_), .A1(new_n1556_), .B0(new_n1535_), .B1(new_n1507_), .Y(new_n1585_));
  AND2X1   g01521(.A(new_n1584_), .B(new_n1556_), .Y(new_n1586_));
  OR4X1    g01522(.A(new_n293_), .B(new_n400_), .C(new_n199_), .D(new_n758_), .Y(new_n1587_));
  OAI21X1  g01523(.A0(new_n115_), .A1(new_n94_), .B0(new_n551_), .Y(new_n1588_));
  OR4X1    g01524(.A(new_n1588_), .B(new_n1021_), .C(new_n884_), .D(new_n307_), .Y(new_n1589_));
  OR2X1    g01525(.A(new_n1589_), .B(new_n1587_), .Y(new_n1590_));
  OR4X1    g01526(.A(new_n1398_), .B(new_n815_), .C(new_n391_), .D(new_n363_), .Y(new_n1591_));
  OAI22X1  g01527(.A0(new_n152_), .A1(new_n125_), .B0(new_n102_), .B1(new_n72_), .Y(new_n1592_));
  OR2X1    g01528(.A(new_n1592_), .B(new_n938_), .Y(new_n1593_));
  OR2X1    g01529(.A(new_n848_), .B(new_n432_), .Y(new_n1594_));
  OAI22X1  g01530(.A0(new_n88_), .A1(new_n81_), .B0(new_n84_), .B1(new_n78_), .Y(new_n1595_));
  OAI22X1  g01531(.A0(new_n143_), .A1(new_n119_), .B0(new_n90_), .B1(new_n75_), .Y(new_n1596_));
  OR4X1    g01532(.A(new_n1596_), .B(new_n1595_), .C(new_n678_), .D(new_n240_), .Y(new_n1597_));
  OR4X1    g01533(.A(new_n494_), .B(new_n398_), .C(new_n536_), .D(new_n183_), .Y(new_n1598_));
  OAI22X1  g01534(.A0(new_n131_), .A1(new_n102_), .B0(new_n127_), .B1(new_n79_), .Y(new_n1599_));
  AOI21X1  g01535(.A0(new_n125_), .A1(new_n105_), .B0(new_n115_), .Y(new_n1600_));
  OR4X1    g01536(.A(new_n1600_), .B(new_n1599_), .C(new_n1598_), .D(new_n1597_), .Y(new_n1601_));
  OR4X1    g01537(.A(new_n1601_), .B(new_n1594_), .C(new_n1593_), .D(new_n1591_), .Y(new_n1602_));
  OR2X1    g01538(.A(new_n1602_), .B(new_n1590_), .Y(new_n1603_));
  OR2X1    g01539(.A(new_n514_), .B(new_n521_), .Y(new_n1604_));
  OR4X1    g01540(.A(new_n968_), .B(new_n354_), .C(new_n615_), .D(new_n274_), .Y(new_n1605_));
  OR4X1    g01541(.A(new_n840_), .B(new_n177_), .C(new_n141_), .D(new_n133_), .Y(new_n1606_));
  OR4X1    g01542(.A(new_n1606_), .B(new_n907_), .C(new_n493_), .D(new_n449_), .Y(new_n1607_));
  AOI21X1  g01543(.A0(new_n161_), .A1(new_n72_), .B0(new_n84_), .Y(new_n1608_));
  OAI22X1  g01544(.A0(new_n99_), .A1(new_n84_), .B0(new_n96_), .B1(new_n94_), .Y(new_n1609_));
  OR4X1    g01545(.A(new_n1609_), .B(new_n1347_), .C(new_n1608_), .D(new_n1100_), .Y(new_n1610_));
  OR4X1    g01546(.A(new_n1610_), .B(new_n1607_), .C(new_n1605_), .D(new_n442_), .Y(new_n1611_));
  OR4X1    g01547(.A(new_n213_), .B(new_n648_), .C(new_n585_), .D(new_n86_), .Y(new_n1612_));
  OAI22X1  g01548(.A0(new_n108_), .A1(new_n75_), .B0(new_n105_), .B1(new_n102_), .Y(new_n1613_));
  OR2X1    g01549(.A(new_n1613_), .B(new_n154_), .Y(new_n1614_));
  OR4X1    g01550(.A(new_n506_), .B(new_n243_), .C(new_n522_), .D(new_n218_), .Y(new_n1615_));
  OR4X1    g01551(.A(new_n634_), .B(new_n370_), .C(new_n176_), .D(new_n303_), .Y(new_n1616_));
  OR4X1    g01552(.A(new_n1616_), .B(new_n1615_), .C(new_n1614_), .D(new_n1612_), .Y(new_n1617_));
  OR4X1    g01553(.A(new_n1256_), .B(new_n676_), .C(new_n641_), .D(new_n607_), .Y(new_n1618_));
  OR4X1    g01554(.A(new_n1618_), .B(new_n285_), .C(new_n189_), .D(new_n1579_), .Y(new_n1619_));
  OR4X1    g01555(.A(new_n1619_), .B(new_n1617_), .C(new_n1611_), .D(new_n1450_), .Y(new_n1620_));
  NOR4X1   g01556(.A(new_n1620_), .B(new_n1604_), .C(new_n1603_), .D(new_n1421_), .Y(new_n1621_));
  OR2X1    g01557(.A(new_n1621_), .B(new_n1586_), .Y(new_n1622_));
  OAI22X1  g01558(.A0(new_n127_), .A1(new_n123_), .B0(new_n81_), .B1(new_n79_), .Y(new_n1623_));
  OR4X1    g01559(.A(new_n1385_), .B(new_n1623_), .C(new_n786_), .D(new_n657_), .Y(new_n1624_));
  OAI22X1  g01560(.A0(new_n129_), .A1(new_n96_), .B0(new_n115_), .B1(new_n99_), .Y(new_n1625_));
  OR4X1    g01561(.A(new_n1625_), .B(new_n511_), .C(new_n451_), .D(new_n785_), .Y(new_n1626_));
  OR4X1    g01562(.A(new_n385_), .B(new_n372_), .C(new_n974_), .D(new_n118_), .Y(new_n1627_));
  OR4X1    g01563(.A(new_n323_), .B(new_n819_), .C(new_n208_), .D(new_n184_), .Y(new_n1628_));
  OR4X1    g01564(.A(new_n1628_), .B(new_n1627_), .C(new_n1626_), .D(new_n1624_), .Y(new_n1629_));
  NOR4X1   g01565(.A(new_n498_), .B(new_n475_), .C(new_n474_), .D(new_n86_), .Y(new_n1630_));
  OR4X1    g01566(.A(new_n642_), .B(new_n539_), .C(new_n410_), .D(new_n156_), .Y(new_n1631_));
  NOR4X1   g01567(.A(new_n1631_), .B(new_n1261_), .C(new_n394_), .D(new_n1579_), .Y(new_n1632_));
  OAI22X1  g01568(.A0(new_n182_), .A1(new_n123_), .B0(new_n119_), .B1(new_n94_), .Y(new_n1633_));
  OAI22X1  g01569(.A0(new_n152_), .A1(new_n129_), .B0(new_n108_), .B1(new_n115_), .Y(new_n1634_));
  OAI22X1  g01570(.A0(new_n127_), .A1(new_n106_), .B0(new_n125_), .B1(new_n84_), .Y(new_n1635_));
  NOR4X1   g01571(.A(new_n1635_), .B(new_n1634_), .C(new_n1633_), .D(new_n632_), .Y(new_n1636_));
  NAND3X1  g01572(.A(new_n1636_), .B(new_n1632_), .C(new_n1630_), .Y(new_n1637_));
  OAI21X1  g01573(.A0(new_n123_), .A1(new_n99_), .B0(new_n776_), .Y(new_n1638_));
  AOI21X1  g01574(.A0(new_n92_), .A1(new_n90_), .B0(new_n123_), .Y(new_n1639_));
  OAI22X1  g01575(.A0(new_n125_), .A1(new_n88_), .B0(new_n108_), .B1(new_n106_), .Y(new_n1640_));
  OR4X1    g01576(.A(new_n1640_), .B(new_n1639_), .C(new_n1638_), .D(new_n714_), .Y(new_n1641_));
  OAI22X1  g01577(.A0(new_n152_), .A1(new_n78_), .B0(new_n96_), .B1(new_n90_), .Y(new_n1642_));
  OR4X1    g01578(.A(new_n354_), .B(new_n202_), .C(new_n196_), .D(new_n426_), .Y(new_n1643_));
  OR4X1    g01579(.A(new_n1643_), .B(new_n1642_), .C(new_n1641_), .D(new_n594_), .Y(new_n1644_));
  OR4X1    g01580(.A(new_n1644_), .B(new_n1637_), .C(new_n1629_), .D(new_n462_), .Y(new_n1645_));
  AOI21X1  g01581(.A0(new_n152_), .A1(new_n75_), .B0(new_n108_), .Y(new_n1646_));
  OAI22X1  g01582(.A0(new_n148_), .A1(new_n108_), .B0(new_n127_), .B1(new_n69_), .Y(new_n1647_));
  OR4X1    g01583(.A(new_n1647_), .B(new_n1646_), .C(new_n386_), .D(new_n535_), .Y(new_n1648_));
  OAI22X1  g01584(.A0(new_n105_), .A1(new_n75_), .B0(new_n84_), .B1(new_n72_), .Y(new_n1649_));
  OAI22X1  g01585(.A0(new_n152_), .A1(new_n94_), .B0(new_n125_), .B1(new_n96_), .Y(new_n1650_));
  OR4X1    g01586(.A(new_n1650_), .B(new_n875_), .C(new_n427_), .D(new_n1649_), .Y(new_n1651_));
  OR4X1    g01587(.A(new_n702_), .B(new_n393_), .C(new_n540_), .D(new_n615_), .Y(new_n1652_));
  OR4X1    g01588(.A(new_n1652_), .B(new_n417_), .C(new_n329_), .D(new_n299_), .Y(new_n1653_));
  OR4X1    g01589(.A(new_n1653_), .B(new_n1651_), .C(new_n1648_), .D(new_n794_), .Y(new_n1654_));
  NOR3X1   g01590(.A(new_n1654_), .B(new_n1645_), .C(new_n1603_), .Y(new_n1655_));
  NOR2X1   g01591(.A(new_n1655_), .B(new_n1621_), .Y(new_n1656_));
  OAI22X1  g01592(.A0(new_n131_), .A1(new_n115_), .B0(new_n129_), .B1(new_n106_), .Y(new_n1657_));
  OR4X1    g01593(.A(new_n1657_), .B(new_n1478_), .C(new_n578_), .D(new_n137_), .Y(new_n1658_));
  OR2X1    g01594(.A(new_n88_), .B(new_n78_), .Y(new_n1659_));
  NAND3X1  g01595(.A(new_n380_), .B(new_n818_), .C(new_n1659_), .Y(new_n1660_));
  OR4X1    g01596(.A(new_n998_), .B(new_n483_), .C(new_n474_), .D(new_n292_), .Y(new_n1661_));
  OR4X1    g01597(.A(new_n1661_), .B(new_n1660_), .C(new_n1658_), .D(new_n1594_), .Y(new_n1662_));
  OAI22X1  g01598(.A0(new_n168_), .A1(new_n99_), .B0(new_n125_), .B1(new_n117_), .Y(new_n1663_));
  OAI22X1  g01599(.A0(new_n152_), .A1(new_n125_), .B0(new_n131_), .B1(new_n88_), .Y(new_n1664_));
  NOR2X1   g01600(.A(new_n1664_), .B(new_n1663_), .Y(new_n1665_));
  NOR3X1   g01601(.A(new_n815_), .B(new_n386_), .C(new_n329_), .Y(new_n1666_));
  NOR3X1   g01602(.A(new_n647_), .B(new_n114_), .C(new_n80_), .Y(new_n1667_));
  NAND3X1  g01603(.A(new_n1667_), .B(new_n1666_), .C(new_n1665_), .Y(new_n1668_));
  OR4X1    g01604(.A(new_n1347_), .B(new_n1090_), .C(new_n814_), .D(new_n196_), .Y(new_n1669_));
  OR4X1    g01605(.A(new_n720_), .B(new_n679_), .C(new_n1166_), .D(new_n358_), .Y(new_n1670_));
  OR4X1    g01606(.A(new_n321_), .B(new_n265_), .C(new_n240_), .D(new_n239_), .Y(new_n1671_));
  OR4X1    g01607(.A(new_n1671_), .B(new_n1670_), .C(new_n1095_), .D(new_n874_), .Y(new_n1672_));
  OR4X1    g01608(.A(new_n1672_), .B(new_n1669_), .C(new_n1668_), .D(new_n1662_), .Y(new_n1673_));
  NOR4X1   g01609(.A(new_n1673_), .B(new_n966_), .C(new_n753_), .D(new_n736_), .Y(new_n1674_));
  OR2X1    g01610(.A(new_n1674_), .B(new_n1655_), .Y(new_n1675_));
  OR4X1    g01611(.A(new_n1673_), .B(new_n966_), .C(new_n753_), .D(new_n736_), .Y(new_n1676_));
  OR4X1    g01612(.A(new_n598_), .B(new_n691_), .C(new_n265_), .D(new_n177_), .Y(new_n1677_));
  OR2X1    g01613(.A(new_n835_), .B(new_n729_), .Y(new_n1678_));
  OR2X1    g01614(.A(new_n125_), .B(new_n91_), .Y(new_n1679_));
  OR2X1    g01615(.A(new_n91_), .B(new_n72_), .Y(new_n1680_));
  NAND3X1  g01616(.A(new_n1680_), .B(new_n1679_), .C(new_n1071_), .Y(new_n1681_));
  OR4X1    g01617(.A(new_n1681_), .B(new_n1678_), .C(new_n1677_), .D(new_n1207_), .Y(new_n1682_));
  OAI22X1  g01618(.A0(new_n168_), .A1(new_n92_), .B0(new_n108_), .B1(new_n79_), .Y(new_n1683_));
  OR4X1    g01619(.A(new_n1683_), .B(new_n523_), .C(new_n412_), .D(new_n329_), .Y(new_n1684_));
  OR4X1    g01620(.A(new_n1639_), .B(new_n1275_), .C(new_n480_), .D(new_n226_), .Y(new_n1685_));
  OR4X1    g01621(.A(new_n1685_), .B(new_n1684_), .C(new_n1682_), .D(new_n1123_), .Y(new_n1686_));
  NOR4X1   g01622(.A(new_n450_), .B(new_n815_), .C(new_n274_), .D(new_n399_), .Y(new_n1687_));
  NOR3X1   g01623(.A(new_n724_), .B(new_n596_), .C(new_n429_), .Y(new_n1688_));
  NOR4X1   g01624(.A(new_n1550_), .B(new_n579_), .C(new_n757_), .D(new_n183_), .Y(new_n1689_));
  NAND3X1  g01625(.A(new_n1689_), .B(new_n1688_), .C(new_n1687_), .Y(new_n1690_));
  NAND3X1  g01626(.A(new_n1469_), .B(new_n526_), .C(new_n366_), .Y(new_n1691_));
  OR4X1    g01627(.A(new_n603_), .B(new_n286_), .C(new_n280_), .D(new_n223_), .Y(new_n1692_));
  OR4X1    g01628(.A(new_n1692_), .B(new_n1691_), .C(new_n479_), .D(new_n219_), .Y(new_n1693_));
  OR4X1    g01629(.A(new_n263_), .B(new_n292_), .C(new_n208_), .D(new_n178_), .Y(new_n1694_));
  OAI22X1  g01630(.A0(new_n148_), .A1(new_n78_), .B0(new_n91_), .B1(new_n90_), .Y(new_n1695_));
  OR2X1    g01631(.A(new_n1695_), .B(new_n209_), .Y(new_n1696_));
  OR4X1    g01632(.A(new_n1082_), .B(new_n383_), .C(new_n356_), .D(new_n681_), .Y(new_n1697_));
  AOI21X1  g01633(.A0(new_n123_), .A1(new_n91_), .B0(new_n127_), .Y(new_n1698_));
  OR2X1    g01634(.A(new_n1698_), .B(new_n496_), .Y(new_n1699_));
  OR4X1    g01635(.A(new_n1699_), .B(new_n1697_), .C(new_n1696_), .D(new_n1694_), .Y(new_n1700_));
  OAI22X1  g01636(.A0(new_n168_), .A1(new_n99_), .B0(new_n123_), .B1(new_n105_), .Y(new_n1701_));
  OR4X1    g01637(.A(new_n1701_), .B(new_n589_), .C(new_n740_), .D(new_n304_), .Y(new_n1702_));
  AOI21X1  g01638(.A0(new_n161_), .A1(new_n94_), .B0(new_n79_), .Y(new_n1703_));
  OR4X1    g01639(.A(new_n1703_), .B(new_n714_), .C(new_n702_), .D(new_n176_), .Y(new_n1704_));
  OR4X1    g01640(.A(new_n1704_), .B(new_n1702_), .C(new_n1700_), .D(new_n1693_), .Y(new_n1705_));
  OR4X1    g01641(.A(new_n1705_), .B(new_n1690_), .C(new_n1686_), .D(new_n167_), .Y(new_n1706_));
  AND2X1   g01642(.A(new_n1706_), .B(new_n1676_), .Y(new_n1707_));
  NOR4X1   g01643(.A(new_n1705_), .B(new_n1690_), .C(new_n1686_), .D(new_n167_), .Y(new_n1708_));
  OR4X1    g01644(.A(new_n1609_), .B(new_n1438_), .C(new_n959_), .D(new_n209_), .Y(new_n1709_));
  OR2X1    g01645(.A(new_n143_), .B(new_n106_), .Y(new_n1710_));
  NAND3X1  g01646(.A(new_n244_), .B(new_n1710_), .C(new_n1330_), .Y(new_n1711_));
  OR4X1    g01647(.A(new_n243_), .B(new_n234_), .C(new_n648_), .D(new_n746_), .Y(new_n1712_));
  OR4X1    g01648(.A(new_n1712_), .B(new_n1711_), .C(new_n1089_), .D(new_n347_), .Y(new_n1713_));
  OR4X1    g01649(.A(new_n586_), .B(new_n444_), .C(new_n385_), .D(new_n981_), .Y(new_n1714_));
  OR4X1    g01650(.A(new_n1714_), .B(new_n506_), .C(new_n301_), .D(new_n196_), .Y(new_n1715_));
  OR4X1    g01651(.A(new_n1715_), .B(new_n1713_), .C(new_n1709_), .D(new_n1573_), .Y(new_n1716_));
  OAI22X1  g01652(.A0(new_n125_), .A1(new_n96_), .B0(new_n102_), .B1(new_n92_), .Y(new_n1717_));
  OR4X1    g01653(.A(new_n1717_), .B(new_n823_), .C(new_n272_), .D(new_n237_), .Y(new_n1718_));
  AOI21X1  g01654(.A0(new_n161_), .A1(new_n108_), .B0(new_n117_), .Y(new_n1719_));
  AOI21X1  g01655(.A0(new_n99_), .A1(new_n72_), .B0(new_n117_), .Y(new_n1720_));
  OR4X1    g01656(.A(new_n1720_), .B(new_n1719_), .C(new_n370_), .D(new_n273_), .Y(new_n1721_));
  OR4X1    g01657(.A(new_n371_), .B(new_n578_), .C(new_n233_), .D(new_n170_), .Y(new_n1722_));
  OR4X1    g01658(.A(new_n1722_), .B(new_n1721_), .C(new_n1718_), .D(new_n1557_), .Y(new_n1723_));
  OAI22X1  g01659(.A0(new_n127_), .A1(new_n84_), .B0(new_n105_), .B1(new_n91_), .Y(new_n1724_));
  OAI22X1  g01660(.A0(new_n127_), .A1(new_n117_), .B0(new_n96_), .B1(new_n90_), .Y(new_n1725_));
  NOR4X1   g01661(.A(new_n1725_), .B(new_n1724_), .C(new_n1640_), .D(new_n1220_), .Y(new_n1726_));
  NOR4X1   g01662(.A(new_n840_), .B(new_n843_), .C(new_n299_), .D(new_n259_), .Y(new_n1727_));
  NOR4X1   g01663(.A(new_n194_), .B(new_n175_), .C(new_n449_), .D(new_n337_), .Y(new_n1728_));
  NAND3X1  g01664(.A(new_n1728_), .B(new_n1727_), .C(new_n1726_), .Y(new_n1729_));
  OR2X1    g01665(.A(new_n127_), .B(new_n69_), .Y(new_n1730_));
  NAND3X1  g01666(.A(new_n719_), .B(new_n1730_), .C(new_n171_), .Y(new_n1731_));
  OR4X1    g01667(.A(new_n328_), .B(new_n261_), .C(new_n291_), .D(new_n884_), .Y(new_n1732_));
  OR4X1    g01668(.A(new_n968_), .B(new_n850_), .C(new_n758_), .D(new_n137_), .Y(new_n1733_));
  OR4X1    g01669(.A(new_n1733_), .B(new_n1732_), .C(new_n1731_), .D(new_n1729_), .Y(new_n1734_));
  NOR4X1   g01670(.A(new_n1734_), .B(new_n1723_), .C(new_n1716_), .D(new_n1686_), .Y(new_n1735_));
  OR4X1    g01671(.A(new_n1271_), .B(new_n293_), .C(new_n282_), .D(new_n256_), .Y(new_n1736_));
  OR4X1    g01672(.A(new_n1736_), .B(new_n594_), .C(new_n627_), .D(new_n263_), .Y(new_n1737_));
  OR4X1    g01673(.A(new_n724_), .B(new_n543_), .C(new_n598_), .D(new_n286_), .Y(new_n1738_));
  OR2X1    g01674(.A(new_n143_), .B(new_n119_), .Y(new_n1739_));
  NAND3X1  g01675(.A(new_n1056_), .B(new_n1739_), .C(new_n326_), .Y(new_n1740_));
  OR2X1    g01676(.A(new_n102_), .B(new_n90_), .Y(new_n1741_));
  OR2X1    g01677(.A(new_n182_), .B(new_n123_), .Y(new_n1742_));
  NAND3X1  g01678(.A(new_n558_), .B(new_n1742_), .C(new_n1741_), .Y(new_n1743_));
  OR4X1    g01679(.A(new_n1743_), .B(new_n1740_), .C(new_n1738_), .D(new_n419_), .Y(new_n1744_));
  OR4X1    g01680(.A(new_n292_), .B(new_n259_), .C(new_n246_), .D(new_n199_), .Y(new_n1745_));
  OR4X1    g01681(.A(new_n1745_), .B(new_n642_), .C(new_n500_), .D(new_n396_), .Y(new_n1746_));
  OR4X1    g01682(.A(new_n659_), .B(new_n1316_), .C(new_n885_), .D(new_n183_), .Y(new_n1747_));
  OR4X1    g01683(.A(new_n1747_), .B(new_n1746_), .C(new_n1744_), .D(new_n1737_), .Y(new_n1748_));
  OAI22X1  g01684(.A0(new_n161_), .A1(new_n69_), .B0(new_n148_), .B1(new_n108_), .Y(new_n1749_));
  OR4X1    g01685(.A(new_n1749_), .B(new_n234_), .C(new_n449_), .D(new_n337_), .Y(new_n1750_));
  AOI21X1  g01686(.A0(new_n108_), .A1(new_n94_), .B0(new_n106_), .Y(new_n1751_));
  OAI22X1  g01687(.A0(new_n182_), .A1(new_n96_), .B0(new_n108_), .B1(new_n102_), .Y(new_n1752_));
  OR4X1    g01688(.A(new_n1752_), .B(new_n1751_), .C(new_n1701_), .D(new_n1657_), .Y(new_n1753_));
  OR4X1    g01689(.A(new_n1753_), .B(new_n285_), .C(new_n189_), .D(new_n1579_), .Y(new_n1754_));
  OR4X1    g01690(.A(new_n243_), .B(new_n133_), .C(new_n126_), .D(new_n1284_), .Y(new_n1755_));
  AOI21X1  g01691(.A0(new_n182_), .A1(new_n78_), .B0(new_n117_), .Y(new_n1756_));
  AOI21X1  g01692(.A0(new_n129_), .A1(new_n81_), .B0(new_n119_), .Y(new_n1757_));
  OR2X1    g01693(.A(new_n1757_), .B(new_n1756_), .Y(new_n1758_));
  OR4X1    g01694(.A(new_n387_), .B(new_n274_), .C(new_n261_), .D(new_n159_), .Y(new_n1759_));
  OR4X1    g01695(.A(new_n723_), .B(new_n329_), .C(new_n323_), .D(new_n138_), .Y(new_n1760_));
  OR4X1    g01696(.A(new_n1760_), .B(new_n1759_), .C(new_n1758_), .D(new_n1755_), .Y(new_n1761_));
  OR4X1    g01697(.A(new_n1082_), .B(new_n219_), .C(new_n200_), .D(new_n124_), .Y(new_n1762_));
  OR2X1    g01698(.A(new_n993_), .B(new_n569_), .Y(new_n1763_));
  OR2X1    g01699(.A(new_n582_), .B(new_n843_), .Y(new_n1764_));
  OR4X1    g01700(.A(new_n586_), .B(new_n612_), .C(new_n460_), .D(new_n394_), .Y(new_n1765_));
  OR4X1    g01701(.A(new_n1765_), .B(new_n1764_), .C(new_n1763_), .D(new_n1762_), .Y(new_n1766_));
  OR4X1    g01702(.A(new_n1766_), .B(new_n1761_), .C(new_n1754_), .D(new_n1750_), .Y(new_n1767_));
  AOI21X1  g01703(.A0(new_n106_), .A1(new_n88_), .B0(new_n131_), .Y(new_n1768_));
  NOR4X1   g01704(.A(new_n1135_), .B(new_n1768_), .C(new_n629_), .D(new_n165_), .Y(new_n1769_));
  NOR3X1   g01705(.A(new_n815_), .B(new_n393_), .C(new_n574_), .Y(new_n1770_));
  NOR4X1   g01706(.A(new_n208_), .B(new_n180_), .C(new_n746_), .D(new_n142_), .Y(new_n1771_));
  NAND3X1  g01707(.A(new_n1771_), .B(new_n1770_), .C(new_n1769_), .Y(new_n1772_));
  OR4X1    g01708(.A(new_n1205_), .B(new_n1002_), .C(new_n560_), .D(new_n333_), .Y(new_n1773_));
  NOR3X1   g01709(.A(new_n1473_), .B(new_n496_), .C(new_n294_), .Y(new_n1774_));
  INVX1    g01710(.A(new_n1774_), .Y(new_n1775_));
  OR4X1    g01711(.A(new_n1398_), .B(new_n421_), .C(new_n455_), .D(new_n494_), .Y(new_n1776_));
  OR2X1    g01712(.A(new_n400_), .B(new_n202_), .Y(new_n1777_));
  OAI22X1  g01713(.A0(new_n161_), .A1(new_n79_), .B0(new_n129_), .B1(new_n88_), .Y(new_n1778_));
  AOI21X1  g01714(.A0(new_n148_), .A1(new_n79_), .B0(new_n72_), .Y(new_n1779_));
  OAI22X1  g01715(.A0(new_n127_), .A1(new_n84_), .B0(new_n123_), .B1(new_n94_), .Y(new_n1780_));
  OR4X1    g01716(.A(new_n1780_), .B(new_n1384_), .C(new_n1296_), .D(new_n1259_), .Y(new_n1781_));
  OR4X1    g01717(.A(new_n1781_), .B(new_n1779_), .C(new_n1778_), .D(new_n1777_), .Y(new_n1782_));
  OR4X1    g01718(.A(new_n1782_), .B(new_n1776_), .C(new_n1775_), .D(new_n1773_), .Y(new_n1783_));
  NOR4X1   g01719(.A(new_n1783_), .B(new_n1772_), .C(new_n1767_), .D(new_n1748_), .Y(new_n1784_));
  AOI21X1  g01720(.A0(new_n1784_), .A1(new_n1708_), .B0(new_n1735_), .Y(new_n1785_));
  XOR2X1   g01721(.A(new_n1706_), .B(new_n1676_), .Y(new_n1786_));
  AOI21X1  g01722(.A0(new_n1786_), .A1(new_n1785_), .B0(new_n1707_), .Y(new_n1787_));
  XOR2X1   g01723(.A(new_n1676_), .B(new_n1655_), .Y(new_n1788_));
  OAI21X1  g01724(.A0(new_n1788_), .A1(new_n1787_), .B0(new_n1675_), .Y(new_n1789_));
  XOR2X1   g01725(.A(new_n1655_), .B(new_n1621_), .Y(new_n1790_));
  AOI21X1  g01726(.A0(new_n1790_), .A1(new_n1789_), .B0(new_n1656_), .Y(new_n1791_));
  XOR2X1   g01727(.A(new_n1621_), .B(new_n1586_), .Y(new_n1792_));
  INVX1    g01728(.A(new_n1792_), .Y(new_n1793_));
  OAI21X1  g01729(.A0(new_n1793_), .A1(new_n1791_), .B0(new_n1622_), .Y(new_n1794_));
  INVX1    g01730(.A(new_n1536_), .Y(new_n1795_));
  XOR2X1   g01731(.A(new_n1586_), .B(new_n1795_), .Y(new_n1796_));
  AOI21X1  g01732(.A0(new_n1796_), .A1(new_n1794_), .B0(new_n1585_), .Y(new_n1797_));
  NOR2X1   g01733(.A(new_n1536_), .B(new_n1490_), .Y(new_n1798_));
  OAI21X1  g01734(.A0(new_n1798_), .A1(new_n1797_), .B0(new_n1537_), .Y(new_n1799_));
  INVX1    g01735(.A(new_n1465_), .Y(new_n1800_));
  XOR2X1   g01736(.A(new_n1490_), .B(new_n1800_), .Y(new_n1801_));
  AND2X1   g01737(.A(new_n1801_), .B(new_n1799_), .Y(new_n1802_));
  XOR2X1   g01738(.A(new_n1465_), .B(new_n1423_), .Y(new_n1803_));
  OAI21X1  g01739(.A0(new_n1802_), .A1(new_n1489_), .B0(new_n1803_), .Y(new_n1804_));
  NAND2X1  g01740(.A(new_n1804_), .B(new_n1466_), .Y(new_n1805_));
  XOR2X1   g01741(.A(new_n1423_), .B(new_n1389_), .Y(new_n1806_));
  AND2X1   g01742(.A(new_n1806_), .B(new_n1805_), .Y(new_n1807_));
  XOR2X1   g01743(.A(new_n1389_), .B(new_n1358_), .Y(new_n1808_));
  OAI21X1  g01744(.A0(new_n1807_), .A1(new_n1424_), .B0(new_n1808_), .Y(new_n1809_));
  OAI21X1  g01745(.A0(new_n1389_), .A1(new_n1358_), .B0(new_n1809_), .Y(new_n1810_));
  XOR2X1   g01746(.A(new_n1358_), .B(new_n1339_), .Y(new_n1811_));
  AOI21X1  g01747(.A0(new_n1811_), .A1(new_n1810_), .B0(new_n1359_), .Y(new_n1812_));
  AND2X1   g01748(.A(new_n1339_), .B(new_n1294_), .Y(new_n1813_));
  OAI21X1  g01749(.A0(new_n1813_), .A1(new_n1812_), .B0(new_n1340_), .Y(new_n1814_));
  XOR2X1   g01750(.A(new_n1294_), .B(new_n1236_), .Y(new_n1815_));
  AND2X1   g01751(.A(new_n1815_), .B(new_n1814_), .Y(new_n1816_));
  XOR2X1   g01752(.A(new_n1236_), .B(new_n1189_), .Y(new_n1817_));
  OAI21X1  g01753(.A0(new_n1816_), .A1(new_n1295_), .B0(new_n1817_), .Y(new_n1818_));
  NAND2X1  g01754(.A(new_n1818_), .B(new_n1237_), .Y(new_n1819_));
  XOR2X1   g01755(.A(new_n1187_), .B(new_n1126_), .Y(new_n1820_));
  AND2X1   g01756(.A(new_n1820_), .B(new_n1819_), .Y(new_n1821_));
  INVX1    g01757(.A(new_n1065_), .Y(new_n1822_));
  XOR2X1   g01758(.A(new_n1126_), .B(new_n1822_), .Y(new_n1823_));
  OAI21X1  g01759(.A0(new_n1821_), .A1(new_n1188_), .B0(new_n1823_), .Y(new_n1824_));
  OAI21X1  g01760(.A0(new_n1127_), .A1(new_n1065_), .B0(new_n1824_), .Y(new_n1825_));
  XOR2X1   g01761(.A(new_n1065_), .B(new_n985_), .Y(new_n1826_));
  AOI21X1  g01762(.A0(new_n1826_), .A1(new_n1825_), .B0(new_n1066_), .Y(new_n1827_));
  AND2X1   g01763(.A(new_n985_), .B(new_n957_), .Y(new_n1828_));
  OAI21X1  g01764(.A0(new_n1828_), .A1(new_n1827_), .B0(new_n986_), .Y(new_n1829_));
  XOR2X1   g01765(.A(new_n957_), .B(new_n903_), .Y(new_n1830_));
  AND2X1   g01766(.A(new_n1830_), .B(new_n1829_), .Y(new_n1831_));
  XOR2X1   g01767(.A(new_n903_), .B(new_n847_), .Y(new_n1832_));
  OAI21X1  g01768(.A0(new_n1831_), .A1(new_n956_), .B0(new_n1832_), .Y(new_n1833_));
  NAND2X1  g01769(.A(new_n1833_), .B(new_n902_), .Y(new_n1834_));
  XOR2X1   g01770(.A(new_n847_), .B(new_n783_), .Y(new_n1835_));
  NAND2X1  g01771(.A(new_n1835_), .B(new_n1834_), .Y(new_n1836_));
  OAI21X1  g01772(.A0(new_n847_), .A1(new_n783_), .B0(new_n1836_), .Y(new_n1837_));
  XOR2X1   g01773(.A(new_n783_), .B(new_n690_), .Y(new_n1838_));
  AOI21X1  g01774(.A0(new_n1838_), .A1(new_n1837_), .B0(new_n784_), .Y(new_n1839_));
  XOR2X1   g01775(.A(new_n690_), .B(new_n623_), .Y(new_n1840_));
  INVX1    g01776(.A(new_n1840_), .Y(new_n1841_));
  OR2X1    g01777(.A(new_n1841_), .B(new_n1839_), .Y(new_n1842_));
  OAI21X1  g01778(.A0(new_n690_), .A1(new_n623_), .B0(new_n1842_), .Y(new_n1843_));
  XOR2X1   g01779(.A(new_n623_), .B(new_n520_), .Y(new_n1844_));
  AOI21X1  g01780(.A0(new_n1844_), .A1(new_n1843_), .B0(new_n624_), .Y(new_n1845_));
  OR4X1    g01781(.A(new_n634_), .B(new_n371_), .C(new_n678_), .D(new_n286_), .Y(new_n1846_));
  OR4X1    g01782(.A(new_n539_), .B(new_n398_), .C(new_n664_), .D(new_n156_), .Y(new_n1847_));
  OR4X1    g01783(.A(new_n497_), .B(new_n475_), .C(new_n304_), .D(new_n86_), .Y(new_n1848_));
  OR4X1    g01784(.A(new_n1848_), .B(new_n1847_), .C(new_n1846_), .D(new_n738_), .Y(new_n1849_));
  OAI22X1  g01785(.A0(new_n161_), .A1(new_n148_), .B0(new_n117_), .B1(new_n72_), .Y(new_n1850_));
  OR4X1    g01786(.A(new_n1752_), .B(new_n1850_), .C(new_n541_), .D(new_n350_), .Y(new_n1851_));
  OR4X1    g01787(.A(new_n1415_), .B(new_n1386_), .C(new_n483_), .D(new_n280_), .Y(new_n1852_));
  OR4X1    g01788(.A(new_n1106_), .B(new_n1002_), .C(new_n514_), .D(new_n311_), .Y(new_n1853_));
  OR4X1    g01789(.A(new_n1853_), .B(new_n1852_), .C(new_n1851_), .D(new_n1849_), .Y(new_n1854_));
  INVX1    g01790(.A(new_n132_), .Y(new_n1855_));
  NOR4X1   g01791(.A(new_n256_), .B(new_n578_), .C(new_n252_), .D(new_n208_), .Y(new_n1856_));
  NOR4X1   g01792(.A(new_n1261_), .B(new_n393_), .C(new_n181_), .D(new_n535_), .Y(new_n1857_));
  NOR4X1   g01793(.A(new_n642_), .B(new_n361_), .C(new_n819_), .D(new_n240_), .Y(new_n1858_));
  NAND4X1  g01794(.A(new_n1858_), .B(new_n1857_), .C(new_n1856_), .D(new_n1855_), .Y(new_n1859_));
  NOR4X1   g01795(.A(new_n724_), .B(new_n496_), .C(new_n459_), .D(new_n261_), .Y(new_n1860_));
  NOR4X1   g01796(.A(new_n758_), .B(new_n825_), .C(new_n139_), .D(new_n884_), .Y(new_n1861_));
  NAND2X1  g01797(.A(new_n1861_), .B(new_n1860_), .Y(new_n1862_));
  OR4X1    g01798(.A(new_n1172_), .B(new_n423_), .C(new_n206_), .D(new_n124_), .Y(new_n1863_));
  OR4X1    g01799(.A(new_n494_), .B(new_n228_), .C(new_n1579_), .D(new_n1284_), .Y(new_n1864_));
  OR4X1    g01800(.A(new_n1864_), .B(new_n1863_), .C(new_n1119_), .D(new_n875_), .Y(new_n1865_));
  OR4X1    g01801(.A(new_n1865_), .B(new_n1862_), .C(new_n1859_), .D(new_n1500_), .Y(new_n1866_));
  OR4X1    g01802(.A(new_n857_), .B(new_n659_), .C(new_n586_), .D(new_n547_), .Y(new_n1867_));
  OR2X1    g01803(.A(new_n1459_), .B(new_n1090_), .Y(new_n1868_));
  OR4X1    g01804(.A(new_n1868_), .B(new_n1332_), .C(new_n1133_), .D(new_n489_), .Y(new_n1869_));
  OAI22X1  g01805(.A0(new_n152_), .A1(new_n108_), .B0(new_n96_), .B1(new_n81_), .Y(new_n1870_));
  OR4X1    g01806(.A(new_n540_), .B(new_n400_), .C(new_n260_), .D(new_n850_), .Y(new_n1871_));
  OR4X1    g01807(.A(new_n1871_), .B(new_n1870_), .C(new_n1615_), .D(new_n308_), .Y(new_n1872_));
  OR4X1    g01808(.A(new_n292_), .B(new_n201_), .C(new_n191_), .D(new_n981_), .Y(new_n1873_));
  OR4X1    g01809(.A(new_n1873_), .B(new_n579_), .C(new_n968_), .D(new_n387_), .Y(new_n1874_));
  OR4X1    g01810(.A(new_n383_), .B(new_n797_), .C(new_n213_), .D(new_n379_), .Y(new_n1875_));
  OR4X1    g01811(.A(new_n412_), .B(new_n928_), .C(new_n120_), .D(new_n100_), .Y(new_n1876_));
  OR4X1    g01812(.A(new_n1876_), .B(new_n1875_), .C(new_n1874_), .D(new_n1872_), .Y(new_n1877_));
  OR4X1    g01813(.A(new_n1877_), .B(new_n1869_), .C(new_n1867_), .D(new_n1866_), .Y(new_n1878_));
  NOR2X1   g01814(.A(new_n1878_), .B(new_n1854_), .Y(new_n1879_));
  XOR2X1   g01815(.A(new_n1879_), .B(new_n520_), .Y(new_n1880_));
  XOR2X1   g01816(.A(new_n1880_), .B(new_n1845_), .Y(new_n1881_));
  INVX1    g01817(.A(new_n1881_), .Y(new_n1882_));
  XOR2X1   g01818(.A(\a[31] ), .B(new_n68_), .Y(new_n1883_));
  NOR2X1   g01819(.A(new_n1883_), .B(new_n406_), .Y(new_n1884_));
  INVX1    g01820(.A(new_n1884_), .Y(new_n1885_));
  INVX1    g01821(.A(new_n623_), .Y(new_n1886_));
  INVX1    g01822(.A(new_n1879_), .Y(new_n1887_));
  INVX1    g01823(.A(\a[31] ), .Y(new_n1888_));
  AND2X1   g01824(.A(new_n406_), .B(new_n1888_), .Y(new_n1889_));
  NOR3X1   g01825(.A(new_n1888_), .B(new_n68_), .C(new_n74_), .Y(new_n1890_));
  AOI22X1  g01826(.A0(new_n1890_), .A1(new_n1886_), .B0(new_n1889_), .B1(new_n1887_), .Y(new_n1891_));
  OAI21X1  g01827(.A0(new_n1885_), .A1(new_n520_), .B0(new_n1891_), .Y(new_n1892_));
  AOI21X1  g01828(.A0(new_n1882_), .A1(new_n407_), .B0(new_n1892_), .Y(new_n1893_));
  OAI22X1  g01829(.A0(new_n161_), .A1(new_n115_), .B0(new_n119_), .B1(new_n94_), .Y(new_n1894_));
  OR2X1    g01830(.A(new_n1894_), .B(new_n720_), .Y(new_n1895_));
  OR4X1    g01831(.A(new_n968_), .B(new_n372_), .C(new_n265_), .D(new_n410_), .Y(new_n1896_));
  OR4X1    g01832(.A(new_n1896_), .B(new_n1895_), .C(new_n850_), .D(new_n228_), .Y(new_n1897_));
  OAI22X1  g01833(.A0(new_n129_), .A1(new_n117_), .B0(new_n78_), .B1(new_n69_), .Y(new_n1898_));
  OR4X1    g01834(.A(new_n1701_), .B(new_n1898_), .C(new_n750_), .D(new_n618_), .Y(new_n1899_));
  OAI22X1  g01835(.A0(new_n182_), .A1(new_n69_), .B0(new_n131_), .B1(new_n117_), .Y(new_n1900_));
  OR4X1    g01836(.A(new_n400_), .B(new_n292_), .C(new_n1087_), .D(new_n884_), .Y(new_n1901_));
  OR4X1    g01837(.A(new_n1901_), .B(new_n1900_), .C(new_n1899_), .D(new_n527_), .Y(new_n1902_));
  OR4X1    g01838(.A(new_n627_), .B(new_n312_), .C(new_n1008_), .D(new_n1284_), .Y(new_n1903_));
  OR4X1    g01839(.A(new_n1903_), .B(new_n1902_), .C(new_n1897_), .D(new_n601_), .Y(new_n1904_));
  INVX1    g01840(.A(new_n286_), .Y(new_n1905_));
  NAND3X1  g01841(.A(new_n503_), .B(new_n1468_), .C(new_n1905_), .Y(new_n1906_));
  AOI21X1  g01842(.A0(new_n152_), .A1(new_n84_), .B0(new_n129_), .Y(new_n1907_));
  OR4X1    g01843(.A(new_n1907_), .B(new_n1906_), .C(new_n1750_), .D(new_n1436_), .Y(new_n1908_));
  OAI22X1  g01844(.A0(new_n161_), .A1(new_n102_), .B0(new_n129_), .B1(new_n123_), .Y(new_n1909_));
  OAI22X1  g01845(.A0(new_n161_), .A1(new_n79_), .B0(new_n131_), .B1(new_n96_), .Y(new_n1910_));
  OAI22X1  g01846(.A0(new_n117_), .A1(new_n78_), .B0(new_n91_), .B1(new_n90_), .Y(new_n1911_));
  AOI21X1  g01847(.A0(new_n152_), .A1(new_n106_), .B0(new_n81_), .Y(new_n1912_));
  OR4X1    g01848(.A(new_n1912_), .B(new_n1911_), .C(new_n1910_), .D(new_n1909_), .Y(new_n1913_));
  OR4X1    g01849(.A(new_n1336_), .B(new_n947_), .C(new_n1002_), .D(new_n513_), .Y(new_n1914_));
  OAI22X1  g01850(.A0(new_n125_), .A1(new_n102_), .B0(new_n81_), .B1(new_n69_), .Y(new_n1915_));
  OR2X1    g01851(.A(new_n1915_), .B(new_n843_), .Y(new_n1916_));
  OR4X1    g01852(.A(new_n1916_), .B(new_n594_), .C(new_n229_), .D(new_n746_), .Y(new_n1917_));
  OR4X1    g01853(.A(new_n1917_), .B(new_n1914_), .C(new_n1913_), .D(new_n1908_), .Y(new_n1918_));
  OR4X1    g01854(.A(new_n1918_), .B(new_n1904_), .C(new_n1569_), .D(new_n822_), .Y(new_n1919_));
  INVX1    g01855(.A(\a[20] ), .Y(new_n1920_));
  OR2X1    g01856(.A(new_n656_), .B(new_n338_), .Y(new_n1921_));
  OR4X1    g01857(.A(new_n1028_), .B(new_n505_), .C(new_n382_), .D(new_n303_), .Y(new_n1922_));
  OAI22X1  g01858(.A0(new_n182_), .A1(new_n123_), .B0(new_n152_), .B1(new_n92_), .Y(new_n1923_));
  NOR4X1   g01859(.A(new_n1923_), .B(new_n1922_), .C(new_n1921_), .D(new_n169_), .Y(new_n1924_));
  OR4X1    g01860(.A(new_n531_), .B(new_n1467_), .C(new_n568_), .D(new_n1057_), .Y(new_n1925_));
  NOR4X1   g01861(.A(new_n1925_), .B(new_n1426_), .C(new_n787_), .D(new_n667_), .Y(new_n1926_));
  NAND4X1  g01862(.A(new_n1926_), .B(new_n1924_), .C(new_n1149_), .D(new_n914_), .Y(new_n1927_));
  OR4X1    g01863(.A(new_n1717_), .B(new_n1703_), .C(new_n617_), .D(new_n342_), .Y(new_n1928_));
  OR4X1    g01864(.A(new_n634_), .B(new_n412_), .C(new_n408_), .D(new_n998_), .Y(new_n1929_));
  OR4X1    g01865(.A(new_n479_), .B(new_n191_), .C(new_n381_), .D(new_n449_), .Y(new_n1930_));
  OR4X1    g01866(.A(new_n1930_), .B(new_n1929_), .C(new_n1894_), .D(new_n720_), .Y(new_n1931_));
  OR4X1    g01867(.A(new_n193_), .B(new_n431_), .C(new_n1008_), .D(new_n1284_), .Y(new_n1932_));
  INVX1    g01868(.A(new_n585_), .Y(new_n1933_));
  NAND3X1  g01869(.A(new_n861_), .B(new_n776_), .C(new_n1933_), .Y(new_n1934_));
  OR4X1    g01870(.A(new_n1934_), .B(new_n460_), .C(new_n386_), .D(new_n615_), .Y(new_n1935_));
  OR4X1    g01871(.A(new_n1935_), .B(new_n1932_), .C(new_n710_), .D(new_n666_), .Y(new_n1936_));
  OR4X1    g01872(.A(new_n1936_), .B(new_n1931_), .C(new_n1928_), .D(new_n1349_), .Y(new_n1937_));
  OR4X1    g01873(.A(new_n1732_), .B(new_n1017_), .C(new_n891_), .D(new_n147_), .Y(new_n1938_));
  OR4X1    g01874(.A(new_n1336_), .B(new_n1105_), .C(new_n239_), .D(new_n648_), .Y(new_n1939_));
  INVX1    g01875(.A(new_n603_), .Y(new_n1940_));
  NAND3X1  g01876(.A(new_n1940_), .B(new_n1343_), .C(new_n818_), .Y(new_n1941_));
  OR4X1    g01877(.A(new_n1941_), .B(new_n1939_), .C(new_n1006_), .D(new_n951_), .Y(new_n1942_));
  OR4X1    g01878(.A(new_n228_), .B(new_n176_), .C(new_n981_), .D(new_n86_), .Y(new_n1943_));
  OR4X1    g01879(.A(new_n1943_), .B(new_n541_), .C(new_n356_), .D(new_n304_), .Y(new_n1944_));
  OR2X1    g01880(.A(new_n1541_), .B(new_n504_), .Y(new_n1945_));
  NOR4X1   g01881(.A(new_n1945_), .B(new_n1944_), .C(new_n1942_), .D(new_n1938_), .Y(new_n1946_));
  INVX1    g01882(.A(new_n1946_), .Y(new_n1947_));
  NOR3X1   g01883(.A(new_n1947_), .B(new_n1937_), .C(new_n1927_), .Y(new_n1948_));
  OR4X1    g01884(.A(new_n1106_), .B(new_n716_), .C(new_n311_), .D(new_n992_), .Y(new_n1949_));
  OAI22X1  g01885(.A0(new_n148_), .A1(new_n129_), .B0(new_n106_), .B1(new_n78_), .Y(new_n1950_));
  OR2X1    g01886(.A(new_n1950_), .B(new_n422_), .Y(new_n1951_));
  OR4X1    g01887(.A(new_n206_), .B(new_n181_), .C(new_n431_), .D(new_n118_), .Y(new_n1952_));
  OR4X1    g01888(.A(new_n1952_), .B(new_n1951_), .C(new_n569_), .D(new_n259_), .Y(new_n1953_));
  OR4X1    g01889(.A(new_n603_), .B(new_n296_), .C(new_n184_), .D(new_n114_), .Y(new_n1954_));
  OR4X1    g01890(.A(new_n418_), .B(new_n382_), .C(new_n691_), .D(new_n175_), .Y(new_n1955_));
  OR4X1    g01891(.A(new_n1955_), .B(new_n509_), .C(new_n506_), .D(new_n468_), .Y(new_n1956_));
  OR4X1    g01892(.A(new_n1956_), .B(new_n1954_), .C(new_n608_), .D(new_n571_), .Y(new_n1957_));
  OR4X1    g01893(.A(new_n1957_), .B(new_n1953_), .C(new_n1949_), .D(new_n1180_), .Y(new_n1958_));
  OR4X1    g01894(.A(new_n636_), .B(new_n354_), .C(new_n483_), .D(new_n191_), .Y(new_n1959_));
  OR4X1    g01895(.A(new_n1959_), .B(new_n312_), .C(new_n1008_), .D(new_n307_), .Y(new_n1960_));
  OR4X1    g01896(.A(new_n1261_), .B(new_n850_), .C(new_n757_), .D(new_n327_), .Y(new_n1961_));
  OAI22X1  g01897(.A0(new_n131_), .A1(new_n119_), .B0(new_n123_), .B1(new_n108_), .Y(new_n1962_));
  OAI22X1  g01898(.A0(new_n161_), .A1(new_n96_), .B0(new_n143_), .B1(new_n91_), .Y(new_n1963_));
  OR4X1    g01899(.A(new_n1963_), .B(new_n1962_), .C(new_n1961_), .D(new_n1960_), .Y(new_n1964_));
  OAI22X1  g01900(.A0(new_n182_), .A1(new_n148_), .B0(new_n152_), .B1(new_n90_), .Y(new_n1965_));
  AOI21X1  g01901(.A0(new_n182_), .A1(new_n161_), .B0(new_n152_), .Y(new_n1966_));
  OR4X1    g01902(.A(new_n1966_), .B(new_n1779_), .C(new_n1965_), .D(new_n565_), .Y(new_n1967_));
  OR4X1    g01903(.A(new_n945_), .B(new_n931_), .C(new_n741_), .D(new_n459_), .Y(new_n1968_));
  OR4X1    g01904(.A(new_n750_), .B(new_n728_), .C(new_n641_), .D(new_n1467_), .Y(new_n1969_));
  NOR4X1   g01905(.A(new_n1969_), .B(new_n1968_), .C(new_n1967_), .D(new_n1964_), .Y(new_n1970_));
  OR2X1    g01906(.A(new_n1576_), .B(new_n197_), .Y(new_n1971_));
  OR4X1    g01907(.A(new_n1646_), .B(new_n444_), .C(new_n381_), .D(new_n158_), .Y(new_n1972_));
  OAI22X1  g01908(.A0(new_n182_), .A1(new_n117_), .B0(new_n106_), .B1(new_n92_), .Y(new_n1973_));
  OR2X1    g01909(.A(new_n1973_), .B(new_n586_), .Y(new_n1974_));
  OAI22X1  g01910(.A0(new_n129_), .A1(new_n79_), .B0(new_n105_), .B1(new_n84_), .Y(new_n1975_));
  OR4X1    g01911(.A(new_n1975_), .B(new_n1974_), .C(new_n1972_), .D(new_n632_), .Y(new_n1976_));
  NOR2X1   g01912(.A(new_n276_), .B(new_n449_), .Y(new_n1977_));
  INVX1    g01913(.A(new_n1977_), .Y(new_n1978_));
  OAI22X1  g01914(.A0(new_n168_), .A1(new_n72_), .B0(new_n117_), .B1(new_n94_), .Y(new_n1979_));
  OR4X1    g01915(.A(new_n1979_), .B(new_n1227_), .C(new_n657_), .D(new_n1978_), .Y(new_n1980_));
  OR4X1    g01916(.A(new_n702_), .B(new_n371_), .C(new_n193_), .D(new_n86_), .Y(new_n1981_));
  NOR4X1   g01917(.A(new_n1981_), .B(new_n1980_), .C(new_n1976_), .D(new_n1971_), .Y(new_n1982_));
  NOR4X1   g01918(.A(new_n251_), .B(new_n200_), .C(new_n199_), .D(new_n187_), .Y(new_n1983_));
  AOI21X1  g01919(.A0(new_n143_), .A1(new_n94_), .B0(new_n69_), .Y(new_n1984_));
  NOR3X1   g01920(.A(new_n1984_), .B(new_n226_), .C(new_n213_), .Y(new_n1985_));
  NOR3X1   g01921(.A(new_n720_), .B(new_n383_), .C(new_n885_), .Y(new_n1986_));
  NOR4X1   g01922(.A(new_n280_), .B(new_n273_), .C(new_n398_), .D(new_n664_), .Y(new_n1987_));
  NAND4X1  g01923(.A(new_n1987_), .B(new_n1986_), .C(new_n1985_), .D(new_n1983_), .Y(new_n1988_));
  OAI22X1  g01924(.A0(new_n127_), .A1(new_n96_), .B0(new_n108_), .B1(new_n84_), .Y(new_n1989_));
  OR4X1    g01925(.A(new_n1142_), .B(new_n1989_), .C(new_n133_), .D(new_n535_), .Y(new_n1990_));
  OR4X1    g01926(.A(new_n1990_), .B(new_n815_), .C(new_n521_), .D(new_n80_), .Y(new_n1991_));
  NOR2X1   g01927(.A(new_n1991_), .B(new_n1988_), .Y(new_n1992_));
  NAND3X1  g01928(.A(new_n1992_), .B(new_n1982_), .C(new_n1970_), .Y(new_n1993_));
  NOR2X1   g01929(.A(new_n1993_), .B(new_n1958_), .Y(new_n1994_));
  NOR2X1   g01930(.A(new_n1994_), .B(new_n1948_), .Y(new_n1995_));
  NAND2X1  g01931(.A(new_n1994_), .B(new_n1948_), .Y(new_n1996_));
  AOI21X1  g01932(.A0(new_n1996_), .A1(new_n1920_), .B0(new_n1995_), .Y(new_n1997_));
  XOR2X1   g01933(.A(new_n1997_), .B(new_n1919_), .Y(new_n1998_));
  XOR2X1   g01934(.A(new_n1998_), .B(new_n1893_), .Y(new_n1999_));
  NOR3X1   g01935(.A(new_n741_), .B(new_n589_), .C(new_n1166_), .Y(new_n2000_));
  NOR2X1   g01936(.A(new_n142_), .B(new_n1008_), .Y(new_n2001_));
  NOR4X1   g01937(.A(new_n612_), .B(new_n361_), .C(new_n758_), .D(new_n175_), .Y(new_n2002_));
  NAND3X1  g01938(.A(new_n2002_), .B(new_n2001_), .C(new_n2000_), .Y(new_n2003_));
  OAI22X1  g01939(.A0(new_n143_), .A1(new_n88_), .B0(new_n108_), .B1(new_n75_), .Y(new_n2004_));
  OR2X1    g01940(.A(new_n2004_), .B(new_n474_), .Y(new_n2005_));
  OR2X1    g01941(.A(new_n444_), .B(new_n313_), .Y(new_n2006_));
  OR4X1    g01942(.A(new_n478_), .B(new_n217_), .C(new_n381_), .D(new_n155_), .Y(new_n2007_));
  NAND3X1  g01943(.A(new_n364_), .B(new_n1905_), .C(new_n279_), .Y(new_n2008_));
  OR4X1    g01944(.A(new_n2008_), .B(new_n2007_), .C(new_n2006_), .D(new_n2005_), .Y(new_n2009_));
  OR4X1    g01945(.A(new_n848_), .B(new_n723_), .C(new_n586_), .D(new_n740_), .Y(new_n2010_));
  OR4X1    g01946(.A(new_n2010_), .B(new_n714_), .C(new_n386_), .D(new_n431_), .Y(new_n2011_));
  OR4X1    g01947(.A(new_n1156_), .B(new_n716_), .C(new_n569_), .D(new_n561_), .Y(new_n2012_));
  OR4X1    g01948(.A(new_n2012_), .B(new_n2011_), .C(new_n2009_), .D(new_n2003_), .Y(new_n2013_));
  OAI22X1  g01949(.A0(new_n131_), .A1(new_n88_), .B0(new_n127_), .B1(new_n69_), .Y(new_n2014_));
  OR4X1    g01950(.A(new_n2014_), .B(new_n968_), .C(new_n1087_), .D(new_n610_), .Y(new_n2015_));
  OR4X1    g01951(.A(new_n547_), .B(new_n615_), .C(new_n814_), .D(new_n251_), .Y(new_n2016_));
  OR4X1    g01952(.A(new_n2016_), .B(new_n2015_), .C(new_n1461_), .D(new_n772_), .Y(new_n2017_));
  OR4X1    g01953(.A(new_n634_), .B(new_n802_), .C(new_n264_), .D(new_n792_), .Y(new_n2018_));
  OR4X1    g01954(.A(new_n931_), .B(new_n243_), .C(new_n133_), .D(new_n114_), .Y(new_n2019_));
  OAI22X1  g01955(.A0(new_n131_), .A1(new_n106_), .B0(new_n105_), .B1(new_n69_), .Y(new_n2020_));
  OR4X1    g01956(.A(new_n240_), .B(new_n296_), .C(new_n187_), .D(new_n928_), .Y(new_n2021_));
  NOR4X1   g01957(.A(new_n2021_), .B(new_n2020_), .C(new_n1725_), .D(new_n636_), .Y(new_n2022_));
  NOR3X1   g01958(.A(new_n537_), .B(new_n505_), .C(new_n158_), .Y(new_n2023_));
  NOR4X1   g01959(.A(new_n594_), .B(new_n439_), .C(new_n379_), .D(new_n651_), .Y(new_n2024_));
  NAND4X1  g01960(.A(new_n2024_), .B(new_n2023_), .C(new_n2022_), .D(new_n1857_), .Y(new_n2025_));
  OR4X1    g01961(.A(new_n2025_), .B(new_n2019_), .C(new_n2018_), .D(new_n2017_), .Y(new_n2026_));
  NOR3X1   g01962(.A(new_n265_), .B(new_n138_), .C(new_n116_), .Y(new_n2027_));
  NOR3X1   g01963(.A(new_n702_), .B(new_n370_), .C(new_n156_), .Y(new_n2028_));
  NAND3X1  g01964(.A(new_n2028_), .B(new_n2027_), .C(new_n841_), .Y(new_n2029_));
  OR4X1    g01965(.A(new_n480_), .B(new_n414_), .C(new_n356_), .D(new_n691_), .Y(new_n2030_));
  OR4X1    g01966(.A(new_n2030_), .B(new_n1361_), .C(new_n750_), .D(new_n803_), .Y(new_n2031_));
  OR4X1    g01967(.A(new_n2031_), .B(new_n2029_), .C(new_n1498_), .D(new_n584_), .Y(new_n2032_));
  NOR3X1   g01968(.A(new_n2032_), .B(new_n2026_), .C(new_n2013_), .Y(new_n2033_));
  NOR4X1   g01969(.A(new_n2033_), .B(new_n1947_), .C(new_n1937_), .D(new_n1927_), .Y(new_n2034_));
  XOR2X1   g01970(.A(new_n1841_), .B(new_n1839_), .Y(new_n2035_));
  INVX1    g01971(.A(new_n783_), .Y(new_n2036_));
  AOI22X1  g01972(.A0(new_n1890_), .A1(new_n2036_), .B0(new_n1889_), .B1(new_n1886_), .Y(new_n2037_));
  OAI21X1  g01973(.A0(new_n1885_), .A1(new_n690_), .B0(new_n2037_), .Y(new_n2038_));
  AOI21X1  g01974(.A0(new_n2035_), .A1(new_n407_), .B0(new_n2038_), .Y(new_n2039_));
  NOR4X1   g01975(.A(new_n2032_), .B(new_n2026_), .C(new_n2013_), .D(new_n1948_), .Y(new_n2040_));
  NOR3X1   g01976(.A(new_n2040_), .B(new_n2039_), .C(new_n2034_), .Y(new_n2041_));
  NOR2X1   g01977(.A(new_n2041_), .B(new_n2034_), .Y(new_n2042_));
  NOR2X1   g01978(.A(new_n1995_), .B(\a[20] ), .Y(new_n2043_));
  AOI21X1  g01979(.A0(new_n2043_), .A1(new_n1996_), .B0(\a[20] ), .Y(new_n2044_));
  AOI21X1  g01980(.A0(new_n1997_), .A1(new_n1996_), .B0(new_n2044_), .Y(new_n2045_));
  NOR2X1   g01981(.A(new_n2045_), .B(new_n2042_), .Y(new_n2046_));
  XOR2X1   g01982(.A(new_n1844_), .B(new_n1843_), .Y(new_n2047_));
  INVX1    g01983(.A(new_n520_), .Y(new_n2048_));
  INVX1    g01984(.A(new_n690_), .Y(new_n2049_));
  AOI22X1  g01985(.A0(new_n1890_), .A1(new_n2049_), .B0(new_n1889_), .B1(new_n2048_), .Y(new_n2050_));
  OAI21X1  g01986(.A0(new_n1885_), .A1(new_n623_), .B0(new_n2050_), .Y(new_n2051_));
  AOI21X1  g01987(.A0(new_n2047_), .A1(new_n407_), .B0(new_n2051_), .Y(new_n2052_));
  INVX1    g01988(.A(new_n2052_), .Y(new_n2053_));
  XOR2X1   g01989(.A(new_n2045_), .B(new_n2042_), .Y(new_n2054_));
  AOI21X1  g01990(.A0(new_n2054_), .A1(new_n2053_), .B0(new_n2046_), .Y(new_n2055_));
  NOR2X1   g01991(.A(new_n2055_), .B(new_n1999_), .Y(new_n2056_));
  INVX1    g01992(.A(new_n2056_), .Y(new_n2057_));
  INVX1    g01993(.A(new_n1999_), .Y(new_n2058_));
  XOR2X1   g01994(.A(new_n2055_), .B(new_n2058_), .Y(new_n2059_));
  XOR2X1   g01995(.A(\a[29] ), .B(new_n95_), .Y(new_n2060_));
  XOR2X1   g01996(.A(\a[27] ), .B(new_n89_), .Y(new_n2061_));
  NOR2X1   g01997(.A(new_n2061_), .B(new_n2060_), .Y(new_n2062_));
  INVX1    g01998(.A(new_n2062_), .Y(new_n2063_));
  OR4X1    g01999(.A(new_n1538_), .B(new_n1407_), .C(new_n252_), .D(new_n213_), .Y(new_n2064_));
  AOI21X1  g02000(.A0(new_n105_), .A1(new_n78_), .B0(new_n91_), .Y(new_n2065_));
  OR2X1    g02001(.A(new_n522_), .B(new_n2065_), .Y(new_n2066_));
  OR4X1    g02002(.A(new_n594_), .B(new_n541_), .C(new_n231_), .D(new_n103_), .Y(new_n2067_));
  OR2X1    g02003(.A(new_n2067_), .B(new_n2066_), .Y(new_n2068_));
  AOI21X1  g02004(.A0(new_n143_), .A1(new_n90_), .B0(new_n117_), .Y(new_n2069_));
  OR4X1    g02005(.A(new_n2069_), .B(new_n579_), .C(new_n372_), .D(new_n840_), .Y(new_n2070_));
  OR4X1    g02006(.A(new_n2070_), .B(new_n2068_), .C(new_n2064_), .D(new_n1508_), .Y(new_n2071_));
  OAI22X1  g02007(.A0(new_n127_), .A1(new_n91_), .B0(new_n125_), .B1(new_n84_), .Y(new_n2072_));
  OAI22X1  g02008(.A0(new_n129_), .A1(new_n106_), .B0(new_n79_), .B1(new_n78_), .Y(new_n2073_));
  OR4X1    g02009(.A(new_n2073_), .B(new_n2072_), .C(new_n1018_), .D(new_n193_), .Y(new_n2074_));
  OR4X1    g02010(.A(new_n1028_), .B(new_n631_), .C(new_n387_), .D(new_n201_), .Y(new_n2075_));
  OR4X1    g02011(.A(new_n2075_), .B(new_n465_), .C(new_n232_), .D(new_n124_), .Y(new_n2076_));
  OR4X1    g02012(.A(new_n328_), .B(new_n286_), .C(new_n398_), .D(new_n224_), .Y(new_n2077_));
  OR4X1    g02013(.A(new_n226_), .B(new_n172_), .C(new_n118_), .D(new_n1284_), .Y(new_n2078_));
  OR4X1    g02014(.A(new_n2078_), .B(new_n2077_), .C(new_n2076_), .D(new_n2074_), .Y(new_n2079_));
  NOR4X1   g02015(.A(new_n678_), .B(new_n261_), .C(new_n256_), .D(new_n234_), .Y(new_n2080_));
  NOR3X1   g02016(.A(new_n500_), .B(new_n740_), .C(new_n819_), .Y(new_n2081_));
  NAND3X1  g02017(.A(new_n2081_), .B(new_n2080_), .C(new_n1368_), .Y(new_n2082_));
  OR4X1    g02018(.A(new_n2082_), .B(new_n2079_), .C(new_n2071_), .D(new_n1247_), .Y(new_n2083_));
  OAI22X1  g02019(.A0(new_n125_), .A1(new_n75_), .B0(new_n90_), .B1(new_n69_), .Y(new_n2084_));
  OR4X1    g02020(.A(new_n2084_), .B(new_n1156_), .C(new_n560_), .D(new_n1166_), .Y(new_n2085_));
  OAI21X1  g02021(.A0(new_n81_), .A1(new_n69_), .B0(new_n776_), .Y(new_n2086_));
  OR4X1    g02022(.A(new_n2086_), .B(new_n358_), .C(new_n348_), .D(new_n300_), .Y(new_n2087_));
  OAI22X1  g02023(.A0(new_n152_), .A1(new_n78_), .B0(new_n131_), .B1(new_n96_), .Y(new_n2088_));
  OAI22X1  g02024(.A0(new_n127_), .A1(new_n115_), .B0(new_n117_), .B1(new_n94_), .Y(new_n2089_));
  OR4X1    g02025(.A(new_n2089_), .B(new_n2088_), .C(new_n1403_), .D(new_n1227_), .Y(new_n2090_));
  OR4X1    g02026(.A(new_n2090_), .B(new_n2087_), .C(new_n2085_), .D(new_n278_), .Y(new_n2091_));
  NOR3X1   g02027(.A(new_n2091_), .B(new_n2083_), .C(new_n438_), .Y(new_n2092_));
  INVX1    g02028(.A(new_n2092_), .Y(new_n2093_));
  XOR2X1   g02029(.A(\a[28] ), .B(\a[27] ), .Y(new_n2094_));
  AND2X1   g02030(.A(new_n2094_), .B(new_n2061_), .Y(new_n2095_));
  OR4X1    g02031(.A(new_n1473_), .B(new_n720_), .C(new_n229_), .D(new_n449_), .Y(new_n2096_));
  OAI22X1  g02032(.A0(new_n182_), .A1(new_n69_), .B0(new_n152_), .B1(new_n94_), .Y(new_n2097_));
  OR4X1    g02033(.A(new_n1923_), .B(new_n951_), .C(new_n714_), .D(new_n837_), .Y(new_n2098_));
  OR4X1    g02034(.A(new_n2098_), .B(new_n2097_), .C(new_n1096_), .D(new_n959_), .Y(new_n2099_));
  OR4X1    g02035(.A(new_n603_), .B(new_n208_), .C(new_n757_), .D(new_n581_), .Y(new_n2100_));
  AOI21X1  g02036(.A0(new_n182_), .A1(new_n78_), .B0(new_n119_), .Y(new_n2101_));
  OR4X1    g02037(.A(new_n2101_), .B(new_n2100_), .C(new_n887_), .D(new_n511_), .Y(new_n2102_));
  INVX1    g02038(.A(new_n2023_), .Y(new_n2103_));
  OR4X1    g02039(.A(new_n500_), .B(new_n480_), .C(new_n1261_), .D(new_n100_), .Y(new_n2104_));
  OR2X1    g02040(.A(new_n1316_), .B(new_n465_), .Y(new_n2105_));
  OR4X1    g02041(.A(new_n2105_), .B(new_n2104_), .C(new_n2103_), .D(new_n897_), .Y(new_n2106_));
  NOR4X1   g02042(.A(new_n2106_), .B(new_n2102_), .C(new_n2099_), .D(new_n2096_), .Y(new_n2107_));
  INVX1    g02043(.A(new_n2107_), .Y(new_n2108_));
  NOR4X1   g02044(.A(new_n1990_), .B(new_n815_), .C(new_n521_), .D(new_n80_), .Y(new_n2109_));
  NOR3X1   g02045(.A(new_n421_), .B(new_n522_), .C(new_n103_), .Y(new_n2110_));
  NOR2X1   g02046(.A(new_n825_), .B(new_n303_), .Y(new_n2111_));
  NOR4X1   g02047(.A(new_n594_), .B(new_n968_), .C(new_n274_), .D(new_n224_), .Y(new_n2112_));
  NAND3X1  g02048(.A(new_n2112_), .B(new_n2111_), .C(new_n2110_), .Y(new_n2113_));
  OR4X1    g02049(.A(new_n547_), .B(new_n615_), .C(new_n252_), .D(new_n159_), .Y(new_n2114_));
  OR4X1    g02050(.A(new_n2114_), .B(new_n1276_), .C(new_n504_), .D(new_n300_), .Y(new_n2115_));
  OR4X1    g02051(.A(new_n280_), .B(new_n539_), .C(new_n207_), .D(new_n1284_), .Y(new_n2116_));
  OR4X1    g02052(.A(new_n2116_), .B(new_n527_), .C(new_n348_), .D(new_n400_), .Y(new_n2117_));
  OR4X1    g02053(.A(new_n1635_), .B(new_n1028_), .C(new_n354_), .D(new_n717_), .Y(new_n2118_));
  OR4X1    g02054(.A(new_n975_), .B(new_n276_), .C(new_n138_), .D(new_n651_), .Y(new_n2119_));
  OR4X1    g02055(.A(new_n2119_), .B(new_n2118_), .C(new_n2117_), .D(new_n2115_), .Y(new_n2120_));
  NOR2X1   g02056(.A(new_n2120_), .B(new_n2113_), .Y(new_n2121_));
  OAI21X1  g02057(.A0(new_n99_), .A1(new_n75_), .B0(new_n341_), .Y(new_n2122_));
  OR4X1    g02058(.A(new_n2122_), .B(new_n602_), .C(new_n490_), .D(new_n335_), .Y(new_n2123_));
  OAI22X1  g02059(.A0(new_n131_), .A1(new_n102_), .B0(new_n123_), .B1(new_n81_), .Y(new_n2124_));
  OR2X1    g02060(.A(new_n2124_), .B(new_n321_), .Y(new_n2125_));
  OR4X1    g02061(.A(new_n632_), .B(new_n541_), .C(new_n509_), .D(new_n328_), .Y(new_n2126_));
  OR4X1    g02062(.A(new_n947_), .B(new_n385_), .C(new_n379_), .D(new_n141_), .Y(new_n2127_));
  OR4X1    g02063(.A(new_n1757_), .B(new_n1384_), .C(new_n873_), .D(new_n728_), .Y(new_n2128_));
  OR2X1    g02064(.A(new_n2128_), .B(new_n2127_), .Y(new_n2129_));
  NOR4X1   g02065(.A(new_n2129_), .B(new_n2126_), .C(new_n2125_), .D(new_n2123_), .Y(new_n2130_));
  OR4X1    g02066(.A(new_n429_), .B(new_n396_), .C(new_n598_), .D(new_n293_), .Y(new_n2131_));
  OR4X1    g02067(.A(new_n457_), .B(new_n203_), .C(new_n327_), .D(new_n585_), .Y(new_n2132_));
  OAI22X1  g02068(.A0(new_n148_), .A1(new_n78_), .B0(new_n129_), .B1(new_n96_), .Y(new_n2133_));
  OR2X1    g02069(.A(new_n2133_), .B(new_n636_), .Y(new_n2134_));
  NOR4X1   g02070(.A(new_n2134_), .B(new_n2132_), .C(new_n2131_), .D(new_n1593_), .Y(new_n2135_));
  NAND4X1  g02071(.A(new_n2135_), .B(new_n2130_), .C(new_n2121_), .D(new_n2109_), .Y(new_n2136_));
  NOR2X1   g02072(.A(new_n2136_), .B(new_n2108_), .Y(new_n2137_));
  INVX1    g02073(.A(new_n2060_), .Y(new_n2138_));
  NOR2X1   g02074(.A(new_n2061_), .B(new_n2138_), .Y(new_n2139_));
  INVX1    g02075(.A(new_n2139_), .Y(new_n2140_));
  OAI22X1  g02076(.A0(new_n117_), .A1(new_n99_), .B0(new_n88_), .B1(new_n78_), .Y(new_n2141_));
  OR4X1    g02077(.A(new_n2141_), .B(new_n1493_), .C(new_n1415_), .D(new_n1402_), .Y(new_n2142_));
  NOR4X1   g02078(.A(new_n280_), .B(new_n797_), .C(new_n264_), .D(new_n223_), .Y(new_n2143_));
  NOR4X1   g02079(.A(new_n1000_), .B(new_n994_), .C(new_n829_), .D(new_n515_), .Y(new_n2144_));
  NAND2X1  g02080(.A(new_n2144_), .B(new_n2143_), .Y(new_n2145_));
  OR4X1    g02081(.A(new_n1459_), .B(new_n1142_), .C(new_n608_), .D(new_n289_), .Y(new_n2146_));
  OR4X1    g02082(.A(new_n2146_), .B(new_n1398_), .C(new_n1261_), .D(new_n840_), .Y(new_n2147_));
  OR4X1    g02083(.A(new_n2147_), .B(new_n2145_), .C(new_n2142_), .D(new_n683_), .Y(new_n2148_));
  INVX1    g02084(.A(new_n338_), .Y(new_n2149_));
  INVX1    g02085(.A(new_n386_), .Y(new_n2150_));
  NAND3X1  g02086(.A(new_n2150_), .B(new_n2149_), .C(new_n1741_), .Y(new_n2151_));
  OR4X1    g02087(.A(new_n408_), .B(new_n396_), .C(new_n260_), .D(new_n80_), .Y(new_n2152_));
  OAI22X1  g02088(.A0(new_n152_), .A1(new_n125_), .B0(new_n119_), .B1(new_n92_), .Y(new_n2153_));
  OAI22X1  g02089(.A0(new_n129_), .A1(new_n117_), .B0(new_n123_), .B1(new_n108_), .Y(new_n2154_));
  OR4X1    g02090(.A(new_n2154_), .B(new_n2153_), .C(new_n891_), .D(new_n723_), .Y(new_n2155_));
  OR4X1    g02091(.A(new_n2155_), .B(new_n2152_), .C(new_n2151_), .D(new_n2148_), .Y(new_n2156_));
  OAI22X1  g02092(.A0(new_n143_), .A1(new_n115_), .B0(new_n131_), .B1(new_n91_), .Y(new_n2157_));
  OR4X1    g02093(.A(new_n2157_), .B(new_n1225_), .C(new_n370_), .D(new_n173_), .Y(new_n2158_));
  OR4X1    g02094(.A(new_n1210_), .B(new_n896_), .C(new_n666_), .D(new_n803_), .Y(new_n2159_));
  INVX1    g02095(.A(new_n220_), .Y(new_n2160_));
  INVX1    g02096(.A(new_n294_), .Y(new_n2161_));
  NAND3X1  g02097(.A(new_n2161_), .B(new_n2160_), .C(new_n326_), .Y(new_n2162_));
  OR4X1    g02098(.A(new_n2162_), .B(new_n1044_), .C(new_n375_), .D(new_n116_), .Y(new_n2163_));
  OR4X1    g02099(.A(new_n1426_), .B(new_n777_), .C(new_n226_), .D(new_n648_), .Y(new_n2164_));
  OR4X1    g02100(.A(new_n2164_), .B(new_n510_), .C(new_n350_), .D(new_n142_), .Y(new_n2165_));
  NOR4X1   g02101(.A(new_n355_), .B(new_n354_), .C(new_n536_), .D(new_n149_), .Y(new_n2166_));
  INVX1    g02102(.A(new_n2166_), .Y(new_n2167_));
  NOR4X1   g02103(.A(new_n455_), .B(new_n233_), .C(new_n118_), .D(new_n86_), .Y(new_n2168_));
  INVX1    g02104(.A(new_n2168_), .Y(new_n2169_));
  OR4X1    g02105(.A(new_n2169_), .B(new_n2167_), .C(new_n2165_), .D(new_n722_), .Y(new_n2170_));
  OR4X1    g02106(.A(new_n2170_), .B(new_n2163_), .C(new_n2159_), .D(new_n2158_), .Y(new_n2171_));
  OAI22X1  g02107(.A0(new_n143_), .A1(new_n75_), .B0(new_n115_), .B1(new_n99_), .Y(new_n2172_));
  OR2X1    g02108(.A(new_n2172_), .B(new_n293_), .Y(new_n2173_));
  NOR4X1   g02109(.A(new_n2173_), .B(new_n1701_), .C(new_n478_), .D(new_n155_), .Y(new_n2174_));
  NAND3X1  g02110(.A(new_n2174_), .B(new_n855_), .C(new_n542_), .Y(new_n2175_));
  OR4X1    g02111(.A(new_n505_), .B(new_n276_), .C(new_n850_), .D(new_n219_), .Y(new_n2176_));
  OR4X1    g02112(.A(new_n2176_), .B(new_n755_), .C(new_n757_), .D(new_n103_), .Y(new_n2177_));
  OAI22X1  g02113(.A0(new_n129_), .A1(new_n123_), .B0(new_n108_), .B1(new_n96_), .Y(new_n2178_));
  OR4X1    g02114(.A(new_n2178_), .B(new_n1211_), .C(new_n2097_), .D(new_n673_), .Y(new_n2179_));
  OAI22X1  g02115(.A0(new_n161_), .A1(new_n123_), .B0(new_n143_), .B1(new_n96_), .Y(new_n2180_));
  OR4X1    g02116(.A(new_n2180_), .B(new_n1166_), .C(new_n334_), .D(new_n332_), .Y(new_n2181_));
  OR4X1    g02117(.A(new_n2181_), .B(new_n2179_), .C(new_n2177_), .D(new_n2175_), .Y(new_n2182_));
  NOR3X1   g02118(.A(new_n2182_), .B(new_n2171_), .C(new_n2156_), .Y(new_n2183_));
  INVX1    g02119(.A(new_n2061_), .Y(new_n2184_));
  NOR3X1   g02120(.A(new_n2094_), .B(new_n2184_), .C(new_n2060_), .Y(new_n2185_));
  INVX1    g02121(.A(new_n2185_), .Y(new_n2186_));
  OAI22X1  g02122(.A0(new_n2186_), .A1(new_n2183_), .B0(new_n2140_), .B1(new_n2137_), .Y(new_n2187_));
  AOI21X1  g02123(.A0(new_n2095_), .A1(new_n2093_), .B0(new_n2187_), .Y(new_n2188_));
  NOR2X1   g02124(.A(new_n2183_), .B(new_n1879_), .Y(new_n2189_));
  INVX1    g02125(.A(new_n1845_), .Y(new_n2190_));
  NOR2X1   g02126(.A(new_n1879_), .B(new_n520_), .Y(new_n2191_));
  AOI21X1  g02127(.A0(new_n1880_), .A1(new_n2190_), .B0(new_n2191_), .Y(new_n2192_));
  INVX1    g02128(.A(new_n2192_), .Y(new_n2193_));
  XOR2X1   g02129(.A(new_n2183_), .B(new_n1879_), .Y(new_n2194_));
  AOI21X1  g02130(.A0(new_n2194_), .A1(new_n2193_), .B0(new_n2189_), .Y(new_n2195_));
  XOR2X1   g02131(.A(new_n2183_), .B(new_n2092_), .Y(new_n2196_));
  INVX1    g02132(.A(new_n2196_), .Y(new_n2197_));
  OR2X1    g02133(.A(new_n2197_), .B(new_n2195_), .Y(new_n2198_));
  OAI21X1  g02134(.A0(new_n2183_), .A1(new_n2092_), .B0(new_n2198_), .Y(new_n2199_));
  XOR2X1   g02135(.A(new_n2137_), .B(new_n2092_), .Y(new_n2200_));
  XOR2X1   g02136(.A(new_n2200_), .B(new_n2199_), .Y(new_n2201_));
  INVX1    g02137(.A(new_n2201_), .Y(new_n2202_));
  OAI21X1  g02138(.A0(new_n2202_), .A1(new_n2063_), .B0(new_n2188_), .Y(new_n2203_));
  XOR2X1   g02139(.A(new_n2203_), .B(new_n74_), .Y(new_n2204_));
  OAI21X1  g02140(.A0(new_n2204_), .A1(new_n2059_), .B0(new_n2057_), .Y(new_n2205_));
  INVX1    g02141(.A(new_n1893_), .Y(new_n2206_));
  NOR2X1   g02142(.A(new_n1997_), .B(new_n1919_), .Y(new_n2207_));
  AOI21X1  g02143(.A0(new_n1998_), .A1(new_n2206_), .B0(new_n2207_), .Y(new_n2208_));
  OAI22X1  g02144(.A0(new_n152_), .A1(new_n78_), .B0(new_n99_), .B1(new_n84_), .Y(new_n2209_));
  OR4X1    g02145(.A(new_n2209_), .B(new_n1119_), .C(new_n814_), .D(new_n974_), .Y(new_n2210_));
  OR4X1    g02146(.A(new_n475_), .B(new_n260_), .C(new_n928_), .D(new_n80_), .Y(new_n2211_));
  OR4X1    g02147(.A(new_n2211_), .B(new_n612_), .C(new_n468_), .D(new_n579_), .Y(new_n2212_));
  OR4X1    g02148(.A(new_n2212_), .B(new_n2210_), .C(new_n2169_), .D(new_n1109_), .Y(new_n2213_));
  OR4X1    g02149(.A(new_n494_), .B(new_n232_), .C(new_n213_), .D(new_n191_), .Y(new_n2214_));
  OAI22X1  g02150(.A0(new_n123_), .A1(new_n108_), .B0(new_n105_), .B1(new_n84_), .Y(new_n2215_));
  OR4X1    g02151(.A(new_n2215_), .B(new_n1142_), .C(new_n393_), .D(new_n137_), .Y(new_n2216_));
  OR4X1    g02152(.A(new_n2216_), .B(new_n2214_), .C(new_n196_), .D(new_n884_), .Y(new_n2217_));
  OR4X1    g02153(.A(new_n938_), .B(new_n636_), .C(new_n282_), .D(new_n274_), .Y(new_n2218_));
  OR4X1    g02154(.A(new_n423_), .B(new_n746_), .C(new_n111_), .D(new_n1046_), .Y(new_n2219_));
  OR4X1    g02155(.A(new_n2219_), .B(new_n2218_), .C(new_n370_), .D(new_n173_), .Y(new_n2220_));
  AOI21X1  g02156(.A0(new_n129_), .A1(new_n125_), .B0(new_n88_), .Y(new_n2221_));
  OR4X1    g02157(.A(new_n2221_), .B(new_n417_), .C(new_n439_), .D(new_n390_), .Y(new_n2222_));
  OR4X1    g02158(.A(new_n2222_), .B(new_n394_), .C(new_n361_), .D(new_n358_), .Y(new_n2223_));
  OR4X1    g02159(.A(new_n2223_), .B(new_n2220_), .C(new_n2217_), .D(new_n1693_), .Y(new_n2224_));
  OR2X1    g02160(.A(new_n2224_), .B(new_n2213_), .Y(new_n2225_));
  NOR4X1   g02161(.A(new_n478_), .B(new_n255_), .C(new_n291_), .D(new_n651_), .Y(new_n2226_));
  INVX1    g02162(.A(new_n2226_), .Y(new_n2227_));
  OR4X1    g02163(.A(new_n399_), .B(new_n208_), .C(new_n303_), .D(new_n981_), .Y(new_n2228_));
  OR4X1    g02164(.A(new_n2228_), .B(new_n543_), .C(new_n504_), .D(new_n329_), .Y(new_n2229_));
  OR4X1    g02165(.A(new_n2229_), .B(new_n1385_), .C(new_n1105_), .D(new_n896_), .Y(new_n2230_));
  NOR2X1   g02166(.A(new_n848_), .B(new_n432_), .Y(new_n2231_));
  NOR4X1   g02167(.A(new_n1261_), .B(new_n365_), .C(new_n420_), .D(new_n144_), .Y(new_n2232_));
  NOR3X1   g02168(.A(new_n710_), .B(new_n449_), .C(new_n338_), .Y(new_n2233_));
  NOR3X1   g02169(.A(new_n1100_), .B(new_n1082_), .C(new_n850_), .Y(new_n2234_));
  NAND4X1  g02170(.A(new_n2234_), .B(new_n2233_), .C(new_n2232_), .D(new_n2231_), .Y(new_n2235_));
  OR4X1    g02171(.A(new_n2235_), .B(new_n2230_), .C(new_n2227_), .D(new_n1039_), .Y(new_n2236_));
  NOR2X1   g02172(.A(new_n2236_), .B(new_n2225_), .Y(new_n2237_));
  NOR2X1   g02173(.A(new_n2237_), .B(new_n1919_), .Y(new_n2238_));
  AND2X1   g02174(.A(new_n2237_), .B(new_n1919_), .Y(new_n2239_));
  NOR3X1   g02175(.A(new_n2239_), .B(new_n2238_), .C(new_n2208_), .Y(new_n2240_));
  OR2X1    g02176(.A(new_n2240_), .B(new_n2239_), .Y(new_n2241_));
  OAI22X1  g02177(.A0(new_n2241_), .A1(new_n2238_), .B0(new_n2240_), .B1(new_n2208_), .Y(new_n2242_));
  XOR2X1   g02178(.A(new_n2194_), .B(new_n2192_), .Y(new_n2243_));
  INVX1    g02179(.A(new_n2243_), .Y(new_n2244_));
  INVX1    g02180(.A(new_n1890_), .Y(new_n2245_));
  INVX1    g02181(.A(new_n2183_), .Y(new_n2246_));
  AOI22X1  g02182(.A0(new_n2246_), .A1(new_n1889_), .B0(new_n1884_), .B1(new_n1887_), .Y(new_n2247_));
  OAI21X1  g02183(.A0(new_n2245_), .A1(new_n520_), .B0(new_n2247_), .Y(new_n2248_));
  AOI21X1  g02184(.A0(new_n2244_), .A1(new_n407_), .B0(new_n2248_), .Y(new_n2249_));
  XOR2X1   g02185(.A(new_n2249_), .B(new_n2242_), .Y(new_n2250_));
  XOR2X1   g02186(.A(new_n2250_), .B(new_n2205_), .Y(new_n2251_));
  INVX1    g02187(.A(new_n2137_), .Y(new_n2252_));
  OR4X1    g02188(.A(new_n395_), .B(new_n474_), .C(new_n190_), .D(new_n177_), .Y(new_n2253_));
  NOR2X1   g02189(.A(new_n2253_), .B(new_n801_), .Y(new_n2254_));
  OR4X1    g02190(.A(new_n285_), .B(new_n180_), .C(new_n159_), .D(new_n158_), .Y(new_n2255_));
  OR4X1    g02191(.A(new_n2255_), .B(new_n1316_), .C(new_n843_), .D(new_n139_), .Y(new_n2256_));
  NOR4X1   g02192(.A(new_n2256_), .B(new_n741_), .C(new_n412_), .D(new_n274_), .Y(new_n2257_));
  OR4X1    g02193(.A(new_n720_), .B(new_n596_), .C(new_n361_), .D(new_n126_), .Y(new_n2258_));
  OR4X1    g02194(.A(new_n2258_), .B(new_n229_), .C(new_n648_), .D(new_n104_), .Y(new_n2259_));
  OR4X1    g02195(.A(new_n372_), .B(new_n423_), .C(new_n203_), .D(new_n144_), .Y(new_n2260_));
  OR4X1    g02196(.A(new_n2260_), .B(new_n740_), .C(new_n426_), .D(new_n120_), .Y(new_n2261_));
  OR4X1    g02197(.A(new_n2157_), .B(new_n1114_), .C(new_n947_), .D(new_n714_), .Y(new_n2262_));
  NOR3X1   g02198(.A(new_n2262_), .B(new_n2261_), .C(new_n2259_), .Y(new_n2263_));
  NAND3X1  g02199(.A(new_n2263_), .B(new_n2257_), .C(new_n2254_), .Y(new_n2264_));
  INVX1    g02200(.A(new_n1636_), .Y(new_n2265_));
  OR2X1    g02201(.A(new_n891_), .B(new_n147_), .Y(new_n2266_));
  OR4X1    g02202(.A(new_n589_), .B(new_n478_), .C(new_n251_), .D(new_n449_), .Y(new_n2267_));
  OR4X1    g02203(.A(new_n2267_), .B(new_n2266_), .C(new_n504_), .D(new_n300_), .Y(new_n2268_));
  OR4X1    g02204(.A(new_n681_), .B(new_n228_), .C(new_n522_), .D(new_n337_), .Y(new_n2269_));
  OR4X1    g02205(.A(new_n2269_), .B(new_n505_), .C(new_n459_), .D(new_n806_), .Y(new_n2270_));
  OR4X1    g02206(.A(new_n2270_), .B(new_n1320_), .C(new_n842_), .D(new_n1087_), .Y(new_n2271_));
  OR4X1    g02207(.A(new_n694_), .B(new_n358_), .C(new_n850_), .D(new_n232_), .Y(new_n2272_));
  OR4X1    g02208(.A(new_n2272_), .B(new_n2271_), .C(new_n2268_), .D(new_n2265_), .Y(new_n2273_));
  OAI22X1  g02209(.A0(new_n125_), .A1(new_n102_), .B0(new_n84_), .B1(new_n81_), .Y(new_n2274_));
  OR2X1    g02210(.A(new_n2274_), .B(new_n747_), .Y(new_n2275_));
  OR4X1    g02211(.A(new_n541_), .B(new_n496_), .C(new_n246_), .D(new_n202_), .Y(new_n2276_));
  OR4X1    g02212(.A(new_n2276_), .B(new_n2275_), .C(new_n823_), .D(new_n566_), .Y(new_n2277_));
  OR4X1    g02213(.A(new_n2277_), .B(new_n1909_), .C(new_n1757_), .D(new_n1608_), .Y(new_n2278_));
  AOI21X1  g02214(.A0(new_n161_), .A1(new_n94_), .B0(new_n96_), .Y(new_n2279_));
  OR4X1    g02215(.A(new_n357_), .B(new_n410_), .C(new_n155_), .D(new_n134_), .Y(new_n2280_));
  OR4X1    g02216(.A(new_n2280_), .B(new_n2279_), .C(new_n1558_), .D(new_n1044_), .Y(new_n2281_));
  INVX1    g02217(.A(new_n586_), .Y(new_n2282_));
  NAND3X1  g02218(.A(new_n719_), .B(new_n2282_), .C(new_n171_), .Y(new_n2283_));
  OR4X1    g02219(.A(new_n245_), .B(new_n231_), .C(new_n114_), .D(new_n1579_), .Y(new_n2284_));
  OR4X1    g02220(.A(new_n2284_), .B(new_n2283_), .C(new_n1205_), .D(new_n1096_), .Y(new_n2285_));
  OR4X1    g02221(.A(new_n2285_), .B(new_n2281_), .C(new_n2278_), .D(new_n2273_), .Y(new_n2286_));
  NOR2X1   g02222(.A(new_n2286_), .B(new_n2264_), .Y(new_n2287_));
  OAI22X1  g02223(.A0(new_n2287_), .A1(new_n2140_), .B0(new_n2186_), .B1(new_n2092_), .Y(new_n2288_));
  AOI21X1  g02224(.A0(new_n2252_), .A1(new_n2095_), .B0(new_n2288_), .Y(new_n2289_));
  NOR2X1   g02225(.A(new_n2137_), .B(new_n2092_), .Y(new_n2290_));
  AOI21X1  g02226(.A0(new_n2200_), .A1(new_n2199_), .B0(new_n2290_), .Y(new_n2291_));
  XOR2X1   g02227(.A(new_n2287_), .B(new_n2137_), .Y(new_n2292_));
  INVX1    g02228(.A(new_n2292_), .Y(new_n2293_));
  XOR2X1   g02229(.A(new_n2293_), .B(new_n2291_), .Y(new_n2294_));
  INVX1    g02230(.A(new_n2294_), .Y(new_n2295_));
  OAI21X1  g02231(.A0(new_n2295_), .A1(new_n2063_), .B0(new_n2289_), .Y(new_n2296_));
  XOR2X1   g02232(.A(new_n2296_), .B(new_n74_), .Y(new_n2297_));
  XOR2X1   g02233(.A(new_n2297_), .B(new_n2251_), .Y(new_n2298_));
  XOR2X1   g02234(.A(\a[24] ), .B(new_n70_), .Y(new_n2299_));
  XOR2X1   g02235(.A(\a[26] ), .B(new_n77_), .Y(new_n2300_));
  NOR2X1   g02236(.A(new_n2300_), .B(new_n2299_), .Y(new_n2301_));
  OAI22X1  g02237(.A0(new_n131_), .A1(new_n79_), .B0(new_n105_), .B1(new_n96_), .Y(new_n2302_));
  OR4X1    g02238(.A(new_n2302_), .B(new_n1609_), .C(new_n459_), .D(new_n133_), .Y(new_n2303_));
  OAI22X1  g02239(.A0(new_n182_), .A1(new_n123_), .B0(new_n106_), .B1(new_n81_), .Y(new_n2304_));
  OR4X1    g02240(.A(new_n2304_), .B(new_n1306_), .C(new_n1156_), .D(new_n312_), .Y(new_n2305_));
  OR4X1    g02241(.A(new_n642_), .B(new_n1044_), .C(new_n408_), .D(new_n382_), .Y(new_n2306_));
  OR4X1    g02242(.A(new_n840_), .B(new_n193_), .C(new_n134_), .D(new_n338_), .Y(new_n2307_));
  NOR4X1   g02243(.A(new_n2307_), .B(new_n2306_), .C(new_n2305_), .D(new_n2303_), .Y(new_n2308_));
  AOI21X1  g02244(.A0(new_n148_), .A1(new_n123_), .B0(new_n105_), .Y(new_n2309_));
  OR4X1    g02245(.A(new_n2309_), .B(new_n300_), .C(new_n243_), .D(new_n337_), .Y(new_n2310_));
  OR4X1    g02246(.A(new_n358_), .B(new_n285_), .C(new_n280_), .D(new_n194_), .Y(new_n2311_));
  OR4X1    g02247(.A(new_n355_), .B(new_n292_), .C(new_n535_), .D(new_n585_), .Y(new_n2312_));
  NOR4X1   g02248(.A(new_n2312_), .B(new_n2311_), .C(new_n2310_), .D(new_n1273_), .Y(new_n2313_));
  OR4X1    g02249(.A(new_n536_), .B(new_n191_), .C(new_n825_), .D(new_n928_), .Y(new_n2314_));
  OR4X1    g02250(.A(new_n2314_), .B(new_n1028_), .C(new_n265_), .D(new_n398_), .Y(new_n2315_));
  NOR3X1   g02251(.A(new_n2315_), .B(new_n767_), .C(new_n208_), .Y(new_n2316_));
  OR4X1    g02252(.A(new_n580_), .B(new_n509_), .C(new_n506_), .D(new_n372_), .Y(new_n2317_));
  NOR3X1   g02253(.A(new_n2317_), .B(new_n873_), .C(new_n694_), .Y(new_n2318_));
  NAND4X1  g02254(.A(new_n2318_), .B(new_n2316_), .C(new_n2313_), .D(new_n2308_), .Y(new_n2319_));
  INVX1    g02255(.A(new_n426_), .Y(new_n2320_));
  NAND3X1  g02256(.A(new_n1570_), .B(new_n2320_), .C(new_n344_), .Y(new_n2321_));
  OR4X1    g02257(.A(new_n2101_), .B(new_n1061_), .C(new_n256_), .D(new_n228_), .Y(new_n2322_));
  AOI21X1  g02258(.A0(new_n143_), .A1(new_n131_), .B0(new_n119_), .Y(new_n2323_));
  OR2X1    g02259(.A(new_n2323_), .B(new_n274_), .Y(new_n2324_));
  NOR4X1   g02260(.A(new_n2324_), .B(new_n2322_), .C(new_n2321_), .D(new_n1079_), .Y(new_n2325_));
  INVX1    g02261(.A(new_n2325_), .Y(new_n2326_));
  OR4X1    g02262(.A(new_n187_), .B(new_n291_), .C(new_n431_), .D(new_n111_), .Y(new_n2327_));
  OR4X1    g02263(.A(new_n399_), .B(new_n220_), .C(new_n183_), .D(new_n1008_), .Y(new_n2328_));
  OAI22X1  g02264(.A0(new_n108_), .A1(new_n102_), .B0(new_n99_), .B1(new_n91_), .Y(new_n2329_));
  OR2X1    g02265(.A(new_n2329_), .B(new_n505_), .Y(new_n2330_));
  OR4X1    g02266(.A(new_n2330_), .B(new_n2328_), .C(new_n2327_), .D(new_n1717_), .Y(new_n2331_));
  OR4X1    g02267(.A(new_n1757_), .B(new_n921_), .C(new_n301_), .D(new_n200_), .Y(new_n2332_));
  OR4X1    g02268(.A(new_n213_), .B(new_n648_), .C(new_n746_), .D(new_n103_), .Y(new_n2333_));
  OR2X1    g02269(.A(new_n714_), .B(new_n582_), .Y(new_n2334_));
  OR4X1    g02270(.A(new_n393_), .B(new_n391_), .C(new_n371_), .D(new_n400_), .Y(new_n2335_));
  OR4X1    g02271(.A(new_n540_), .B(new_n365_), .C(new_n350_), .D(new_n259_), .Y(new_n2336_));
  OR4X1    g02272(.A(new_n2336_), .B(new_n2335_), .C(new_n2334_), .D(new_n2333_), .Y(new_n2337_));
  OR4X1    g02273(.A(new_n2337_), .B(new_n2332_), .C(new_n2331_), .D(new_n2326_), .Y(new_n2338_));
  NOR2X1   g02274(.A(new_n2338_), .B(new_n2319_), .Y(new_n2339_));
  AOI21X1  g02275(.A0(new_n161_), .A1(new_n81_), .B0(new_n106_), .Y(new_n2340_));
  OR4X1    g02276(.A(new_n259_), .B(new_n184_), .C(new_n178_), .D(new_n177_), .Y(new_n2341_));
  OAI22X1  g02277(.A0(new_n119_), .A1(new_n81_), .B0(new_n106_), .B1(new_n92_), .Y(new_n2342_));
  OR4X1    g02278(.A(new_n2342_), .B(new_n1921_), .C(new_n429_), .D(new_n396_), .Y(new_n2343_));
  NOR4X1   g02279(.A(new_n2343_), .B(new_n2341_), .C(new_n2340_), .D(new_n2328_), .Y(new_n2344_));
  NAND3X1  g02280(.A(new_n2344_), .B(new_n2325_), .C(new_n2316_), .Y(new_n2345_));
  OR4X1    g02281(.A(new_n679_), .B(new_n226_), .C(new_n201_), .D(new_n379_), .Y(new_n2346_));
  OR2X1    g02282(.A(new_n1438_), .B(new_n1090_), .Y(new_n2347_));
  NOR4X1   g02283(.A(new_n2347_), .B(new_n2346_), .C(new_n1756_), .D(new_n1721_), .Y(new_n2348_));
  INVX1    g02284(.A(new_n2348_), .Y(new_n2349_));
  OR4X1    g02285(.A(new_n500_), .B(new_n480_), .C(new_n423_), .D(new_n156_), .Y(new_n2350_));
  OR4X1    g02286(.A(new_n1386_), .B(new_n374_), .C(new_n246_), .D(new_n126_), .Y(new_n2351_));
  OR2X1    g02287(.A(new_n2351_), .B(new_n2350_), .Y(new_n2352_));
  NOR3X1   g02288(.A(new_n314_), .B(new_n180_), .C(new_n610_), .Y(new_n2353_));
  NOR4X1   g02289(.A(new_n843_), .B(new_n282_), .C(new_n247_), .D(new_n234_), .Y(new_n2354_));
  NAND2X1  g02290(.A(new_n2354_), .B(new_n2353_), .Y(new_n2355_));
  OR4X1    g02291(.A(new_n540_), .B(new_n400_), .C(new_n218_), .D(new_n116_), .Y(new_n2356_));
  OR4X1    g02292(.A(new_n2356_), .B(new_n2355_), .C(new_n2352_), .D(new_n566_), .Y(new_n2357_));
  OR4X1    g02293(.A(new_n504_), .B(new_n412_), .C(new_n354_), .D(new_n100_), .Y(new_n2358_));
  OR4X1    g02294(.A(new_n2358_), .B(new_n1320_), .C(new_n560_), .D(new_n233_), .Y(new_n2359_));
  OR4X1    g02295(.A(new_n2359_), .B(new_n2357_), .C(new_n2349_), .D(new_n2096_), .Y(new_n2360_));
  AOI21X1  g02296(.A0(new_n161_), .A1(new_n78_), .B0(new_n168_), .Y(new_n2361_));
  NOR4X1   g02297(.A(new_n2361_), .B(new_n1663_), .C(new_n1274_), .D(new_n723_), .Y(new_n2362_));
  NAND2X1  g02298(.A(new_n2362_), .B(new_n1164_), .Y(new_n2363_));
  OR2X1    g02299(.A(new_n206_), .B(new_n199_), .Y(new_n2364_));
  OR4X1    g02300(.A(new_n2364_), .B(new_n2363_), .C(new_n2360_), .D(new_n2345_), .Y(new_n2365_));
  OR4X1    g02301(.A(new_n1703_), .B(new_n444_), .C(new_n286_), .D(new_n276_), .Y(new_n2366_));
  OR2X1    g02302(.A(new_n2366_), .B(new_n1528_), .Y(new_n2367_));
  OR2X1    g02303(.A(new_n815_), .B(new_n433_), .Y(new_n2368_));
  OR4X1    g02304(.A(new_n1623_), .B(new_n676_), .C(new_n301_), .D(new_n200_), .Y(new_n2369_));
  OR4X1    g02305(.A(new_n2369_), .B(new_n2368_), .C(new_n2367_), .D(new_n2285_), .Y(new_n2370_));
  OR4X1    g02306(.A(new_n386_), .B(new_n565_), .C(new_n757_), .D(new_n137_), .Y(new_n2371_));
  OR4X1    g02307(.A(new_n2371_), .B(new_n691_), .C(new_n207_), .D(new_n664_), .Y(new_n2372_));
  OR4X1    g02308(.A(new_n2372_), .B(new_n417_), .C(new_n329_), .D(new_n299_), .Y(new_n2373_));
  AOI21X1  g02309(.A0(new_n182_), .A1(new_n105_), .B0(new_n123_), .Y(new_n2374_));
  NOR4X1   g02310(.A(new_n2374_), .B(new_n755_), .C(new_n631_), .D(new_n285_), .Y(new_n2375_));
  INVX1    g02311(.A(new_n2375_), .Y(new_n2376_));
  OR4X1    g02312(.A(new_n2376_), .B(new_n2373_), .C(new_n537_), .D(new_n307_), .Y(new_n2377_));
  OR2X1    g02313(.A(new_n2377_), .B(new_n2370_), .Y(new_n2378_));
  NOR2X1   g02314(.A(new_n2378_), .B(new_n2365_), .Y(new_n2379_));
  NOR2X1   g02315(.A(new_n2339_), .B(new_n2287_), .Y(new_n2380_));
  OR2X1    g02316(.A(new_n2293_), .B(new_n2291_), .Y(new_n2381_));
  OAI21X1  g02317(.A0(new_n2287_), .A1(new_n2137_), .B0(new_n2381_), .Y(new_n2382_));
  XOR2X1   g02318(.A(new_n2339_), .B(new_n2287_), .Y(new_n2383_));
  AOI21X1  g02319(.A0(new_n2383_), .A1(new_n2382_), .B0(new_n2380_), .Y(new_n2384_));
  XOR2X1   g02320(.A(new_n2379_), .B(new_n2339_), .Y(new_n2385_));
  INVX1    g02321(.A(new_n2385_), .Y(new_n2386_));
  OR2X1    g02322(.A(new_n2386_), .B(new_n2384_), .Y(new_n2387_));
  OAI21X1  g02323(.A0(new_n2379_), .A1(new_n2339_), .B0(new_n2387_), .Y(new_n2388_));
  NOR3X1   g02324(.A(new_n1134_), .B(new_n743_), .C(new_n537_), .Y(new_n2389_));
  NOR4X1   g02325(.A(new_n496_), .B(new_n348_), .C(new_n329_), .D(new_n664_), .Y(new_n2390_));
  NOR3X1   g02326(.A(new_n271_), .B(new_n133_), .C(new_n1579_), .Y(new_n2391_));
  NAND3X1  g02327(.A(new_n2391_), .B(new_n2390_), .C(new_n2389_), .Y(new_n2392_));
  AOI21X1  g02328(.A0(new_n143_), .A1(new_n81_), .B0(new_n79_), .Y(new_n2393_));
  OR4X1    g02329(.A(new_n2393_), .B(new_n2392_), .C(new_n2367_), .D(new_n1513_), .Y(new_n2394_));
  OR2X1    g02330(.A(new_n108_), .B(new_n91_), .Y(new_n2395_));
  INVX1    g02331(.A(new_n814_), .Y(new_n2396_));
  OR2X1    g02332(.A(new_n647_), .B(new_n441_), .Y(new_n2397_));
  AOI21X1  g02333(.A0(new_n99_), .A1(new_n92_), .B0(new_n69_), .Y(new_n2398_));
  OR4X1    g02334(.A(new_n2398_), .B(new_n547_), .C(new_n332_), .D(new_n209_), .Y(new_n2399_));
  NOR4X1   g02335(.A(new_n2399_), .B(new_n2397_), .C(new_n1984_), .D(new_n1848_), .Y(new_n2400_));
  NOR4X1   g02336(.A(new_n478_), .B(new_n474_), .C(new_n251_), .D(new_n521_), .Y(new_n2401_));
  NAND4X1  g02337(.A(new_n2401_), .B(new_n2400_), .C(new_n2396_), .D(new_n2395_), .Y(new_n2402_));
  OR4X1    g02338(.A(new_n2066_), .B(new_n1158_), .C(new_n891_), .D(new_n391_), .Y(new_n2403_));
  NOR3X1   g02339(.A(new_n2403_), .B(new_n2402_), .C(new_n2394_), .Y(new_n2404_));
  INVX1    g02340(.A(new_n2404_), .Y(new_n2405_));
  AOI21X1  g02341(.A0(new_n129_), .A1(new_n99_), .B0(new_n123_), .Y(new_n2406_));
  OR4X1    g02342(.A(new_n2406_), .B(new_n232_), .C(new_n187_), .D(new_n111_), .Y(new_n2407_));
  OR2X1    g02343(.A(new_n2407_), .B(new_n2125_), .Y(new_n2408_));
  AOI21X1  g02344(.A0(new_n182_), .A1(new_n78_), .B0(new_n102_), .Y(new_n2409_));
  OR4X1    g02345(.A(new_n2409_), .B(new_n641_), .C(new_n365_), .D(new_n233_), .Y(new_n2410_));
  OR4X1    g02346(.A(new_n802_), .B(new_n427_), .C(new_n400_), .D(new_n206_), .Y(new_n2411_));
  NOR3X1   g02347(.A(new_n2411_), .B(new_n2410_), .C(new_n2408_), .Y(new_n2412_));
  INVX1    g02348(.A(new_n2412_), .Y(new_n2413_));
  NOR4X1   g02349(.A(new_n2413_), .B(new_n2405_), .C(new_n510_), .D(new_n460_), .Y(new_n2414_));
  XOR2X1   g02350(.A(new_n2414_), .B(new_n2379_), .Y(new_n2415_));
  XOR2X1   g02351(.A(new_n2415_), .B(new_n2388_), .Y(new_n2416_));
  XOR2X1   g02352(.A(\a[25] ), .B(\a[24] ), .Y(new_n2417_));
  AND2X1   g02353(.A(new_n2417_), .B(new_n2299_), .Y(new_n2418_));
  INVX1    g02354(.A(new_n2418_), .Y(new_n2419_));
  INVX1    g02355(.A(new_n2339_), .Y(new_n2420_));
  INVX1    g02356(.A(new_n2414_), .Y(new_n2421_));
  INVX1    g02357(.A(new_n2299_), .Y(new_n2422_));
  AND2X1   g02358(.A(new_n2300_), .B(new_n2422_), .Y(new_n2423_));
  NOR3X1   g02359(.A(new_n2417_), .B(new_n2300_), .C(new_n2422_), .Y(new_n2424_));
  AOI22X1  g02360(.A0(new_n2424_), .A1(new_n2420_), .B0(new_n2423_), .B1(new_n2421_), .Y(new_n2425_));
  OAI21X1  g02361(.A0(new_n2419_), .A1(new_n2379_), .B0(new_n2425_), .Y(new_n2426_));
  AOI21X1  g02362(.A0(new_n2416_), .A1(new_n2301_), .B0(new_n2426_), .Y(new_n2427_));
  XOR2X1   g02363(.A(new_n2427_), .B(\a[26] ), .Y(new_n2428_));
  XOR2X1   g02364(.A(new_n2428_), .B(new_n2298_), .Y(new_n2429_));
  XOR2X1   g02365(.A(new_n2197_), .B(new_n2195_), .Y(new_n2430_));
  INVX1    g02366(.A(new_n2095_), .Y(new_n2431_));
  AOI22X1  g02367(.A0(new_n2185_), .A1(new_n1887_), .B0(new_n2139_), .B1(new_n2093_), .Y(new_n2432_));
  OAI21X1  g02368(.A0(new_n2183_), .A1(new_n2431_), .B0(new_n2432_), .Y(new_n2433_));
  AOI21X1  g02369(.A0(new_n2430_), .A1(new_n2062_), .B0(new_n2433_), .Y(new_n2434_));
  XOR2X1   g02370(.A(new_n2434_), .B(\a[29] ), .Y(new_n2435_));
  XOR2X1   g02371(.A(new_n2054_), .B(new_n2052_), .Y(new_n2436_));
  NOR2X1   g02372(.A(new_n2436_), .B(new_n2435_), .Y(new_n2437_));
  INVX1    g02373(.A(new_n2437_), .Y(new_n2438_));
  XOR2X1   g02374(.A(new_n2436_), .B(new_n2435_), .Y(new_n2439_));
  INVX1    g02375(.A(new_n2439_), .Y(new_n2440_));
  INVX1    g02376(.A(new_n2040_), .Y(new_n2441_));
  NOR2X1   g02377(.A(new_n2041_), .B(new_n2039_), .Y(new_n2442_));
  AOI21X1  g02378(.A0(new_n2042_), .A1(new_n2441_), .B0(new_n2442_), .Y(new_n2443_));
  INVX1    g02379(.A(new_n1948_), .Y(new_n2444_));
  INVX1    g02380(.A(\a[17] ), .Y(new_n2445_));
  INVX1    g02381(.A(new_n2308_), .Y(new_n2446_));
  NOR4X1   g02382(.A(new_n777_), .B(new_n569_), .C(new_n484_), .D(new_n272_), .Y(new_n2447_));
  NOR4X1   g02383(.A(new_n412_), .B(new_n282_), .C(new_n259_), .D(new_n792_), .Y(new_n2448_));
  NOR4X1   g02384(.A(new_n546_), .B(new_n245_), .C(new_n218_), .D(new_n181_), .Y(new_n2449_));
  AOI21X1  g02385(.A0(new_n131_), .A1(new_n125_), .B0(new_n69_), .Y(new_n2450_));
  OAI22X1  g02386(.A0(new_n168_), .A1(new_n72_), .B0(new_n131_), .B1(new_n115_), .Y(new_n2451_));
  OR4X1    g02387(.A(new_n2451_), .B(new_n1514_), .C(new_n2450_), .D(new_n827_), .Y(new_n2452_));
  NOR2X1   g02388(.A(new_n2452_), .B(new_n1863_), .Y(new_n2453_));
  NAND4X1  g02389(.A(new_n2453_), .B(new_n2449_), .C(new_n2448_), .D(new_n2447_), .Y(new_n2454_));
  OR4X1    g02390(.A(new_n2454_), .B(new_n2446_), .C(new_n1629_), .D(new_n1533_), .Y(new_n2455_));
  NOR3X1   g02391(.A(new_n2455_), .B(new_n2120_), .C(new_n2113_), .Y(new_n2456_));
  OR4X1    g02392(.A(new_n589_), .B(new_n1166_), .C(new_n968_), .D(new_n224_), .Y(new_n2457_));
  OR4X1    g02393(.A(new_n245_), .B(new_n226_), .C(new_n177_), .D(new_n156_), .Y(new_n2458_));
  OR4X1    g02394(.A(new_n543_), .B(new_n422_), .C(new_n246_), .D(new_n381_), .Y(new_n2459_));
  OR4X1    g02395(.A(new_n2459_), .B(new_n2458_), .C(new_n2457_), .D(new_n897_), .Y(new_n2460_));
  OR4X1    g02396(.A(new_n1255_), .B(new_n947_), .C(new_n1443_), .D(new_n602_), .Y(new_n2461_));
  OR2X1    g02397(.A(new_n2461_), .B(new_n1011_), .Y(new_n2462_));
  OR4X1    g02398(.A(new_n848_), .B(new_n414_), .C(new_n350_), .D(new_n300_), .Y(new_n2463_));
  OR4X1    g02399(.A(new_n2463_), .B(new_n935_), .C(new_n173_), .D(new_n172_), .Y(new_n2464_));
  OR4X1    g02400(.A(new_n1336_), .B(new_n945_), .C(new_n627_), .D(new_n183_), .Y(new_n2465_));
  OR4X1    g02401(.A(new_n2465_), .B(new_n2464_), .C(new_n2462_), .D(new_n2460_), .Y(new_n2466_));
  OR4X1    g02402(.A(new_n523_), .B(new_n387_), .C(new_n265_), .D(new_n1087_), .Y(new_n2467_));
  OR4X1    g02403(.A(new_n251_), .B(new_n194_), .C(new_n147_), .D(new_n981_), .Y(new_n2468_));
  OR4X1    g02404(.A(new_n497_), .B(new_n496_), .C(new_n307_), .D(new_n337_), .Y(new_n2469_));
  OR4X1    g02405(.A(new_n2469_), .B(new_n2468_), .C(new_n2467_), .D(new_n477_), .Y(new_n2470_));
  OR4X1    g02406(.A(new_n1550_), .B(new_n882_), .C(new_n421_), .D(new_n299_), .Y(new_n2471_));
  OR4X1    g02407(.A(new_n181_), .B(new_n792_), .C(new_n610_), .D(new_n138_), .Y(new_n2472_));
  OR4X1    g02408(.A(new_n2472_), .B(new_n772_), .C(new_n365_), .D(new_n233_), .Y(new_n2473_));
  OR4X1    g02409(.A(new_n2473_), .B(new_n2471_), .C(new_n2470_), .D(new_n2096_), .Y(new_n2474_));
  NOR3X1   g02410(.A(new_n2474_), .B(new_n2466_), .C(new_n2156_), .Y(new_n2475_));
  NOR2X1   g02411(.A(new_n2475_), .B(new_n2456_), .Y(new_n2476_));
  NAND2X1  g02412(.A(new_n2475_), .B(new_n2456_), .Y(new_n2477_));
  AOI21X1  g02413(.A0(new_n2477_), .A1(new_n2445_), .B0(new_n2476_), .Y(new_n2478_));
  NOR2X1   g02414(.A(new_n2478_), .B(new_n2444_), .Y(new_n2479_));
  XOR2X1   g02415(.A(new_n1838_), .B(new_n1837_), .Y(new_n2480_));
  INVX1    g02416(.A(new_n847_), .Y(new_n2481_));
  AOI22X1  g02417(.A0(new_n1890_), .A1(new_n2481_), .B0(new_n1889_), .B1(new_n2049_), .Y(new_n2482_));
  OAI21X1  g02418(.A0(new_n1885_), .A1(new_n783_), .B0(new_n2482_), .Y(new_n2483_));
  AOI21X1  g02419(.A0(new_n2480_), .A1(new_n407_), .B0(new_n2483_), .Y(new_n2484_));
  INVX1    g02420(.A(new_n2484_), .Y(new_n2485_));
  XOR2X1   g02421(.A(new_n2478_), .B(new_n2444_), .Y(new_n2486_));
  AOI21X1  g02422(.A0(new_n2486_), .A1(new_n2485_), .B0(new_n2479_), .Y(new_n2487_));
  NOR2X1   g02423(.A(new_n2487_), .B(new_n2443_), .Y(new_n2488_));
  XOR2X1   g02424(.A(new_n2487_), .B(new_n2443_), .Y(new_n2489_));
  XOR2X1   g02425(.A(new_n2486_), .B(new_n2484_), .Y(new_n2490_));
  NOR2X1   g02426(.A(new_n2476_), .B(\a[17] ), .Y(new_n2491_));
  AOI21X1  g02427(.A0(new_n2491_), .A1(new_n2477_), .B0(\a[17] ), .Y(new_n2492_));
  AOI21X1  g02428(.A0(new_n2478_), .A1(new_n2477_), .B0(new_n2492_), .Y(new_n2493_));
  XOR2X1   g02429(.A(new_n1835_), .B(new_n1834_), .Y(new_n2494_));
  AOI22X1  g02430(.A0(new_n1889_), .A1(new_n2036_), .B0(new_n1884_), .B1(new_n2481_), .Y(new_n2495_));
  OAI21X1  g02431(.A0(new_n2245_), .A1(new_n903_), .B0(new_n2495_), .Y(new_n2496_));
  AOI21X1  g02432(.A0(new_n2494_), .A1(new_n407_), .B0(new_n2496_), .Y(new_n2497_));
  NOR2X1   g02433(.A(new_n2497_), .B(new_n2493_), .Y(new_n2498_));
  INVX1    g02434(.A(new_n1561_), .Y(new_n2499_));
  OAI22X1  g02435(.A0(new_n127_), .A1(new_n119_), .B0(new_n94_), .B1(new_n75_), .Y(new_n2500_));
  OR2X1    g02436(.A(new_n2500_), .B(new_n1087_), .Y(new_n2501_));
  OR4X1    g02437(.A(new_n480_), .B(new_n229_), .C(new_n191_), .D(new_n114_), .Y(new_n2502_));
  OAI22X1  g02438(.A0(new_n131_), .A1(new_n96_), .B0(new_n105_), .B1(new_n91_), .Y(new_n2503_));
  OR2X1    g02439(.A(new_n2503_), .B(new_n398_), .Y(new_n2504_));
  OR4X1    g02440(.A(new_n2504_), .B(new_n2502_), .C(new_n2501_), .D(new_n1934_), .Y(new_n2505_));
  OAI22X1  g02441(.A0(new_n152_), .A1(new_n94_), .B0(new_n123_), .B1(new_n92_), .Y(new_n2506_));
  OR4X1    g02442(.A(new_n2506_), .B(new_n786_), .C(new_n751_), .D(new_n607_), .Y(new_n2507_));
  OR2X1    g02443(.A(new_n2507_), .B(new_n1437_), .Y(new_n2508_));
  OR4X1    g02444(.A(new_n2508_), .B(new_n2505_), .C(new_n2499_), .D(new_n1520_), .Y(new_n2509_));
  OR4X1    g02445(.A(new_n393_), .B(new_n479_), .C(new_n199_), .D(new_n303_), .Y(new_n2510_));
  OR4X1    g02446(.A(new_n2510_), .B(new_n1640_), .C(new_n1502_), .D(new_n567_), .Y(new_n2511_));
  NOR3X1   g02447(.A(new_n523_), .B(new_n412_), .C(new_n329_), .Y(new_n2512_));
  NOR4X1   g02448(.A(new_n724_), .B(new_n634_), .C(new_n527_), .D(new_n387_), .Y(new_n2513_));
  NOR4X1   g02449(.A(new_n328_), .B(new_n819_), .C(new_n194_), .D(new_n173_), .Y(new_n2514_));
  NAND3X1  g02450(.A(new_n2514_), .B(new_n2513_), .C(new_n2512_), .Y(new_n2515_));
  OR4X1    g02451(.A(new_n2515_), .B(new_n2511_), .C(new_n1715_), .D(new_n1581_), .Y(new_n2516_));
  NOR3X1   g02452(.A(new_n391_), .B(new_n158_), .C(new_n80_), .Y(new_n2517_));
  NOR3X1   g02453(.A(new_n1538_), .B(new_n132_), .C(new_n93_), .Y(new_n2518_));
  NAND3X1  g02454(.A(new_n2518_), .B(new_n2517_), .C(new_n1630_), .Y(new_n2519_));
  OR4X1    g02455(.A(new_n755_), .B(new_n243_), .C(new_n224_), .D(new_n223_), .Y(new_n2520_));
  OR4X1    g02456(.A(new_n370_), .B(new_n285_), .C(new_n439_), .D(new_n206_), .Y(new_n2521_));
  OR4X1    g02457(.A(new_n578_), .B(new_n758_), .C(new_n177_), .D(new_n120_), .Y(new_n2522_));
  OR2X1    g02458(.A(new_n2522_), .B(new_n2521_), .Y(new_n2523_));
  OR4X1    g02459(.A(new_n2406_), .B(new_n1757_), .C(new_n769_), .D(new_n432_), .Y(new_n2524_));
  OR4X1    g02460(.A(new_n2524_), .B(new_n2523_), .C(new_n2520_), .D(new_n1409_), .Y(new_n2525_));
  NOR4X1   g02461(.A(new_n2525_), .B(new_n2519_), .C(new_n2516_), .D(new_n2509_), .Y(new_n2526_));
  OR4X1    g02462(.A(new_n2526_), .B(new_n2455_), .C(new_n2120_), .D(new_n2113_), .Y(new_n2527_));
  INVX1    g02463(.A(new_n2526_), .Y(new_n2528_));
  INVX1    g02464(.A(\a[14] ), .Y(new_n2529_));
  OAI22X1  g02465(.A0(new_n152_), .A1(new_n108_), .B0(new_n125_), .B1(new_n69_), .Y(new_n2530_));
  OR2X1    g02466(.A(new_n2530_), .B(new_n848_), .Y(new_n2531_));
  OR4X1    g02467(.A(new_n968_), .B(new_n421_), .C(new_n885_), .D(new_n292_), .Y(new_n2532_));
  OR4X1    g02468(.A(new_n2532_), .B(new_n2531_), .C(new_n1367_), .D(new_n347_), .Y(new_n2533_));
  OR4X1    g02469(.A(new_n892_), .B(new_n625_), .C(new_n162_), .D(new_n610_), .Y(new_n2534_));
  OR4X1    g02470(.A(new_n720_), .B(new_n631_), .C(new_n246_), .D(new_n522_), .Y(new_n2535_));
  AOI21X1  g02471(.A0(new_n119_), .A1(new_n115_), .B0(new_n90_), .Y(new_n2536_));
  OR4X1    g02472(.A(new_n2536_), .B(new_n2535_), .C(new_n371_), .D(new_n273_), .Y(new_n2537_));
  OR4X1    g02473(.A(new_n2537_), .B(new_n1384_), .C(new_n772_), .D(new_n1057_), .Y(new_n2538_));
  OR4X1    g02474(.A(new_n2538_), .B(new_n2534_), .C(new_n2533_), .D(new_n2519_), .Y(new_n2539_));
  OR4X1    g02475(.A(new_n678_), .B(new_n220_), .C(new_n206_), .D(new_n176_), .Y(new_n2540_));
  OR4X1    g02476(.A(new_n2540_), .B(new_n2504_), .C(new_n896_), .D(new_n382_), .Y(new_n2541_));
  OR4X1    g02477(.A(new_n423_), .B(new_n263_), .C(new_n177_), .D(new_n291_), .Y(new_n2542_));
  OAI22X1  g02478(.A0(new_n152_), .A1(new_n81_), .B0(new_n131_), .B1(new_n88_), .Y(new_n2543_));
  OR2X1    g02479(.A(new_n2543_), .B(new_n596_), .Y(new_n2544_));
  OR4X1    g02480(.A(new_n2544_), .B(new_n2542_), .C(new_n1751_), .D(new_n216_), .Y(new_n2545_));
  NOR4X1   g02481(.A(new_n2545_), .B(new_n2541_), .C(new_n2177_), .D(new_n1684_), .Y(new_n2546_));
  INVX1    g02482(.A(new_n2546_), .Y(new_n2547_));
  OR4X1    g02483(.A(new_n829_), .B(new_n234_), .C(new_n165_), .D(new_n100_), .Y(new_n2548_));
  OR4X1    g02484(.A(new_n387_), .B(new_n840_), .C(new_n717_), .D(new_n285_), .Y(new_n2549_));
  OR4X1    g02485(.A(new_n565_), .B(new_n187_), .C(new_n156_), .D(new_n137_), .Y(new_n2550_));
  OR4X1    g02486(.A(new_n2550_), .B(new_n2549_), .C(new_n2548_), .D(new_n368_), .Y(new_n2551_));
  OAI22X1  g02487(.A0(new_n119_), .A1(new_n108_), .B0(new_n75_), .B1(new_n72_), .Y(new_n2552_));
  OR4X1    g02488(.A(new_n2552_), .B(new_n1550_), .C(new_n1473_), .D(new_n636_), .Y(new_n2553_));
  OR4X1    g02489(.A(new_n2553_), .B(new_n494_), .C(new_n814_), .D(new_n256_), .Y(new_n2554_));
  OR4X1    g02490(.A(new_n642_), .B(new_n496_), .C(new_n224_), .D(new_n172_), .Y(new_n2555_));
  OR4X1    g02491(.A(new_n372_), .B(new_n286_), .C(new_n251_), .D(new_n449_), .Y(new_n2556_));
  OR4X1    g02492(.A(new_n2556_), .B(new_n2555_), .C(new_n1485_), .D(new_n298_), .Y(new_n2557_));
  OR4X1    g02493(.A(new_n1757_), .B(new_n959_), .C(new_n723_), .D(new_n370_), .Y(new_n2558_));
  OR4X1    g02494(.A(new_n2558_), .B(new_n2557_), .C(new_n2554_), .D(new_n1945_), .Y(new_n2559_));
  NOR4X1   g02495(.A(new_n2559_), .B(new_n2551_), .C(new_n2547_), .D(new_n2539_), .Y(new_n2560_));
  OAI22X1  g02496(.A0(new_n168_), .A1(new_n161_), .B0(new_n125_), .B1(new_n79_), .Y(new_n2561_));
  OR4X1    g02497(.A(new_n2561_), .B(new_n1778_), .C(new_n296_), .D(new_n180_), .Y(new_n2562_));
  OAI22X1  g02498(.A0(new_n108_), .A1(new_n115_), .B0(new_n106_), .B1(new_n81_), .Y(new_n2563_));
  OR2X1    g02499(.A(new_n2563_), .B(new_n144_), .Y(new_n2564_));
  OR2X1    g02500(.A(new_n1407_), .B(new_n1965_), .Y(new_n2565_));
  NOR4X1   g02501(.A(new_n2565_), .B(new_n2564_), .C(new_n2562_), .D(new_n2469_), .Y(new_n2566_));
  OR4X1    g02502(.A(new_n1516_), .B(new_n531_), .C(new_n717_), .D(new_n118_), .Y(new_n2567_));
  OR4X1    g02503(.A(new_n527_), .B(new_n510_), .C(new_n505_), .D(new_n523_), .Y(new_n2568_));
  OR4X1    g02504(.A(new_n383_), .B(new_n421_), .C(new_n371_), .D(new_n350_), .Y(new_n2569_));
  NOR4X1   g02505(.A(new_n2569_), .B(new_n2568_), .C(new_n2567_), .D(new_n2520_), .Y(new_n2570_));
  NAND3X1  g02506(.A(new_n2570_), .B(new_n2566_), .C(new_n2135_), .Y(new_n2571_));
  INVX1    g02507(.A(new_n1559_), .Y(new_n2572_));
  OR4X1    g02508(.A(new_n478_), .B(new_n251_), .C(new_n229_), .D(new_n213_), .Y(new_n2573_));
  NOR4X1   g02509(.A(new_n679_), .B(new_n422_), .C(new_n385_), .D(new_n274_), .Y(new_n2574_));
  NOR4X1   g02510(.A(new_n261_), .B(new_n240_), .C(new_n197_), .D(new_n156_), .Y(new_n2575_));
  NAND2X1  g02511(.A(new_n2575_), .B(new_n2574_), .Y(new_n2576_));
  OR4X1    g02512(.A(new_n2576_), .B(new_n2573_), .C(new_n778_), .D(new_n666_), .Y(new_n2577_));
  OR4X1    g02513(.A(new_n873_), .B(new_n743_), .C(new_n194_), .D(new_n338_), .Y(new_n2578_));
  OR4X1    g02514(.A(new_n2578_), .B(new_n2577_), .C(new_n2011_), .D(new_n2572_), .Y(new_n2579_));
  OAI22X1  g02515(.A0(new_n148_), .A1(new_n94_), .B0(new_n108_), .B1(new_n84_), .Y(new_n2580_));
  OR4X1    g02516(.A(new_n2580_), .B(new_n882_), .C(new_n400_), .D(new_n196_), .Y(new_n2581_));
  OR4X1    g02517(.A(new_n475_), .B(new_n418_), .C(new_n483_), .D(new_n323_), .Y(new_n2582_));
  OR4X1    g02518(.A(new_n2582_), .B(new_n2581_), .C(new_n1575_), .D(new_n943_), .Y(new_n2583_));
  OAI22X1  g02519(.A0(new_n152_), .A1(new_n143_), .B0(new_n125_), .B1(new_n91_), .Y(new_n2584_));
  OR4X1    g02520(.A(new_n2584_), .B(new_n547_), .C(new_n158_), .D(new_n1008_), .Y(new_n2585_));
  OR2X1    g02521(.A(new_n2585_), .B(new_n1241_), .Y(new_n2586_));
  OAI22X1  g02522(.A0(new_n182_), .A1(new_n79_), .B0(new_n148_), .B1(new_n143_), .Y(new_n2587_));
  OR4X1    g02523(.A(new_n2587_), .B(new_n2105_), .C(new_n868_), .D(new_n594_), .Y(new_n2588_));
  OR2X1    g02524(.A(new_n1408_), .B(new_n1319_), .Y(new_n2589_));
  OR4X1    g02525(.A(new_n1398_), .B(new_n540_), .C(new_n265_), .D(new_n139_), .Y(new_n2590_));
  OR2X1    g02526(.A(new_n1062_), .B(new_n766_), .Y(new_n2591_));
  OR4X1    g02527(.A(new_n2591_), .B(new_n2590_), .C(new_n2589_), .D(new_n1717_), .Y(new_n2592_));
  OR4X1    g02528(.A(new_n2592_), .B(new_n2588_), .C(new_n2586_), .D(new_n2583_), .Y(new_n2593_));
  NOR3X1   g02529(.A(new_n2593_), .B(new_n2579_), .C(new_n2571_), .Y(new_n2594_));
  NOR2X1   g02530(.A(new_n2594_), .B(new_n2560_), .Y(new_n2595_));
  NAND2X1  g02531(.A(new_n2594_), .B(new_n2560_), .Y(new_n2596_));
  AOI21X1  g02532(.A0(new_n2596_), .A1(new_n2529_), .B0(new_n2595_), .Y(new_n2597_));
  NOR2X1   g02533(.A(new_n2597_), .B(new_n2528_), .Y(new_n2598_));
  INVX1    g02534(.A(new_n1830_), .Y(new_n2599_));
  XOR2X1   g02535(.A(new_n2599_), .B(new_n1829_), .Y(new_n2600_));
  INVX1    g02536(.A(new_n2600_), .Y(new_n2601_));
  INVX1    g02537(.A(new_n903_), .Y(new_n2602_));
  INVX1    g02538(.A(new_n985_), .Y(new_n2603_));
  AOI22X1  g02539(.A0(new_n1890_), .A1(new_n2603_), .B0(new_n1889_), .B1(new_n2602_), .Y(new_n2604_));
  OAI21X1  g02540(.A0(new_n1885_), .A1(new_n957_), .B0(new_n2604_), .Y(new_n2605_));
  AOI21X1  g02541(.A0(new_n2601_), .A1(new_n407_), .B0(new_n2605_), .Y(new_n2606_));
  INVX1    g02542(.A(new_n2606_), .Y(new_n2607_));
  XOR2X1   g02543(.A(new_n2597_), .B(new_n2528_), .Y(new_n2608_));
  AOI21X1  g02544(.A0(new_n2608_), .A1(new_n2607_), .B0(new_n2598_), .Y(new_n2609_));
  NOR2X1   g02545(.A(new_n2528_), .B(new_n2456_), .Y(new_n2610_));
  OAI21X1  g02546(.A0(new_n2610_), .A1(new_n2609_), .B0(new_n2527_), .Y(new_n2611_));
  XOR2X1   g02547(.A(new_n2497_), .B(new_n2493_), .Y(new_n2612_));
  AOI21X1  g02548(.A0(new_n2612_), .A1(new_n2611_), .B0(new_n2498_), .Y(new_n2613_));
  OR2X1    g02549(.A(new_n2613_), .B(new_n2490_), .Y(new_n2614_));
  INVX1    g02550(.A(new_n2490_), .Y(new_n2615_));
  XOR2X1   g02551(.A(new_n2613_), .B(new_n2615_), .Y(new_n2616_));
  OAI22X1  g02552(.A0(new_n2186_), .A1(new_n623_), .B0(new_n2140_), .B1(new_n1879_), .Y(new_n2617_));
  AOI21X1  g02553(.A0(new_n2095_), .A1(new_n2048_), .B0(new_n2617_), .Y(new_n2618_));
  OAI21X1  g02554(.A0(new_n2063_), .A1(new_n1881_), .B0(new_n2618_), .Y(new_n2619_));
  XOR2X1   g02555(.A(new_n2619_), .B(new_n74_), .Y(new_n2620_));
  OAI21X1  g02556(.A0(new_n2620_), .A1(new_n2616_), .B0(new_n2614_), .Y(new_n2621_));
  AOI21X1  g02557(.A0(new_n2621_), .A1(new_n2489_), .B0(new_n2488_), .Y(new_n2622_));
  OAI21X1  g02558(.A0(new_n2622_), .A1(new_n2440_), .B0(new_n2438_), .Y(new_n2623_));
  XOR2X1   g02559(.A(new_n2204_), .B(new_n2059_), .Y(new_n2624_));
  XOR2X1   g02560(.A(new_n2386_), .B(new_n2384_), .Y(new_n2625_));
  INVX1    g02561(.A(new_n2423_), .Y(new_n2626_));
  INVX1    g02562(.A(new_n2287_), .Y(new_n2627_));
  AOI22X1  g02563(.A0(new_n2424_), .A1(new_n2627_), .B0(new_n2418_), .B1(new_n2420_), .Y(new_n2628_));
  OAI21X1  g02564(.A0(new_n2626_), .A1(new_n2379_), .B0(new_n2628_), .Y(new_n2629_));
  AOI21X1  g02565(.A0(new_n2625_), .A1(new_n2301_), .B0(new_n2629_), .Y(new_n2630_));
  XOR2X1   g02566(.A(new_n2630_), .B(\a[26] ), .Y(new_n2631_));
  INVX1    g02567(.A(new_n2623_), .Y(new_n2632_));
  XOR2X1   g02568(.A(new_n2624_), .B(new_n2632_), .Y(new_n2633_));
  NOR2X1   g02569(.A(new_n2633_), .B(new_n2631_), .Y(new_n2634_));
  AOI21X1  g02570(.A0(new_n2624_), .A1(new_n2623_), .B0(new_n2634_), .Y(new_n2635_));
  NOR3X1   g02571(.A(new_n1478_), .B(new_n1319_), .C(new_n1096_), .Y(new_n2636_));
  NOR4X1   g02572(.A(new_n356_), .B(new_n300_), .C(new_n176_), .D(new_n85_), .Y(new_n2637_));
  NOR3X1   g02573(.A(new_n676_), .B(new_n578_), .C(new_n337_), .Y(new_n2638_));
  NAND3X1  g02574(.A(new_n2638_), .B(new_n2637_), .C(new_n2636_), .Y(new_n2639_));
  AOI21X1  g02575(.A0(new_n182_), .A1(new_n105_), .B0(new_n84_), .Y(new_n2640_));
  AOI21X1  g02576(.A0(new_n94_), .A1(new_n78_), .B0(new_n84_), .Y(new_n2641_));
  OR4X1    g02577(.A(new_n2641_), .B(new_n2640_), .C(new_n1408_), .D(new_n724_), .Y(new_n2642_));
  OR4X1    g02578(.A(new_n1608_), .B(new_n1114_), .C(new_n594_), .D(new_n160_), .Y(new_n2643_));
  OR4X1    g02579(.A(new_n815_), .B(new_n301_), .C(new_n231_), .D(new_n200_), .Y(new_n2644_));
  OR4X1    g02580(.A(new_n2644_), .B(new_n494_), .C(new_n535_), .D(new_n307_), .Y(new_n2645_));
  OR4X1    g02581(.A(new_n2645_), .B(new_n2643_), .C(new_n2642_), .D(new_n2639_), .Y(new_n2646_));
  NOR4X1   g02582(.A(new_n2646_), .B(new_n2376_), .C(new_n510_), .D(new_n197_), .Y(new_n2647_));
  AND2X1   g02583(.A(new_n2647_), .B(new_n2412_), .Y(new_n2648_));
  INVX1    g02584(.A(new_n2648_), .Y(new_n2649_));
  NOR2X1   g02585(.A(new_n2414_), .B(new_n2379_), .Y(new_n2650_));
  AOI21X1  g02586(.A0(new_n2415_), .A1(new_n2388_), .B0(new_n2650_), .Y(new_n2651_));
  AOI21X1  g02587(.A0(new_n2651_), .A1(new_n2414_), .B0(new_n2648_), .Y(new_n2652_));
  XOR2X1   g02588(.A(new_n70_), .B(\a[22] ), .Y(new_n2653_));
  XOR2X1   g02589(.A(\a[22] ), .B(\a[21] ), .Y(new_n2654_));
  XOR2X1   g02590(.A(\a[21] ), .B(new_n1920_), .Y(new_n2655_));
  INVX1    g02591(.A(new_n2655_), .Y(new_n2656_));
  NOR3X1   g02592(.A(new_n2656_), .B(new_n2654_), .C(new_n2653_), .Y(new_n2657_));
  NOR2X1   g02593(.A(new_n2655_), .B(new_n2653_), .Y(new_n2658_));
  AOI22X1  g02594(.A0(new_n2658_), .A1(new_n2652_), .B0(new_n2657_), .B1(new_n2649_), .Y(new_n2659_));
  XOR2X1   g02595(.A(new_n2659_), .B(\a[23] ), .Y(new_n2660_));
  XOR2X1   g02596(.A(new_n2660_), .B(new_n2635_), .Y(new_n2661_));
  XOR2X1   g02597(.A(new_n2661_), .B(new_n2429_), .Y(new_n2662_));
  XOR2X1   g02598(.A(new_n2622_), .B(new_n2440_), .Y(new_n2663_));
  INVX1    g02599(.A(new_n2663_), .Y(new_n2664_));
  INVX1    g02600(.A(new_n2301_), .Y(new_n2665_));
  INVX1    g02601(.A(new_n2424_), .Y(new_n2666_));
  OAI22X1  g02602(.A0(new_n2666_), .A1(new_n2137_), .B0(new_n2626_), .B1(new_n2339_), .Y(new_n2667_));
  AOI21X1  g02603(.A0(new_n2418_), .A1(new_n2627_), .B0(new_n2667_), .Y(new_n2668_));
  XOR2X1   g02604(.A(new_n2383_), .B(new_n2382_), .Y(new_n2669_));
  INVX1    g02605(.A(new_n2669_), .Y(new_n2670_));
  OAI21X1  g02606(.A0(new_n2670_), .A1(new_n2665_), .B0(new_n2668_), .Y(new_n2671_));
  XOR2X1   g02607(.A(new_n2671_), .B(new_n89_), .Y(new_n2672_));
  OR2X1    g02608(.A(new_n2672_), .B(new_n2664_), .Y(new_n2673_));
  INVX1    g02609(.A(new_n2489_), .Y(new_n2674_));
  XOR2X1   g02610(.A(new_n2621_), .B(new_n2674_), .Y(new_n2675_));
  OAI22X1  g02611(.A0(new_n2186_), .A1(new_n520_), .B0(new_n2183_), .B1(new_n2140_), .Y(new_n2676_));
  AOI21X1  g02612(.A0(new_n2095_), .A1(new_n1887_), .B0(new_n2676_), .Y(new_n2677_));
  OAI21X1  g02613(.A0(new_n2243_), .A1(new_n2063_), .B0(new_n2677_), .Y(new_n2678_));
  XOR2X1   g02614(.A(new_n2678_), .B(new_n74_), .Y(new_n2679_));
  NOR2X1   g02615(.A(new_n2679_), .B(new_n2675_), .Y(new_n2680_));
  AOI22X1  g02616(.A0(new_n2424_), .A1(new_n2093_), .B0(new_n2423_), .B1(new_n2627_), .Y(new_n2681_));
  OAI21X1  g02617(.A0(new_n2419_), .A1(new_n2137_), .B0(new_n2681_), .Y(new_n2682_));
  AOI21X1  g02618(.A0(new_n2301_), .A1(new_n2294_), .B0(new_n2682_), .Y(new_n2683_));
  XOR2X1   g02619(.A(new_n2683_), .B(\a[26] ), .Y(new_n2684_));
  INVX1    g02620(.A(new_n2684_), .Y(new_n2685_));
  XOR2X1   g02621(.A(new_n2679_), .B(new_n2675_), .Y(new_n2686_));
  AOI21X1  g02622(.A0(new_n2686_), .A1(new_n2685_), .B0(new_n2680_), .Y(new_n2687_));
  XOR2X1   g02623(.A(new_n2672_), .B(new_n2663_), .Y(new_n2688_));
  OAI21X1  g02624(.A0(new_n2688_), .A1(new_n2687_), .B0(new_n2673_), .Y(new_n2689_));
  XOR2X1   g02625(.A(new_n2633_), .B(new_n2631_), .Y(new_n2690_));
  AND2X1   g02626(.A(new_n2690_), .B(new_n2689_), .Y(new_n2691_));
  INVX1    g02627(.A(new_n2658_), .Y(new_n2692_));
  INVX1    g02628(.A(new_n2652_), .Y(new_n2693_));
  OAI21X1  g02629(.A0(new_n2651_), .A1(new_n2414_), .B0(new_n2648_), .Y(new_n2694_));
  NAND2X1  g02630(.A(new_n2694_), .B(new_n2693_), .Y(new_n2695_));
  AND2X1   g02631(.A(new_n2655_), .B(new_n2654_), .Y(new_n2696_));
  AOI22X1  g02632(.A0(new_n2696_), .A1(new_n2649_), .B0(new_n2657_), .B1(new_n2421_), .Y(new_n2697_));
  OAI21X1  g02633(.A0(new_n2695_), .A1(new_n2692_), .B0(new_n2697_), .Y(new_n2698_));
  XOR2X1   g02634(.A(new_n2698_), .B(\a[23] ), .Y(new_n2699_));
  XOR2X1   g02635(.A(new_n2690_), .B(new_n2689_), .Y(new_n2700_));
  AOI21X1  g02636(.A0(new_n2700_), .A1(new_n2699_), .B0(new_n2691_), .Y(new_n2701_));
  XOR2X1   g02637(.A(new_n2701_), .B(new_n2662_), .Y(new_n2702_));
  INVX1    g02638(.A(new_n2702_), .Y(new_n2703_));
  XOR2X1   g02639(.A(new_n2686_), .B(new_n2684_), .Y(new_n2704_));
  XOR2X1   g02640(.A(new_n2528_), .B(new_n2456_), .Y(new_n2705_));
  OAI22X1  g02641(.A0(new_n2611_), .A1(new_n2610_), .B0(new_n2705_), .B1(new_n2609_), .Y(new_n2706_));
  AOI21X1  g02642(.A0(new_n1830_), .A1(new_n1829_), .B0(new_n956_), .Y(new_n2707_));
  XOR2X1   g02643(.A(new_n1832_), .B(new_n2707_), .Y(new_n2708_));
  INVX1    g02644(.A(new_n2708_), .Y(new_n2709_));
  AOI22X1  g02645(.A0(new_n1889_), .A1(new_n2481_), .B0(new_n1884_), .B1(new_n2602_), .Y(new_n2710_));
  OAI21X1  g02646(.A0(new_n2245_), .A1(new_n957_), .B0(new_n2710_), .Y(new_n2711_));
  AOI21X1  g02647(.A0(new_n2709_), .A1(new_n407_), .B0(new_n2711_), .Y(new_n2712_));
  INVX1    g02648(.A(new_n2712_), .Y(new_n2713_));
  NAND2X1  g02649(.A(new_n2713_), .B(new_n2706_), .Y(new_n2714_));
  AOI22X1  g02650(.A0(new_n2185_), .A1(new_n2036_), .B0(new_n2139_), .B1(new_n1886_), .Y(new_n2715_));
  OAI21X1  g02651(.A0(new_n2431_), .A1(new_n690_), .B0(new_n2715_), .Y(new_n2716_));
  AOI21X1  g02652(.A0(new_n2062_), .A1(new_n2035_), .B0(new_n2716_), .Y(new_n2717_));
  XOR2X1   g02653(.A(new_n2717_), .B(\a[29] ), .Y(new_n2718_));
  XOR2X1   g02654(.A(new_n2712_), .B(new_n2706_), .Y(new_n2719_));
  OAI21X1  g02655(.A0(new_n2719_), .A1(new_n2718_), .B0(new_n2714_), .Y(new_n2720_));
  XOR2X1   g02656(.A(new_n2612_), .B(new_n2611_), .Y(new_n2721_));
  AND2X1   g02657(.A(new_n2721_), .B(new_n2720_), .Y(new_n2722_));
  AOI22X1  g02658(.A0(new_n2185_), .A1(new_n2049_), .B0(new_n2139_), .B1(new_n2048_), .Y(new_n2723_));
  OAI21X1  g02659(.A0(new_n2431_), .A1(new_n623_), .B0(new_n2723_), .Y(new_n2724_));
  AOI21X1  g02660(.A0(new_n2062_), .A1(new_n2047_), .B0(new_n2724_), .Y(new_n2725_));
  XOR2X1   g02661(.A(new_n2725_), .B(\a[29] ), .Y(new_n2726_));
  INVX1    g02662(.A(new_n2726_), .Y(new_n2727_));
  XOR2X1   g02663(.A(new_n2721_), .B(new_n2720_), .Y(new_n2728_));
  AOI21X1  g02664(.A0(new_n2728_), .A1(new_n2727_), .B0(new_n2722_), .Y(new_n2729_));
  INVX1    g02665(.A(new_n2729_), .Y(new_n2730_));
  XOR2X1   g02666(.A(new_n2620_), .B(new_n2616_), .Y(new_n2731_));
  AND2X1   g02667(.A(new_n2731_), .B(new_n2730_), .Y(new_n2732_));
  XOR2X1   g02668(.A(new_n2731_), .B(new_n2730_), .Y(new_n2733_));
  AOI22X1  g02669(.A0(new_n2424_), .A1(new_n2246_), .B0(new_n2423_), .B1(new_n2252_), .Y(new_n2734_));
  OAI21X1  g02670(.A0(new_n2419_), .A1(new_n2092_), .B0(new_n2734_), .Y(new_n2735_));
  AOI21X1  g02671(.A0(new_n2301_), .A1(new_n2201_), .B0(new_n2735_), .Y(new_n2736_));
  XOR2X1   g02672(.A(new_n2736_), .B(new_n89_), .Y(new_n2737_));
  AOI21X1  g02673(.A0(new_n2737_), .A1(new_n2733_), .B0(new_n2732_), .Y(new_n2738_));
  NOR2X1   g02674(.A(new_n2738_), .B(new_n2704_), .Y(new_n2739_));
  INVX1    g02675(.A(new_n2739_), .Y(new_n2740_));
  XOR2X1   g02676(.A(new_n2738_), .B(new_n2704_), .Y(new_n2741_));
  INVX1    g02677(.A(new_n2741_), .Y(new_n2742_));
  INVX1    g02678(.A(new_n2696_), .Y(new_n2743_));
  INVX1    g02679(.A(new_n2653_), .Y(new_n2744_));
  NOR2X1   g02680(.A(new_n2655_), .B(new_n2744_), .Y(new_n2745_));
  AOI22X1  g02681(.A0(new_n2745_), .A1(new_n2421_), .B0(new_n2657_), .B1(new_n2420_), .Y(new_n2746_));
  OAI21X1  g02682(.A0(new_n2743_), .A1(new_n2379_), .B0(new_n2746_), .Y(new_n2747_));
  AOI21X1  g02683(.A0(new_n2658_), .A1(new_n2416_), .B0(new_n2747_), .Y(new_n2748_));
  XOR2X1   g02684(.A(new_n2748_), .B(\a[23] ), .Y(new_n2749_));
  OAI21X1  g02685(.A0(new_n2749_), .A1(new_n2742_), .B0(new_n2740_), .Y(new_n2750_));
  INVX1    g02686(.A(new_n2750_), .Y(new_n2751_));
  INVX1    g02687(.A(new_n2379_), .Y(new_n2752_));
  INVX1    g02688(.A(new_n2745_), .Y(new_n2753_));
  OAI22X1  g02689(.A0(new_n2753_), .A1(new_n2648_), .B0(new_n2743_), .B1(new_n2414_), .Y(new_n2754_));
  AOI21X1  g02690(.A0(new_n2657_), .A1(new_n2752_), .B0(new_n2754_), .Y(new_n2755_));
  XOR2X1   g02691(.A(new_n2648_), .B(new_n2414_), .Y(new_n2756_));
  XOR2X1   g02692(.A(new_n2756_), .B(new_n2651_), .Y(new_n2757_));
  OAI21X1  g02693(.A0(new_n2757_), .A1(new_n2692_), .B0(new_n2755_), .Y(new_n2758_));
  XOR2X1   g02694(.A(new_n2758_), .B(new_n70_), .Y(new_n2759_));
  NOR2X1   g02695(.A(new_n2759_), .B(new_n2751_), .Y(new_n2760_));
  INVX1    g02696(.A(new_n2760_), .Y(new_n2761_));
  XOR2X1   g02697(.A(new_n2759_), .B(new_n2751_), .Y(new_n2762_));
  INVX1    g02698(.A(new_n2762_), .Y(new_n2763_));
  INVX1    g02699(.A(new_n2687_), .Y(new_n2764_));
  XOR2X1   g02700(.A(new_n2688_), .B(new_n2764_), .Y(new_n2765_));
  OAI21X1  g02701(.A0(new_n2765_), .A1(new_n2763_), .B0(new_n2761_), .Y(new_n2766_));
  XOR2X1   g02702(.A(new_n2700_), .B(new_n2699_), .Y(new_n2767_));
  AND2X1   g02703(.A(new_n2767_), .B(new_n2766_), .Y(new_n2768_));
  XOR2X1   g02704(.A(new_n2765_), .B(new_n2762_), .Y(new_n2769_));
  XOR2X1   g02705(.A(new_n2736_), .B(\a[26] ), .Y(new_n2770_));
  XOR2X1   g02706(.A(new_n2770_), .B(new_n2733_), .Y(new_n2771_));
  XOR2X1   g02707(.A(new_n2728_), .B(new_n2726_), .Y(new_n2772_));
  AOI22X1  g02708(.A0(new_n2424_), .A1(new_n1887_), .B0(new_n2423_), .B1(new_n2093_), .Y(new_n2773_));
  OAI21X1  g02709(.A0(new_n2419_), .A1(new_n2183_), .B0(new_n2773_), .Y(new_n2774_));
  AOI21X1  g02710(.A0(new_n2430_), .A1(new_n2301_), .B0(new_n2774_), .Y(new_n2775_));
  XOR2X1   g02711(.A(new_n2775_), .B(\a[26] ), .Y(new_n2776_));
  NOR2X1   g02712(.A(new_n2776_), .B(new_n2772_), .Y(new_n2777_));
  XOR2X1   g02713(.A(new_n2719_), .B(new_n2718_), .Y(new_n2778_));
  INVX1    g02714(.A(new_n2778_), .Y(new_n2779_));
  XOR2X1   g02715(.A(new_n2608_), .B(new_n2606_), .Y(new_n2780_));
  NOR2X1   g02716(.A(new_n2595_), .B(\a[14] ), .Y(new_n2781_));
  AOI21X1  g02717(.A0(new_n2781_), .A1(new_n2596_), .B0(\a[14] ), .Y(new_n2782_));
  AOI21X1  g02718(.A0(new_n2597_), .A1(new_n2596_), .B0(new_n2782_), .Y(new_n2783_));
  INVX1    g02719(.A(new_n2560_), .Y(new_n2784_));
  OAI22X1  g02720(.A0(new_n143_), .A1(new_n84_), .B0(new_n102_), .B1(new_n81_), .Y(new_n2785_));
  OR4X1    g02721(.A(new_n2785_), .B(new_n642_), .C(new_n596_), .D(new_n968_), .Y(new_n2786_));
  OR4X1    g02722(.A(new_n1274_), .B(new_n803_), .C(new_n535_), .D(new_n928_), .Y(new_n2787_));
  OR4X1    g02723(.A(new_n615_), .B(new_n598_), .C(new_n301_), .D(new_n259_), .Y(new_n2788_));
  OR4X1    g02724(.A(new_n2788_), .B(new_n2787_), .C(new_n2786_), .D(new_n1731_), .Y(new_n2789_));
  NOR2X1   g02725(.A(new_n394_), .B(new_n540_), .Y(new_n2790_));
  NOR4X1   g02726(.A(new_n691_), .B(new_n229_), .C(new_n217_), .D(new_n103_), .Y(new_n2791_));
  NAND4X1  g02727(.A(new_n2791_), .B(new_n2790_), .C(new_n1368_), .D(new_n551_), .Y(new_n2792_));
  OR4X1    g02728(.A(new_n634_), .B(new_n460_), .C(new_n717_), .D(new_n280_), .Y(new_n2793_));
  OR4X1    g02729(.A(new_n2793_), .B(new_n1912_), .C(new_n651_), .D(new_n337_), .Y(new_n2794_));
  OAI22X1  g02730(.A0(new_n127_), .A1(new_n115_), .B0(new_n123_), .B1(new_n94_), .Y(new_n2795_));
  OR4X1    g02731(.A(new_n2795_), .B(new_n1646_), .C(new_n1210_), .D(new_n561_), .Y(new_n2796_));
  OR4X1    g02732(.A(new_n2796_), .B(new_n2794_), .C(new_n2792_), .D(new_n1383_), .Y(new_n2797_));
  OR4X1    g02733(.A(new_n891_), .B(new_n831_), .C(new_n342_), .D(new_n164_), .Y(new_n2798_));
  OR4X1    g02734(.A(new_n263_), .B(new_n239_), .C(new_n194_), .D(new_n176_), .Y(new_n2799_));
  OR4X1    g02735(.A(new_n546_), .B(new_n329_), .C(new_n144_), .D(new_n307_), .Y(new_n2800_));
  NOR3X1   g02736(.A(new_n1090_), .B(new_n671_), .C(new_n391_), .Y(new_n2801_));
  NOR4X1   g02737(.A(new_n2451_), .B(new_n2209_), .C(new_n1547_), .D(new_n975_), .Y(new_n2802_));
  NAND3X1  g02738(.A(new_n2802_), .B(new_n2801_), .C(new_n448_), .Y(new_n2803_));
  OR4X1    g02739(.A(new_n2803_), .B(new_n2800_), .C(new_n2799_), .D(new_n2798_), .Y(new_n2804_));
  OR4X1    g02740(.A(new_n1608_), .B(new_n723_), .C(new_n885_), .D(new_n202_), .Y(new_n2805_));
  OAI22X1  g02741(.A0(new_n152_), .A1(new_n72_), .B0(new_n119_), .B1(new_n78_), .Y(new_n2806_));
  OR4X1    g02742(.A(new_n2806_), .B(new_n848_), .C(new_n531_), .D(new_n1044_), .Y(new_n2807_));
  OR4X1    g02743(.A(new_n681_), .B(new_n228_), .C(new_n536_), .D(new_n187_), .Y(new_n2808_));
  OR4X1    g02744(.A(new_n2808_), .B(new_n2807_), .C(new_n1390_), .D(new_n1467_), .Y(new_n2809_));
  OAI22X1  g02745(.A0(new_n99_), .A1(new_n96_), .B0(new_n94_), .B1(new_n88_), .Y(new_n2810_));
  NOR2X1   g02746(.A(new_n2810_), .B(new_n274_), .Y(new_n2811_));
  NOR3X1   g02747(.A(new_n1028_), .B(new_n370_), .C(new_n265_), .Y(new_n2812_));
  NOR3X1   g02748(.A(new_n1474_), .B(new_n426_), .C(new_n410_), .Y(new_n2813_));
  NAND3X1  g02749(.A(new_n2813_), .B(new_n2812_), .C(new_n2811_), .Y(new_n2814_));
  OAI22X1  g02750(.A0(new_n129_), .A1(new_n91_), .B0(new_n115_), .B1(new_n72_), .Y(new_n2815_));
  NOR3X1   g02751(.A(new_n2815_), .B(new_n386_), .C(new_n155_), .Y(new_n2816_));
  INVX1    g02752(.A(new_n2816_), .Y(new_n2817_));
  OR4X1    g02753(.A(new_n543_), .B(new_n395_), .C(new_n361_), .D(new_n603_), .Y(new_n2818_));
  OR4X1    g02754(.A(new_n2818_), .B(new_n2817_), .C(new_n1499_), .D(new_n429_), .Y(new_n2819_));
  NOR4X1   g02755(.A(new_n2819_), .B(new_n2814_), .C(new_n2809_), .D(new_n2805_), .Y(new_n2820_));
  INVX1    g02756(.A(new_n2820_), .Y(new_n2821_));
  NOR4X1   g02757(.A(new_n2821_), .B(new_n2804_), .C(new_n2797_), .D(new_n2789_), .Y(new_n2822_));
  NOR2X1   g02758(.A(new_n2822_), .B(new_n2784_), .Y(new_n2823_));
  XOR2X1   g02759(.A(new_n1826_), .B(new_n1825_), .Y(new_n2824_));
  AOI22X1  g02760(.A0(new_n1890_), .A1(new_n1126_), .B0(new_n1889_), .B1(new_n2603_), .Y(new_n2825_));
  OAI21X1  g02761(.A0(new_n1885_), .A1(new_n1065_), .B0(new_n2825_), .Y(new_n2826_));
  AOI21X1  g02762(.A0(new_n2824_), .A1(new_n407_), .B0(new_n2826_), .Y(new_n2827_));
  AND2X1   g02763(.A(new_n2822_), .B(new_n2784_), .Y(new_n2828_));
  NOR3X1   g02764(.A(new_n2828_), .B(new_n2827_), .C(new_n2823_), .Y(new_n2829_));
  NOR2X1   g02765(.A(new_n2829_), .B(new_n2823_), .Y(new_n2830_));
  NOR2X1   g02766(.A(new_n2830_), .B(new_n2783_), .Y(new_n2831_));
  XOR2X1   g02767(.A(new_n985_), .B(new_n957_), .Y(new_n2832_));
  XOR2X1   g02768(.A(new_n2832_), .B(new_n1827_), .Y(new_n2833_));
  INVX1    g02769(.A(new_n2833_), .Y(new_n2834_));
  INVX1    g02770(.A(new_n957_), .Y(new_n2835_));
  AOI22X1  g02771(.A0(new_n1889_), .A1(new_n2835_), .B0(new_n1884_), .B1(new_n2603_), .Y(new_n2836_));
  OAI21X1  g02772(.A0(new_n2245_), .A1(new_n1065_), .B0(new_n2836_), .Y(new_n2837_));
  AOI21X1  g02773(.A0(new_n2834_), .A1(new_n407_), .B0(new_n2837_), .Y(new_n2838_));
  INVX1    g02774(.A(new_n2838_), .Y(new_n2839_));
  XOR2X1   g02775(.A(new_n2830_), .B(new_n2783_), .Y(new_n2840_));
  AOI21X1  g02776(.A0(new_n2840_), .A1(new_n2839_), .B0(new_n2831_), .Y(new_n2841_));
  OR2X1    g02777(.A(new_n2841_), .B(new_n2780_), .Y(new_n2842_));
  INVX1    g02778(.A(new_n2780_), .Y(new_n2843_));
  XOR2X1   g02779(.A(new_n2841_), .B(new_n2843_), .Y(new_n2844_));
  INVX1    g02780(.A(new_n2480_), .Y(new_n2845_));
  OAI22X1  g02781(.A0(new_n2186_), .A1(new_n847_), .B0(new_n2140_), .B1(new_n690_), .Y(new_n2846_));
  AOI21X1  g02782(.A0(new_n2095_), .A1(new_n2036_), .B0(new_n2846_), .Y(new_n2847_));
  OAI21X1  g02783(.A0(new_n2845_), .A1(new_n2063_), .B0(new_n2847_), .Y(new_n2848_));
  XOR2X1   g02784(.A(new_n2848_), .B(new_n74_), .Y(new_n2849_));
  OR2X1    g02785(.A(new_n2849_), .B(new_n2844_), .Y(new_n2850_));
  AND2X1   g02786(.A(new_n2850_), .B(new_n2842_), .Y(new_n2851_));
  OR2X1    g02787(.A(new_n2851_), .B(new_n2779_), .Y(new_n2852_));
  XOR2X1   g02788(.A(new_n2851_), .B(new_n2779_), .Y(new_n2853_));
  INVX1    g02789(.A(new_n2853_), .Y(new_n2854_));
  AOI22X1  g02790(.A0(new_n2424_), .A1(new_n2048_), .B0(new_n2423_), .B1(new_n2246_), .Y(new_n2855_));
  OAI21X1  g02791(.A0(new_n2419_), .A1(new_n1879_), .B0(new_n2855_), .Y(new_n2856_));
  AOI21X1  g02792(.A0(new_n2301_), .A1(new_n2244_), .B0(new_n2856_), .Y(new_n2857_));
  XOR2X1   g02793(.A(new_n2857_), .B(\a[26] ), .Y(new_n2858_));
  OAI21X1  g02794(.A0(new_n2858_), .A1(new_n2854_), .B0(new_n2852_), .Y(new_n2859_));
  XOR2X1   g02795(.A(new_n2776_), .B(new_n2772_), .Y(new_n2860_));
  AOI21X1  g02796(.A0(new_n2860_), .A1(new_n2859_), .B0(new_n2777_), .Y(new_n2861_));
  NOR2X1   g02797(.A(new_n2861_), .B(new_n2771_), .Y(new_n2862_));
  XOR2X1   g02798(.A(new_n2861_), .B(new_n2771_), .Y(new_n2863_));
  AOI22X1  g02799(.A0(new_n2696_), .A1(new_n2420_), .B0(new_n2657_), .B1(new_n2627_), .Y(new_n2864_));
  OAI21X1  g02800(.A0(new_n2753_), .A1(new_n2379_), .B0(new_n2864_), .Y(new_n2865_));
  AOI21X1  g02801(.A0(new_n2658_), .A1(new_n2625_), .B0(new_n2865_), .Y(new_n2866_));
  XOR2X1   g02802(.A(new_n2866_), .B(new_n70_), .Y(new_n2867_));
  AOI21X1  g02803(.A0(new_n2867_), .A1(new_n2863_), .B0(new_n2862_), .Y(new_n2868_));
  XOR2X1   g02804(.A(\a[18] ), .B(new_n2445_), .Y(new_n2869_));
  INVX1    g02805(.A(new_n2869_), .Y(new_n2870_));
  INVX1    g02806(.A(\a[19] ), .Y(new_n2871_));
  XOR2X1   g02807(.A(new_n2871_), .B(\a[18] ), .Y(new_n2872_));
  INVX1    g02808(.A(new_n2872_), .Y(new_n2873_));
  XOR2X1   g02809(.A(\a[20] ), .B(new_n2871_), .Y(new_n2874_));
  NOR3X1   g02810(.A(new_n2874_), .B(new_n2873_), .C(new_n2870_), .Y(new_n2875_));
  NOR2X1   g02811(.A(new_n2874_), .B(new_n2869_), .Y(new_n2876_));
  AOI22X1  g02812(.A0(new_n2876_), .A1(new_n2652_), .B0(new_n2875_), .B1(new_n2649_), .Y(new_n2877_));
  XOR2X1   g02813(.A(new_n2877_), .B(\a[20] ), .Y(new_n2878_));
  NOR2X1   g02814(.A(new_n2878_), .B(new_n2868_), .Y(new_n2879_));
  XOR2X1   g02815(.A(new_n2749_), .B(new_n2741_), .Y(new_n2880_));
  INVX1    g02816(.A(new_n2880_), .Y(new_n2881_));
  XOR2X1   g02817(.A(new_n2878_), .B(new_n2868_), .Y(new_n2882_));
  AOI21X1  g02818(.A0(new_n2882_), .A1(new_n2881_), .B0(new_n2879_), .Y(new_n2883_));
  NOR2X1   g02819(.A(new_n2883_), .B(new_n2769_), .Y(new_n2884_));
  INVX1    g02820(.A(new_n2884_), .Y(new_n2885_));
  XOR2X1   g02821(.A(new_n2883_), .B(new_n2769_), .Y(new_n2886_));
  INVX1    g02822(.A(new_n2886_), .Y(new_n2887_));
  XOR2X1   g02823(.A(new_n2882_), .B(new_n2880_), .Y(new_n2888_));
  XOR2X1   g02824(.A(new_n2867_), .B(new_n2863_), .Y(new_n2889_));
  INVX1    g02825(.A(new_n2889_), .Y(new_n2890_));
  AOI22X1  g02826(.A0(new_n2745_), .A1(new_n2420_), .B0(new_n2657_), .B1(new_n2252_), .Y(new_n2891_));
  OAI21X1  g02827(.A0(new_n2743_), .A1(new_n2287_), .B0(new_n2891_), .Y(new_n2892_));
  AOI21X1  g02828(.A0(new_n2669_), .A1(new_n2658_), .B0(new_n2892_), .Y(new_n2893_));
  XOR2X1   g02829(.A(new_n2893_), .B(\a[23] ), .Y(new_n2894_));
  INVX1    g02830(.A(new_n2894_), .Y(new_n2895_));
  XOR2X1   g02831(.A(new_n2860_), .B(new_n2859_), .Y(new_n2896_));
  XOR2X1   g02832(.A(new_n2896_), .B(new_n2894_), .Y(new_n2897_));
  XOR2X1   g02833(.A(new_n2858_), .B(new_n2853_), .Y(new_n2898_));
  AOI22X1  g02834(.A0(new_n2185_), .A1(new_n2602_), .B0(new_n2139_), .B1(new_n2036_), .Y(new_n2899_));
  OAI21X1  g02835(.A0(new_n2431_), .A1(new_n847_), .B0(new_n2899_), .Y(new_n2900_));
  AOI21X1  g02836(.A0(new_n2494_), .A1(new_n2062_), .B0(new_n2900_), .Y(new_n2901_));
  XOR2X1   g02837(.A(new_n2901_), .B(\a[29] ), .Y(new_n2902_));
  XOR2X1   g02838(.A(new_n2840_), .B(new_n2838_), .Y(new_n2903_));
  NOR2X1   g02839(.A(new_n2903_), .B(new_n2902_), .Y(new_n2904_));
  INVX1    g02840(.A(new_n2904_), .Y(new_n2905_));
  XOR2X1   g02841(.A(new_n2903_), .B(new_n2902_), .Y(new_n2906_));
  INVX1    g02842(.A(new_n2906_), .Y(new_n2907_));
  INVX1    g02843(.A(new_n2828_), .Y(new_n2908_));
  NOR2X1   g02844(.A(new_n2829_), .B(new_n2827_), .Y(new_n2909_));
  AOI21X1  g02845(.A0(new_n2830_), .A1(new_n2908_), .B0(new_n2909_), .Y(new_n2910_));
  INVX1    g02846(.A(\a[11] ), .Y(new_n2911_));
  OR4X1    g02847(.A(new_n720_), .B(new_n523_), .C(new_n627_), .D(new_n226_), .Y(new_n2912_));
  OR4X1    g02848(.A(new_n2912_), .B(new_n1443_), .C(new_n631_), .D(new_n234_), .Y(new_n2913_));
  OAI22X1  g02849(.A0(new_n152_), .A1(new_n90_), .B0(new_n129_), .B1(new_n79_), .Y(new_n2914_));
  OR2X1    g02850(.A(new_n2914_), .B(new_n328_), .Y(new_n2915_));
  NOR3X1   g02851(.A(new_n540_), .B(new_n457_), .C(new_n928_), .Y(new_n2916_));
  INVX1    g02852(.A(new_n2916_), .Y(new_n2917_));
  OR4X1    g02853(.A(new_n2917_), .B(new_n2915_), .C(new_n2913_), .D(new_n210_), .Y(new_n2918_));
  OR2X1    g02854(.A(new_n2554_), .B(new_n1193_), .Y(new_n2919_));
  OAI22X1  g02855(.A0(new_n129_), .A1(new_n117_), .B0(new_n90_), .B1(new_n88_), .Y(new_n2920_));
  NOR3X1   g02856(.A(new_n2920_), .B(new_n2580_), .C(new_n2302_), .Y(new_n2921_));
  OR4X1    g02857(.A(new_n265_), .B(new_n264_), .C(new_n243_), .D(new_n535_), .Y(new_n2922_));
  NOR3X1   g02858(.A(new_n2922_), .B(new_n560_), .C(new_n335_), .Y(new_n2923_));
  NOR4X1   g02859(.A(new_n1660_), .B(new_n500_), .C(new_n327_), .D(new_n307_), .Y(new_n2924_));
  NAND3X1  g02860(.A(new_n2924_), .B(new_n2923_), .C(new_n2921_), .Y(new_n2925_));
  OR4X1    g02861(.A(new_n615_), .B(new_n717_), .C(new_n474_), .D(new_n224_), .Y(new_n2926_));
  OR4X1    g02862(.A(new_n2926_), .B(new_n691_), .C(new_n194_), .D(new_n338_), .Y(new_n2927_));
  NAND4X1  g02863(.A(new_n1327_), .B(new_n989_), .C(new_n1151_), .D(new_n804_), .Y(new_n2928_));
  OR4X1    g02864(.A(new_n459_), .B(new_n815_), .C(new_n702_), .D(new_n100_), .Y(new_n2929_));
  OR4X1    g02865(.A(new_n2929_), .B(new_n1259_), .C(new_n232_), .D(new_n149_), .Y(new_n2930_));
  OR4X1    g02866(.A(new_n246_), .B(new_n974_), .C(new_n1087_), .D(new_n1284_), .Y(new_n2931_));
  OR4X1    g02867(.A(new_n2931_), .B(new_n1962_), .C(new_n1398_), .D(new_n395_), .Y(new_n2932_));
  OR4X1    g02868(.A(new_n2932_), .B(new_n2930_), .C(new_n2928_), .D(new_n2927_), .Y(new_n2933_));
  OR4X1    g02869(.A(new_n2933_), .B(new_n2925_), .C(new_n2919_), .D(new_n2918_), .Y(new_n2934_));
  NOR2X1   g02870(.A(new_n2934_), .B(new_n1854_), .Y(new_n2935_));
  OR4X1    g02871(.A(new_n1912_), .B(new_n657_), .C(new_n785_), .D(new_n153_), .Y(new_n2936_));
  OR4X1    g02872(.A(new_n396_), .B(new_n540_), .C(new_n627_), .D(new_n274_), .Y(new_n2937_));
  OAI22X1  g02873(.A0(new_n152_), .A1(new_n92_), .B0(new_n84_), .B1(new_n81_), .Y(new_n2938_));
  OR4X1    g02874(.A(new_n2938_), .B(new_n2937_), .C(new_n2936_), .D(new_n543_), .Y(new_n2939_));
  NOR4X1   g02875(.A(new_n300_), .B(new_n144_), .C(new_n139_), .D(new_n981_), .Y(new_n2940_));
  NOR2X1   g02876(.A(new_n441_), .B(new_n238_), .Y(new_n2941_));
  NOR3X1   g02877(.A(new_n740_), .B(new_n246_), .C(new_n338_), .Y(new_n2942_));
  NOR4X1   g02878(.A(new_n741_), .B(new_n702_), .C(new_n319_), .D(new_n280_), .Y(new_n2943_));
  NAND4X1  g02879(.A(new_n2943_), .B(new_n2942_), .C(new_n2941_), .D(new_n2940_), .Y(new_n2944_));
  OAI22X1  g02880(.A0(new_n123_), .A1(new_n72_), .B0(new_n99_), .B1(new_n75_), .Y(new_n2945_));
  OR4X1    g02881(.A(new_n2945_), .B(new_n1256_), .C(new_n1238_), .D(new_n882_), .Y(new_n2946_));
  OR4X1    g02882(.A(new_n2946_), .B(new_n2944_), .C(new_n2939_), .D(new_n639_), .Y(new_n2947_));
  OR4X1    g02883(.A(new_n201_), .B(new_n156_), .C(new_n134_), .D(new_n521_), .Y(new_n2948_));
  OR4X1    g02884(.A(new_n2948_), .B(new_n848_), .C(new_n546_), .D(new_n497_), .Y(new_n2949_));
  OR4X1    g02885(.A(new_n1082_), .B(new_n815_), .C(new_n565_), .D(new_n199_), .Y(new_n2950_));
  OR4X1    g02886(.A(new_n2950_), .B(new_n1134_), .C(new_n385_), .D(new_n819_), .Y(new_n2951_));
  OR4X1    g02887(.A(new_n1478_), .B(new_n1461_), .C(new_n729_), .D(new_n570_), .Y(new_n2952_));
  AOI21X1  g02888(.A0(new_n91_), .A1(new_n84_), .B0(new_n161_), .Y(new_n2953_));
  OR4X1    g02889(.A(new_n2953_), .B(new_n559_), .C(new_n465_), .D(new_n333_), .Y(new_n2954_));
  OR4X1    g02890(.A(new_n2954_), .B(new_n2952_), .C(new_n2951_), .D(new_n2949_), .Y(new_n2955_));
  OR4X1    g02891(.A(new_n2955_), .B(new_n2925_), .C(new_n2213_), .D(new_n1936_), .Y(new_n2956_));
  NOR2X1   g02892(.A(new_n2956_), .B(new_n2947_), .Y(new_n2957_));
  NOR2X1   g02893(.A(new_n2957_), .B(new_n2935_), .Y(new_n2958_));
  OR4X1    g02894(.A(new_n2956_), .B(new_n2947_), .C(new_n2934_), .D(new_n1854_), .Y(new_n2959_));
  AOI21X1  g02895(.A0(new_n2959_), .A1(new_n2911_), .B0(new_n2958_), .Y(new_n2960_));
  NOR2X1   g02896(.A(new_n2960_), .B(new_n2784_), .Y(new_n2961_));
  OR2X1    g02897(.A(new_n1821_), .B(new_n1188_), .Y(new_n2962_));
  XOR2X1   g02898(.A(new_n1823_), .B(new_n2962_), .Y(new_n2963_));
  AOI22X1  g02899(.A0(new_n1889_), .A1(new_n1822_), .B0(new_n1884_), .B1(new_n1126_), .Y(new_n2964_));
  OAI21X1  g02900(.A0(new_n2245_), .A1(new_n1189_), .B0(new_n2964_), .Y(new_n2965_));
  AOI21X1  g02901(.A0(new_n2963_), .A1(new_n407_), .B0(new_n2965_), .Y(new_n2966_));
  INVX1    g02902(.A(new_n2966_), .Y(new_n2967_));
  XOR2X1   g02903(.A(new_n2960_), .B(new_n2784_), .Y(new_n2968_));
  AOI21X1  g02904(.A0(new_n2968_), .A1(new_n2967_), .B0(new_n2961_), .Y(new_n2969_));
  NOR2X1   g02905(.A(new_n2969_), .B(new_n2910_), .Y(new_n2970_));
  XOR2X1   g02906(.A(new_n2969_), .B(new_n2910_), .Y(new_n2971_));
  XOR2X1   g02907(.A(new_n2968_), .B(new_n2966_), .Y(new_n2972_));
  NOR2X1   g02908(.A(new_n2958_), .B(\a[11] ), .Y(new_n2973_));
  AOI21X1  g02909(.A0(new_n2973_), .A1(new_n2959_), .B0(\a[11] ), .Y(new_n2974_));
  AOI21X1  g02910(.A0(new_n2960_), .A1(new_n2959_), .B0(new_n2974_), .Y(new_n2975_));
  XOR2X1   g02911(.A(new_n1820_), .B(new_n1819_), .Y(new_n2976_));
  INVX1    g02912(.A(new_n1236_), .Y(new_n2977_));
  AOI22X1  g02913(.A0(new_n1890_), .A1(new_n2977_), .B0(new_n1889_), .B1(new_n1126_), .Y(new_n2978_));
  OAI21X1  g02914(.A0(new_n1885_), .A1(new_n1189_), .B0(new_n2978_), .Y(new_n2979_));
  AOI21X1  g02915(.A0(new_n2976_), .A1(new_n407_), .B0(new_n2979_), .Y(new_n2980_));
  NOR2X1   g02916(.A(new_n2980_), .B(new_n2975_), .Y(new_n2981_));
  INVX1    g02917(.A(new_n2935_), .Y(new_n2982_));
  OAI22X1  g02918(.A0(new_n152_), .A1(new_n105_), .B0(new_n148_), .B1(new_n90_), .Y(new_n2983_));
  OR2X1    g02919(.A(new_n2983_), .B(new_n459_), .Y(new_n2984_));
  OR4X1    g02920(.A(new_n565_), .B(new_n423_), .C(new_n522_), .D(new_n175_), .Y(new_n2985_));
  OR4X1    g02921(.A(new_n329_), .B(new_n194_), .C(new_n147_), .D(new_n338_), .Y(new_n2986_));
  OR4X1    g02922(.A(new_n2986_), .B(new_n2985_), .C(new_n2984_), .D(new_n816_), .Y(new_n2987_));
  OAI22X1  g02923(.A0(new_n152_), .A1(new_n127_), .B0(new_n96_), .B1(new_n94_), .Y(new_n2988_));
  OR4X1    g02924(.A(new_n2988_), .B(new_n272_), .C(new_n155_), .D(new_n120_), .Y(new_n2989_));
  OR4X1    g02925(.A(new_n199_), .B(new_n160_), .C(new_n141_), .D(new_n118_), .Y(new_n2990_));
  OR4X1    g02926(.A(new_n2990_), .B(new_n2989_), .C(new_n1639_), .D(new_n1385_), .Y(new_n2991_));
  OR4X1    g02927(.A(new_n2991_), .B(new_n2987_), .C(new_n2223_), .D(new_n1209_), .Y(new_n2992_));
  NOR3X1   g02928(.A(new_n2992_), .B(new_n1204_), .C(new_n727_), .Y(new_n2993_));
  NOR2X1   g02929(.A(new_n2993_), .B(new_n2982_), .Y(new_n2994_));
  INVX1    g02930(.A(\a[8] ), .Y(new_n2995_));
  INVX1    g02931(.A(new_n541_), .Y(new_n2996_));
  NAND3X1  g02932(.A(new_n2996_), .B(new_n862_), .C(new_n1710_), .Y(new_n2997_));
  OR4X1    g02933(.A(new_n2997_), .B(new_n1599_), .C(new_n259_), .D(new_n181_), .Y(new_n2998_));
  OAI22X1  g02934(.A0(new_n117_), .A1(new_n92_), .B0(new_n81_), .B1(new_n69_), .Y(new_n2999_));
  OR4X1    g02935(.A(new_n293_), .B(new_n252_), .C(new_n457_), .D(new_n521_), .Y(new_n3000_));
  OR4X1    g02936(.A(new_n3000_), .B(new_n2999_), .C(new_n2998_), .D(new_n1335_), .Y(new_n3001_));
  OR4X1    g02937(.A(new_n1438_), .B(new_n1269_), .C(new_n702_), .D(new_n483_), .Y(new_n3002_));
  OR4X1    g02938(.A(new_n3002_), .B(new_n589_), .C(new_n612_), .D(new_n475_), .Y(new_n3003_));
  NOR3X1   g02939(.A(new_n1752_), .B(new_n1114_), .C(new_n921_), .Y(new_n3004_));
  NOR4X1   g02940(.A(new_n815_), .B(new_n565_), .C(new_n757_), .D(new_n585_), .Y(new_n3005_));
  NOR4X1   g02941(.A(new_n586_), .B(new_n494_), .C(new_n220_), .D(new_n1046_), .Y(new_n3006_));
  NAND3X1  g02942(.A(new_n3006_), .B(new_n3005_), .C(new_n3004_), .Y(new_n3007_));
  NOR2X1   g02943(.A(new_n659_), .B(new_n309_), .Y(new_n3008_));
  NOR3X1   g02944(.A(new_n634_), .B(new_n523_), .C(new_n681_), .Y(new_n3009_));
  NAND3X1  g02945(.A(new_n3009_), .B(new_n2942_), .C(new_n3008_), .Y(new_n3010_));
  OR4X1    g02946(.A(new_n3010_), .B(new_n3007_), .C(new_n3003_), .D(new_n3001_), .Y(new_n3011_));
  OR4X1    g02947(.A(new_n460_), .B(new_n998_), .C(new_n243_), .D(new_n133_), .Y(new_n3012_));
  OR4X1    g02948(.A(new_n509_), .B(new_n480_), .C(new_n350_), .D(new_n239_), .Y(new_n3013_));
  OR4X1    g02949(.A(new_n1962_), .B(new_n787_), .C(new_n869_), .D(new_n177_), .Y(new_n3014_));
  OR4X1    g02950(.A(new_n968_), .B(new_n493_), .C(new_n234_), .D(new_n758_), .Y(new_n3015_));
  OR4X1    g02951(.A(new_n3015_), .B(new_n3014_), .C(new_n441_), .D(new_n568_), .Y(new_n3016_));
  OR4X1    g02952(.A(new_n3016_), .B(new_n3013_), .C(new_n3012_), .D(new_n1522_), .Y(new_n3017_));
  OR4X1    g02953(.A(new_n3017_), .B(new_n2586_), .C(new_n403_), .D(new_n378_), .Y(new_n3018_));
  NOR2X1   g02954(.A(new_n3018_), .B(new_n3011_), .Y(new_n3019_));
  OAI22X1  g02955(.A0(new_n92_), .A1(new_n84_), .B0(new_n91_), .B1(new_n90_), .Y(new_n3020_));
  OR4X1    g02956(.A(new_n3020_), .B(new_n2815_), .C(new_n823_), .D(new_n659_), .Y(new_n3021_));
  OR4X1    g02957(.A(new_n1540_), .B(new_n1224_), .C(new_n657_), .D(new_n375_), .Y(new_n3022_));
  OR2X1    g02958(.A(new_n3022_), .B(new_n2019_), .Y(new_n3023_));
  NOR3X1   g02959(.A(new_n1909_), .B(new_n1600_), .C(new_n1415_), .Y(new_n3024_));
  NOR4X1   g02960(.A(new_n422_), .B(new_n391_), .C(new_n603_), .D(new_n806_), .Y(new_n3025_));
  NOR4X1   g02961(.A(new_n261_), .B(new_n245_), .C(new_n149_), .D(new_n120_), .Y(new_n3026_));
  NAND3X1  g02962(.A(new_n3026_), .B(new_n3025_), .C(new_n3024_), .Y(new_n3027_));
  OR4X1    g02963(.A(new_n1028_), .B(new_n632_), .C(new_n1398_), .D(new_n285_), .Y(new_n3028_));
  OR4X1    g02964(.A(new_n578_), .B(new_n176_), .C(new_n86_), .D(new_n85_), .Y(new_n3029_));
  OR4X1    g02965(.A(new_n523_), .B(new_n968_), .C(new_n522_), .D(new_n581_), .Y(new_n3030_));
  OR4X1    g02966(.A(new_n3030_), .B(new_n3029_), .C(new_n3028_), .D(new_n842_), .Y(new_n3031_));
  NOR4X1   g02967(.A(new_n3031_), .B(new_n3027_), .C(new_n3023_), .D(new_n3021_), .Y(new_n3032_));
  INVX1    g02968(.A(new_n3032_), .Y(new_n3033_));
  INVX1    g02969(.A(new_n1688_), .Y(new_n3034_));
  OR4X1    g02970(.A(new_n510_), .B(new_n296_), .C(new_n139_), .D(new_n521_), .Y(new_n3035_));
  OR4X1    g02971(.A(new_n3035_), .B(new_n332_), .C(new_n246_), .D(new_n199_), .Y(new_n3036_));
  OR4X1    g02972(.A(new_n1205_), .B(new_n666_), .C(new_n490_), .D(new_n463_), .Y(new_n3037_));
  OR4X1    g02973(.A(new_n3037_), .B(new_n3036_), .C(new_n2018_), .D(new_n3034_), .Y(new_n3038_));
  NOR4X1   g02974(.A(new_n1635_), .B(new_n1191_), .C(new_n904_), .D(new_n641_), .Y(new_n3039_));
  NOR3X1   g02975(.A(new_n500_), .B(new_n496_), .C(new_n679_), .Y(new_n3040_));
  NOR4X1   g02976(.A(new_n372_), .B(new_n998_), .C(new_n300_), .D(new_n177_), .Y(new_n3041_));
  NAND3X1  g02977(.A(new_n3041_), .B(new_n3040_), .C(new_n3039_), .Y(new_n3042_));
  OR4X1    g02978(.A(new_n497_), .B(new_n717_), .C(new_n263_), .D(new_n757_), .Y(new_n3043_));
  OR4X1    g02979(.A(new_n229_), .B(new_n213_), .C(new_n193_), .D(new_n307_), .Y(new_n3044_));
  OR4X1    g02980(.A(new_n3044_), .B(new_n3043_), .C(new_n226_), .D(new_n379_), .Y(new_n3045_));
  OR4X1    g02981(.A(new_n3045_), .B(new_n3042_), .C(new_n3038_), .D(new_n2013_), .Y(new_n3046_));
  NOR2X1   g02982(.A(new_n3046_), .B(new_n3033_), .Y(new_n3047_));
  NOR2X1   g02983(.A(new_n3047_), .B(new_n3019_), .Y(new_n3048_));
  OR4X1    g02984(.A(new_n3046_), .B(new_n3033_), .C(new_n3018_), .D(new_n3011_), .Y(new_n3049_));
  AOI21X1  g02985(.A0(new_n3049_), .A1(new_n2995_), .B0(new_n3048_), .Y(new_n3050_));
  NOR2X1   g02986(.A(new_n3050_), .B(new_n2982_), .Y(new_n3051_));
  INVX1    g02987(.A(new_n1815_), .Y(new_n3052_));
  XOR2X1   g02988(.A(new_n3052_), .B(new_n1814_), .Y(new_n3053_));
  INVX1    g02989(.A(new_n3053_), .Y(new_n3054_));
  INVX1    g02990(.A(new_n1339_), .Y(new_n3055_));
  AOI22X1  g02991(.A0(new_n1890_), .A1(new_n3055_), .B0(new_n1889_), .B1(new_n2977_), .Y(new_n3056_));
  OAI21X1  g02992(.A0(new_n1885_), .A1(new_n1294_), .B0(new_n3056_), .Y(new_n3057_));
  AOI21X1  g02993(.A0(new_n3054_), .A1(new_n407_), .B0(new_n3057_), .Y(new_n3058_));
  INVX1    g02994(.A(new_n3058_), .Y(new_n3059_));
  XOR2X1   g02995(.A(new_n3050_), .B(new_n2982_), .Y(new_n3060_));
  AOI21X1  g02996(.A0(new_n3060_), .A1(new_n3059_), .B0(new_n3051_), .Y(new_n3061_));
  INVX1    g02997(.A(new_n3061_), .Y(new_n3062_));
  XOR2X1   g02998(.A(new_n2993_), .B(new_n2982_), .Y(new_n3063_));
  AOI21X1  g02999(.A0(new_n3063_), .A1(new_n3062_), .B0(new_n2994_), .Y(new_n3064_));
  INVX1    g03000(.A(new_n3064_), .Y(new_n3065_));
  XOR2X1   g03001(.A(new_n2980_), .B(new_n2975_), .Y(new_n3066_));
  AOI21X1  g03002(.A0(new_n3066_), .A1(new_n3065_), .B0(new_n2981_), .Y(new_n3067_));
  OR2X1    g03003(.A(new_n3067_), .B(new_n2972_), .Y(new_n3068_));
  INVX1    g03004(.A(new_n2972_), .Y(new_n3069_));
  XOR2X1   g03005(.A(new_n3067_), .B(new_n3069_), .Y(new_n3070_));
  OAI22X1  g03006(.A0(new_n2186_), .A1(new_n985_), .B0(new_n2140_), .B1(new_n903_), .Y(new_n3071_));
  AOI21X1  g03007(.A0(new_n2095_), .A1(new_n2835_), .B0(new_n3071_), .Y(new_n3072_));
  OAI21X1  g03008(.A0(new_n2600_), .A1(new_n2063_), .B0(new_n3072_), .Y(new_n3073_));
  XOR2X1   g03009(.A(new_n3073_), .B(new_n74_), .Y(new_n3074_));
  OAI21X1  g03010(.A0(new_n3074_), .A1(new_n3070_), .B0(new_n3068_), .Y(new_n3075_));
  AOI21X1  g03011(.A0(new_n3075_), .A1(new_n2971_), .B0(new_n2970_), .Y(new_n3076_));
  OAI21X1  g03012(.A0(new_n3076_), .A1(new_n2907_), .B0(new_n2905_), .Y(new_n3077_));
  XOR2X1   g03013(.A(new_n2849_), .B(new_n2844_), .Y(new_n3078_));
  AND2X1   g03014(.A(new_n3078_), .B(new_n3077_), .Y(new_n3079_));
  XOR2X1   g03015(.A(new_n3078_), .B(new_n3077_), .Y(new_n3080_));
  AOI22X1  g03016(.A0(new_n2424_), .A1(new_n1886_), .B0(new_n2423_), .B1(new_n1887_), .Y(new_n3081_));
  OAI21X1  g03017(.A0(new_n2419_), .A1(new_n520_), .B0(new_n3081_), .Y(new_n3082_));
  AOI21X1  g03018(.A0(new_n2301_), .A1(new_n1882_), .B0(new_n3082_), .Y(new_n3083_));
  XOR2X1   g03019(.A(new_n3083_), .B(new_n89_), .Y(new_n3084_));
  AOI21X1  g03020(.A0(new_n3084_), .A1(new_n3080_), .B0(new_n3079_), .Y(new_n3085_));
  NOR2X1   g03021(.A(new_n3085_), .B(new_n2898_), .Y(new_n3086_));
  XOR2X1   g03022(.A(new_n3085_), .B(new_n2898_), .Y(new_n3087_));
  AOI22X1  g03023(.A0(new_n2745_), .A1(new_n2627_), .B0(new_n2657_), .B1(new_n2093_), .Y(new_n3088_));
  OAI21X1  g03024(.A0(new_n2743_), .A1(new_n2137_), .B0(new_n3088_), .Y(new_n3089_));
  AOI21X1  g03025(.A0(new_n2658_), .A1(new_n2294_), .B0(new_n3089_), .Y(new_n3090_));
  XOR2X1   g03026(.A(new_n3090_), .B(new_n70_), .Y(new_n3091_));
  AOI21X1  g03027(.A0(new_n3091_), .A1(new_n3087_), .B0(new_n3086_), .Y(new_n3092_));
  NOR2X1   g03028(.A(new_n3092_), .B(new_n2897_), .Y(new_n3093_));
  AOI21X1  g03029(.A0(new_n2896_), .A1(new_n2895_), .B0(new_n3093_), .Y(new_n3094_));
  OR2X1    g03030(.A(new_n3094_), .B(new_n2890_), .Y(new_n3095_));
  XOR2X1   g03031(.A(new_n3094_), .B(new_n2890_), .Y(new_n3096_));
  INVX1    g03032(.A(new_n3096_), .Y(new_n3097_));
  INVX1    g03033(.A(new_n2876_), .Y(new_n3098_));
  AND2X1   g03034(.A(new_n2873_), .B(new_n2869_), .Y(new_n3099_));
  AOI22X1  g03035(.A0(new_n3099_), .A1(new_n2649_), .B0(new_n2875_), .B1(new_n2421_), .Y(new_n3100_));
  OAI21X1  g03036(.A0(new_n3098_), .A1(new_n2695_), .B0(new_n3100_), .Y(new_n3101_));
  XOR2X1   g03037(.A(new_n3101_), .B(new_n1920_), .Y(new_n3102_));
  OR2X1    g03038(.A(new_n3102_), .B(new_n3097_), .Y(new_n3103_));
  AOI21X1  g03039(.A0(new_n3103_), .A1(new_n3095_), .B0(new_n2888_), .Y(new_n3104_));
  INVX1    g03040(.A(new_n2888_), .Y(new_n3105_));
  OAI21X1  g03041(.A0(new_n3102_), .A1(new_n3097_), .B0(new_n3095_), .Y(new_n3106_));
  XOR2X1   g03042(.A(new_n3106_), .B(new_n3105_), .Y(new_n3107_));
  XOR2X1   g03043(.A(new_n3102_), .B(new_n3096_), .Y(new_n3108_));
  XOR2X1   g03044(.A(new_n3091_), .B(new_n3087_), .Y(new_n3109_));
  INVX1    g03045(.A(new_n3109_), .Y(new_n3110_));
  XOR2X1   g03046(.A(new_n3083_), .B(\a[26] ), .Y(new_n3111_));
  XOR2X1   g03047(.A(new_n3111_), .B(new_n3080_), .Y(new_n3112_));
  XOR2X1   g03048(.A(new_n3076_), .B(new_n2906_), .Y(new_n3113_));
  INVX1    g03049(.A(new_n2047_), .Y(new_n3114_));
  OAI22X1  g03050(.A0(new_n2666_), .A1(new_n690_), .B0(new_n2626_), .B1(new_n520_), .Y(new_n3115_));
  AOI21X1  g03051(.A0(new_n2418_), .A1(new_n1886_), .B0(new_n3115_), .Y(new_n3116_));
  OAI21X1  g03052(.A0(new_n2665_), .A1(new_n3114_), .B0(new_n3116_), .Y(new_n3117_));
  XOR2X1   g03053(.A(new_n3117_), .B(new_n89_), .Y(new_n3118_));
  NOR2X1   g03054(.A(new_n3118_), .B(new_n3113_), .Y(new_n3119_));
  INVX1    g03055(.A(new_n2971_), .Y(new_n3120_));
  XOR2X1   g03056(.A(new_n3075_), .B(new_n3120_), .Y(new_n3121_));
  OAI22X1  g03057(.A0(new_n2186_), .A1(new_n957_), .B0(new_n2140_), .B1(new_n847_), .Y(new_n3122_));
  AOI21X1  g03058(.A0(new_n2095_), .A1(new_n2602_), .B0(new_n3122_), .Y(new_n3123_));
  OAI21X1  g03059(.A0(new_n2708_), .A1(new_n2063_), .B0(new_n3123_), .Y(new_n3124_));
  XOR2X1   g03060(.A(new_n3124_), .B(new_n74_), .Y(new_n3125_));
  OR2X1    g03061(.A(new_n3125_), .B(new_n3121_), .Y(new_n3126_));
  AOI22X1  g03062(.A0(new_n2424_), .A1(new_n2036_), .B0(new_n2423_), .B1(new_n1886_), .Y(new_n3127_));
  OAI21X1  g03063(.A0(new_n2419_), .A1(new_n690_), .B0(new_n3127_), .Y(new_n3128_));
  AOI21X1  g03064(.A0(new_n2301_), .A1(new_n2035_), .B0(new_n3128_), .Y(new_n3129_));
  XOR2X1   g03065(.A(new_n3129_), .B(\a[26] ), .Y(new_n3130_));
  AND2X1   g03066(.A(new_n3125_), .B(new_n3121_), .Y(new_n3131_));
  OAI21X1  g03067(.A0(new_n3131_), .A1(new_n3130_), .B0(new_n3126_), .Y(new_n3132_));
  XOR2X1   g03068(.A(new_n3118_), .B(new_n3113_), .Y(new_n3133_));
  AOI21X1  g03069(.A0(new_n3133_), .A1(new_n3132_), .B0(new_n3119_), .Y(new_n3134_));
  NOR2X1   g03070(.A(new_n3134_), .B(new_n3112_), .Y(new_n3135_));
  XOR2X1   g03071(.A(new_n3134_), .B(new_n3112_), .Y(new_n3136_));
  AOI22X1  g03072(.A0(new_n2745_), .A1(new_n2252_), .B0(new_n2657_), .B1(new_n2246_), .Y(new_n3137_));
  OAI21X1  g03073(.A0(new_n2743_), .A1(new_n2092_), .B0(new_n3137_), .Y(new_n3138_));
  AOI21X1  g03074(.A0(new_n2658_), .A1(new_n2201_), .B0(new_n3138_), .Y(new_n3139_));
  XOR2X1   g03075(.A(new_n3139_), .B(new_n70_), .Y(new_n3140_));
  AOI21X1  g03076(.A0(new_n3140_), .A1(new_n3136_), .B0(new_n3135_), .Y(new_n3141_));
  NOR2X1   g03077(.A(new_n3141_), .B(new_n3110_), .Y(new_n3142_));
  XOR2X1   g03078(.A(new_n3141_), .B(new_n3110_), .Y(new_n3143_));
  INVX1    g03079(.A(new_n3099_), .Y(new_n3144_));
  INVX1    g03080(.A(new_n2874_), .Y(new_n3145_));
  NOR2X1   g03081(.A(new_n3145_), .B(new_n2869_), .Y(new_n3146_));
  AOI22X1  g03082(.A0(new_n3146_), .A1(new_n2421_), .B0(new_n2875_), .B1(new_n2420_), .Y(new_n3147_));
  OAI21X1  g03083(.A0(new_n3144_), .A1(new_n2379_), .B0(new_n3147_), .Y(new_n3148_));
  AOI21X1  g03084(.A0(new_n2876_), .A1(new_n2416_), .B0(new_n3148_), .Y(new_n3149_));
  XOR2X1   g03085(.A(new_n3149_), .B(new_n1920_), .Y(new_n3150_));
  AOI21X1  g03086(.A0(new_n3150_), .A1(new_n3143_), .B0(new_n3142_), .Y(new_n3151_));
  INVX1    g03087(.A(new_n3146_), .Y(new_n3152_));
  OAI22X1  g03088(.A0(new_n3152_), .A1(new_n2648_), .B0(new_n3144_), .B1(new_n2414_), .Y(new_n3153_));
  AOI21X1  g03089(.A0(new_n2875_), .A1(new_n2752_), .B0(new_n3153_), .Y(new_n3154_));
  OAI21X1  g03090(.A0(new_n3098_), .A1(new_n2757_), .B0(new_n3154_), .Y(new_n3155_));
  XOR2X1   g03091(.A(new_n3155_), .B(new_n1920_), .Y(new_n3156_));
  NOR2X1   g03092(.A(new_n3156_), .B(new_n3151_), .Y(new_n3157_));
  XOR2X1   g03093(.A(new_n3092_), .B(new_n2897_), .Y(new_n3158_));
  XOR2X1   g03094(.A(new_n3156_), .B(new_n3151_), .Y(new_n3159_));
  AOI21X1  g03095(.A0(new_n3159_), .A1(new_n3158_), .B0(new_n3157_), .Y(new_n3160_));
  NOR2X1   g03096(.A(new_n3160_), .B(new_n3108_), .Y(new_n3161_));
  INVX1    g03097(.A(new_n3161_), .Y(new_n3162_));
  XOR2X1   g03098(.A(new_n3160_), .B(new_n3108_), .Y(new_n3163_));
  INVX1    g03099(.A(new_n3163_), .Y(new_n3164_));
  XOR2X1   g03100(.A(new_n3140_), .B(new_n3136_), .Y(new_n3165_));
  INVX1    g03101(.A(new_n3165_), .Y(new_n3166_));
  AOI22X1  g03102(.A0(new_n2745_), .A1(new_n2093_), .B0(new_n2657_), .B1(new_n1887_), .Y(new_n3167_));
  OAI21X1  g03103(.A0(new_n2743_), .A1(new_n2183_), .B0(new_n3167_), .Y(new_n3168_));
  AOI21X1  g03104(.A0(new_n2658_), .A1(new_n2430_), .B0(new_n3168_), .Y(new_n3169_));
  XOR2X1   g03105(.A(new_n3169_), .B(\a[23] ), .Y(new_n3170_));
  INVX1    g03106(.A(new_n3170_), .Y(new_n3171_));
  XOR2X1   g03107(.A(new_n3133_), .B(new_n3132_), .Y(new_n3172_));
  XOR2X1   g03108(.A(new_n3172_), .B(new_n3170_), .Y(new_n3173_));
  XOR2X1   g03109(.A(new_n3125_), .B(new_n3121_), .Y(new_n3174_));
  XOR2X1   g03110(.A(new_n3174_), .B(new_n3130_), .Y(new_n3175_));
  NOR4X1   g03111(.A(new_n2992_), .B(new_n2935_), .C(new_n1204_), .D(new_n727_), .Y(new_n3176_));
  OAI22X1  g03112(.A0(new_n3065_), .A1(new_n3176_), .B0(new_n3063_), .B1(new_n3061_), .Y(new_n3177_));
  INVX1    g03113(.A(new_n407_), .Y(new_n3178_));
  AOI21X1  g03114(.A0(new_n1815_), .A1(new_n1814_), .B0(new_n1295_), .Y(new_n3179_));
  XOR2X1   g03115(.A(new_n1817_), .B(new_n3179_), .Y(new_n3180_));
  NOR2X1   g03116(.A(new_n3180_), .B(new_n3178_), .Y(new_n3181_));
  AOI22X1  g03117(.A0(new_n1889_), .A1(new_n1187_), .B0(new_n1884_), .B1(new_n2977_), .Y(new_n3182_));
  OAI21X1  g03118(.A0(new_n2245_), .A1(new_n1294_), .B0(new_n3182_), .Y(new_n3183_));
  OAI21X1  g03119(.A0(new_n3183_), .A1(new_n3181_), .B0(new_n3177_), .Y(new_n3184_));
  AOI22X1  g03120(.A0(new_n2185_), .A1(new_n1126_), .B0(new_n2139_), .B1(new_n2603_), .Y(new_n3185_));
  OAI21X1  g03121(.A0(new_n2431_), .A1(new_n1065_), .B0(new_n3185_), .Y(new_n3186_));
  AOI21X1  g03122(.A0(new_n2824_), .A1(new_n2062_), .B0(new_n3186_), .Y(new_n3187_));
  XOR2X1   g03123(.A(new_n3187_), .B(\a[29] ), .Y(new_n3188_));
  INVX1    g03124(.A(new_n3180_), .Y(new_n3189_));
  AOI21X1  g03125(.A0(new_n3189_), .A1(new_n407_), .B0(new_n3183_), .Y(new_n3190_));
  XOR2X1   g03126(.A(new_n3190_), .B(new_n3177_), .Y(new_n3191_));
  OAI21X1  g03127(.A0(new_n3191_), .A1(new_n3188_), .B0(new_n3184_), .Y(new_n3192_));
  XOR2X1   g03128(.A(new_n3066_), .B(new_n3065_), .Y(new_n3193_));
  AND2X1   g03129(.A(new_n3193_), .B(new_n3192_), .Y(new_n3194_));
  AOI22X1  g03130(.A0(new_n2139_), .A1(new_n2835_), .B0(new_n2095_), .B1(new_n2603_), .Y(new_n3195_));
  OAI21X1  g03131(.A0(new_n2186_), .A1(new_n1065_), .B0(new_n3195_), .Y(new_n3196_));
  AOI21X1  g03132(.A0(new_n2834_), .A1(new_n2062_), .B0(new_n3196_), .Y(new_n3197_));
  XOR2X1   g03133(.A(new_n3197_), .B(\a[29] ), .Y(new_n3198_));
  INVX1    g03134(.A(new_n3198_), .Y(new_n3199_));
  XOR2X1   g03135(.A(new_n3193_), .B(new_n3192_), .Y(new_n3200_));
  AOI21X1  g03136(.A0(new_n3200_), .A1(new_n3199_), .B0(new_n3194_), .Y(new_n3201_));
  INVX1    g03137(.A(new_n3201_), .Y(new_n3202_));
  XOR2X1   g03138(.A(new_n3074_), .B(new_n3070_), .Y(new_n3203_));
  AND2X1   g03139(.A(new_n3203_), .B(new_n3202_), .Y(new_n3204_));
  XOR2X1   g03140(.A(new_n3203_), .B(new_n3202_), .Y(new_n3205_));
  AOI22X1  g03141(.A0(new_n2424_), .A1(new_n2481_), .B0(new_n2423_), .B1(new_n2049_), .Y(new_n3206_));
  OAI21X1  g03142(.A0(new_n2419_), .A1(new_n783_), .B0(new_n3206_), .Y(new_n3207_));
  AOI21X1  g03143(.A0(new_n2480_), .A1(new_n2301_), .B0(new_n3207_), .Y(new_n3208_));
  XOR2X1   g03144(.A(new_n3208_), .B(new_n89_), .Y(new_n3209_));
  AOI21X1  g03145(.A0(new_n3209_), .A1(new_n3205_), .B0(new_n3204_), .Y(new_n3210_));
  NOR2X1   g03146(.A(new_n3210_), .B(new_n3175_), .Y(new_n3211_));
  XOR2X1   g03147(.A(new_n3210_), .B(new_n3175_), .Y(new_n3212_));
  AOI22X1  g03148(.A0(new_n2745_), .A1(new_n2246_), .B0(new_n2657_), .B1(new_n2048_), .Y(new_n3213_));
  OAI21X1  g03149(.A0(new_n2743_), .A1(new_n1879_), .B0(new_n3213_), .Y(new_n3214_));
  AOI21X1  g03150(.A0(new_n2658_), .A1(new_n2244_), .B0(new_n3214_), .Y(new_n3215_));
  XOR2X1   g03151(.A(new_n3215_), .B(new_n70_), .Y(new_n3216_));
  AOI21X1  g03152(.A0(new_n3216_), .A1(new_n3212_), .B0(new_n3211_), .Y(new_n3217_));
  NOR2X1   g03153(.A(new_n3217_), .B(new_n3173_), .Y(new_n3218_));
  AOI21X1  g03154(.A0(new_n3172_), .A1(new_n3171_), .B0(new_n3218_), .Y(new_n3219_));
  NOR2X1   g03155(.A(new_n3219_), .B(new_n3166_), .Y(new_n3220_));
  XOR2X1   g03156(.A(new_n3219_), .B(new_n3166_), .Y(new_n3221_));
  AOI22X1  g03157(.A0(new_n3099_), .A1(new_n2420_), .B0(new_n2875_), .B1(new_n2627_), .Y(new_n3222_));
  OAI21X1  g03158(.A0(new_n3152_), .A1(new_n2379_), .B0(new_n3222_), .Y(new_n3223_));
  AOI21X1  g03159(.A0(new_n2876_), .A1(new_n2625_), .B0(new_n3223_), .Y(new_n3224_));
  XOR2X1   g03160(.A(new_n3224_), .B(new_n1920_), .Y(new_n3225_));
  AOI21X1  g03161(.A0(new_n3225_), .A1(new_n3221_), .B0(new_n3220_), .Y(new_n3226_));
  XOR2X1   g03162(.A(\a[17] ), .B(\a[16] ), .Y(new_n3227_));
  XOR2X1   g03163(.A(\a[16] ), .B(\a[15] ), .Y(new_n3228_));
  INVX1    g03164(.A(new_n3228_), .Y(new_n3229_));
  XOR2X1   g03165(.A(\a[15] ), .B(new_n2529_), .Y(new_n3230_));
  NAND3X1  g03166(.A(new_n3230_), .B(new_n3229_), .C(new_n3227_), .Y(new_n3231_));
  INVX1    g03167(.A(new_n3231_), .Y(new_n3232_));
  INVX1    g03168(.A(new_n3227_), .Y(new_n3233_));
  NOR2X1   g03169(.A(new_n3230_), .B(new_n3233_), .Y(new_n3234_));
  AOI22X1  g03170(.A0(new_n3234_), .A1(new_n2652_), .B0(new_n3232_), .B1(new_n2649_), .Y(new_n3235_));
  XOR2X1   g03171(.A(new_n3235_), .B(\a[17] ), .Y(new_n3236_));
  NOR2X1   g03172(.A(new_n3236_), .B(new_n3226_), .Y(new_n3237_));
  XOR2X1   g03173(.A(new_n3150_), .B(new_n3143_), .Y(new_n3238_));
  XOR2X1   g03174(.A(new_n3236_), .B(new_n3226_), .Y(new_n3239_));
  AOI21X1  g03175(.A0(new_n3239_), .A1(new_n3238_), .B0(new_n3237_), .Y(new_n3240_));
  INVX1    g03176(.A(new_n3240_), .Y(new_n3241_));
  XOR2X1   g03177(.A(new_n3159_), .B(new_n3158_), .Y(new_n3242_));
  AND2X1   g03178(.A(new_n3242_), .B(new_n3241_), .Y(new_n3243_));
  XOR2X1   g03179(.A(new_n3239_), .B(new_n3238_), .Y(new_n3244_));
  INVX1    g03180(.A(new_n3244_), .Y(new_n3245_));
  XOR2X1   g03181(.A(new_n3225_), .B(new_n3221_), .Y(new_n3246_));
  INVX1    g03182(.A(new_n3246_), .Y(new_n3247_));
  INVX1    g03183(.A(new_n3173_), .Y(new_n3248_));
  XOR2X1   g03184(.A(new_n3217_), .B(new_n3248_), .Y(new_n3249_));
  INVX1    g03185(.A(new_n2875_), .Y(new_n3250_));
  OAI22X1  g03186(.A0(new_n3152_), .A1(new_n2339_), .B0(new_n3250_), .B1(new_n2137_), .Y(new_n3251_));
  AOI21X1  g03187(.A0(new_n3099_), .A1(new_n2627_), .B0(new_n3251_), .Y(new_n3252_));
  OAI21X1  g03188(.A0(new_n3098_), .A1(new_n2670_), .B0(new_n3252_), .Y(new_n3253_));
  XOR2X1   g03189(.A(new_n3253_), .B(new_n1920_), .Y(new_n3254_));
  NOR2X1   g03190(.A(new_n3254_), .B(new_n3249_), .Y(new_n3255_));
  XOR2X1   g03191(.A(new_n3216_), .B(new_n3212_), .Y(new_n3256_));
  INVX1    g03192(.A(new_n3256_), .Y(new_n3257_));
  XOR2X1   g03193(.A(new_n3208_), .B(\a[26] ), .Y(new_n3258_));
  XOR2X1   g03194(.A(new_n3258_), .B(new_n3205_), .Y(new_n3259_));
  XOR2X1   g03195(.A(new_n3200_), .B(new_n3198_), .Y(new_n3260_));
  INVX1    g03196(.A(new_n2494_), .Y(new_n3261_));
  OAI22X1  g03197(.A0(new_n2666_), .A1(new_n903_), .B0(new_n2626_), .B1(new_n783_), .Y(new_n3262_));
  AOI21X1  g03198(.A0(new_n2418_), .A1(new_n2481_), .B0(new_n3262_), .Y(new_n3263_));
  OAI21X1  g03199(.A0(new_n3261_), .A1(new_n2665_), .B0(new_n3263_), .Y(new_n3264_));
  XOR2X1   g03200(.A(new_n3264_), .B(new_n89_), .Y(new_n3265_));
  NOR2X1   g03201(.A(new_n3265_), .B(new_n3260_), .Y(new_n3266_));
  XOR2X1   g03202(.A(new_n3191_), .B(new_n3188_), .Y(new_n3267_));
  INVX1    g03203(.A(new_n3267_), .Y(new_n3268_));
  XOR2X1   g03204(.A(new_n3060_), .B(new_n3058_), .Y(new_n3269_));
  NOR2X1   g03205(.A(new_n3048_), .B(\a[8] ), .Y(new_n3270_));
  AOI21X1  g03206(.A0(new_n3270_), .A1(new_n3049_), .B0(\a[8] ), .Y(new_n3271_));
  AOI21X1  g03207(.A0(new_n3050_), .A1(new_n3049_), .B0(new_n3271_), .Y(new_n3272_));
  NOR3X1   g03208(.A(new_n547_), .B(new_n998_), .C(new_n149_), .Y(new_n3273_));
  NOR4X1   g03209(.A(new_n594_), .B(new_n579_), .C(new_n412_), .D(new_n540_), .Y(new_n3274_));
  NOR4X1   g03210(.A(new_n356_), .B(new_n197_), .C(new_n792_), .D(new_n120_), .Y(new_n3275_));
  NAND3X1  g03211(.A(new_n3275_), .B(new_n3274_), .C(new_n3273_), .Y(new_n3276_));
  OR4X1    g03212(.A(new_n638_), .B(new_n803_), .C(new_n464_), .D(new_n312_), .Y(new_n3277_));
  OR4X1    g03213(.A(new_n3277_), .B(new_n3276_), .C(new_n3021_), .D(new_n3003_), .Y(new_n3278_));
  OR4X1    g03214(.A(new_n393_), .B(new_n391_), .C(new_n806_), .D(new_n141_), .Y(new_n3279_));
  OR4X1    g03215(.A(new_n3279_), .B(new_n536_), .C(new_n981_), .D(new_n93_), .Y(new_n3280_));
  NAND2X1  g03216(.A(new_n2234_), .B(new_n2080_), .Y(new_n3281_));
  OR4X1    g03217(.A(new_n1002_), .B(new_n510_), .C(new_n429_), .D(new_n372_), .Y(new_n3282_));
  OAI22X1  g03218(.A0(new_n161_), .A1(new_n79_), .B0(new_n119_), .B1(new_n105_), .Y(new_n3283_));
  OR4X1    g03219(.A(new_n3283_), .B(new_n1224_), .C(new_n414_), .D(new_n299_), .Y(new_n3284_));
  OR4X1    g03220(.A(new_n3284_), .B(new_n3282_), .C(new_n3281_), .D(new_n3280_), .Y(new_n3285_));
  NOR4X1   g03221(.A(new_n3285_), .B(new_n3278_), .C(new_n1958_), .D(new_n736_), .Y(new_n3286_));
  NOR3X1   g03222(.A(new_n3286_), .B(new_n3018_), .C(new_n3011_), .Y(new_n3287_));
  INVX1    g03223(.A(new_n3019_), .Y(new_n3288_));
  INVX1    g03224(.A(\a[5] ), .Y(new_n3289_));
  NAND3X1  g03225(.A(new_n988_), .B(new_n2150_), .C(new_n807_), .Y(new_n3290_));
  OR4X1    g03226(.A(new_n998_), .B(new_n183_), .C(new_n172_), .D(new_n147_), .Y(new_n3291_));
  OAI22X1  g03227(.A0(new_n148_), .A1(new_n125_), .B0(new_n131_), .B1(new_n79_), .Y(new_n3292_));
  NOR2X1   g03228(.A(new_n3292_), .B(new_n631_), .Y(new_n3293_));
  INVX1    g03229(.A(new_n3293_), .Y(new_n3294_));
  INVX1    g03230(.A(new_n304_), .Y(new_n3295_));
  INVX1    g03231(.A(new_n460_), .Y(new_n3296_));
  NAND3X1  g03232(.A(new_n3296_), .B(new_n861_), .C(new_n3295_), .Y(new_n3297_));
  OR4X1    g03233(.A(new_n3297_), .B(new_n3294_), .C(new_n3291_), .D(new_n3290_), .Y(new_n3298_));
  AOI21X1  g03234(.A0(new_n127_), .A1(new_n125_), .B0(new_n119_), .Y(new_n3299_));
  OR2X1    g03235(.A(new_n3299_), .B(new_n420_), .Y(new_n3300_));
  OAI22X1  g03236(.A0(new_n182_), .A1(new_n88_), .B0(new_n129_), .B1(new_n69_), .Y(new_n3301_));
  OR4X1    g03237(.A(new_n201_), .B(new_n133_), .C(new_n100_), .D(new_n85_), .Y(new_n3302_));
  OR4X1    g03238(.A(new_n3302_), .B(new_n3301_), .C(new_n3300_), .D(new_n589_), .Y(new_n3303_));
  OAI22X1  g03239(.A0(new_n108_), .A1(new_n75_), .B0(new_n91_), .B1(new_n78_), .Y(new_n3304_));
  OR2X1    g03240(.A(new_n3304_), .B(new_n848_), .Y(new_n3305_));
  OAI22X1  g03241(.A0(new_n168_), .A1(new_n81_), .B0(new_n148_), .B1(new_n131_), .Y(new_n3306_));
  OR4X1    g03242(.A(new_n3306_), .B(new_n3305_), .C(new_n504_), .D(new_n274_), .Y(new_n3307_));
  OR4X1    g03243(.A(new_n1749_), .B(new_n878_), .C(new_n463_), .D(new_n1057_), .Y(new_n3308_));
  OR4X1    g03244(.A(new_n3308_), .B(new_n3307_), .C(new_n3303_), .D(new_n3298_), .Y(new_n3309_));
  OR4X1    g03245(.A(new_n260_), .B(new_n539_), .C(new_n1046_), .D(new_n86_), .Y(new_n3310_));
  OR4X1    g03246(.A(new_n3310_), .B(new_n455_), .C(new_n474_), .D(new_n301_), .Y(new_n3311_));
  OAI22X1  g03247(.A0(new_n143_), .A1(new_n91_), .B0(new_n106_), .B1(new_n78_), .Y(new_n3312_));
  OR2X1    g03248(.A(new_n3312_), .B(new_n391_), .Y(new_n3313_));
  OR4X1    g03249(.A(new_n1701_), .B(new_n582_), .C(new_n648_), .D(new_n338_), .Y(new_n3314_));
  OR2X1    g03250(.A(new_n3314_), .B(new_n1867_), .Y(new_n3315_));
  OR4X1    g03251(.A(new_n3315_), .B(new_n3313_), .C(new_n3311_), .D(new_n686_), .Y(new_n3316_));
  OR4X1    g03252(.A(new_n2178_), .B(new_n1159_), .C(new_n155_), .D(new_n141_), .Y(new_n3317_));
  OR4X1    g03253(.A(new_n3317_), .B(new_n634_), .C(new_n398_), .D(new_n291_), .Y(new_n3318_));
  OR2X1    g03254(.A(new_n3318_), .B(new_n1859_), .Y(new_n3319_));
  NOR4X1   g03255(.A(new_n3319_), .B(new_n3316_), .C(new_n3309_), .D(new_n2571_), .Y(new_n3320_));
  NOR2X1   g03256(.A(new_n3320_), .B(\a[2] ), .Y(new_n3321_));
  XOR2X1   g03257(.A(new_n3320_), .B(\a[2] ), .Y(new_n3322_));
  AOI21X1  g03258(.A0(new_n3322_), .A1(new_n3289_), .B0(new_n3321_), .Y(new_n3323_));
  NOR2X1   g03259(.A(new_n3323_), .B(new_n3288_), .Y(new_n3324_));
  OR2X1    g03260(.A(new_n1807_), .B(new_n1424_), .Y(new_n3325_));
  XOR2X1   g03261(.A(new_n1808_), .B(new_n3325_), .Y(new_n3326_));
  INVX1    g03262(.A(new_n1423_), .Y(new_n3327_));
  AOI22X1  g03263(.A0(new_n1890_), .A1(new_n3327_), .B0(new_n1889_), .B1(new_n1357_), .Y(new_n3328_));
  OAI21X1  g03264(.A0(new_n1885_), .A1(new_n1389_), .B0(new_n3328_), .Y(new_n3329_));
  AOI21X1  g03265(.A0(new_n3326_), .A1(new_n407_), .B0(new_n3329_), .Y(new_n3330_));
  INVX1    g03266(.A(new_n3330_), .Y(new_n3331_));
  XOR2X1   g03267(.A(new_n3323_), .B(new_n3288_), .Y(new_n3332_));
  AOI21X1  g03268(.A0(new_n3332_), .A1(new_n3331_), .B0(new_n3324_), .Y(new_n3333_));
  INVX1    g03269(.A(new_n3333_), .Y(new_n3334_));
  AND2X1   g03270(.A(new_n3286_), .B(new_n3288_), .Y(new_n3335_));
  INVX1    g03271(.A(new_n3335_), .Y(new_n3336_));
  AOI21X1  g03272(.A0(new_n3336_), .A1(new_n3334_), .B0(new_n3287_), .Y(new_n3337_));
  NOR2X1   g03273(.A(new_n3337_), .B(new_n3272_), .Y(new_n3338_));
  XOR2X1   g03274(.A(new_n1339_), .B(new_n1294_), .Y(new_n3339_));
  XOR2X1   g03275(.A(new_n3339_), .B(new_n1812_), .Y(new_n3340_));
  INVX1    g03276(.A(new_n3340_), .Y(new_n3341_));
  INVX1    g03277(.A(new_n1294_), .Y(new_n3342_));
  AOI22X1  g03278(.A0(new_n1890_), .A1(new_n1357_), .B0(new_n1889_), .B1(new_n3342_), .Y(new_n3343_));
  OAI21X1  g03279(.A0(new_n1885_), .A1(new_n1339_), .B0(new_n3343_), .Y(new_n3344_));
  AOI21X1  g03280(.A0(new_n3341_), .A1(new_n407_), .B0(new_n3344_), .Y(new_n3345_));
  INVX1    g03281(.A(new_n3345_), .Y(new_n3346_));
  XOR2X1   g03282(.A(new_n3337_), .B(new_n3272_), .Y(new_n3347_));
  AOI21X1  g03283(.A0(new_n3347_), .A1(new_n3346_), .B0(new_n3338_), .Y(new_n3348_));
  OR2X1    g03284(.A(new_n3348_), .B(new_n3269_), .Y(new_n3349_));
  INVX1    g03285(.A(new_n3269_), .Y(new_n3350_));
  XOR2X1   g03286(.A(new_n3348_), .B(new_n3350_), .Y(new_n3351_));
  INVX1    g03287(.A(new_n2963_), .Y(new_n3352_));
  OAI22X1  g03288(.A0(new_n2140_), .A1(new_n1065_), .B0(new_n2431_), .B1(new_n1127_), .Y(new_n3353_));
  AOI21X1  g03289(.A0(new_n2185_), .A1(new_n1187_), .B0(new_n3353_), .Y(new_n3354_));
  OAI21X1  g03290(.A0(new_n3352_), .A1(new_n2063_), .B0(new_n3354_), .Y(new_n3355_));
  XOR2X1   g03291(.A(new_n3355_), .B(new_n74_), .Y(new_n3356_));
  OR2X1    g03292(.A(new_n3356_), .B(new_n3351_), .Y(new_n3357_));
  AND2X1   g03293(.A(new_n3357_), .B(new_n3349_), .Y(new_n3358_));
  OR2X1    g03294(.A(new_n3358_), .B(new_n3268_), .Y(new_n3359_));
  AND2X1   g03295(.A(new_n3358_), .B(new_n3268_), .Y(new_n3360_));
  AOI22X1  g03296(.A0(new_n2424_), .A1(new_n2835_), .B0(new_n2423_), .B1(new_n2481_), .Y(new_n3361_));
  OAI21X1  g03297(.A0(new_n2419_), .A1(new_n903_), .B0(new_n3361_), .Y(new_n3362_));
  AOI21X1  g03298(.A0(new_n2709_), .A1(new_n2301_), .B0(new_n3362_), .Y(new_n3363_));
  XOR2X1   g03299(.A(new_n3363_), .B(\a[26] ), .Y(new_n3364_));
  OAI21X1  g03300(.A0(new_n3364_), .A1(new_n3360_), .B0(new_n3359_), .Y(new_n3365_));
  XOR2X1   g03301(.A(new_n3265_), .B(new_n3260_), .Y(new_n3366_));
  AOI21X1  g03302(.A0(new_n3366_), .A1(new_n3365_), .B0(new_n3266_), .Y(new_n3367_));
  NOR2X1   g03303(.A(new_n3367_), .B(new_n3259_), .Y(new_n3368_));
  XOR2X1   g03304(.A(new_n3367_), .B(new_n3259_), .Y(new_n3369_));
  AOI22X1  g03305(.A0(new_n2745_), .A1(new_n1887_), .B0(new_n2657_), .B1(new_n1886_), .Y(new_n3370_));
  OAI21X1  g03306(.A0(new_n2743_), .A1(new_n520_), .B0(new_n3370_), .Y(new_n3371_));
  AOI21X1  g03307(.A0(new_n2658_), .A1(new_n1882_), .B0(new_n3371_), .Y(new_n3372_));
  XOR2X1   g03308(.A(new_n3372_), .B(new_n70_), .Y(new_n3373_));
  AOI21X1  g03309(.A0(new_n3373_), .A1(new_n3369_), .B0(new_n3368_), .Y(new_n3374_));
  OR2X1    g03310(.A(new_n3374_), .B(new_n3257_), .Y(new_n3375_));
  XOR2X1   g03311(.A(new_n3374_), .B(new_n3257_), .Y(new_n3376_));
  INVX1    g03312(.A(new_n3376_), .Y(new_n3377_));
  AOI22X1  g03313(.A0(new_n3146_), .A1(new_n2627_), .B0(new_n2875_), .B1(new_n2093_), .Y(new_n3378_));
  OAI21X1  g03314(.A0(new_n3144_), .A1(new_n2137_), .B0(new_n3378_), .Y(new_n3379_));
  AOI21X1  g03315(.A0(new_n2876_), .A1(new_n2294_), .B0(new_n3379_), .Y(new_n3380_));
  XOR2X1   g03316(.A(new_n3380_), .B(\a[20] ), .Y(new_n3381_));
  OAI21X1  g03317(.A0(new_n3381_), .A1(new_n3377_), .B0(new_n3375_), .Y(new_n3382_));
  XOR2X1   g03318(.A(new_n3254_), .B(new_n3249_), .Y(new_n3383_));
  AOI21X1  g03319(.A0(new_n3383_), .A1(new_n3382_), .B0(new_n3255_), .Y(new_n3384_));
  OR2X1    g03320(.A(new_n3384_), .B(new_n3247_), .Y(new_n3385_));
  XOR2X1   g03321(.A(new_n3384_), .B(new_n3247_), .Y(new_n3386_));
  INVX1    g03322(.A(new_n3386_), .Y(new_n3387_));
  INVX1    g03323(.A(new_n3234_), .Y(new_n3388_));
  NAND2X1  g03324(.A(new_n3230_), .B(new_n3228_), .Y(new_n3389_));
  INVX1    g03325(.A(new_n3389_), .Y(new_n3390_));
  AOI22X1  g03326(.A0(new_n3390_), .A1(new_n2649_), .B0(new_n3232_), .B1(new_n2421_), .Y(new_n3391_));
  OAI21X1  g03327(.A0(new_n3388_), .A1(new_n2695_), .B0(new_n3391_), .Y(new_n3392_));
  XOR2X1   g03328(.A(new_n3392_), .B(new_n2445_), .Y(new_n3393_));
  OR2X1    g03329(.A(new_n3393_), .B(new_n3387_), .Y(new_n3394_));
  AOI21X1  g03330(.A0(new_n3394_), .A1(new_n3385_), .B0(new_n3245_), .Y(new_n3395_));
  INVX1    g03331(.A(new_n3395_), .Y(new_n3396_));
  AND2X1   g03332(.A(new_n3394_), .B(new_n3385_), .Y(new_n3397_));
  XOR2X1   g03333(.A(new_n3397_), .B(new_n3245_), .Y(new_n3398_));
  INVX1    g03334(.A(new_n3398_), .Y(new_n3399_));
  XOR2X1   g03335(.A(new_n3393_), .B(new_n3386_), .Y(new_n3400_));
  XOR2X1   g03336(.A(new_n3381_), .B(new_n3376_), .Y(new_n3401_));
  XOR2X1   g03337(.A(new_n3373_), .B(new_n3369_), .Y(new_n3402_));
  INVX1    g03338(.A(new_n3402_), .Y(new_n3403_));
  AOI22X1  g03339(.A0(new_n2745_), .A1(new_n2048_), .B0(new_n2657_), .B1(new_n2049_), .Y(new_n3404_));
  OAI21X1  g03340(.A0(new_n2743_), .A1(new_n623_), .B0(new_n3404_), .Y(new_n3405_));
  AOI21X1  g03341(.A0(new_n2658_), .A1(new_n2047_), .B0(new_n3405_), .Y(new_n3406_));
  XOR2X1   g03342(.A(new_n3406_), .B(\a[23] ), .Y(new_n3407_));
  INVX1    g03343(.A(new_n3407_), .Y(new_n3408_));
  XOR2X1   g03344(.A(new_n3366_), .B(new_n3365_), .Y(new_n3409_));
  XOR2X1   g03345(.A(new_n3409_), .B(new_n3407_), .Y(new_n3410_));
  XOR2X1   g03346(.A(new_n3358_), .B(new_n3268_), .Y(new_n3411_));
  XOR2X1   g03347(.A(new_n3364_), .B(new_n3411_), .Y(new_n3412_));
  AOI22X1  g03348(.A0(new_n2185_), .A1(new_n2977_), .B0(new_n2139_), .B1(new_n1126_), .Y(new_n3413_));
  OAI21X1  g03349(.A0(new_n2431_), .A1(new_n1189_), .B0(new_n3413_), .Y(new_n3414_));
  AOI21X1  g03350(.A0(new_n2976_), .A1(new_n2062_), .B0(new_n3414_), .Y(new_n3415_));
  XOR2X1   g03351(.A(new_n3415_), .B(\a[29] ), .Y(new_n3416_));
  XOR2X1   g03352(.A(new_n3347_), .B(new_n3345_), .Y(new_n3417_));
  NOR2X1   g03353(.A(new_n3417_), .B(new_n3416_), .Y(new_n3418_));
  INVX1    g03354(.A(new_n3418_), .Y(new_n3419_));
  XOR2X1   g03355(.A(new_n3417_), .B(new_n3416_), .Y(new_n3420_));
  INVX1    g03356(.A(new_n3420_), .Y(new_n3421_));
  XOR2X1   g03357(.A(new_n3286_), .B(new_n3288_), .Y(new_n3422_));
  NOR2X1   g03358(.A(new_n3422_), .B(new_n3333_), .Y(new_n3423_));
  AOI21X1  g03359(.A0(new_n3337_), .A1(new_n3336_), .B0(new_n3423_), .Y(new_n3424_));
  XOR2X1   g03360(.A(new_n1811_), .B(new_n1810_), .Y(new_n3425_));
  AOI22X1  g03361(.A0(new_n1889_), .A1(new_n3055_), .B0(new_n1884_), .B1(new_n1357_), .Y(new_n3426_));
  OAI21X1  g03362(.A0(new_n2245_), .A1(new_n1389_), .B0(new_n3426_), .Y(new_n3427_));
  AOI21X1  g03363(.A0(new_n3425_), .A1(new_n407_), .B0(new_n3427_), .Y(new_n3428_));
  OR2X1    g03364(.A(new_n3428_), .B(new_n3424_), .Y(new_n3429_));
  XOR2X1   g03365(.A(new_n3332_), .B(new_n3330_), .Y(new_n3430_));
  INVX1    g03366(.A(\a[2] ), .Y(new_n3431_));
  OR4X1    g03367(.A(new_n422_), .B(new_n227_), .C(new_n379_), .D(new_n337_), .Y(new_n3432_));
  OR4X1    g03368(.A(new_n3432_), .B(new_n547_), .C(new_n385_), .D(new_n357_), .Y(new_n3433_));
  OAI22X1  g03369(.A0(new_n168_), .A1(new_n129_), .B0(new_n117_), .B1(new_n94_), .Y(new_n3434_));
  OR4X1    g03370(.A(new_n2806_), .B(new_n3434_), .C(new_n925_), .D(new_n656_), .Y(new_n3435_));
  OR4X1    g03371(.A(new_n1725_), .B(new_n2157_), .C(new_n1271_), .D(new_n1244_), .Y(new_n3436_));
  OR4X1    g03372(.A(new_n3436_), .B(new_n747_), .C(new_n220_), .D(new_n175_), .Y(new_n3437_));
  INVX1    g03373(.A(new_n855_), .Y(new_n3438_));
  OR4X1    g03374(.A(new_n632_), .B(new_n394_), .C(new_n574_), .D(new_n1046_), .Y(new_n3439_));
  OR4X1    g03375(.A(new_n3439_), .B(new_n2986_), .C(new_n2937_), .D(new_n3438_), .Y(new_n3440_));
  OR4X1    g03376(.A(new_n3440_), .B(new_n3437_), .C(new_n3435_), .D(new_n3433_), .Y(new_n3441_));
  NOR4X1   g03377(.A(new_n3441_), .B(new_n2071_), .C(new_n1603_), .D(new_n1464_), .Y(new_n3442_));
  NOR2X1   g03378(.A(new_n3442_), .B(new_n3431_), .Y(new_n3443_));
  OR4X1    g03379(.A(new_n2795_), .B(new_n1095_), .C(new_n293_), .D(new_n239_), .Y(new_n3444_));
  OR4X1    g03380(.A(new_n667_), .B(new_n656_), .C(new_n480_), .D(new_n356_), .Y(new_n3445_));
  OR4X1    g03381(.A(new_n3445_), .B(new_n3444_), .C(new_n2537_), .D(new_n1851_), .Y(new_n3446_));
  NOR4X1   g03382(.A(new_n553_), .B(new_n285_), .C(new_n249_), .D(new_n296_), .Y(new_n3447_));
  NOR4X1   g03383(.A(new_n938_), .B(new_n724_), .C(new_n594_), .D(new_n543_), .Y(new_n3448_));
  NOR4X1   g03384(.A(new_n394_), .B(new_n383_), .C(new_n354_), .D(new_n843_), .Y(new_n3449_));
  NAND3X1  g03385(.A(new_n3449_), .B(new_n3448_), .C(new_n3447_), .Y(new_n3450_));
  OR4X1    g03386(.A(new_n1082_), .B(new_n385_), .C(new_n365_), .D(new_n233_), .Y(new_n3451_));
  OR4X1    g03387(.A(new_n3451_), .B(new_n561_), .C(new_n194_), .D(new_n187_), .Y(new_n3452_));
  OR4X1    g03388(.A(new_n391_), .B(new_n423_), .C(new_n301_), .D(new_n664_), .Y(new_n3453_));
  OR4X1    g03389(.A(new_n3453_), .B(new_n3452_), .C(new_n3450_), .D(new_n419_), .Y(new_n3454_));
  NOR4X1   g03390(.A(new_n3454_), .B(new_n3446_), .C(new_n518_), .D(new_n167_), .Y(new_n3455_));
  NOR2X1   g03391(.A(new_n3455_), .B(new_n3431_), .Y(new_n3456_));
  OAI22X1  g03392(.A0(new_n168_), .A1(new_n72_), .B0(new_n96_), .B1(new_n90_), .Y(new_n3457_));
  OR4X1    g03393(.A(new_n3457_), .B(new_n1225_), .C(new_n1898_), .D(new_n834_), .Y(new_n3458_));
  OAI22X1  g03394(.A0(new_n152_), .A1(new_n78_), .B0(new_n115_), .B1(new_n72_), .Y(new_n3459_));
  OR2X1    g03395(.A(new_n3459_), .B(new_n720_), .Y(new_n3460_));
  OR4X1    g03396(.A(new_n264_), .B(new_n357_), .C(new_n439_), .D(new_n207_), .Y(new_n3461_));
  OR4X1    g03397(.A(new_n3461_), .B(new_n3460_), .C(new_n3458_), .D(new_n2998_), .Y(new_n3462_));
  OR4X1    g03398(.A(new_n3462_), .B(new_n2985_), .C(new_n3438_), .D(new_n113_), .Y(new_n3463_));
  OR4X1    g03399(.A(new_n385_), .B(new_n885_), .C(new_n202_), .D(new_n184_), .Y(new_n3464_));
  OR4X1    g03400(.A(new_n523_), .B(new_n286_), .C(new_n263_), .D(new_n194_), .Y(new_n3465_));
  OR4X1    g03401(.A(new_n3465_), .B(new_n3464_), .C(new_n1502_), .D(new_n671_), .Y(new_n3466_));
  OR4X1    g03402(.A(new_n478_), .B(new_n251_), .C(new_n224_), .D(new_n208_), .Y(new_n3467_));
  OR4X1    g03403(.A(new_n3467_), .B(new_n724_), .C(new_n1261_), .D(new_n355_), .Y(new_n3468_));
  OR4X1    g03404(.A(new_n2806_), .B(new_n2536_), .C(new_n459_), .D(new_n231_), .Y(new_n3469_));
  OR4X1    g03405(.A(new_n500_), .B(new_n815_), .C(new_n240_), .D(new_n196_), .Y(new_n3470_));
  OR4X1    g03406(.A(new_n1223_), .B(new_n1135_), .C(new_n850_), .D(new_n227_), .Y(new_n3471_));
  OR2X1    g03407(.A(new_n3471_), .B(new_n3470_), .Y(new_n3472_));
  OR2X1    g03408(.A(new_n3472_), .B(new_n1761_), .Y(new_n3473_));
  OR4X1    g03409(.A(new_n3473_), .B(new_n3469_), .C(new_n3468_), .D(new_n3466_), .Y(new_n3474_));
  NOR3X1   g03410(.A(new_n3474_), .B(new_n3463_), .C(new_n1015_), .Y(new_n3475_));
  NOR2X1   g03411(.A(new_n3475_), .B(new_n3431_), .Y(new_n3476_));
  XOR2X1   g03412(.A(new_n1536_), .B(new_n1490_), .Y(new_n3477_));
  XOR2X1   g03413(.A(new_n3477_), .B(new_n1797_), .Y(new_n3478_));
  INVX1    g03414(.A(new_n3478_), .Y(new_n3479_));
  INVX1    g03415(.A(new_n1586_), .Y(new_n3480_));
  AOI22X1  g03416(.A0(new_n1890_), .A1(new_n3480_), .B0(new_n1889_), .B1(new_n1490_), .Y(new_n3481_));
  OAI21X1  g03417(.A0(new_n1885_), .A1(new_n1795_), .B0(new_n3481_), .Y(new_n3482_));
  AOI21X1  g03418(.A0(new_n3479_), .A1(new_n407_), .B0(new_n3482_), .Y(new_n3483_));
  NOR4X1   g03419(.A(new_n3474_), .B(new_n3463_), .C(new_n1015_), .D(\a[2] ), .Y(new_n3484_));
  NOR3X1   g03420(.A(new_n3484_), .B(new_n3483_), .C(new_n3476_), .Y(new_n3485_));
  NOR2X1   g03421(.A(new_n3485_), .B(new_n3476_), .Y(new_n3486_));
  INVX1    g03422(.A(new_n3486_), .Y(new_n3487_));
  AND2X1   g03423(.A(new_n3455_), .B(new_n3431_), .Y(new_n3488_));
  INVX1    g03424(.A(new_n3488_), .Y(new_n3489_));
  AOI21X1  g03425(.A0(new_n3489_), .A1(new_n3487_), .B0(new_n3456_), .Y(new_n3490_));
  INVX1    g03426(.A(new_n3490_), .Y(new_n3491_));
  XOR2X1   g03427(.A(new_n3442_), .B(new_n3431_), .Y(new_n3492_));
  AOI21X1  g03428(.A0(new_n3492_), .A1(new_n3491_), .B0(new_n3443_), .Y(new_n3493_));
  INVX1    g03429(.A(new_n3493_), .Y(new_n3494_));
  XOR2X1   g03430(.A(new_n3322_), .B(new_n3289_), .Y(new_n3495_));
  AND2X1   g03431(.A(new_n3495_), .B(new_n3494_), .Y(new_n3496_));
  XOR2X1   g03432(.A(new_n1806_), .B(new_n1805_), .Y(new_n3497_));
  INVX1    g03433(.A(new_n1889_), .Y(new_n3498_));
  AOI22X1  g03434(.A0(new_n1890_), .A1(new_n1800_), .B0(new_n1884_), .B1(new_n3327_), .Y(new_n3499_));
  OAI21X1  g03435(.A0(new_n3498_), .A1(new_n1389_), .B0(new_n3499_), .Y(new_n3500_));
  AOI21X1  g03436(.A0(new_n3497_), .A1(new_n407_), .B0(new_n3500_), .Y(new_n3501_));
  INVX1    g03437(.A(new_n3501_), .Y(new_n3502_));
  XOR2X1   g03438(.A(new_n3495_), .B(new_n3494_), .Y(new_n3503_));
  AOI21X1  g03439(.A0(new_n3503_), .A1(new_n3502_), .B0(new_n3496_), .Y(new_n3504_));
  NOR2X1   g03440(.A(new_n3504_), .B(new_n3430_), .Y(new_n3505_));
  INVX1    g03441(.A(new_n3430_), .Y(new_n3506_));
  XOR2X1   g03442(.A(new_n3504_), .B(new_n3506_), .Y(new_n3507_));
  OAI22X1  g03443(.A0(new_n2186_), .A1(new_n1339_), .B0(new_n2140_), .B1(new_n1236_), .Y(new_n3508_));
  AOI21X1  g03444(.A0(new_n2095_), .A1(new_n3342_), .B0(new_n3508_), .Y(new_n3509_));
  OAI21X1  g03445(.A0(new_n3053_), .A1(new_n2063_), .B0(new_n3509_), .Y(new_n3510_));
  XOR2X1   g03446(.A(new_n3510_), .B(new_n74_), .Y(new_n3511_));
  NOR2X1   g03447(.A(new_n3511_), .B(new_n3507_), .Y(new_n3512_));
  NOR2X1   g03448(.A(new_n3512_), .B(new_n3505_), .Y(new_n3513_));
  INVX1    g03449(.A(new_n3424_), .Y(new_n3514_));
  XOR2X1   g03450(.A(new_n3428_), .B(new_n3514_), .Y(new_n3515_));
  OR2X1    g03451(.A(new_n3515_), .B(new_n3513_), .Y(new_n3516_));
  AND2X1   g03452(.A(new_n3516_), .B(new_n3429_), .Y(new_n3517_));
  OAI21X1  g03453(.A0(new_n3517_), .A1(new_n3421_), .B0(new_n3419_), .Y(new_n3518_));
  XOR2X1   g03454(.A(new_n3356_), .B(new_n3351_), .Y(new_n3519_));
  AND2X1   g03455(.A(new_n3519_), .B(new_n3518_), .Y(new_n3520_));
  XOR2X1   g03456(.A(new_n3519_), .B(new_n3518_), .Y(new_n3521_));
  AOI22X1  g03457(.A0(new_n2424_), .A1(new_n2603_), .B0(new_n2423_), .B1(new_n2602_), .Y(new_n3522_));
  OAI21X1  g03458(.A0(new_n2419_), .A1(new_n957_), .B0(new_n3522_), .Y(new_n3523_));
  AOI21X1  g03459(.A0(new_n2601_), .A1(new_n2301_), .B0(new_n3523_), .Y(new_n3524_));
  XOR2X1   g03460(.A(new_n3524_), .B(new_n89_), .Y(new_n3525_));
  AOI21X1  g03461(.A0(new_n3525_), .A1(new_n3521_), .B0(new_n3520_), .Y(new_n3526_));
  NOR2X1   g03462(.A(new_n3526_), .B(new_n3412_), .Y(new_n3527_));
  XOR2X1   g03463(.A(new_n3526_), .B(new_n3412_), .Y(new_n3528_));
  AOI22X1  g03464(.A0(new_n2745_), .A1(new_n1886_), .B0(new_n2657_), .B1(new_n2036_), .Y(new_n3529_));
  OAI21X1  g03465(.A0(new_n2743_), .A1(new_n690_), .B0(new_n3529_), .Y(new_n3530_));
  AOI21X1  g03466(.A0(new_n2658_), .A1(new_n2035_), .B0(new_n3530_), .Y(new_n3531_));
  XOR2X1   g03467(.A(new_n3531_), .B(new_n70_), .Y(new_n3532_));
  AOI21X1  g03468(.A0(new_n3532_), .A1(new_n3528_), .B0(new_n3527_), .Y(new_n3533_));
  NOR2X1   g03469(.A(new_n3533_), .B(new_n3410_), .Y(new_n3534_));
  AOI21X1  g03470(.A0(new_n3409_), .A1(new_n3408_), .B0(new_n3534_), .Y(new_n3535_));
  NOR2X1   g03471(.A(new_n3535_), .B(new_n3403_), .Y(new_n3536_));
  XOR2X1   g03472(.A(new_n3535_), .B(new_n3403_), .Y(new_n3537_));
  AOI22X1  g03473(.A0(new_n3146_), .A1(new_n2252_), .B0(new_n2875_), .B1(new_n2246_), .Y(new_n3538_));
  OAI21X1  g03474(.A0(new_n3144_), .A1(new_n2092_), .B0(new_n3538_), .Y(new_n3539_));
  AOI21X1  g03475(.A0(new_n2876_), .A1(new_n2201_), .B0(new_n3539_), .Y(new_n3540_));
  XOR2X1   g03476(.A(new_n3540_), .B(new_n1920_), .Y(new_n3541_));
  AOI21X1  g03477(.A0(new_n3541_), .A1(new_n3537_), .B0(new_n3536_), .Y(new_n3542_));
  NOR2X1   g03478(.A(new_n3542_), .B(new_n3401_), .Y(new_n3543_));
  XOR2X1   g03479(.A(new_n3542_), .B(new_n3401_), .Y(new_n3544_));
  OR2X1    g03480(.A(new_n3230_), .B(new_n3227_), .Y(new_n3545_));
  INVX1    g03481(.A(new_n3545_), .Y(new_n3546_));
  AOI22X1  g03482(.A0(new_n3546_), .A1(new_n2421_), .B0(new_n3232_), .B1(new_n2420_), .Y(new_n3547_));
  OAI21X1  g03483(.A0(new_n3389_), .A1(new_n2379_), .B0(new_n3547_), .Y(new_n3548_));
  AOI21X1  g03484(.A0(new_n3234_), .A1(new_n2416_), .B0(new_n3548_), .Y(new_n3549_));
  XOR2X1   g03485(.A(new_n3549_), .B(new_n2445_), .Y(new_n3550_));
  AOI21X1  g03486(.A0(new_n3550_), .A1(new_n3544_), .B0(new_n3543_), .Y(new_n3551_));
  OAI22X1  g03487(.A0(new_n3545_), .A1(new_n2648_), .B0(new_n3389_), .B1(new_n2414_), .Y(new_n3552_));
  AOI21X1  g03488(.A0(new_n3232_), .A1(new_n2752_), .B0(new_n3552_), .Y(new_n3553_));
  OAI21X1  g03489(.A0(new_n3388_), .A1(new_n2757_), .B0(new_n3553_), .Y(new_n3554_));
  XOR2X1   g03490(.A(new_n3554_), .B(new_n2445_), .Y(new_n3555_));
  NOR2X1   g03491(.A(new_n3555_), .B(new_n3551_), .Y(new_n3556_));
  XOR2X1   g03492(.A(new_n3555_), .B(new_n3551_), .Y(new_n3557_));
  XOR2X1   g03493(.A(new_n3383_), .B(new_n3382_), .Y(new_n3558_));
  AOI21X1  g03494(.A0(new_n3558_), .A1(new_n3557_), .B0(new_n3556_), .Y(new_n3559_));
  NOR2X1   g03495(.A(new_n3559_), .B(new_n3400_), .Y(new_n3560_));
  XOR2X1   g03496(.A(new_n3559_), .B(new_n3400_), .Y(new_n3561_));
  XOR2X1   g03497(.A(new_n3541_), .B(new_n3537_), .Y(new_n3562_));
  INVX1    g03498(.A(new_n3410_), .Y(new_n3563_));
  XOR2X1   g03499(.A(new_n3533_), .B(new_n3563_), .Y(new_n3564_));
  AOI22X1  g03500(.A0(new_n3146_), .A1(new_n2093_), .B0(new_n2875_), .B1(new_n1887_), .Y(new_n3565_));
  OAI21X1  g03501(.A0(new_n3144_), .A1(new_n2183_), .B0(new_n3565_), .Y(new_n3566_));
  AOI21X1  g03502(.A0(new_n2876_), .A1(new_n2430_), .B0(new_n3566_), .Y(new_n3567_));
  XOR2X1   g03503(.A(new_n3567_), .B(\a[20] ), .Y(new_n3568_));
  NOR2X1   g03504(.A(new_n3568_), .B(new_n3564_), .Y(new_n3569_));
  XOR2X1   g03505(.A(new_n3532_), .B(new_n3528_), .Y(new_n3570_));
  INVX1    g03506(.A(new_n3570_), .Y(new_n3571_));
  XOR2X1   g03507(.A(new_n3524_), .B(\a[26] ), .Y(new_n3572_));
  XOR2X1   g03508(.A(new_n3572_), .B(new_n3521_), .Y(new_n3573_));
  XOR2X1   g03509(.A(new_n3517_), .B(new_n3420_), .Y(new_n3574_));
  OAI22X1  g03510(.A0(new_n2626_), .A1(new_n957_), .B0(new_n2419_), .B1(new_n985_), .Y(new_n3575_));
  AOI21X1  g03511(.A0(new_n2424_), .A1(new_n1822_), .B0(new_n3575_), .Y(new_n3576_));
  OAI21X1  g03512(.A0(new_n2833_), .A1(new_n2665_), .B0(new_n3576_), .Y(new_n3577_));
  XOR2X1   g03513(.A(new_n3577_), .B(new_n89_), .Y(new_n3578_));
  NOR2X1   g03514(.A(new_n3578_), .B(new_n3574_), .Y(new_n3579_));
  XOR2X1   g03515(.A(new_n3515_), .B(new_n3513_), .Y(new_n3580_));
  INVX1    g03516(.A(new_n3580_), .Y(new_n3581_));
  OAI22X1  g03517(.A0(new_n2140_), .A1(new_n1189_), .B0(new_n2431_), .B1(new_n1236_), .Y(new_n3582_));
  AOI21X1  g03518(.A0(new_n2185_), .A1(new_n3342_), .B0(new_n3582_), .Y(new_n3583_));
  OAI21X1  g03519(.A0(new_n3180_), .A1(new_n2063_), .B0(new_n3583_), .Y(new_n3584_));
  XOR2X1   g03520(.A(new_n3584_), .B(new_n74_), .Y(new_n3585_));
  OR2X1    g03521(.A(new_n3585_), .B(new_n3581_), .Y(new_n3586_));
  AND2X1   g03522(.A(new_n3585_), .B(new_n3581_), .Y(new_n3587_));
  AOI22X1  g03523(.A0(new_n2424_), .A1(new_n1126_), .B0(new_n2423_), .B1(new_n2603_), .Y(new_n3588_));
  OAI21X1  g03524(.A0(new_n2419_), .A1(new_n1065_), .B0(new_n3588_), .Y(new_n3589_));
  AOI21X1  g03525(.A0(new_n2824_), .A1(new_n2301_), .B0(new_n3589_), .Y(new_n3590_));
  XOR2X1   g03526(.A(new_n3590_), .B(\a[26] ), .Y(new_n3591_));
  OAI21X1  g03527(.A0(new_n3591_), .A1(new_n3587_), .B0(new_n3586_), .Y(new_n3592_));
  XOR2X1   g03528(.A(new_n3578_), .B(new_n3574_), .Y(new_n3593_));
  AOI21X1  g03529(.A0(new_n3593_), .A1(new_n3592_), .B0(new_n3579_), .Y(new_n3594_));
  NOR2X1   g03530(.A(new_n3594_), .B(new_n3573_), .Y(new_n3595_));
  XOR2X1   g03531(.A(new_n3594_), .B(new_n3573_), .Y(new_n3596_));
  AOI22X1  g03532(.A0(new_n2745_), .A1(new_n2049_), .B0(new_n2657_), .B1(new_n2481_), .Y(new_n3597_));
  OAI21X1  g03533(.A0(new_n2743_), .A1(new_n783_), .B0(new_n3597_), .Y(new_n3598_));
  AOI21X1  g03534(.A0(new_n2658_), .A1(new_n2480_), .B0(new_n3598_), .Y(new_n3599_));
  XOR2X1   g03535(.A(new_n3599_), .B(new_n70_), .Y(new_n3600_));
  AOI21X1  g03536(.A0(new_n3600_), .A1(new_n3596_), .B0(new_n3595_), .Y(new_n3601_));
  OR2X1    g03537(.A(new_n3601_), .B(new_n3571_), .Y(new_n3602_));
  XOR2X1   g03538(.A(new_n3601_), .B(new_n3571_), .Y(new_n3603_));
  INVX1    g03539(.A(new_n3603_), .Y(new_n3604_));
  AOI22X1  g03540(.A0(new_n3146_), .A1(new_n2246_), .B0(new_n2875_), .B1(new_n2048_), .Y(new_n3605_));
  OAI21X1  g03541(.A0(new_n3144_), .A1(new_n1879_), .B0(new_n3605_), .Y(new_n3606_));
  AOI21X1  g03542(.A0(new_n2876_), .A1(new_n2244_), .B0(new_n3606_), .Y(new_n3607_));
  XOR2X1   g03543(.A(new_n3607_), .B(\a[20] ), .Y(new_n3608_));
  OAI21X1  g03544(.A0(new_n3608_), .A1(new_n3604_), .B0(new_n3602_), .Y(new_n3609_));
  XOR2X1   g03545(.A(new_n3568_), .B(new_n3564_), .Y(new_n3610_));
  AND2X1   g03546(.A(new_n3610_), .B(new_n3609_), .Y(new_n3611_));
  OAI21X1  g03547(.A0(new_n3611_), .A1(new_n3569_), .B0(new_n3562_), .Y(new_n3612_));
  AOI21X1  g03548(.A0(new_n3610_), .A1(new_n3609_), .B0(new_n3569_), .Y(new_n3613_));
  XOR2X1   g03549(.A(new_n3613_), .B(new_n3562_), .Y(new_n3614_));
  AOI22X1  g03550(.A0(new_n3390_), .A1(new_n2420_), .B0(new_n3232_), .B1(new_n2627_), .Y(new_n3615_));
  OAI21X1  g03551(.A0(new_n3545_), .A1(new_n2379_), .B0(new_n3615_), .Y(new_n3616_));
  AOI21X1  g03552(.A0(new_n3234_), .A1(new_n2625_), .B0(new_n3616_), .Y(new_n3617_));
  XOR2X1   g03553(.A(new_n3617_), .B(\a[17] ), .Y(new_n3618_));
  OR2X1    g03554(.A(new_n3618_), .B(new_n3614_), .Y(new_n3619_));
  AND2X1   g03555(.A(new_n3619_), .B(new_n3612_), .Y(new_n3620_));
  XOR2X1   g03556(.A(\a[12] ), .B(new_n2911_), .Y(new_n3621_));
  XOR2X1   g03557(.A(\a[14] ), .B(\a[13] ), .Y(new_n3622_));
  INVX1    g03558(.A(new_n3622_), .Y(new_n3623_));
  NOR2X1   g03559(.A(new_n3623_), .B(new_n3621_), .Y(new_n3624_));
  XOR2X1   g03560(.A(\a[13] ), .B(\a[12] ), .Y(new_n3625_));
  INVX1    g03561(.A(new_n3625_), .Y(new_n3626_));
  NAND3X1  g03562(.A(new_n3626_), .B(new_n3622_), .C(new_n3621_), .Y(new_n3627_));
  INVX1    g03563(.A(new_n3627_), .Y(new_n3628_));
  AOI22X1  g03564(.A0(new_n3628_), .A1(new_n2649_), .B0(new_n3624_), .B1(new_n2652_), .Y(new_n3629_));
  XOR2X1   g03565(.A(new_n3629_), .B(\a[14] ), .Y(new_n3630_));
  NOR2X1   g03566(.A(new_n3630_), .B(new_n3620_), .Y(new_n3631_));
  XOR2X1   g03567(.A(new_n3550_), .B(new_n3544_), .Y(new_n3632_));
  XOR2X1   g03568(.A(new_n3630_), .B(new_n3620_), .Y(new_n3633_));
  AOI21X1  g03569(.A0(new_n3633_), .A1(new_n3632_), .B0(new_n3631_), .Y(new_n3634_));
  INVX1    g03570(.A(new_n3634_), .Y(new_n3635_));
  XOR2X1   g03571(.A(new_n3558_), .B(new_n3557_), .Y(new_n3636_));
  AND2X1   g03572(.A(new_n3636_), .B(new_n3635_), .Y(new_n3637_));
  INVX1    g03573(.A(new_n3637_), .Y(new_n3638_));
  XOR2X1   g03574(.A(new_n3636_), .B(new_n3635_), .Y(new_n3639_));
  INVX1    g03575(.A(new_n3639_), .Y(new_n3640_));
  XOR2X1   g03576(.A(new_n3633_), .B(new_n3632_), .Y(new_n3641_));
  INVX1    g03577(.A(new_n3641_), .Y(new_n3642_));
  AOI22X1  g03578(.A0(new_n3546_), .A1(new_n2420_), .B0(new_n3232_), .B1(new_n2252_), .Y(new_n3643_));
  OAI21X1  g03579(.A0(new_n3389_), .A1(new_n2287_), .B0(new_n3643_), .Y(new_n3644_));
  AOI21X1  g03580(.A0(new_n3234_), .A1(new_n2669_), .B0(new_n3644_), .Y(new_n3645_));
  XOR2X1   g03581(.A(new_n3645_), .B(\a[17] ), .Y(new_n3646_));
  INVX1    g03582(.A(new_n3646_), .Y(new_n3647_));
  XOR2X1   g03583(.A(new_n3610_), .B(new_n3609_), .Y(new_n3648_));
  XOR2X1   g03584(.A(new_n3648_), .B(new_n3646_), .Y(new_n3649_));
  XOR2X1   g03585(.A(new_n3608_), .B(new_n3603_), .Y(new_n3650_));
  XOR2X1   g03586(.A(new_n3600_), .B(new_n3596_), .Y(new_n3651_));
  INVX1    g03587(.A(new_n3651_), .Y(new_n3652_));
  AOI22X1  g03588(.A0(new_n2745_), .A1(new_n2036_), .B0(new_n2657_), .B1(new_n2602_), .Y(new_n3653_));
  OAI21X1  g03589(.A0(new_n2743_), .A1(new_n847_), .B0(new_n3653_), .Y(new_n3654_));
  AOI21X1  g03590(.A0(new_n2658_), .A1(new_n2494_), .B0(new_n3654_), .Y(new_n3655_));
  XOR2X1   g03591(.A(new_n3655_), .B(\a[23] ), .Y(new_n3656_));
  INVX1    g03592(.A(new_n3656_), .Y(new_n3657_));
  XOR2X1   g03593(.A(new_n3593_), .B(new_n3592_), .Y(new_n3658_));
  XOR2X1   g03594(.A(new_n3658_), .B(new_n3656_), .Y(new_n3659_));
  XOR2X1   g03595(.A(new_n3585_), .B(new_n3581_), .Y(new_n3660_));
  XOR2X1   g03596(.A(new_n3591_), .B(new_n3660_), .Y(new_n3661_));
  XOR2X1   g03597(.A(new_n3503_), .B(new_n3501_), .Y(new_n3662_));
  INVX1    g03598(.A(new_n3662_), .Y(new_n3663_));
  AND2X1   g03599(.A(new_n3442_), .B(new_n3431_), .Y(new_n3664_));
  OAI22X1  g03600(.A0(new_n3494_), .A1(new_n3664_), .B0(new_n3492_), .B1(new_n3490_), .Y(new_n3665_));
  AOI21X1  g03601(.A0(new_n1801_), .A1(new_n1799_), .B0(new_n1489_), .Y(new_n3666_));
  XOR2X1   g03602(.A(new_n1803_), .B(new_n3666_), .Y(new_n3667_));
  NOR2X1   g03603(.A(new_n3667_), .B(new_n3178_), .Y(new_n3668_));
  INVX1    g03604(.A(new_n1490_), .Y(new_n3669_));
  AOI22X1  g03605(.A0(new_n1889_), .A1(new_n3327_), .B0(new_n1884_), .B1(new_n1800_), .Y(new_n3670_));
  OAI21X1  g03606(.A0(new_n2245_), .A1(new_n3669_), .B0(new_n3670_), .Y(new_n3671_));
  OAI21X1  g03607(.A0(new_n3671_), .A1(new_n3668_), .B0(new_n3665_), .Y(new_n3672_));
  OAI22X1  g03608(.A0(new_n3488_), .A1(new_n3456_), .B0(new_n3485_), .B1(new_n3476_), .Y(new_n3673_));
  OAI21X1  g03609(.A0(new_n3491_), .A1(new_n3488_), .B0(new_n3673_), .Y(new_n3674_));
  INVX1    g03610(.A(new_n1801_), .Y(new_n3675_));
  XOR2X1   g03611(.A(new_n3675_), .B(new_n1799_), .Y(new_n3676_));
  NOR2X1   g03612(.A(new_n3676_), .B(new_n3178_), .Y(new_n3677_));
  AOI22X1  g03613(.A0(new_n1889_), .A1(new_n1800_), .B0(new_n1884_), .B1(new_n1490_), .Y(new_n3678_));
  OAI21X1  g03614(.A0(new_n2245_), .A1(new_n1795_), .B0(new_n3678_), .Y(new_n3679_));
  OAI21X1  g03615(.A0(new_n3679_), .A1(new_n3677_), .B0(new_n3674_), .Y(new_n3680_));
  OAI22X1  g03616(.A0(new_n3487_), .A1(new_n3484_), .B0(new_n3485_), .B1(new_n3483_), .Y(new_n3681_));
  INVX1    g03617(.A(new_n3681_), .Y(new_n3682_));
  INVX1    g03618(.A(new_n2566_), .Y(new_n3683_));
  NAND3X1  g03619(.A(new_n3293_), .B(new_n1164_), .C(new_n179_), .Y(new_n3684_));
  OR4X1    g03620(.A(new_n2999_), .B(new_n1261_), .C(new_n393_), .D(new_n390_), .Y(new_n3685_));
  OR4X1    g03621(.A(new_n2178_), .B(new_n1259_), .C(new_n716_), .D(new_n668_), .Y(new_n3686_));
  OR4X1    g03622(.A(new_n365_), .B(new_n565_), .C(new_n233_), .D(new_n191_), .Y(new_n3687_));
  OR4X1    g03623(.A(new_n3687_), .B(new_n1044_), .C(new_n506_), .D(new_n273_), .Y(new_n3688_));
  OR4X1    g03624(.A(new_n3688_), .B(new_n3686_), .C(new_n3685_), .D(new_n3684_), .Y(new_n3689_));
  OR4X1    g03625(.A(new_n1061_), .B(new_n945_), .C(new_n831_), .D(new_n465_), .Y(new_n3690_));
  NOR3X1   g03626(.A(new_n219_), .B(new_n187_), .C(new_n153_), .Y(new_n3691_));
  NAND4X1  g03627(.A(new_n3691_), .B(new_n469_), .C(new_n324_), .D(new_n281_), .Y(new_n3692_));
  OR4X1    g03628(.A(new_n2795_), .B(new_n2580_), .C(new_n412_), .D(new_n100_), .Y(new_n3693_));
  OR4X1    g03629(.A(new_n3693_), .B(new_n3692_), .C(new_n3690_), .D(new_n2534_), .Y(new_n3694_));
  OR2X1    g03630(.A(new_n3694_), .B(new_n1325_), .Y(new_n3695_));
  NOR4X1   g03631(.A(new_n3695_), .B(new_n3689_), .C(new_n2579_), .D(new_n3683_), .Y(new_n3696_));
  XOR2X1   g03632(.A(new_n1796_), .B(new_n1794_), .Y(new_n3697_));
  AOI22X1  g03633(.A0(new_n1889_), .A1(new_n1536_), .B0(new_n1884_), .B1(new_n3480_), .Y(new_n3698_));
  OAI21X1  g03634(.A0(new_n2245_), .A1(new_n1621_), .B0(new_n3698_), .Y(new_n3699_));
  AOI21X1  g03635(.A0(new_n3697_), .A1(new_n407_), .B0(new_n3699_), .Y(new_n3700_));
  NOR2X1   g03636(.A(new_n3700_), .B(new_n3696_), .Y(new_n3701_));
  OAI22X1  g03637(.A0(new_n182_), .A1(new_n102_), .B0(new_n125_), .B1(new_n96_), .Y(new_n3702_));
  OR4X1    g03638(.A(new_n3702_), .B(new_n938_), .C(new_n561_), .D(new_n806_), .Y(new_n3703_));
  OR2X1    g03639(.A(new_n1493_), .B(new_n1608_), .Y(new_n3704_));
  OR4X1    g03640(.A(new_n1277_), .B(new_n1259_), .C(new_n1255_), .D(new_n827_), .Y(new_n3705_));
  OR4X1    g03641(.A(new_n3705_), .B(new_n3704_), .C(new_n3703_), .D(new_n2561_), .Y(new_n3706_));
  OR4X1    g03642(.A(new_n1082_), .B(new_n429_), .C(new_n968_), .D(new_n420_), .Y(new_n3707_));
  OR4X1    g03643(.A(new_n3707_), .B(new_n552_), .C(new_n504_), .D(new_n356_), .Y(new_n3708_));
  OR4X1    g03644(.A(new_n1398_), .B(new_n243_), .C(new_n539_), .D(new_n133_), .Y(new_n3709_));
  OR4X1    g03645(.A(new_n3709_), .B(new_n3708_), .C(new_n2939_), .D(new_n2105_), .Y(new_n3710_));
  OR4X1    g03646(.A(new_n229_), .B(new_n426_), .C(new_n651_), .D(new_n1046_), .Y(new_n3711_));
  OR4X1    g03647(.A(new_n3711_), .B(new_n679_), .C(new_n840_), .D(new_n263_), .Y(new_n3712_));
  OAI22X1  g03648(.A0(new_n152_), .A1(new_n94_), .B0(new_n96_), .B1(new_n92_), .Y(new_n3713_));
  OR2X1    g03649(.A(new_n3713_), .B(new_n497_), .Y(new_n3714_));
  OR4X1    g03650(.A(new_n3714_), .B(new_n632_), .C(new_n408_), .D(new_n199_), .Y(new_n3715_));
  OR4X1    g03651(.A(new_n1319_), .B(new_n1211_), .C(new_n463_), .D(new_n164_), .Y(new_n3716_));
  OR4X1    g03652(.A(new_n3716_), .B(new_n3715_), .C(new_n3712_), .D(new_n2464_), .Y(new_n3717_));
  NOR4X1   g03653(.A(new_n3717_), .B(new_n3710_), .C(new_n3706_), .D(new_n492_), .Y(new_n3718_));
  XOR2X1   g03654(.A(new_n1792_), .B(new_n1791_), .Y(new_n3719_));
  INVX1    g03655(.A(new_n3719_), .Y(new_n3720_));
  INVX1    g03656(.A(new_n1655_), .Y(new_n3721_));
  AOI22X1  g03657(.A0(new_n1890_), .A1(new_n3721_), .B0(new_n1889_), .B1(new_n3480_), .Y(new_n3722_));
  OAI21X1  g03658(.A0(new_n1885_), .A1(new_n1621_), .B0(new_n3722_), .Y(new_n3723_));
  AOI21X1  g03659(.A0(new_n3720_), .A1(new_n407_), .B0(new_n3723_), .Y(new_n3724_));
  OR2X1    g03660(.A(new_n3724_), .B(new_n3718_), .Y(new_n3725_));
  NOR3X1   g03661(.A(new_n402_), .B(new_n389_), .C(new_n378_), .Y(new_n3726_));
  OR4X1    g03662(.A(new_n1485_), .B(new_n596_), .C(new_n457_), .D(new_n181_), .Y(new_n3727_));
  OR4X1    g03663(.A(new_n1044_), .B(new_n603_), .C(new_n282_), .D(new_n439_), .Y(new_n3728_));
  OR4X1    g03664(.A(new_n408_), .B(new_n260_), .C(new_n199_), .D(new_n114_), .Y(new_n3729_));
  OR4X1    g03665(.A(new_n3729_), .B(new_n3728_), .C(new_n3727_), .D(new_n1159_), .Y(new_n3730_));
  OAI22X1  g03666(.A0(new_n125_), .A1(new_n69_), .B0(new_n105_), .B1(new_n96_), .Y(new_n3731_));
  OR4X1    g03667(.A(new_n747_), .B(new_n301_), .C(new_n206_), .D(new_n80_), .Y(new_n3732_));
  OR4X1    g03668(.A(new_n1451_), .B(new_n741_), .C(new_n642_), .D(new_n547_), .Y(new_n3733_));
  OR4X1    g03669(.A(new_n3733_), .B(new_n3732_), .C(new_n1515_), .D(new_n3731_), .Y(new_n3734_));
  NOR4X1   g03670(.A(new_n3734_), .B(new_n3730_), .C(new_n2268_), .D(new_n1549_), .Y(new_n3735_));
  OR4X1    g03671(.A(new_n422_), .B(new_n840_), .C(new_n757_), .D(new_n928_), .Y(new_n3736_));
  OR4X1    g03672(.A(new_n3736_), .B(new_n1216_), .C(new_n1197_), .D(new_n848_), .Y(new_n3737_));
  OR4X1    g03673(.A(new_n814_), .B(new_n493_), .C(new_n792_), .D(new_n162_), .Y(new_n3738_));
  OR4X1    g03674(.A(new_n3738_), .B(new_n2989_), .C(new_n1067_), .D(new_n714_), .Y(new_n3739_));
  OR4X1    g03675(.A(new_n1316_), .B(new_n460_), .C(new_n234_), .D(new_n535_), .Y(new_n3740_));
  OR4X1    g03676(.A(new_n1306_), .B(new_n720_), .C(new_n321_), .D(new_n286_), .Y(new_n3741_));
  NOR4X1   g03677(.A(new_n3741_), .B(new_n3740_), .C(new_n3739_), .D(new_n3737_), .Y(new_n3742_));
  NAND3X1  g03678(.A(new_n3742_), .B(new_n3735_), .C(new_n3726_), .Y(new_n3743_));
  INVX1    g03679(.A(new_n3743_), .Y(new_n3744_));
  XOR2X1   g03680(.A(new_n1790_), .B(new_n1789_), .Y(new_n3745_));
  AOI22X1  g03681(.A0(new_n1890_), .A1(new_n1676_), .B0(new_n1884_), .B1(new_n3721_), .Y(new_n3746_));
  OAI21X1  g03682(.A0(new_n3498_), .A1(new_n1621_), .B0(new_n3746_), .Y(new_n3747_));
  AOI21X1  g03683(.A0(new_n3745_), .A1(new_n407_), .B0(new_n3747_), .Y(new_n3748_));
  NOR2X1   g03684(.A(new_n3748_), .B(new_n3744_), .Y(new_n3749_));
  INVX1    g03685(.A(new_n3749_), .Y(new_n3750_));
  INVX1    g03686(.A(new_n1507_), .Y(new_n3751_));
  INVX1    g03687(.A(new_n2027_), .Y(new_n3752_));
  OR4X1    g03688(.A(new_n2101_), .B(new_n2088_), .C(new_n1134_), .D(new_n313_), .Y(new_n3753_));
  OAI22X1  g03689(.A0(new_n148_), .A1(new_n92_), .B0(new_n119_), .B1(new_n99_), .Y(new_n3754_));
  OR2X1    g03690(.A(new_n3754_), .B(new_n631_), .Y(new_n3755_));
  OR4X1    g03691(.A(new_n319_), .B(new_n246_), .C(new_n177_), .D(new_n134_), .Y(new_n3756_));
  NOR4X1   g03692(.A(new_n3756_), .B(new_n3755_), .C(new_n3753_), .D(new_n3752_), .Y(new_n3757_));
  INVX1    g03693(.A(new_n3757_), .Y(new_n3758_));
  OR4X1    g03694(.A(new_n612_), .B(new_n372_), .C(new_n294_), .D(new_n439_), .Y(new_n3759_));
  OR4X1    g03695(.A(new_n586_), .B(new_n478_), .C(new_n328_), .D(new_n410_), .Y(new_n3760_));
  NOR3X1   g03696(.A(new_n676_), .B(new_n740_), .C(new_n348_), .Y(new_n3761_));
  INVX1    g03697(.A(new_n3761_), .Y(new_n3762_));
  OR4X1    g03698(.A(new_n3762_), .B(new_n3760_), .C(new_n3759_), .D(new_n1207_), .Y(new_n3763_));
  OAI22X1  g03699(.A0(new_n182_), .A1(new_n91_), .B0(new_n108_), .B1(new_n79_), .Y(new_n3764_));
  OAI22X1  g03700(.A0(new_n108_), .A1(new_n88_), .B0(new_n92_), .B1(new_n79_), .Y(new_n3765_));
  OR4X1    g03701(.A(new_n3765_), .B(new_n3764_), .C(new_n743_), .D(new_n178_), .Y(new_n3766_));
  OR4X1    g03702(.A(new_n2536_), .B(new_n1703_), .C(new_n1142_), .D(new_n947_), .Y(new_n3767_));
  OR4X1    g03703(.A(new_n603_), .B(new_n648_), .C(new_n535_), .D(new_n124_), .Y(new_n3768_));
  OR2X1    g03704(.A(new_n873_), .B(new_n751_), .Y(new_n3769_));
  OR4X1    g03705(.A(new_n3769_), .B(new_n3768_), .C(new_n3767_), .D(new_n3766_), .Y(new_n3770_));
  NOR4X1   g03706(.A(new_n3770_), .B(new_n3763_), .C(new_n3758_), .D(new_n3751_), .Y(new_n3771_));
  XOR2X1   g03707(.A(new_n1674_), .B(new_n1655_), .Y(new_n3772_));
  XOR2X1   g03708(.A(new_n3772_), .B(new_n1787_), .Y(new_n3773_));
  INVX1    g03709(.A(new_n3773_), .Y(new_n3774_));
  AOI22X1  g03710(.A0(new_n1889_), .A1(new_n3721_), .B0(new_n1884_), .B1(new_n1676_), .Y(new_n3775_));
  OAI21X1  g03711(.A0(new_n2245_), .A1(new_n1708_), .B0(new_n3775_), .Y(new_n3776_));
  AOI21X1  g03712(.A0(new_n3774_), .A1(new_n407_), .B0(new_n3776_), .Y(new_n3777_));
  NOR2X1   g03713(.A(new_n3777_), .B(new_n3771_), .Y(new_n3778_));
  OR4X1    g03714(.A(new_n510_), .B(new_n370_), .C(new_n172_), .D(new_n85_), .Y(new_n3779_));
  AOI21X1  g03715(.A0(new_n143_), .A1(new_n94_), .B0(new_n84_), .Y(new_n3780_));
  NOR2X1   g03716(.A(new_n3780_), .B(new_n103_), .Y(new_n3781_));
  INVX1    g03717(.A(new_n3781_), .Y(new_n3782_));
  OR4X1    g03718(.A(new_n612_), .B(new_n565_), .C(new_n825_), .D(new_n1087_), .Y(new_n3783_));
  OR4X1    g03719(.A(new_n3783_), .B(new_n418_), .C(new_n387_), .D(new_n998_), .Y(new_n3784_));
  OR4X1    g03720(.A(new_n393_), .B(new_n627_), .C(new_n455_), .D(new_n207_), .Y(new_n3785_));
  OR4X1    g03721(.A(new_n382_), .B(new_n321_), .C(new_n493_), .D(new_n245_), .Y(new_n3786_));
  OR4X1    g03722(.A(new_n3786_), .B(new_n3785_), .C(new_n3784_), .D(new_n1201_), .Y(new_n3787_));
  OR4X1    g03723(.A(new_n3787_), .B(new_n3782_), .C(new_n3779_), .D(new_n973_), .Y(new_n3788_));
  NOR3X1   g03724(.A(new_n2302_), .B(new_n2097_), .C(new_n312_), .Y(new_n3789_));
  NOR4X1   g03725(.A(new_n723_), .B(new_n400_), .C(new_n814_), .D(new_n223_), .Y(new_n3790_));
  NAND3X1  g03726(.A(new_n3790_), .B(new_n3789_), .C(new_n1196_), .Y(new_n3791_));
  OR4X1    g03727(.A(new_n480_), .B(new_n226_), .C(new_n114_), .D(new_n585_), .Y(new_n3792_));
  OR2X1    g03728(.A(new_n744_), .B(new_n641_), .Y(new_n3793_));
  OR4X1    g03729(.A(new_n523_), .B(new_n261_), .C(new_n256_), .D(new_n231_), .Y(new_n3794_));
  OR4X1    g03730(.A(new_n848_), .B(new_n355_), .C(new_n296_), .D(new_n178_), .Y(new_n3795_));
  OR4X1    g03731(.A(new_n3795_), .B(new_n3794_), .C(new_n3793_), .D(new_n3792_), .Y(new_n3796_));
  OR4X1    g03732(.A(new_n361_), .B(new_n536_), .C(new_n522_), .D(new_n149_), .Y(new_n3797_));
  OR4X1    g03733(.A(new_n1599_), .B(new_n1171_), .C(new_n1142_), .D(new_n787_), .Y(new_n3798_));
  OR4X1    g03734(.A(new_n3798_), .B(new_n3797_), .C(new_n3796_), .D(new_n3791_), .Y(new_n3799_));
  OR4X1    g03735(.A(new_n3799_), .B(new_n3788_), .C(new_n1690_), .D(new_n1085_), .Y(new_n3800_));
  OR4X1    g03736(.A(new_n1028_), .B(new_n594_), .C(new_n455_), .D(new_n292_), .Y(new_n3801_));
  OR4X1    g03737(.A(new_n1724_), .B(new_n511_), .C(new_n974_), .D(new_n184_), .Y(new_n3802_));
  OR2X1    g03738(.A(new_n3802_), .B(new_n3801_), .Y(new_n3803_));
  NOR4X1   g03739(.A(new_n728_), .B(new_n701_), .C(new_n571_), .D(new_n514_), .Y(new_n3804_));
  NOR4X1   g03740(.A(new_n547_), .B(new_n418_), .C(new_n282_), .D(new_n274_), .Y(new_n3805_));
  NOR4X1   g03741(.A(new_n840_), .B(new_n301_), .C(new_n398_), .D(new_n219_), .Y(new_n3806_));
  NAND3X1  g03742(.A(new_n3806_), .B(new_n3805_), .C(new_n3804_), .Y(new_n3807_));
  OR4X1    g03743(.A(new_n1142_), .B(new_n814_), .C(new_n137_), .D(new_n133_), .Y(new_n3808_));
  OR4X1    g03744(.A(new_n1647_), .B(new_n1238_), .C(new_n1211_), .D(new_n830_), .Y(new_n3809_));
  OR4X1    g03745(.A(new_n3809_), .B(new_n3808_), .C(new_n3807_), .D(new_n3803_), .Y(new_n3810_));
  NAND4X1  g03746(.A(new_n392_), .B(new_n1564_), .C(new_n322_), .D(new_n1033_), .Y(new_n3811_));
  OR4X1    g03747(.A(new_n1473_), .B(new_n1306_), .C(new_n399_), .D(new_n1008_), .Y(new_n3812_));
  OR4X1    g03748(.A(new_n243_), .B(new_n232_), .C(new_n86_), .D(new_n85_), .Y(new_n3813_));
  OR2X1    g03749(.A(new_n768_), .B(new_n553_), .Y(new_n3814_));
  OR4X1    g03750(.A(new_n3814_), .B(new_n3813_), .C(new_n3812_), .D(new_n1403_), .Y(new_n3815_));
  NOR4X1   g03751(.A(new_n3815_), .B(new_n3811_), .C(new_n3760_), .D(new_n3300_), .Y(new_n3816_));
  INVX1    g03752(.A(new_n3816_), .Y(new_n3817_));
  NOR4X1   g03753(.A(new_n3817_), .B(new_n3810_), .C(new_n2466_), .D(new_n1431_), .Y(new_n3818_));
  OR4X1    g03754(.A(new_n1734_), .B(new_n1723_), .C(new_n1716_), .D(new_n1686_), .Y(new_n3819_));
  AOI21X1  g03755(.A0(new_n1784_), .A1(new_n3819_), .B0(new_n1706_), .Y(new_n3820_));
  OR4X1    g03756(.A(new_n1783_), .B(new_n1772_), .C(new_n1767_), .D(new_n1748_), .Y(new_n3821_));
  NOR3X1   g03757(.A(new_n3821_), .B(new_n1735_), .C(new_n1708_), .Y(new_n3822_));
  NOR3X1   g03758(.A(new_n3822_), .B(new_n3820_), .C(new_n3178_), .Y(new_n3823_));
  AOI22X1  g03759(.A0(new_n1890_), .A1(new_n3821_), .B0(new_n1884_), .B1(new_n3819_), .Y(new_n3824_));
  OAI21X1  g03760(.A0(new_n3498_), .A1(new_n1708_), .B0(new_n3824_), .Y(new_n3825_));
  NOR2X1   g03761(.A(new_n3825_), .B(new_n3823_), .Y(new_n3826_));
  NOR2X1   g03762(.A(new_n3826_), .B(new_n3818_), .Y(new_n3827_));
  AND2X1   g03763(.A(new_n3827_), .B(new_n3800_), .Y(new_n3828_));
  XOR2X1   g03764(.A(new_n1786_), .B(new_n1785_), .Y(new_n3829_));
  AOI22X1  g03765(.A0(new_n1890_), .A1(new_n3819_), .B0(new_n1889_), .B1(new_n1676_), .Y(new_n3830_));
  OAI21X1  g03766(.A0(new_n1885_), .A1(new_n1708_), .B0(new_n3830_), .Y(new_n3831_));
  AOI21X1  g03767(.A0(new_n3829_), .A1(new_n407_), .B0(new_n3831_), .Y(new_n3832_));
  INVX1    g03768(.A(new_n3832_), .Y(new_n3833_));
  XOR2X1   g03769(.A(new_n3827_), .B(new_n3800_), .Y(new_n3834_));
  AOI21X1  g03770(.A0(new_n3834_), .A1(new_n3833_), .B0(new_n3828_), .Y(new_n3835_));
  INVX1    g03771(.A(new_n3835_), .Y(new_n3836_));
  XOR2X1   g03772(.A(new_n3777_), .B(new_n3771_), .Y(new_n3837_));
  AOI21X1  g03773(.A0(new_n3837_), .A1(new_n3836_), .B0(new_n3778_), .Y(new_n3838_));
  XOR2X1   g03774(.A(new_n3748_), .B(new_n3743_), .Y(new_n3839_));
  OAI21X1  g03775(.A0(new_n3839_), .A1(new_n3838_), .B0(new_n3750_), .Y(new_n3840_));
  INVX1    g03776(.A(new_n3840_), .Y(new_n3841_));
  INVX1    g03777(.A(new_n3718_), .Y(new_n3842_));
  XOR2X1   g03778(.A(new_n3724_), .B(new_n3842_), .Y(new_n3843_));
  OAI21X1  g03779(.A0(new_n3843_), .A1(new_n3841_), .B0(new_n3725_), .Y(new_n3844_));
  XOR2X1   g03780(.A(new_n3700_), .B(new_n3696_), .Y(new_n3845_));
  AOI21X1  g03781(.A0(new_n3845_), .A1(new_n3844_), .B0(new_n3701_), .Y(new_n3846_));
  NOR2X1   g03782(.A(new_n3846_), .B(new_n3682_), .Y(new_n3847_));
  XOR2X1   g03783(.A(new_n3846_), .B(new_n3681_), .Y(new_n3848_));
  INVX1    g03784(.A(new_n3497_), .Y(new_n3849_));
  INVX1    g03785(.A(new_n1389_), .Y(new_n3850_));
  OAI22X1  g03786(.A0(new_n2186_), .A1(new_n1465_), .B0(new_n2431_), .B1(new_n1423_), .Y(new_n3851_));
  AOI21X1  g03787(.A0(new_n2139_), .A1(new_n3850_), .B0(new_n3851_), .Y(new_n3852_));
  OAI21X1  g03788(.A0(new_n3849_), .A1(new_n2063_), .B0(new_n3852_), .Y(new_n3853_));
  XOR2X1   g03789(.A(new_n3853_), .B(new_n74_), .Y(new_n3854_));
  NOR2X1   g03790(.A(new_n3854_), .B(new_n3848_), .Y(new_n3855_));
  NOR2X1   g03791(.A(new_n3855_), .B(new_n3847_), .Y(new_n3856_));
  NOR2X1   g03792(.A(new_n3679_), .B(new_n3677_), .Y(new_n3857_));
  XOR2X1   g03793(.A(new_n3857_), .B(new_n3674_), .Y(new_n3858_));
  OAI21X1  g03794(.A0(new_n3858_), .A1(new_n3856_), .B0(new_n3680_), .Y(new_n3859_));
  INVX1    g03795(.A(new_n3859_), .Y(new_n3860_));
  NOR2X1   g03796(.A(new_n3671_), .B(new_n3668_), .Y(new_n3861_));
  XOR2X1   g03797(.A(new_n3861_), .B(new_n3665_), .Y(new_n3862_));
  OAI21X1  g03798(.A0(new_n3862_), .A1(new_n3860_), .B0(new_n3672_), .Y(new_n3863_));
  AND2X1   g03799(.A(new_n3863_), .B(new_n3663_), .Y(new_n3864_));
  INVX1    g03800(.A(new_n3864_), .Y(new_n3865_));
  XOR2X1   g03801(.A(new_n3863_), .B(new_n3663_), .Y(new_n3866_));
  INVX1    g03802(.A(new_n3866_), .Y(new_n3867_));
  AOI22X1  g03803(.A0(new_n2185_), .A1(new_n1357_), .B0(new_n2139_), .B1(new_n3342_), .Y(new_n3868_));
  OAI21X1  g03804(.A0(new_n2431_), .A1(new_n1339_), .B0(new_n3868_), .Y(new_n3869_));
  AOI21X1  g03805(.A0(new_n3341_), .A1(new_n2062_), .B0(new_n3869_), .Y(new_n3870_));
  XOR2X1   g03806(.A(new_n3870_), .B(\a[29] ), .Y(new_n3871_));
  OAI21X1  g03807(.A0(new_n3871_), .A1(new_n3867_), .B0(new_n3865_), .Y(new_n3872_));
  XOR2X1   g03808(.A(new_n3511_), .B(new_n3507_), .Y(new_n3873_));
  AND2X1   g03809(.A(new_n3873_), .B(new_n3872_), .Y(new_n3874_));
  XOR2X1   g03810(.A(new_n3873_), .B(new_n3872_), .Y(new_n3875_));
  AOI22X1  g03811(.A0(new_n2423_), .A1(new_n1822_), .B0(new_n2418_), .B1(new_n1126_), .Y(new_n3876_));
  OAI21X1  g03812(.A0(new_n2666_), .A1(new_n1189_), .B0(new_n3876_), .Y(new_n3877_));
  AOI21X1  g03813(.A0(new_n2963_), .A1(new_n2301_), .B0(new_n3877_), .Y(new_n3878_));
  XOR2X1   g03814(.A(new_n3878_), .B(new_n89_), .Y(new_n3879_));
  AOI21X1  g03815(.A0(new_n3879_), .A1(new_n3875_), .B0(new_n3874_), .Y(new_n3880_));
  NOR2X1   g03816(.A(new_n3880_), .B(new_n3661_), .Y(new_n3881_));
  XOR2X1   g03817(.A(new_n3880_), .B(new_n3661_), .Y(new_n3882_));
  AOI22X1  g03818(.A0(new_n2745_), .A1(new_n2481_), .B0(new_n2657_), .B1(new_n2835_), .Y(new_n3883_));
  OAI21X1  g03819(.A0(new_n2743_), .A1(new_n903_), .B0(new_n3883_), .Y(new_n3884_));
  AOI21X1  g03820(.A0(new_n2709_), .A1(new_n2658_), .B0(new_n3884_), .Y(new_n3885_));
  XOR2X1   g03821(.A(new_n3885_), .B(new_n70_), .Y(new_n3886_));
  AOI21X1  g03822(.A0(new_n3886_), .A1(new_n3882_), .B0(new_n3881_), .Y(new_n3887_));
  NOR2X1   g03823(.A(new_n3887_), .B(new_n3659_), .Y(new_n3888_));
  AOI21X1  g03824(.A0(new_n3658_), .A1(new_n3657_), .B0(new_n3888_), .Y(new_n3889_));
  NOR2X1   g03825(.A(new_n3889_), .B(new_n3652_), .Y(new_n3890_));
  XOR2X1   g03826(.A(new_n3889_), .B(new_n3652_), .Y(new_n3891_));
  AOI22X1  g03827(.A0(new_n3146_), .A1(new_n1887_), .B0(new_n2875_), .B1(new_n1886_), .Y(new_n3892_));
  OAI21X1  g03828(.A0(new_n3144_), .A1(new_n520_), .B0(new_n3892_), .Y(new_n3893_));
  AOI21X1  g03829(.A0(new_n2876_), .A1(new_n1882_), .B0(new_n3893_), .Y(new_n3894_));
  XOR2X1   g03830(.A(new_n3894_), .B(new_n1920_), .Y(new_n3895_));
  AOI21X1  g03831(.A0(new_n3895_), .A1(new_n3891_), .B0(new_n3890_), .Y(new_n3896_));
  NOR2X1   g03832(.A(new_n3896_), .B(new_n3650_), .Y(new_n3897_));
  XOR2X1   g03833(.A(new_n3896_), .B(new_n3650_), .Y(new_n3898_));
  AOI22X1  g03834(.A0(new_n3546_), .A1(new_n2627_), .B0(new_n3232_), .B1(new_n2093_), .Y(new_n3899_));
  OAI21X1  g03835(.A0(new_n3389_), .A1(new_n2137_), .B0(new_n3899_), .Y(new_n3900_));
  AOI21X1  g03836(.A0(new_n3234_), .A1(new_n2294_), .B0(new_n3900_), .Y(new_n3901_));
  XOR2X1   g03837(.A(new_n3901_), .B(new_n2445_), .Y(new_n3902_));
  AOI21X1  g03838(.A0(new_n3902_), .A1(new_n3898_), .B0(new_n3897_), .Y(new_n3903_));
  NOR2X1   g03839(.A(new_n3903_), .B(new_n3649_), .Y(new_n3904_));
  AOI21X1  g03840(.A0(new_n3648_), .A1(new_n3647_), .B0(new_n3904_), .Y(new_n3905_));
  INVX1    g03841(.A(new_n3624_), .Y(new_n3906_));
  NAND2X1  g03842(.A(new_n3625_), .B(new_n3621_), .Y(new_n3907_));
  INVX1    g03843(.A(new_n3907_), .Y(new_n3908_));
  AOI22X1  g03844(.A0(new_n3908_), .A1(new_n2649_), .B0(new_n3628_), .B1(new_n2421_), .Y(new_n3909_));
  OAI21X1  g03845(.A0(new_n3906_), .A1(new_n2695_), .B0(new_n3909_), .Y(new_n3910_));
  XOR2X1   g03846(.A(new_n3910_), .B(new_n2529_), .Y(new_n3911_));
  NOR2X1   g03847(.A(new_n3911_), .B(new_n3905_), .Y(new_n3912_));
  XOR2X1   g03848(.A(new_n3618_), .B(new_n3614_), .Y(new_n3913_));
  XOR2X1   g03849(.A(new_n3911_), .B(new_n3905_), .Y(new_n3914_));
  AOI21X1  g03850(.A0(new_n3914_), .A1(new_n3913_), .B0(new_n3912_), .Y(new_n3915_));
  NOR2X1   g03851(.A(new_n3915_), .B(new_n3642_), .Y(new_n3916_));
  XOR2X1   g03852(.A(new_n3915_), .B(new_n3642_), .Y(new_n3917_));
  XOR2X1   g03853(.A(new_n3902_), .B(new_n3898_), .Y(new_n3918_));
  INVX1    g03854(.A(new_n3918_), .Y(new_n3919_));
  XOR2X1   g03855(.A(new_n3895_), .B(new_n3891_), .Y(new_n3920_));
  INVX1    g03856(.A(new_n3920_), .Y(new_n3921_));
  INVX1    g03857(.A(new_n3659_), .Y(new_n3922_));
  XOR2X1   g03858(.A(new_n3887_), .B(new_n3922_), .Y(new_n3923_));
  OAI22X1  g03859(.A0(new_n3152_), .A1(new_n520_), .B0(new_n3250_), .B1(new_n690_), .Y(new_n3924_));
  AOI21X1  g03860(.A0(new_n3099_), .A1(new_n1886_), .B0(new_n3924_), .Y(new_n3925_));
  OAI21X1  g03861(.A0(new_n3098_), .A1(new_n3114_), .B0(new_n3925_), .Y(new_n3926_));
  XOR2X1   g03862(.A(new_n3926_), .B(new_n1920_), .Y(new_n3927_));
  NOR2X1   g03863(.A(new_n3927_), .B(new_n3923_), .Y(new_n3928_));
  XOR2X1   g03864(.A(new_n3886_), .B(new_n3882_), .Y(new_n3929_));
  INVX1    g03865(.A(new_n3929_), .Y(new_n3930_));
  XOR2X1   g03866(.A(new_n3878_), .B(\a[26] ), .Y(new_n3931_));
  XOR2X1   g03867(.A(new_n3931_), .B(new_n3875_), .Y(new_n3932_));
  XOR2X1   g03868(.A(new_n3871_), .B(new_n3866_), .Y(new_n3933_));
  INVX1    g03869(.A(new_n2976_), .Y(new_n3934_));
  OAI22X1  g03870(.A0(new_n2666_), .A1(new_n1236_), .B0(new_n2626_), .B1(new_n1127_), .Y(new_n3935_));
  AOI21X1  g03871(.A0(new_n2418_), .A1(new_n1187_), .B0(new_n3935_), .Y(new_n3936_));
  OAI21X1  g03872(.A0(new_n3934_), .A1(new_n2665_), .B0(new_n3936_), .Y(new_n3937_));
  XOR2X1   g03873(.A(new_n3937_), .B(new_n89_), .Y(new_n3938_));
  NOR2X1   g03874(.A(new_n3938_), .B(new_n3933_), .Y(new_n3939_));
  XOR2X1   g03875(.A(new_n3862_), .B(new_n3859_), .Y(new_n3940_));
  INVX1    g03876(.A(new_n3425_), .Y(new_n3941_));
  OAI22X1  g03877(.A0(new_n2140_), .A1(new_n1339_), .B0(new_n2431_), .B1(new_n1358_), .Y(new_n3942_));
  AOI21X1  g03878(.A0(new_n2185_), .A1(new_n3850_), .B0(new_n3942_), .Y(new_n3943_));
  OAI21X1  g03879(.A0(new_n3941_), .A1(new_n2063_), .B0(new_n3943_), .Y(new_n3944_));
  XOR2X1   g03880(.A(new_n3944_), .B(new_n74_), .Y(new_n3945_));
  OR2X1    g03881(.A(new_n3945_), .B(new_n3940_), .Y(new_n3946_));
  AND2X1   g03882(.A(new_n3945_), .B(new_n3940_), .Y(new_n3947_));
  AOI22X1  g03883(.A0(new_n2423_), .A1(new_n1187_), .B0(new_n2418_), .B1(new_n2977_), .Y(new_n3948_));
  OAI21X1  g03884(.A0(new_n2666_), .A1(new_n1294_), .B0(new_n3948_), .Y(new_n3949_));
  AOI21X1  g03885(.A0(new_n3189_), .A1(new_n2301_), .B0(new_n3949_), .Y(new_n3950_));
  XOR2X1   g03886(.A(new_n3950_), .B(\a[26] ), .Y(new_n3951_));
  OAI21X1  g03887(.A0(new_n3951_), .A1(new_n3947_), .B0(new_n3946_), .Y(new_n3952_));
  XOR2X1   g03888(.A(new_n3938_), .B(new_n3933_), .Y(new_n3953_));
  AOI21X1  g03889(.A0(new_n3953_), .A1(new_n3952_), .B0(new_n3939_), .Y(new_n3954_));
  NOR2X1   g03890(.A(new_n3954_), .B(new_n3932_), .Y(new_n3955_));
  XOR2X1   g03891(.A(new_n3954_), .B(new_n3932_), .Y(new_n3956_));
  AOI22X1  g03892(.A0(new_n2745_), .A1(new_n2602_), .B0(new_n2657_), .B1(new_n2603_), .Y(new_n3957_));
  OAI21X1  g03893(.A0(new_n2743_), .A1(new_n957_), .B0(new_n3957_), .Y(new_n3958_));
  AOI21X1  g03894(.A0(new_n2658_), .A1(new_n2601_), .B0(new_n3958_), .Y(new_n3959_));
  XOR2X1   g03895(.A(new_n3959_), .B(new_n70_), .Y(new_n3960_));
  AOI21X1  g03896(.A0(new_n3960_), .A1(new_n3956_), .B0(new_n3955_), .Y(new_n3961_));
  OR2X1    g03897(.A(new_n3961_), .B(new_n3930_), .Y(new_n3962_));
  XOR2X1   g03898(.A(new_n3961_), .B(new_n3930_), .Y(new_n3963_));
  INVX1    g03899(.A(new_n3963_), .Y(new_n3964_));
  AOI22X1  g03900(.A0(new_n3146_), .A1(new_n1886_), .B0(new_n2875_), .B1(new_n2036_), .Y(new_n3965_));
  OAI21X1  g03901(.A0(new_n3144_), .A1(new_n690_), .B0(new_n3965_), .Y(new_n3966_));
  AOI21X1  g03902(.A0(new_n2876_), .A1(new_n2035_), .B0(new_n3966_), .Y(new_n3967_));
  XOR2X1   g03903(.A(new_n3967_), .B(\a[20] ), .Y(new_n3968_));
  OAI21X1  g03904(.A0(new_n3968_), .A1(new_n3964_), .B0(new_n3962_), .Y(new_n3969_));
  XOR2X1   g03905(.A(new_n3927_), .B(new_n3923_), .Y(new_n3970_));
  AOI21X1  g03906(.A0(new_n3970_), .A1(new_n3969_), .B0(new_n3928_), .Y(new_n3971_));
  NOR2X1   g03907(.A(new_n3971_), .B(new_n3921_), .Y(new_n3972_));
  XOR2X1   g03908(.A(new_n3971_), .B(new_n3921_), .Y(new_n3973_));
  AOI22X1  g03909(.A0(new_n3546_), .A1(new_n2252_), .B0(new_n3232_), .B1(new_n2246_), .Y(new_n3974_));
  OAI21X1  g03910(.A0(new_n3389_), .A1(new_n2092_), .B0(new_n3974_), .Y(new_n3975_));
  AOI21X1  g03911(.A0(new_n3234_), .A1(new_n2201_), .B0(new_n3975_), .Y(new_n3976_));
  XOR2X1   g03912(.A(new_n3976_), .B(new_n2445_), .Y(new_n3977_));
  AOI21X1  g03913(.A0(new_n3977_), .A1(new_n3973_), .B0(new_n3972_), .Y(new_n3978_));
  NOR2X1   g03914(.A(new_n3978_), .B(new_n3919_), .Y(new_n3979_));
  INVX1    g03915(.A(new_n3979_), .Y(new_n3980_));
  XOR2X1   g03916(.A(new_n3978_), .B(new_n3919_), .Y(new_n3981_));
  INVX1    g03917(.A(new_n3981_), .Y(new_n3982_));
  OR2X1    g03918(.A(new_n3622_), .B(new_n3621_), .Y(new_n3983_));
  INVX1    g03919(.A(new_n3983_), .Y(new_n3984_));
  AOI22X1  g03920(.A0(new_n3984_), .A1(new_n2421_), .B0(new_n3628_), .B1(new_n2420_), .Y(new_n3985_));
  OAI21X1  g03921(.A0(new_n3907_), .A1(new_n2379_), .B0(new_n3985_), .Y(new_n3986_));
  AOI21X1  g03922(.A0(new_n3624_), .A1(new_n2416_), .B0(new_n3986_), .Y(new_n3987_));
  XOR2X1   g03923(.A(new_n3987_), .B(\a[14] ), .Y(new_n3988_));
  OAI21X1  g03924(.A0(new_n3988_), .A1(new_n3982_), .B0(new_n3980_), .Y(new_n3989_));
  OAI22X1  g03925(.A0(new_n3983_), .A1(new_n2648_), .B0(new_n3907_), .B1(new_n2414_), .Y(new_n3990_));
  AOI21X1  g03926(.A0(new_n3628_), .A1(new_n2752_), .B0(new_n3990_), .Y(new_n3991_));
  OAI21X1  g03927(.A0(new_n3906_), .A1(new_n2757_), .B0(new_n3991_), .Y(new_n3992_));
  XOR2X1   g03928(.A(new_n3992_), .B(\a[14] ), .Y(new_n3993_));
  XOR2X1   g03929(.A(new_n3903_), .B(new_n3649_), .Y(new_n3994_));
  INVX1    g03930(.A(new_n3994_), .Y(new_n3995_));
  XOR2X1   g03931(.A(new_n3992_), .B(new_n2529_), .Y(new_n3996_));
  XOR2X1   g03932(.A(new_n3996_), .B(new_n3989_), .Y(new_n3997_));
  NOR2X1   g03933(.A(new_n3997_), .B(new_n3995_), .Y(new_n3998_));
  AOI21X1  g03934(.A0(new_n3993_), .A1(new_n3989_), .B0(new_n3998_), .Y(new_n3999_));
  INVX1    g03935(.A(new_n3999_), .Y(new_n4000_));
  XOR2X1   g03936(.A(new_n3914_), .B(new_n3913_), .Y(new_n4001_));
  AND2X1   g03937(.A(new_n4001_), .B(new_n4000_), .Y(new_n4002_));
  INVX1    g03938(.A(new_n4002_), .Y(new_n4003_));
  XOR2X1   g03939(.A(new_n3977_), .B(new_n3973_), .Y(new_n4004_));
  AOI22X1  g03940(.A0(new_n3546_), .A1(new_n2093_), .B0(new_n3232_), .B1(new_n1887_), .Y(new_n4005_));
  OAI21X1  g03941(.A0(new_n3389_), .A1(new_n2183_), .B0(new_n4005_), .Y(new_n4006_));
  AOI21X1  g03942(.A0(new_n3234_), .A1(new_n2430_), .B0(new_n4006_), .Y(new_n4007_));
  XOR2X1   g03943(.A(new_n4007_), .B(\a[17] ), .Y(new_n4008_));
  INVX1    g03944(.A(new_n4008_), .Y(new_n4009_));
  XOR2X1   g03945(.A(new_n3970_), .B(new_n3969_), .Y(new_n4010_));
  AND2X1   g03946(.A(new_n4010_), .B(new_n4009_), .Y(new_n4011_));
  XOR2X1   g03947(.A(new_n4010_), .B(new_n4008_), .Y(new_n4012_));
  XOR2X1   g03948(.A(new_n3968_), .B(new_n3963_), .Y(new_n4013_));
  XOR2X1   g03949(.A(new_n3960_), .B(new_n3956_), .Y(new_n4014_));
  INVX1    g03950(.A(new_n4014_), .Y(new_n4015_));
  INVX1    g03951(.A(new_n2657_), .Y(new_n4016_));
  AOI22X1  g03952(.A0(new_n2745_), .A1(new_n2835_), .B0(new_n2696_), .B1(new_n2603_), .Y(new_n4017_));
  OAI21X1  g03953(.A0(new_n4016_), .A1(new_n1065_), .B0(new_n4017_), .Y(new_n4018_));
  AOI21X1  g03954(.A0(new_n2834_), .A1(new_n2658_), .B0(new_n4018_), .Y(new_n4019_));
  XOR2X1   g03955(.A(new_n4019_), .B(\a[23] ), .Y(new_n4020_));
  INVX1    g03956(.A(new_n4020_), .Y(new_n4021_));
  XOR2X1   g03957(.A(new_n3953_), .B(new_n3952_), .Y(new_n4022_));
  XOR2X1   g03958(.A(new_n4022_), .B(new_n4020_), .Y(new_n4023_));
  XOR2X1   g03959(.A(new_n3945_), .B(new_n3940_), .Y(new_n4024_));
  XOR2X1   g03960(.A(new_n3951_), .B(new_n4024_), .Y(new_n4025_));
  XOR2X1   g03961(.A(new_n3858_), .B(new_n3856_), .Y(new_n4026_));
  INVX1    g03962(.A(new_n4026_), .Y(new_n4027_));
  INVX1    g03963(.A(new_n3326_), .Y(new_n4028_));
  OAI22X1  g03964(.A0(new_n2186_), .A1(new_n1423_), .B0(new_n2140_), .B1(new_n1358_), .Y(new_n4029_));
  AOI21X1  g03965(.A0(new_n2095_), .A1(new_n3850_), .B0(new_n4029_), .Y(new_n4030_));
  OAI21X1  g03966(.A0(new_n4028_), .A1(new_n2063_), .B0(new_n4030_), .Y(new_n4031_));
  XOR2X1   g03967(.A(new_n4031_), .B(new_n74_), .Y(new_n4032_));
  NOR2X1   g03968(.A(new_n4032_), .B(new_n4027_), .Y(new_n4033_));
  XOR2X1   g03969(.A(new_n4032_), .B(new_n4027_), .Y(new_n4034_));
  AOI22X1  g03970(.A0(new_n2424_), .A1(new_n3055_), .B0(new_n2423_), .B1(new_n2977_), .Y(new_n4035_));
  OAI21X1  g03971(.A0(new_n2419_), .A1(new_n1294_), .B0(new_n4035_), .Y(new_n4036_));
  AOI21X1  g03972(.A0(new_n3054_), .A1(new_n2301_), .B0(new_n4036_), .Y(new_n4037_));
  XOR2X1   g03973(.A(new_n4037_), .B(new_n89_), .Y(new_n4038_));
  AOI21X1  g03974(.A0(new_n4038_), .A1(new_n4034_), .B0(new_n4033_), .Y(new_n4039_));
  NOR2X1   g03975(.A(new_n4039_), .B(new_n4025_), .Y(new_n4040_));
  XOR2X1   g03976(.A(new_n4039_), .B(new_n4025_), .Y(new_n4041_));
  AOI22X1  g03977(.A0(new_n2745_), .A1(new_n2603_), .B0(new_n2657_), .B1(new_n1126_), .Y(new_n4042_));
  OAI21X1  g03978(.A0(new_n2743_), .A1(new_n1065_), .B0(new_n4042_), .Y(new_n4043_));
  AOI21X1  g03979(.A0(new_n2824_), .A1(new_n2658_), .B0(new_n4043_), .Y(new_n4044_));
  XOR2X1   g03980(.A(new_n4044_), .B(new_n70_), .Y(new_n4045_));
  AOI21X1  g03981(.A0(new_n4045_), .A1(new_n4041_), .B0(new_n4040_), .Y(new_n4046_));
  NOR2X1   g03982(.A(new_n4046_), .B(new_n4023_), .Y(new_n4047_));
  AOI21X1  g03983(.A0(new_n4022_), .A1(new_n4021_), .B0(new_n4047_), .Y(new_n4048_));
  NOR2X1   g03984(.A(new_n4048_), .B(new_n4015_), .Y(new_n4049_));
  XOR2X1   g03985(.A(new_n4048_), .B(new_n4015_), .Y(new_n4050_));
  AOI22X1  g03986(.A0(new_n3146_), .A1(new_n2049_), .B0(new_n2875_), .B1(new_n2481_), .Y(new_n4051_));
  OAI21X1  g03987(.A0(new_n3144_), .A1(new_n783_), .B0(new_n4051_), .Y(new_n4052_));
  AOI21X1  g03988(.A0(new_n2876_), .A1(new_n2480_), .B0(new_n4052_), .Y(new_n4053_));
  XOR2X1   g03989(.A(new_n4053_), .B(new_n1920_), .Y(new_n4054_));
  AOI21X1  g03990(.A0(new_n4054_), .A1(new_n4050_), .B0(new_n4049_), .Y(new_n4055_));
  NOR2X1   g03991(.A(new_n4055_), .B(new_n4013_), .Y(new_n4056_));
  XOR2X1   g03992(.A(new_n4055_), .B(new_n4013_), .Y(new_n4057_));
  AOI22X1  g03993(.A0(new_n3546_), .A1(new_n2246_), .B0(new_n3232_), .B1(new_n2048_), .Y(new_n4058_));
  OAI21X1  g03994(.A0(new_n3389_), .A1(new_n1879_), .B0(new_n4058_), .Y(new_n4059_));
  AOI21X1  g03995(.A0(new_n3234_), .A1(new_n2244_), .B0(new_n4059_), .Y(new_n4060_));
  XOR2X1   g03996(.A(new_n4060_), .B(new_n2445_), .Y(new_n4061_));
  AOI21X1  g03997(.A0(new_n4061_), .A1(new_n4057_), .B0(new_n4056_), .Y(new_n4062_));
  NOR2X1   g03998(.A(new_n4062_), .B(new_n4012_), .Y(new_n4063_));
  OAI21X1  g03999(.A0(new_n4063_), .A1(new_n4011_), .B0(new_n4004_), .Y(new_n4064_));
  NOR2X1   g04000(.A(new_n4063_), .B(new_n4011_), .Y(new_n4065_));
  XOR2X1   g04001(.A(new_n4065_), .B(new_n4004_), .Y(new_n4066_));
  AOI22X1  g04002(.A0(new_n3908_), .A1(new_n2420_), .B0(new_n3628_), .B1(new_n2627_), .Y(new_n4067_));
  OAI21X1  g04003(.A0(new_n3983_), .A1(new_n2379_), .B0(new_n4067_), .Y(new_n4068_));
  AOI21X1  g04004(.A0(new_n3624_), .A1(new_n2625_), .B0(new_n4068_), .Y(new_n4069_));
  XOR2X1   g04005(.A(new_n4069_), .B(\a[14] ), .Y(new_n4070_));
  OR2X1    g04006(.A(new_n4070_), .B(new_n4066_), .Y(new_n4071_));
  AND2X1   g04007(.A(new_n4071_), .B(new_n4064_), .Y(new_n4072_));
  XOR2X1   g04008(.A(\a[9] ), .B(new_n2995_), .Y(new_n4073_));
  XOR2X1   g04009(.A(\a[10] ), .B(\a[9] ), .Y(new_n4074_));
  INVX1    g04010(.A(new_n4074_), .Y(new_n4075_));
  XOR2X1   g04011(.A(\a[11] ), .B(\a[10] ), .Y(new_n4076_));
  NAND3X1  g04012(.A(new_n4076_), .B(new_n4075_), .C(new_n4073_), .Y(new_n4077_));
  INVX1    g04013(.A(new_n4077_), .Y(new_n4078_));
  INVX1    g04014(.A(new_n4073_), .Y(new_n4079_));
  AND2X1   g04015(.A(new_n4076_), .B(new_n4079_), .Y(new_n4080_));
  AOI22X1  g04016(.A0(new_n4080_), .A1(new_n2652_), .B0(new_n4078_), .B1(new_n2649_), .Y(new_n4081_));
  XOR2X1   g04017(.A(new_n4081_), .B(\a[11] ), .Y(new_n4082_));
  NOR2X1   g04018(.A(new_n4082_), .B(new_n4072_), .Y(new_n4083_));
  XOR2X1   g04019(.A(new_n3988_), .B(new_n3981_), .Y(new_n4084_));
  INVX1    g04020(.A(new_n4084_), .Y(new_n4085_));
  XOR2X1   g04021(.A(new_n4082_), .B(new_n4072_), .Y(new_n4086_));
  AOI21X1  g04022(.A0(new_n4086_), .A1(new_n4085_), .B0(new_n4083_), .Y(new_n4087_));
  INVX1    g04023(.A(new_n4087_), .Y(new_n4088_));
  OR2X1    g04024(.A(new_n3996_), .B(new_n3989_), .Y(new_n4089_));
  AOI21X1  g04025(.A0(new_n3996_), .A1(new_n3989_), .B0(new_n3994_), .Y(new_n4090_));
  AOI21X1  g04026(.A0(new_n4090_), .A1(new_n4089_), .B0(new_n3998_), .Y(new_n4091_));
  AND2X1   g04027(.A(new_n4091_), .B(new_n4088_), .Y(new_n4092_));
  XOR2X1   g04028(.A(new_n4086_), .B(new_n4084_), .Y(new_n4093_));
  XOR2X1   g04029(.A(new_n4062_), .B(new_n4012_), .Y(new_n4094_));
  INVX1    g04030(.A(new_n4094_), .Y(new_n4095_));
  OAI22X1  g04031(.A0(new_n3983_), .A1(new_n2339_), .B0(new_n3627_), .B1(new_n2137_), .Y(new_n4096_));
  AOI21X1  g04032(.A0(new_n3908_), .A1(new_n2627_), .B0(new_n4096_), .Y(new_n4097_));
  OAI21X1  g04033(.A0(new_n3906_), .A1(new_n2670_), .B0(new_n4097_), .Y(new_n4098_));
  XOR2X1   g04034(.A(new_n4098_), .B(new_n2529_), .Y(new_n4099_));
  NOR2X1   g04035(.A(new_n4099_), .B(new_n4095_), .Y(new_n4100_));
  XOR2X1   g04036(.A(new_n4061_), .B(new_n4057_), .Y(new_n4101_));
  INVX1    g04037(.A(new_n4101_), .Y(new_n4102_));
  XOR2X1   g04038(.A(new_n4054_), .B(new_n4050_), .Y(new_n4103_));
  INVX1    g04039(.A(new_n4103_), .Y(new_n4104_));
  INVX1    g04040(.A(new_n4023_), .Y(new_n4105_));
  XOR2X1   g04041(.A(new_n4046_), .B(new_n4105_), .Y(new_n4106_));
  OAI22X1  g04042(.A0(new_n3152_), .A1(new_n783_), .B0(new_n3250_), .B1(new_n903_), .Y(new_n4107_));
  AOI21X1  g04043(.A0(new_n3099_), .A1(new_n2481_), .B0(new_n4107_), .Y(new_n4108_));
  OAI21X1  g04044(.A0(new_n3098_), .A1(new_n3261_), .B0(new_n4108_), .Y(new_n4109_));
  XOR2X1   g04045(.A(new_n4109_), .B(new_n1920_), .Y(new_n4110_));
  NOR2X1   g04046(.A(new_n4110_), .B(new_n4106_), .Y(new_n4111_));
  XOR2X1   g04047(.A(new_n4045_), .B(new_n4041_), .Y(new_n4112_));
  INVX1    g04048(.A(new_n4112_), .Y(new_n4113_));
  XOR2X1   g04049(.A(new_n4038_), .B(new_n4034_), .Y(new_n4114_));
  INVX1    g04050(.A(new_n4114_), .Y(new_n4115_));
  INVX1    g04051(.A(new_n3845_), .Y(new_n4116_));
  XOR2X1   g04052(.A(new_n4116_), .B(new_n3844_), .Y(new_n4117_));
  OAI22X1  g04053(.A0(new_n2186_), .A1(new_n3669_), .B0(new_n2140_), .B1(new_n1423_), .Y(new_n4118_));
  AOI21X1  g04054(.A0(new_n2095_), .A1(new_n1800_), .B0(new_n4118_), .Y(new_n4119_));
  OAI21X1  g04055(.A0(new_n3667_), .A1(new_n2063_), .B0(new_n4119_), .Y(new_n4120_));
  XOR2X1   g04056(.A(new_n4120_), .B(new_n74_), .Y(new_n4121_));
  XOR2X1   g04057(.A(new_n3843_), .B(new_n3840_), .Y(new_n4122_));
  OAI22X1  g04058(.A0(new_n2140_), .A1(new_n1465_), .B0(new_n2431_), .B1(new_n3669_), .Y(new_n4123_));
  AOI21X1  g04059(.A0(new_n2185_), .A1(new_n1536_), .B0(new_n4123_), .Y(new_n4124_));
  OAI21X1  g04060(.A0(new_n3676_), .A1(new_n2063_), .B0(new_n4124_), .Y(new_n4125_));
  XOR2X1   g04061(.A(new_n4125_), .B(new_n74_), .Y(new_n4126_));
  NOR2X1   g04062(.A(new_n4126_), .B(new_n4122_), .Y(new_n4127_));
  AOI22X1  g04063(.A0(new_n2185_), .A1(new_n3480_), .B0(new_n2139_), .B1(new_n1490_), .Y(new_n4128_));
  OAI21X1  g04064(.A0(new_n2431_), .A1(new_n1795_), .B0(new_n4128_), .Y(new_n4129_));
  AOI21X1  g04065(.A0(new_n3479_), .A1(new_n2062_), .B0(new_n4129_), .Y(new_n4130_));
  XOR2X1   g04066(.A(new_n4130_), .B(\a[29] ), .Y(new_n4131_));
  INVX1    g04067(.A(new_n3839_), .Y(new_n4132_));
  XOR2X1   g04068(.A(new_n4132_), .B(new_n3838_), .Y(new_n4133_));
  NOR2X1   g04069(.A(new_n4133_), .B(new_n4131_), .Y(new_n4134_));
  INVX1    g04070(.A(new_n4134_), .Y(new_n4135_));
  XOR2X1   g04071(.A(new_n4133_), .B(new_n4131_), .Y(new_n4136_));
  INVX1    g04072(.A(new_n4136_), .Y(new_n4137_));
  AOI22X1  g04073(.A0(new_n2139_), .A1(new_n1536_), .B0(new_n2095_), .B1(new_n3480_), .Y(new_n4138_));
  OAI21X1  g04074(.A0(new_n2186_), .A1(new_n1621_), .B0(new_n4138_), .Y(new_n4139_));
  AOI21X1  g04075(.A0(new_n3697_), .A1(new_n2062_), .B0(new_n4139_), .Y(new_n4140_));
  XOR2X1   g04076(.A(new_n4140_), .B(\a[29] ), .Y(new_n4141_));
  XOR2X1   g04077(.A(new_n3837_), .B(new_n3835_), .Y(new_n4142_));
  NOR2X1   g04078(.A(new_n4142_), .B(new_n4141_), .Y(new_n4143_));
  XOR2X1   g04079(.A(new_n4142_), .B(new_n4141_), .Y(new_n4144_));
  AOI22X1  g04080(.A0(new_n2185_), .A1(new_n3721_), .B0(new_n2139_), .B1(new_n3480_), .Y(new_n4145_));
  OAI21X1  g04081(.A0(new_n2431_), .A1(new_n1621_), .B0(new_n4145_), .Y(new_n4146_));
  AOI21X1  g04082(.A0(new_n3720_), .A1(new_n2062_), .B0(new_n4146_), .Y(new_n4147_));
  XOR2X1   g04083(.A(new_n4147_), .B(\a[29] ), .Y(new_n4148_));
  XOR2X1   g04084(.A(new_n3834_), .B(new_n3832_), .Y(new_n4149_));
  OR2X1    g04085(.A(new_n4149_), .B(new_n4148_), .Y(new_n4150_));
  XOR2X1   g04086(.A(new_n4149_), .B(new_n4148_), .Y(new_n4151_));
  INVX1    g04087(.A(new_n4151_), .Y(new_n4152_));
  AOI22X1  g04088(.A0(new_n2185_), .A1(new_n1676_), .B0(new_n2095_), .B1(new_n3721_), .Y(new_n4153_));
  OAI21X1  g04089(.A0(new_n2140_), .A1(new_n1621_), .B0(new_n4153_), .Y(new_n4154_));
  AOI21X1  g04090(.A0(new_n3745_), .A1(new_n2062_), .B0(new_n4154_), .Y(new_n4155_));
  XOR2X1   g04091(.A(new_n4155_), .B(\a[29] ), .Y(new_n4156_));
  INVX1    g04092(.A(new_n3818_), .Y(new_n4157_));
  XOR2X1   g04093(.A(new_n3826_), .B(new_n4157_), .Y(new_n4158_));
  NOR2X1   g04094(.A(new_n4158_), .B(new_n4156_), .Y(new_n4159_));
  XOR2X1   g04095(.A(new_n4158_), .B(new_n4156_), .Y(new_n4160_));
  AOI22X1  g04096(.A0(new_n2139_), .A1(new_n3721_), .B0(new_n2095_), .B1(new_n1676_), .Y(new_n4161_));
  OAI21X1  g04097(.A0(new_n2186_), .A1(new_n1708_), .B0(new_n4161_), .Y(new_n4162_));
  AOI21X1  g04098(.A0(new_n3774_), .A1(new_n2062_), .B0(new_n4162_), .Y(new_n4163_));
  XOR2X1   g04099(.A(new_n4163_), .B(\a[29] ), .Y(new_n4164_));
  XOR2X1   g04100(.A(new_n1784_), .B(new_n1735_), .Y(new_n4165_));
  OAI22X1  g04101(.A0(new_n3498_), .A1(new_n1735_), .B0(new_n1885_), .B1(new_n1784_), .Y(new_n4166_));
  AOI21X1  g04102(.A0(new_n4165_), .A1(new_n407_), .B0(new_n4166_), .Y(new_n4167_));
  OR2X1    g04103(.A(new_n4167_), .B(new_n4164_), .Y(new_n4168_));
  XOR2X1   g04104(.A(new_n4167_), .B(new_n4164_), .Y(new_n4169_));
  INVX1    g04105(.A(new_n4169_), .Y(new_n4170_));
  XOR2X1   g04106(.A(\a[30] ), .B(new_n74_), .Y(new_n4171_));
  NOR2X1   g04107(.A(new_n4171_), .B(new_n1784_), .Y(new_n4172_));
  OAI22X1  g04108(.A0(new_n2140_), .A1(new_n1735_), .B0(new_n2431_), .B1(new_n1784_), .Y(new_n4173_));
  AOI21X1  g04109(.A0(new_n4165_), .A1(new_n2062_), .B0(new_n4173_), .Y(new_n4174_));
  XOR2X1   g04110(.A(new_n4174_), .B(\a[29] ), .Y(new_n4175_));
  AND2X1   g04111(.A(new_n2184_), .B(new_n3821_), .Y(new_n4176_));
  OR2X1    g04112(.A(new_n3822_), .B(new_n3820_), .Y(new_n4177_));
  OAI22X1  g04113(.A0(new_n2186_), .A1(new_n1784_), .B0(new_n2431_), .B1(new_n1735_), .Y(new_n4178_));
  AOI21X1  g04114(.A0(new_n2139_), .A1(new_n1706_), .B0(new_n4178_), .Y(new_n4179_));
  OAI21X1  g04115(.A0(new_n4177_), .A1(new_n2063_), .B0(new_n4179_), .Y(new_n4180_));
  NOR4X1   g04116(.A(new_n4180_), .B(new_n4176_), .C(new_n4175_), .D(new_n74_), .Y(new_n4181_));
  AOI22X1  g04117(.A0(new_n2185_), .A1(new_n3819_), .B0(new_n2139_), .B1(new_n1676_), .Y(new_n4182_));
  OAI21X1  g04118(.A0(new_n2431_), .A1(new_n1708_), .B0(new_n4182_), .Y(new_n4183_));
  AOI21X1  g04119(.A0(new_n3829_), .A1(new_n2062_), .B0(new_n4183_), .Y(new_n4184_));
  XOR2X1   g04120(.A(new_n4184_), .B(\a[29] ), .Y(new_n4185_));
  INVX1    g04121(.A(new_n4172_), .Y(new_n4186_));
  XOR2X1   g04122(.A(new_n4181_), .B(new_n4186_), .Y(new_n4187_));
  NOR2X1   g04123(.A(new_n4187_), .B(new_n4185_), .Y(new_n4188_));
  AOI21X1  g04124(.A0(new_n4181_), .A1(new_n4172_), .B0(new_n4188_), .Y(new_n4189_));
  OAI21X1  g04125(.A0(new_n4189_), .A1(new_n4170_), .B0(new_n4168_), .Y(new_n4190_));
  AOI21X1  g04126(.A0(new_n4190_), .A1(new_n4160_), .B0(new_n4159_), .Y(new_n4191_));
  OAI21X1  g04127(.A0(new_n4191_), .A1(new_n4152_), .B0(new_n4150_), .Y(new_n4192_));
  AOI21X1  g04128(.A0(new_n4192_), .A1(new_n4144_), .B0(new_n4143_), .Y(new_n4193_));
  OAI21X1  g04129(.A0(new_n4193_), .A1(new_n4137_), .B0(new_n4135_), .Y(new_n4194_));
  XOR2X1   g04130(.A(new_n4126_), .B(new_n4122_), .Y(new_n4195_));
  AOI21X1  g04131(.A0(new_n4195_), .A1(new_n4194_), .B0(new_n4127_), .Y(new_n4196_));
  INVX1    g04132(.A(new_n4196_), .Y(new_n4197_));
  XOR2X1   g04133(.A(new_n4121_), .B(new_n4117_), .Y(new_n4198_));
  NAND2X1  g04134(.A(new_n4198_), .B(new_n4197_), .Y(new_n4199_));
  OAI21X1  g04135(.A0(new_n4121_), .A1(new_n4117_), .B0(new_n4199_), .Y(new_n4200_));
  XOR2X1   g04136(.A(new_n3854_), .B(new_n3848_), .Y(new_n4201_));
  AND2X1   g04137(.A(new_n4201_), .B(new_n4200_), .Y(new_n4202_));
  AOI22X1  g04138(.A0(new_n2424_), .A1(new_n1357_), .B0(new_n2423_), .B1(new_n3342_), .Y(new_n4203_));
  OAI21X1  g04139(.A0(new_n2419_), .A1(new_n1339_), .B0(new_n4203_), .Y(new_n4204_));
  AOI21X1  g04140(.A0(new_n3341_), .A1(new_n2301_), .B0(new_n4204_), .Y(new_n4205_));
  XOR2X1   g04141(.A(new_n4205_), .B(new_n89_), .Y(new_n4206_));
  XOR2X1   g04142(.A(new_n4201_), .B(new_n4200_), .Y(new_n4207_));
  AOI21X1  g04143(.A0(new_n4207_), .A1(new_n4206_), .B0(new_n4202_), .Y(new_n4208_));
  NOR2X1   g04144(.A(new_n4208_), .B(new_n4115_), .Y(new_n4209_));
  XOR2X1   g04145(.A(new_n4208_), .B(new_n4115_), .Y(new_n4210_));
  AOI22X1  g04146(.A0(new_n2745_), .A1(new_n1822_), .B0(new_n2696_), .B1(new_n1126_), .Y(new_n4211_));
  OAI21X1  g04147(.A0(new_n4016_), .A1(new_n1189_), .B0(new_n4211_), .Y(new_n4212_));
  AOI21X1  g04148(.A0(new_n2963_), .A1(new_n2658_), .B0(new_n4212_), .Y(new_n4213_));
  XOR2X1   g04149(.A(new_n4213_), .B(\a[23] ), .Y(new_n4214_));
  INVX1    g04150(.A(new_n4214_), .Y(new_n4215_));
  AOI21X1  g04151(.A0(new_n4215_), .A1(new_n4210_), .B0(new_n4209_), .Y(new_n4216_));
  OR2X1    g04152(.A(new_n4216_), .B(new_n4113_), .Y(new_n4217_));
  XOR2X1   g04153(.A(new_n4216_), .B(new_n4113_), .Y(new_n4218_));
  INVX1    g04154(.A(new_n4218_), .Y(new_n4219_));
  AOI22X1  g04155(.A0(new_n3146_), .A1(new_n2481_), .B0(new_n2875_), .B1(new_n2835_), .Y(new_n4220_));
  OAI21X1  g04156(.A0(new_n3144_), .A1(new_n903_), .B0(new_n4220_), .Y(new_n4221_));
  AOI21X1  g04157(.A0(new_n2876_), .A1(new_n2709_), .B0(new_n4221_), .Y(new_n4222_));
  XOR2X1   g04158(.A(new_n4222_), .B(\a[20] ), .Y(new_n4223_));
  OAI21X1  g04159(.A0(new_n4223_), .A1(new_n4219_), .B0(new_n4217_), .Y(new_n4224_));
  XOR2X1   g04160(.A(new_n4110_), .B(new_n4106_), .Y(new_n4225_));
  AOI21X1  g04161(.A0(new_n4225_), .A1(new_n4224_), .B0(new_n4111_), .Y(new_n4226_));
  NOR2X1   g04162(.A(new_n4226_), .B(new_n4104_), .Y(new_n4227_));
  XOR2X1   g04163(.A(new_n4226_), .B(new_n4104_), .Y(new_n4228_));
  AOI22X1  g04164(.A0(new_n3546_), .A1(new_n1887_), .B0(new_n3232_), .B1(new_n1886_), .Y(new_n4229_));
  OAI21X1  g04165(.A0(new_n3389_), .A1(new_n520_), .B0(new_n4229_), .Y(new_n4230_));
  AOI21X1  g04166(.A0(new_n3234_), .A1(new_n1882_), .B0(new_n4230_), .Y(new_n4231_));
  XOR2X1   g04167(.A(new_n4231_), .B(new_n2445_), .Y(new_n4232_));
  AOI21X1  g04168(.A0(new_n4232_), .A1(new_n4228_), .B0(new_n4227_), .Y(new_n4233_));
  OR2X1    g04169(.A(new_n4233_), .B(new_n4102_), .Y(new_n4234_));
  XOR2X1   g04170(.A(new_n4233_), .B(new_n4102_), .Y(new_n4235_));
  INVX1    g04171(.A(new_n4235_), .Y(new_n4236_));
  AOI22X1  g04172(.A0(new_n3984_), .A1(new_n2627_), .B0(new_n3628_), .B1(new_n2093_), .Y(new_n4237_));
  OAI21X1  g04173(.A0(new_n3907_), .A1(new_n2137_), .B0(new_n4237_), .Y(new_n4238_));
  AOI21X1  g04174(.A0(new_n3624_), .A1(new_n2294_), .B0(new_n4238_), .Y(new_n4239_));
  XOR2X1   g04175(.A(new_n4239_), .B(\a[14] ), .Y(new_n4240_));
  OAI21X1  g04176(.A0(new_n4240_), .A1(new_n4236_), .B0(new_n4234_), .Y(new_n4241_));
  XOR2X1   g04177(.A(new_n4099_), .B(new_n4094_), .Y(new_n4242_));
  INVX1    g04178(.A(new_n4242_), .Y(new_n4243_));
  AOI21X1  g04179(.A0(new_n4243_), .A1(new_n4241_), .B0(new_n4100_), .Y(new_n4244_));
  INVX1    g04180(.A(new_n4080_), .Y(new_n4245_));
  NAND2X1  g04181(.A(new_n4074_), .B(new_n4073_), .Y(new_n4246_));
  INVX1    g04182(.A(new_n4246_), .Y(new_n4247_));
  AOI22X1  g04183(.A0(new_n4247_), .A1(new_n2649_), .B0(new_n4078_), .B1(new_n2421_), .Y(new_n4248_));
  OAI21X1  g04184(.A0(new_n4245_), .A1(new_n2695_), .B0(new_n4248_), .Y(new_n4249_));
  XOR2X1   g04185(.A(new_n4249_), .B(new_n2911_), .Y(new_n4250_));
  NOR2X1   g04186(.A(new_n4250_), .B(new_n4244_), .Y(new_n4251_));
  XOR2X1   g04187(.A(new_n4070_), .B(new_n4066_), .Y(new_n4252_));
  XOR2X1   g04188(.A(new_n4250_), .B(new_n4244_), .Y(new_n4253_));
  AOI21X1  g04189(.A0(new_n4253_), .A1(new_n4252_), .B0(new_n4251_), .Y(new_n4254_));
  NOR2X1   g04190(.A(new_n4254_), .B(new_n4093_), .Y(new_n4255_));
  INVX1    g04191(.A(new_n4255_), .Y(new_n4256_));
  XOR2X1   g04192(.A(new_n4254_), .B(new_n4093_), .Y(new_n4257_));
  INVX1    g04193(.A(new_n4257_), .Y(new_n4258_));
  XOR2X1   g04194(.A(new_n4240_), .B(new_n4235_), .Y(new_n4259_));
  XOR2X1   g04195(.A(new_n4232_), .B(new_n4228_), .Y(new_n4260_));
  INVX1    g04196(.A(new_n4260_), .Y(new_n4261_));
  AOI22X1  g04197(.A0(new_n3546_), .A1(new_n2048_), .B0(new_n3232_), .B1(new_n2049_), .Y(new_n4262_));
  OAI21X1  g04198(.A0(new_n3389_), .A1(new_n623_), .B0(new_n4262_), .Y(new_n4263_));
  AOI21X1  g04199(.A0(new_n3234_), .A1(new_n2047_), .B0(new_n4263_), .Y(new_n4264_));
  XOR2X1   g04200(.A(new_n4264_), .B(\a[17] ), .Y(new_n4265_));
  INVX1    g04201(.A(new_n4265_), .Y(new_n4266_));
  XOR2X1   g04202(.A(new_n4225_), .B(new_n4224_), .Y(new_n4267_));
  XOR2X1   g04203(.A(new_n4267_), .B(new_n4265_), .Y(new_n4268_));
  XOR2X1   g04204(.A(new_n4223_), .B(new_n4218_), .Y(new_n4269_));
  XOR2X1   g04205(.A(new_n4214_), .B(new_n4210_), .Y(new_n4270_));
  XOR2X1   g04206(.A(new_n4198_), .B(new_n4197_), .Y(new_n4271_));
  INVX1    g04207(.A(new_n4271_), .Y(new_n4272_));
  OAI22X1  g04208(.A0(new_n2626_), .A1(new_n1339_), .B0(new_n2419_), .B1(new_n1358_), .Y(new_n4273_));
  AOI21X1  g04209(.A0(new_n2424_), .A1(new_n3850_), .B0(new_n4273_), .Y(new_n4274_));
  OAI21X1  g04210(.A0(new_n3941_), .A1(new_n2665_), .B0(new_n4274_), .Y(new_n4275_));
  XOR2X1   g04211(.A(new_n4275_), .B(new_n89_), .Y(new_n4276_));
  OR2X1    g04212(.A(new_n4276_), .B(new_n4272_), .Y(new_n4277_));
  XOR2X1   g04213(.A(new_n4195_), .B(new_n4194_), .Y(new_n4278_));
  INVX1    g04214(.A(new_n4278_), .Y(new_n4279_));
  OAI22X1  g04215(.A0(new_n2666_), .A1(new_n1423_), .B0(new_n2626_), .B1(new_n1358_), .Y(new_n4280_));
  AOI21X1  g04216(.A0(new_n2418_), .A1(new_n3850_), .B0(new_n4280_), .Y(new_n4281_));
  OAI21X1  g04217(.A0(new_n4028_), .A1(new_n2665_), .B0(new_n4281_), .Y(new_n4282_));
  XOR2X1   g04218(.A(new_n4282_), .B(new_n89_), .Y(new_n4283_));
  NOR2X1   g04219(.A(new_n4283_), .B(new_n4279_), .Y(new_n4284_));
  INVX1    g04220(.A(new_n4284_), .Y(new_n4285_));
  XOR2X1   g04221(.A(new_n4193_), .B(new_n4137_), .Y(new_n4286_));
  INVX1    g04222(.A(new_n4286_), .Y(new_n4287_));
  OAI22X1  g04223(.A0(new_n2666_), .A1(new_n1465_), .B0(new_n2419_), .B1(new_n1423_), .Y(new_n4288_));
  AOI21X1  g04224(.A0(new_n2423_), .A1(new_n3850_), .B0(new_n4288_), .Y(new_n4289_));
  OAI21X1  g04225(.A0(new_n3849_), .A1(new_n2665_), .B0(new_n4289_), .Y(new_n4290_));
  XOR2X1   g04226(.A(new_n4290_), .B(new_n89_), .Y(new_n4291_));
  NOR2X1   g04227(.A(new_n4291_), .B(new_n4287_), .Y(new_n4292_));
  INVX1    g04228(.A(new_n4292_), .Y(new_n4293_));
  XOR2X1   g04229(.A(new_n4192_), .B(new_n4144_), .Y(new_n4294_));
  OAI22X1  g04230(.A0(new_n2666_), .A1(new_n3669_), .B0(new_n2626_), .B1(new_n1423_), .Y(new_n4295_));
  AOI21X1  g04231(.A0(new_n2418_), .A1(new_n1800_), .B0(new_n4295_), .Y(new_n4296_));
  OAI21X1  g04232(.A0(new_n3667_), .A1(new_n2665_), .B0(new_n4296_), .Y(new_n4297_));
  XOR2X1   g04233(.A(new_n4297_), .B(\a[26] ), .Y(new_n4298_));
  AND2X1   g04234(.A(new_n4298_), .B(new_n4294_), .Y(new_n4299_));
  INVX1    g04235(.A(new_n4299_), .Y(new_n4300_));
  XOR2X1   g04236(.A(new_n4191_), .B(new_n4152_), .Y(new_n4301_));
  OAI22X1  g04237(.A0(new_n2626_), .A1(new_n1465_), .B0(new_n2419_), .B1(new_n3669_), .Y(new_n4302_));
  AOI21X1  g04238(.A0(new_n2424_), .A1(new_n1536_), .B0(new_n4302_), .Y(new_n4303_));
  OAI21X1  g04239(.A0(new_n3676_), .A1(new_n2665_), .B0(new_n4303_), .Y(new_n4304_));
  XOR2X1   g04240(.A(new_n4304_), .B(\a[26] ), .Y(new_n4305_));
  AND2X1   g04241(.A(new_n4305_), .B(new_n4301_), .Y(new_n4306_));
  INVX1    g04242(.A(new_n4306_), .Y(new_n4307_));
  XOR2X1   g04243(.A(new_n4190_), .B(new_n4160_), .Y(new_n4308_));
  OAI22X1  g04244(.A0(new_n2666_), .A1(new_n1586_), .B0(new_n2626_), .B1(new_n3669_), .Y(new_n4309_));
  AOI21X1  g04245(.A0(new_n2418_), .A1(new_n1536_), .B0(new_n4309_), .Y(new_n4310_));
  OAI21X1  g04246(.A0(new_n3478_), .A1(new_n2665_), .B0(new_n4310_), .Y(new_n4311_));
  XOR2X1   g04247(.A(new_n4311_), .B(\a[26] ), .Y(new_n4312_));
  AND2X1   g04248(.A(new_n4312_), .B(new_n4308_), .Y(new_n4313_));
  INVX1    g04249(.A(new_n4313_), .Y(new_n4314_));
  XOR2X1   g04250(.A(new_n4189_), .B(new_n4169_), .Y(new_n4315_));
  AOI22X1  g04251(.A0(new_n2423_), .A1(new_n1536_), .B0(new_n2418_), .B1(new_n3480_), .Y(new_n4316_));
  OAI21X1  g04252(.A0(new_n2666_), .A1(new_n1621_), .B0(new_n4316_), .Y(new_n4317_));
  AOI21X1  g04253(.A0(new_n3697_), .A1(new_n2301_), .B0(new_n4317_), .Y(new_n4318_));
  XOR2X1   g04254(.A(new_n4318_), .B(\a[26] ), .Y(new_n4319_));
  NOR2X1   g04255(.A(new_n4319_), .B(new_n4315_), .Y(new_n4320_));
  INVX1    g04256(.A(new_n4320_), .Y(new_n4321_));
  AOI22X1  g04257(.A0(new_n2424_), .A1(new_n3721_), .B0(new_n2423_), .B1(new_n3480_), .Y(new_n4322_));
  OAI21X1  g04258(.A0(new_n2419_), .A1(new_n1621_), .B0(new_n4322_), .Y(new_n4323_));
  AOI21X1  g04259(.A0(new_n3720_), .A1(new_n2301_), .B0(new_n4323_), .Y(new_n4324_));
  XOR2X1   g04260(.A(new_n4324_), .B(\a[26] ), .Y(new_n4325_));
  INVX1    g04261(.A(new_n4325_), .Y(new_n4326_));
  XOR2X1   g04262(.A(new_n4187_), .B(new_n4185_), .Y(new_n4327_));
  XOR2X1   g04263(.A(new_n4327_), .B(new_n4325_), .Y(new_n4328_));
  AOI22X1  g04264(.A0(new_n2424_), .A1(new_n1676_), .B0(new_n2418_), .B1(new_n3721_), .Y(new_n4329_));
  OAI21X1  g04265(.A0(new_n2626_), .A1(new_n1621_), .B0(new_n4329_), .Y(new_n4330_));
  AOI21X1  g04266(.A0(new_n3745_), .A1(new_n2301_), .B0(new_n4330_), .Y(new_n4331_));
  XOR2X1   g04267(.A(new_n4331_), .B(\a[26] ), .Y(new_n4332_));
  INVX1    g04268(.A(new_n4332_), .Y(new_n4333_));
  INVX1    g04269(.A(new_n4176_), .Y(new_n4334_));
  NAND3X1  g04270(.A(new_n4334_), .B(new_n4174_), .C(\a[29] ), .Y(new_n4335_));
  XOR2X1   g04271(.A(new_n4180_), .B(new_n74_), .Y(new_n4336_));
  XOR2X1   g04272(.A(new_n4336_), .B(new_n4335_), .Y(new_n4337_));
  XOR2X1   g04273(.A(new_n4337_), .B(new_n4332_), .Y(new_n4338_));
  AOI21X1  g04274(.A0(new_n2184_), .A1(new_n3821_), .B0(new_n74_), .Y(new_n4339_));
  XOR2X1   g04275(.A(new_n4339_), .B(new_n4175_), .Y(new_n4340_));
  OAI22X1  g04276(.A0(new_n2626_), .A1(new_n1655_), .B0(new_n2419_), .B1(new_n1674_), .Y(new_n4341_));
  AOI21X1  g04277(.A0(new_n2424_), .A1(new_n1706_), .B0(new_n4341_), .Y(new_n4342_));
  OAI21X1  g04278(.A0(new_n3773_), .A1(new_n2665_), .B0(new_n4342_), .Y(new_n4343_));
  XOR2X1   g04279(.A(new_n4343_), .B(new_n89_), .Y(new_n4344_));
  NOR2X1   g04280(.A(new_n4344_), .B(new_n4340_), .Y(new_n4345_));
  OAI22X1  g04281(.A0(new_n2626_), .A1(new_n1735_), .B0(new_n2419_), .B1(new_n1784_), .Y(new_n4346_));
  AOI21X1  g04282(.A0(new_n4165_), .A1(new_n2301_), .B0(new_n4346_), .Y(new_n4347_));
  XOR2X1   g04283(.A(new_n4347_), .B(\a[26] ), .Y(new_n4348_));
  AND2X1   g04284(.A(new_n2422_), .B(new_n3821_), .Y(new_n4349_));
  OAI22X1  g04285(.A0(new_n2666_), .A1(new_n1784_), .B0(new_n2419_), .B1(new_n1735_), .Y(new_n4350_));
  AOI21X1  g04286(.A0(new_n2423_), .A1(new_n1706_), .B0(new_n4350_), .Y(new_n4351_));
  OAI21X1  g04287(.A0(new_n4177_), .A1(new_n2665_), .B0(new_n4351_), .Y(new_n4352_));
  NOR4X1   g04288(.A(new_n4352_), .B(new_n4349_), .C(new_n4348_), .D(new_n89_), .Y(new_n4353_));
  NAND2X1  g04289(.A(new_n4353_), .B(new_n4176_), .Y(new_n4354_));
  XOR2X1   g04290(.A(new_n4353_), .B(new_n4334_), .Y(new_n4355_));
  AOI22X1  g04291(.A0(new_n2424_), .A1(new_n3819_), .B0(new_n2423_), .B1(new_n1676_), .Y(new_n4356_));
  OAI21X1  g04292(.A0(new_n2419_), .A1(new_n1708_), .B0(new_n4356_), .Y(new_n4357_));
  AOI21X1  g04293(.A0(new_n3829_), .A1(new_n2301_), .B0(new_n4357_), .Y(new_n4358_));
  XOR2X1   g04294(.A(new_n4358_), .B(\a[26] ), .Y(new_n4359_));
  OAI21X1  g04295(.A0(new_n4359_), .A1(new_n4355_), .B0(new_n4354_), .Y(new_n4360_));
  XOR2X1   g04296(.A(new_n4344_), .B(new_n4340_), .Y(new_n4361_));
  AOI21X1  g04297(.A0(new_n4361_), .A1(new_n4360_), .B0(new_n4345_), .Y(new_n4362_));
  NOR2X1   g04298(.A(new_n4362_), .B(new_n4338_), .Y(new_n4363_));
  AOI21X1  g04299(.A0(new_n4337_), .A1(new_n4333_), .B0(new_n4363_), .Y(new_n4364_));
  NOR2X1   g04300(.A(new_n4364_), .B(new_n4328_), .Y(new_n4365_));
  AOI21X1  g04301(.A0(new_n4327_), .A1(new_n4326_), .B0(new_n4365_), .Y(new_n4366_));
  XOR2X1   g04302(.A(new_n4319_), .B(new_n4315_), .Y(new_n4367_));
  INVX1    g04303(.A(new_n4367_), .Y(new_n4368_));
  OAI21X1  g04304(.A0(new_n4368_), .A1(new_n4366_), .B0(new_n4321_), .Y(new_n4369_));
  INVX1    g04305(.A(new_n4369_), .Y(new_n4370_));
  XOR2X1   g04306(.A(new_n4311_), .B(new_n89_), .Y(new_n4371_));
  XOR2X1   g04307(.A(new_n4371_), .B(new_n4308_), .Y(new_n4372_));
  OAI21X1  g04308(.A0(new_n4372_), .A1(new_n4370_), .B0(new_n4314_), .Y(new_n4373_));
  INVX1    g04309(.A(new_n4373_), .Y(new_n4374_));
  XOR2X1   g04310(.A(new_n4304_), .B(new_n89_), .Y(new_n4375_));
  XOR2X1   g04311(.A(new_n4375_), .B(new_n4301_), .Y(new_n4376_));
  OAI21X1  g04312(.A0(new_n4376_), .A1(new_n4374_), .B0(new_n4307_), .Y(new_n4377_));
  INVX1    g04313(.A(new_n4377_), .Y(new_n4378_));
  XOR2X1   g04314(.A(new_n4297_), .B(new_n89_), .Y(new_n4379_));
  XOR2X1   g04315(.A(new_n4379_), .B(new_n4294_), .Y(new_n4380_));
  OAI21X1  g04316(.A0(new_n4380_), .A1(new_n4378_), .B0(new_n4300_), .Y(new_n4381_));
  INVX1    g04317(.A(new_n4381_), .Y(new_n4382_));
  XOR2X1   g04318(.A(new_n4291_), .B(new_n4286_), .Y(new_n4383_));
  OAI21X1  g04319(.A0(new_n4383_), .A1(new_n4382_), .B0(new_n4293_), .Y(new_n4384_));
  INVX1    g04320(.A(new_n4384_), .Y(new_n4385_));
  XOR2X1   g04321(.A(new_n4283_), .B(new_n4278_), .Y(new_n4386_));
  OAI21X1  g04322(.A0(new_n4386_), .A1(new_n4385_), .B0(new_n4285_), .Y(new_n4387_));
  INVX1    g04323(.A(new_n4387_), .Y(new_n4388_));
  XOR2X1   g04324(.A(new_n4276_), .B(new_n4271_), .Y(new_n4389_));
  OAI21X1  g04325(.A0(new_n4389_), .A1(new_n4388_), .B0(new_n4277_), .Y(new_n4390_));
  XOR2X1   g04326(.A(new_n4207_), .B(new_n4206_), .Y(new_n4391_));
  AND2X1   g04327(.A(new_n4391_), .B(new_n4390_), .Y(new_n4392_));
  AOI22X1  g04328(.A0(new_n2745_), .A1(new_n1126_), .B0(new_n2657_), .B1(new_n2977_), .Y(new_n4393_));
  OAI21X1  g04329(.A0(new_n2743_), .A1(new_n1189_), .B0(new_n4393_), .Y(new_n4394_));
  AOI21X1  g04330(.A0(new_n2976_), .A1(new_n2658_), .B0(new_n4394_), .Y(new_n4395_));
  XOR2X1   g04331(.A(new_n4395_), .B(new_n70_), .Y(new_n4396_));
  XOR2X1   g04332(.A(new_n4391_), .B(new_n4390_), .Y(new_n4397_));
  AOI21X1  g04333(.A0(new_n4397_), .A1(new_n4396_), .B0(new_n4392_), .Y(new_n4398_));
  NOR2X1   g04334(.A(new_n4398_), .B(new_n4270_), .Y(new_n4399_));
  XOR2X1   g04335(.A(new_n4398_), .B(new_n4270_), .Y(new_n4400_));
  AOI22X1  g04336(.A0(new_n3146_), .A1(new_n2602_), .B0(new_n2875_), .B1(new_n2603_), .Y(new_n4401_));
  OAI21X1  g04337(.A0(new_n3144_), .A1(new_n957_), .B0(new_n4401_), .Y(new_n4402_));
  AOI21X1  g04338(.A0(new_n2876_), .A1(new_n2601_), .B0(new_n4402_), .Y(new_n4403_));
  XOR2X1   g04339(.A(new_n4403_), .B(\a[20] ), .Y(new_n4404_));
  INVX1    g04340(.A(new_n4404_), .Y(new_n4405_));
  AOI21X1  g04341(.A0(new_n4405_), .A1(new_n4400_), .B0(new_n4399_), .Y(new_n4406_));
  NOR2X1   g04342(.A(new_n4406_), .B(new_n4269_), .Y(new_n4407_));
  XOR2X1   g04343(.A(new_n4406_), .B(new_n4269_), .Y(new_n4408_));
  AOI22X1  g04344(.A0(new_n3546_), .A1(new_n1886_), .B0(new_n3232_), .B1(new_n2036_), .Y(new_n4409_));
  OAI21X1  g04345(.A0(new_n3389_), .A1(new_n690_), .B0(new_n4409_), .Y(new_n4410_));
  AOI21X1  g04346(.A0(new_n3234_), .A1(new_n2035_), .B0(new_n4410_), .Y(new_n4411_));
  XOR2X1   g04347(.A(new_n4411_), .B(new_n2445_), .Y(new_n4412_));
  AOI21X1  g04348(.A0(new_n4412_), .A1(new_n4408_), .B0(new_n4407_), .Y(new_n4413_));
  NOR2X1   g04349(.A(new_n4413_), .B(new_n4268_), .Y(new_n4414_));
  AOI21X1  g04350(.A0(new_n4267_), .A1(new_n4266_), .B0(new_n4414_), .Y(new_n4415_));
  NOR2X1   g04351(.A(new_n4415_), .B(new_n4261_), .Y(new_n4416_));
  XOR2X1   g04352(.A(new_n4415_), .B(new_n4261_), .Y(new_n4417_));
  AOI22X1  g04353(.A0(new_n3984_), .A1(new_n2252_), .B0(new_n3628_), .B1(new_n2246_), .Y(new_n4418_));
  OAI21X1  g04354(.A0(new_n3907_), .A1(new_n2092_), .B0(new_n4418_), .Y(new_n4419_));
  AOI21X1  g04355(.A0(new_n3624_), .A1(new_n2201_), .B0(new_n4419_), .Y(new_n4420_));
  XOR2X1   g04356(.A(new_n4420_), .B(new_n2529_), .Y(new_n4421_));
  AOI21X1  g04357(.A0(new_n4421_), .A1(new_n4417_), .B0(new_n4416_), .Y(new_n4422_));
  NOR2X1   g04358(.A(new_n4422_), .B(new_n4259_), .Y(new_n4423_));
  INVX1    g04359(.A(new_n4423_), .Y(new_n4424_));
  XOR2X1   g04360(.A(new_n4422_), .B(new_n4259_), .Y(new_n4425_));
  INVX1    g04361(.A(new_n4425_), .Y(new_n4426_));
  OR2X1    g04362(.A(new_n4076_), .B(new_n4073_), .Y(new_n4427_));
  INVX1    g04363(.A(new_n4427_), .Y(new_n4428_));
  AOI22X1  g04364(.A0(new_n4428_), .A1(new_n2421_), .B0(new_n4078_), .B1(new_n2420_), .Y(new_n4429_));
  OAI21X1  g04365(.A0(new_n4246_), .A1(new_n2379_), .B0(new_n4429_), .Y(new_n4430_));
  AOI21X1  g04366(.A0(new_n4080_), .A1(new_n2416_), .B0(new_n4430_), .Y(new_n4431_));
  XOR2X1   g04367(.A(new_n4431_), .B(\a[11] ), .Y(new_n4432_));
  OAI21X1  g04368(.A0(new_n4432_), .A1(new_n4426_), .B0(new_n4424_), .Y(new_n4433_));
  INVX1    g04369(.A(new_n4433_), .Y(new_n4434_));
  OAI22X1  g04370(.A0(new_n4427_), .A1(new_n2648_), .B0(new_n4246_), .B1(new_n2414_), .Y(new_n4435_));
  AOI21X1  g04371(.A0(new_n4078_), .A1(new_n2752_), .B0(new_n4435_), .Y(new_n4436_));
  OAI21X1  g04372(.A0(new_n4245_), .A1(new_n2757_), .B0(new_n4436_), .Y(new_n4437_));
  XOR2X1   g04373(.A(new_n4437_), .B(new_n2911_), .Y(new_n4438_));
  NOR2X1   g04374(.A(new_n4438_), .B(new_n4434_), .Y(new_n4439_));
  INVX1    g04375(.A(new_n4439_), .Y(new_n4440_));
  XOR2X1   g04376(.A(new_n4438_), .B(new_n4434_), .Y(new_n4441_));
  INVX1    g04377(.A(new_n4441_), .Y(new_n4442_));
  XOR2X1   g04378(.A(new_n4242_), .B(new_n4241_), .Y(new_n4443_));
  OAI21X1  g04379(.A0(new_n4443_), .A1(new_n4442_), .B0(new_n4440_), .Y(new_n4444_));
  XOR2X1   g04380(.A(new_n4253_), .B(new_n4252_), .Y(new_n4445_));
  AND2X1   g04381(.A(new_n4445_), .B(new_n4444_), .Y(new_n4446_));
  XOR2X1   g04382(.A(new_n4443_), .B(new_n4441_), .Y(new_n4447_));
  XOR2X1   g04383(.A(new_n4421_), .B(new_n4417_), .Y(new_n4448_));
  INVX1    g04384(.A(new_n4268_), .Y(new_n4449_));
  XOR2X1   g04385(.A(new_n4413_), .B(new_n4449_), .Y(new_n4450_));
  AOI22X1  g04386(.A0(new_n3984_), .A1(new_n2093_), .B0(new_n3628_), .B1(new_n1887_), .Y(new_n4451_));
  OAI21X1  g04387(.A0(new_n3907_), .A1(new_n2183_), .B0(new_n4451_), .Y(new_n4452_));
  AOI21X1  g04388(.A0(new_n3624_), .A1(new_n2430_), .B0(new_n4452_), .Y(new_n4453_));
  XOR2X1   g04389(.A(new_n4453_), .B(\a[14] ), .Y(new_n4454_));
  NOR2X1   g04390(.A(new_n4454_), .B(new_n4450_), .Y(new_n4455_));
  XOR2X1   g04391(.A(new_n4412_), .B(new_n4408_), .Y(new_n4456_));
  INVX1    g04392(.A(new_n4456_), .Y(new_n4457_));
  XOR2X1   g04393(.A(new_n4404_), .B(new_n4400_), .Y(new_n4458_));
  AOI22X1  g04394(.A0(new_n2745_), .A1(new_n1187_), .B0(new_n2696_), .B1(new_n2977_), .Y(new_n4459_));
  OAI21X1  g04395(.A0(new_n4016_), .A1(new_n1294_), .B0(new_n4459_), .Y(new_n4460_));
  AOI21X1  g04396(.A0(new_n3189_), .A1(new_n2658_), .B0(new_n4460_), .Y(new_n4461_));
  XOR2X1   g04397(.A(new_n4461_), .B(\a[23] ), .Y(new_n4462_));
  XOR2X1   g04398(.A(new_n4389_), .B(new_n4387_), .Y(new_n4463_));
  OR2X1    g04399(.A(new_n4463_), .B(new_n4462_), .Y(new_n4464_));
  XOR2X1   g04400(.A(new_n4463_), .B(new_n4462_), .Y(new_n4465_));
  INVX1    g04401(.A(new_n4465_), .Y(new_n4466_));
  AOI22X1  g04402(.A0(new_n2745_), .A1(new_n2977_), .B0(new_n2657_), .B1(new_n3055_), .Y(new_n4467_));
  OAI21X1  g04403(.A0(new_n2743_), .A1(new_n1294_), .B0(new_n4467_), .Y(new_n4468_));
  AOI21X1  g04404(.A0(new_n3054_), .A1(new_n2658_), .B0(new_n4468_), .Y(new_n4469_));
  XOR2X1   g04405(.A(new_n4469_), .B(\a[23] ), .Y(new_n4470_));
  XOR2X1   g04406(.A(new_n4386_), .B(new_n4384_), .Y(new_n4471_));
  NOR2X1   g04407(.A(new_n4471_), .B(new_n4470_), .Y(new_n4472_));
  XOR2X1   g04408(.A(new_n4471_), .B(new_n4470_), .Y(new_n4473_));
  AOI22X1  g04409(.A0(new_n2745_), .A1(new_n3342_), .B0(new_n2657_), .B1(new_n1357_), .Y(new_n4474_));
  OAI21X1  g04410(.A0(new_n2743_), .A1(new_n1339_), .B0(new_n4474_), .Y(new_n4475_));
  AOI21X1  g04411(.A0(new_n3341_), .A1(new_n2658_), .B0(new_n4475_), .Y(new_n4476_));
  XOR2X1   g04412(.A(new_n4476_), .B(\a[23] ), .Y(new_n4477_));
  XOR2X1   g04413(.A(new_n4383_), .B(new_n4381_), .Y(new_n4478_));
  OR2X1    g04414(.A(new_n4478_), .B(new_n4477_), .Y(new_n4479_));
  XOR2X1   g04415(.A(new_n4478_), .B(new_n4477_), .Y(new_n4480_));
  INVX1    g04416(.A(new_n4480_), .Y(new_n4481_));
  AOI22X1  g04417(.A0(new_n2745_), .A1(new_n3055_), .B0(new_n2696_), .B1(new_n1357_), .Y(new_n4482_));
  OAI21X1  g04418(.A0(new_n4016_), .A1(new_n1389_), .B0(new_n4482_), .Y(new_n4483_));
  AOI21X1  g04419(.A0(new_n3425_), .A1(new_n2658_), .B0(new_n4483_), .Y(new_n4484_));
  XOR2X1   g04420(.A(new_n4484_), .B(\a[23] ), .Y(new_n4485_));
  XOR2X1   g04421(.A(new_n4380_), .B(new_n4377_), .Y(new_n4486_));
  NOR2X1   g04422(.A(new_n4486_), .B(new_n4485_), .Y(new_n4487_));
  XOR2X1   g04423(.A(new_n4486_), .B(new_n4485_), .Y(new_n4488_));
  AOI22X1  g04424(.A0(new_n2745_), .A1(new_n1357_), .B0(new_n2657_), .B1(new_n3327_), .Y(new_n4489_));
  OAI21X1  g04425(.A0(new_n2743_), .A1(new_n1389_), .B0(new_n4489_), .Y(new_n4490_));
  AOI21X1  g04426(.A0(new_n3326_), .A1(new_n2658_), .B0(new_n4490_), .Y(new_n4491_));
  XOR2X1   g04427(.A(new_n4491_), .B(\a[23] ), .Y(new_n4492_));
  XOR2X1   g04428(.A(new_n4376_), .B(new_n4373_), .Y(new_n4493_));
  OR2X1    g04429(.A(new_n4493_), .B(new_n4492_), .Y(new_n4494_));
  XOR2X1   g04430(.A(new_n4493_), .B(new_n4492_), .Y(new_n4495_));
  INVX1    g04431(.A(new_n4495_), .Y(new_n4496_));
  AOI22X1  g04432(.A0(new_n2696_), .A1(new_n3327_), .B0(new_n2657_), .B1(new_n1800_), .Y(new_n4497_));
  OAI21X1  g04433(.A0(new_n2753_), .A1(new_n1389_), .B0(new_n4497_), .Y(new_n4498_));
  AOI21X1  g04434(.A0(new_n3497_), .A1(new_n2658_), .B0(new_n4498_), .Y(new_n4499_));
  XOR2X1   g04435(.A(new_n4499_), .B(\a[23] ), .Y(new_n4500_));
  XOR2X1   g04436(.A(new_n4372_), .B(new_n4369_), .Y(new_n4501_));
  NOR2X1   g04437(.A(new_n4501_), .B(new_n4500_), .Y(new_n4502_));
  XOR2X1   g04438(.A(new_n4501_), .B(new_n4500_), .Y(new_n4503_));
  NOR2X1   g04439(.A(new_n3667_), .B(new_n2692_), .Y(new_n4504_));
  AOI22X1  g04440(.A0(new_n2745_), .A1(new_n3327_), .B0(new_n2657_), .B1(new_n1490_), .Y(new_n4505_));
  OAI21X1  g04441(.A0(new_n2743_), .A1(new_n1465_), .B0(new_n4505_), .Y(new_n4506_));
  NOR2X1   g04442(.A(new_n4506_), .B(new_n4504_), .Y(new_n4507_));
  XOR2X1   g04443(.A(new_n4507_), .B(\a[23] ), .Y(new_n4508_));
  XOR2X1   g04444(.A(new_n4367_), .B(new_n4366_), .Y(new_n4509_));
  OR2X1    g04445(.A(new_n4509_), .B(new_n4508_), .Y(new_n4510_));
  XOR2X1   g04446(.A(new_n4509_), .B(new_n4508_), .Y(new_n4511_));
  INVX1    g04447(.A(new_n4511_), .Y(new_n4512_));
  INVX1    g04448(.A(new_n4328_), .Y(new_n4513_));
  XOR2X1   g04449(.A(new_n4364_), .B(new_n4513_), .Y(new_n4514_));
  OAI22X1  g04450(.A0(new_n2753_), .A1(new_n1465_), .B0(new_n2743_), .B1(new_n3669_), .Y(new_n4515_));
  AOI21X1  g04451(.A0(new_n2657_), .A1(new_n1536_), .B0(new_n4515_), .Y(new_n4516_));
  OAI21X1  g04452(.A0(new_n3676_), .A1(new_n2692_), .B0(new_n4516_), .Y(new_n4517_));
  XOR2X1   g04453(.A(new_n4517_), .B(new_n70_), .Y(new_n4518_));
  NOR2X1   g04454(.A(new_n4518_), .B(new_n4514_), .Y(new_n4519_));
  XOR2X1   g04455(.A(new_n4362_), .B(new_n4338_), .Y(new_n4520_));
  INVX1    g04456(.A(new_n4520_), .Y(new_n4521_));
  OAI22X1  g04457(.A0(new_n2753_), .A1(new_n3669_), .B0(new_n4016_), .B1(new_n1586_), .Y(new_n4522_));
  AOI21X1  g04458(.A0(new_n2696_), .A1(new_n1536_), .B0(new_n4522_), .Y(new_n4523_));
  OAI21X1  g04459(.A0(new_n3478_), .A1(new_n2692_), .B0(new_n4523_), .Y(new_n4524_));
  XOR2X1   g04460(.A(new_n4524_), .B(new_n70_), .Y(new_n4525_));
  OR2X1    g04461(.A(new_n4525_), .B(new_n4521_), .Y(new_n4526_));
  AOI22X1  g04462(.A0(new_n2745_), .A1(new_n1536_), .B0(new_n2696_), .B1(new_n3480_), .Y(new_n4527_));
  OAI21X1  g04463(.A0(new_n4016_), .A1(new_n1621_), .B0(new_n4527_), .Y(new_n4528_));
  AOI21X1  g04464(.A0(new_n3697_), .A1(new_n2658_), .B0(new_n4528_), .Y(new_n4529_));
  XOR2X1   g04465(.A(new_n4529_), .B(\a[23] ), .Y(new_n4530_));
  INVX1    g04466(.A(new_n4530_), .Y(new_n4531_));
  XOR2X1   g04467(.A(new_n4361_), .B(new_n4360_), .Y(new_n4532_));
  AND2X1   g04468(.A(new_n4532_), .B(new_n4531_), .Y(new_n4533_));
  INVX1    g04469(.A(new_n4533_), .Y(new_n4534_));
  XOR2X1   g04470(.A(new_n4532_), .B(new_n4530_), .Y(new_n4535_));
  INVX1    g04471(.A(new_n4359_), .Y(new_n4536_));
  XOR2X1   g04472(.A(new_n4536_), .B(new_n4355_), .Y(new_n4537_));
  INVX1    g04473(.A(new_n1621_), .Y(new_n4538_));
  OAI22X1  g04474(.A0(new_n2753_), .A1(new_n1586_), .B0(new_n4016_), .B1(new_n1655_), .Y(new_n4539_));
  AOI21X1  g04475(.A0(new_n2696_), .A1(new_n4538_), .B0(new_n4539_), .Y(new_n4540_));
  OAI21X1  g04476(.A0(new_n3719_), .A1(new_n2692_), .B0(new_n4540_), .Y(new_n4541_));
  XOR2X1   g04477(.A(new_n4541_), .B(new_n70_), .Y(new_n4542_));
  NOR2X1   g04478(.A(new_n4542_), .B(new_n4537_), .Y(new_n4543_));
  AOI22X1  g04479(.A0(new_n2696_), .A1(new_n3721_), .B0(new_n2657_), .B1(new_n1676_), .Y(new_n4544_));
  OAI21X1  g04480(.A0(new_n2753_), .A1(new_n1621_), .B0(new_n4544_), .Y(new_n4545_));
  AOI21X1  g04481(.A0(new_n3745_), .A1(new_n2658_), .B0(new_n4545_), .Y(new_n4546_));
  XOR2X1   g04482(.A(new_n4546_), .B(\a[23] ), .Y(new_n4547_));
  INVX1    g04483(.A(new_n4547_), .Y(new_n4548_));
  INVX1    g04484(.A(new_n4349_), .Y(new_n4549_));
  NAND3X1  g04485(.A(new_n4549_), .B(new_n4347_), .C(\a[26] ), .Y(new_n4550_));
  XOR2X1   g04486(.A(new_n4352_), .B(new_n89_), .Y(new_n4551_));
  XOR2X1   g04487(.A(new_n4551_), .B(new_n4550_), .Y(new_n4552_));
  XOR2X1   g04488(.A(new_n4552_), .B(new_n4547_), .Y(new_n4553_));
  AOI21X1  g04489(.A0(new_n2422_), .A1(new_n3821_), .B0(new_n89_), .Y(new_n4554_));
  XOR2X1   g04490(.A(new_n4554_), .B(new_n4348_), .Y(new_n4555_));
  OAI22X1  g04491(.A0(new_n2753_), .A1(new_n1655_), .B0(new_n2743_), .B1(new_n1674_), .Y(new_n4556_));
  AOI21X1  g04492(.A0(new_n2657_), .A1(new_n1706_), .B0(new_n4556_), .Y(new_n4557_));
  OAI21X1  g04493(.A0(new_n3773_), .A1(new_n2692_), .B0(new_n4557_), .Y(new_n4558_));
  XOR2X1   g04494(.A(new_n4558_), .B(new_n70_), .Y(new_n4559_));
  NOR2X1   g04495(.A(new_n4559_), .B(new_n4555_), .Y(new_n4560_));
  OAI22X1  g04496(.A0(new_n2753_), .A1(new_n1735_), .B0(new_n2743_), .B1(new_n1784_), .Y(new_n4561_));
  AOI21X1  g04497(.A0(new_n4165_), .A1(new_n2658_), .B0(new_n4561_), .Y(new_n4562_));
  XOR2X1   g04498(.A(new_n4562_), .B(\a[23] ), .Y(new_n4563_));
  AND2X1   g04499(.A(new_n2656_), .B(new_n3821_), .Y(new_n4564_));
  OAI22X1  g04500(.A0(new_n2743_), .A1(new_n1735_), .B0(new_n4016_), .B1(new_n1784_), .Y(new_n4565_));
  AOI21X1  g04501(.A0(new_n2745_), .A1(new_n1706_), .B0(new_n4565_), .Y(new_n4566_));
  OAI21X1  g04502(.A0(new_n4177_), .A1(new_n2692_), .B0(new_n4566_), .Y(new_n4567_));
  NOR4X1   g04503(.A(new_n4567_), .B(new_n4564_), .C(new_n4563_), .D(new_n70_), .Y(new_n4568_));
  NAND2X1  g04504(.A(new_n4568_), .B(new_n4349_), .Y(new_n4569_));
  XOR2X1   g04505(.A(new_n4568_), .B(new_n4549_), .Y(new_n4570_));
  AOI22X1  g04506(.A0(new_n2745_), .A1(new_n1676_), .B0(new_n2657_), .B1(new_n3819_), .Y(new_n4571_));
  OAI21X1  g04507(.A0(new_n2743_), .A1(new_n1708_), .B0(new_n4571_), .Y(new_n4572_));
  AOI21X1  g04508(.A0(new_n3829_), .A1(new_n2658_), .B0(new_n4572_), .Y(new_n4573_));
  XOR2X1   g04509(.A(new_n4573_), .B(\a[23] ), .Y(new_n4574_));
  OAI21X1  g04510(.A0(new_n4574_), .A1(new_n4570_), .B0(new_n4569_), .Y(new_n4575_));
  XOR2X1   g04511(.A(new_n4559_), .B(new_n4555_), .Y(new_n4576_));
  AOI21X1  g04512(.A0(new_n4576_), .A1(new_n4575_), .B0(new_n4560_), .Y(new_n4577_));
  NOR2X1   g04513(.A(new_n4577_), .B(new_n4553_), .Y(new_n4578_));
  AOI21X1  g04514(.A0(new_n4552_), .A1(new_n4548_), .B0(new_n4578_), .Y(new_n4579_));
  INVX1    g04515(.A(new_n4579_), .Y(new_n4580_));
  XOR2X1   g04516(.A(new_n4542_), .B(new_n4537_), .Y(new_n4581_));
  AOI21X1  g04517(.A0(new_n4581_), .A1(new_n4580_), .B0(new_n4543_), .Y(new_n4582_));
  OAI21X1  g04518(.A0(new_n4582_), .A1(new_n4535_), .B0(new_n4534_), .Y(new_n4583_));
  INVX1    g04519(.A(new_n4583_), .Y(new_n4584_));
  XOR2X1   g04520(.A(new_n4525_), .B(new_n4520_), .Y(new_n4585_));
  OAI21X1  g04521(.A0(new_n4585_), .A1(new_n4584_), .B0(new_n4526_), .Y(new_n4586_));
  XOR2X1   g04522(.A(new_n4518_), .B(new_n4514_), .Y(new_n4587_));
  AOI21X1  g04523(.A0(new_n4587_), .A1(new_n4586_), .B0(new_n4519_), .Y(new_n4588_));
  OAI21X1  g04524(.A0(new_n4588_), .A1(new_n4512_), .B0(new_n4510_), .Y(new_n4589_));
  AOI21X1  g04525(.A0(new_n4589_), .A1(new_n4503_), .B0(new_n4502_), .Y(new_n4590_));
  OAI21X1  g04526(.A0(new_n4590_), .A1(new_n4496_), .B0(new_n4494_), .Y(new_n4591_));
  AOI21X1  g04527(.A0(new_n4591_), .A1(new_n4488_), .B0(new_n4487_), .Y(new_n4592_));
  OAI21X1  g04528(.A0(new_n4592_), .A1(new_n4481_), .B0(new_n4479_), .Y(new_n4593_));
  AOI21X1  g04529(.A0(new_n4593_), .A1(new_n4473_), .B0(new_n4472_), .Y(new_n4594_));
  OAI21X1  g04530(.A0(new_n4594_), .A1(new_n4466_), .B0(new_n4464_), .Y(new_n4595_));
  XOR2X1   g04531(.A(new_n4397_), .B(new_n4396_), .Y(new_n4596_));
  AND2X1   g04532(.A(new_n4596_), .B(new_n4595_), .Y(new_n4597_));
  AOI22X1  g04533(.A0(new_n3146_), .A1(new_n2835_), .B0(new_n3099_), .B1(new_n2603_), .Y(new_n4598_));
  OAI21X1  g04534(.A0(new_n3250_), .A1(new_n1065_), .B0(new_n4598_), .Y(new_n4599_));
  AOI21X1  g04535(.A0(new_n2876_), .A1(new_n2834_), .B0(new_n4599_), .Y(new_n4600_));
  XOR2X1   g04536(.A(new_n4600_), .B(new_n1920_), .Y(new_n4601_));
  XOR2X1   g04537(.A(new_n4596_), .B(new_n4595_), .Y(new_n4602_));
  AOI21X1  g04538(.A0(new_n4602_), .A1(new_n4601_), .B0(new_n4597_), .Y(new_n4603_));
  NOR2X1   g04539(.A(new_n4603_), .B(new_n4458_), .Y(new_n4604_));
  XOR2X1   g04540(.A(new_n4603_), .B(new_n4458_), .Y(new_n4605_));
  AOI22X1  g04541(.A0(new_n3546_), .A1(new_n2049_), .B0(new_n3232_), .B1(new_n2481_), .Y(new_n4606_));
  OAI21X1  g04542(.A0(new_n3389_), .A1(new_n783_), .B0(new_n4606_), .Y(new_n4607_));
  AOI21X1  g04543(.A0(new_n3234_), .A1(new_n2480_), .B0(new_n4607_), .Y(new_n4608_));
  XOR2X1   g04544(.A(new_n4608_), .B(new_n2445_), .Y(new_n4609_));
  AOI21X1  g04545(.A0(new_n4609_), .A1(new_n4605_), .B0(new_n4604_), .Y(new_n4610_));
  OR2X1    g04546(.A(new_n4610_), .B(new_n4457_), .Y(new_n4611_));
  XOR2X1   g04547(.A(new_n4610_), .B(new_n4457_), .Y(new_n4612_));
  INVX1    g04548(.A(new_n4612_), .Y(new_n4613_));
  AOI22X1  g04549(.A0(new_n3984_), .A1(new_n2246_), .B0(new_n3628_), .B1(new_n2048_), .Y(new_n4614_));
  OAI21X1  g04550(.A0(new_n3907_), .A1(new_n1879_), .B0(new_n4614_), .Y(new_n4615_));
  AOI21X1  g04551(.A0(new_n3624_), .A1(new_n2244_), .B0(new_n4615_), .Y(new_n4616_));
  XOR2X1   g04552(.A(new_n4616_), .B(\a[14] ), .Y(new_n4617_));
  OAI21X1  g04553(.A0(new_n4617_), .A1(new_n4613_), .B0(new_n4611_), .Y(new_n4618_));
  XOR2X1   g04554(.A(new_n4454_), .B(new_n4450_), .Y(new_n4619_));
  AND2X1   g04555(.A(new_n4619_), .B(new_n4618_), .Y(new_n4620_));
  OAI21X1  g04556(.A0(new_n4620_), .A1(new_n4455_), .B0(new_n4448_), .Y(new_n4621_));
  AOI21X1  g04557(.A0(new_n4619_), .A1(new_n4618_), .B0(new_n4455_), .Y(new_n4622_));
  XOR2X1   g04558(.A(new_n4622_), .B(new_n4448_), .Y(new_n4623_));
  AOI22X1  g04559(.A0(new_n4247_), .A1(new_n2420_), .B0(new_n4078_), .B1(new_n2627_), .Y(new_n4624_));
  OAI21X1  g04560(.A0(new_n4427_), .A1(new_n2379_), .B0(new_n4624_), .Y(new_n4625_));
  AOI21X1  g04561(.A0(new_n4080_), .A1(new_n2625_), .B0(new_n4625_), .Y(new_n4626_));
  XOR2X1   g04562(.A(new_n4626_), .B(\a[11] ), .Y(new_n4627_));
  OR2X1    g04563(.A(new_n4627_), .B(new_n4623_), .Y(new_n4628_));
  AND2X1   g04564(.A(new_n4628_), .B(new_n4621_), .Y(new_n4629_));
  XOR2X1   g04565(.A(\a[6] ), .B(new_n3289_), .Y(new_n4630_));
  XOR2X1   g04566(.A(\a[7] ), .B(\a[6] ), .Y(new_n4631_));
  INVX1    g04567(.A(new_n4631_), .Y(new_n4632_));
  XOR2X1   g04568(.A(\a[8] ), .B(\a[7] ), .Y(new_n4633_));
  NAND3X1  g04569(.A(new_n4633_), .B(new_n4632_), .C(new_n4630_), .Y(new_n4634_));
  INVX1    g04570(.A(new_n4634_), .Y(new_n4635_));
  INVX1    g04571(.A(new_n4630_), .Y(new_n4636_));
  AND2X1   g04572(.A(new_n4633_), .B(new_n4636_), .Y(new_n4637_));
  AOI22X1  g04573(.A0(new_n4637_), .A1(new_n2652_), .B0(new_n4635_), .B1(new_n2649_), .Y(new_n4638_));
  XOR2X1   g04574(.A(new_n4638_), .B(\a[8] ), .Y(new_n4639_));
  NOR2X1   g04575(.A(new_n4639_), .B(new_n4629_), .Y(new_n4640_));
  XOR2X1   g04576(.A(new_n4432_), .B(new_n4425_), .Y(new_n4641_));
  INVX1    g04577(.A(new_n4641_), .Y(new_n4642_));
  XOR2X1   g04578(.A(new_n4639_), .B(new_n4629_), .Y(new_n4643_));
  AOI21X1  g04579(.A0(new_n4643_), .A1(new_n4642_), .B0(new_n4640_), .Y(new_n4644_));
  NOR2X1   g04580(.A(new_n4644_), .B(new_n4447_), .Y(new_n4645_));
  INVX1    g04581(.A(new_n4645_), .Y(new_n4646_));
  XOR2X1   g04582(.A(new_n4644_), .B(new_n4447_), .Y(new_n4647_));
  INVX1    g04583(.A(new_n4647_), .Y(new_n4648_));
  XOR2X1   g04584(.A(new_n4643_), .B(new_n4641_), .Y(new_n4649_));
  XOR2X1   g04585(.A(new_n4617_), .B(new_n4612_), .Y(new_n4650_));
  XOR2X1   g04586(.A(new_n4609_), .B(new_n4605_), .Y(new_n4651_));
  INVX1    g04587(.A(new_n4651_), .Y(new_n4652_));
  XOR2X1   g04588(.A(new_n4594_), .B(new_n4466_), .Y(new_n4653_));
  INVX1    g04589(.A(new_n2824_), .Y(new_n4654_));
  OAI22X1  g04590(.A0(new_n3152_), .A1(new_n985_), .B0(new_n3250_), .B1(new_n1127_), .Y(new_n4655_));
  AOI21X1  g04591(.A0(new_n3099_), .A1(new_n1822_), .B0(new_n4655_), .Y(new_n4656_));
  OAI21X1  g04592(.A0(new_n3098_), .A1(new_n4654_), .B0(new_n4656_), .Y(new_n4657_));
  XOR2X1   g04593(.A(new_n4657_), .B(\a[20] ), .Y(new_n4658_));
  NAND2X1  g04594(.A(new_n4658_), .B(new_n4653_), .Y(new_n4659_));
  XOR2X1   g04595(.A(new_n4593_), .B(new_n4473_), .Y(new_n4660_));
  INVX1    g04596(.A(new_n4660_), .Y(new_n4661_));
  OAI22X1  g04597(.A0(new_n3152_), .A1(new_n1065_), .B0(new_n3144_), .B1(new_n1127_), .Y(new_n4662_));
  AOI21X1  g04598(.A0(new_n2875_), .A1(new_n1187_), .B0(new_n4662_), .Y(new_n4663_));
  OAI21X1  g04599(.A0(new_n3352_), .A1(new_n3098_), .B0(new_n4663_), .Y(new_n4664_));
  XOR2X1   g04600(.A(new_n4664_), .B(new_n1920_), .Y(new_n4665_));
  NOR2X1   g04601(.A(new_n4665_), .B(new_n4661_), .Y(new_n4666_));
  INVX1    g04602(.A(new_n4666_), .Y(new_n4667_));
  XOR2X1   g04603(.A(new_n4592_), .B(new_n4481_), .Y(new_n4668_));
  OAI22X1  g04604(.A0(new_n3152_), .A1(new_n1127_), .B0(new_n3250_), .B1(new_n1236_), .Y(new_n4669_));
  AOI21X1  g04605(.A0(new_n3099_), .A1(new_n1187_), .B0(new_n4669_), .Y(new_n4670_));
  OAI21X1  g04606(.A0(new_n3934_), .A1(new_n3098_), .B0(new_n4670_), .Y(new_n4671_));
  XOR2X1   g04607(.A(new_n4671_), .B(\a[20] ), .Y(new_n4672_));
  AND2X1   g04608(.A(new_n4672_), .B(new_n4668_), .Y(new_n4673_));
  INVX1    g04609(.A(new_n4673_), .Y(new_n4674_));
  XOR2X1   g04610(.A(new_n4591_), .B(new_n4488_), .Y(new_n4675_));
  OAI22X1  g04611(.A0(new_n3152_), .A1(new_n1189_), .B0(new_n3144_), .B1(new_n1236_), .Y(new_n4676_));
  AOI21X1  g04612(.A0(new_n2875_), .A1(new_n3342_), .B0(new_n4676_), .Y(new_n4677_));
  OAI21X1  g04613(.A0(new_n3180_), .A1(new_n3098_), .B0(new_n4677_), .Y(new_n4678_));
  XOR2X1   g04614(.A(new_n4678_), .B(\a[20] ), .Y(new_n4679_));
  AND2X1   g04615(.A(new_n4679_), .B(new_n4675_), .Y(new_n4680_));
  INVX1    g04616(.A(new_n4680_), .Y(new_n4681_));
  XOR2X1   g04617(.A(new_n4590_), .B(new_n4496_), .Y(new_n4682_));
  OAI22X1  g04618(.A0(new_n3152_), .A1(new_n1236_), .B0(new_n3250_), .B1(new_n1339_), .Y(new_n4683_));
  AOI21X1  g04619(.A0(new_n3099_), .A1(new_n3342_), .B0(new_n4683_), .Y(new_n4684_));
  OAI21X1  g04620(.A0(new_n3053_), .A1(new_n3098_), .B0(new_n4684_), .Y(new_n4685_));
  XOR2X1   g04621(.A(new_n4685_), .B(\a[20] ), .Y(new_n4686_));
  AND2X1   g04622(.A(new_n4686_), .B(new_n4682_), .Y(new_n4687_));
  INVX1    g04623(.A(new_n4687_), .Y(new_n4688_));
  XOR2X1   g04624(.A(new_n4589_), .B(new_n4503_), .Y(new_n4689_));
  OAI22X1  g04625(.A0(new_n3152_), .A1(new_n1294_), .B0(new_n3250_), .B1(new_n1358_), .Y(new_n4690_));
  AOI21X1  g04626(.A0(new_n3099_), .A1(new_n3055_), .B0(new_n4690_), .Y(new_n4691_));
  OAI21X1  g04627(.A0(new_n3340_), .A1(new_n3098_), .B0(new_n4691_), .Y(new_n4692_));
  XOR2X1   g04628(.A(new_n4692_), .B(\a[20] ), .Y(new_n4693_));
  AND2X1   g04629(.A(new_n4693_), .B(new_n4689_), .Y(new_n4694_));
  INVX1    g04630(.A(new_n4694_), .Y(new_n4695_));
  XOR2X1   g04631(.A(new_n4588_), .B(new_n4512_), .Y(new_n4696_));
  INVX1    g04632(.A(new_n4696_), .Y(new_n4697_));
  OAI22X1  g04633(.A0(new_n3152_), .A1(new_n1339_), .B0(new_n3144_), .B1(new_n1358_), .Y(new_n4698_));
  AOI21X1  g04634(.A0(new_n2875_), .A1(new_n3850_), .B0(new_n4698_), .Y(new_n4699_));
  OAI21X1  g04635(.A0(new_n3941_), .A1(new_n3098_), .B0(new_n4699_), .Y(new_n4700_));
  XOR2X1   g04636(.A(new_n4700_), .B(new_n1920_), .Y(new_n4701_));
  NOR2X1   g04637(.A(new_n4701_), .B(new_n4697_), .Y(new_n4702_));
  INVX1    g04638(.A(new_n4702_), .Y(new_n4703_));
  AOI22X1  g04639(.A0(new_n3146_), .A1(new_n1357_), .B0(new_n2875_), .B1(new_n3327_), .Y(new_n4704_));
  OAI21X1  g04640(.A0(new_n3144_), .A1(new_n1389_), .B0(new_n4704_), .Y(new_n4705_));
  AOI21X1  g04641(.A0(new_n3326_), .A1(new_n2876_), .B0(new_n4705_), .Y(new_n4706_));
  XOR2X1   g04642(.A(new_n4706_), .B(\a[20] ), .Y(new_n4707_));
  INVX1    g04643(.A(new_n4707_), .Y(new_n4708_));
  XOR2X1   g04644(.A(new_n4587_), .B(new_n4586_), .Y(new_n4709_));
  AND2X1   g04645(.A(new_n4709_), .B(new_n4708_), .Y(new_n4710_));
  XOR2X1   g04646(.A(new_n4709_), .B(new_n4707_), .Y(new_n4711_));
  INVX1    g04647(.A(new_n4711_), .Y(new_n4712_));
  AOI22X1  g04648(.A0(new_n3099_), .A1(new_n3327_), .B0(new_n2875_), .B1(new_n1800_), .Y(new_n4713_));
  OAI21X1  g04649(.A0(new_n3152_), .A1(new_n1389_), .B0(new_n4713_), .Y(new_n4714_));
  AOI21X1  g04650(.A0(new_n3497_), .A1(new_n2876_), .B0(new_n4714_), .Y(new_n4715_));
  XOR2X1   g04651(.A(new_n4715_), .B(\a[20] ), .Y(new_n4716_));
  XOR2X1   g04652(.A(new_n4585_), .B(new_n4583_), .Y(new_n4717_));
  OR2X1    g04653(.A(new_n4717_), .B(new_n4716_), .Y(new_n4718_));
  XOR2X1   g04654(.A(new_n4717_), .B(new_n4716_), .Y(new_n4719_));
  INVX1    g04655(.A(new_n4719_), .Y(new_n4720_));
  INVX1    g04656(.A(new_n4535_), .Y(new_n4721_));
  XOR2X1   g04657(.A(new_n4582_), .B(new_n4721_), .Y(new_n4722_));
  OAI22X1  g04658(.A0(new_n3152_), .A1(new_n1423_), .B0(new_n3250_), .B1(new_n3669_), .Y(new_n4723_));
  AOI21X1  g04659(.A0(new_n3099_), .A1(new_n1800_), .B0(new_n4723_), .Y(new_n4724_));
  OAI21X1  g04660(.A0(new_n3667_), .A1(new_n3098_), .B0(new_n4724_), .Y(new_n4725_));
  XOR2X1   g04661(.A(new_n4725_), .B(new_n1920_), .Y(new_n4726_));
  NOR2X1   g04662(.A(new_n4726_), .B(new_n4722_), .Y(new_n4727_));
  XOR2X1   g04663(.A(new_n4581_), .B(new_n4580_), .Y(new_n4728_));
  OAI22X1  g04664(.A0(new_n3152_), .A1(new_n1465_), .B0(new_n3144_), .B1(new_n3669_), .Y(new_n4729_));
  AOI21X1  g04665(.A0(new_n2875_), .A1(new_n1536_), .B0(new_n4729_), .Y(new_n4730_));
  OAI21X1  g04666(.A0(new_n3676_), .A1(new_n3098_), .B0(new_n4730_), .Y(new_n4731_));
  XOR2X1   g04667(.A(new_n4731_), .B(\a[20] ), .Y(new_n4732_));
  NAND2X1  g04668(.A(new_n4732_), .B(new_n4728_), .Y(new_n4733_));
  XOR2X1   g04669(.A(new_n4577_), .B(new_n4553_), .Y(new_n4734_));
  INVX1    g04670(.A(new_n4734_), .Y(new_n4735_));
  OAI22X1  g04671(.A0(new_n3152_), .A1(new_n3669_), .B0(new_n3250_), .B1(new_n1586_), .Y(new_n4736_));
  AOI21X1  g04672(.A0(new_n3099_), .A1(new_n1536_), .B0(new_n4736_), .Y(new_n4737_));
  OAI21X1  g04673(.A0(new_n3478_), .A1(new_n3098_), .B0(new_n4737_), .Y(new_n4738_));
  XOR2X1   g04674(.A(new_n4738_), .B(new_n1920_), .Y(new_n4739_));
  NOR2X1   g04675(.A(new_n4739_), .B(new_n4735_), .Y(new_n4740_));
  INVX1    g04676(.A(new_n4740_), .Y(new_n4741_));
  AOI22X1  g04677(.A0(new_n3146_), .A1(new_n1536_), .B0(new_n3099_), .B1(new_n3480_), .Y(new_n4742_));
  OAI21X1  g04678(.A0(new_n3250_), .A1(new_n1621_), .B0(new_n4742_), .Y(new_n4743_));
  AOI21X1  g04679(.A0(new_n3697_), .A1(new_n2876_), .B0(new_n4743_), .Y(new_n4744_));
  XOR2X1   g04680(.A(new_n4744_), .B(\a[20] ), .Y(new_n4745_));
  INVX1    g04681(.A(new_n4745_), .Y(new_n4746_));
  XOR2X1   g04682(.A(new_n4576_), .B(new_n4575_), .Y(new_n4747_));
  AND2X1   g04683(.A(new_n4747_), .B(new_n4746_), .Y(new_n4748_));
  INVX1    g04684(.A(new_n4748_), .Y(new_n4749_));
  XOR2X1   g04685(.A(new_n4747_), .B(new_n4745_), .Y(new_n4750_));
  INVX1    g04686(.A(new_n4574_), .Y(new_n4751_));
  XOR2X1   g04687(.A(new_n4751_), .B(new_n4570_), .Y(new_n4752_));
  OAI22X1  g04688(.A0(new_n3152_), .A1(new_n1586_), .B0(new_n3250_), .B1(new_n1655_), .Y(new_n4753_));
  AOI21X1  g04689(.A0(new_n3099_), .A1(new_n4538_), .B0(new_n4753_), .Y(new_n4754_));
  OAI21X1  g04690(.A0(new_n3719_), .A1(new_n3098_), .B0(new_n4754_), .Y(new_n4755_));
  XOR2X1   g04691(.A(new_n4755_), .B(new_n1920_), .Y(new_n4756_));
  NOR2X1   g04692(.A(new_n4756_), .B(new_n4752_), .Y(new_n4757_));
  AOI22X1  g04693(.A0(new_n3099_), .A1(new_n3721_), .B0(new_n2875_), .B1(new_n1676_), .Y(new_n4758_));
  OAI21X1  g04694(.A0(new_n3152_), .A1(new_n1621_), .B0(new_n4758_), .Y(new_n4759_));
  AOI21X1  g04695(.A0(new_n3745_), .A1(new_n2876_), .B0(new_n4759_), .Y(new_n4760_));
  XOR2X1   g04696(.A(new_n4760_), .B(\a[20] ), .Y(new_n4761_));
  INVX1    g04697(.A(new_n4761_), .Y(new_n4762_));
  INVX1    g04698(.A(new_n4564_), .Y(new_n4763_));
  NAND3X1  g04699(.A(new_n4763_), .B(new_n4562_), .C(\a[23] ), .Y(new_n4764_));
  XOR2X1   g04700(.A(new_n4567_), .B(new_n70_), .Y(new_n4765_));
  XOR2X1   g04701(.A(new_n4765_), .B(new_n4764_), .Y(new_n4766_));
  XOR2X1   g04702(.A(new_n4766_), .B(new_n4761_), .Y(new_n4767_));
  AOI21X1  g04703(.A0(new_n2656_), .A1(new_n3821_), .B0(new_n70_), .Y(new_n4768_));
  XOR2X1   g04704(.A(new_n4768_), .B(new_n4563_), .Y(new_n4769_));
  OAI22X1  g04705(.A0(new_n3152_), .A1(new_n1655_), .B0(new_n3144_), .B1(new_n1674_), .Y(new_n4770_));
  AOI21X1  g04706(.A0(new_n2875_), .A1(new_n1706_), .B0(new_n4770_), .Y(new_n4771_));
  OAI21X1  g04707(.A0(new_n3773_), .A1(new_n3098_), .B0(new_n4771_), .Y(new_n4772_));
  XOR2X1   g04708(.A(new_n4772_), .B(new_n1920_), .Y(new_n4773_));
  NOR2X1   g04709(.A(new_n4773_), .B(new_n4769_), .Y(new_n4774_));
  OAI22X1  g04710(.A0(new_n3152_), .A1(new_n1735_), .B0(new_n3144_), .B1(new_n1784_), .Y(new_n4775_));
  AOI21X1  g04711(.A0(new_n4165_), .A1(new_n2876_), .B0(new_n4775_), .Y(new_n4776_));
  XOR2X1   g04712(.A(new_n4776_), .B(\a[20] ), .Y(new_n4777_));
  AND2X1   g04713(.A(new_n2870_), .B(new_n3821_), .Y(new_n4778_));
  OAI22X1  g04714(.A0(new_n3144_), .A1(new_n1735_), .B0(new_n3250_), .B1(new_n1784_), .Y(new_n4779_));
  AOI21X1  g04715(.A0(new_n3146_), .A1(new_n1706_), .B0(new_n4779_), .Y(new_n4780_));
  OAI21X1  g04716(.A0(new_n4177_), .A1(new_n3098_), .B0(new_n4780_), .Y(new_n4781_));
  NOR4X1   g04717(.A(new_n4781_), .B(new_n4778_), .C(new_n4777_), .D(new_n1920_), .Y(new_n4782_));
  NAND2X1  g04718(.A(new_n4782_), .B(new_n4564_), .Y(new_n4783_));
  XOR2X1   g04719(.A(new_n4782_), .B(new_n4763_), .Y(new_n4784_));
  AOI22X1  g04720(.A0(new_n3146_), .A1(new_n1676_), .B0(new_n2875_), .B1(new_n3819_), .Y(new_n4785_));
  OAI21X1  g04721(.A0(new_n3144_), .A1(new_n1708_), .B0(new_n4785_), .Y(new_n4786_));
  AOI21X1  g04722(.A0(new_n3829_), .A1(new_n2876_), .B0(new_n4786_), .Y(new_n4787_));
  XOR2X1   g04723(.A(new_n4787_), .B(\a[20] ), .Y(new_n4788_));
  OAI21X1  g04724(.A0(new_n4788_), .A1(new_n4784_), .B0(new_n4783_), .Y(new_n4789_));
  XOR2X1   g04725(.A(new_n4773_), .B(new_n4769_), .Y(new_n4790_));
  AOI21X1  g04726(.A0(new_n4790_), .A1(new_n4789_), .B0(new_n4774_), .Y(new_n4791_));
  NOR2X1   g04727(.A(new_n4791_), .B(new_n4767_), .Y(new_n4792_));
  AOI21X1  g04728(.A0(new_n4766_), .A1(new_n4762_), .B0(new_n4792_), .Y(new_n4793_));
  INVX1    g04729(.A(new_n4793_), .Y(new_n4794_));
  XOR2X1   g04730(.A(new_n4756_), .B(new_n4752_), .Y(new_n4795_));
  AOI21X1  g04731(.A0(new_n4795_), .A1(new_n4794_), .B0(new_n4757_), .Y(new_n4796_));
  OAI21X1  g04732(.A0(new_n4796_), .A1(new_n4750_), .B0(new_n4749_), .Y(new_n4797_));
  INVX1    g04733(.A(new_n4797_), .Y(new_n4798_));
  XOR2X1   g04734(.A(new_n4739_), .B(new_n4734_), .Y(new_n4799_));
  OAI21X1  g04735(.A0(new_n4799_), .A1(new_n4798_), .B0(new_n4741_), .Y(new_n4800_));
  INVX1    g04736(.A(new_n4800_), .Y(new_n4801_));
  XOR2X1   g04737(.A(new_n4731_), .B(new_n1920_), .Y(new_n4802_));
  XOR2X1   g04738(.A(new_n4802_), .B(new_n4728_), .Y(new_n4803_));
  OAI21X1  g04739(.A0(new_n4803_), .A1(new_n4801_), .B0(new_n4733_), .Y(new_n4804_));
  XOR2X1   g04740(.A(new_n4726_), .B(new_n4722_), .Y(new_n4805_));
  AOI21X1  g04741(.A0(new_n4805_), .A1(new_n4804_), .B0(new_n4727_), .Y(new_n4806_));
  OAI21X1  g04742(.A0(new_n4806_), .A1(new_n4720_), .B0(new_n4718_), .Y(new_n4807_));
  AOI21X1  g04743(.A0(new_n4807_), .A1(new_n4712_), .B0(new_n4710_), .Y(new_n4808_));
  XOR2X1   g04744(.A(new_n4701_), .B(new_n4696_), .Y(new_n4809_));
  OAI21X1  g04745(.A0(new_n4809_), .A1(new_n4808_), .B0(new_n4703_), .Y(new_n4810_));
  INVX1    g04746(.A(new_n4810_), .Y(new_n4811_));
  XOR2X1   g04747(.A(new_n4692_), .B(new_n1920_), .Y(new_n4812_));
  XOR2X1   g04748(.A(new_n4812_), .B(new_n4689_), .Y(new_n4813_));
  OAI21X1  g04749(.A0(new_n4813_), .A1(new_n4811_), .B0(new_n4695_), .Y(new_n4814_));
  INVX1    g04750(.A(new_n4814_), .Y(new_n4815_));
  XOR2X1   g04751(.A(new_n4685_), .B(new_n1920_), .Y(new_n4816_));
  XOR2X1   g04752(.A(new_n4816_), .B(new_n4682_), .Y(new_n4817_));
  OAI21X1  g04753(.A0(new_n4817_), .A1(new_n4815_), .B0(new_n4688_), .Y(new_n4818_));
  INVX1    g04754(.A(new_n4818_), .Y(new_n4819_));
  XOR2X1   g04755(.A(new_n4678_), .B(new_n1920_), .Y(new_n4820_));
  XOR2X1   g04756(.A(new_n4820_), .B(new_n4675_), .Y(new_n4821_));
  OAI21X1  g04757(.A0(new_n4821_), .A1(new_n4819_), .B0(new_n4681_), .Y(new_n4822_));
  INVX1    g04758(.A(new_n4822_), .Y(new_n4823_));
  XOR2X1   g04759(.A(new_n4671_), .B(new_n1920_), .Y(new_n4824_));
  XOR2X1   g04760(.A(new_n4824_), .B(new_n4668_), .Y(new_n4825_));
  OAI21X1  g04761(.A0(new_n4825_), .A1(new_n4823_), .B0(new_n4674_), .Y(new_n4826_));
  INVX1    g04762(.A(new_n4826_), .Y(new_n4827_));
  XOR2X1   g04763(.A(new_n4665_), .B(new_n4660_), .Y(new_n4828_));
  OAI21X1  g04764(.A0(new_n4828_), .A1(new_n4827_), .B0(new_n4667_), .Y(new_n4829_));
  INVX1    g04765(.A(new_n4829_), .Y(new_n4830_));
  XOR2X1   g04766(.A(new_n4657_), .B(new_n1920_), .Y(new_n4831_));
  XOR2X1   g04767(.A(new_n4831_), .B(new_n4653_), .Y(new_n4832_));
  OAI21X1  g04768(.A0(new_n4832_), .A1(new_n4830_), .B0(new_n4659_), .Y(new_n4833_));
  XOR2X1   g04769(.A(new_n4602_), .B(new_n4601_), .Y(new_n4834_));
  AND2X1   g04770(.A(new_n4834_), .B(new_n4833_), .Y(new_n4835_));
  AOI22X1  g04771(.A0(new_n3546_), .A1(new_n2036_), .B0(new_n3232_), .B1(new_n2602_), .Y(new_n4836_));
  OAI21X1  g04772(.A0(new_n3389_), .A1(new_n847_), .B0(new_n4836_), .Y(new_n4837_));
  AOI21X1  g04773(.A0(new_n3234_), .A1(new_n2494_), .B0(new_n4837_), .Y(new_n4838_));
  XOR2X1   g04774(.A(new_n4838_), .B(\a[17] ), .Y(new_n4839_));
  INVX1    g04775(.A(new_n4839_), .Y(new_n4840_));
  XOR2X1   g04776(.A(new_n4834_), .B(new_n4833_), .Y(new_n4841_));
  AOI21X1  g04777(.A0(new_n4841_), .A1(new_n4840_), .B0(new_n4835_), .Y(new_n4842_));
  NOR2X1   g04778(.A(new_n4842_), .B(new_n4652_), .Y(new_n4843_));
  XOR2X1   g04779(.A(new_n4842_), .B(new_n4652_), .Y(new_n4844_));
  AOI22X1  g04780(.A0(new_n3984_), .A1(new_n1887_), .B0(new_n3628_), .B1(new_n1886_), .Y(new_n4845_));
  OAI21X1  g04781(.A0(new_n3907_), .A1(new_n520_), .B0(new_n4845_), .Y(new_n4846_));
  AOI21X1  g04782(.A0(new_n3624_), .A1(new_n1882_), .B0(new_n4846_), .Y(new_n4847_));
  XOR2X1   g04783(.A(new_n4847_), .B(new_n2529_), .Y(new_n4848_));
  AOI21X1  g04784(.A0(new_n4848_), .A1(new_n4844_), .B0(new_n4843_), .Y(new_n4849_));
  NOR2X1   g04785(.A(new_n4849_), .B(new_n4650_), .Y(new_n4850_));
  INVX1    g04786(.A(new_n4850_), .Y(new_n4851_));
  XOR2X1   g04787(.A(new_n4849_), .B(new_n4650_), .Y(new_n4852_));
  INVX1    g04788(.A(new_n4852_), .Y(new_n4853_));
  AOI22X1  g04789(.A0(new_n4428_), .A1(new_n2627_), .B0(new_n4078_), .B1(new_n2093_), .Y(new_n4854_));
  OAI21X1  g04790(.A0(new_n4246_), .A1(new_n2137_), .B0(new_n4854_), .Y(new_n4855_));
  AOI21X1  g04791(.A0(new_n4080_), .A1(new_n2294_), .B0(new_n4855_), .Y(new_n4856_));
  XOR2X1   g04792(.A(new_n4856_), .B(\a[11] ), .Y(new_n4857_));
  OAI21X1  g04793(.A0(new_n4857_), .A1(new_n4853_), .B0(new_n4851_), .Y(new_n4858_));
  INVX1    g04794(.A(new_n4858_), .Y(new_n4859_));
  OAI22X1  g04795(.A0(new_n4427_), .A1(new_n2339_), .B0(new_n4077_), .B1(new_n2137_), .Y(new_n4860_));
  AOI21X1  g04796(.A0(new_n4247_), .A1(new_n2627_), .B0(new_n4860_), .Y(new_n4861_));
  OAI21X1  g04797(.A0(new_n4245_), .A1(new_n2670_), .B0(new_n4861_), .Y(new_n4862_));
  XOR2X1   g04798(.A(new_n4862_), .B(new_n2911_), .Y(new_n4863_));
  NOR2X1   g04799(.A(new_n4863_), .B(new_n4859_), .Y(new_n4864_));
  XOR2X1   g04800(.A(new_n4863_), .B(new_n4859_), .Y(new_n4865_));
  XOR2X1   g04801(.A(new_n4619_), .B(new_n4618_), .Y(new_n4866_));
  AOI21X1  g04802(.A0(new_n4866_), .A1(new_n4865_), .B0(new_n4864_), .Y(new_n4867_));
  INVX1    g04803(.A(new_n4637_), .Y(new_n4868_));
  NAND2X1  g04804(.A(new_n4631_), .B(new_n4630_), .Y(new_n4869_));
  INVX1    g04805(.A(new_n4869_), .Y(new_n4870_));
  AOI22X1  g04806(.A0(new_n4870_), .A1(new_n2649_), .B0(new_n4635_), .B1(new_n2421_), .Y(new_n4871_));
  OAI21X1  g04807(.A0(new_n4868_), .A1(new_n2695_), .B0(new_n4871_), .Y(new_n4872_));
  XOR2X1   g04808(.A(new_n4872_), .B(new_n2995_), .Y(new_n4873_));
  NOR2X1   g04809(.A(new_n4873_), .B(new_n4867_), .Y(new_n4874_));
  XOR2X1   g04810(.A(new_n4627_), .B(new_n4623_), .Y(new_n4875_));
  XOR2X1   g04811(.A(new_n4873_), .B(new_n4867_), .Y(new_n4876_));
  AOI21X1  g04812(.A0(new_n4876_), .A1(new_n4875_), .B0(new_n4874_), .Y(new_n4877_));
  NOR2X1   g04813(.A(new_n4877_), .B(new_n4649_), .Y(new_n4878_));
  XOR2X1   g04814(.A(new_n4877_), .B(new_n4649_), .Y(new_n4879_));
  XOR2X1   g04815(.A(new_n4857_), .B(new_n4852_), .Y(new_n4880_));
  XOR2X1   g04816(.A(new_n4848_), .B(new_n4844_), .Y(new_n4881_));
  INVX1    g04817(.A(new_n4881_), .Y(new_n4882_));
  AOI22X1  g04818(.A0(new_n3546_), .A1(new_n2481_), .B0(new_n3232_), .B1(new_n2835_), .Y(new_n4883_));
  OAI21X1  g04819(.A0(new_n3389_), .A1(new_n903_), .B0(new_n4883_), .Y(new_n4884_));
  AOI21X1  g04820(.A0(new_n3234_), .A1(new_n2709_), .B0(new_n4884_), .Y(new_n4885_));
  XOR2X1   g04821(.A(new_n4885_), .B(\a[17] ), .Y(new_n4886_));
  XOR2X1   g04822(.A(new_n4832_), .B(new_n4829_), .Y(new_n4887_));
  OR2X1    g04823(.A(new_n4887_), .B(new_n4886_), .Y(new_n4888_));
  XOR2X1   g04824(.A(new_n4887_), .B(new_n4886_), .Y(new_n4889_));
  INVX1    g04825(.A(new_n4889_), .Y(new_n4890_));
  AOI22X1  g04826(.A0(new_n3546_), .A1(new_n2602_), .B0(new_n3232_), .B1(new_n2603_), .Y(new_n4891_));
  OAI21X1  g04827(.A0(new_n3389_), .A1(new_n957_), .B0(new_n4891_), .Y(new_n4892_));
  AOI21X1  g04828(.A0(new_n3234_), .A1(new_n2601_), .B0(new_n4892_), .Y(new_n4893_));
  XOR2X1   g04829(.A(new_n4893_), .B(\a[17] ), .Y(new_n4894_));
  XOR2X1   g04830(.A(new_n4828_), .B(new_n4826_), .Y(new_n4895_));
  NOR2X1   g04831(.A(new_n4895_), .B(new_n4894_), .Y(new_n4896_));
  XOR2X1   g04832(.A(new_n4895_), .B(new_n4894_), .Y(new_n4897_));
  AOI22X1  g04833(.A0(new_n3546_), .A1(new_n2835_), .B0(new_n3390_), .B1(new_n2603_), .Y(new_n4898_));
  OAI21X1  g04834(.A0(new_n3231_), .A1(new_n1065_), .B0(new_n4898_), .Y(new_n4899_));
  AOI21X1  g04835(.A0(new_n3234_), .A1(new_n2834_), .B0(new_n4899_), .Y(new_n4900_));
  XOR2X1   g04836(.A(new_n4900_), .B(\a[17] ), .Y(new_n4901_));
  XOR2X1   g04837(.A(new_n4825_), .B(new_n4822_), .Y(new_n4902_));
  NOR2X1   g04838(.A(new_n4902_), .B(new_n4901_), .Y(new_n4903_));
  XOR2X1   g04839(.A(new_n4902_), .B(new_n4901_), .Y(new_n4904_));
  AOI22X1  g04840(.A0(new_n3546_), .A1(new_n2603_), .B0(new_n3232_), .B1(new_n1126_), .Y(new_n4905_));
  OAI21X1  g04841(.A0(new_n3389_), .A1(new_n1065_), .B0(new_n4905_), .Y(new_n4906_));
  AOI21X1  g04842(.A0(new_n3234_), .A1(new_n2824_), .B0(new_n4906_), .Y(new_n4907_));
  XOR2X1   g04843(.A(new_n4907_), .B(\a[17] ), .Y(new_n4908_));
  XOR2X1   g04844(.A(new_n4821_), .B(new_n4818_), .Y(new_n4909_));
  NOR2X1   g04845(.A(new_n4909_), .B(new_n4908_), .Y(new_n4910_));
  INVX1    g04846(.A(new_n4910_), .Y(new_n4911_));
  XOR2X1   g04847(.A(new_n4909_), .B(new_n4908_), .Y(new_n4912_));
  INVX1    g04848(.A(new_n4912_), .Y(new_n4913_));
  AOI22X1  g04849(.A0(new_n3546_), .A1(new_n1822_), .B0(new_n3390_), .B1(new_n1126_), .Y(new_n4914_));
  OAI21X1  g04850(.A0(new_n3231_), .A1(new_n1189_), .B0(new_n4914_), .Y(new_n4915_));
  AOI21X1  g04851(.A0(new_n3234_), .A1(new_n2963_), .B0(new_n4915_), .Y(new_n4916_));
  XOR2X1   g04852(.A(new_n4916_), .B(\a[17] ), .Y(new_n4917_));
  XOR2X1   g04853(.A(new_n4817_), .B(new_n4814_), .Y(new_n4918_));
  OR2X1    g04854(.A(new_n4918_), .B(new_n4917_), .Y(new_n4919_));
  XOR2X1   g04855(.A(new_n4918_), .B(new_n4917_), .Y(new_n4920_));
  INVX1    g04856(.A(new_n4920_), .Y(new_n4921_));
  AOI22X1  g04857(.A0(new_n3546_), .A1(new_n1126_), .B0(new_n3232_), .B1(new_n2977_), .Y(new_n4922_));
  OAI21X1  g04858(.A0(new_n3389_), .A1(new_n1189_), .B0(new_n4922_), .Y(new_n4923_));
  AOI21X1  g04859(.A0(new_n3234_), .A1(new_n2976_), .B0(new_n4923_), .Y(new_n4924_));
  XOR2X1   g04860(.A(new_n4924_), .B(\a[17] ), .Y(new_n4925_));
  XOR2X1   g04861(.A(new_n4813_), .B(new_n4810_), .Y(new_n4926_));
  NOR2X1   g04862(.A(new_n4926_), .B(new_n4925_), .Y(new_n4927_));
  XOR2X1   g04863(.A(new_n4926_), .B(new_n4925_), .Y(new_n4928_));
  AOI22X1  g04864(.A0(new_n3546_), .A1(new_n1187_), .B0(new_n3390_), .B1(new_n2977_), .Y(new_n4929_));
  OAI21X1  g04865(.A0(new_n3231_), .A1(new_n1294_), .B0(new_n4929_), .Y(new_n4930_));
  AOI21X1  g04866(.A0(new_n3234_), .A1(new_n3189_), .B0(new_n4930_), .Y(new_n4931_));
  XOR2X1   g04867(.A(new_n4931_), .B(\a[17] ), .Y(new_n4932_));
  INVX1    g04868(.A(new_n4809_), .Y(new_n4933_));
  XOR2X1   g04869(.A(new_n4933_), .B(new_n4808_), .Y(new_n4934_));
  OR2X1    g04870(.A(new_n4934_), .B(new_n4932_), .Y(new_n4935_));
  XOR2X1   g04871(.A(new_n4934_), .B(new_n4932_), .Y(new_n4936_));
  INVX1    g04872(.A(new_n4936_), .Y(new_n4937_));
  XOR2X1   g04873(.A(new_n4807_), .B(new_n4711_), .Y(new_n4938_));
  OAI22X1  g04874(.A0(new_n3545_), .A1(new_n1236_), .B0(new_n3231_), .B1(new_n1339_), .Y(new_n4939_));
  AOI21X1  g04875(.A0(new_n3390_), .A1(new_n3342_), .B0(new_n4939_), .Y(new_n4940_));
  OAI21X1  g04876(.A0(new_n3388_), .A1(new_n3053_), .B0(new_n4940_), .Y(new_n4941_));
  XOR2X1   g04877(.A(new_n4941_), .B(new_n2445_), .Y(new_n4942_));
  NOR2X1   g04878(.A(new_n4942_), .B(new_n4938_), .Y(new_n4943_));
  XOR2X1   g04879(.A(new_n4806_), .B(new_n4720_), .Y(new_n4944_));
  OAI22X1  g04880(.A0(new_n3545_), .A1(new_n1294_), .B0(new_n3231_), .B1(new_n1358_), .Y(new_n4945_));
  AOI21X1  g04881(.A0(new_n3390_), .A1(new_n3055_), .B0(new_n4945_), .Y(new_n4946_));
  OAI21X1  g04882(.A0(new_n3340_), .A1(new_n3388_), .B0(new_n4946_), .Y(new_n4947_));
  XOR2X1   g04883(.A(new_n4947_), .B(\a[17] ), .Y(new_n4948_));
  NAND2X1  g04884(.A(new_n4948_), .B(new_n4944_), .Y(new_n4949_));
  AOI22X1  g04885(.A0(new_n3546_), .A1(new_n3055_), .B0(new_n3390_), .B1(new_n1357_), .Y(new_n4950_));
  OAI21X1  g04886(.A0(new_n3231_), .A1(new_n1389_), .B0(new_n4950_), .Y(new_n4951_));
  AOI21X1  g04887(.A0(new_n3425_), .A1(new_n3234_), .B0(new_n4951_), .Y(new_n4952_));
  XOR2X1   g04888(.A(new_n4952_), .B(\a[17] ), .Y(new_n4953_));
  INVX1    g04889(.A(new_n4953_), .Y(new_n4954_));
  XOR2X1   g04890(.A(new_n4805_), .B(new_n4804_), .Y(new_n4955_));
  AND2X1   g04891(.A(new_n4955_), .B(new_n4954_), .Y(new_n4956_));
  XOR2X1   g04892(.A(new_n4955_), .B(new_n4953_), .Y(new_n4957_));
  AOI22X1  g04893(.A0(new_n3546_), .A1(new_n1357_), .B0(new_n3232_), .B1(new_n3327_), .Y(new_n4958_));
  OAI21X1  g04894(.A0(new_n3389_), .A1(new_n1389_), .B0(new_n4958_), .Y(new_n4959_));
  AOI21X1  g04895(.A0(new_n3326_), .A1(new_n3234_), .B0(new_n4959_), .Y(new_n4960_));
  XOR2X1   g04896(.A(new_n4960_), .B(\a[17] ), .Y(new_n4961_));
  XOR2X1   g04897(.A(new_n4803_), .B(new_n4800_), .Y(new_n4962_));
  NOR2X1   g04898(.A(new_n4962_), .B(new_n4961_), .Y(new_n4963_));
  XOR2X1   g04899(.A(new_n4962_), .B(new_n4961_), .Y(new_n4964_));
  AOI22X1  g04900(.A0(new_n3390_), .A1(new_n3327_), .B0(new_n3232_), .B1(new_n1800_), .Y(new_n4965_));
  OAI21X1  g04901(.A0(new_n3545_), .A1(new_n1389_), .B0(new_n4965_), .Y(new_n4966_));
  AOI21X1  g04902(.A0(new_n3497_), .A1(new_n3234_), .B0(new_n4966_), .Y(new_n4967_));
  XOR2X1   g04903(.A(new_n4967_), .B(\a[17] ), .Y(new_n4968_));
  XOR2X1   g04904(.A(new_n4799_), .B(new_n4797_), .Y(new_n4969_));
  OR2X1    g04905(.A(new_n4969_), .B(new_n4968_), .Y(new_n4970_));
  XOR2X1   g04906(.A(new_n4969_), .B(new_n4968_), .Y(new_n4971_));
  INVX1    g04907(.A(new_n4971_), .Y(new_n4972_));
  INVX1    g04908(.A(new_n4750_), .Y(new_n4973_));
  XOR2X1   g04909(.A(new_n4796_), .B(new_n4973_), .Y(new_n4974_));
  OAI22X1  g04910(.A0(new_n3545_), .A1(new_n1423_), .B0(new_n3231_), .B1(new_n3669_), .Y(new_n4975_));
  AOI21X1  g04911(.A0(new_n3390_), .A1(new_n1800_), .B0(new_n4975_), .Y(new_n4976_));
  OAI21X1  g04912(.A0(new_n3667_), .A1(new_n3388_), .B0(new_n4976_), .Y(new_n4977_));
  XOR2X1   g04913(.A(new_n4977_), .B(new_n2445_), .Y(new_n4978_));
  NOR2X1   g04914(.A(new_n4978_), .B(new_n4974_), .Y(new_n4979_));
  XOR2X1   g04915(.A(new_n4795_), .B(new_n4794_), .Y(new_n4980_));
  OAI22X1  g04916(.A0(new_n3545_), .A1(new_n1465_), .B0(new_n3389_), .B1(new_n3669_), .Y(new_n4981_));
  AOI21X1  g04917(.A0(new_n3232_), .A1(new_n1536_), .B0(new_n4981_), .Y(new_n4982_));
  OAI21X1  g04918(.A0(new_n3676_), .A1(new_n3388_), .B0(new_n4982_), .Y(new_n4983_));
  XOR2X1   g04919(.A(new_n4983_), .B(\a[17] ), .Y(new_n4984_));
  NAND2X1  g04920(.A(new_n4984_), .B(new_n4980_), .Y(new_n4985_));
  XOR2X1   g04921(.A(new_n4791_), .B(new_n4767_), .Y(new_n4986_));
  INVX1    g04922(.A(new_n4986_), .Y(new_n4987_));
  OAI22X1  g04923(.A0(new_n3545_), .A1(new_n3669_), .B0(new_n3231_), .B1(new_n1586_), .Y(new_n4988_));
  AOI21X1  g04924(.A0(new_n3390_), .A1(new_n1536_), .B0(new_n4988_), .Y(new_n4989_));
  OAI21X1  g04925(.A0(new_n3478_), .A1(new_n3388_), .B0(new_n4989_), .Y(new_n4990_));
  XOR2X1   g04926(.A(new_n4990_), .B(new_n2445_), .Y(new_n4991_));
  NOR2X1   g04927(.A(new_n4991_), .B(new_n4987_), .Y(new_n4992_));
  AOI22X1  g04928(.A0(new_n3546_), .A1(new_n1536_), .B0(new_n3390_), .B1(new_n3480_), .Y(new_n4993_));
  OAI21X1  g04929(.A0(new_n3231_), .A1(new_n1621_), .B0(new_n4993_), .Y(new_n4994_));
  AOI21X1  g04930(.A0(new_n3697_), .A1(new_n3234_), .B0(new_n4994_), .Y(new_n4995_));
  XOR2X1   g04931(.A(new_n4995_), .B(\a[17] ), .Y(new_n4996_));
  INVX1    g04932(.A(new_n4996_), .Y(new_n4997_));
  XOR2X1   g04933(.A(new_n4790_), .B(new_n4789_), .Y(new_n4998_));
  AND2X1   g04934(.A(new_n4998_), .B(new_n4997_), .Y(new_n4999_));
  INVX1    g04935(.A(new_n4999_), .Y(new_n5000_));
  XOR2X1   g04936(.A(new_n4998_), .B(new_n4996_), .Y(new_n5001_));
  INVX1    g04937(.A(new_n4788_), .Y(new_n5002_));
  XOR2X1   g04938(.A(new_n5002_), .B(new_n4784_), .Y(new_n5003_));
  OAI22X1  g04939(.A0(new_n3545_), .A1(new_n1586_), .B0(new_n3231_), .B1(new_n1655_), .Y(new_n5004_));
  AOI21X1  g04940(.A0(new_n3390_), .A1(new_n4538_), .B0(new_n5004_), .Y(new_n5005_));
  OAI21X1  g04941(.A0(new_n3719_), .A1(new_n3388_), .B0(new_n5005_), .Y(new_n5006_));
  XOR2X1   g04942(.A(new_n5006_), .B(new_n2445_), .Y(new_n5007_));
  NOR2X1   g04943(.A(new_n5007_), .B(new_n5003_), .Y(new_n5008_));
  AOI22X1  g04944(.A0(new_n3390_), .A1(new_n3721_), .B0(new_n3232_), .B1(new_n1676_), .Y(new_n5009_));
  OAI21X1  g04945(.A0(new_n3545_), .A1(new_n1621_), .B0(new_n5009_), .Y(new_n5010_));
  AOI21X1  g04946(.A0(new_n3745_), .A1(new_n3234_), .B0(new_n5010_), .Y(new_n5011_));
  XOR2X1   g04947(.A(new_n5011_), .B(\a[17] ), .Y(new_n5012_));
  INVX1    g04948(.A(new_n4778_), .Y(new_n5013_));
  NAND3X1  g04949(.A(new_n5013_), .B(new_n4776_), .C(\a[20] ), .Y(new_n5014_));
  XOR2X1   g04950(.A(new_n4781_), .B(new_n1920_), .Y(new_n5015_));
  AND2X1   g04951(.A(new_n5015_), .B(new_n5014_), .Y(new_n5016_));
  NOR3X1   g04952(.A(new_n5016_), .B(new_n5012_), .C(new_n4782_), .Y(new_n5017_));
  XOR2X1   g04953(.A(new_n5015_), .B(new_n5014_), .Y(new_n5018_));
  XOR2X1   g04954(.A(new_n5018_), .B(new_n5012_), .Y(new_n5019_));
  AOI21X1  g04955(.A0(new_n2870_), .A1(new_n3821_), .B0(new_n1920_), .Y(new_n5020_));
  XOR2X1   g04956(.A(new_n5020_), .B(new_n4777_), .Y(new_n5021_));
  OAI22X1  g04957(.A0(new_n3545_), .A1(new_n1655_), .B0(new_n3389_), .B1(new_n1674_), .Y(new_n5022_));
  AOI21X1  g04958(.A0(new_n3232_), .A1(new_n1706_), .B0(new_n5022_), .Y(new_n5023_));
  OAI21X1  g04959(.A0(new_n3773_), .A1(new_n3388_), .B0(new_n5023_), .Y(new_n5024_));
  XOR2X1   g04960(.A(new_n5024_), .B(new_n2445_), .Y(new_n5025_));
  NOR2X1   g04961(.A(new_n5025_), .B(new_n5021_), .Y(new_n5026_));
  OAI22X1  g04962(.A0(new_n3545_), .A1(new_n1735_), .B0(new_n3389_), .B1(new_n1784_), .Y(new_n5027_));
  AOI21X1  g04963(.A0(new_n4165_), .A1(new_n3234_), .B0(new_n5027_), .Y(new_n5028_));
  XOR2X1   g04964(.A(new_n5028_), .B(\a[17] ), .Y(new_n5029_));
  INVX1    g04965(.A(new_n3230_), .Y(new_n5030_));
  AND2X1   g04966(.A(new_n5030_), .B(new_n3821_), .Y(new_n5031_));
  OAI22X1  g04967(.A0(new_n3389_), .A1(new_n1735_), .B0(new_n3231_), .B1(new_n1784_), .Y(new_n5032_));
  AOI21X1  g04968(.A0(new_n3546_), .A1(new_n1706_), .B0(new_n5032_), .Y(new_n5033_));
  OAI21X1  g04969(.A0(new_n4177_), .A1(new_n3388_), .B0(new_n5033_), .Y(new_n5034_));
  NOR4X1   g04970(.A(new_n5034_), .B(new_n5031_), .C(new_n5029_), .D(new_n2445_), .Y(new_n5035_));
  NAND2X1  g04971(.A(new_n5035_), .B(new_n4778_), .Y(new_n5036_));
  XOR2X1   g04972(.A(new_n5035_), .B(new_n5013_), .Y(new_n5037_));
  AOI22X1  g04973(.A0(new_n3546_), .A1(new_n1676_), .B0(new_n3232_), .B1(new_n3819_), .Y(new_n5038_));
  OAI21X1  g04974(.A0(new_n3389_), .A1(new_n1708_), .B0(new_n5038_), .Y(new_n5039_));
  AOI21X1  g04975(.A0(new_n3829_), .A1(new_n3234_), .B0(new_n5039_), .Y(new_n5040_));
  XOR2X1   g04976(.A(new_n5040_), .B(\a[17] ), .Y(new_n5041_));
  OAI21X1  g04977(.A0(new_n5041_), .A1(new_n5037_), .B0(new_n5036_), .Y(new_n5042_));
  XOR2X1   g04978(.A(new_n5025_), .B(new_n5021_), .Y(new_n5043_));
  AOI21X1  g04979(.A0(new_n5043_), .A1(new_n5042_), .B0(new_n5026_), .Y(new_n5044_));
  NOR2X1   g04980(.A(new_n5044_), .B(new_n5019_), .Y(new_n5045_));
  OR2X1    g04981(.A(new_n5045_), .B(new_n5017_), .Y(new_n5046_));
  XOR2X1   g04982(.A(new_n5007_), .B(new_n5003_), .Y(new_n5047_));
  AOI21X1  g04983(.A0(new_n5047_), .A1(new_n5046_), .B0(new_n5008_), .Y(new_n5048_));
  OR2X1    g04984(.A(new_n5048_), .B(new_n5001_), .Y(new_n5049_));
  XOR2X1   g04985(.A(new_n4991_), .B(new_n4986_), .Y(new_n5050_));
  AOI21X1  g04986(.A0(new_n5049_), .A1(new_n5000_), .B0(new_n5050_), .Y(new_n5051_));
  NOR2X1   g04987(.A(new_n5051_), .B(new_n4992_), .Y(new_n5052_));
  XOR2X1   g04988(.A(new_n4983_), .B(new_n2445_), .Y(new_n5053_));
  XOR2X1   g04989(.A(new_n5053_), .B(new_n4980_), .Y(new_n5054_));
  OAI21X1  g04990(.A0(new_n5054_), .A1(new_n5052_), .B0(new_n4985_), .Y(new_n5055_));
  XOR2X1   g04991(.A(new_n4978_), .B(new_n4974_), .Y(new_n5056_));
  AOI21X1  g04992(.A0(new_n5056_), .A1(new_n5055_), .B0(new_n4979_), .Y(new_n5057_));
  OAI21X1  g04993(.A0(new_n5057_), .A1(new_n4972_), .B0(new_n4970_), .Y(new_n5058_));
  AOI21X1  g04994(.A0(new_n5058_), .A1(new_n4964_), .B0(new_n4963_), .Y(new_n5059_));
  NOR2X1   g04995(.A(new_n5059_), .B(new_n4957_), .Y(new_n5060_));
  NOR2X1   g04996(.A(new_n5060_), .B(new_n4956_), .Y(new_n5061_));
  XOR2X1   g04997(.A(new_n4947_), .B(new_n2445_), .Y(new_n5062_));
  XOR2X1   g04998(.A(new_n5062_), .B(new_n4944_), .Y(new_n5063_));
  OAI21X1  g04999(.A0(new_n5063_), .A1(new_n5061_), .B0(new_n4949_), .Y(new_n5064_));
  XOR2X1   g05000(.A(new_n4942_), .B(new_n4938_), .Y(new_n5065_));
  AOI21X1  g05001(.A0(new_n5065_), .A1(new_n5064_), .B0(new_n4943_), .Y(new_n5066_));
  OAI21X1  g05002(.A0(new_n5066_), .A1(new_n4937_), .B0(new_n4935_), .Y(new_n5067_));
  AOI21X1  g05003(.A0(new_n5067_), .A1(new_n4928_), .B0(new_n4927_), .Y(new_n5068_));
  OR2X1    g05004(.A(new_n5068_), .B(new_n4921_), .Y(new_n5069_));
  AND2X1   g05005(.A(new_n5069_), .B(new_n4919_), .Y(new_n5070_));
  OAI21X1  g05006(.A0(new_n5070_), .A1(new_n4913_), .B0(new_n4911_), .Y(new_n5071_));
  AOI21X1  g05007(.A0(new_n5071_), .A1(new_n4904_), .B0(new_n4903_), .Y(new_n5072_));
  INVX1    g05008(.A(new_n5072_), .Y(new_n5073_));
  AOI21X1  g05009(.A0(new_n5073_), .A1(new_n4897_), .B0(new_n4896_), .Y(new_n5074_));
  OAI21X1  g05010(.A0(new_n5074_), .A1(new_n4890_), .B0(new_n4888_), .Y(new_n5075_));
  XOR2X1   g05011(.A(new_n4841_), .B(new_n4840_), .Y(new_n5076_));
  AND2X1   g05012(.A(new_n5076_), .B(new_n5075_), .Y(new_n5077_));
  AOI22X1  g05013(.A0(new_n3984_), .A1(new_n2048_), .B0(new_n3628_), .B1(new_n2049_), .Y(new_n5078_));
  OAI21X1  g05014(.A0(new_n3907_), .A1(new_n623_), .B0(new_n5078_), .Y(new_n5079_));
  AOI21X1  g05015(.A0(new_n3624_), .A1(new_n2047_), .B0(new_n5079_), .Y(new_n5080_));
  XOR2X1   g05016(.A(new_n5080_), .B(\a[14] ), .Y(new_n5081_));
  INVX1    g05017(.A(new_n5081_), .Y(new_n5082_));
  XOR2X1   g05018(.A(new_n5076_), .B(new_n5075_), .Y(new_n5083_));
  AOI21X1  g05019(.A0(new_n5083_), .A1(new_n5082_), .B0(new_n5077_), .Y(new_n5084_));
  NOR2X1   g05020(.A(new_n5084_), .B(new_n4882_), .Y(new_n5085_));
  XOR2X1   g05021(.A(new_n5084_), .B(new_n4882_), .Y(new_n5086_));
  AOI22X1  g05022(.A0(new_n4428_), .A1(new_n2252_), .B0(new_n4078_), .B1(new_n2246_), .Y(new_n5087_));
  OAI21X1  g05023(.A0(new_n4246_), .A1(new_n2092_), .B0(new_n5087_), .Y(new_n5088_));
  AOI21X1  g05024(.A0(new_n4080_), .A1(new_n2201_), .B0(new_n5088_), .Y(new_n5089_));
  XOR2X1   g05025(.A(new_n5089_), .B(new_n2911_), .Y(new_n5090_));
  AOI21X1  g05026(.A0(new_n5090_), .A1(new_n5086_), .B0(new_n5085_), .Y(new_n5091_));
  NOR2X1   g05027(.A(new_n5091_), .B(new_n4880_), .Y(new_n5092_));
  INVX1    g05028(.A(new_n5092_), .Y(new_n5093_));
  XOR2X1   g05029(.A(new_n5091_), .B(new_n4880_), .Y(new_n5094_));
  INVX1    g05030(.A(new_n5094_), .Y(new_n5095_));
  OR2X1    g05031(.A(new_n4633_), .B(new_n4630_), .Y(new_n5096_));
  INVX1    g05032(.A(new_n5096_), .Y(new_n5097_));
  AOI22X1  g05033(.A0(new_n5097_), .A1(new_n2421_), .B0(new_n4635_), .B1(new_n2420_), .Y(new_n5098_));
  OAI21X1  g05034(.A0(new_n4869_), .A1(new_n2379_), .B0(new_n5098_), .Y(new_n5099_));
  AOI21X1  g05035(.A0(new_n4637_), .A1(new_n2416_), .B0(new_n5099_), .Y(new_n5100_));
  XOR2X1   g05036(.A(new_n5100_), .B(\a[8] ), .Y(new_n5101_));
  OAI21X1  g05037(.A0(new_n5101_), .A1(new_n5095_), .B0(new_n5093_), .Y(new_n5102_));
  OAI22X1  g05038(.A0(new_n5096_), .A1(new_n2648_), .B0(new_n4869_), .B1(new_n2414_), .Y(new_n5103_));
  AOI21X1  g05039(.A0(new_n4635_), .A1(new_n2752_), .B0(new_n5103_), .Y(new_n5104_));
  OAI21X1  g05040(.A0(new_n4868_), .A1(new_n2757_), .B0(new_n5104_), .Y(new_n5105_));
  XOR2X1   g05041(.A(new_n5105_), .B(\a[8] ), .Y(new_n5106_));
  AND2X1   g05042(.A(new_n5106_), .B(new_n5102_), .Y(new_n5107_));
  XOR2X1   g05043(.A(new_n5105_), .B(new_n2995_), .Y(new_n5108_));
  XOR2X1   g05044(.A(new_n5108_), .B(new_n5102_), .Y(new_n5109_));
  INVX1    g05045(.A(new_n5109_), .Y(new_n5110_));
  XOR2X1   g05046(.A(new_n4866_), .B(new_n4865_), .Y(new_n5111_));
  AOI21X1  g05047(.A0(new_n5111_), .A1(new_n5110_), .B0(new_n5107_), .Y(new_n5112_));
  INVX1    g05048(.A(new_n5112_), .Y(new_n5113_));
  XOR2X1   g05049(.A(new_n4876_), .B(new_n4875_), .Y(new_n5114_));
  AND2X1   g05050(.A(new_n5114_), .B(new_n5113_), .Y(new_n5115_));
  INVX1    g05051(.A(new_n5115_), .Y(new_n5116_));
  XOR2X1   g05052(.A(new_n5090_), .B(new_n5086_), .Y(new_n5117_));
  INVX1    g05053(.A(new_n5117_), .Y(new_n5118_));
  XOR2X1   g05054(.A(new_n5074_), .B(new_n4890_), .Y(new_n5119_));
  INVX1    g05055(.A(new_n2035_), .Y(new_n5120_));
  OAI22X1  g05056(.A0(new_n3983_), .A1(new_n623_), .B0(new_n3627_), .B1(new_n783_), .Y(new_n5121_));
  AOI21X1  g05057(.A0(new_n3908_), .A1(new_n2049_), .B0(new_n5121_), .Y(new_n5122_));
  OAI21X1  g05058(.A0(new_n3906_), .A1(new_n5120_), .B0(new_n5122_), .Y(new_n5123_));
  XOR2X1   g05059(.A(new_n5123_), .B(\a[14] ), .Y(new_n5124_));
  AND2X1   g05060(.A(new_n5124_), .B(new_n5119_), .Y(new_n5125_));
  XOR2X1   g05061(.A(new_n5073_), .B(new_n4897_), .Y(new_n5126_));
  INVX1    g05062(.A(new_n5126_), .Y(new_n5127_));
  OAI22X1  g05063(.A0(new_n3983_), .A1(new_n690_), .B0(new_n3627_), .B1(new_n847_), .Y(new_n5128_));
  AOI21X1  g05064(.A0(new_n3908_), .A1(new_n2036_), .B0(new_n5128_), .Y(new_n5129_));
  OAI21X1  g05065(.A0(new_n3906_), .A1(new_n2845_), .B0(new_n5129_), .Y(new_n5130_));
  XOR2X1   g05066(.A(new_n5130_), .B(new_n2529_), .Y(new_n5131_));
  NOR2X1   g05067(.A(new_n5131_), .B(new_n5127_), .Y(new_n5132_));
  INVX1    g05068(.A(new_n5132_), .Y(new_n5133_));
  XOR2X1   g05069(.A(new_n5071_), .B(new_n4904_), .Y(new_n5134_));
  OAI22X1  g05070(.A0(new_n3983_), .A1(new_n783_), .B0(new_n3627_), .B1(new_n903_), .Y(new_n5135_));
  AOI21X1  g05071(.A0(new_n3908_), .A1(new_n2481_), .B0(new_n5135_), .Y(new_n5136_));
  OAI21X1  g05072(.A0(new_n3906_), .A1(new_n3261_), .B0(new_n5136_), .Y(new_n5137_));
  XOR2X1   g05073(.A(new_n5137_), .B(\a[14] ), .Y(new_n5138_));
  XOR2X1   g05074(.A(new_n5070_), .B(new_n4913_), .Y(new_n5139_));
  OAI22X1  g05075(.A0(new_n3983_), .A1(new_n847_), .B0(new_n3627_), .B1(new_n957_), .Y(new_n5140_));
  AOI21X1  g05076(.A0(new_n3908_), .A1(new_n2602_), .B0(new_n5140_), .Y(new_n5141_));
  OAI21X1  g05077(.A0(new_n3906_), .A1(new_n2708_), .B0(new_n5141_), .Y(new_n5142_));
  XOR2X1   g05078(.A(new_n5142_), .B(\a[14] ), .Y(new_n5143_));
  AND2X1   g05079(.A(new_n5143_), .B(new_n5139_), .Y(new_n5144_));
  INVX1    g05080(.A(new_n5144_), .Y(new_n5145_));
  XOR2X1   g05081(.A(new_n5068_), .B(new_n4921_), .Y(new_n5146_));
  OAI22X1  g05082(.A0(new_n3983_), .A1(new_n903_), .B0(new_n3627_), .B1(new_n985_), .Y(new_n5147_));
  AOI21X1  g05083(.A0(new_n3908_), .A1(new_n2835_), .B0(new_n5147_), .Y(new_n5148_));
  OAI21X1  g05084(.A0(new_n3906_), .A1(new_n2600_), .B0(new_n5148_), .Y(new_n5149_));
  XOR2X1   g05085(.A(new_n5149_), .B(\a[14] ), .Y(new_n5150_));
  AND2X1   g05086(.A(new_n5150_), .B(new_n5146_), .Y(new_n5151_));
  XOR2X1   g05087(.A(new_n5067_), .B(new_n4928_), .Y(new_n5152_));
  OAI22X1  g05088(.A0(new_n3983_), .A1(new_n957_), .B0(new_n3907_), .B1(new_n985_), .Y(new_n5153_));
  AOI21X1  g05089(.A0(new_n3628_), .A1(new_n1822_), .B0(new_n5153_), .Y(new_n5154_));
  OAI21X1  g05090(.A0(new_n3906_), .A1(new_n2833_), .B0(new_n5154_), .Y(new_n5155_));
  XOR2X1   g05091(.A(new_n5155_), .B(\a[14] ), .Y(new_n5156_));
  XOR2X1   g05092(.A(new_n5066_), .B(new_n4937_), .Y(new_n5157_));
  INVX1    g05093(.A(new_n5157_), .Y(new_n5158_));
  OAI22X1  g05094(.A0(new_n3983_), .A1(new_n985_), .B0(new_n3627_), .B1(new_n1127_), .Y(new_n5159_));
  AOI21X1  g05095(.A0(new_n3908_), .A1(new_n1822_), .B0(new_n5159_), .Y(new_n5160_));
  OAI21X1  g05096(.A0(new_n3906_), .A1(new_n4654_), .B0(new_n5160_), .Y(new_n5161_));
  XOR2X1   g05097(.A(new_n5161_), .B(new_n2529_), .Y(new_n5162_));
  NOR2X1   g05098(.A(new_n5162_), .B(new_n5158_), .Y(new_n5163_));
  INVX1    g05099(.A(new_n5163_), .Y(new_n5164_));
  AOI22X1  g05100(.A0(new_n3984_), .A1(new_n1822_), .B0(new_n3908_), .B1(new_n1126_), .Y(new_n5165_));
  OAI21X1  g05101(.A0(new_n3627_), .A1(new_n1189_), .B0(new_n5165_), .Y(new_n5166_));
  AOI21X1  g05102(.A0(new_n3624_), .A1(new_n2963_), .B0(new_n5166_), .Y(new_n5167_));
  XOR2X1   g05103(.A(new_n5167_), .B(\a[14] ), .Y(new_n5168_));
  INVX1    g05104(.A(new_n5168_), .Y(new_n5169_));
  XOR2X1   g05105(.A(new_n5065_), .B(new_n5064_), .Y(new_n5170_));
  AND2X1   g05106(.A(new_n5170_), .B(new_n5169_), .Y(new_n5171_));
  XOR2X1   g05107(.A(new_n5170_), .B(new_n5168_), .Y(new_n5172_));
  INVX1    g05108(.A(new_n5172_), .Y(new_n5173_));
  AOI22X1  g05109(.A0(new_n3984_), .A1(new_n1126_), .B0(new_n3628_), .B1(new_n2977_), .Y(new_n5174_));
  OAI21X1  g05110(.A0(new_n3907_), .A1(new_n1189_), .B0(new_n5174_), .Y(new_n5175_));
  AOI21X1  g05111(.A0(new_n3624_), .A1(new_n2976_), .B0(new_n5175_), .Y(new_n5176_));
  XOR2X1   g05112(.A(new_n5176_), .B(\a[14] ), .Y(new_n5177_));
  XOR2X1   g05113(.A(new_n4948_), .B(new_n4944_), .Y(new_n5178_));
  XOR2X1   g05114(.A(new_n5178_), .B(new_n5061_), .Y(new_n5179_));
  OR2X1    g05115(.A(new_n5179_), .B(new_n5177_), .Y(new_n5180_));
  XOR2X1   g05116(.A(new_n5179_), .B(new_n5177_), .Y(new_n5181_));
  INVX1    g05117(.A(new_n5181_), .Y(new_n5182_));
  INVX1    g05118(.A(new_n4957_), .Y(new_n5183_));
  XOR2X1   g05119(.A(new_n5059_), .B(new_n5183_), .Y(new_n5184_));
  OAI22X1  g05120(.A0(new_n3983_), .A1(new_n1189_), .B0(new_n3907_), .B1(new_n1236_), .Y(new_n5185_));
  AOI21X1  g05121(.A0(new_n3628_), .A1(new_n3342_), .B0(new_n5185_), .Y(new_n5186_));
  OAI21X1  g05122(.A0(new_n3906_), .A1(new_n3180_), .B0(new_n5186_), .Y(new_n5187_));
  XOR2X1   g05123(.A(new_n5187_), .B(new_n2529_), .Y(new_n5188_));
  NOR2X1   g05124(.A(new_n5188_), .B(new_n5184_), .Y(new_n5189_));
  XOR2X1   g05125(.A(new_n5058_), .B(new_n4964_), .Y(new_n5190_));
  INVX1    g05126(.A(new_n5190_), .Y(new_n5191_));
  OAI22X1  g05127(.A0(new_n3983_), .A1(new_n1236_), .B0(new_n3627_), .B1(new_n1339_), .Y(new_n5192_));
  AOI21X1  g05128(.A0(new_n3908_), .A1(new_n3342_), .B0(new_n5192_), .Y(new_n5193_));
  OAI21X1  g05129(.A0(new_n3906_), .A1(new_n3053_), .B0(new_n5193_), .Y(new_n5194_));
  XOR2X1   g05130(.A(new_n5194_), .B(new_n2529_), .Y(new_n5195_));
  OR2X1    g05131(.A(new_n5195_), .B(new_n5191_), .Y(new_n5196_));
  XOR2X1   g05132(.A(new_n5057_), .B(new_n4972_), .Y(new_n5197_));
  INVX1    g05133(.A(new_n5197_), .Y(new_n5198_));
  OAI22X1  g05134(.A0(new_n3983_), .A1(new_n1294_), .B0(new_n3627_), .B1(new_n1358_), .Y(new_n5199_));
  AOI21X1  g05135(.A0(new_n3908_), .A1(new_n3055_), .B0(new_n5199_), .Y(new_n5200_));
  OAI21X1  g05136(.A0(new_n3906_), .A1(new_n3340_), .B0(new_n5200_), .Y(new_n5201_));
  XOR2X1   g05137(.A(new_n5201_), .B(new_n2529_), .Y(new_n5202_));
  NOR2X1   g05138(.A(new_n5202_), .B(new_n5198_), .Y(new_n5203_));
  INVX1    g05139(.A(new_n5203_), .Y(new_n5204_));
  AOI22X1  g05140(.A0(new_n3984_), .A1(new_n3055_), .B0(new_n3908_), .B1(new_n1357_), .Y(new_n5205_));
  OAI21X1  g05141(.A0(new_n3627_), .A1(new_n1389_), .B0(new_n5205_), .Y(new_n5206_));
  AOI21X1  g05142(.A0(new_n3624_), .A1(new_n3425_), .B0(new_n5206_), .Y(new_n5207_));
  XOR2X1   g05143(.A(new_n5207_), .B(\a[14] ), .Y(new_n5208_));
  INVX1    g05144(.A(new_n5208_), .Y(new_n5209_));
  XOR2X1   g05145(.A(new_n5056_), .B(new_n5055_), .Y(new_n5210_));
  XOR2X1   g05146(.A(new_n5210_), .B(new_n5208_), .Y(new_n5211_));
  AOI22X1  g05147(.A0(new_n3984_), .A1(new_n1357_), .B0(new_n3628_), .B1(new_n3327_), .Y(new_n5212_));
  OAI21X1  g05148(.A0(new_n3907_), .A1(new_n1389_), .B0(new_n5212_), .Y(new_n5213_));
  AOI21X1  g05149(.A0(new_n3624_), .A1(new_n3326_), .B0(new_n5213_), .Y(new_n5214_));
  XOR2X1   g05150(.A(new_n5214_), .B(\a[14] ), .Y(new_n5215_));
  XOR2X1   g05151(.A(new_n4984_), .B(new_n4980_), .Y(new_n5216_));
  XOR2X1   g05152(.A(new_n5216_), .B(new_n5052_), .Y(new_n5217_));
  NOR2X1   g05153(.A(new_n5217_), .B(new_n5215_), .Y(new_n5218_));
  XOR2X1   g05154(.A(new_n5217_), .B(new_n5215_), .Y(new_n5219_));
  AOI22X1  g05155(.A0(new_n3908_), .A1(new_n3327_), .B0(new_n3628_), .B1(new_n1800_), .Y(new_n5220_));
  OAI21X1  g05156(.A0(new_n3983_), .A1(new_n1389_), .B0(new_n5220_), .Y(new_n5221_));
  AOI21X1  g05157(.A0(new_n3624_), .A1(new_n3497_), .B0(new_n5221_), .Y(new_n5222_));
  XOR2X1   g05158(.A(new_n5222_), .B(\a[14] ), .Y(new_n5223_));
  AND2X1   g05159(.A(new_n5049_), .B(new_n5000_), .Y(new_n5224_));
  INVX1    g05160(.A(new_n5050_), .Y(new_n5225_));
  XOR2X1   g05161(.A(new_n5225_), .B(new_n5224_), .Y(new_n5226_));
  OR2X1    g05162(.A(new_n5226_), .B(new_n5223_), .Y(new_n5227_));
  XOR2X1   g05163(.A(new_n5226_), .B(new_n5223_), .Y(new_n5228_));
  INVX1    g05164(.A(new_n5228_), .Y(new_n5229_));
  INVX1    g05165(.A(new_n5001_), .Y(new_n5230_));
  XOR2X1   g05166(.A(new_n5048_), .B(new_n5230_), .Y(new_n5231_));
  OAI22X1  g05167(.A0(new_n3983_), .A1(new_n1423_), .B0(new_n3627_), .B1(new_n3669_), .Y(new_n5232_));
  AOI21X1  g05168(.A0(new_n3908_), .A1(new_n1800_), .B0(new_n5232_), .Y(new_n5233_));
  OAI21X1  g05169(.A0(new_n3667_), .A1(new_n3906_), .B0(new_n5233_), .Y(new_n5234_));
  XOR2X1   g05170(.A(new_n5234_), .B(new_n2529_), .Y(new_n5235_));
  NOR2X1   g05171(.A(new_n5235_), .B(new_n5231_), .Y(new_n5236_));
  XOR2X1   g05172(.A(new_n5047_), .B(new_n5046_), .Y(new_n5237_));
  INVX1    g05173(.A(new_n5237_), .Y(new_n5238_));
  OAI22X1  g05174(.A0(new_n3983_), .A1(new_n1465_), .B0(new_n3907_), .B1(new_n3669_), .Y(new_n5239_));
  AOI21X1  g05175(.A0(new_n3628_), .A1(new_n1536_), .B0(new_n5239_), .Y(new_n5240_));
  OAI21X1  g05176(.A0(new_n3676_), .A1(new_n3906_), .B0(new_n5240_), .Y(new_n5241_));
  XOR2X1   g05177(.A(new_n5241_), .B(new_n2529_), .Y(new_n5242_));
  OR2X1    g05178(.A(new_n5242_), .B(new_n5238_), .Y(new_n5243_));
  XOR2X1   g05179(.A(new_n5044_), .B(new_n5019_), .Y(new_n5244_));
  OAI22X1  g05180(.A0(new_n3983_), .A1(new_n3669_), .B0(new_n3627_), .B1(new_n1586_), .Y(new_n5245_));
  AOI21X1  g05181(.A0(new_n3908_), .A1(new_n1536_), .B0(new_n5245_), .Y(new_n5246_));
  OAI21X1  g05182(.A0(new_n3906_), .A1(new_n3478_), .B0(new_n5246_), .Y(new_n5247_));
  XOR2X1   g05183(.A(new_n5247_), .B(\a[14] ), .Y(new_n5248_));
  AOI22X1  g05184(.A0(new_n3984_), .A1(new_n1536_), .B0(new_n3908_), .B1(new_n3480_), .Y(new_n5249_));
  OAI21X1  g05185(.A0(new_n3627_), .A1(new_n1621_), .B0(new_n5249_), .Y(new_n5250_));
  AOI21X1  g05186(.A0(new_n3697_), .A1(new_n3624_), .B0(new_n5250_), .Y(new_n5251_));
  XOR2X1   g05187(.A(new_n5251_), .B(\a[14] ), .Y(new_n5252_));
  INVX1    g05188(.A(new_n5252_), .Y(new_n5253_));
  XOR2X1   g05189(.A(new_n5043_), .B(new_n5042_), .Y(new_n5254_));
  AND2X1   g05190(.A(new_n5254_), .B(new_n5253_), .Y(new_n5255_));
  INVX1    g05191(.A(new_n5255_), .Y(new_n5256_));
  XOR2X1   g05192(.A(new_n5254_), .B(new_n5252_), .Y(new_n5257_));
  INVX1    g05193(.A(new_n5041_), .Y(new_n5258_));
  XOR2X1   g05194(.A(new_n5258_), .B(new_n5037_), .Y(new_n5259_));
  OAI22X1  g05195(.A0(new_n3983_), .A1(new_n1586_), .B0(new_n3627_), .B1(new_n1655_), .Y(new_n5260_));
  AOI21X1  g05196(.A0(new_n3908_), .A1(new_n4538_), .B0(new_n5260_), .Y(new_n5261_));
  OAI21X1  g05197(.A0(new_n3719_), .A1(new_n3906_), .B0(new_n5261_), .Y(new_n5262_));
  XOR2X1   g05198(.A(new_n5262_), .B(new_n2529_), .Y(new_n5263_));
  NOR2X1   g05199(.A(new_n5263_), .B(new_n5259_), .Y(new_n5264_));
  AOI22X1  g05200(.A0(new_n3908_), .A1(new_n3721_), .B0(new_n3628_), .B1(new_n1676_), .Y(new_n5265_));
  OAI21X1  g05201(.A0(new_n3983_), .A1(new_n1621_), .B0(new_n5265_), .Y(new_n5266_));
  AOI21X1  g05202(.A0(new_n3745_), .A1(new_n3624_), .B0(new_n5266_), .Y(new_n5267_));
  XOR2X1   g05203(.A(new_n5267_), .B(\a[14] ), .Y(new_n5268_));
  INVX1    g05204(.A(new_n5031_), .Y(new_n5269_));
  NAND3X1  g05205(.A(new_n5269_), .B(new_n5028_), .C(\a[17] ), .Y(new_n5270_));
  XOR2X1   g05206(.A(new_n5034_), .B(new_n2445_), .Y(new_n5271_));
  AND2X1   g05207(.A(new_n5271_), .B(new_n5270_), .Y(new_n5272_));
  NOR3X1   g05208(.A(new_n5272_), .B(new_n5268_), .C(new_n5035_), .Y(new_n5273_));
  XOR2X1   g05209(.A(new_n5271_), .B(new_n5270_), .Y(new_n5274_));
  XOR2X1   g05210(.A(new_n5274_), .B(new_n5268_), .Y(new_n5275_));
  AOI21X1  g05211(.A0(new_n5030_), .A1(new_n3821_), .B0(new_n2445_), .Y(new_n5276_));
  XOR2X1   g05212(.A(new_n5276_), .B(new_n5029_), .Y(new_n5277_));
  OAI22X1  g05213(.A0(new_n3983_), .A1(new_n1655_), .B0(new_n3907_), .B1(new_n1674_), .Y(new_n5278_));
  AOI21X1  g05214(.A0(new_n3628_), .A1(new_n1706_), .B0(new_n5278_), .Y(new_n5279_));
  OAI21X1  g05215(.A0(new_n3773_), .A1(new_n3906_), .B0(new_n5279_), .Y(new_n5280_));
  XOR2X1   g05216(.A(new_n5280_), .B(new_n2529_), .Y(new_n5281_));
  NOR2X1   g05217(.A(new_n5281_), .B(new_n5277_), .Y(new_n5282_));
  OAI22X1  g05218(.A0(new_n3983_), .A1(new_n1735_), .B0(new_n3907_), .B1(new_n1784_), .Y(new_n5283_));
  AOI21X1  g05219(.A0(new_n4165_), .A1(new_n3624_), .B0(new_n5283_), .Y(new_n5284_));
  XOR2X1   g05220(.A(new_n5284_), .B(\a[14] ), .Y(new_n5285_));
  INVX1    g05221(.A(new_n3621_), .Y(new_n5286_));
  AND2X1   g05222(.A(new_n5286_), .B(new_n3821_), .Y(new_n5287_));
  OAI22X1  g05223(.A0(new_n3907_), .A1(new_n1735_), .B0(new_n3627_), .B1(new_n1784_), .Y(new_n5288_));
  AOI21X1  g05224(.A0(new_n3984_), .A1(new_n1706_), .B0(new_n5288_), .Y(new_n5289_));
  OAI21X1  g05225(.A0(new_n4177_), .A1(new_n3906_), .B0(new_n5289_), .Y(new_n5290_));
  NOR4X1   g05226(.A(new_n5290_), .B(new_n5287_), .C(new_n5285_), .D(new_n2529_), .Y(new_n5291_));
  NAND2X1  g05227(.A(new_n5291_), .B(new_n5031_), .Y(new_n5292_));
  XOR2X1   g05228(.A(new_n5291_), .B(new_n5269_), .Y(new_n5293_));
  AOI22X1  g05229(.A0(new_n3984_), .A1(new_n1676_), .B0(new_n3628_), .B1(new_n3819_), .Y(new_n5294_));
  OAI21X1  g05230(.A0(new_n3907_), .A1(new_n1708_), .B0(new_n5294_), .Y(new_n5295_));
  AOI21X1  g05231(.A0(new_n3829_), .A1(new_n3624_), .B0(new_n5295_), .Y(new_n5296_));
  XOR2X1   g05232(.A(new_n5296_), .B(\a[14] ), .Y(new_n5297_));
  OAI21X1  g05233(.A0(new_n5297_), .A1(new_n5293_), .B0(new_n5292_), .Y(new_n5298_));
  XOR2X1   g05234(.A(new_n5281_), .B(new_n5277_), .Y(new_n5299_));
  AOI21X1  g05235(.A0(new_n5299_), .A1(new_n5298_), .B0(new_n5282_), .Y(new_n5300_));
  NOR2X1   g05236(.A(new_n5300_), .B(new_n5275_), .Y(new_n5301_));
  OR2X1    g05237(.A(new_n5301_), .B(new_n5273_), .Y(new_n5302_));
  XOR2X1   g05238(.A(new_n5263_), .B(new_n5259_), .Y(new_n5303_));
  AOI21X1  g05239(.A0(new_n5303_), .A1(new_n5302_), .B0(new_n5264_), .Y(new_n5304_));
  OR2X1    g05240(.A(new_n5304_), .B(new_n5257_), .Y(new_n5305_));
  XOR2X1   g05241(.A(new_n5247_), .B(new_n2529_), .Y(new_n5306_));
  XOR2X1   g05242(.A(new_n5306_), .B(new_n5244_), .Y(new_n5307_));
  AOI21X1  g05243(.A0(new_n5305_), .A1(new_n5256_), .B0(new_n5307_), .Y(new_n5308_));
  AOI21X1  g05244(.A0(new_n5248_), .A1(new_n5244_), .B0(new_n5308_), .Y(new_n5309_));
  XOR2X1   g05245(.A(new_n5242_), .B(new_n5237_), .Y(new_n5310_));
  OAI21X1  g05246(.A0(new_n5310_), .A1(new_n5309_), .B0(new_n5243_), .Y(new_n5311_));
  XOR2X1   g05247(.A(new_n5235_), .B(new_n5231_), .Y(new_n5312_));
  AOI21X1  g05248(.A0(new_n5312_), .A1(new_n5311_), .B0(new_n5236_), .Y(new_n5313_));
  OAI21X1  g05249(.A0(new_n5313_), .A1(new_n5229_), .B0(new_n5227_), .Y(new_n5314_));
  AOI21X1  g05250(.A0(new_n5314_), .A1(new_n5219_), .B0(new_n5218_), .Y(new_n5315_));
  NOR2X1   g05251(.A(new_n5315_), .B(new_n5211_), .Y(new_n5316_));
  AOI21X1  g05252(.A0(new_n5210_), .A1(new_n5209_), .B0(new_n5316_), .Y(new_n5317_));
  XOR2X1   g05253(.A(new_n5202_), .B(new_n5197_), .Y(new_n5318_));
  OAI21X1  g05254(.A0(new_n5318_), .A1(new_n5317_), .B0(new_n5204_), .Y(new_n5319_));
  INVX1    g05255(.A(new_n5319_), .Y(new_n5320_));
  XOR2X1   g05256(.A(new_n5195_), .B(new_n5190_), .Y(new_n5321_));
  OAI21X1  g05257(.A0(new_n5321_), .A1(new_n5320_), .B0(new_n5196_), .Y(new_n5322_));
  XOR2X1   g05258(.A(new_n5188_), .B(new_n5184_), .Y(new_n5323_));
  AOI21X1  g05259(.A0(new_n5323_), .A1(new_n5322_), .B0(new_n5189_), .Y(new_n5324_));
  OAI21X1  g05260(.A0(new_n5324_), .A1(new_n5182_), .B0(new_n5180_), .Y(new_n5325_));
  AOI21X1  g05261(.A0(new_n5325_), .A1(new_n5173_), .B0(new_n5171_), .Y(new_n5326_));
  XOR2X1   g05262(.A(new_n5162_), .B(new_n5157_), .Y(new_n5327_));
  OR2X1    g05263(.A(new_n5327_), .B(new_n5326_), .Y(new_n5328_));
  XOR2X1   g05264(.A(new_n5155_), .B(new_n2529_), .Y(new_n5329_));
  XOR2X1   g05265(.A(new_n5329_), .B(new_n5152_), .Y(new_n5330_));
  AOI21X1  g05266(.A0(new_n5328_), .A1(new_n5164_), .B0(new_n5330_), .Y(new_n5331_));
  AOI21X1  g05267(.A0(new_n5156_), .A1(new_n5152_), .B0(new_n5331_), .Y(new_n5332_));
  XOR2X1   g05268(.A(new_n5149_), .B(new_n2529_), .Y(new_n5333_));
  XOR2X1   g05269(.A(new_n5333_), .B(new_n5146_), .Y(new_n5334_));
  NOR2X1   g05270(.A(new_n5334_), .B(new_n5332_), .Y(new_n5335_));
  XOR2X1   g05271(.A(new_n5142_), .B(new_n2529_), .Y(new_n5336_));
  XOR2X1   g05272(.A(new_n5336_), .B(new_n5139_), .Y(new_n5337_));
  INVX1    g05273(.A(new_n5337_), .Y(new_n5338_));
  OAI21X1  g05274(.A0(new_n5335_), .A1(new_n5151_), .B0(new_n5338_), .Y(new_n5339_));
  XOR2X1   g05275(.A(new_n5137_), .B(new_n2529_), .Y(new_n5340_));
  XOR2X1   g05276(.A(new_n5340_), .B(new_n5134_), .Y(new_n5341_));
  AOI21X1  g05277(.A0(new_n5339_), .A1(new_n5145_), .B0(new_n5341_), .Y(new_n5342_));
  AOI21X1  g05278(.A0(new_n5138_), .A1(new_n5134_), .B0(new_n5342_), .Y(new_n5343_));
  XOR2X1   g05279(.A(new_n5131_), .B(new_n5126_), .Y(new_n5344_));
  OR2X1    g05280(.A(new_n5344_), .B(new_n5343_), .Y(new_n5345_));
  AND2X1   g05281(.A(new_n5345_), .B(new_n5133_), .Y(new_n5346_));
  XOR2X1   g05282(.A(new_n5123_), .B(new_n2529_), .Y(new_n5347_));
  XOR2X1   g05283(.A(new_n5347_), .B(new_n5119_), .Y(new_n5348_));
  NOR2X1   g05284(.A(new_n5348_), .B(new_n5346_), .Y(new_n5349_));
  XOR2X1   g05285(.A(new_n5083_), .B(new_n5082_), .Y(new_n5350_));
  OAI21X1  g05286(.A0(new_n5349_), .A1(new_n5125_), .B0(new_n5350_), .Y(new_n5351_));
  AOI22X1  g05287(.A0(new_n4428_), .A1(new_n2093_), .B0(new_n4078_), .B1(new_n1887_), .Y(new_n5352_));
  OAI21X1  g05288(.A0(new_n4246_), .A1(new_n2183_), .B0(new_n5352_), .Y(new_n5353_));
  AOI21X1  g05289(.A0(new_n4080_), .A1(new_n2430_), .B0(new_n5353_), .Y(new_n5354_));
  XOR2X1   g05290(.A(new_n5354_), .B(\a[11] ), .Y(new_n5355_));
  NOR2X1   g05291(.A(new_n5349_), .B(new_n5125_), .Y(new_n5356_));
  XOR2X1   g05292(.A(new_n5350_), .B(new_n5356_), .Y(new_n5357_));
  OR2X1    g05293(.A(new_n5357_), .B(new_n5355_), .Y(new_n5358_));
  AND2X1   g05294(.A(new_n5358_), .B(new_n5351_), .Y(new_n5359_));
  OR2X1    g05295(.A(new_n5359_), .B(new_n5118_), .Y(new_n5360_));
  XOR2X1   g05296(.A(new_n5359_), .B(new_n5118_), .Y(new_n5361_));
  INVX1    g05297(.A(new_n5361_), .Y(new_n5362_));
  AOI22X1  g05298(.A0(new_n4870_), .A1(new_n2420_), .B0(new_n4635_), .B1(new_n2627_), .Y(new_n5363_));
  OAI21X1  g05299(.A0(new_n5096_), .A1(new_n2379_), .B0(new_n5363_), .Y(new_n5364_));
  AOI21X1  g05300(.A0(new_n4637_), .A1(new_n2625_), .B0(new_n5364_), .Y(new_n5365_));
  XOR2X1   g05301(.A(new_n5365_), .B(\a[8] ), .Y(new_n5366_));
  OR2X1    g05302(.A(new_n5366_), .B(new_n5362_), .Y(new_n5367_));
  AND2X1   g05303(.A(new_n5367_), .B(new_n5360_), .Y(new_n5368_));
  INVX1    g05304(.A(new_n66_), .Y(new_n5369_));
  XOR2X1   g05305(.A(\a[4] ), .B(\a[3] ), .Y(new_n5370_));
  INVX1    g05306(.A(new_n5370_), .Y(new_n5371_));
  NAND3X1  g05307(.A(new_n5371_), .B(new_n5369_), .C(new_n65_), .Y(new_n5372_));
  INVX1    g05308(.A(new_n5372_), .Y(new_n5373_));
  AOI22X1  g05309(.A0(new_n5373_), .A1(new_n2649_), .B0(new_n2652_), .B1(new_n67_), .Y(new_n5374_));
  XOR2X1   g05310(.A(new_n5374_), .B(\a[5] ), .Y(new_n5375_));
  NOR2X1   g05311(.A(new_n5375_), .B(new_n5368_), .Y(new_n5376_));
  XOR2X1   g05312(.A(new_n5101_), .B(new_n5094_), .Y(new_n5377_));
  INVX1    g05313(.A(new_n5377_), .Y(new_n5378_));
  XOR2X1   g05314(.A(new_n5375_), .B(new_n5368_), .Y(new_n5379_));
  AOI21X1  g05315(.A0(new_n5379_), .A1(new_n5378_), .B0(new_n5376_), .Y(new_n5380_));
  INVX1    g05316(.A(new_n5380_), .Y(new_n5381_));
  OR2X1    g05317(.A(new_n5108_), .B(new_n5102_), .Y(new_n5382_));
  AOI21X1  g05318(.A0(new_n5108_), .A1(new_n5102_), .B0(new_n5111_), .Y(new_n5383_));
  AOI22X1  g05319(.A0(new_n5383_), .A1(new_n5382_), .B0(new_n5111_), .B1(new_n5110_), .Y(new_n5384_));
  AND2X1   g05320(.A(new_n5384_), .B(new_n5381_), .Y(new_n5385_));
  XOR2X1   g05321(.A(new_n5379_), .B(new_n5377_), .Y(new_n5386_));
  AOI22X1  g05322(.A0(new_n4428_), .A1(new_n2246_), .B0(new_n4078_), .B1(new_n2048_), .Y(new_n5387_));
  OAI21X1  g05323(.A0(new_n4246_), .A1(new_n1879_), .B0(new_n5387_), .Y(new_n5388_));
  AOI21X1  g05324(.A0(new_n4080_), .A1(new_n2244_), .B0(new_n5388_), .Y(new_n5389_));
  XOR2X1   g05325(.A(new_n5389_), .B(\a[11] ), .Y(new_n5390_));
  XOR2X1   g05326(.A(new_n5124_), .B(new_n5119_), .Y(new_n5391_));
  XOR2X1   g05327(.A(new_n5391_), .B(new_n5346_), .Y(new_n5392_));
  OR2X1    g05328(.A(new_n5392_), .B(new_n5390_), .Y(new_n5393_));
  XOR2X1   g05329(.A(new_n5392_), .B(new_n5390_), .Y(new_n5394_));
  AOI22X1  g05330(.A0(new_n4428_), .A1(new_n1887_), .B0(new_n4078_), .B1(new_n1886_), .Y(new_n5395_));
  OAI21X1  g05331(.A0(new_n4246_), .A1(new_n520_), .B0(new_n5395_), .Y(new_n5396_));
  AOI21X1  g05332(.A0(new_n4080_), .A1(new_n1882_), .B0(new_n5396_), .Y(new_n5397_));
  XOR2X1   g05333(.A(new_n5397_), .B(new_n2911_), .Y(new_n5398_));
  XOR2X1   g05334(.A(new_n5344_), .B(new_n5343_), .Y(new_n5399_));
  AND2X1   g05335(.A(new_n5399_), .B(new_n5398_), .Y(new_n5400_));
  XOR2X1   g05336(.A(new_n5399_), .B(new_n5398_), .Y(new_n5401_));
  INVX1    g05337(.A(new_n5401_), .Y(new_n5402_));
  AOI22X1  g05338(.A0(new_n4428_), .A1(new_n2048_), .B0(new_n4078_), .B1(new_n2049_), .Y(new_n5403_));
  OAI21X1  g05339(.A0(new_n4246_), .A1(new_n623_), .B0(new_n5403_), .Y(new_n5404_));
  AOI21X1  g05340(.A0(new_n4080_), .A1(new_n2047_), .B0(new_n5404_), .Y(new_n5405_));
  XOR2X1   g05341(.A(new_n5405_), .B(\a[11] ), .Y(new_n5406_));
  AND2X1   g05342(.A(new_n5339_), .B(new_n5145_), .Y(new_n5407_));
  INVX1    g05343(.A(new_n5341_), .Y(new_n5408_));
  XOR2X1   g05344(.A(new_n5408_), .B(new_n5407_), .Y(new_n5409_));
  OR2X1    g05345(.A(new_n5409_), .B(new_n5406_), .Y(new_n5410_));
  XOR2X1   g05346(.A(new_n5409_), .B(new_n5406_), .Y(new_n5411_));
  INVX1    g05347(.A(new_n5411_), .Y(new_n5412_));
  AOI22X1  g05348(.A0(new_n4428_), .A1(new_n1886_), .B0(new_n4078_), .B1(new_n2036_), .Y(new_n5413_));
  OAI21X1  g05349(.A0(new_n4246_), .A1(new_n690_), .B0(new_n5413_), .Y(new_n5414_));
  AOI21X1  g05350(.A0(new_n4080_), .A1(new_n2035_), .B0(new_n5414_), .Y(new_n5415_));
  XOR2X1   g05351(.A(new_n5415_), .B(\a[11] ), .Y(new_n5416_));
  NOR2X1   g05352(.A(new_n5335_), .B(new_n5151_), .Y(new_n5417_));
  XOR2X1   g05353(.A(new_n5338_), .B(new_n5417_), .Y(new_n5418_));
  NOR2X1   g05354(.A(new_n5418_), .B(new_n5416_), .Y(new_n5419_));
  XOR2X1   g05355(.A(new_n5418_), .B(new_n5416_), .Y(new_n5420_));
  AOI22X1  g05356(.A0(new_n4428_), .A1(new_n2049_), .B0(new_n4078_), .B1(new_n2481_), .Y(new_n5421_));
  OAI21X1  g05357(.A0(new_n4246_), .A1(new_n783_), .B0(new_n5421_), .Y(new_n5422_));
  AOI21X1  g05358(.A0(new_n4080_), .A1(new_n2480_), .B0(new_n5422_), .Y(new_n5423_));
  XOR2X1   g05359(.A(new_n5423_), .B(\a[11] ), .Y(new_n5424_));
  INVX1    g05360(.A(new_n5334_), .Y(new_n5425_));
  XOR2X1   g05361(.A(new_n5425_), .B(new_n5332_), .Y(new_n5426_));
  NOR2X1   g05362(.A(new_n5426_), .B(new_n5424_), .Y(new_n5427_));
  XOR2X1   g05363(.A(new_n5426_), .B(new_n5424_), .Y(new_n5428_));
  INVX1    g05364(.A(new_n5428_), .Y(new_n5429_));
  AOI22X1  g05365(.A0(new_n4428_), .A1(new_n2036_), .B0(new_n4078_), .B1(new_n2602_), .Y(new_n5430_));
  OAI21X1  g05366(.A0(new_n4246_), .A1(new_n847_), .B0(new_n5430_), .Y(new_n5431_));
  AOI21X1  g05367(.A0(new_n4080_), .A1(new_n2494_), .B0(new_n5431_), .Y(new_n5432_));
  XOR2X1   g05368(.A(new_n5432_), .B(\a[11] ), .Y(new_n5433_));
  AND2X1   g05369(.A(new_n5328_), .B(new_n5164_), .Y(new_n5434_));
  INVX1    g05370(.A(new_n5330_), .Y(new_n5435_));
  XOR2X1   g05371(.A(new_n5435_), .B(new_n5434_), .Y(new_n5436_));
  NOR2X1   g05372(.A(new_n5436_), .B(new_n5433_), .Y(new_n5437_));
  INVX1    g05373(.A(new_n5437_), .Y(new_n5438_));
  XOR2X1   g05374(.A(new_n5436_), .B(new_n5433_), .Y(new_n5439_));
  INVX1    g05375(.A(new_n5439_), .Y(new_n5440_));
  AOI22X1  g05376(.A0(new_n4428_), .A1(new_n2481_), .B0(new_n4078_), .B1(new_n2835_), .Y(new_n5441_));
  OAI21X1  g05377(.A0(new_n4246_), .A1(new_n903_), .B0(new_n5441_), .Y(new_n5442_));
  AOI21X1  g05378(.A0(new_n4080_), .A1(new_n2709_), .B0(new_n5442_), .Y(new_n5443_));
  XOR2X1   g05379(.A(new_n5443_), .B(\a[11] ), .Y(new_n5444_));
  INVX1    g05380(.A(new_n5327_), .Y(new_n5445_));
  XOR2X1   g05381(.A(new_n5445_), .B(new_n5326_), .Y(new_n5446_));
  NOR2X1   g05382(.A(new_n5446_), .B(new_n5444_), .Y(new_n5447_));
  XOR2X1   g05383(.A(new_n5446_), .B(new_n5444_), .Y(new_n5448_));
  XOR2X1   g05384(.A(new_n5325_), .B(new_n5173_), .Y(new_n5449_));
  INVX1    g05385(.A(new_n5449_), .Y(new_n5450_));
  OAI22X1  g05386(.A0(new_n4427_), .A1(new_n903_), .B0(new_n4077_), .B1(new_n985_), .Y(new_n5451_));
  AOI21X1  g05387(.A0(new_n4247_), .A1(new_n2835_), .B0(new_n5451_), .Y(new_n5452_));
  OAI21X1  g05388(.A0(new_n4245_), .A1(new_n2600_), .B0(new_n5452_), .Y(new_n5453_));
  XOR2X1   g05389(.A(new_n5453_), .B(new_n2911_), .Y(new_n5454_));
  NOR2X1   g05390(.A(new_n5454_), .B(new_n5450_), .Y(new_n5455_));
  XOR2X1   g05391(.A(new_n5324_), .B(new_n5182_), .Y(new_n5456_));
  INVX1    g05392(.A(new_n5456_), .Y(new_n5457_));
  OAI22X1  g05393(.A0(new_n4427_), .A1(new_n957_), .B0(new_n4246_), .B1(new_n985_), .Y(new_n5458_));
  AOI21X1  g05394(.A0(new_n4078_), .A1(new_n1822_), .B0(new_n5458_), .Y(new_n5459_));
  OAI21X1  g05395(.A0(new_n4245_), .A1(new_n2833_), .B0(new_n5459_), .Y(new_n5460_));
  XOR2X1   g05396(.A(new_n5460_), .B(new_n2911_), .Y(new_n5461_));
  NOR2X1   g05397(.A(new_n5461_), .B(new_n5457_), .Y(new_n5462_));
  AOI22X1  g05398(.A0(new_n4428_), .A1(new_n2603_), .B0(new_n4078_), .B1(new_n1126_), .Y(new_n5463_));
  OAI21X1  g05399(.A0(new_n4246_), .A1(new_n1065_), .B0(new_n5463_), .Y(new_n5464_));
  AOI21X1  g05400(.A0(new_n4080_), .A1(new_n2824_), .B0(new_n5464_), .Y(new_n5465_));
  XOR2X1   g05401(.A(new_n5465_), .B(\a[11] ), .Y(new_n5466_));
  INVX1    g05402(.A(new_n5466_), .Y(new_n5467_));
  XOR2X1   g05403(.A(new_n5323_), .B(new_n5322_), .Y(new_n5468_));
  NAND2X1  g05404(.A(new_n5468_), .B(new_n5467_), .Y(new_n5469_));
  XOR2X1   g05405(.A(new_n5468_), .B(new_n5466_), .Y(new_n5470_));
  AOI22X1  g05406(.A0(new_n4428_), .A1(new_n1822_), .B0(new_n4247_), .B1(new_n1126_), .Y(new_n5471_));
  OAI21X1  g05407(.A0(new_n4077_), .A1(new_n1189_), .B0(new_n5471_), .Y(new_n5472_));
  AOI21X1  g05408(.A0(new_n4080_), .A1(new_n2963_), .B0(new_n5472_), .Y(new_n5473_));
  XOR2X1   g05409(.A(new_n5473_), .B(\a[11] ), .Y(new_n5474_));
  XOR2X1   g05410(.A(new_n5321_), .B(new_n5319_), .Y(new_n5475_));
  NOR2X1   g05411(.A(new_n5475_), .B(new_n5474_), .Y(new_n5476_));
  XOR2X1   g05412(.A(new_n5475_), .B(new_n5474_), .Y(new_n5477_));
  AOI22X1  g05413(.A0(new_n4428_), .A1(new_n1126_), .B0(new_n4078_), .B1(new_n2977_), .Y(new_n5478_));
  OAI21X1  g05414(.A0(new_n4246_), .A1(new_n1189_), .B0(new_n5478_), .Y(new_n5479_));
  AOI21X1  g05415(.A0(new_n4080_), .A1(new_n2976_), .B0(new_n5479_), .Y(new_n5480_));
  XOR2X1   g05416(.A(new_n5480_), .B(\a[11] ), .Y(new_n5481_));
  INVX1    g05417(.A(new_n5318_), .Y(new_n5482_));
  XOR2X1   g05418(.A(new_n5482_), .B(new_n5317_), .Y(new_n5483_));
  OR2X1    g05419(.A(new_n5483_), .B(new_n5481_), .Y(new_n5484_));
  XOR2X1   g05420(.A(new_n5483_), .B(new_n5481_), .Y(new_n5485_));
  INVX1    g05421(.A(new_n5485_), .Y(new_n5486_));
  INVX1    g05422(.A(new_n5211_), .Y(new_n5487_));
  XOR2X1   g05423(.A(new_n5315_), .B(new_n5487_), .Y(new_n5488_));
  OAI22X1  g05424(.A0(new_n4427_), .A1(new_n1189_), .B0(new_n4246_), .B1(new_n1236_), .Y(new_n5489_));
  AOI21X1  g05425(.A0(new_n4078_), .A1(new_n3342_), .B0(new_n5489_), .Y(new_n5490_));
  OAI21X1  g05426(.A0(new_n4245_), .A1(new_n3180_), .B0(new_n5490_), .Y(new_n5491_));
  XOR2X1   g05427(.A(new_n5491_), .B(new_n2911_), .Y(new_n5492_));
  NOR2X1   g05428(.A(new_n5492_), .B(new_n5488_), .Y(new_n5493_));
  XOR2X1   g05429(.A(new_n5314_), .B(new_n5219_), .Y(new_n5494_));
  INVX1    g05430(.A(new_n5494_), .Y(new_n5495_));
  OAI22X1  g05431(.A0(new_n4427_), .A1(new_n1236_), .B0(new_n4077_), .B1(new_n1339_), .Y(new_n5496_));
  AOI21X1  g05432(.A0(new_n4247_), .A1(new_n3342_), .B0(new_n5496_), .Y(new_n5497_));
  OAI21X1  g05433(.A0(new_n4245_), .A1(new_n3053_), .B0(new_n5497_), .Y(new_n5498_));
  XOR2X1   g05434(.A(new_n5498_), .B(new_n2911_), .Y(new_n5499_));
  OR2X1    g05435(.A(new_n5499_), .B(new_n5495_), .Y(new_n5500_));
  XOR2X1   g05436(.A(new_n5313_), .B(new_n5229_), .Y(new_n5501_));
  INVX1    g05437(.A(new_n5501_), .Y(new_n5502_));
  OAI22X1  g05438(.A0(new_n4427_), .A1(new_n1294_), .B0(new_n4077_), .B1(new_n1358_), .Y(new_n5503_));
  AOI21X1  g05439(.A0(new_n4247_), .A1(new_n3055_), .B0(new_n5503_), .Y(new_n5504_));
  OAI21X1  g05440(.A0(new_n4245_), .A1(new_n3340_), .B0(new_n5504_), .Y(new_n5505_));
  XOR2X1   g05441(.A(new_n5505_), .B(new_n2911_), .Y(new_n5506_));
  NOR2X1   g05442(.A(new_n5506_), .B(new_n5502_), .Y(new_n5507_));
  INVX1    g05443(.A(new_n5507_), .Y(new_n5508_));
  AOI22X1  g05444(.A0(new_n4428_), .A1(new_n3055_), .B0(new_n4247_), .B1(new_n1357_), .Y(new_n5509_));
  OAI21X1  g05445(.A0(new_n4077_), .A1(new_n1389_), .B0(new_n5509_), .Y(new_n5510_));
  AOI21X1  g05446(.A0(new_n4080_), .A1(new_n3425_), .B0(new_n5510_), .Y(new_n5511_));
  XOR2X1   g05447(.A(new_n5511_), .B(\a[11] ), .Y(new_n5512_));
  INVX1    g05448(.A(new_n5512_), .Y(new_n5513_));
  XOR2X1   g05449(.A(new_n5312_), .B(new_n5311_), .Y(new_n5514_));
  XOR2X1   g05450(.A(new_n5514_), .B(new_n5512_), .Y(new_n5515_));
  AOI22X1  g05451(.A0(new_n4428_), .A1(new_n1357_), .B0(new_n4078_), .B1(new_n3327_), .Y(new_n5516_));
  OAI21X1  g05452(.A0(new_n4246_), .A1(new_n1389_), .B0(new_n5516_), .Y(new_n5517_));
  AOI21X1  g05453(.A0(new_n4080_), .A1(new_n3326_), .B0(new_n5517_), .Y(new_n5518_));
  XOR2X1   g05454(.A(new_n5518_), .B(\a[11] ), .Y(new_n5519_));
  INVX1    g05455(.A(new_n5310_), .Y(new_n5520_));
  XOR2X1   g05456(.A(new_n5520_), .B(new_n5309_), .Y(new_n5521_));
  NOR2X1   g05457(.A(new_n5521_), .B(new_n5519_), .Y(new_n5522_));
  XOR2X1   g05458(.A(new_n5521_), .B(new_n5519_), .Y(new_n5523_));
  AOI22X1  g05459(.A0(new_n4247_), .A1(new_n3327_), .B0(new_n4078_), .B1(new_n1800_), .Y(new_n5524_));
  OAI21X1  g05460(.A0(new_n4427_), .A1(new_n1389_), .B0(new_n5524_), .Y(new_n5525_));
  AOI21X1  g05461(.A0(new_n4080_), .A1(new_n3497_), .B0(new_n5525_), .Y(new_n5526_));
  XOR2X1   g05462(.A(new_n5526_), .B(\a[11] ), .Y(new_n5527_));
  AND2X1   g05463(.A(new_n5305_), .B(new_n5256_), .Y(new_n5528_));
  INVX1    g05464(.A(new_n5307_), .Y(new_n5529_));
  XOR2X1   g05465(.A(new_n5529_), .B(new_n5528_), .Y(new_n5530_));
  OR2X1    g05466(.A(new_n5530_), .B(new_n5527_), .Y(new_n5531_));
  XOR2X1   g05467(.A(new_n5530_), .B(new_n5527_), .Y(new_n5532_));
  INVX1    g05468(.A(new_n5532_), .Y(new_n5533_));
  INVX1    g05469(.A(new_n5257_), .Y(new_n5534_));
  XOR2X1   g05470(.A(new_n5304_), .B(new_n5534_), .Y(new_n5535_));
  OAI22X1  g05471(.A0(new_n4427_), .A1(new_n1423_), .B0(new_n4077_), .B1(new_n3669_), .Y(new_n5536_));
  AOI21X1  g05472(.A0(new_n4247_), .A1(new_n1800_), .B0(new_n5536_), .Y(new_n5537_));
  OAI21X1  g05473(.A0(new_n4245_), .A1(new_n3667_), .B0(new_n5537_), .Y(new_n5538_));
  XOR2X1   g05474(.A(new_n5538_), .B(new_n2911_), .Y(new_n5539_));
  NOR2X1   g05475(.A(new_n5539_), .B(new_n5535_), .Y(new_n5540_));
  XOR2X1   g05476(.A(new_n5303_), .B(new_n5302_), .Y(new_n5541_));
  INVX1    g05477(.A(new_n5541_), .Y(new_n5542_));
  OAI22X1  g05478(.A0(new_n4427_), .A1(new_n1465_), .B0(new_n4246_), .B1(new_n3669_), .Y(new_n5543_));
  AOI21X1  g05479(.A0(new_n4078_), .A1(new_n1536_), .B0(new_n5543_), .Y(new_n5544_));
  OAI21X1  g05480(.A0(new_n4245_), .A1(new_n3676_), .B0(new_n5544_), .Y(new_n5545_));
  XOR2X1   g05481(.A(new_n5545_), .B(new_n2911_), .Y(new_n5546_));
  OR2X1    g05482(.A(new_n5546_), .B(new_n5542_), .Y(new_n5547_));
  XOR2X1   g05483(.A(new_n5300_), .B(new_n5275_), .Y(new_n5548_));
  OAI22X1  g05484(.A0(new_n4427_), .A1(new_n3669_), .B0(new_n4077_), .B1(new_n1586_), .Y(new_n5549_));
  AOI21X1  g05485(.A0(new_n4247_), .A1(new_n1536_), .B0(new_n5549_), .Y(new_n5550_));
  OAI21X1  g05486(.A0(new_n4245_), .A1(new_n3478_), .B0(new_n5550_), .Y(new_n5551_));
  XOR2X1   g05487(.A(new_n5551_), .B(\a[11] ), .Y(new_n5552_));
  AOI22X1  g05488(.A0(new_n4428_), .A1(new_n1536_), .B0(new_n4247_), .B1(new_n3480_), .Y(new_n5553_));
  OAI21X1  g05489(.A0(new_n4077_), .A1(new_n1621_), .B0(new_n5553_), .Y(new_n5554_));
  AOI21X1  g05490(.A0(new_n4080_), .A1(new_n3697_), .B0(new_n5554_), .Y(new_n5555_));
  XOR2X1   g05491(.A(new_n5555_), .B(\a[11] ), .Y(new_n5556_));
  INVX1    g05492(.A(new_n5556_), .Y(new_n5557_));
  XOR2X1   g05493(.A(new_n5299_), .B(new_n5298_), .Y(new_n5558_));
  AND2X1   g05494(.A(new_n5558_), .B(new_n5557_), .Y(new_n5559_));
  INVX1    g05495(.A(new_n5559_), .Y(new_n5560_));
  XOR2X1   g05496(.A(new_n5558_), .B(new_n5556_), .Y(new_n5561_));
  INVX1    g05497(.A(new_n5297_), .Y(new_n5562_));
  XOR2X1   g05498(.A(new_n5562_), .B(new_n5293_), .Y(new_n5563_));
  OAI22X1  g05499(.A0(new_n4427_), .A1(new_n1586_), .B0(new_n4077_), .B1(new_n1655_), .Y(new_n5564_));
  AOI21X1  g05500(.A0(new_n4247_), .A1(new_n4538_), .B0(new_n5564_), .Y(new_n5565_));
  OAI21X1  g05501(.A0(new_n4245_), .A1(new_n3719_), .B0(new_n5565_), .Y(new_n5566_));
  XOR2X1   g05502(.A(new_n5566_), .B(new_n2911_), .Y(new_n5567_));
  NOR2X1   g05503(.A(new_n5567_), .B(new_n5563_), .Y(new_n5568_));
  AOI22X1  g05504(.A0(new_n4247_), .A1(new_n3721_), .B0(new_n4078_), .B1(new_n1676_), .Y(new_n5569_));
  OAI21X1  g05505(.A0(new_n4427_), .A1(new_n1621_), .B0(new_n5569_), .Y(new_n5570_));
  AOI21X1  g05506(.A0(new_n4080_), .A1(new_n3745_), .B0(new_n5570_), .Y(new_n5571_));
  XOR2X1   g05507(.A(new_n5571_), .B(\a[11] ), .Y(new_n5572_));
  INVX1    g05508(.A(new_n5287_), .Y(new_n5573_));
  NAND3X1  g05509(.A(new_n5573_), .B(new_n5284_), .C(\a[14] ), .Y(new_n5574_));
  XOR2X1   g05510(.A(new_n5290_), .B(new_n2529_), .Y(new_n5575_));
  AND2X1   g05511(.A(new_n5575_), .B(new_n5574_), .Y(new_n5576_));
  NOR3X1   g05512(.A(new_n5576_), .B(new_n5572_), .C(new_n5291_), .Y(new_n5577_));
  XOR2X1   g05513(.A(new_n5575_), .B(new_n5574_), .Y(new_n5578_));
  XOR2X1   g05514(.A(new_n5578_), .B(new_n5572_), .Y(new_n5579_));
  AOI21X1  g05515(.A0(new_n5286_), .A1(new_n3821_), .B0(new_n2529_), .Y(new_n5580_));
  XOR2X1   g05516(.A(new_n5580_), .B(new_n5285_), .Y(new_n5581_));
  OAI22X1  g05517(.A0(new_n4427_), .A1(new_n1655_), .B0(new_n4246_), .B1(new_n1674_), .Y(new_n5582_));
  AOI21X1  g05518(.A0(new_n4078_), .A1(new_n1706_), .B0(new_n5582_), .Y(new_n5583_));
  OAI21X1  g05519(.A0(new_n4245_), .A1(new_n3773_), .B0(new_n5583_), .Y(new_n5584_));
  XOR2X1   g05520(.A(new_n5584_), .B(new_n2911_), .Y(new_n5585_));
  NOR2X1   g05521(.A(new_n5585_), .B(new_n5581_), .Y(new_n5586_));
  OAI22X1  g05522(.A0(new_n4427_), .A1(new_n1735_), .B0(new_n4246_), .B1(new_n1784_), .Y(new_n5587_));
  AOI21X1  g05523(.A0(new_n4165_), .A1(new_n4080_), .B0(new_n5587_), .Y(new_n5588_));
  XOR2X1   g05524(.A(new_n5588_), .B(\a[11] ), .Y(new_n5589_));
  AND2X1   g05525(.A(new_n4079_), .B(new_n3821_), .Y(new_n5590_));
  OAI22X1  g05526(.A0(new_n4246_), .A1(new_n1735_), .B0(new_n4077_), .B1(new_n1784_), .Y(new_n5591_));
  AOI21X1  g05527(.A0(new_n4428_), .A1(new_n1706_), .B0(new_n5591_), .Y(new_n5592_));
  OAI21X1  g05528(.A0(new_n4245_), .A1(new_n4177_), .B0(new_n5592_), .Y(new_n5593_));
  NOR4X1   g05529(.A(new_n5593_), .B(new_n5590_), .C(new_n5589_), .D(new_n2911_), .Y(new_n5594_));
  NAND2X1  g05530(.A(new_n5594_), .B(new_n5287_), .Y(new_n5595_));
  XOR2X1   g05531(.A(new_n5594_), .B(new_n5573_), .Y(new_n5596_));
  AOI22X1  g05532(.A0(new_n4428_), .A1(new_n1676_), .B0(new_n4078_), .B1(new_n3819_), .Y(new_n5597_));
  OAI21X1  g05533(.A0(new_n4246_), .A1(new_n1708_), .B0(new_n5597_), .Y(new_n5598_));
  AOI21X1  g05534(.A0(new_n4080_), .A1(new_n3829_), .B0(new_n5598_), .Y(new_n5599_));
  XOR2X1   g05535(.A(new_n5599_), .B(\a[11] ), .Y(new_n5600_));
  OAI21X1  g05536(.A0(new_n5600_), .A1(new_n5596_), .B0(new_n5595_), .Y(new_n5601_));
  XOR2X1   g05537(.A(new_n5585_), .B(new_n5581_), .Y(new_n5602_));
  AOI21X1  g05538(.A0(new_n5602_), .A1(new_n5601_), .B0(new_n5586_), .Y(new_n5603_));
  NOR2X1   g05539(.A(new_n5603_), .B(new_n5579_), .Y(new_n5604_));
  OR2X1    g05540(.A(new_n5604_), .B(new_n5577_), .Y(new_n5605_));
  XOR2X1   g05541(.A(new_n5567_), .B(new_n5563_), .Y(new_n5606_));
  AOI21X1  g05542(.A0(new_n5606_), .A1(new_n5605_), .B0(new_n5568_), .Y(new_n5607_));
  OR2X1    g05543(.A(new_n5607_), .B(new_n5561_), .Y(new_n5608_));
  XOR2X1   g05544(.A(new_n5551_), .B(new_n2911_), .Y(new_n5609_));
  XOR2X1   g05545(.A(new_n5609_), .B(new_n5548_), .Y(new_n5610_));
  AOI21X1  g05546(.A0(new_n5608_), .A1(new_n5560_), .B0(new_n5610_), .Y(new_n5611_));
  AOI21X1  g05547(.A0(new_n5552_), .A1(new_n5548_), .B0(new_n5611_), .Y(new_n5612_));
  XOR2X1   g05548(.A(new_n5546_), .B(new_n5541_), .Y(new_n5613_));
  OAI21X1  g05549(.A0(new_n5613_), .A1(new_n5612_), .B0(new_n5547_), .Y(new_n5614_));
  XOR2X1   g05550(.A(new_n5539_), .B(new_n5535_), .Y(new_n5615_));
  AOI21X1  g05551(.A0(new_n5615_), .A1(new_n5614_), .B0(new_n5540_), .Y(new_n5616_));
  OAI21X1  g05552(.A0(new_n5616_), .A1(new_n5533_), .B0(new_n5531_), .Y(new_n5617_));
  AOI21X1  g05553(.A0(new_n5617_), .A1(new_n5523_), .B0(new_n5522_), .Y(new_n5618_));
  NOR2X1   g05554(.A(new_n5618_), .B(new_n5515_), .Y(new_n5619_));
  AOI21X1  g05555(.A0(new_n5514_), .A1(new_n5513_), .B0(new_n5619_), .Y(new_n5620_));
  XOR2X1   g05556(.A(new_n5506_), .B(new_n5501_), .Y(new_n5621_));
  OAI21X1  g05557(.A0(new_n5621_), .A1(new_n5620_), .B0(new_n5508_), .Y(new_n5622_));
  INVX1    g05558(.A(new_n5622_), .Y(new_n5623_));
  XOR2X1   g05559(.A(new_n5499_), .B(new_n5494_), .Y(new_n5624_));
  OAI21X1  g05560(.A0(new_n5624_), .A1(new_n5623_), .B0(new_n5500_), .Y(new_n5625_));
  XOR2X1   g05561(.A(new_n5492_), .B(new_n5488_), .Y(new_n5626_));
  AOI21X1  g05562(.A0(new_n5626_), .A1(new_n5625_), .B0(new_n5493_), .Y(new_n5627_));
  OAI21X1  g05563(.A0(new_n5627_), .A1(new_n5486_), .B0(new_n5484_), .Y(new_n5628_));
  AOI21X1  g05564(.A0(new_n5628_), .A1(new_n5477_), .B0(new_n5476_), .Y(new_n5629_));
  OAI21X1  g05565(.A0(new_n5629_), .A1(new_n5470_), .B0(new_n5469_), .Y(new_n5630_));
  XOR2X1   g05566(.A(new_n5461_), .B(new_n5456_), .Y(new_n5631_));
  INVX1    g05567(.A(new_n5631_), .Y(new_n5632_));
  AOI21X1  g05568(.A0(new_n5632_), .A1(new_n5630_), .B0(new_n5462_), .Y(new_n5633_));
  INVX1    g05569(.A(new_n5633_), .Y(new_n5634_));
  XOR2X1   g05570(.A(new_n5454_), .B(new_n5450_), .Y(new_n5635_));
  AOI21X1  g05571(.A0(new_n5635_), .A1(new_n5634_), .B0(new_n5455_), .Y(new_n5636_));
  INVX1    g05572(.A(new_n5636_), .Y(new_n5637_));
  AOI21X1  g05573(.A0(new_n5637_), .A1(new_n5448_), .B0(new_n5447_), .Y(new_n5638_));
  OR2X1    g05574(.A(new_n5638_), .B(new_n5440_), .Y(new_n5639_));
  AOI21X1  g05575(.A0(new_n5639_), .A1(new_n5438_), .B0(new_n5429_), .Y(new_n5640_));
  NOR2X1   g05576(.A(new_n5640_), .B(new_n5427_), .Y(new_n5641_));
  INVX1    g05577(.A(new_n5641_), .Y(new_n5642_));
  AOI21X1  g05578(.A0(new_n5642_), .A1(new_n5420_), .B0(new_n5419_), .Y(new_n5643_));
  OR2X1    g05579(.A(new_n5643_), .B(new_n5412_), .Y(new_n5644_));
  AOI21X1  g05580(.A0(new_n5644_), .A1(new_n5410_), .B0(new_n5402_), .Y(new_n5645_));
  OAI21X1  g05581(.A0(new_n5645_), .A1(new_n5400_), .B0(new_n5394_), .Y(new_n5646_));
  AND2X1   g05582(.A(new_n5646_), .B(new_n5393_), .Y(new_n5647_));
  INVX1    g05583(.A(new_n5647_), .Y(new_n5648_));
  XOR2X1   g05584(.A(new_n5357_), .B(new_n5355_), .Y(new_n5649_));
  AOI22X1  g05585(.A0(new_n5097_), .A1(new_n2420_), .B0(new_n4635_), .B1(new_n2252_), .Y(new_n5650_));
  OAI21X1  g05586(.A0(new_n4869_), .A1(new_n2287_), .B0(new_n5650_), .Y(new_n5651_));
  AOI21X1  g05587(.A0(new_n4637_), .A1(new_n2669_), .B0(new_n5651_), .Y(new_n5652_));
  XOR2X1   g05588(.A(new_n5652_), .B(\a[8] ), .Y(new_n5653_));
  XOR2X1   g05589(.A(new_n5649_), .B(new_n5647_), .Y(new_n5654_));
  NOR2X1   g05590(.A(new_n5654_), .B(new_n5653_), .Y(new_n5655_));
  AOI21X1  g05591(.A0(new_n5649_), .A1(new_n5648_), .B0(new_n5655_), .Y(new_n5656_));
  INVX1    g05592(.A(new_n67_), .Y(new_n5657_));
  OR2X1    g05593(.A(new_n5371_), .B(new_n66_), .Y(new_n5658_));
  INVX1    g05594(.A(new_n5658_), .Y(new_n5659_));
  AOI22X1  g05595(.A0(new_n5659_), .A1(new_n2649_), .B0(new_n5373_), .B1(new_n2421_), .Y(new_n5660_));
  OAI21X1  g05596(.A0(new_n2695_), .A1(new_n5657_), .B0(new_n5660_), .Y(new_n5661_));
  XOR2X1   g05597(.A(new_n5661_), .B(new_n3289_), .Y(new_n5662_));
  NOR2X1   g05598(.A(new_n5662_), .B(new_n5656_), .Y(new_n5663_));
  XOR2X1   g05599(.A(new_n5366_), .B(new_n5362_), .Y(new_n5664_));
  XOR2X1   g05600(.A(new_n5662_), .B(new_n5656_), .Y(new_n5665_));
  AOI21X1  g05601(.A0(new_n5665_), .A1(new_n5664_), .B0(new_n5663_), .Y(new_n5666_));
  NOR2X1   g05602(.A(new_n5666_), .B(new_n5386_), .Y(new_n5667_));
  INVX1    g05603(.A(new_n5667_), .Y(new_n5668_));
  XOR2X1   g05604(.A(new_n5666_), .B(new_n5386_), .Y(new_n5669_));
  INVX1    g05605(.A(new_n5669_), .Y(new_n5670_));
  NOR2X1   g05606(.A(new_n5645_), .B(new_n5400_), .Y(new_n5671_));
  XOR2X1   g05607(.A(new_n5671_), .B(new_n5394_), .Y(new_n5672_));
  OAI22X1  g05608(.A0(new_n5096_), .A1(new_n2287_), .B0(new_n4634_), .B1(new_n2092_), .Y(new_n5673_));
  AOI21X1  g05609(.A0(new_n4870_), .A1(new_n2252_), .B0(new_n5673_), .Y(new_n5674_));
  OAI21X1  g05610(.A0(new_n4868_), .A1(new_n2295_), .B0(new_n5674_), .Y(new_n5675_));
  XOR2X1   g05611(.A(new_n5675_), .B(new_n2995_), .Y(new_n5676_));
  NOR2X1   g05612(.A(new_n5676_), .B(new_n5672_), .Y(new_n5677_));
  AND2X1   g05613(.A(new_n5644_), .B(new_n5410_), .Y(new_n5678_));
  XOR2X1   g05614(.A(new_n5678_), .B(new_n5402_), .Y(new_n5679_));
  INVX1    g05615(.A(new_n5679_), .Y(new_n5680_));
  OAI22X1  g05616(.A0(new_n5096_), .A1(new_n2137_), .B0(new_n4634_), .B1(new_n2183_), .Y(new_n5681_));
  AOI21X1  g05617(.A0(new_n4870_), .A1(new_n2093_), .B0(new_n5681_), .Y(new_n5682_));
  OAI21X1  g05618(.A0(new_n4868_), .A1(new_n2202_), .B0(new_n5682_), .Y(new_n5683_));
  XOR2X1   g05619(.A(new_n5683_), .B(new_n2995_), .Y(new_n5684_));
  OR2X1    g05620(.A(new_n5684_), .B(new_n5680_), .Y(new_n5685_));
  XOR2X1   g05621(.A(new_n5643_), .B(new_n5412_), .Y(new_n5686_));
  AOI22X1  g05622(.A0(new_n5097_), .A1(new_n2093_), .B0(new_n4635_), .B1(new_n1887_), .Y(new_n5687_));
  OAI21X1  g05623(.A0(new_n4869_), .A1(new_n2183_), .B0(new_n5687_), .Y(new_n5688_));
  AOI21X1  g05624(.A0(new_n4637_), .A1(new_n2430_), .B0(new_n5688_), .Y(new_n5689_));
  XOR2X1   g05625(.A(new_n5689_), .B(new_n2995_), .Y(new_n5690_));
  XOR2X1   g05626(.A(new_n5641_), .B(new_n5420_), .Y(new_n5691_));
  OAI22X1  g05627(.A0(new_n5096_), .A1(new_n2183_), .B0(new_n4634_), .B1(new_n520_), .Y(new_n5692_));
  AOI21X1  g05628(.A0(new_n4870_), .A1(new_n1887_), .B0(new_n5692_), .Y(new_n5693_));
  OAI21X1  g05629(.A0(new_n4868_), .A1(new_n2243_), .B0(new_n5693_), .Y(new_n5694_));
  XOR2X1   g05630(.A(new_n5694_), .B(new_n2995_), .Y(new_n5695_));
  NOR2X1   g05631(.A(new_n5695_), .B(new_n5691_), .Y(new_n5696_));
  INVX1    g05632(.A(new_n5696_), .Y(new_n5697_));
  AND2X1   g05633(.A(new_n5639_), .B(new_n5438_), .Y(new_n5698_));
  XOR2X1   g05634(.A(new_n5698_), .B(new_n5429_), .Y(new_n5699_));
  OAI22X1  g05635(.A0(new_n5096_), .A1(new_n1879_), .B0(new_n4634_), .B1(new_n623_), .Y(new_n5700_));
  AOI21X1  g05636(.A0(new_n4870_), .A1(new_n2048_), .B0(new_n5700_), .Y(new_n5701_));
  OAI21X1  g05637(.A0(new_n4868_), .A1(new_n1881_), .B0(new_n5701_), .Y(new_n5702_));
  XOR2X1   g05638(.A(new_n5702_), .B(\a[8] ), .Y(new_n5703_));
  AND2X1   g05639(.A(new_n5703_), .B(new_n5699_), .Y(new_n5704_));
  XOR2X1   g05640(.A(new_n5638_), .B(new_n5440_), .Y(new_n5705_));
  INVX1    g05641(.A(new_n5705_), .Y(new_n5706_));
  OAI22X1  g05642(.A0(new_n5096_), .A1(new_n520_), .B0(new_n4634_), .B1(new_n690_), .Y(new_n5707_));
  AOI21X1  g05643(.A0(new_n4870_), .A1(new_n1886_), .B0(new_n5707_), .Y(new_n5708_));
  OAI21X1  g05644(.A0(new_n4868_), .A1(new_n3114_), .B0(new_n5708_), .Y(new_n5709_));
  XOR2X1   g05645(.A(new_n5709_), .B(new_n2995_), .Y(new_n5710_));
  NOR2X1   g05646(.A(new_n5710_), .B(new_n5706_), .Y(new_n5711_));
  INVX1    g05647(.A(new_n5711_), .Y(new_n5712_));
  XOR2X1   g05648(.A(new_n5637_), .B(new_n5448_), .Y(new_n5713_));
  OAI22X1  g05649(.A0(new_n5096_), .A1(new_n623_), .B0(new_n4634_), .B1(new_n783_), .Y(new_n5714_));
  AOI21X1  g05650(.A0(new_n4870_), .A1(new_n2049_), .B0(new_n5714_), .Y(new_n5715_));
  OAI21X1  g05651(.A0(new_n4868_), .A1(new_n5120_), .B0(new_n5715_), .Y(new_n5716_));
  XOR2X1   g05652(.A(new_n5716_), .B(\a[8] ), .Y(new_n5717_));
  AOI22X1  g05653(.A0(new_n5097_), .A1(new_n2049_), .B0(new_n4635_), .B1(new_n2481_), .Y(new_n5718_));
  OAI21X1  g05654(.A0(new_n4869_), .A1(new_n783_), .B0(new_n5718_), .Y(new_n5719_));
  AOI21X1  g05655(.A0(new_n4637_), .A1(new_n2480_), .B0(new_n5719_), .Y(new_n5720_));
  XOR2X1   g05656(.A(new_n5720_), .B(\a[8] ), .Y(new_n5721_));
  XOR2X1   g05657(.A(new_n5635_), .B(new_n5633_), .Y(new_n5722_));
  NOR2X1   g05658(.A(new_n5722_), .B(new_n5721_), .Y(new_n5723_));
  XOR2X1   g05659(.A(new_n5635_), .B(new_n5634_), .Y(new_n5724_));
  XOR2X1   g05660(.A(new_n5724_), .B(new_n5721_), .Y(new_n5725_));
  INVX1    g05661(.A(new_n5725_), .Y(new_n5726_));
  AOI22X1  g05662(.A0(new_n5097_), .A1(new_n2036_), .B0(new_n4635_), .B1(new_n2602_), .Y(new_n5727_));
  OAI21X1  g05663(.A0(new_n4869_), .A1(new_n847_), .B0(new_n5727_), .Y(new_n5728_));
  AOI21X1  g05664(.A0(new_n4637_), .A1(new_n2494_), .B0(new_n5728_), .Y(new_n5729_));
  XOR2X1   g05665(.A(new_n5729_), .B(\a[8] ), .Y(new_n5730_));
  XOR2X1   g05666(.A(new_n5631_), .B(new_n5630_), .Y(new_n5731_));
  NOR2X1   g05667(.A(new_n5731_), .B(new_n5730_), .Y(new_n5732_));
  INVX1    g05668(.A(new_n5732_), .Y(new_n5733_));
  XOR2X1   g05669(.A(new_n5731_), .B(new_n5730_), .Y(new_n5734_));
  INVX1    g05670(.A(new_n5734_), .Y(new_n5735_));
  INVX1    g05671(.A(new_n5470_), .Y(new_n5736_));
  XOR2X1   g05672(.A(new_n5629_), .B(new_n5736_), .Y(new_n5737_));
  OAI22X1  g05673(.A0(new_n5096_), .A1(new_n847_), .B0(new_n4634_), .B1(new_n957_), .Y(new_n5738_));
  AOI21X1  g05674(.A0(new_n4870_), .A1(new_n2602_), .B0(new_n5738_), .Y(new_n5739_));
  OAI21X1  g05675(.A0(new_n4868_), .A1(new_n2708_), .B0(new_n5739_), .Y(new_n5740_));
  XOR2X1   g05676(.A(new_n5740_), .B(new_n2995_), .Y(new_n5741_));
  NOR2X1   g05677(.A(new_n5741_), .B(new_n5737_), .Y(new_n5742_));
  XOR2X1   g05678(.A(new_n5628_), .B(new_n5477_), .Y(new_n5743_));
  INVX1    g05679(.A(new_n5743_), .Y(new_n5744_));
  OAI22X1  g05680(.A0(new_n5096_), .A1(new_n903_), .B0(new_n4634_), .B1(new_n985_), .Y(new_n5745_));
  AOI21X1  g05681(.A0(new_n4870_), .A1(new_n2835_), .B0(new_n5745_), .Y(new_n5746_));
  OAI21X1  g05682(.A0(new_n4868_), .A1(new_n2600_), .B0(new_n5746_), .Y(new_n5747_));
  XOR2X1   g05683(.A(new_n5747_), .B(new_n2995_), .Y(new_n5748_));
  OR2X1    g05684(.A(new_n5748_), .B(new_n5744_), .Y(new_n5749_));
  XOR2X1   g05685(.A(new_n5627_), .B(new_n5486_), .Y(new_n5750_));
  INVX1    g05686(.A(new_n5750_), .Y(new_n5751_));
  OAI22X1  g05687(.A0(new_n5096_), .A1(new_n957_), .B0(new_n4869_), .B1(new_n985_), .Y(new_n5752_));
  AOI21X1  g05688(.A0(new_n4635_), .A1(new_n1822_), .B0(new_n5752_), .Y(new_n5753_));
  OAI21X1  g05689(.A0(new_n4868_), .A1(new_n2833_), .B0(new_n5753_), .Y(new_n5754_));
  XOR2X1   g05690(.A(new_n5754_), .B(new_n2995_), .Y(new_n5755_));
  NOR2X1   g05691(.A(new_n5755_), .B(new_n5751_), .Y(new_n5756_));
  AOI22X1  g05692(.A0(new_n5097_), .A1(new_n2603_), .B0(new_n4635_), .B1(new_n1126_), .Y(new_n5757_));
  OAI21X1  g05693(.A0(new_n4869_), .A1(new_n1065_), .B0(new_n5757_), .Y(new_n5758_));
  AOI21X1  g05694(.A0(new_n4637_), .A1(new_n2824_), .B0(new_n5758_), .Y(new_n5759_));
  XOR2X1   g05695(.A(new_n5759_), .B(\a[8] ), .Y(new_n5760_));
  INVX1    g05696(.A(new_n5760_), .Y(new_n5761_));
  XOR2X1   g05697(.A(new_n5626_), .B(new_n5625_), .Y(new_n5762_));
  NAND2X1  g05698(.A(new_n5762_), .B(new_n5761_), .Y(new_n5763_));
  XOR2X1   g05699(.A(new_n5762_), .B(new_n5760_), .Y(new_n5764_));
  AOI22X1  g05700(.A0(new_n5097_), .A1(new_n1822_), .B0(new_n4870_), .B1(new_n1126_), .Y(new_n5765_));
  OAI21X1  g05701(.A0(new_n4634_), .A1(new_n1189_), .B0(new_n5765_), .Y(new_n5766_));
  AOI21X1  g05702(.A0(new_n4637_), .A1(new_n2963_), .B0(new_n5766_), .Y(new_n5767_));
  XOR2X1   g05703(.A(new_n5767_), .B(\a[8] ), .Y(new_n5768_));
  XOR2X1   g05704(.A(new_n5624_), .B(new_n5622_), .Y(new_n5769_));
  NOR2X1   g05705(.A(new_n5769_), .B(new_n5768_), .Y(new_n5770_));
  XOR2X1   g05706(.A(new_n5769_), .B(new_n5768_), .Y(new_n5771_));
  AOI22X1  g05707(.A0(new_n5097_), .A1(new_n1126_), .B0(new_n4635_), .B1(new_n2977_), .Y(new_n5772_));
  OAI21X1  g05708(.A0(new_n4869_), .A1(new_n1189_), .B0(new_n5772_), .Y(new_n5773_));
  AOI21X1  g05709(.A0(new_n4637_), .A1(new_n2976_), .B0(new_n5773_), .Y(new_n5774_));
  XOR2X1   g05710(.A(new_n5774_), .B(\a[8] ), .Y(new_n5775_));
  INVX1    g05711(.A(new_n5621_), .Y(new_n5776_));
  XOR2X1   g05712(.A(new_n5776_), .B(new_n5620_), .Y(new_n5777_));
  NOR2X1   g05713(.A(new_n5777_), .B(new_n5775_), .Y(new_n5778_));
  INVX1    g05714(.A(new_n5778_), .Y(new_n5779_));
  XOR2X1   g05715(.A(new_n5777_), .B(new_n5775_), .Y(new_n5780_));
  INVX1    g05716(.A(new_n5780_), .Y(new_n5781_));
  INVX1    g05717(.A(new_n5515_), .Y(new_n5782_));
  XOR2X1   g05718(.A(new_n5618_), .B(new_n5782_), .Y(new_n5783_));
  OAI22X1  g05719(.A0(new_n5096_), .A1(new_n1189_), .B0(new_n4869_), .B1(new_n1236_), .Y(new_n5784_));
  AOI21X1  g05720(.A0(new_n4635_), .A1(new_n3342_), .B0(new_n5784_), .Y(new_n5785_));
  OAI21X1  g05721(.A0(new_n4868_), .A1(new_n3180_), .B0(new_n5785_), .Y(new_n5786_));
  XOR2X1   g05722(.A(new_n5786_), .B(new_n2995_), .Y(new_n5787_));
  NOR2X1   g05723(.A(new_n5787_), .B(new_n5783_), .Y(new_n5788_));
  XOR2X1   g05724(.A(new_n5617_), .B(new_n5523_), .Y(new_n5789_));
  INVX1    g05725(.A(new_n5789_), .Y(new_n5790_));
  OAI22X1  g05726(.A0(new_n5096_), .A1(new_n1236_), .B0(new_n4634_), .B1(new_n1339_), .Y(new_n5791_));
  AOI21X1  g05727(.A0(new_n4870_), .A1(new_n3342_), .B0(new_n5791_), .Y(new_n5792_));
  OAI21X1  g05728(.A0(new_n4868_), .A1(new_n3053_), .B0(new_n5792_), .Y(new_n5793_));
  XOR2X1   g05729(.A(new_n5793_), .B(new_n2995_), .Y(new_n5794_));
  OR2X1    g05730(.A(new_n5794_), .B(new_n5790_), .Y(new_n5795_));
  XOR2X1   g05731(.A(new_n5616_), .B(new_n5533_), .Y(new_n5796_));
  INVX1    g05732(.A(new_n5796_), .Y(new_n5797_));
  OAI22X1  g05733(.A0(new_n5096_), .A1(new_n1294_), .B0(new_n4634_), .B1(new_n1358_), .Y(new_n5798_));
  AOI21X1  g05734(.A0(new_n4870_), .A1(new_n3055_), .B0(new_n5798_), .Y(new_n5799_));
  OAI21X1  g05735(.A0(new_n4868_), .A1(new_n3340_), .B0(new_n5799_), .Y(new_n5800_));
  XOR2X1   g05736(.A(new_n5800_), .B(new_n2995_), .Y(new_n5801_));
  NOR2X1   g05737(.A(new_n5801_), .B(new_n5797_), .Y(new_n5802_));
  AOI22X1  g05738(.A0(new_n5097_), .A1(new_n3055_), .B0(new_n4870_), .B1(new_n1357_), .Y(new_n5803_));
  OAI21X1  g05739(.A0(new_n4634_), .A1(new_n1389_), .B0(new_n5803_), .Y(new_n5804_));
  AOI21X1  g05740(.A0(new_n4637_), .A1(new_n3425_), .B0(new_n5804_), .Y(new_n5805_));
  XOR2X1   g05741(.A(new_n5805_), .B(\a[8] ), .Y(new_n5806_));
  INVX1    g05742(.A(new_n5806_), .Y(new_n5807_));
  XOR2X1   g05743(.A(new_n5615_), .B(new_n5614_), .Y(new_n5808_));
  NAND2X1  g05744(.A(new_n5808_), .B(new_n5807_), .Y(new_n5809_));
  XOR2X1   g05745(.A(new_n5808_), .B(new_n5806_), .Y(new_n5810_));
  AOI22X1  g05746(.A0(new_n5097_), .A1(new_n1357_), .B0(new_n4635_), .B1(new_n3327_), .Y(new_n5811_));
  OAI21X1  g05747(.A0(new_n4869_), .A1(new_n1389_), .B0(new_n5811_), .Y(new_n5812_));
  AOI21X1  g05748(.A0(new_n4637_), .A1(new_n3326_), .B0(new_n5812_), .Y(new_n5813_));
  XOR2X1   g05749(.A(new_n5813_), .B(\a[8] ), .Y(new_n5814_));
  INVX1    g05750(.A(new_n5613_), .Y(new_n5815_));
  XOR2X1   g05751(.A(new_n5815_), .B(new_n5612_), .Y(new_n5816_));
  NOR2X1   g05752(.A(new_n5816_), .B(new_n5814_), .Y(new_n5817_));
  XOR2X1   g05753(.A(new_n5816_), .B(new_n5814_), .Y(new_n5818_));
  AOI22X1  g05754(.A0(new_n4870_), .A1(new_n3327_), .B0(new_n4635_), .B1(new_n1800_), .Y(new_n5819_));
  OAI21X1  g05755(.A0(new_n5096_), .A1(new_n1389_), .B0(new_n5819_), .Y(new_n5820_));
  AOI21X1  g05756(.A0(new_n4637_), .A1(new_n3497_), .B0(new_n5820_), .Y(new_n5821_));
  XOR2X1   g05757(.A(new_n5821_), .B(\a[8] ), .Y(new_n5822_));
  AND2X1   g05758(.A(new_n5608_), .B(new_n5560_), .Y(new_n5823_));
  INVX1    g05759(.A(new_n5610_), .Y(new_n5824_));
  XOR2X1   g05760(.A(new_n5824_), .B(new_n5823_), .Y(new_n5825_));
  NOR2X1   g05761(.A(new_n5825_), .B(new_n5822_), .Y(new_n5826_));
  INVX1    g05762(.A(new_n5826_), .Y(new_n5827_));
  XOR2X1   g05763(.A(new_n5825_), .B(new_n5822_), .Y(new_n5828_));
  INVX1    g05764(.A(new_n5828_), .Y(new_n5829_));
  INVX1    g05765(.A(new_n5561_), .Y(new_n5830_));
  XOR2X1   g05766(.A(new_n5607_), .B(new_n5830_), .Y(new_n5831_));
  OAI22X1  g05767(.A0(new_n5096_), .A1(new_n1423_), .B0(new_n4634_), .B1(new_n3669_), .Y(new_n5832_));
  AOI21X1  g05768(.A0(new_n4870_), .A1(new_n1800_), .B0(new_n5832_), .Y(new_n5833_));
  OAI21X1  g05769(.A0(new_n4868_), .A1(new_n3667_), .B0(new_n5833_), .Y(new_n5834_));
  XOR2X1   g05770(.A(new_n5834_), .B(new_n2995_), .Y(new_n5835_));
  NOR2X1   g05771(.A(new_n5835_), .B(new_n5831_), .Y(new_n5836_));
  XOR2X1   g05772(.A(new_n5606_), .B(new_n5605_), .Y(new_n5837_));
  INVX1    g05773(.A(new_n5837_), .Y(new_n5838_));
  OAI22X1  g05774(.A0(new_n5096_), .A1(new_n1465_), .B0(new_n4869_), .B1(new_n3669_), .Y(new_n5839_));
  AOI21X1  g05775(.A0(new_n4635_), .A1(new_n1536_), .B0(new_n5839_), .Y(new_n5840_));
  OAI21X1  g05776(.A0(new_n4868_), .A1(new_n3676_), .B0(new_n5840_), .Y(new_n5841_));
  XOR2X1   g05777(.A(new_n5841_), .B(new_n2995_), .Y(new_n5842_));
  OR2X1    g05778(.A(new_n5842_), .B(new_n5838_), .Y(new_n5843_));
  XOR2X1   g05779(.A(new_n5603_), .B(new_n5579_), .Y(new_n5844_));
  OAI22X1  g05780(.A0(new_n5096_), .A1(new_n3669_), .B0(new_n4634_), .B1(new_n1586_), .Y(new_n5845_));
  AOI21X1  g05781(.A0(new_n4870_), .A1(new_n1536_), .B0(new_n5845_), .Y(new_n5846_));
  OAI21X1  g05782(.A0(new_n4868_), .A1(new_n3478_), .B0(new_n5846_), .Y(new_n5847_));
  XOR2X1   g05783(.A(new_n5847_), .B(\a[8] ), .Y(new_n5848_));
  AOI22X1  g05784(.A0(new_n5097_), .A1(new_n1536_), .B0(new_n4870_), .B1(new_n3480_), .Y(new_n5849_));
  OAI21X1  g05785(.A0(new_n4634_), .A1(new_n1621_), .B0(new_n5849_), .Y(new_n5850_));
  AOI21X1  g05786(.A0(new_n4637_), .A1(new_n3697_), .B0(new_n5850_), .Y(new_n5851_));
  XOR2X1   g05787(.A(new_n5851_), .B(\a[8] ), .Y(new_n5852_));
  INVX1    g05788(.A(new_n5852_), .Y(new_n5853_));
  XOR2X1   g05789(.A(new_n5602_), .B(new_n5601_), .Y(new_n5854_));
  AND2X1   g05790(.A(new_n5854_), .B(new_n5853_), .Y(new_n5855_));
  INVX1    g05791(.A(new_n5855_), .Y(new_n5856_));
  XOR2X1   g05792(.A(new_n5854_), .B(new_n5852_), .Y(new_n5857_));
  INVX1    g05793(.A(new_n5600_), .Y(new_n5858_));
  XOR2X1   g05794(.A(new_n5858_), .B(new_n5596_), .Y(new_n5859_));
  OAI22X1  g05795(.A0(new_n5096_), .A1(new_n1586_), .B0(new_n4634_), .B1(new_n1655_), .Y(new_n5860_));
  AOI21X1  g05796(.A0(new_n4870_), .A1(new_n4538_), .B0(new_n5860_), .Y(new_n5861_));
  OAI21X1  g05797(.A0(new_n4868_), .A1(new_n3719_), .B0(new_n5861_), .Y(new_n5862_));
  XOR2X1   g05798(.A(new_n5862_), .B(new_n2995_), .Y(new_n5863_));
  NOR2X1   g05799(.A(new_n5863_), .B(new_n5859_), .Y(new_n5864_));
  AOI22X1  g05800(.A0(new_n4870_), .A1(new_n3721_), .B0(new_n4635_), .B1(new_n1676_), .Y(new_n5865_));
  OAI21X1  g05801(.A0(new_n5096_), .A1(new_n1621_), .B0(new_n5865_), .Y(new_n5866_));
  AOI21X1  g05802(.A0(new_n4637_), .A1(new_n3745_), .B0(new_n5866_), .Y(new_n5867_));
  XOR2X1   g05803(.A(new_n5867_), .B(\a[8] ), .Y(new_n5868_));
  INVX1    g05804(.A(new_n5590_), .Y(new_n5869_));
  NAND3X1  g05805(.A(new_n5869_), .B(new_n5588_), .C(\a[11] ), .Y(new_n5870_));
  XOR2X1   g05806(.A(new_n5593_), .B(new_n2911_), .Y(new_n5871_));
  AND2X1   g05807(.A(new_n5871_), .B(new_n5870_), .Y(new_n5872_));
  NOR3X1   g05808(.A(new_n5872_), .B(new_n5868_), .C(new_n5594_), .Y(new_n5873_));
  XOR2X1   g05809(.A(new_n5871_), .B(new_n5870_), .Y(new_n5874_));
  XOR2X1   g05810(.A(new_n5874_), .B(new_n5868_), .Y(new_n5875_));
  AOI21X1  g05811(.A0(new_n4079_), .A1(new_n3821_), .B0(new_n2911_), .Y(new_n5876_));
  XOR2X1   g05812(.A(new_n5876_), .B(new_n5589_), .Y(new_n5877_));
  OAI22X1  g05813(.A0(new_n5096_), .A1(new_n1655_), .B0(new_n4869_), .B1(new_n1674_), .Y(new_n5878_));
  AOI21X1  g05814(.A0(new_n4635_), .A1(new_n1706_), .B0(new_n5878_), .Y(new_n5879_));
  OAI21X1  g05815(.A0(new_n4868_), .A1(new_n3773_), .B0(new_n5879_), .Y(new_n5880_));
  XOR2X1   g05816(.A(new_n5880_), .B(new_n2995_), .Y(new_n5881_));
  NOR2X1   g05817(.A(new_n5881_), .B(new_n5877_), .Y(new_n5882_));
  OAI22X1  g05818(.A0(new_n5096_), .A1(new_n1735_), .B0(new_n4869_), .B1(new_n1784_), .Y(new_n5883_));
  AOI21X1  g05819(.A0(new_n4637_), .A1(new_n4165_), .B0(new_n5883_), .Y(new_n5884_));
  XOR2X1   g05820(.A(new_n5884_), .B(\a[8] ), .Y(new_n5885_));
  AND2X1   g05821(.A(new_n4636_), .B(new_n3821_), .Y(new_n5886_));
  OAI22X1  g05822(.A0(new_n4869_), .A1(new_n1735_), .B0(new_n4634_), .B1(new_n1784_), .Y(new_n5887_));
  AOI21X1  g05823(.A0(new_n5097_), .A1(new_n1706_), .B0(new_n5887_), .Y(new_n5888_));
  OAI21X1  g05824(.A0(new_n4868_), .A1(new_n4177_), .B0(new_n5888_), .Y(new_n5889_));
  NOR4X1   g05825(.A(new_n5889_), .B(new_n5886_), .C(new_n5885_), .D(new_n2995_), .Y(new_n5890_));
  NAND2X1  g05826(.A(new_n5890_), .B(new_n5590_), .Y(new_n5891_));
  XOR2X1   g05827(.A(new_n5890_), .B(new_n5869_), .Y(new_n5892_));
  AOI22X1  g05828(.A0(new_n5097_), .A1(new_n1676_), .B0(new_n4635_), .B1(new_n3819_), .Y(new_n5893_));
  OAI21X1  g05829(.A0(new_n4869_), .A1(new_n1708_), .B0(new_n5893_), .Y(new_n5894_));
  AOI21X1  g05830(.A0(new_n4637_), .A1(new_n3829_), .B0(new_n5894_), .Y(new_n5895_));
  XOR2X1   g05831(.A(new_n5895_), .B(\a[8] ), .Y(new_n5896_));
  OAI21X1  g05832(.A0(new_n5896_), .A1(new_n5892_), .B0(new_n5891_), .Y(new_n5897_));
  XOR2X1   g05833(.A(new_n5881_), .B(new_n5877_), .Y(new_n5898_));
  AOI21X1  g05834(.A0(new_n5898_), .A1(new_n5897_), .B0(new_n5882_), .Y(new_n5899_));
  NOR2X1   g05835(.A(new_n5899_), .B(new_n5875_), .Y(new_n5900_));
  OR2X1    g05836(.A(new_n5900_), .B(new_n5873_), .Y(new_n5901_));
  XOR2X1   g05837(.A(new_n5863_), .B(new_n5859_), .Y(new_n5902_));
  AOI21X1  g05838(.A0(new_n5902_), .A1(new_n5901_), .B0(new_n5864_), .Y(new_n5903_));
  OR2X1    g05839(.A(new_n5903_), .B(new_n5857_), .Y(new_n5904_));
  XOR2X1   g05840(.A(new_n5847_), .B(new_n2995_), .Y(new_n5905_));
  XOR2X1   g05841(.A(new_n5905_), .B(new_n5844_), .Y(new_n5906_));
  AOI21X1  g05842(.A0(new_n5904_), .A1(new_n5856_), .B0(new_n5906_), .Y(new_n5907_));
  AOI21X1  g05843(.A0(new_n5848_), .A1(new_n5844_), .B0(new_n5907_), .Y(new_n5908_));
  XOR2X1   g05844(.A(new_n5842_), .B(new_n5837_), .Y(new_n5909_));
  OAI21X1  g05845(.A0(new_n5909_), .A1(new_n5908_), .B0(new_n5843_), .Y(new_n5910_));
  XOR2X1   g05846(.A(new_n5835_), .B(new_n5831_), .Y(new_n5911_));
  AOI21X1  g05847(.A0(new_n5911_), .A1(new_n5910_), .B0(new_n5836_), .Y(new_n5912_));
  OAI21X1  g05848(.A0(new_n5912_), .A1(new_n5829_), .B0(new_n5827_), .Y(new_n5913_));
  AOI21X1  g05849(.A0(new_n5913_), .A1(new_n5818_), .B0(new_n5817_), .Y(new_n5914_));
  OAI21X1  g05850(.A0(new_n5914_), .A1(new_n5810_), .B0(new_n5809_), .Y(new_n5915_));
  XOR2X1   g05851(.A(new_n5801_), .B(new_n5796_), .Y(new_n5916_));
  INVX1    g05852(.A(new_n5916_), .Y(new_n5917_));
  AOI21X1  g05853(.A0(new_n5917_), .A1(new_n5915_), .B0(new_n5802_), .Y(new_n5918_));
  XOR2X1   g05854(.A(new_n5794_), .B(new_n5789_), .Y(new_n5919_));
  OAI21X1  g05855(.A0(new_n5919_), .A1(new_n5918_), .B0(new_n5795_), .Y(new_n5920_));
  XOR2X1   g05856(.A(new_n5787_), .B(new_n5783_), .Y(new_n5921_));
  AOI21X1  g05857(.A0(new_n5921_), .A1(new_n5920_), .B0(new_n5788_), .Y(new_n5922_));
  OAI21X1  g05858(.A0(new_n5922_), .A1(new_n5781_), .B0(new_n5779_), .Y(new_n5923_));
  AOI21X1  g05859(.A0(new_n5923_), .A1(new_n5771_), .B0(new_n5770_), .Y(new_n5924_));
  OAI21X1  g05860(.A0(new_n5924_), .A1(new_n5764_), .B0(new_n5763_), .Y(new_n5925_));
  XOR2X1   g05861(.A(new_n5755_), .B(new_n5750_), .Y(new_n5926_));
  INVX1    g05862(.A(new_n5926_), .Y(new_n5927_));
  AOI21X1  g05863(.A0(new_n5927_), .A1(new_n5925_), .B0(new_n5756_), .Y(new_n5928_));
  XOR2X1   g05864(.A(new_n5748_), .B(new_n5743_), .Y(new_n5929_));
  OAI21X1  g05865(.A0(new_n5929_), .A1(new_n5928_), .B0(new_n5749_), .Y(new_n5930_));
  XOR2X1   g05866(.A(new_n5741_), .B(new_n5737_), .Y(new_n5931_));
  AOI21X1  g05867(.A0(new_n5931_), .A1(new_n5930_), .B0(new_n5742_), .Y(new_n5932_));
  OAI21X1  g05868(.A0(new_n5932_), .A1(new_n5735_), .B0(new_n5733_), .Y(new_n5933_));
  AOI21X1  g05869(.A0(new_n5933_), .A1(new_n5726_), .B0(new_n5723_), .Y(new_n5934_));
  XOR2X1   g05870(.A(new_n5716_), .B(new_n2995_), .Y(new_n5935_));
  XOR2X1   g05871(.A(new_n5935_), .B(new_n5713_), .Y(new_n5936_));
  NOR2X1   g05872(.A(new_n5936_), .B(new_n5934_), .Y(new_n5937_));
  AOI21X1  g05873(.A0(new_n5717_), .A1(new_n5713_), .B0(new_n5937_), .Y(new_n5938_));
  XOR2X1   g05874(.A(new_n5710_), .B(new_n5705_), .Y(new_n5939_));
  OR2X1    g05875(.A(new_n5939_), .B(new_n5938_), .Y(new_n5940_));
  XOR2X1   g05876(.A(new_n5702_), .B(new_n2995_), .Y(new_n5941_));
  XOR2X1   g05877(.A(new_n5941_), .B(new_n5699_), .Y(new_n5942_));
  AOI21X1  g05878(.A0(new_n5940_), .A1(new_n5712_), .B0(new_n5942_), .Y(new_n5943_));
  XOR2X1   g05879(.A(new_n5695_), .B(new_n5691_), .Y(new_n5944_));
  OAI21X1  g05880(.A0(new_n5943_), .A1(new_n5704_), .B0(new_n5944_), .Y(new_n5945_));
  AND2X1   g05881(.A(new_n5945_), .B(new_n5697_), .Y(new_n5946_));
  XOR2X1   g05882(.A(new_n5689_), .B(\a[8] ), .Y(new_n5947_));
  XOR2X1   g05883(.A(new_n5947_), .B(new_n5686_), .Y(new_n5948_));
  NOR2X1   g05884(.A(new_n5948_), .B(new_n5946_), .Y(new_n5949_));
  AOI21X1  g05885(.A0(new_n5690_), .A1(new_n5686_), .B0(new_n5949_), .Y(new_n5950_));
  XOR2X1   g05886(.A(new_n5684_), .B(new_n5679_), .Y(new_n5951_));
  OAI21X1  g05887(.A0(new_n5951_), .A1(new_n5950_), .B0(new_n5685_), .Y(new_n5952_));
  XOR2X1   g05888(.A(new_n5676_), .B(new_n5672_), .Y(new_n5953_));
  AND2X1   g05889(.A(new_n5953_), .B(new_n5952_), .Y(new_n5954_));
  XOR2X1   g05890(.A(new_n5654_), .B(new_n5653_), .Y(new_n5955_));
  OAI21X1  g05891(.A0(new_n5954_), .A1(new_n5677_), .B0(new_n5955_), .Y(new_n5956_));
  INVX1    g05892(.A(new_n2757_), .Y(new_n5957_));
  INVX1    g05893(.A(new_n65_), .Y(new_n5958_));
  NAND2X1  g05894(.A(new_n66_), .B(new_n5958_), .Y(new_n5959_));
  INVX1    g05895(.A(new_n5959_), .Y(new_n5960_));
  AOI22X1  g05896(.A0(new_n5960_), .A1(new_n2649_), .B0(new_n5659_), .B1(new_n2421_), .Y(new_n5961_));
  OAI21X1  g05897(.A0(new_n5372_), .A1(new_n2379_), .B0(new_n5961_), .Y(new_n5962_));
  AOI21X1  g05898(.A0(new_n5957_), .A1(new_n67_), .B0(new_n5962_), .Y(new_n5963_));
  XOR2X1   g05899(.A(new_n5963_), .B(\a[5] ), .Y(new_n5964_));
  AOI21X1  g05900(.A0(new_n5953_), .A1(new_n5952_), .B0(new_n5677_), .Y(new_n5965_));
  XOR2X1   g05901(.A(new_n5955_), .B(new_n5965_), .Y(new_n5966_));
  OAI21X1  g05902(.A0(new_n5966_), .A1(new_n5964_), .B0(new_n5956_), .Y(new_n5967_));
  XOR2X1   g05903(.A(new_n5665_), .B(new_n5664_), .Y(new_n5968_));
  AND2X1   g05904(.A(new_n5968_), .B(new_n5967_), .Y(new_n5969_));
  NOR3X1   g05905(.A(new_n3431_), .B(\a[1] ), .C(\a[0] ), .Y(new_n5970_));
  XOR2X1   g05906(.A(\a[2] ), .B(\a[1] ), .Y(new_n5971_));
  AND2X1   g05907(.A(new_n5971_), .B(\a[0] ), .Y(new_n5972_));
  AOI22X1  g05908(.A0(new_n5972_), .A1(new_n2652_), .B0(new_n5970_), .B1(new_n2649_), .Y(new_n5973_));
  XOR2X1   g05909(.A(new_n5973_), .B(\a[2] ), .Y(new_n5974_));
  AOI22X1  g05910(.A0(new_n5960_), .A1(new_n2421_), .B0(new_n5373_), .B1(new_n2420_), .Y(new_n5975_));
  OAI21X1  g05911(.A0(new_n5658_), .A1(new_n2379_), .B0(new_n5975_), .Y(new_n5976_));
  AOI21X1  g05912(.A0(new_n2416_), .A1(new_n67_), .B0(new_n5976_), .Y(new_n5977_));
  XOR2X1   g05913(.A(new_n5977_), .B(\a[5] ), .Y(new_n5978_));
  NOR2X1   g05914(.A(new_n5978_), .B(new_n5974_), .Y(new_n5979_));
  XOR2X1   g05915(.A(new_n5978_), .B(new_n5974_), .Y(new_n5980_));
  XOR2X1   g05916(.A(new_n5953_), .B(new_n5952_), .Y(new_n5981_));
  AOI21X1  g05917(.A0(new_n5981_), .A1(new_n5980_), .B0(new_n5979_), .Y(new_n5982_));
  INVX1    g05918(.A(new_n5982_), .Y(new_n5983_));
  XOR2X1   g05919(.A(new_n5966_), .B(new_n5964_), .Y(new_n5984_));
  AND2X1   g05920(.A(new_n5984_), .B(new_n5983_), .Y(new_n5985_));
  INVX1    g05921(.A(new_n5985_), .Y(new_n5986_));
  XOR2X1   g05922(.A(new_n5981_), .B(new_n5980_), .Y(new_n5987_));
  INVX1    g05923(.A(new_n5987_), .Y(new_n5988_));
  AOI22X1  g05924(.A0(new_n5659_), .A1(new_n2420_), .B0(new_n5373_), .B1(new_n2627_), .Y(new_n5989_));
  OAI21X1  g05925(.A0(new_n5959_), .A1(new_n2379_), .B0(new_n5989_), .Y(new_n5990_));
  AOI21X1  g05926(.A0(new_n2625_), .A1(new_n67_), .B0(new_n5990_), .Y(new_n5991_));
  XOR2X1   g05927(.A(new_n5991_), .B(\a[5] ), .Y(new_n5992_));
  INVX1    g05928(.A(new_n5992_), .Y(new_n5993_));
  XOR2X1   g05929(.A(new_n5951_), .B(new_n5950_), .Y(new_n5994_));
  XOR2X1   g05930(.A(new_n5994_), .B(new_n5992_), .Y(new_n5995_));
  AOI22X1  g05931(.A0(new_n5960_), .A1(new_n2420_), .B0(new_n5373_), .B1(new_n2252_), .Y(new_n5996_));
  OAI21X1  g05932(.A0(new_n5658_), .A1(new_n2287_), .B0(new_n5996_), .Y(new_n5997_));
  AOI21X1  g05933(.A0(new_n2669_), .A1(new_n67_), .B0(new_n5997_), .Y(new_n5998_));
  XOR2X1   g05934(.A(new_n5998_), .B(\a[5] ), .Y(new_n5999_));
  INVX1    g05935(.A(new_n5948_), .Y(new_n6000_));
  XOR2X1   g05936(.A(new_n6000_), .B(new_n5946_), .Y(new_n6001_));
  NOR2X1   g05937(.A(new_n6001_), .B(new_n5999_), .Y(new_n6002_));
  XOR2X1   g05938(.A(new_n6001_), .B(new_n5999_), .Y(new_n6003_));
  AOI22X1  g05939(.A0(new_n5960_), .A1(new_n2627_), .B0(new_n5373_), .B1(new_n2093_), .Y(new_n6004_));
  OAI21X1  g05940(.A0(new_n5658_), .A1(new_n2137_), .B0(new_n6004_), .Y(new_n6005_));
  AOI21X1  g05941(.A0(new_n2294_), .A1(new_n67_), .B0(new_n6005_), .Y(new_n6006_));
  XOR2X1   g05942(.A(new_n6006_), .B(\a[5] ), .Y(new_n6007_));
  NOR2X1   g05943(.A(new_n5943_), .B(new_n5704_), .Y(new_n6008_));
  XOR2X1   g05944(.A(new_n5944_), .B(new_n6008_), .Y(new_n6009_));
  XOR2X1   g05945(.A(new_n6009_), .B(new_n6007_), .Y(new_n6010_));
  INVX1    g05946(.A(new_n6010_), .Y(new_n6011_));
  AOI22X1  g05947(.A0(new_n5960_), .A1(new_n2252_), .B0(new_n5373_), .B1(new_n2246_), .Y(new_n6012_));
  OAI21X1  g05948(.A0(new_n5658_), .A1(new_n2092_), .B0(new_n6012_), .Y(new_n6013_));
  AOI21X1  g05949(.A0(new_n2201_), .A1(new_n67_), .B0(new_n6013_), .Y(new_n6014_));
  XOR2X1   g05950(.A(new_n6014_), .B(\a[5] ), .Y(new_n6015_));
  AND2X1   g05951(.A(new_n5940_), .B(new_n5712_), .Y(new_n6016_));
  INVX1    g05952(.A(new_n5942_), .Y(new_n6017_));
  XOR2X1   g05953(.A(new_n6017_), .B(new_n6016_), .Y(new_n6018_));
  NOR2X1   g05954(.A(new_n6018_), .B(new_n6015_), .Y(new_n6019_));
  XOR2X1   g05955(.A(new_n6018_), .B(new_n6015_), .Y(new_n6020_));
  AOI22X1  g05956(.A0(new_n5960_), .A1(new_n2093_), .B0(new_n5373_), .B1(new_n1887_), .Y(new_n6021_));
  OAI21X1  g05957(.A0(new_n5658_), .A1(new_n2183_), .B0(new_n6021_), .Y(new_n6022_));
  AOI21X1  g05958(.A0(new_n2430_), .A1(new_n67_), .B0(new_n6022_), .Y(new_n6023_));
  XOR2X1   g05959(.A(new_n6023_), .B(\a[5] ), .Y(new_n6024_));
  INVX1    g05960(.A(new_n5939_), .Y(new_n6025_));
  XOR2X1   g05961(.A(new_n6025_), .B(new_n5938_), .Y(new_n6026_));
  XOR2X1   g05962(.A(new_n6026_), .B(new_n6024_), .Y(new_n6027_));
  INVX1    g05963(.A(new_n6027_), .Y(new_n6028_));
  AOI22X1  g05964(.A0(new_n5960_), .A1(new_n2246_), .B0(new_n5373_), .B1(new_n2048_), .Y(new_n6029_));
  OAI21X1  g05965(.A0(new_n5658_), .A1(new_n1879_), .B0(new_n6029_), .Y(new_n6030_));
  AOI21X1  g05966(.A0(new_n2244_), .A1(new_n67_), .B0(new_n6030_), .Y(new_n6031_));
  XOR2X1   g05967(.A(new_n6031_), .B(\a[5] ), .Y(new_n6032_));
  INVX1    g05968(.A(new_n5934_), .Y(new_n6033_));
  XOR2X1   g05969(.A(new_n5936_), .B(new_n6033_), .Y(new_n6034_));
  NOR2X1   g05970(.A(new_n6034_), .B(new_n6032_), .Y(new_n6035_));
  XOR2X1   g05971(.A(new_n6034_), .B(new_n6032_), .Y(new_n6036_));
  XOR2X1   g05972(.A(new_n5933_), .B(new_n5726_), .Y(new_n6037_));
  INVX1    g05973(.A(new_n6037_), .Y(new_n6038_));
  OAI22X1  g05974(.A0(new_n5959_), .A1(new_n1879_), .B0(new_n5372_), .B1(new_n623_), .Y(new_n6039_));
  AOI21X1  g05975(.A0(new_n5659_), .A1(new_n2048_), .B0(new_n6039_), .Y(new_n6040_));
  OAI21X1  g05976(.A0(new_n1881_), .A1(new_n5657_), .B0(new_n6040_), .Y(new_n6041_));
  XOR2X1   g05977(.A(new_n6041_), .B(new_n3289_), .Y(new_n6042_));
  NOR2X1   g05978(.A(new_n6042_), .B(new_n6038_), .Y(new_n6043_));
  XOR2X1   g05979(.A(new_n5932_), .B(new_n5735_), .Y(new_n6044_));
  INVX1    g05980(.A(new_n6044_), .Y(new_n6045_));
  OAI22X1  g05981(.A0(new_n5959_), .A1(new_n520_), .B0(new_n5372_), .B1(new_n690_), .Y(new_n6046_));
  AOI21X1  g05982(.A0(new_n5659_), .A1(new_n1886_), .B0(new_n6046_), .Y(new_n6047_));
  OAI21X1  g05983(.A0(new_n3114_), .A1(new_n5657_), .B0(new_n6047_), .Y(new_n6048_));
  XOR2X1   g05984(.A(new_n6048_), .B(new_n3289_), .Y(new_n6049_));
  NOR2X1   g05985(.A(new_n6049_), .B(new_n6045_), .Y(new_n6050_));
  INVX1    g05986(.A(new_n6050_), .Y(new_n6051_));
  AOI22X1  g05987(.A0(new_n5960_), .A1(new_n1886_), .B0(new_n5373_), .B1(new_n2036_), .Y(new_n6052_));
  OAI21X1  g05988(.A0(new_n5658_), .A1(new_n690_), .B0(new_n6052_), .Y(new_n6053_));
  AOI21X1  g05989(.A0(new_n2035_), .A1(new_n67_), .B0(new_n6053_), .Y(new_n6054_));
  XOR2X1   g05990(.A(new_n6054_), .B(\a[5] ), .Y(new_n6055_));
  INVX1    g05991(.A(new_n6055_), .Y(new_n6056_));
  XOR2X1   g05992(.A(new_n5931_), .B(new_n5930_), .Y(new_n6057_));
  XOR2X1   g05993(.A(new_n6057_), .B(new_n6055_), .Y(new_n6058_));
  AOI22X1  g05994(.A0(new_n5960_), .A1(new_n2049_), .B0(new_n5373_), .B1(new_n2481_), .Y(new_n6059_));
  OAI21X1  g05995(.A0(new_n5658_), .A1(new_n783_), .B0(new_n6059_), .Y(new_n6060_));
  AOI21X1  g05996(.A0(new_n2480_), .A1(new_n67_), .B0(new_n6060_), .Y(new_n6061_));
  XOR2X1   g05997(.A(new_n6061_), .B(\a[5] ), .Y(new_n6062_));
  INVX1    g05998(.A(new_n5929_), .Y(new_n6063_));
  XOR2X1   g05999(.A(new_n6063_), .B(new_n5928_), .Y(new_n6064_));
  NOR2X1   g06000(.A(new_n6064_), .B(new_n6062_), .Y(new_n6065_));
  XOR2X1   g06001(.A(new_n6064_), .B(new_n6062_), .Y(new_n6066_));
  AOI22X1  g06002(.A0(new_n5960_), .A1(new_n2036_), .B0(new_n5373_), .B1(new_n2602_), .Y(new_n6067_));
  OAI21X1  g06003(.A0(new_n5658_), .A1(new_n847_), .B0(new_n6067_), .Y(new_n6068_));
  AOI21X1  g06004(.A0(new_n2494_), .A1(new_n67_), .B0(new_n6068_), .Y(new_n6069_));
  XOR2X1   g06005(.A(new_n6069_), .B(\a[5] ), .Y(new_n6070_));
  XOR2X1   g06006(.A(new_n5926_), .B(new_n5925_), .Y(new_n6071_));
  NOR2X1   g06007(.A(new_n6071_), .B(new_n6070_), .Y(new_n6072_));
  INVX1    g06008(.A(new_n6072_), .Y(new_n6073_));
  XOR2X1   g06009(.A(new_n6071_), .B(new_n6070_), .Y(new_n6074_));
  INVX1    g06010(.A(new_n6074_), .Y(new_n6075_));
  INVX1    g06011(.A(new_n5764_), .Y(new_n6076_));
  XOR2X1   g06012(.A(new_n5924_), .B(new_n6076_), .Y(new_n6077_));
  OAI22X1  g06013(.A0(new_n5959_), .A1(new_n847_), .B0(new_n5372_), .B1(new_n957_), .Y(new_n6078_));
  AOI21X1  g06014(.A0(new_n5659_), .A1(new_n2602_), .B0(new_n6078_), .Y(new_n6079_));
  OAI21X1  g06015(.A0(new_n2708_), .A1(new_n5657_), .B0(new_n6079_), .Y(new_n6080_));
  XOR2X1   g06016(.A(new_n6080_), .B(new_n3289_), .Y(new_n6081_));
  NOR2X1   g06017(.A(new_n6081_), .B(new_n6077_), .Y(new_n6082_));
  XOR2X1   g06018(.A(new_n5923_), .B(new_n5771_), .Y(new_n6083_));
  INVX1    g06019(.A(new_n6083_), .Y(new_n6084_));
  OAI22X1  g06020(.A0(new_n5959_), .A1(new_n903_), .B0(new_n5372_), .B1(new_n985_), .Y(new_n6085_));
  AOI21X1  g06021(.A0(new_n5659_), .A1(new_n2835_), .B0(new_n6085_), .Y(new_n6086_));
  OAI21X1  g06022(.A0(new_n2600_), .A1(new_n5657_), .B0(new_n6086_), .Y(new_n6087_));
  XOR2X1   g06023(.A(new_n6087_), .B(new_n3289_), .Y(new_n6088_));
  NOR2X1   g06024(.A(new_n6088_), .B(new_n6084_), .Y(new_n6089_));
  XOR2X1   g06025(.A(new_n5922_), .B(new_n5781_), .Y(new_n6090_));
  INVX1    g06026(.A(new_n6090_), .Y(new_n6091_));
  OAI22X1  g06027(.A0(new_n5959_), .A1(new_n957_), .B0(new_n5658_), .B1(new_n985_), .Y(new_n6092_));
  AOI21X1  g06028(.A0(new_n5373_), .A1(new_n1822_), .B0(new_n6092_), .Y(new_n6093_));
  OAI21X1  g06029(.A0(new_n2833_), .A1(new_n5657_), .B0(new_n6093_), .Y(new_n6094_));
  XOR2X1   g06030(.A(new_n6094_), .B(new_n3289_), .Y(new_n6095_));
  AOI22X1  g06031(.A0(new_n5960_), .A1(new_n2603_), .B0(new_n5373_), .B1(new_n1126_), .Y(new_n6096_));
  OAI21X1  g06032(.A0(new_n5658_), .A1(new_n1065_), .B0(new_n6096_), .Y(new_n6097_));
  AOI21X1  g06033(.A0(new_n2824_), .A1(new_n67_), .B0(new_n6097_), .Y(new_n6098_));
  XOR2X1   g06034(.A(new_n6098_), .B(\a[5] ), .Y(new_n6099_));
  INVX1    g06035(.A(new_n6099_), .Y(new_n6100_));
  XOR2X1   g06036(.A(new_n5921_), .B(new_n5920_), .Y(new_n6101_));
  AND2X1   g06037(.A(new_n6101_), .B(new_n6100_), .Y(new_n6102_));
  XOR2X1   g06038(.A(new_n6101_), .B(new_n6099_), .Y(new_n6103_));
  AOI22X1  g06039(.A0(new_n5960_), .A1(new_n1822_), .B0(new_n5659_), .B1(new_n1126_), .Y(new_n6104_));
  OAI21X1  g06040(.A0(new_n5372_), .A1(new_n1189_), .B0(new_n6104_), .Y(new_n6105_));
  AOI21X1  g06041(.A0(new_n2963_), .A1(new_n67_), .B0(new_n6105_), .Y(new_n6106_));
  XOR2X1   g06042(.A(new_n6106_), .B(\a[5] ), .Y(new_n6107_));
  INVX1    g06043(.A(new_n5919_), .Y(new_n6108_));
  XOR2X1   g06044(.A(new_n6108_), .B(new_n5918_), .Y(new_n6109_));
  NOR2X1   g06045(.A(new_n6109_), .B(new_n6107_), .Y(new_n6110_));
  XOR2X1   g06046(.A(new_n6109_), .B(new_n6107_), .Y(new_n6111_));
  AOI22X1  g06047(.A0(new_n5960_), .A1(new_n1126_), .B0(new_n5373_), .B1(new_n2977_), .Y(new_n6112_));
  OAI21X1  g06048(.A0(new_n5658_), .A1(new_n1189_), .B0(new_n6112_), .Y(new_n6113_));
  AOI21X1  g06049(.A0(new_n2976_), .A1(new_n67_), .B0(new_n6113_), .Y(new_n6114_));
  XOR2X1   g06050(.A(new_n6114_), .B(\a[5] ), .Y(new_n6115_));
  XOR2X1   g06051(.A(new_n5916_), .B(new_n5915_), .Y(new_n6116_));
  XOR2X1   g06052(.A(new_n6116_), .B(new_n6115_), .Y(new_n6117_));
  INVX1    g06053(.A(new_n6117_), .Y(new_n6118_));
  INVX1    g06054(.A(new_n5810_), .Y(new_n6119_));
  XOR2X1   g06055(.A(new_n5914_), .B(new_n6119_), .Y(new_n6120_));
  OAI22X1  g06056(.A0(new_n5959_), .A1(new_n1189_), .B0(new_n5658_), .B1(new_n1236_), .Y(new_n6121_));
  AOI21X1  g06057(.A0(new_n5373_), .A1(new_n3342_), .B0(new_n6121_), .Y(new_n6122_));
  OAI21X1  g06058(.A0(new_n3180_), .A1(new_n5657_), .B0(new_n6122_), .Y(new_n6123_));
  XOR2X1   g06059(.A(new_n6123_), .B(new_n3289_), .Y(new_n6124_));
  NOR2X1   g06060(.A(new_n6124_), .B(new_n6120_), .Y(new_n6125_));
  XOR2X1   g06061(.A(new_n5913_), .B(new_n5818_), .Y(new_n6126_));
  INVX1    g06062(.A(new_n6126_), .Y(new_n6127_));
  OAI22X1  g06063(.A0(new_n5959_), .A1(new_n1236_), .B0(new_n5372_), .B1(new_n1339_), .Y(new_n6128_));
  AOI21X1  g06064(.A0(new_n5659_), .A1(new_n3342_), .B0(new_n6128_), .Y(new_n6129_));
  OAI21X1  g06065(.A0(new_n3053_), .A1(new_n5657_), .B0(new_n6129_), .Y(new_n6130_));
  XOR2X1   g06066(.A(new_n6130_), .B(new_n3289_), .Y(new_n6131_));
  NOR2X1   g06067(.A(new_n6131_), .B(new_n6127_), .Y(new_n6132_));
  XOR2X1   g06068(.A(new_n5912_), .B(new_n5829_), .Y(new_n6133_));
  INVX1    g06069(.A(new_n6133_), .Y(new_n6134_));
  OAI22X1  g06070(.A0(new_n5959_), .A1(new_n1294_), .B0(new_n5372_), .B1(new_n1358_), .Y(new_n6135_));
  AOI21X1  g06071(.A0(new_n5659_), .A1(new_n3055_), .B0(new_n6135_), .Y(new_n6136_));
  OAI21X1  g06072(.A0(new_n3340_), .A1(new_n5657_), .B0(new_n6136_), .Y(new_n6137_));
  XOR2X1   g06073(.A(new_n6137_), .B(new_n3289_), .Y(new_n6138_));
  NOR2X1   g06074(.A(new_n6138_), .B(new_n6134_), .Y(new_n6139_));
  AOI22X1  g06075(.A0(new_n5960_), .A1(new_n3055_), .B0(new_n5659_), .B1(new_n1357_), .Y(new_n6140_));
  OAI21X1  g06076(.A0(new_n5372_), .A1(new_n1389_), .B0(new_n6140_), .Y(new_n6141_));
  AOI21X1  g06077(.A0(new_n3425_), .A1(new_n67_), .B0(new_n6141_), .Y(new_n6142_));
  XOR2X1   g06078(.A(new_n6142_), .B(\a[5] ), .Y(new_n6143_));
  INVX1    g06079(.A(new_n6143_), .Y(new_n6144_));
  XOR2X1   g06080(.A(new_n5911_), .B(new_n5910_), .Y(new_n6145_));
  NAND2X1  g06081(.A(new_n6145_), .B(new_n6144_), .Y(new_n6146_));
  XOR2X1   g06082(.A(new_n6145_), .B(new_n6143_), .Y(new_n6147_));
  AOI22X1  g06083(.A0(new_n5960_), .A1(new_n1357_), .B0(new_n5373_), .B1(new_n3327_), .Y(new_n6148_));
  OAI21X1  g06084(.A0(new_n5658_), .A1(new_n1389_), .B0(new_n6148_), .Y(new_n6149_));
  AOI21X1  g06085(.A0(new_n3326_), .A1(new_n67_), .B0(new_n6149_), .Y(new_n6150_));
  XOR2X1   g06086(.A(new_n6150_), .B(\a[5] ), .Y(new_n6151_));
  INVX1    g06087(.A(new_n5909_), .Y(new_n6152_));
  XOR2X1   g06088(.A(new_n6152_), .B(new_n5908_), .Y(new_n6153_));
  NOR2X1   g06089(.A(new_n6153_), .B(new_n6151_), .Y(new_n6154_));
  XOR2X1   g06090(.A(new_n6153_), .B(new_n6151_), .Y(new_n6155_));
  AOI22X1  g06091(.A0(new_n5659_), .A1(new_n3327_), .B0(new_n5373_), .B1(new_n1800_), .Y(new_n6156_));
  OAI21X1  g06092(.A0(new_n5959_), .A1(new_n1389_), .B0(new_n6156_), .Y(new_n6157_));
  AOI21X1  g06093(.A0(new_n3497_), .A1(new_n67_), .B0(new_n6157_), .Y(new_n6158_));
  XOR2X1   g06094(.A(new_n6158_), .B(\a[5] ), .Y(new_n6159_));
  AND2X1   g06095(.A(new_n5904_), .B(new_n5856_), .Y(new_n6160_));
  INVX1    g06096(.A(new_n5906_), .Y(new_n6161_));
  XOR2X1   g06097(.A(new_n6161_), .B(new_n6160_), .Y(new_n6162_));
  NOR2X1   g06098(.A(new_n6162_), .B(new_n6159_), .Y(new_n6163_));
  INVX1    g06099(.A(new_n6163_), .Y(new_n6164_));
  XOR2X1   g06100(.A(new_n6162_), .B(new_n6159_), .Y(new_n6165_));
  INVX1    g06101(.A(new_n6165_), .Y(new_n6166_));
  XOR2X1   g06102(.A(new_n5903_), .B(new_n5857_), .Y(new_n6167_));
  INVX1    g06103(.A(new_n6167_), .Y(new_n6168_));
  OAI22X1  g06104(.A0(new_n5959_), .A1(new_n1423_), .B0(new_n5372_), .B1(new_n3669_), .Y(new_n6169_));
  AOI21X1  g06105(.A0(new_n5659_), .A1(new_n1800_), .B0(new_n6169_), .Y(new_n6170_));
  OAI21X1  g06106(.A0(new_n3667_), .A1(new_n5657_), .B0(new_n6170_), .Y(new_n6171_));
  XOR2X1   g06107(.A(new_n6171_), .B(new_n3289_), .Y(new_n6172_));
  NOR2X1   g06108(.A(new_n6172_), .B(new_n6168_), .Y(new_n6173_));
  XOR2X1   g06109(.A(new_n5902_), .B(new_n5901_), .Y(new_n6174_));
  OAI22X1  g06110(.A0(new_n5959_), .A1(new_n1465_), .B0(new_n5658_), .B1(new_n3669_), .Y(new_n6175_));
  AOI21X1  g06111(.A0(new_n5373_), .A1(new_n1536_), .B0(new_n6175_), .Y(new_n6176_));
  OAI21X1  g06112(.A0(new_n3676_), .A1(new_n5657_), .B0(new_n6176_), .Y(new_n6177_));
  XOR2X1   g06113(.A(new_n6177_), .B(\a[5] ), .Y(new_n6178_));
  NAND2X1  g06114(.A(new_n6178_), .B(new_n6174_), .Y(new_n6179_));
  XOR2X1   g06115(.A(new_n5899_), .B(new_n5875_), .Y(new_n6180_));
  INVX1    g06116(.A(new_n6180_), .Y(new_n6181_));
  OAI22X1  g06117(.A0(new_n5959_), .A1(new_n3669_), .B0(new_n5372_), .B1(new_n1586_), .Y(new_n6182_));
  AOI21X1  g06118(.A0(new_n5659_), .A1(new_n1536_), .B0(new_n6182_), .Y(new_n6183_));
  OAI21X1  g06119(.A0(new_n3478_), .A1(new_n5657_), .B0(new_n6183_), .Y(new_n6184_));
  XOR2X1   g06120(.A(new_n6184_), .B(new_n3289_), .Y(new_n6185_));
  NOR2X1   g06121(.A(new_n6185_), .B(new_n6181_), .Y(new_n6186_));
  AOI22X1  g06122(.A0(new_n5960_), .A1(new_n1536_), .B0(new_n5659_), .B1(new_n3480_), .Y(new_n6187_));
  OAI21X1  g06123(.A0(new_n5372_), .A1(new_n1621_), .B0(new_n6187_), .Y(new_n6188_));
  AOI21X1  g06124(.A0(new_n3697_), .A1(new_n67_), .B0(new_n6188_), .Y(new_n6189_));
  XOR2X1   g06125(.A(new_n6189_), .B(\a[5] ), .Y(new_n6190_));
  INVX1    g06126(.A(new_n6190_), .Y(new_n6191_));
  XOR2X1   g06127(.A(new_n5898_), .B(new_n5897_), .Y(new_n6192_));
  NAND2X1  g06128(.A(new_n6192_), .B(new_n6191_), .Y(new_n6193_));
  XOR2X1   g06129(.A(new_n6192_), .B(new_n6190_), .Y(new_n6194_));
  XOR2X1   g06130(.A(new_n5896_), .B(new_n5892_), .Y(new_n6195_));
  INVX1    g06131(.A(new_n6195_), .Y(new_n6196_));
  OAI22X1  g06132(.A0(new_n5959_), .A1(new_n1586_), .B0(new_n5372_), .B1(new_n1655_), .Y(new_n6197_));
  AOI21X1  g06133(.A0(new_n5659_), .A1(new_n4538_), .B0(new_n6197_), .Y(new_n6198_));
  OAI21X1  g06134(.A0(new_n3719_), .A1(new_n5657_), .B0(new_n6198_), .Y(new_n6199_));
  XOR2X1   g06135(.A(new_n6199_), .B(new_n3289_), .Y(new_n6200_));
  NOR2X1   g06136(.A(new_n6200_), .B(new_n6196_), .Y(new_n6201_));
  AOI22X1  g06137(.A0(new_n5659_), .A1(new_n3721_), .B0(new_n5373_), .B1(new_n1676_), .Y(new_n6202_));
  OAI21X1  g06138(.A0(new_n5959_), .A1(new_n1621_), .B0(new_n6202_), .Y(new_n6203_));
  AOI21X1  g06139(.A0(new_n3745_), .A1(new_n67_), .B0(new_n6203_), .Y(new_n6204_));
  XOR2X1   g06140(.A(new_n6204_), .B(\a[5] ), .Y(new_n6205_));
  INVX1    g06141(.A(new_n6205_), .Y(new_n6206_));
  INVX1    g06142(.A(new_n5886_), .Y(new_n6207_));
  NAND3X1  g06143(.A(new_n6207_), .B(new_n5884_), .C(\a[8] ), .Y(new_n6208_));
  XOR2X1   g06144(.A(new_n5889_), .B(new_n2995_), .Y(new_n6209_));
  XOR2X1   g06145(.A(new_n6209_), .B(new_n6208_), .Y(new_n6210_));
  NAND2X1  g06146(.A(new_n6210_), .B(new_n6206_), .Y(new_n6211_));
  XOR2X1   g06147(.A(new_n6210_), .B(new_n6205_), .Y(new_n6212_));
  AOI21X1  g06148(.A0(new_n4636_), .A1(new_n3821_), .B0(new_n2995_), .Y(new_n6213_));
  XOR2X1   g06149(.A(new_n6213_), .B(new_n5885_), .Y(new_n6214_));
  OAI22X1  g06150(.A0(new_n5959_), .A1(new_n1655_), .B0(new_n5658_), .B1(new_n1674_), .Y(new_n6215_));
  AOI21X1  g06151(.A0(new_n5373_), .A1(new_n1706_), .B0(new_n6215_), .Y(new_n6216_));
  OAI21X1  g06152(.A0(new_n3773_), .A1(new_n5657_), .B0(new_n6216_), .Y(new_n6217_));
  XOR2X1   g06153(.A(new_n6217_), .B(new_n3289_), .Y(new_n6218_));
  NOR2X1   g06154(.A(new_n6218_), .B(new_n6214_), .Y(new_n6219_));
  OAI22X1  g06155(.A0(new_n5959_), .A1(new_n1735_), .B0(new_n5658_), .B1(new_n1784_), .Y(new_n6220_));
  AOI21X1  g06156(.A0(new_n4165_), .A1(new_n67_), .B0(new_n6220_), .Y(new_n6221_));
  XOR2X1   g06157(.A(new_n6221_), .B(\a[5] ), .Y(new_n6222_));
  AND2X1   g06158(.A(new_n3821_), .B(new_n66_), .Y(new_n6223_));
  OAI22X1  g06159(.A0(new_n5658_), .A1(new_n1735_), .B0(new_n5372_), .B1(new_n1784_), .Y(new_n6224_));
  AOI21X1  g06160(.A0(new_n5960_), .A1(new_n1706_), .B0(new_n6224_), .Y(new_n6225_));
  OAI21X1  g06161(.A0(new_n4177_), .A1(new_n5657_), .B0(new_n6225_), .Y(new_n6226_));
  NOR4X1   g06162(.A(new_n6226_), .B(new_n6223_), .C(new_n6222_), .D(new_n3289_), .Y(new_n6227_));
  NAND2X1  g06163(.A(new_n6227_), .B(new_n5886_), .Y(new_n6228_));
  XOR2X1   g06164(.A(new_n6227_), .B(new_n6207_), .Y(new_n6229_));
  AOI22X1  g06165(.A0(new_n5960_), .A1(new_n1676_), .B0(new_n5373_), .B1(new_n3819_), .Y(new_n6230_));
  OAI21X1  g06166(.A0(new_n5658_), .A1(new_n1708_), .B0(new_n6230_), .Y(new_n6231_));
  AOI21X1  g06167(.A0(new_n3829_), .A1(new_n67_), .B0(new_n6231_), .Y(new_n6232_));
  XOR2X1   g06168(.A(new_n6232_), .B(\a[5] ), .Y(new_n6233_));
  OAI21X1  g06169(.A0(new_n6233_), .A1(new_n6229_), .B0(new_n6228_), .Y(new_n6234_));
  XOR2X1   g06170(.A(new_n6218_), .B(new_n6214_), .Y(new_n6235_));
  AOI21X1  g06171(.A0(new_n6235_), .A1(new_n6234_), .B0(new_n6219_), .Y(new_n6236_));
  OAI21X1  g06172(.A0(new_n6236_), .A1(new_n6212_), .B0(new_n6211_), .Y(new_n6237_));
  XOR2X1   g06173(.A(new_n6200_), .B(new_n6196_), .Y(new_n6238_));
  AOI21X1  g06174(.A0(new_n6238_), .A1(new_n6237_), .B0(new_n6201_), .Y(new_n6239_));
  OAI21X1  g06175(.A0(new_n6239_), .A1(new_n6194_), .B0(new_n6193_), .Y(new_n6240_));
  XOR2X1   g06176(.A(new_n6185_), .B(new_n6180_), .Y(new_n6241_));
  INVX1    g06177(.A(new_n6241_), .Y(new_n6242_));
  AOI21X1  g06178(.A0(new_n6242_), .A1(new_n6240_), .B0(new_n6186_), .Y(new_n6243_));
  XOR2X1   g06179(.A(new_n6177_), .B(new_n3289_), .Y(new_n6244_));
  XOR2X1   g06180(.A(new_n6244_), .B(new_n6174_), .Y(new_n6245_));
  OAI21X1  g06181(.A0(new_n6245_), .A1(new_n6243_), .B0(new_n6179_), .Y(new_n6246_));
  XOR2X1   g06182(.A(new_n6172_), .B(new_n6168_), .Y(new_n6247_));
  AOI21X1  g06183(.A0(new_n6247_), .A1(new_n6246_), .B0(new_n6173_), .Y(new_n6248_));
  OAI21X1  g06184(.A0(new_n6248_), .A1(new_n6166_), .B0(new_n6164_), .Y(new_n6249_));
  AOI21X1  g06185(.A0(new_n6249_), .A1(new_n6155_), .B0(new_n6154_), .Y(new_n6250_));
  OAI21X1  g06186(.A0(new_n6250_), .A1(new_n6147_), .B0(new_n6146_), .Y(new_n6251_));
  XOR2X1   g06187(.A(new_n6138_), .B(new_n6133_), .Y(new_n6252_));
  INVX1    g06188(.A(new_n6252_), .Y(new_n6253_));
  AOI21X1  g06189(.A0(new_n6253_), .A1(new_n6251_), .B0(new_n6139_), .Y(new_n6254_));
  XOR2X1   g06190(.A(new_n6131_), .B(new_n6126_), .Y(new_n6255_));
  NOR2X1   g06191(.A(new_n6255_), .B(new_n6254_), .Y(new_n6256_));
  NOR2X1   g06192(.A(new_n6256_), .B(new_n6132_), .Y(new_n6257_));
  INVX1    g06193(.A(new_n6257_), .Y(new_n6258_));
  XOR2X1   g06194(.A(new_n6124_), .B(new_n6120_), .Y(new_n6259_));
  AOI21X1  g06195(.A0(new_n6259_), .A1(new_n6258_), .B0(new_n6125_), .Y(new_n6260_));
  OR2X1    g06196(.A(new_n6260_), .B(new_n6118_), .Y(new_n6261_));
  OAI21X1  g06197(.A0(new_n6116_), .A1(new_n6115_), .B0(new_n6261_), .Y(new_n6262_));
  AOI21X1  g06198(.A0(new_n6262_), .A1(new_n6111_), .B0(new_n6110_), .Y(new_n6263_));
  NOR2X1   g06199(.A(new_n6263_), .B(new_n6103_), .Y(new_n6264_));
  NOR2X1   g06200(.A(new_n6264_), .B(new_n6102_), .Y(new_n6265_));
  XOR2X1   g06201(.A(new_n6095_), .B(new_n6090_), .Y(new_n6266_));
  OR2X1    g06202(.A(new_n6266_), .B(new_n6265_), .Y(new_n6267_));
  OAI21X1  g06203(.A0(new_n6095_), .A1(new_n6091_), .B0(new_n6267_), .Y(new_n6268_));
  XOR2X1   g06204(.A(new_n6088_), .B(new_n6083_), .Y(new_n6269_));
  INVX1    g06205(.A(new_n6269_), .Y(new_n6270_));
  AOI21X1  g06206(.A0(new_n6270_), .A1(new_n6268_), .B0(new_n6089_), .Y(new_n6271_));
  INVX1    g06207(.A(new_n6271_), .Y(new_n6272_));
  XOR2X1   g06208(.A(new_n6081_), .B(new_n6077_), .Y(new_n6273_));
  AOI21X1  g06209(.A0(new_n6273_), .A1(new_n6272_), .B0(new_n6082_), .Y(new_n6274_));
  OAI21X1  g06210(.A0(new_n6274_), .A1(new_n6075_), .B0(new_n6073_), .Y(new_n6275_));
  AOI21X1  g06211(.A0(new_n6275_), .A1(new_n6066_), .B0(new_n6065_), .Y(new_n6276_));
  NOR2X1   g06212(.A(new_n6276_), .B(new_n6058_), .Y(new_n6277_));
  AOI21X1  g06213(.A0(new_n6057_), .A1(new_n6056_), .B0(new_n6277_), .Y(new_n6278_));
  XOR2X1   g06214(.A(new_n6049_), .B(new_n6044_), .Y(new_n6279_));
  OAI21X1  g06215(.A0(new_n6279_), .A1(new_n6278_), .B0(new_n6051_), .Y(new_n6280_));
  XOR2X1   g06216(.A(new_n6042_), .B(new_n6038_), .Y(new_n6281_));
  AOI21X1  g06217(.A0(new_n6281_), .A1(new_n6280_), .B0(new_n6043_), .Y(new_n6282_));
  INVX1    g06218(.A(new_n6282_), .Y(new_n6283_));
  AOI21X1  g06219(.A0(new_n6283_), .A1(new_n6036_), .B0(new_n6035_), .Y(new_n6284_));
  OR2X1    g06220(.A(new_n6284_), .B(new_n6028_), .Y(new_n6285_));
  OAI21X1  g06221(.A0(new_n6026_), .A1(new_n6024_), .B0(new_n6285_), .Y(new_n6286_));
  AOI21X1  g06222(.A0(new_n6286_), .A1(new_n6020_), .B0(new_n6019_), .Y(new_n6287_));
  OR2X1    g06223(.A(new_n6287_), .B(new_n6011_), .Y(new_n6288_));
  OAI21X1  g06224(.A0(new_n6009_), .A1(new_n6007_), .B0(new_n6288_), .Y(new_n6289_));
  AOI21X1  g06225(.A0(new_n6289_), .A1(new_n6003_), .B0(new_n6002_), .Y(new_n6290_));
  NOR2X1   g06226(.A(new_n6290_), .B(new_n5995_), .Y(new_n6291_));
  AOI21X1  g06227(.A0(new_n5994_), .A1(new_n5993_), .B0(new_n6291_), .Y(new_n6292_));
  NOR2X1   g06228(.A(new_n6292_), .B(new_n5988_), .Y(new_n6293_));
  XOR2X1   g06229(.A(new_n6292_), .B(new_n5987_), .Y(new_n6294_));
  INVX1    g06230(.A(new_n6294_), .Y(new_n6295_));
  XOR2X1   g06231(.A(new_n6290_), .B(new_n5995_), .Y(new_n6296_));
  INVX1    g06232(.A(new_n6296_), .Y(new_n6297_));
  INVX1    g06233(.A(new_n5972_), .Y(new_n6298_));
  INVX1    g06234(.A(\a[0] ), .Y(new_n6299_));
  AND2X1   g06235(.A(\a[1] ), .B(new_n6299_), .Y(new_n6300_));
  AOI22X1  g06236(.A0(new_n6300_), .A1(new_n2649_), .B0(new_n5970_), .B1(new_n2421_), .Y(new_n6301_));
  OAI21X1  g06237(.A0(new_n6298_), .A1(new_n2695_), .B0(new_n6301_), .Y(new_n6302_));
  XOR2X1   g06238(.A(new_n6302_), .B(new_n3431_), .Y(new_n6303_));
  OR2X1    g06239(.A(new_n6303_), .B(new_n6297_), .Y(new_n6304_));
  XOR2X1   g06240(.A(new_n6289_), .B(new_n6003_), .Y(new_n6305_));
  INVX1    g06241(.A(new_n6305_), .Y(new_n6306_));
  INVX1    g06242(.A(new_n6300_), .Y(new_n6307_));
  NOR2X1   g06243(.A(new_n5971_), .B(new_n6299_), .Y(new_n6308_));
  INVX1    g06244(.A(new_n6308_), .Y(new_n6309_));
  OAI22X1  g06245(.A0(new_n6309_), .A1(new_n2648_), .B0(new_n6307_), .B1(new_n2414_), .Y(new_n6310_));
  AOI21X1  g06246(.A0(new_n5970_), .A1(new_n2752_), .B0(new_n6310_), .Y(new_n6311_));
  OAI21X1  g06247(.A0(new_n6298_), .A1(new_n2757_), .B0(new_n6311_), .Y(new_n6312_));
  XOR2X1   g06248(.A(new_n6312_), .B(new_n3431_), .Y(new_n6313_));
  NOR2X1   g06249(.A(new_n6313_), .B(new_n6306_), .Y(new_n6314_));
  XOR2X1   g06250(.A(new_n6287_), .B(new_n6011_), .Y(new_n6315_));
  INVX1    g06251(.A(new_n6315_), .Y(new_n6316_));
  AOI22X1  g06252(.A0(new_n6308_), .A1(new_n2421_), .B0(new_n5970_), .B1(new_n2420_), .Y(new_n6317_));
  OAI21X1  g06253(.A0(new_n6307_), .A1(new_n2379_), .B0(new_n6317_), .Y(new_n6318_));
  AOI21X1  g06254(.A0(new_n5972_), .A1(new_n2416_), .B0(new_n6318_), .Y(new_n6319_));
  XOR2X1   g06255(.A(new_n6319_), .B(\a[2] ), .Y(new_n6320_));
  OR2X1    g06256(.A(new_n6320_), .B(new_n6316_), .Y(new_n6321_));
  XOR2X1   g06257(.A(new_n6286_), .B(new_n6020_), .Y(new_n6322_));
  INVX1    g06258(.A(new_n6322_), .Y(new_n6323_));
  INVX1    g06259(.A(new_n2625_), .Y(new_n6324_));
  INVX1    g06260(.A(new_n5970_), .Y(new_n6325_));
  OAI22X1  g06261(.A0(new_n6307_), .A1(new_n2339_), .B0(new_n6325_), .B1(new_n2287_), .Y(new_n6326_));
  AOI21X1  g06262(.A0(new_n6308_), .A1(new_n2752_), .B0(new_n6326_), .Y(new_n6327_));
  OAI21X1  g06263(.A0(new_n6298_), .A1(new_n6324_), .B0(new_n6327_), .Y(new_n6328_));
  XOR2X1   g06264(.A(new_n6328_), .B(new_n3431_), .Y(new_n6329_));
  NOR2X1   g06265(.A(new_n6329_), .B(new_n6323_), .Y(new_n6330_));
  XOR2X1   g06266(.A(new_n6284_), .B(new_n6028_), .Y(new_n6331_));
  INVX1    g06267(.A(new_n6331_), .Y(new_n6332_));
  OAI22X1  g06268(.A0(new_n6309_), .A1(new_n2339_), .B0(new_n6325_), .B1(new_n2137_), .Y(new_n6333_));
  AOI21X1  g06269(.A0(new_n6300_), .A1(new_n2627_), .B0(new_n6333_), .Y(new_n6334_));
  OAI21X1  g06270(.A0(new_n6298_), .A1(new_n2670_), .B0(new_n6334_), .Y(new_n6335_));
  XOR2X1   g06271(.A(new_n6335_), .B(new_n3431_), .Y(new_n6336_));
  OR2X1    g06272(.A(new_n6336_), .B(new_n6332_), .Y(new_n6337_));
  XOR2X1   g06273(.A(new_n6281_), .B(new_n6280_), .Y(new_n6338_));
  INVX1    g06274(.A(new_n6338_), .Y(new_n6339_));
  XOR2X1   g06275(.A(new_n6273_), .B(new_n6271_), .Y(new_n6340_));
  XOR2X1   g06276(.A(new_n6259_), .B(new_n6258_), .Y(new_n6341_));
  INVX1    g06277(.A(new_n6341_), .Y(new_n6342_));
  XOR2X1   g06278(.A(new_n6247_), .B(new_n6246_), .Y(new_n6343_));
  XOR2X1   g06279(.A(new_n6235_), .B(new_n6234_), .Y(new_n6344_));
  INVX1    g06280(.A(new_n6344_), .Y(new_n6345_));
  INVX1    g06281(.A(new_n6223_), .Y(new_n6346_));
  NAND3X1  g06282(.A(new_n6346_), .B(new_n6221_), .C(\a[5] ), .Y(new_n6347_));
  XOR2X1   g06283(.A(new_n6226_), .B(new_n3289_), .Y(new_n6348_));
  XOR2X1   g06284(.A(new_n6348_), .B(new_n6347_), .Y(new_n6349_));
  NOR3X1   g06285(.A(new_n3431_), .B(\a[1] ), .C(new_n6299_), .Y(new_n6350_));
  INVX1    g06286(.A(new_n6350_), .Y(new_n6351_));
  NOR3X1   g06287(.A(new_n6351_), .B(new_n3822_), .C(new_n3820_), .Y(new_n6352_));
  NAND2X1  g06288(.A(new_n6308_), .B(new_n1706_), .Y(new_n6353_));
  AOI22X1  g06289(.A0(new_n6300_), .A1(new_n3819_), .B0(new_n5970_), .B1(new_n3821_), .Y(new_n6354_));
  AOI21X1  g06290(.A0(new_n6354_), .A1(new_n6353_), .B0(new_n3431_), .Y(new_n6355_));
  AND2X1   g06291(.A(new_n6350_), .B(new_n4165_), .Y(new_n6356_));
  NOR2X1   g06292(.A(new_n6308_), .B(new_n5972_), .Y(new_n6357_));
  OAI21X1  g06293(.A0(new_n6357_), .A1(new_n1784_), .B0(\a[2] ), .Y(new_n6358_));
  INVX1    g06294(.A(\a[1] ), .Y(new_n6359_));
  NOR3X1   g06295(.A(new_n3431_), .B(new_n6359_), .C(\a[0] ), .Y(new_n6360_));
  INVX1    g06296(.A(new_n6360_), .Y(new_n6361_));
  NAND3X1  g06297(.A(\a[2] ), .B(\a[1] ), .C(\a[0] ), .Y(new_n6362_));
  OAI22X1  g06298(.A0(new_n6362_), .A1(new_n1735_), .B0(new_n6361_), .B1(new_n1784_), .Y(new_n6363_));
  OR4X1    g06299(.A(new_n6363_), .B(new_n6358_), .C(new_n6356_), .D(new_n6355_), .Y(new_n6364_));
  NOR3X1   g06300(.A(new_n6364_), .B(new_n6352_), .C(new_n6346_), .Y(new_n6365_));
  OAI21X1  g06301(.A0(new_n6364_), .A1(new_n6352_), .B0(new_n6346_), .Y(new_n6366_));
  AOI22X1  g06302(.A0(new_n6308_), .A1(new_n1676_), .B0(new_n5970_), .B1(new_n3819_), .Y(new_n6367_));
  OAI21X1  g06303(.A0(new_n6307_), .A1(new_n1708_), .B0(new_n6367_), .Y(new_n6368_));
  AOI21X1  g06304(.A0(new_n5972_), .A1(new_n3829_), .B0(new_n6368_), .Y(new_n6369_));
  XOR2X1   g06305(.A(new_n6369_), .B(new_n3431_), .Y(new_n6370_));
  AOI21X1  g06306(.A0(new_n6370_), .A1(new_n6366_), .B0(new_n6365_), .Y(new_n6371_));
  OAI22X1  g06307(.A0(new_n6309_), .A1(new_n1655_), .B0(new_n6307_), .B1(new_n1674_), .Y(new_n6372_));
  AOI21X1  g06308(.A0(new_n5970_), .A1(new_n1706_), .B0(new_n6372_), .Y(new_n6373_));
  OAI21X1  g06309(.A0(new_n6298_), .A1(new_n3773_), .B0(new_n6373_), .Y(new_n6374_));
  XOR2X1   g06310(.A(new_n6374_), .B(new_n3431_), .Y(new_n6375_));
  AOI21X1  g06311(.A0(new_n3821_), .A1(new_n66_), .B0(new_n3289_), .Y(new_n6376_));
  XOR2X1   g06312(.A(new_n6376_), .B(new_n6222_), .Y(new_n6377_));
  AOI21X1  g06313(.A0(new_n6375_), .A1(new_n6371_), .B0(new_n6377_), .Y(new_n6378_));
  NOR2X1   g06314(.A(new_n6375_), .B(new_n6371_), .Y(new_n6379_));
  OAI21X1  g06315(.A0(new_n6379_), .A1(new_n6378_), .B0(new_n6349_), .Y(new_n6380_));
  NOR3X1   g06316(.A(new_n6379_), .B(new_n6378_), .C(new_n6349_), .Y(new_n6381_));
  AOI22X1  g06317(.A0(new_n6300_), .A1(new_n3721_), .B0(new_n5970_), .B1(new_n1676_), .Y(new_n6382_));
  OAI21X1  g06318(.A0(new_n6309_), .A1(new_n1621_), .B0(new_n6382_), .Y(new_n6383_));
  AOI21X1  g06319(.A0(new_n5972_), .A1(new_n3745_), .B0(new_n6383_), .Y(new_n6384_));
  XOR2X1   g06320(.A(new_n6384_), .B(\a[2] ), .Y(new_n6385_));
  OAI21X1  g06321(.A0(new_n6385_), .A1(new_n6381_), .B0(new_n6380_), .Y(new_n6386_));
  OAI22X1  g06322(.A0(new_n6309_), .A1(new_n1586_), .B0(new_n6325_), .B1(new_n1655_), .Y(new_n6387_));
  AOI21X1  g06323(.A0(new_n6300_), .A1(new_n4538_), .B0(new_n6387_), .Y(new_n6388_));
  OAI21X1  g06324(.A0(new_n6298_), .A1(new_n3719_), .B0(new_n6388_), .Y(new_n6389_));
  XOR2X1   g06325(.A(new_n6389_), .B(\a[2] ), .Y(new_n6390_));
  NAND2X1  g06326(.A(new_n6390_), .B(new_n6386_), .Y(new_n6391_));
  XOR2X1   g06327(.A(new_n6233_), .B(new_n6229_), .Y(new_n6392_));
  OAI21X1  g06328(.A0(new_n6390_), .A1(new_n6386_), .B0(new_n6392_), .Y(new_n6393_));
  AOI21X1  g06329(.A0(new_n6393_), .A1(new_n6391_), .B0(new_n6345_), .Y(new_n6394_));
  NAND3X1  g06330(.A(new_n6393_), .B(new_n6391_), .C(new_n6345_), .Y(new_n6395_));
  AOI22X1  g06331(.A0(new_n6308_), .A1(new_n1536_), .B0(new_n6300_), .B1(new_n3480_), .Y(new_n6396_));
  OAI21X1  g06332(.A0(new_n6325_), .A1(new_n1621_), .B0(new_n6396_), .Y(new_n6397_));
  AOI21X1  g06333(.A0(new_n5972_), .A1(new_n3697_), .B0(new_n6397_), .Y(new_n6398_));
  XOR2X1   g06334(.A(new_n6398_), .B(\a[2] ), .Y(new_n6399_));
  INVX1    g06335(.A(new_n6399_), .Y(new_n6400_));
  AOI21X1  g06336(.A0(new_n6400_), .A1(new_n6395_), .B0(new_n6394_), .Y(new_n6401_));
  OAI22X1  g06337(.A0(new_n6309_), .A1(new_n3669_), .B0(new_n6325_), .B1(new_n1586_), .Y(new_n6402_));
  AOI21X1  g06338(.A0(new_n6300_), .A1(new_n1536_), .B0(new_n6402_), .Y(new_n6403_));
  OAI21X1  g06339(.A0(new_n6298_), .A1(new_n3478_), .B0(new_n6403_), .Y(new_n6404_));
  XOR2X1   g06340(.A(new_n6404_), .B(new_n3431_), .Y(new_n6405_));
  XOR2X1   g06341(.A(new_n6236_), .B(new_n6212_), .Y(new_n6406_));
  INVX1    g06342(.A(new_n6406_), .Y(new_n6407_));
  AOI21X1  g06343(.A0(new_n6405_), .A1(new_n6401_), .B0(new_n6407_), .Y(new_n6408_));
  NOR2X1   g06344(.A(new_n6405_), .B(new_n6401_), .Y(new_n6409_));
  OAI22X1  g06345(.A0(new_n6309_), .A1(new_n1465_), .B0(new_n6307_), .B1(new_n3669_), .Y(new_n6410_));
  AOI21X1  g06346(.A0(new_n5970_), .A1(new_n1536_), .B0(new_n6410_), .Y(new_n6411_));
  OAI21X1  g06347(.A0(new_n6298_), .A1(new_n3676_), .B0(new_n6411_), .Y(new_n6412_));
  XOR2X1   g06348(.A(new_n6412_), .B(new_n3431_), .Y(new_n6413_));
  INVX1    g06349(.A(new_n6413_), .Y(new_n6414_));
  NOR3X1   g06350(.A(new_n6414_), .B(new_n6409_), .C(new_n6408_), .Y(new_n6415_));
  XOR2X1   g06351(.A(new_n6238_), .B(new_n6237_), .Y(new_n6416_));
  INVX1    g06352(.A(new_n6416_), .Y(new_n6417_));
  OAI21X1  g06353(.A0(new_n6409_), .A1(new_n6408_), .B0(new_n6414_), .Y(new_n6418_));
  OAI21X1  g06354(.A0(new_n6417_), .A1(new_n6415_), .B0(new_n6418_), .Y(new_n6419_));
  OAI22X1  g06355(.A0(new_n6309_), .A1(new_n1423_), .B0(new_n6325_), .B1(new_n3669_), .Y(new_n6420_));
  AOI21X1  g06356(.A0(new_n6300_), .A1(new_n1800_), .B0(new_n6420_), .Y(new_n6421_));
  OAI21X1  g06357(.A0(new_n6298_), .A1(new_n3667_), .B0(new_n6421_), .Y(new_n6422_));
  XOR2X1   g06358(.A(new_n6422_), .B(new_n3431_), .Y(new_n6423_));
  INVX1    g06359(.A(new_n6423_), .Y(new_n6424_));
  XOR2X1   g06360(.A(new_n6239_), .B(new_n6194_), .Y(new_n6425_));
  OAI21X1  g06361(.A0(new_n6424_), .A1(new_n6419_), .B0(new_n6425_), .Y(new_n6426_));
  NAND2X1  g06362(.A(new_n6424_), .B(new_n6419_), .Y(new_n6427_));
  XOR2X1   g06363(.A(new_n6242_), .B(new_n6240_), .Y(new_n6428_));
  INVX1    g06364(.A(new_n6428_), .Y(new_n6429_));
  AOI21X1  g06365(.A0(new_n6427_), .A1(new_n6426_), .B0(new_n6429_), .Y(new_n6430_));
  NAND3X1  g06366(.A(new_n6429_), .B(new_n6427_), .C(new_n6426_), .Y(new_n6431_));
  AOI22X1  g06367(.A0(new_n6300_), .A1(new_n3327_), .B0(new_n5970_), .B1(new_n1800_), .Y(new_n6432_));
  OAI21X1  g06368(.A0(new_n6309_), .A1(new_n1389_), .B0(new_n6432_), .Y(new_n6433_));
  AOI21X1  g06369(.A0(new_n5972_), .A1(new_n3497_), .B0(new_n6433_), .Y(new_n6434_));
  XOR2X1   g06370(.A(new_n6434_), .B(\a[2] ), .Y(new_n6435_));
  INVX1    g06371(.A(new_n6435_), .Y(new_n6436_));
  AOI21X1  g06372(.A0(new_n6436_), .A1(new_n6431_), .B0(new_n6430_), .Y(new_n6437_));
  XOR2X1   g06373(.A(new_n6245_), .B(new_n6243_), .Y(new_n6438_));
  INVX1    g06374(.A(new_n6438_), .Y(new_n6439_));
  NOR2X1   g06375(.A(new_n6439_), .B(new_n6437_), .Y(new_n6440_));
  AOI22X1  g06376(.A0(new_n6308_), .A1(new_n1357_), .B0(new_n5970_), .B1(new_n3327_), .Y(new_n6441_));
  OAI21X1  g06377(.A0(new_n6307_), .A1(new_n1389_), .B0(new_n6441_), .Y(new_n6442_));
  AOI21X1  g06378(.A0(new_n5972_), .A1(new_n3326_), .B0(new_n6442_), .Y(new_n6443_));
  XOR2X1   g06379(.A(new_n6443_), .B(\a[2] ), .Y(new_n6444_));
  AOI21X1  g06380(.A0(new_n6439_), .A1(new_n6437_), .B0(new_n6444_), .Y(new_n6445_));
  OAI21X1  g06381(.A0(new_n6445_), .A1(new_n6440_), .B0(new_n6343_), .Y(new_n6446_));
  NOR3X1   g06382(.A(new_n6445_), .B(new_n6440_), .C(new_n6343_), .Y(new_n6447_));
  AOI22X1  g06383(.A0(new_n6308_), .A1(new_n3055_), .B0(new_n6300_), .B1(new_n1357_), .Y(new_n6448_));
  OAI21X1  g06384(.A0(new_n6325_), .A1(new_n1389_), .B0(new_n6448_), .Y(new_n6449_));
  AOI21X1  g06385(.A0(new_n5972_), .A1(new_n3425_), .B0(new_n6449_), .Y(new_n6450_));
  XOR2X1   g06386(.A(new_n6450_), .B(\a[2] ), .Y(new_n6451_));
  OAI21X1  g06387(.A0(new_n6451_), .A1(new_n6447_), .B0(new_n6446_), .Y(new_n6452_));
  OAI22X1  g06388(.A0(new_n6309_), .A1(new_n1294_), .B0(new_n6325_), .B1(new_n1358_), .Y(new_n6453_));
  AOI21X1  g06389(.A0(new_n6300_), .A1(new_n3055_), .B0(new_n6453_), .Y(new_n6454_));
  OAI21X1  g06390(.A0(new_n6298_), .A1(new_n3340_), .B0(new_n6454_), .Y(new_n6455_));
  XOR2X1   g06391(.A(new_n6455_), .B(new_n3431_), .Y(new_n6456_));
  INVX1    g06392(.A(new_n6456_), .Y(new_n6457_));
  XOR2X1   g06393(.A(new_n6248_), .B(new_n6166_), .Y(new_n6458_));
  OAI21X1  g06394(.A0(new_n6457_), .A1(new_n6452_), .B0(new_n6458_), .Y(new_n6459_));
  NAND2X1  g06395(.A(new_n6457_), .B(new_n6452_), .Y(new_n6460_));
  OAI22X1  g06396(.A0(new_n6309_), .A1(new_n1236_), .B0(new_n6325_), .B1(new_n1339_), .Y(new_n6461_));
  AOI21X1  g06397(.A0(new_n6300_), .A1(new_n3342_), .B0(new_n6461_), .Y(new_n6462_));
  OAI21X1  g06398(.A0(new_n6298_), .A1(new_n3053_), .B0(new_n6462_), .Y(new_n6463_));
  XOR2X1   g06399(.A(new_n6463_), .B(new_n3431_), .Y(new_n6464_));
  NAND3X1  g06400(.A(new_n6464_), .B(new_n6460_), .C(new_n6459_), .Y(new_n6465_));
  XOR2X1   g06401(.A(new_n6249_), .B(new_n6155_), .Y(new_n6466_));
  AOI21X1  g06402(.A0(new_n6460_), .A1(new_n6459_), .B0(new_n6464_), .Y(new_n6467_));
  AOI21X1  g06403(.A0(new_n6466_), .A1(new_n6465_), .B0(new_n6467_), .Y(new_n6468_));
  OAI22X1  g06404(.A0(new_n6309_), .A1(new_n1189_), .B0(new_n6307_), .B1(new_n1236_), .Y(new_n6469_));
  AOI21X1  g06405(.A0(new_n5970_), .A1(new_n3342_), .B0(new_n6469_), .Y(new_n6470_));
  OAI21X1  g06406(.A0(new_n6298_), .A1(new_n3180_), .B0(new_n6470_), .Y(new_n6471_));
  XOR2X1   g06407(.A(new_n6471_), .B(new_n3431_), .Y(new_n6472_));
  XOR2X1   g06408(.A(new_n6250_), .B(new_n6147_), .Y(new_n6473_));
  INVX1    g06409(.A(new_n6473_), .Y(new_n6474_));
  AOI21X1  g06410(.A0(new_n6472_), .A1(new_n6468_), .B0(new_n6474_), .Y(new_n6475_));
  NOR2X1   g06411(.A(new_n6472_), .B(new_n6468_), .Y(new_n6476_));
  XOR2X1   g06412(.A(new_n6253_), .B(new_n6251_), .Y(new_n6477_));
  OAI21X1  g06413(.A0(new_n6476_), .A1(new_n6475_), .B0(new_n6477_), .Y(new_n6478_));
  NOR3X1   g06414(.A(new_n6477_), .B(new_n6476_), .C(new_n6475_), .Y(new_n6479_));
  AOI22X1  g06415(.A0(new_n6308_), .A1(new_n1126_), .B0(new_n5970_), .B1(new_n2977_), .Y(new_n6480_));
  OAI21X1  g06416(.A0(new_n6307_), .A1(new_n1189_), .B0(new_n6480_), .Y(new_n6481_));
  AOI21X1  g06417(.A0(new_n5972_), .A1(new_n2976_), .B0(new_n6481_), .Y(new_n6482_));
  XOR2X1   g06418(.A(new_n6482_), .B(\a[2] ), .Y(new_n6483_));
  OAI21X1  g06419(.A0(new_n6483_), .A1(new_n6479_), .B0(new_n6478_), .Y(new_n6484_));
  XOR2X1   g06420(.A(new_n6255_), .B(new_n6254_), .Y(new_n6485_));
  NAND2X1  g06421(.A(new_n6485_), .B(new_n6484_), .Y(new_n6486_));
  AOI22X1  g06422(.A0(new_n6308_), .A1(new_n1822_), .B0(new_n6300_), .B1(new_n1126_), .Y(new_n6487_));
  OAI21X1  g06423(.A0(new_n6325_), .A1(new_n1189_), .B0(new_n6487_), .Y(new_n6488_));
  AOI21X1  g06424(.A0(new_n5972_), .A1(new_n2963_), .B0(new_n6488_), .Y(new_n6489_));
  XOR2X1   g06425(.A(new_n6489_), .B(\a[2] ), .Y(new_n6490_));
  INVX1    g06426(.A(new_n6490_), .Y(new_n6491_));
  OAI21X1  g06427(.A0(new_n6485_), .A1(new_n6484_), .B0(new_n6491_), .Y(new_n6492_));
  AOI21X1  g06428(.A0(new_n6492_), .A1(new_n6486_), .B0(new_n6342_), .Y(new_n6493_));
  NAND3X1  g06429(.A(new_n6492_), .B(new_n6486_), .C(new_n6342_), .Y(new_n6494_));
  AOI22X1  g06430(.A0(new_n6308_), .A1(new_n2603_), .B0(new_n5970_), .B1(new_n1126_), .Y(new_n6495_));
  OAI21X1  g06431(.A0(new_n6307_), .A1(new_n1065_), .B0(new_n6495_), .Y(new_n6496_));
  AOI21X1  g06432(.A0(new_n5972_), .A1(new_n2824_), .B0(new_n6496_), .Y(new_n6497_));
  XOR2X1   g06433(.A(new_n6497_), .B(\a[2] ), .Y(new_n6498_));
  INVX1    g06434(.A(new_n6498_), .Y(new_n6499_));
  AOI21X1  g06435(.A0(new_n6499_), .A1(new_n6494_), .B0(new_n6493_), .Y(new_n6500_));
  OAI22X1  g06436(.A0(new_n6309_), .A1(new_n957_), .B0(new_n6307_), .B1(new_n985_), .Y(new_n6501_));
  AOI21X1  g06437(.A0(new_n5970_), .A1(new_n1822_), .B0(new_n6501_), .Y(new_n6502_));
  OAI21X1  g06438(.A0(new_n6298_), .A1(new_n2833_), .B0(new_n6502_), .Y(new_n6503_));
  XOR2X1   g06439(.A(new_n6503_), .B(new_n3431_), .Y(new_n6504_));
  XOR2X1   g06440(.A(new_n6260_), .B(new_n6117_), .Y(new_n6505_));
  AOI21X1  g06441(.A0(new_n6504_), .A1(new_n6500_), .B0(new_n6505_), .Y(new_n6506_));
  AND2X1   g06442(.A(new_n6485_), .B(new_n6484_), .Y(new_n6507_));
  INVX1    g06443(.A(new_n6343_), .Y(new_n6508_));
  OR2X1    g06444(.A(new_n6439_), .B(new_n6437_), .Y(new_n6509_));
  AND2X1   g06445(.A(new_n6390_), .B(new_n6386_), .Y(new_n6510_));
  INVX1    g06446(.A(new_n6347_), .Y(new_n6511_));
  XOR2X1   g06447(.A(new_n6348_), .B(new_n6511_), .Y(new_n6512_));
  OR4X1    g06448(.A(new_n6298_), .B(new_n3822_), .C(new_n3820_), .D(new_n3431_), .Y(new_n6513_));
  NOR4X1   g06449(.A(new_n6363_), .B(new_n6358_), .C(new_n6356_), .D(new_n6355_), .Y(new_n6514_));
  NAND3X1  g06450(.A(new_n6514_), .B(new_n6513_), .C(new_n6223_), .Y(new_n6515_));
  AOI21X1  g06451(.A0(new_n6514_), .A1(new_n6513_), .B0(new_n6223_), .Y(new_n6516_));
  XOR2X1   g06452(.A(new_n6369_), .B(\a[2] ), .Y(new_n6517_));
  OAI21X1  g06453(.A0(new_n6517_), .A1(new_n6516_), .B0(new_n6515_), .Y(new_n6518_));
  XOR2X1   g06454(.A(new_n6374_), .B(\a[2] ), .Y(new_n6519_));
  INVX1    g06455(.A(new_n6376_), .Y(new_n6520_));
  XOR2X1   g06456(.A(new_n6520_), .B(new_n6222_), .Y(new_n6521_));
  OAI21X1  g06457(.A0(new_n6519_), .A1(new_n6518_), .B0(new_n6521_), .Y(new_n6522_));
  OR2X1    g06458(.A(new_n6375_), .B(new_n6371_), .Y(new_n6523_));
  AOI21X1  g06459(.A0(new_n6523_), .A1(new_n6522_), .B0(new_n6512_), .Y(new_n6524_));
  NAND3X1  g06460(.A(new_n6523_), .B(new_n6522_), .C(new_n6512_), .Y(new_n6525_));
  XOR2X1   g06461(.A(new_n6384_), .B(new_n3431_), .Y(new_n6526_));
  AOI21X1  g06462(.A0(new_n6526_), .A1(new_n6525_), .B0(new_n6524_), .Y(new_n6527_));
  XOR2X1   g06463(.A(new_n6389_), .B(new_n3431_), .Y(new_n6528_));
  INVX1    g06464(.A(new_n6392_), .Y(new_n6529_));
  AOI21X1  g06465(.A0(new_n6528_), .A1(new_n6527_), .B0(new_n6529_), .Y(new_n6530_));
  OAI21X1  g06466(.A0(new_n6530_), .A1(new_n6510_), .B0(new_n6344_), .Y(new_n6531_));
  NOR3X1   g06467(.A(new_n6530_), .B(new_n6510_), .C(new_n6344_), .Y(new_n6532_));
  OAI21X1  g06468(.A0(new_n6399_), .A1(new_n6532_), .B0(new_n6531_), .Y(new_n6533_));
  INVX1    g06469(.A(new_n6405_), .Y(new_n6534_));
  OAI21X1  g06470(.A0(new_n6534_), .A1(new_n6533_), .B0(new_n6406_), .Y(new_n6535_));
  OR2X1    g06471(.A(new_n6405_), .B(new_n6401_), .Y(new_n6536_));
  NAND3X1  g06472(.A(new_n6413_), .B(new_n6536_), .C(new_n6535_), .Y(new_n6537_));
  AOI21X1  g06473(.A0(new_n6536_), .A1(new_n6535_), .B0(new_n6413_), .Y(new_n6538_));
  AOI21X1  g06474(.A0(new_n6416_), .A1(new_n6537_), .B0(new_n6538_), .Y(new_n6539_));
  INVX1    g06475(.A(new_n6425_), .Y(new_n6540_));
  AOI21X1  g06476(.A0(new_n6423_), .A1(new_n6539_), .B0(new_n6540_), .Y(new_n6541_));
  AND2X1   g06477(.A(new_n6424_), .B(new_n6419_), .Y(new_n6542_));
  OAI21X1  g06478(.A0(new_n6542_), .A1(new_n6541_), .B0(new_n6428_), .Y(new_n6543_));
  NOR3X1   g06479(.A(new_n6428_), .B(new_n6542_), .C(new_n6541_), .Y(new_n6544_));
  OAI21X1  g06480(.A0(new_n6435_), .A1(new_n6544_), .B0(new_n6543_), .Y(new_n6545_));
  INVX1    g06481(.A(new_n6444_), .Y(new_n6546_));
  OAI21X1  g06482(.A0(new_n6438_), .A1(new_n6545_), .B0(new_n6546_), .Y(new_n6547_));
  AOI21X1  g06483(.A0(new_n6547_), .A1(new_n6509_), .B0(new_n6508_), .Y(new_n6548_));
  NAND3X1  g06484(.A(new_n6547_), .B(new_n6509_), .C(new_n6508_), .Y(new_n6549_));
  INVX1    g06485(.A(new_n6451_), .Y(new_n6550_));
  AOI21X1  g06486(.A0(new_n6550_), .A1(new_n6549_), .B0(new_n6548_), .Y(new_n6551_));
  INVX1    g06487(.A(new_n6458_), .Y(new_n6552_));
  AOI21X1  g06488(.A0(new_n6456_), .A1(new_n6551_), .B0(new_n6552_), .Y(new_n6553_));
  AND2X1   g06489(.A(new_n6457_), .B(new_n6452_), .Y(new_n6554_));
  INVX1    g06490(.A(new_n6464_), .Y(new_n6555_));
  NOR3X1   g06491(.A(new_n6555_), .B(new_n6554_), .C(new_n6553_), .Y(new_n6556_));
  INVX1    g06492(.A(new_n6466_), .Y(new_n6557_));
  OAI21X1  g06493(.A0(new_n6554_), .A1(new_n6553_), .B0(new_n6555_), .Y(new_n6558_));
  OAI21X1  g06494(.A0(new_n6557_), .A1(new_n6556_), .B0(new_n6558_), .Y(new_n6559_));
  INVX1    g06495(.A(new_n6472_), .Y(new_n6560_));
  OAI21X1  g06496(.A0(new_n6560_), .A1(new_n6559_), .B0(new_n6473_), .Y(new_n6561_));
  OR2X1    g06497(.A(new_n6472_), .B(new_n6468_), .Y(new_n6562_));
  INVX1    g06498(.A(new_n6477_), .Y(new_n6563_));
  AOI21X1  g06499(.A0(new_n6562_), .A1(new_n6561_), .B0(new_n6563_), .Y(new_n6564_));
  NAND3X1  g06500(.A(new_n6563_), .B(new_n6562_), .C(new_n6561_), .Y(new_n6565_));
  INVX1    g06501(.A(new_n6483_), .Y(new_n6566_));
  AOI21X1  g06502(.A0(new_n6566_), .A1(new_n6565_), .B0(new_n6564_), .Y(new_n6567_));
  INVX1    g06503(.A(new_n6485_), .Y(new_n6568_));
  AOI21X1  g06504(.A0(new_n6568_), .A1(new_n6567_), .B0(new_n6490_), .Y(new_n6569_));
  OAI21X1  g06505(.A0(new_n6569_), .A1(new_n6507_), .B0(new_n6341_), .Y(new_n6570_));
  NOR3X1   g06506(.A(new_n6569_), .B(new_n6507_), .C(new_n6341_), .Y(new_n6571_));
  OAI21X1  g06507(.A0(new_n6498_), .A1(new_n6571_), .B0(new_n6570_), .Y(new_n6572_));
  INVX1    g06508(.A(new_n6504_), .Y(new_n6573_));
  AND2X1   g06509(.A(new_n6573_), .B(new_n6572_), .Y(new_n6574_));
  OAI22X1  g06510(.A0(new_n6309_), .A1(new_n903_), .B0(new_n6325_), .B1(new_n985_), .Y(new_n6575_));
  AOI21X1  g06511(.A0(new_n6300_), .A1(new_n2835_), .B0(new_n6575_), .Y(new_n6576_));
  OAI21X1  g06512(.A0(new_n6298_), .A1(new_n2600_), .B0(new_n6576_), .Y(new_n6577_));
  XOR2X1   g06513(.A(new_n6577_), .B(new_n3431_), .Y(new_n6578_));
  INVX1    g06514(.A(new_n6578_), .Y(new_n6579_));
  NOR3X1   g06515(.A(new_n6579_), .B(new_n6574_), .C(new_n6506_), .Y(new_n6580_));
  XOR2X1   g06516(.A(new_n6262_), .B(new_n6111_), .Y(new_n6581_));
  INVX1    g06517(.A(new_n6581_), .Y(new_n6582_));
  OAI21X1  g06518(.A0(new_n6574_), .A1(new_n6506_), .B0(new_n6579_), .Y(new_n6583_));
  OAI21X1  g06519(.A0(new_n6582_), .A1(new_n6580_), .B0(new_n6583_), .Y(new_n6584_));
  OAI22X1  g06520(.A0(new_n6309_), .A1(new_n847_), .B0(new_n6325_), .B1(new_n957_), .Y(new_n6585_));
  AOI21X1  g06521(.A0(new_n6300_), .A1(new_n2602_), .B0(new_n6585_), .Y(new_n6586_));
  OAI21X1  g06522(.A0(new_n6298_), .A1(new_n2708_), .B0(new_n6586_), .Y(new_n6587_));
  XOR2X1   g06523(.A(new_n6587_), .B(new_n3431_), .Y(new_n6588_));
  INVX1    g06524(.A(new_n6588_), .Y(new_n6589_));
  XOR2X1   g06525(.A(new_n6263_), .B(new_n6103_), .Y(new_n6590_));
  OAI21X1  g06526(.A0(new_n6589_), .A1(new_n6584_), .B0(new_n6590_), .Y(new_n6591_));
  INVX1    g06527(.A(new_n6505_), .Y(new_n6592_));
  OAI21X1  g06528(.A0(new_n6573_), .A1(new_n6572_), .B0(new_n6592_), .Y(new_n6593_));
  NAND2X1  g06529(.A(new_n6573_), .B(new_n6572_), .Y(new_n6594_));
  NAND3X1  g06530(.A(new_n6578_), .B(new_n6594_), .C(new_n6593_), .Y(new_n6595_));
  AOI21X1  g06531(.A0(new_n6594_), .A1(new_n6593_), .B0(new_n6578_), .Y(new_n6596_));
  AOI21X1  g06532(.A0(new_n6581_), .A1(new_n6595_), .B0(new_n6596_), .Y(new_n6597_));
  OR2X1    g06533(.A(new_n6588_), .B(new_n6597_), .Y(new_n6598_));
  XOR2X1   g06534(.A(new_n6266_), .B(new_n6265_), .Y(new_n6599_));
  INVX1    g06535(.A(new_n6599_), .Y(new_n6600_));
  AOI21X1  g06536(.A0(new_n6598_), .A1(new_n6591_), .B0(new_n6600_), .Y(new_n6601_));
  NAND3X1  g06537(.A(new_n6600_), .B(new_n6598_), .C(new_n6591_), .Y(new_n6602_));
  AOI22X1  g06538(.A0(new_n6308_), .A1(new_n2036_), .B0(new_n5970_), .B1(new_n2602_), .Y(new_n6603_));
  OAI21X1  g06539(.A0(new_n6307_), .A1(new_n847_), .B0(new_n6603_), .Y(new_n6604_));
  AOI21X1  g06540(.A0(new_n5972_), .A1(new_n2494_), .B0(new_n6604_), .Y(new_n6605_));
  XOR2X1   g06541(.A(new_n6605_), .B(\a[2] ), .Y(new_n6606_));
  INVX1    g06542(.A(new_n6606_), .Y(new_n6607_));
  AOI21X1  g06543(.A0(new_n6607_), .A1(new_n6602_), .B0(new_n6601_), .Y(new_n6608_));
  XOR2X1   g06544(.A(new_n6270_), .B(new_n6268_), .Y(new_n6609_));
  INVX1    g06545(.A(new_n6609_), .Y(new_n6610_));
  OR2X1    g06546(.A(new_n6610_), .B(new_n6608_), .Y(new_n6611_));
  INVX1    g06547(.A(new_n6590_), .Y(new_n6612_));
  AOI21X1  g06548(.A0(new_n6588_), .A1(new_n6597_), .B0(new_n6612_), .Y(new_n6613_));
  NOR2X1   g06549(.A(new_n6588_), .B(new_n6597_), .Y(new_n6614_));
  OAI21X1  g06550(.A0(new_n6614_), .A1(new_n6613_), .B0(new_n6599_), .Y(new_n6615_));
  NOR3X1   g06551(.A(new_n6599_), .B(new_n6614_), .C(new_n6613_), .Y(new_n6616_));
  OAI21X1  g06552(.A0(new_n6606_), .A1(new_n6616_), .B0(new_n6615_), .Y(new_n6617_));
  AOI22X1  g06553(.A0(new_n6308_), .A1(new_n2049_), .B0(new_n5970_), .B1(new_n2481_), .Y(new_n6618_));
  OAI21X1  g06554(.A0(new_n6307_), .A1(new_n783_), .B0(new_n6618_), .Y(new_n6619_));
  AOI21X1  g06555(.A0(new_n5972_), .A1(new_n2480_), .B0(new_n6619_), .Y(new_n6620_));
  XOR2X1   g06556(.A(new_n6620_), .B(\a[2] ), .Y(new_n6621_));
  INVX1    g06557(.A(new_n6621_), .Y(new_n6622_));
  OAI21X1  g06558(.A0(new_n6609_), .A1(new_n6617_), .B0(new_n6622_), .Y(new_n6623_));
  AOI21X1  g06559(.A0(new_n6623_), .A1(new_n6611_), .B0(new_n6340_), .Y(new_n6624_));
  NAND3X1  g06560(.A(new_n6623_), .B(new_n6611_), .C(new_n6340_), .Y(new_n6625_));
  AOI22X1  g06561(.A0(new_n6308_), .A1(new_n1886_), .B0(new_n5970_), .B1(new_n2036_), .Y(new_n6626_));
  OAI21X1  g06562(.A0(new_n6307_), .A1(new_n690_), .B0(new_n6626_), .Y(new_n6627_));
  AOI21X1  g06563(.A0(new_n5972_), .A1(new_n2035_), .B0(new_n6627_), .Y(new_n6628_));
  XOR2X1   g06564(.A(new_n6628_), .B(\a[2] ), .Y(new_n6629_));
  INVX1    g06565(.A(new_n6629_), .Y(new_n6630_));
  AOI21X1  g06566(.A0(new_n6630_), .A1(new_n6625_), .B0(new_n6624_), .Y(new_n6631_));
  OAI22X1  g06567(.A0(new_n6309_), .A1(new_n520_), .B0(new_n6325_), .B1(new_n690_), .Y(new_n6632_));
  AOI21X1  g06568(.A0(new_n6300_), .A1(new_n1886_), .B0(new_n6632_), .Y(new_n6633_));
  OAI21X1  g06569(.A0(new_n6298_), .A1(new_n3114_), .B0(new_n6633_), .Y(new_n6634_));
  XOR2X1   g06570(.A(new_n6634_), .B(new_n3431_), .Y(new_n6635_));
  XOR2X1   g06571(.A(new_n6274_), .B(new_n6075_), .Y(new_n6636_));
  INVX1    g06572(.A(new_n6636_), .Y(new_n6637_));
  AOI21X1  g06573(.A0(new_n6635_), .A1(new_n6631_), .B0(new_n6637_), .Y(new_n6638_));
  INVX1    g06574(.A(new_n6340_), .Y(new_n6639_));
  NOR2X1   g06575(.A(new_n6610_), .B(new_n6608_), .Y(new_n6640_));
  AOI21X1  g06576(.A0(new_n6610_), .A1(new_n6608_), .B0(new_n6621_), .Y(new_n6641_));
  OAI21X1  g06577(.A0(new_n6641_), .A1(new_n6640_), .B0(new_n6639_), .Y(new_n6642_));
  NOR3X1   g06578(.A(new_n6641_), .B(new_n6640_), .C(new_n6639_), .Y(new_n6643_));
  OAI21X1  g06579(.A0(new_n6629_), .A1(new_n6643_), .B0(new_n6642_), .Y(new_n6644_));
  INVX1    g06580(.A(new_n6635_), .Y(new_n6645_));
  AND2X1   g06581(.A(new_n6645_), .B(new_n6644_), .Y(new_n6646_));
  OAI22X1  g06582(.A0(new_n6309_), .A1(new_n1879_), .B0(new_n6325_), .B1(new_n623_), .Y(new_n6647_));
  AOI21X1  g06583(.A0(new_n6300_), .A1(new_n2048_), .B0(new_n6647_), .Y(new_n6648_));
  OAI21X1  g06584(.A0(new_n6298_), .A1(new_n1881_), .B0(new_n6648_), .Y(new_n6649_));
  XOR2X1   g06585(.A(new_n6649_), .B(new_n3431_), .Y(new_n6650_));
  INVX1    g06586(.A(new_n6650_), .Y(new_n6651_));
  NOR3X1   g06587(.A(new_n6651_), .B(new_n6646_), .C(new_n6638_), .Y(new_n6652_));
  XOR2X1   g06588(.A(new_n6275_), .B(new_n6066_), .Y(new_n6653_));
  INVX1    g06589(.A(new_n6653_), .Y(new_n6654_));
  OAI21X1  g06590(.A0(new_n6646_), .A1(new_n6638_), .B0(new_n6651_), .Y(new_n6655_));
  OAI21X1  g06591(.A0(new_n6654_), .A1(new_n6652_), .B0(new_n6655_), .Y(new_n6656_));
  OAI22X1  g06592(.A0(new_n6309_), .A1(new_n2183_), .B0(new_n6325_), .B1(new_n520_), .Y(new_n6657_));
  AOI21X1  g06593(.A0(new_n6300_), .A1(new_n1887_), .B0(new_n6657_), .Y(new_n6658_));
  OAI21X1  g06594(.A0(new_n6298_), .A1(new_n2243_), .B0(new_n6658_), .Y(new_n6659_));
  XOR2X1   g06595(.A(new_n6659_), .B(new_n3431_), .Y(new_n6660_));
  INVX1    g06596(.A(new_n6660_), .Y(new_n6661_));
  XOR2X1   g06597(.A(new_n6276_), .B(new_n6058_), .Y(new_n6662_));
  OAI21X1  g06598(.A0(new_n6661_), .A1(new_n6656_), .B0(new_n6662_), .Y(new_n6663_));
  OAI21X1  g06599(.A0(new_n6645_), .A1(new_n6644_), .B0(new_n6636_), .Y(new_n6664_));
  NAND2X1  g06600(.A(new_n6645_), .B(new_n6644_), .Y(new_n6665_));
  NAND3X1  g06601(.A(new_n6650_), .B(new_n6665_), .C(new_n6664_), .Y(new_n6666_));
  AOI21X1  g06602(.A0(new_n6665_), .A1(new_n6664_), .B0(new_n6650_), .Y(new_n6667_));
  AOI21X1  g06603(.A0(new_n6653_), .A1(new_n6666_), .B0(new_n6667_), .Y(new_n6668_));
  OR2X1    g06604(.A(new_n6660_), .B(new_n6668_), .Y(new_n6669_));
  XOR2X1   g06605(.A(new_n6279_), .B(new_n6278_), .Y(new_n6670_));
  INVX1    g06606(.A(new_n6670_), .Y(new_n6671_));
  AOI21X1  g06607(.A0(new_n6669_), .A1(new_n6663_), .B0(new_n6671_), .Y(new_n6672_));
  NAND3X1  g06608(.A(new_n6671_), .B(new_n6669_), .C(new_n6663_), .Y(new_n6673_));
  AOI22X1  g06609(.A0(new_n6308_), .A1(new_n2093_), .B0(new_n5970_), .B1(new_n1887_), .Y(new_n6674_));
  OAI21X1  g06610(.A0(new_n6307_), .A1(new_n2183_), .B0(new_n6674_), .Y(new_n6675_));
  AOI21X1  g06611(.A0(new_n5972_), .A1(new_n2430_), .B0(new_n6675_), .Y(new_n6676_));
  XOR2X1   g06612(.A(new_n6676_), .B(\a[2] ), .Y(new_n6677_));
  INVX1    g06613(.A(new_n6677_), .Y(new_n6678_));
  AOI21X1  g06614(.A0(new_n6678_), .A1(new_n6673_), .B0(new_n6672_), .Y(new_n6679_));
  OR2X1    g06615(.A(new_n6679_), .B(new_n6339_), .Y(new_n6680_));
  INVX1    g06616(.A(new_n6662_), .Y(new_n6681_));
  AOI21X1  g06617(.A0(new_n6660_), .A1(new_n6668_), .B0(new_n6681_), .Y(new_n6682_));
  NOR2X1   g06618(.A(new_n6660_), .B(new_n6668_), .Y(new_n6683_));
  OAI21X1  g06619(.A0(new_n6683_), .A1(new_n6682_), .B0(new_n6670_), .Y(new_n6684_));
  NOR3X1   g06620(.A(new_n6670_), .B(new_n6683_), .C(new_n6682_), .Y(new_n6685_));
  OAI21X1  g06621(.A0(new_n6677_), .A1(new_n6685_), .B0(new_n6684_), .Y(new_n6686_));
  AOI22X1  g06622(.A0(new_n6308_), .A1(new_n2252_), .B0(new_n5970_), .B1(new_n2246_), .Y(new_n6687_));
  OAI21X1  g06623(.A0(new_n6307_), .A1(new_n2092_), .B0(new_n6687_), .Y(new_n6688_));
  AOI21X1  g06624(.A0(new_n5972_), .A1(new_n2201_), .B0(new_n6688_), .Y(new_n6689_));
  XOR2X1   g06625(.A(new_n6689_), .B(\a[2] ), .Y(new_n6690_));
  INVX1    g06626(.A(new_n6690_), .Y(new_n6691_));
  OAI21X1  g06627(.A0(new_n6686_), .A1(new_n6338_), .B0(new_n6691_), .Y(new_n6692_));
  OAI22X1  g06628(.A0(new_n6309_), .A1(new_n2287_), .B0(new_n6325_), .B1(new_n2092_), .Y(new_n6693_));
  AOI21X1  g06629(.A0(new_n6300_), .A1(new_n2252_), .B0(new_n6693_), .Y(new_n6694_));
  OAI21X1  g06630(.A0(new_n6298_), .A1(new_n2295_), .B0(new_n6694_), .Y(new_n6695_));
  XOR2X1   g06631(.A(new_n6695_), .B(new_n3431_), .Y(new_n6696_));
  NAND3X1  g06632(.A(new_n6696_), .B(new_n6692_), .C(new_n6680_), .Y(new_n6697_));
  XOR2X1   g06633(.A(new_n6283_), .B(new_n6036_), .Y(new_n6698_));
  AOI21X1  g06634(.A0(new_n6692_), .A1(new_n6680_), .B0(new_n6696_), .Y(new_n6699_));
  AOI21X1  g06635(.A0(new_n6698_), .A1(new_n6697_), .B0(new_n6699_), .Y(new_n6700_));
  XOR2X1   g06636(.A(new_n6336_), .B(new_n6331_), .Y(new_n6701_));
  OAI21X1  g06637(.A0(new_n6701_), .A1(new_n6700_), .B0(new_n6337_), .Y(new_n6702_));
  XOR2X1   g06638(.A(new_n6329_), .B(new_n6323_), .Y(new_n6703_));
  AOI21X1  g06639(.A0(new_n6703_), .A1(new_n6702_), .B0(new_n6330_), .Y(new_n6704_));
  XOR2X1   g06640(.A(new_n6320_), .B(new_n6315_), .Y(new_n6705_));
  OAI21X1  g06641(.A0(new_n6705_), .A1(new_n6704_), .B0(new_n6321_), .Y(new_n6706_));
  XOR2X1   g06642(.A(new_n6313_), .B(new_n6305_), .Y(new_n6707_));
  INVX1    g06643(.A(new_n6707_), .Y(new_n6708_));
  AOI21X1  g06644(.A0(new_n6708_), .A1(new_n6706_), .B0(new_n6314_), .Y(new_n6709_));
  XOR2X1   g06645(.A(new_n6303_), .B(new_n6296_), .Y(new_n6710_));
  OAI21X1  g06646(.A0(new_n6710_), .A1(new_n6709_), .B0(new_n6304_), .Y(new_n6711_));
  AOI21X1  g06647(.A0(new_n6711_), .A1(new_n6295_), .B0(new_n6293_), .Y(new_n6712_));
  XOR2X1   g06648(.A(new_n5984_), .B(new_n5983_), .Y(new_n6713_));
  INVX1    g06649(.A(new_n6713_), .Y(new_n6714_));
  OAI21X1  g06650(.A0(new_n6714_), .A1(new_n6712_), .B0(new_n5986_), .Y(new_n6715_));
  XOR2X1   g06651(.A(new_n5968_), .B(new_n5967_), .Y(new_n6716_));
  AOI21X1  g06652(.A0(new_n6716_), .A1(new_n6715_), .B0(new_n5969_), .Y(new_n6717_));
  OAI21X1  g06653(.A0(new_n6717_), .A1(new_n5670_), .B0(new_n5668_), .Y(new_n6718_));
  XOR2X1   g06654(.A(new_n5384_), .B(new_n5381_), .Y(new_n6719_));
  AOI21X1  g06655(.A0(new_n6719_), .A1(new_n6718_), .B0(new_n5385_), .Y(new_n6720_));
  XOR2X1   g06656(.A(new_n5114_), .B(new_n5113_), .Y(new_n6721_));
  INVX1    g06657(.A(new_n6721_), .Y(new_n6722_));
  OAI21X1  g06658(.A0(new_n6722_), .A1(new_n6720_), .B0(new_n5116_), .Y(new_n6723_));
  AOI21X1  g06659(.A0(new_n6723_), .A1(new_n4879_), .B0(new_n4878_), .Y(new_n6724_));
  OAI21X1  g06660(.A0(new_n6724_), .A1(new_n4648_), .B0(new_n4646_), .Y(new_n6725_));
  XOR2X1   g06661(.A(new_n4445_), .B(new_n4444_), .Y(new_n6726_));
  AOI21X1  g06662(.A0(new_n6726_), .A1(new_n6725_), .B0(new_n4446_), .Y(new_n6727_));
  OAI21X1  g06663(.A0(new_n6727_), .A1(new_n4258_), .B0(new_n4256_), .Y(new_n6728_));
  XOR2X1   g06664(.A(new_n4091_), .B(new_n4088_), .Y(new_n6729_));
  AOI21X1  g06665(.A0(new_n6729_), .A1(new_n6728_), .B0(new_n4092_), .Y(new_n6730_));
  XOR2X1   g06666(.A(new_n4001_), .B(new_n4000_), .Y(new_n6731_));
  INVX1    g06667(.A(new_n6731_), .Y(new_n6732_));
  OAI21X1  g06668(.A0(new_n6732_), .A1(new_n6730_), .B0(new_n4003_), .Y(new_n6733_));
  AOI21X1  g06669(.A0(new_n6733_), .A1(new_n3917_), .B0(new_n3916_), .Y(new_n6734_));
  OAI21X1  g06670(.A0(new_n6734_), .A1(new_n3640_), .B0(new_n3638_), .Y(new_n6735_));
  AOI21X1  g06671(.A0(new_n6735_), .A1(new_n3561_), .B0(new_n3560_), .Y(new_n6736_));
  OAI21X1  g06672(.A0(new_n6736_), .A1(new_n3399_), .B0(new_n3396_), .Y(new_n6737_));
  XOR2X1   g06673(.A(new_n3242_), .B(new_n3241_), .Y(new_n6738_));
  AOI21X1  g06674(.A0(new_n6738_), .A1(new_n6737_), .B0(new_n3243_), .Y(new_n6739_));
  OAI21X1  g06675(.A0(new_n6739_), .A1(new_n3164_), .B0(new_n3162_), .Y(new_n6740_));
  AOI21X1  g06676(.A0(new_n6740_), .A1(new_n3107_), .B0(new_n3104_), .Y(new_n6741_));
  OAI21X1  g06677(.A0(new_n6741_), .A1(new_n2887_), .B0(new_n2885_), .Y(new_n6742_));
  XOR2X1   g06678(.A(new_n2767_), .B(new_n2766_), .Y(new_n6743_));
  AOI21X1  g06679(.A0(new_n6743_), .A1(new_n6742_), .B0(new_n2768_), .Y(new_n6744_));
  XOR2X1   g06680(.A(new_n6744_), .B(new_n2703_), .Y(new_n6745_));
  NOR2X1   g06681(.A(new_n2701_), .B(new_n2662_), .Y(new_n6746_));
  INVX1    g06682(.A(new_n6746_), .Y(new_n6747_));
  OAI21X1  g06683(.A0(new_n6744_), .A1(new_n2703_), .B0(new_n6747_), .Y(new_n6748_));
  INVX1    g06684(.A(new_n2429_), .Y(new_n6749_));
  NOR2X1   g06685(.A(new_n2660_), .B(new_n2635_), .Y(new_n6750_));
  AOI21X1  g06686(.A0(new_n2661_), .A1(new_n6749_), .B0(new_n6750_), .Y(new_n6751_));
  INVX1    g06687(.A(new_n6751_), .Y(new_n6752_));
  NOR2X1   g06688(.A(new_n2297_), .B(new_n2251_), .Y(new_n6753_));
  INVX1    g06689(.A(new_n6753_), .Y(new_n6754_));
  INVX1    g06690(.A(new_n2298_), .Y(new_n6755_));
  OAI21X1  g06691(.A0(new_n2428_), .A1(new_n6755_), .B0(new_n6754_), .Y(new_n6756_));
  OAI22X1  g06692(.A0(new_n2648_), .A1(new_n2626_), .B0(new_n2419_), .B1(new_n2414_), .Y(new_n6757_));
  AOI21X1  g06693(.A0(new_n2424_), .A1(new_n2752_), .B0(new_n6757_), .Y(new_n6758_));
  OAI21X1  g06694(.A0(new_n2757_), .A1(new_n2665_), .B0(new_n6758_), .Y(new_n6759_));
  XOR2X1   g06695(.A(new_n6759_), .B(new_n89_), .Y(new_n6760_));
  OR2X1    g06696(.A(new_n6760_), .B(new_n6756_), .Y(new_n6761_));
  INVX1    g06697(.A(new_n2205_), .Y(new_n6762_));
  INVX1    g06698(.A(new_n2249_), .Y(new_n6763_));
  AND2X1   g06699(.A(new_n6763_), .B(new_n2242_), .Y(new_n6764_));
  INVX1    g06700(.A(new_n6764_), .Y(new_n6765_));
  OAI21X1  g06701(.A0(new_n2250_), .A1(new_n6762_), .B0(new_n6765_), .Y(new_n6766_));
  OR4X1    g06702(.A(new_n570_), .B(new_n299_), .C(new_n282_), .D(new_n155_), .Y(new_n6767_));
  OR4X1    g06703(.A(new_n1780_), .B(new_n514_), .C(new_n474_), .D(new_n177_), .Y(new_n6768_));
  OAI22X1  g06704(.A0(new_n129_), .A1(new_n119_), .B0(new_n115_), .B1(new_n99_), .Y(new_n6769_));
  OR2X1    g06705(.A(new_n6769_), .B(new_n382_), .Y(new_n6770_));
  OR2X1    g06706(.A(new_n2065_), .B(new_n130_), .Y(new_n6771_));
  OR4X1    g06707(.A(new_n6771_), .B(new_n6770_), .C(new_n6768_), .D(new_n6767_), .Y(new_n6772_));
  OR4X1    g06708(.A(new_n848_), .B(new_n547_), .C(new_n505_), .D(new_n678_), .Y(new_n6773_));
  OR4X1    g06709(.A(new_n596_), .B(new_n494_), .C(new_n256_), .D(new_n184_), .Y(new_n6774_));
  OR4X1    g06710(.A(new_n6774_), .B(new_n6773_), .C(new_n843_), .D(new_n981_), .Y(new_n6775_));
  INVX1    g06711(.A(new_n1028_), .Y(new_n6776_));
  NAND3X1  g06712(.A(new_n6776_), .B(new_n972_), .C(new_n1468_), .Y(new_n6777_));
  OR4X1    g06713(.A(new_n475_), .B(new_n358_), .C(new_n276_), .D(new_n239_), .Y(new_n6778_));
  OR4X1    g06714(.A(new_n263_), .B(new_n814_), .C(new_n825_), .D(new_n431_), .Y(new_n6779_));
  OR4X1    g06715(.A(new_n6779_), .B(new_n6778_), .C(new_n6777_), .D(new_n708_), .Y(new_n6780_));
  OR4X1    g06716(.A(new_n1962_), .B(new_n485_), .C(new_n292_), .D(new_n521_), .Y(new_n6781_));
  OR4X1    g06717(.A(new_n6781_), .B(new_n6780_), .C(new_n6775_), .D(new_n920_), .Y(new_n6782_));
  OR4X1    g06718(.A(new_n3811_), .B(new_n3760_), .C(new_n3299_), .D(new_n420_), .Y(new_n6783_));
  OR4X1    g06719(.A(new_n1223_), .B(new_n993_), .C(new_n786_), .D(new_n729_), .Y(new_n6784_));
  OR4X1    g06720(.A(new_n429_), .B(new_n418_), .C(new_n180_), .D(new_n610_), .Y(new_n6785_));
  OR4X1    g06721(.A(new_n6785_), .B(new_n1002_), .C(new_n414_), .D(new_n691_), .Y(new_n6786_));
  OR4X1    g06722(.A(new_n1540_), .B(new_n365_), .C(new_n615_), .D(new_n578_), .Y(new_n6787_));
  OR4X1    g06723(.A(new_n6787_), .B(new_n6786_), .C(new_n6784_), .D(new_n1851_), .Y(new_n6788_));
  OR4X1    g06724(.A(new_n217_), .B(new_n162_), .C(new_n338_), .D(new_n1046_), .Y(new_n6789_));
  OR4X1    g06725(.A(new_n6789_), .B(new_n766_), .C(new_n1087_), .D(new_n327_), .Y(new_n6790_));
  NOR4X1   g06726(.A(new_n6790_), .B(new_n261_), .C(new_n228_), .D(new_n207_), .Y(new_n6791_));
  NAND2X1  g06727(.A(new_n6791_), .B(new_n1155_), .Y(new_n6792_));
  OR4X1    g06728(.A(new_n6792_), .B(new_n6788_), .C(new_n3815_), .D(new_n6783_), .Y(new_n6793_));
  NOR3X1   g06729(.A(new_n6793_), .B(new_n6782_), .C(new_n6772_), .Y(new_n6794_));
  AND2X1   g06730(.A(new_n6794_), .B(new_n2237_), .Y(new_n6795_));
  INVX1    g06731(.A(new_n6795_), .Y(new_n6796_));
  NOR2X1   g06732(.A(new_n6794_), .B(new_n2237_), .Y(new_n6797_));
  INVX1    g06733(.A(new_n6797_), .Y(new_n6798_));
  AOI21X1  g06734(.A0(new_n6798_), .A1(new_n6796_), .B0(\a[23] ), .Y(new_n6799_));
  AOI21X1  g06735(.A0(new_n6796_), .A1(new_n70_), .B0(new_n6797_), .Y(new_n6800_));
  AOI21X1  g06736(.A0(new_n6800_), .A1(new_n6796_), .B0(new_n6799_), .Y(new_n6801_));
  AOI22X1  g06737(.A0(new_n2246_), .A1(new_n1884_), .B0(new_n2093_), .B1(new_n1889_), .Y(new_n6802_));
  OAI21X1  g06738(.A0(new_n2245_), .A1(new_n1879_), .B0(new_n6802_), .Y(new_n6803_));
  AOI21X1  g06739(.A0(new_n2430_), .A1(new_n407_), .B0(new_n6803_), .Y(new_n6804_));
  XOR2X1   g06740(.A(new_n6804_), .B(new_n6801_), .Y(new_n6805_));
  XOR2X1   g06741(.A(new_n6805_), .B(new_n2241_), .Y(new_n6806_));
  XOR2X1   g06742(.A(new_n6806_), .B(new_n6766_), .Y(new_n6807_));
  AOI22X1  g06743(.A0(new_n2420_), .A1(new_n2139_), .B0(new_n2185_), .B1(new_n2252_), .Y(new_n6808_));
  OAI21X1  g06744(.A0(new_n2287_), .A1(new_n2431_), .B0(new_n6808_), .Y(new_n6809_));
  AOI21X1  g06745(.A0(new_n2669_), .A1(new_n2062_), .B0(new_n6809_), .Y(new_n6810_));
  XOR2X1   g06746(.A(new_n6810_), .B(\a[29] ), .Y(new_n6811_));
  XOR2X1   g06747(.A(new_n6811_), .B(new_n6807_), .Y(new_n6812_));
  NAND2X1  g06748(.A(new_n6760_), .B(new_n6756_), .Y(new_n6813_));
  AOI21X1  g06749(.A0(new_n6761_), .A1(new_n6813_), .B0(new_n6812_), .Y(new_n6814_));
  AND2X1   g06750(.A(new_n6813_), .B(new_n6812_), .Y(new_n6815_));
  AOI21X1  g06751(.A0(new_n6815_), .A1(new_n6761_), .B0(new_n6814_), .Y(new_n6816_));
  XOR2X1   g06752(.A(new_n6816_), .B(new_n6752_), .Y(new_n6817_));
  XOR2X1   g06753(.A(new_n6817_), .B(new_n6748_), .Y(new_n6818_));
  AND2X1   g06754(.A(new_n6818_), .B(new_n6745_), .Y(new_n6819_));
  XOR2X1   g06755(.A(new_n6743_), .B(new_n6742_), .Y(new_n6820_));
  AND2X1   g06756(.A(new_n6820_), .B(new_n6745_), .Y(new_n6821_));
  XOR2X1   g06757(.A(new_n6741_), .B(new_n2887_), .Y(new_n6822_));
  AND2X1   g06758(.A(new_n6822_), .B(new_n6820_), .Y(new_n6823_));
  INVX1    g06759(.A(new_n6823_), .Y(new_n6824_));
  INVX1    g06760(.A(new_n3107_), .Y(new_n6825_));
  INVX1    g06761(.A(new_n3243_), .Y(new_n6826_));
  INVX1    g06762(.A(new_n3560_), .Y(new_n6827_));
  INVX1    g06763(.A(new_n3561_), .Y(new_n6828_));
  INVX1    g06764(.A(new_n3916_), .Y(new_n6829_));
  INVX1    g06765(.A(new_n3917_), .Y(new_n6830_));
  INVX1    g06766(.A(new_n4092_), .Y(new_n6831_));
  INVX1    g06767(.A(new_n4446_), .Y(new_n6832_));
  INVX1    g06768(.A(new_n4878_), .Y(new_n6833_));
  INVX1    g06769(.A(new_n4879_), .Y(new_n6834_));
  INVX1    g06770(.A(new_n5385_), .Y(new_n6835_));
  INVX1    g06771(.A(new_n5969_), .Y(new_n6836_));
  OR2X1    g06772(.A(new_n6292_), .B(new_n5988_), .Y(new_n6837_));
  NOR2X1   g06773(.A(new_n6303_), .B(new_n6297_), .Y(new_n6838_));
  OR2X1    g06774(.A(new_n6313_), .B(new_n6306_), .Y(new_n6839_));
  NOR2X1   g06775(.A(new_n6320_), .B(new_n6316_), .Y(new_n6840_));
  OR2X1    g06776(.A(new_n6329_), .B(new_n6323_), .Y(new_n6841_));
  NOR2X1   g06777(.A(new_n6336_), .B(new_n6332_), .Y(new_n6842_));
  NOR2X1   g06778(.A(new_n6679_), .B(new_n6339_), .Y(new_n6843_));
  AOI21X1  g06779(.A0(new_n6679_), .A1(new_n6339_), .B0(new_n6690_), .Y(new_n6844_));
  INVX1    g06780(.A(new_n6696_), .Y(new_n6845_));
  NOR3X1   g06781(.A(new_n6845_), .B(new_n6844_), .C(new_n6843_), .Y(new_n6846_));
  INVX1    g06782(.A(new_n6698_), .Y(new_n6847_));
  OAI21X1  g06783(.A0(new_n6844_), .A1(new_n6843_), .B0(new_n6845_), .Y(new_n6848_));
  OAI21X1  g06784(.A0(new_n6847_), .A1(new_n6846_), .B0(new_n6848_), .Y(new_n6849_));
  XOR2X1   g06785(.A(new_n6336_), .B(new_n6332_), .Y(new_n6850_));
  AOI21X1  g06786(.A0(new_n6850_), .A1(new_n6849_), .B0(new_n6842_), .Y(new_n6851_));
  XOR2X1   g06787(.A(new_n6329_), .B(new_n6322_), .Y(new_n6852_));
  OAI21X1  g06788(.A0(new_n6852_), .A1(new_n6851_), .B0(new_n6841_), .Y(new_n6853_));
  INVX1    g06789(.A(new_n6705_), .Y(new_n6854_));
  AOI21X1  g06790(.A0(new_n6854_), .A1(new_n6853_), .B0(new_n6840_), .Y(new_n6855_));
  OAI21X1  g06791(.A0(new_n6707_), .A1(new_n6855_), .B0(new_n6839_), .Y(new_n6856_));
  XOR2X1   g06792(.A(new_n6303_), .B(new_n6297_), .Y(new_n6857_));
  AOI21X1  g06793(.A0(new_n6857_), .A1(new_n6856_), .B0(new_n6838_), .Y(new_n6858_));
  OAI21X1  g06794(.A0(new_n6858_), .A1(new_n6294_), .B0(new_n6837_), .Y(new_n6859_));
  AOI21X1  g06795(.A0(new_n6713_), .A1(new_n6859_), .B0(new_n5985_), .Y(new_n6860_));
  INVX1    g06796(.A(new_n6716_), .Y(new_n6861_));
  OAI21X1  g06797(.A0(new_n6861_), .A1(new_n6860_), .B0(new_n6836_), .Y(new_n6862_));
  AOI21X1  g06798(.A0(new_n6862_), .A1(new_n5669_), .B0(new_n5667_), .Y(new_n6863_));
  INVX1    g06799(.A(new_n6719_), .Y(new_n6864_));
  OAI21X1  g06800(.A0(new_n6864_), .A1(new_n6863_), .B0(new_n6835_), .Y(new_n6865_));
  AOI21X1  g06801(.A0(new_n6721_), .A1(new_n6865_), .B0(new_n5115_), .Y(new_n6866_));
  OAI21X1  g06802(.A0(new_n6866_), .A1(new_n6834_), .B0(new_n6833_), .Y(new_n6867_));
  AOI21X1  g06803(.A0(new_n6867_), .A1(new_n4647_), .B0(new_n4645_), .Y(new_n6868_));
  INVX1    g06804(.A(new_n6726_), .Y(new_n6869_));
  OAI21X1  g06805(.A0(new_n6869_), .A1(new_n6868_), .B0(new_n6832_), .Y(new_n6870_));
  AOI21X1  g06806(.A0(new_n6870_), .A1(new_n4257_), .B0(new_n4255_), .Y(new_n6871_));
  INVX1    g06807(.A(new_n6729_), .Y(new_n6872_));
  OAI21X1  g06808(.A0(new_n6872_), .A1(new_n6871_), .B0(new_n6831_), .Y(new_n6873_));
  AOI21X1  g06809(.A0(new_n6731_), .A1(new_n6873_), .B0(new_n4002_), .Y(new_n6874_));
  OAI21X1  g06810(.A0(new_n6874_), .A1(new_n6830_), .B0(new_n6829_), .Y(new_n6875_));
  AOI21X1  g06811(.A0(new_n6875_), .A1(new_n3639_), .B0(new_n3637_), .Y(new_n6876_));
  OAI21X1  g06812(.A0(new_n6876_), .A1(new_n6828_), .B0(new_n6827_), .Y(new_n6877_));
  AOI21X1  g06813(.A0(new_n6877_), .A1(new_n3398_), .B0(new_n3395_), .Y(new_n6878_));
  INVX1    g06814(.A(new_n6738_), .Y(new_n6879_));
  OAI21X1  g06815(.A0(new_n6879_), .A1(new_n6878_), .B0(new_n6826_), .Y(new_n6880_));
  AOI21X1  g06816(.A0(new_n6880_), .A1(new_n3163_), .B0(new_n3161_), .Y(new_n6881_));
  XOR2X1   g06817(.A(new_n6881_), .B(new_n6825_), .Y(new_n6882_));
  AND2X1   g06818(.A(new_n6882_), .B(new_n6822_), .Y(new_n6883_));
  INVX1    g06819(.A(new_n6882_), .Y(new_n6884_));
  XOR2X1   g06820(.A(new_n6739_), .B(new_n3164_), .Y(new_n6885_));
  INVX1    g06821(.A(new_n6885_), .Y(new_n6886_));
  XOR2X1   g06822(.A(new_n6738_), .B(new_n6737_), .Y(new_n6887_));
  AND2X1   g06823(.A(new_n6887_), .B(new_n6885_), .Y(new_n6888_));
  INVX1    g06824(.A(new_n6888_), .Y(new_n6889_));
  XOR2X1   g06825(.A(new_n6736_), .B(new_n3399_), .Y(new_n6890_));
  AND2X1   g06826(.A(new_n6890_), .B(new_n6887_), .Y(new_n6891_));
  XOR2X1   g06827(.A(new_n6876_), .B(new_n6828_), .Y(new_n6892_));
  NAND2X1  g06828(.A(new_n6892_), .B(new_n6890_), .Y(new_n6893_));
  XOR2X1   g06829(.A(new_n6734_), .B(new_n3640_), .Y(new_n6894_));
  AND2X1   g06830(.A(new_n6894_), .B(new_n6892_), .Y(new_n6895_));
  INVX1    g06831(.A(new_n6894_), .Y(new_n6896_));
  XOR2X1   g06832(.A(new_n6874_), .B(new_n6830_), .Y(new_n6897_));
  INVX1    g06833(.A(new_n6897_), .Y(new_n6898_));
  XOR2X1   g06834(.A(new_n6732_), .B(new_n6730_), .Y(new_n6899_));
  AND2X1   g06835(.A(new_n6899_), .B(new_n6897_), .Y(new_n6900_));
  INVX1    g06836(.A(new_n6900_), .Y(new_n6901_));
  XOR2X1   g06837(.A(new_n6729_), .B(new_n6728_), .Y(new_n6902_));
  AND2X1   g06838(.A(new_n6902_), .B(new_n6899_), .Y(new_n6903_));
  XOR2X1   g06839(.A(new_n6727_), .B(new_n4258_), .Y(new_n6904_));
  AND2X1   g06840(.A(new_n6904_), .B(new_n6902_), .Y(new_n6905_));
  XOR2X1   g06841(.A(new_n6726_), .B(new_n6725_), .Y(new_n6906_));
  AND2X1   g06842(.A(new_n6906_), .B(new_n6904_), .Y(new_n6907_));
  INVX1    g06843(.A(new_n6907_), .Y(new_n6908_));
  XOR2X1   g06844(.A(new_n6724_), .B(new_n4648_), .Y(new_n6909_));
  AND2X1   g06845(.A(new_n6909_), .B(new_n6906_), .Y(new_n6910_));
  XOR2X1   g06846(.A(new_n6866_), .B(new_n6834_), .Y(new_n6911_));
  NAND2X1  g06847(.A(new_n6911_), .B(new_n6909_), .Y(new_n6912_));
  XOR2X1   g06848(.A(new_n6722_), .B(new_n6720_), .Y(new_n6913_));
  NAND2X1  g06849(.A(new_n6913_), .B(new_n6911_), .Y(new_n6914_));
  XOR2X1   g06850(.A(new_n6719_), .B(new_n6718_), .Y(new_n6915_));
  NAND2X1  g06851(.A(new_n6915_), .B(new_n6913_), .Y(new_n6916_));
  XOR2X1   g06852(.A(new_n6719_), .B(new_n6863_), .Y(new_n6917_));
  XOR2X1   g06853(.A(new_n6717_), .B(new_n5669_), .Y(new_n6918_));
  OR2X1    g06854(.A(new_n6918_), .B(new_n6917_), .Y(new_n6919_));
  XOR2X1   g06855(.A(new_n6716_), .B(new_n6860_), .Y(new_n6920_));
  NOR2X1   g06856(.A(new_n6920_), .B(new_n6918_), .Y(new_n6921_));
  XOR2X1   g06857(.A(new_n6861_), .B(new_n6860_), .Y(new_n6922_));
  XOR2X1   g06858(.A(new_n6713_), .B(new_n6859_), .Y(new_n6923_));
  NAND2X1  g06859(.A(new_n6923_), .B(new_n6922_), .Y(new_n6924_));
  XOR2X1   g06860(.A(new_n6858_), .B(new_n6294_), .Y(new_n6925_));
  AND2X1   g06861(.A(new_n6925_), .B(new_n6923_), .Y(new_n6926_));
  XOR2X1   g06862(.A(new_n6857_), .B(new_n6856_), .Y(new_n6927_));
  NAND2X1  g06863(.A(new_n6927_), .B(new_n6925_), .Y(new_n6928_));
  XOR2X1   g06864(.A(new_n6857_), .B(new_n6709_), .Y(new_n6929_));
  XOR2X1   g06865(.A(new_n6708_), .B(new_n6855_), .Y(new_n6930_));
  NOR2X1   g06866(.A(new_n6930_), .B(new_n6929_), .Y(new_n6931_));
  XOR2X1   g06867(.A(new_n6708_), .B(new_n6706_), .Y(new_n6932_));
  XOR2X1   g06868(.A(new_n6854_), .B(new_n6853_), .Y(new_n6933_));
  NAND2X1  g06869(.A(new_n6933_), .B(new_n6932_), .Y(new_n6934_));
  XOR2X1   g06870(.A(new_n6703_), .B(new_n6702_), .Y(new_n6935_));
  XOR2X1   g06871(.A(new_n6701_), .B(new_n6849_), .Y(new_n6936_));
  INVX1    g06872(.A(new_n6936_), .Y(new_n6937_));
  OAI21X1  g06873(.A0(new_n6937_), .A1(new_n6933_), .B0(new_n6935_), .Y(new_n6938_));
  XOR2X1   g06874(.A(new_n6933_), .B(new_n6930_), .Y(new_n6939_));
  OAI21X1  g06875(.A0(new_n6939_), .A1(new_n6938_), .B0(new_n6934_), .Y(new_n6940_));
  XOR2X1   g06876(.A(new_n6930_), .B(new_n6929_), .Y(new_n6941_));
  AOI21X1  g06877(.A0(new_n6941_), .A1(new_n6940_), .B0(new_n6931_), .Y(new_n6942_));
  NOR2X1   g06878(.A(new_n6927_), .B(new_n6925_), .Y(new_n6943_));
  OAI21X1  g06879(.A0(new_n6943_), .A1(new_n6942_), .B0(new_n6928_), .Y(new_n6944_));
  OR2X1    g06880(.A(new_n6925_), .B(new_n6923_), .Y(new_n6945_));
  AOI21X1  g06881(.A0(new_n6945_), .A1(new_n6944_), .B0(new_n6926_), .Y(new_n6946_));
  XOR2X1   g06882(.A(new_n6923_), .B(new_n6920_), .Y(new_n6947_));
  OAI21X1  g06883(.A0(new_n6947_), .A1(new_n6946_), .B0(new_n6924_), .Y(new_n6948_));
  NAND2X1  g06884(.A(new_n6920_), .B(new_n6918_), .Y(new_n6949_));
  AOI21X1  g06885(.A0(new_n6949_), .A1(new_n6948_), .B0(new_n6921_), .Y(new_n6950_));
  XOR2X1   g06886(.A(new_n6918_), .B(new_n6915_), .Y(new_n6951_));
  OAI21X1  g06887(.A0(new_n6951_), .A1(new_n6950_), .B0(new_n6919_), .Y(new_n6952_));
  XOR2X1   g06888(.A(new_n6915_), .B(new_n6913_), .Y(new_n6953_));
  NAND2X1  g06889(.A(new_n6953_), .B(new_n6952_), .Y(new_n6954_));
  AND2X1   g06890(.A(new_n6954_), .B(new_n6916_), .Y(new_n6955_));
  NOR2X1   g06891(.A(new_n6913_), .B(new_n6911_), .Y(new_n6956_));
  OAI21X1  g06892(.A0(new_n6956_), .A1(new_n6955_), .B0(new_n6914_), .Y(new_n6957_));
  XOR2X1   g06893(.A(new_n6911_), .B(new_n6909_), .Y(new_n6958_));
  NAND2X1  g06894(.A(new_n6958_), .B(new_n6957_), .Y(new_n6959_));
  INVX1    g06895(.A(new_n6909_), .Y(new_n6960_));
  XOR2X1   g06896(.A(new_n6960_), .B(new_n6906_), .Y(new_n6961_));
  AOI21X1  g06897(.A0(new_n6959_), .A1(new_n6912_), .B0(new_n6961_), .Y(new_n6962_));
  NOR2X1   g06898(.A(new_n6962_), .B(new_n6910_), .Y(new_n6963_));
  INVX1    g06899(.A(new_n6906_), .Y(new_n6964_));
  XOR2X1   g06900(.A(new_n6964_), .B(new_n6904_), .Y(new_n6965_));
  OAI21X1  g06901(.A0(new_n6965_), .A1(new_n6963_), .B0(new_n6908_), .Y(new_n6966_));
  OR2X1    g06902(.A(new_n6904_), .B(new_n6902_), .Y(new_n6967_));
  AOI21X1  g06903(.A0(new_n6967_), .A1(new_n6966_), .B0(new_n6905_), .Y(new_n6968_));
  INVX1    g06904(.A(new_n6968_), .Y(new_n6969_));
  XOR2X1   g06905(.A(new_n6902_), .B(new_n6899_), .Y(new_n6970_));
  AOI21X1  g06906(.A0(new_n6970_), .A1(new_n6969_), .B0(new_n6903_), .Y(new_n6971_));
  NOR2X1   g06907(.A(new_n6899_), .B(new_n6897_), .Y(new_n6972_));
  OAI21X1  g06908(.A0(new_n6972_), .A1(new_n6971_), .B0(new_n6901_), .Y(new_n6973_));
  XOR2X1   g06909(.A(new_n6897_), .B(new_n6894_), .Y(new_n6974_));
  NAND2X1  g06910(.A(new_n6974_), .B(new_n6973_), .Y(new_n6975_));
  OAI21X1  g06911(.A0(new_n6898_), .A1(new_n6896_), .B0(new_n6975_), .Y(new_n6976_));
  XOR2X1   g06912(.A(new_n6894_), .B(new_n6892_), .Y(new_n6977_));
  AOI21X1  g06913(.A0(new_n6977_), .A1(new_n6976_), .B0(new_n6895_), .Y(new_n6978_));
  XOR2X1   g06914(.A(new_n6892_), .B(new_n6890_), .Y(new_n6979_));
  INVX1    g06915(.A(new_n6979_), .Y(new_n6980_));
  OAI21X1  g06916(.A0(new_n6980_), .A1(new_n6978_), .B0(new_n6893_), .Y(new_n6981_));
  XOR2X1   g06917(.A(new_n6890_), .B(new_n6887_), .Y(new_n6982_));
  AOI21X1  g06918(.A0(new_n6982_), .A1(new_n6981_), .B0(new_n6891_), .Y(new_n6983_));
  NOR2X1   g06919(.A(new_n6887_), .B(new_n6885_), .Y(new_n6984_));
  OAI21X1  g06920(.A0(new_n6984_), .A1(new_n6983_), .B0(new_n6889_), .Y(new_n6985_));
  XOR2X1   g06921(.A(new_n6885_), .B(new_n6882_), .Y(new_n6986_));
  NAND2X1  g06922(.A(new_n6986_), .B(new_n6985_), .Y(new_n6987_));
  OAI21X1  g06923(.A0(new_n6886_), .A1(new_n6884_), .B0(new_n6987_), .Y(new_n6988_));
  XOR2X1   g06924(.A(new_n6882_), .B(new_n6822_), .Y(new_n6989_));
  AOI21X1  g06925(.A0(new_n6989_), .A1(new_n6988_), .B0(new_n6883_), .Y(new_n6990_));
  NOR2X1   g06926(.A(new_n6822_), .B(new_n6820_), .Y(new_n6991_));
  OAI21X1  g06927(.A0(new_n6991_), .A1(new_n6990_), .B0(new_n6824_), .Y(new_n6992_));
  XOR2X1   g06928(.A(new_n6820_), .B(new_n6745_), .Y(new_n6993_));
  AOI21X1  g06929(.A0(new_n6993_), .A1(new_n6992_), .B0(new_n6821_), .Y(new_n6994_));
  NOR2X1   g06930(.A(new_n6818_), .B(new_n6745_), .Y(new_n6995_));
  NOR3X1   g06931(.A(new_n6995_), .B(new_n6994_), .C(new_n6819_), .Y(new_n6996_));
  NOR2X1   g06932(.A(new_n6996_), .B(new_n6819_), .Y(new_n6997_));
  INVX1    g06933(.A(new_n6997_), .Y(new_n6998_));
  AND2X1   g06934(.A(new_n6816_), .B(new_n6752_), .Y(new_n6999_));
  AOI21X1  g06935(.A0(new_n6817_), .A1(new_n6748_), .B0(new_n6999_), .Y(new_n7000_));
  XOR2X1   g06936(.A(new_n6759_), .B(\a[26] ), .Y(new_n7001_));
  AOI21X1  g06937(.A0(new_n7001_), .A1(new_n6756_), .B0(new_n6814_), .Y(new_n7002_));
  INVX1    g06938(.A(new_n7002_), .Y(new_n7003_));
  AOI22X1  g06939(.A0(new_n2649_), .A1(new_n2418_), .B0(new_n2424_), .B1(new_n2421_), .Y(new_n7004_));
  OAI21X1  g06940(.A0(new_n2695_), .A1(new_n2665_), .B0(new_n7004_), .Y(new_n7005_));
  XOR2X1   g06941(.A(new_n7005_), .B(new_n89_), .Y(new_n7006_));
  AND2X1   g06942(.A(new_n6806_), .B(new_n6766_), .Y(new_n7007_));
  INVX1    g06943(.A(new_n7007_), .Y(new_n7008_));
  INVX1    g06944(.A(new_n6807_), .Y(new_n7009_));
  OAI21X1  g06945(.A0(new_n6811_), .A1(new_n7009_), .B0(new_n7008_), .Y(new_n7010_));
  INVX1    g06946(.A(new_n7010_), .Y(new_n7011_));
  AOI22X1  g06947(.A0(new_n2246_), .A1(new_n1890_), .B0(new_n2252_), .B1(new_n1889_), .Y(new_n7012_));
  OAI21X1  g06948(.A0(new_n2092_), .A1(new_n1885_), .B0(new_n7012_), .Y(new_n7013_));
  AOI21X1  g06949(.A0(new_n2201_), .A1(new_n407_), .B0(new_n7013_), .Y(new_n7014_));
  INVX1    g06950(.A(new_n1145_), .Y(new_n7015_));
  OR4X1    g06951(.A(new_n741_), .B(new_n429_), .C(new_n797_), .D(new_n144_), .Y(new_n7016_));
  OR4X1    g06952(.A(new_n226_), .B(new_n410_), .C(new_n337_), .D(new_n1579_), .Y(new_n7017_));
  OR4X1    g06953(.A(new_n2806_), .B(new_n1703_), .C(new_n1640_), .D(new_n1547_), .Y(new_n7018_));
  OR4X1    g06954(.A(new_n1347_), .B(new_n1205_), .C(new_n1978_), .D(new_n441_), .Y(new_n7019_));
  OR4X1    g06955(.A(new_n7019_), .B(new_n7018_), .C(new_n7017_), .D(new_n7016_), .Y(new_n7020_));
  OAI22X1  g06956(.A0(new_n143_), .A1(new_n88_), .B0(new_n131_), .B1(new_n69_), .Y(new_n7021_));
  OR2X1    g06957(.A(new_n7021_), .B(new_n523_), .Y(new_n7022_));
  OAI22X1  g06958(.A0(new_n131_), .A1(new_n106_), .B0(new_n105_), .B1(new_n96_), .Y(new_n7023_));
  OR4X1    g06959(.A(new_n885_), .B(new_n184_), .C(new_n175_), .D(new_n120_), .Y(new_n7024_));
  OR4X1    g06960(.A(new_n7024_), .B(new_n7023_), .C(new_n7022_), .D(new_n723_), .Y(new_n7025_));
  OR4X1    g06961(.A(new_n7025_), .B(new_n7020_), .C(new_n3450_), .D(new_n3309_), .Y(new_n7026_));
  NOR2X1   g06962(.A(new_n7026_), .B(new_n7015_), .Y(new_n7027_));
  INVX1    g06963(.A(new_n7027_), .Y(new_n7028_));
  XOR2X1   g06964(.A(new_n7028_), .B(new_n6800_), .Y(new_n7029_));
  XOR2X1   g06965(.A(new_n7029_), .B(new_n7014_), .Y(new_n7030_));
  INVX1    g06966(.A(new_n7030_), .Y(new_n7031_));
  NOR2X1   g06967(.A(new_n6804_), .B(new_n6801_), .Y(new_n7032_));
  AOI21X1  g06968(.A0(new_n6805_), .A1(new_n2241_), .B0(new_n7032_), .Y(new_n7033_));
  XOR2X1   g06969(.A(new_n7033_), .B(new_n7031_), .Y(new_n7034_));
  OAI22X1  g06970(.A0(new_n2339_), .A1(new_n2431_), .B0(new_n2287_), .B1(new_n2186_), .Y(new_n7035_));
  AOI21X1  g06971(.A0(new_n2752_), .A1(new_n2139_), .B0(new_n7035_), .Y(new_n7036_));
  OAI21X1  g06972(.A0(new_n6324_), .A1(new_n2063_), .B0(new_n7036_), .Y(new_n7037_));
  XOR2X1   g06973(.A(new_n7037_), .B(new_n74_), .Y(new_n7038_));
  XOR2X1   g06974(.A(new_n7038_), .B(new_n7034_), .Y(new_n7039_));
  XOR2X1   g06975(.A(new_n7039_), .B(new_n7011_), .Y(new_n7040_));
  XOR2X1   g06976(.A(new_n7040_), .B(new_n7006_), .Y(new_n7041_));
  XOR2X1   g06977(.A(new_n7041_), .B(new_n7003_), .Y(new_n7042_));
  INVX1    g06978(.A(new_n7042_), .Y(new_n7043_));
  XOR2X1   g06979(.A(new_n7043_), .B(new_n7000_), .Y(new_n7044_));
  XOR2X1   g06980(.A(new_n7044_), .B(new_n6818_), .Y(new_n7045_));
  XOR2X1   g06981(.A(new_n7045_), .B(new_n6998_), .Y(new_n7046_));
  INVX1    g06982(.A(new_n7044_), .Y(new_n7047_));
  AOI22X1  g06983(.A0(new_n6818_), .A1(new_n1884_), .B0(new_n6745_), .B1(new_n1890_), .Y(new_n7048_));
  OAI21X1  g06984(.A0(new_n7047_), .A1(new_n3498_), .B0(new_n7048_), .Y(new_n7049_));
  AOI21X1  g06985(.A0(new_n7046_), .A1(new_n407_), .B0(new_n7049_), .Y(new_n7050_));
  AND2X1   g06986(.A(new_n404_), .B(new_n270_), .Y(new_n7051_));
  NOR3X1   g06987(.A(new_n7051_), .B(new_n7050_), .C(new_n405_), .Y(new_n7052_));
  NOR2X1   g06988(.A(new_n7052_), .B(new_n405_), .Y(new_n7053_));
  INVX1    g06989(.A(new_n7053_), .Y(new_n7054_));
  OR4X1    g06990(.A(new_n539_), .B(new_n228_), .C(new_n757_), .D(new_n114_), .Y(new_n7055_));
  OR2X1    g06991(.A(new_n1703_), .B(new_n2065_), .Y(new_n7056_));
  OAI22X1  g06992(.A0(new_n152_), .A1(new_n108_), .B0(new_n143_), .B1(new_n69_), .Y(new_n7057_));
  OR2X1    g06993(.A(new_n7057_), .B(new_n724_), .Y(new_n7058_));
  OR4X1    g06994(.A(new_n7058_), .B(new_n848_), .C(new_n506_), .D(new_n474_), .Y(new_n7059_));
  NOR4X1   g06995(.A(new_n7059_), .B(new_n7056_), .C(new_n7055_), .D(new_n662_), .Y(new_n7060_));
  OR4X1    g06996(.A(new_n1044_), .B(new_n497_), .C(new_n825_), .D(new_n291_), .Y(new_n7061_));
  OR4X1    g06997(.A(new_n840_), .B(new_n747_), .C(new_n217_), .D(new_n120_), .Y(new_n7062_));
  NAND3X1  g06998(.A(new_n749_), .B(new_n762_), .C(new_n2149_), .Y(new_n7063_));
  OAI22X1  g06999(.A0(new_n105_), .A1(new_n115_), .B0(new_n84_), .B1(new_n72_), .Y(new_n7064_));
  OR2X1    g07000(.A(new_n7064_), .B(new_n1082_), .Y(new_n7065_));
  OR4X1    g07001(.A(new_n7065_), .B(new_n7063_), .C(new_n7062_), .D(new_n7061_), .Y(new_n7066_));
  OR4X1    g07002(.A(new_n487_), .B(new_n276_), .C(new_n144_), .D(new_n118_), .Y(new_n7067_));
  OR4X1    g07003(.A(new_n1640_), .B(new_n1006_), .C(new_n612_), .D(new_n191_), .Y(new_n7068_));
  NOR4X1   g07004(.A(new_n7068_), .B(new_n7067_), .C(new_n7066_), .D(new_n1737_), .Y(new_n7069_));
  NAND3X1  g07005(.A(new_n7069_), .B(new_n7060_), .C(new_n1170_), .Y(new_n7070_));
  OR4X1    g07006(.A(new_n1478_), .B(new_n1005_), .C(new_n475_), .D(new_n348_), .Y(new_n7071_));
  OR4X1    g07007(.A(new_n586_), .B(new_n1261_), .C(new_n245_), .D(new_n160_), .Y(new_n7072_));
  OR4X1    g07008(.A(new_n7072_), .B(new_n891_), .C(new_n740_), .D(new_n304_), .Y(new_n7073_));
  OR4X1    g07009(.A(new_n7073_), .B(new_n7071_), .C(new_n3313_), .D(new_n597_), .Y(new_n7074_));
  OAI22X1  g07010(.A0(new_n129_), .A1(new_n117_), .B0(new_n90_), .B1(new_n79_), .Y(new_n7075_));
  OR4X1    g07011(.A(new_n7075_), .B(new_n2342_), .C(new_n229_), .D(new_n207_), .Y(new_n7076_));
  OR4X1    g07012(.A(new_n246_), .B(new_n227_), .C(new_n100_), .D(new_n521_), .Y(new_n7077_));
  OR4X1    g07013(.A(new_n7077_), .B(new_n7076_), .C(new_n1141_), .D(new_n417_), .Y(new_n7078_));
  NOR3X1   g07014(.A(new_n201_), .B(new_n197_), .C(new_n610_), .Y(new_n7079_));
  NOR3X1   g07015(.A(new_n632_), .B(new_n505_), .C(new_n394_), .Y(new_n7080_));
  NOR4X1   g07016(.A(new_n998_), .B(new_n483_), .C(new_n196_), .D(new_n327_), .Y(new_n7081_));
  NAND3X1  g07017(.A(new_n7081_), .B(new_n7080_), .C(new_n7079_), .Y(new_n7082_));
  OR4X1    g07018(.A(new_n7082_), .B(new_n7078_), .C(new_n7074_), .D(new_n2814_), .Y(new_n7083_));
  OAI22X1  g07019(.A0(new_n152_), .A1(new_n81_), .B0(new_n90_), .B1(new_n84_), .Y(new_n7084_));
  OR4X1    g07020(.A(new_n636_), .B(new_n354_), .C(new_n202_), .D(new_n156_), .Y(new_n7085_));
  OR4X1    g07021(.A(new_n7085_), .B(new_n7084_), .C(new_n2468_), .D(new_n642_), .Y(new_n7086_));
  OR4X1    g07022(.A(new_n7086_), .B(new_n1172_), .C(new_n787_), .D(new_n673_), .Y(new_n7087_));
  OR4X1    g07023(.A(new_n1090_), .B(new_n945_), .C(new_n383_), .D(new_n301_), .Y(new_n7088_));
  OR4X1    g07024(.A(new_n479_), .B(new_n664_), .C(new_n1087_), .D(new_n133_), .Y(new_n7089_));
  OR4X1    g07025(.A(new_n7089_), .B(new_n7088_), .C(new_n515_), .D(new_n1467_), .Y(new_n7090_));
  NOR2X1   g07026(.A(new_n3764_), .B(new_n178_), .Y(new_n7091_));
  NAND3X1  g07027(.A(new_n7091_), .B(new_n1397_), .C(new_n855_), .Y(new_n7092_));
  OR4X1    g07028(.A(new_n7092_), .B(new_n7090_), .C(new_n3740_), .D(new_n1185_), .Y(new_n7093_));
  OR4X1    g07029(.A(new_n7093_), .B(new_n7087_), .C(new_n7083_), .D(new_n7070_), .Y(new_n7094_));
  NOR4X1   g07030(.A(new_n7094_), .B(new_n2408_), .C(new_n427_), .D(new_n365_), .Y(new_n7095_));
  INVX1    g07031(.A(new_n7095_), .Y(new_n7096_));
  OR4X1    g07032(.A(new_n1751_), .B(new_n183_), .C(new_n178_), .D(new_n164_), .Y(new_n7097_));
  OR4X1    g07033(.A(new_n7097_), .B(new_n1510_), .C(new_n873_), .D(new_n694_), .Y(new_n7098_));
  OR4X1    g07034(.A(new_n7098_), .B(new_n3007_), .C(new_n2639_), .D(new_n2392_), .Y(new_n7099_));
  NOR4X1   g07035(.A(new_n1336_), .B(new_n994_), .C(new_n391_), .D(new_n307_), .Y(new_n7100_));
  NAND3X1  g07036(.A(new_n7100_), .B(new_n2362_), .C(new_n1164_), .Y(new_n7101_));
  NOR4X1   g07037(.A(new_n7101_), .B(new_n7099_), .C(new_n2360_), .D(new_n2071_), .Y(new_n7102_));
  OR4X1    g07038(.A(new_n2070_), .B(new_n873_), .C(new_n1261_), .D(new_n327_), .Y(new_n7103_));
  OR4X1    g07039(.A(new_n2409_), .B(new_n460_), .C(new_n203_), .D(new_n103_), .Y(new_n7104_));
  NOR4X1   g07040(.A(new_n7104_), .B(new_n7103_), .C(new_n2402_), .D(new_n2365_), .Y(new_n7105_));
  AND2X1   g07041(.A(new_n7105_), .B(new_n7102_), .Y(new_n7106_));
  INVX1    g07042(.A(new_n7106_), .Y(new_n7107_));
  OR4X1    g07043(.A(new_n891_), .B(new_n386_), .C(new_n565_), .D(new_n233_), .Y(new_n7108_));
  OR4X1    g07044(.A(new_n7108_), .B(new_n802_), .C(new_n522_), .D(new_n2065_), .Y(new_n7109_));
  AOI21X1  g07045(.A0(new_n127_), .A1(new_n108_), .B0(new_n84_), .Y(new_n7110_));
  OR4X1    g07046(.A(new_n7110_), .B(new_n1608_), .C(new_n641_), .D(new_n206_), .Y(new_n7111_));
  OR4X1    g07047(.A(new_n7111_), .B(new_n7109_), .C(new_n2642_), .D(new_n2335_), .Y(new_n7112_));
  OR2X1    g07048(.A(new_n7112_), .B(new_n2394_), .Y(new_n7113_));
  AND2X1   g07049(.A(new_n7113_), .B(new_n7102_), .Y(new_n7114_));
  AOI22X1  g07050(.A0(new_n2652_), .A1(new_n407_), .B0(new_n2649_), .B1(new_n1890_), .Y(new_n7115_));
  NOR2X1   g07051(.A(new_n7113_), .B(new_n7102_), .Y(new_n7116_));
  NOR3X1   g07052(.A(new_n7116_), .B(new_n7115_), .C(new_n7114_), .Y(new_n7117_));
  NOR2X1   g07053(.A(new_n7117_), .B(new_n7114_), .Y(new_n7118_));
  XOR2X1   g07054(.A(new_n7105_), .B(new_n7102_), .Y(new_n7119_));
  NOR2X1   g07055(.A(new_n7119_), .B(new_n7118_), .Y(new_n7120_));
  INVX1    g07056(.A(new_n7120_), .Y(new_n7121_));
  INVX1    g07057(.A(new_n7118_), .Y(new_n7122_));
  XOR2X1   g07058(.A(new_n7119_), .B(new_n7122_), .Y(new_n7123_));
  OAI22X1  g07059(.A0(new_n7122_), .A1(new_n7116_), .B0(new_n7117_), .B1(new_n7115_), .Y(new_n7124_));
  INVX1    g07060(.A(new_n7124_), .Y(new_n7125_));
  INVX1    g07061(.A(new_n7102_), .Y(new_n7126_));
  OR4X1    g07062(.A(new_n1647_), .B(new_n1105_), .C(new_n156_), .D(new_n928_), .Y(new_n7127_));
  OR4X1    g07063(.A(new_n494_), .B(new_n218_), .C(new_n142_), .D(new_n338_), .Y(new_n7128_));
  OR4X1    g07064(.A(new_n387_), .B(new_n292_), .C(new_n758_), .D(new_n291_), .Y(new_n7129_));
  OR4X1    g07065(.A(new_n7129_), .B(new_n7128_), .C(new_n7127_), .D(new_n1270_), .Y(new_n7130_));
  OR4X1    g07066(.A(new_n589_), .B(new_n202_), .C(new_n196_), .D(new_n610_), .Y(new_n7131_));
  OR4X1    g07067(.A(new_n631_), .B(new_n843_), .C(new_n234_), .D(new_n981_), .Y(new_n7132_));
  AOI21X1  g07068(.A0(new_n102_), .A1(new_n91_), .B0(new_n129_), .Y(new_n7133_));
  OR2X1    g07069(.A(new_n7133_), .B(new_n1028_), .Y(new_n7134_));
  OR4X1    g07070(.A(new_n632_), .B(new_n500_), .C(new_n869_), .D(new_n301_), .Y(new_n7135_));
  OR4X1    g07071(.A(new_n7135_), .B(new_n7134_), .C(new_n7132_), .D(new_n7131_), .Y(new_n7136_));
  INVX1    g07072(.A(new_n2512_), .Y(new_n7137_));
  OR4X1    g07073(.A(new_n642_), .B(new_n1398_), .C(new_n282_), .D(new_n177_), .Y(new_n7138_));
  OR4X1    g07074(.A(new_n7138_), .B(new_n2950_), .C(new_n7137_), .D(new_n917_), .Y(new_n7139_));
  OR4X1    g07075(.A(new_n7139_), .B(new_n7136_), .C(new_n7130_), .D(new_n712_), .Y(new_n7140_));
  OR4X1    g07076(.A(new_n1757_), .B(new_n334_), .C(new_n172_), .D(new_n648_), .Y(new_n7141_));
  OR4X1    g07077(.A(new_n755_), .B(new_n547_), .C(new_n480_), .D(new_n475_), .Y(new_n7142_));
  OR4X1    g07078(.A(new_n372_), .B(new_n423_), .C(new_n819_), .D(new_n176_), .Y(new_n7143_));
  OR4X1    g07079(.A(new_n7143_), .B(new_n7142_), .C(new_n7141_), .D(new_n2066_), .Y(new_n7144_));
  OR4X1    g07080(.A(new_n7144_), .B(new_n702_), .C(new_n414_), .D(new_n200_), .Y(new_n7145_));
  NOR3X1   g07081(.A(new_n7145_), .B(new_n7140_), .C(new_n966_), .Y(new_n7146_));
  OR4X1    g07082(.A(new_n2945_), .B(new_n2319_), .C(new_n786_), .D(new_n85_), .Y(new_n7147_));
  AOI21X1  g07083(.A0(new_n96_), .A1(new_n79_), .B0(new_n125_), .Y(new_n7148_));
  OAI22X1  g07084(.A0(new_n117_), .A1(new_n90_), .B0(new_n99_), .B1(new_n91_), .Y(new_n7149_));
  OR4X1    g07085(.A(new_n1277_), .B(new_n7149_), .C(new_n896_), .D(new_n238_), .Y(new_n7150_));
  OR4X1    g07086(.A(new_n7150_), .B(new_n7148_), .C(new_n7109_), .D(new_n203_), .Y(new_n7151_));
  OR4X1    g07087(.A(new_n7151_), .B(new_n7101_), .C(new_n2349_), .D(new_n2326_), .Y(new_n7152_));
  NOR2X1   g07088(.A(new_n7152_), .B(new_n7147_), .Y(new_n7153_));
  NOR2X1   g07089(.A(new_n7153_), .B(new_n7146_), .Y(new_n7154_));
  NAND2X1  g07090(.A(new_n7153_), .B(new_n7146_), .Y(new_n7155_));
  AOI21X1  g07091(.A0(new_n7155_), .A1(new_n74_), .B0(new_n7154_), .Y(new_n7156_));
  NOR2X1   g07092(.A(new_n7156_), .B(new_n7126_), .Y(new_n7157_));
  AOI22X1  g07093(.A0(new_n2649_), .A1(new_n1884_), .B0(new_n2421_), .B1(new_n1890_), .Y(new_n7158_));
  OAI21X1  g07094(.A0(new_n2695_), .A1(new_n3178_), .B0(new_n7158_), .Y(new_n7159_));
  XOR2X1   g07095(.A(new_n7156_), .B(new_n7126_), .Y(new_n7160_));
  AOI21X1  g07096(.A0(new_n7160_), .A1(new_n7159_), .B0(new_n7157_), .Y(new_n7161_));
  NOR2X1   g07097(.A(new_n7161_), .B(new_n7125_), .Y(new_n7162_));
  XOR2X1   g07098(.A(new_n7161_), .B(new_n7125_), .Y(new_n7163_));
  XOR2X1   g07099(.A(new_n7160_), .B(new_n7159_), .Y(new_n7164_));
  INVX1    g07100(.A(new_n7164_), .Y(new_n7165_));
  NOR2X1   g07101(.A(new_n7154_), .B(\a[29] ), .Y(new_n7166_));
  AOI21X1  g07102(.A0(new_n7166_), .A1(new_n7155_), .B0(\a[29] ), .Y(new_n7167_));
  AOI21X1  g07103(.A0(new_n7156_), .A1(new_n7155_), .B0(new_n7167_), .Y(new_n7168_));
  OR4X1    g07104(.A(new_n720_), .B(new_n386_), .C(new_n348_), .D(new_n747_), .Y(new_n7169_));
  OR4X1    g07105(.A(new_n1274_), .B(new_n767_), .C(new_n361_), .D(new_n328_), .Y(new_n7170_));
  OR4X1    g07106(.A(new_n246_), .B(new_n381_), .C(new_n792_), .D(new_n80_), .Y(new_n7171_));
  OR4X1    g07107(.A(new_n7171_), .B(new_n7170_), .C(new_n537_), .D(new_n514_), .Y(new_n7172_));
  OR4X1    g07108(.A(new_n7172_), .B(new_n7169_), .C(new_n2008_), .D(new_n944_), .Y(new_n7173_));
  OR4X1    g07109(.A(new_n3305_), .B(new_n2266_), .C(new_n3780_), .D(new_n103_), .Y(new_n7174_));
  NOR4X1   g07110(.A(new_n1142_), .B(new_n647_), .C(new_n618_), .D(new_n332_), .Y(new_n7175_));
  NOR3X1   g07111(.A(new_n723_), .B(new_n408_), .C(new_n264_), .Y(new_n7176_));
  NOR4X1   g07112(.A(new_n616_), .B(new_n233_), .C(new_n291_), .D(new_n124_), .Y(new_n7177_));
  NAND3X1  g07113(.A(new_n7177_), .B(new_n7176_), .C(new_n7175_), .Y(new_n7178_));
  AOI21X1  g07114(.A0(new_n127_), .A1(new_n99_), .B0(new_n79_), .Y(new_n7179_));
  OR4X1    g07115(.A(new_n231_), .B(new_n217_), .C(new_n357_), .D(new_n137_), .Y(new_n7180_));
  OR4X1    g07116(.A(new_n393_), .B(new_n354_), .C(new_n282_), .D(new_n86_), .Y(new_n7181_));
  OR4X1    g07117(.A(new_n7181_), .B(new_n460_), .C(new_n968_), .D(new_n420_), .Y(new_n7182_));
  OR4X1    g07118(.A(new_n7182_), .B(new_n7180_), .C(new_n7179_), .D(new_n744_), .Y(new_n7183_));
  OR4X1    g07119(.A(new_n7183_), .B(new_n7178_), .C(new_n7174_), .D(new_n1872_), .Y(new_n7184_));
  NOR3X1   g07120(.A(new_n7184_), .B(new_n7173_), .C(new_n2509_), .Y(new_n7185_));
  NOR4X1   g07121(.A(new_n7185_), .B(new_n7145_), .C(new_n7140_), .D(new_n966_), .Y(new_n7186_));
  NOR3X1   g07122(.A(new_n421_), .B(new_n574_), .C(new_n86_), .Y(new_n7187_));
  NOR4X1   g07123(.A(new_n1028_), .B(new_n634_), .C(new_n372_), .D(new_n998_), .Y(new_n7188_));
  NOR4X1   g07124(.A(new_n301_), .B(new_n296_), .C(new_n398_), .D(new_n1087_), .Y(new_n7189_));
  NAND3X1  g07125(.A(new_n7189_), .B(new_n7188_), .C(new_n7187_), .Y(new_n7190_));
  OR4X1    g07126(.A(new_n2089_), .B(new_n1105_), .C(new_n509_), .D(new_n173_), .Y(new_n7191_));
  OR4X1    g07127(.A(new_n1061_), .B(new_n668_), .C(new_n513_), .D(new_n311_), .Y(new_n7192_));
  OR4X1    g07128(.A(new_n7192_), .B(new_n7191_), .C(new_n7190_), .D(new_n3472_), .Y(new_n7193_));
  OR4X1    g07129(.A(new_n459_), .B(new_n391_), .C(new_n379_), .D(new_n85_), .Y(new_n7194_));
  OR4X1    g07130(.A(new_n354_), .B(new_n474_), .C(new_n291_), .D(new_n149_), .Y(new_n7195_));
  OR4X1    g07131(.A(new_n7195_), .B(new_n7194_), .C(new_n6787_), .D(new_n2817_), .Y(new_n7196_));
  OR4X1    g07132(.A(new_n3731_), .B(new_n432_), .C(new_n1613_), .D(new_n132_), .Y(new_n7197_));
  OR4X1    g07133(.A(new_n475_), .B(new_n414_), .C(new_n293_), .D(new_n181_), .Y(new_n7198_));
  OR2X1    g07134(.A(new_n7198_), .B(new_n3464_), .Y(new_n7199_));
  OR4X1    g07135(.A(new_n1133_), .B(new_n869_), .C(new_n223_), .D(new_n522_), .Y(new_n7200_));
  OR4X1    g07136(.A(new_n1173_), .B(new_n1018_), .C(new_n382_), .D(new_n231_), .Y(new_n7201_));
  OR4X1    g07137(.A(new_n7201_), .B(new_n7200_), .C(new_n7199_), .D(new_n7197_), .Y(new_n7202_));
  NOR4X1   g07138(.A(new_n7202_), .B(new_n7196_), .C(new_n7193_), .D(new_n1767_), .Y(new_n7203_));
  NOR2X1   g07139(.A(new_n7203_), .B(new_n7027_), .Y(new_n7204_));
  AND2X1   g07140(.A(new_n7203_), .B(new_n7027_), .Y(new_n7205_));
  INVX1    g07141(.A(new_n7205_), .Y(new_n7206_));
  AOI21X1  g07142(.A0(new_n7206_), .A1(new_n89_), .B0(new_n7204_), .Y(new_n7207_));
  NOR4X1   g07143(.A(new_n7207_), .B(new_n7184_), .C(new_n7173_), .D(new_n2509_), .Y(new_n7208_));
  AOI22X1  g07144(.A0(new_n2420_), .A1(new_n1884_), .B0(new_n2627_), .B1(new_n1890_), .Y(new_n7209_));
  OAI21X1  g07145(.A0(new_n2379_), .A1(new_n3498_), .B0(new_n7209_), .Y(new_n7210_));
  AOI21X1  g07146(.A0(new_n2625_), .A1(new_n407_), .B0(new_n7210_), .Y(new_n7211_));
  INVX1    g07147(.A(new_n7211_), .Y(new_n7212_));
  INVX1    g07148(.A(new_n7207_), .Y(new_n7213_));
  XOR2X1   g07149(.A(new_n7213_), .B(new_n7185_), .Y(new_n7214_));
  AOI21X1  g07150(.A0(new_n7214_), .A1(new_n7212_), .B0(new_n7208_), .Y(new_n7215_));
  INVX1    g07151(.A(new_n7215_), .Y(new_n7216_));
  NOR4X1   g07152(.A(new_n7184_), .B(new_n7173_), .C(new_n7146_), .D(new_n2509_), .Y(new_n7217_));
  INVX1    g07153(.A(new_n7217_), .Y(new_n7218_));
  AOI21X1  g07154(.A0(new_n7218_), .A1(new_n7216_), .B0(new_n7186_), .Y(new_n7219_));
  NOR2X1   g07155(.A(new_n7219_), .B(new_n7168_), .Y(new_n7220_));
  OAI22X1  g07156(.A0(new_n2648_), .A1(new_n3498_), .B0(new_n2414_), .B1(new_n1885_), .Y(new_n7221_));
  AOI21X1  g07157(.A0(new_n2752_), .A1(new_n1890_), .B0(new_n7221_), .Y(new_n7222_));
  OAI21X1  g07158(.A0(new_n2757_), .A1(new_n3178_), .B0(new_n7222_), .Y(new_n7223_));
  XOR2X1   g07159(.A(new_n7219_), .B(new_n7168_), .Y(new_n7224_));
  AOI21X1  g07160(.A0(new_n7224_), .A1(new_n7223_), .B0(new_n7220_), .Y(new_n7225_));
  NOR2X1   g07161(.A(new_n7225_), .B(new_n7165_), .Y(new_n7226_));
  INVX1    g07162(.A(new_n7226_), .Y(new_n7227_));
  XOR2X1   g07163(.A(new_n7225_), .B(new_n7165_), .Y(new_n7228_));
  INVX1    g07164(.A(new_n7228_), .Y(new_n7229_));
  AOI22X1  g07165(.A0(new_n2652_), .A1(new_n2062_), .B0(new_n2649_), .B1(new_n2185_), .Y(new_n7230_));
  XOR2X1   g07166(.A(new_n7230_), .B(\a[29] ), .Y(new_n7231_));
  AOI22X1  g07167(.A0(new_n2421_), .A1(new_n1889_), .B0(new_n2420_), .B1(new_n1890_), .Y(new_n7232_));
  OAI21X1  g07168(.A0(new_n2379_), .A1(new_n1885_), .B0(new_n7232_), .Y(new_n7233_));
  AOI21X1  g07169(.A0(new_n2416_), .A1(new_n407_), .B0(new_n7233_), .Y(new_n7234_));
  NOR2X1   g07170(.A(new_n7234_), .B(new_n7231_), .Y(new_n7235_));
  XOR2X1   g07171(.A(new_n7234_), .B(new_n7231_), .Y(new_n7236_));
  NOR2X1   g07172(.A(new_n7217_), .B(new_n7186_), .Y(new_n7237_));
  NOR2X1   g07173(.A(new_n7237_), .B(new_n7215_), .Y(new_n7238_));
  AOI21X1  g07174(.A0(new_n7219_), .A1(new_n7218_), .B0(new_n7238_), .Y(new_n7239_));
  INVX1    g07175(.A(new_n7239_), .Y(new_n7240_));
  AOI21X1  g07176(.A0(new_n7240_), .A1(new_n7236_), .B0(new_n7235_), .Y(new_n7241_));
  INVX1    g07177(.A(new_n7241_), .Y(new_n7242_));
  XOR2X1   g07178(.A(new_n7224_), .B(new_n7223_), .Y(new_n7243_));
  AND2X1   g07179(.A(new_n7243_), .B(new_n7242_), .Y(new_n7244_));
  XOR2X1   g07180(.A(new_n7214_), .B(new_n7211_), .Y(new_n7245_));
  INVX1    g07181(.A(new_n7060_), .Y(new_n7246_));
  OR4X1    g07182(.A(new_n3457_), .B(new_n2406_), .C(new_n1256_), .D(new_n1156_), .Y(new_n7247_));
  OAI22X1  g07183(.A0(new_n127_), .A1(new_n75_), .B0(new_n108_), .B1(new_n115_), .Y(new_n7248_));
  OR2X1    g07184(.A(new_n7248_), .B(new_n1166_), .Y(new_n7249_));
  OR4X1    g07185(.A(new_n1398_), .B(new_n365_), .C(new_n355_), .D(new_n603_), .Y(new_n7250_));
  OR4X1    g07186(.A(new_n7250_), .B(new_n7249_), .C(new_n803_), .D(new_n433_), .Y(new_n7251_));
  NOR4X1   g07187(.A(new_n7251_), .B(new_n7247_), .C(new_n7083_), .D(new_n7246_), .Y(new_n7252_));
  NOR2X1   g07188(.A(new_n7252_), .B(new_n7028_), .Y(new_n7253_));
  AOI22X1  g07189(.A0(new_n2627_), .A1(new_n1889_), .B0(new_n2093_), .B1(new_n1890_), .Y(new_n7254_));
  OAI21X1  g07190(.A0(new_n2137_), .A1(new_n1885_), .B0(new_n7254_), .Y(new_n7255_));
  AOI21X1  g07191(.A0(new_n2294_), .A1(new_n407_), .B0(new_n7255_), .Y(new_n7256_));
  AND2X1   g07192(.A(new_n7252_), .B(new_n7028_), .Y(new_n7257_));
  NOR3X1   g07193(.A(new_n7257_), .B(new_n7256_), .C(new_n7253_), .Y(new_n7258_));
  NOR2X1   g07194(.A(new_n7258_), .B(new_n7253_), .Y(new_n7259_));
  INVX1    g07195(.A(new_n7204_), .Y(new_n7260_));
  AOI21X1  g07196(.A0(new_n7206_), .A1(new_n7260_), .B0(\a[26] ), .Y(new_n7261_));
  AOI21X1  g07197(.A0(new_n7207_), .A1(new_n7206_), .B0(new_n7261_), .Y(new_n7262_));
  NOR2X1   g07198(.A(new_n7262_), .B(new_n7259_), .Y(new_n7263_));
  AOI22X1  g07199(.A0(new_n2420_), .A1(new_n1889_), .B0(new_n2252_), .B1(new_n1890_), .Y(new_n7264_));
  OAI21X1  g07200(.A0(new_n2287_), .A1(new_n1885_), .B0(new_n7264_), .Y(new_n7265_));
  AOI21X1  g07201(.A0(new_n2669_), .A1(new_n407_), .B0(new_n7265_), .Y(new_n7266_));
  INVX1    g07202(.A(new_n7266_), .Y(new_n7267_));
  XOR2X1   g07203(.A(new_n7262_), .B(new_n7259_), .Y(new_n7268_));
  AOI21X1  g07204(.A0(new_n7268_), .A1(new_n7267_), .B0(new_n7263_), .Y(new_n7269_));
  NOR2X1   g07205(.A(new_n7269_), .B(new_n7245_), .Y(new_n7270_));
  INVX1    g07206(.A(new_n7270_), .Y(new_n7271_));
  XOR2X1   g07207(.A(new_n7269_), .B(new_n7245_), .Y(new_n7272_));
  INVX1    g07208(.A(new_n7272_), .Y(new_n7273_));
  AOI22X1  g07209(.A0(new_n2649_), .A1(new_n2095_), .B0(new_n2421_), .B1(new_n2185_), .Y(new_n7274_));
  OAI21X1  g07210(.A0(new_n2695_), .A1(new_n2063_), .B0(new_n7274_), .Y(new_n7275_));
  XOR2X1   g07211(.A(new_n7275_), .B(new_n74_), .Y(new_n7276_));
  OAI21X1  g07212(.A0(new_n7276_), .A1(new_n7273_), .B0(new_n7271_), .Y(new_n7277_));
  INVX1    g07213(.A(new_n7277_), .Y(new_n7278_));
  XOR2X1   g07214(.A(new_n7239_), .B(new_n7236_), .Y(new_n7279_));
  NOR2X1   g07215(.A(new_n7279_), .B(new_n7278_), .Y(new_n7280_));
  INVX1    g07216(.A(new_n7280_), .Y(new_n7281_));
  XOR2X1   g07217(.A(new_n7276_), .B(new_n7272_), .Y(new_n7282_));
  INVX1    g07218(.A(new_n7257_), .Y(new_n7283_));
  NOR2X1   g07219(.A(new_n7258_), .B(new_n7256_), .Y(new_n7284_));
  AOI21X1  g07220(.A0(new_n7259_), .A1(new_n7283_), .B0(new_n7284_), .Y(new_n7285_));
  INVX1    g07221(.A(new_n7014_), .Y(new_n7286_));
  NOR2X1   g07222(.A(new_n7028_), .B(new_n6800_), .Y(new_n7287_));
  AOI21X1  g07223(.A0(new_n7029_), .A1(new_n7286_), .B0(new_n7287_), .Y(new_n7288_));
  NOR2X1   g07224(.A(new_n7288_), .B(new_n7285_), .Y(new_n7289_));
  XOR2X1   g07225(.A(new_n7288_), .B(new_n7285_), .Y(new_n7290_));
  OR2X1    g07226(.A(new_n7033_), .B(new_n7030_), .Y(new_n7291_));
  OAI21X1  g07227(.A0(new_n7038_), .A1(new_n7034_), .B0(new_n7291_), .Y(new_n7292_));
  AOI21X1  g07228(.A0(new_n7292_), .A1(new_n7290_), .B0(new_n7289_), .Y(new_n7293_));
  XOR2X1   g07229(.A(new_n7268_), .B(new_n7266_), .Y(new_n7294_));
  NOR2X1   g07230(.A(new_n7294_), .B(new_n7293_), .Y(new_n7295_));
  XOR2X1   g07231(.A(new_n7294_), .B(new_n7293_), .Y(new_n7296_));
  AOI22X1  g07232(.A0(new_n2649_), .A1(new_n2139_), .B0(new_n2421_), .B1(new_n2095_), .Y(new_n7297_));
  OAI21X1  g07233(.A0(new_n2379_), .A1(new_n2186_), .B0(new_n7297_), .Y(new_n7298_));
  AOI21X1  g07234(.A0(new_n5957_), .A1(new_n2062_), .B0(new_n7298_), .Y(new_n7299_));
  XOR2X1   g07235(.A(new_n7299_), .B(new_n74_), .Y(new_n7300_));
  AOI21X1  g07236(.A0(new_n7300_), .A1(new_n7296_), .B0(new_n7295_), .Y(new_n7301_));
  NOR2X1   g07237(.A(new_n7301_), .B(new_n7282_), .Y(new_n7302_));
  XOR2X1   g07238(.A(new_n7301_), .B(new_n7282_), .Y(new_n7303_));
  XOR2X1   g07239(.A(new_n7300_), .B(new_n7296_), .Y(new_n7304_));
  INVX1    g07240(.A(new_n7304_), .Y(new_n7305_));
  AOI22X1  g07241(.A0(new_n2652_), .A1(new_n2301_), .B0(new_n2649_), .B1(new_n2424_), .Y(new_n7306_));
  XOR2X1   g07242(.A(new_n7306_), .B(\a[26] ), .Y(new_n7307_));
  INVX1    g07243(.A(new_n7307_), .Y(new_n7308_));
  AOI22X1  g07244(.A0(new_n2421_), .A1(new_n2139_), .B0(new_n2420_), .B1(new_n2185_), .Y(new_n7309_));
  OAI21X1  g07245(.A0(new_n2379_), .A1(new_n2431_), .B0(new_n7309_), .Y(new_n7310_));
  AOI21X1  g07246(.A0(new_n2416_), .A1(new_n2062_), .B0(new_n7310_), .Y(new_n7311_));
  XOR2X1   g07247(.A(new_n7311_), .B(new_n74_), .Y(new_n7312_));
  INVX1    g07248(.A(new_n7290_), .Y(new_n7313_));
  XOR2X1   g07249(.A(new_n7292_), .B(new_n7313_), .Y(new_n7314_));
  XOR2X1   g07250(.A(new_n7312_), .B(new_n7307_), .Y(new_n7315_));
  NOR2X1   g07251(.A(new_n7315_), .B(new_n7314_), .Y(new_n7316_));
  AOI21X1  g07252(.A0(new_n7312_), .A1(new_n7308_), .B0(new_n7316_), .Y(new_n7317_));
  NOR2X1   g07253(.A(new_n7317_), .B(new_n7305_), .Y(new_n7318_));
  INVX1    g07254(.A(new_n7318_), .Y(new_n7319_));
  XOR2X1   g07255(.A(new_n7317_), .B(new_n7304_), .Y(new_n7320_));
  AND2X1   g07256(.A(new_n7039_), .B(new_n7010_), .Y(new_n7321_));
  INVX1    g07257(.A(new_n7321_), .Y(new_n7322_));
  OAI21X1  g07258(.A0(new_n7040_), .A1(new_n7006_), .B0(new_n7322_), .Y(new_n7323_));
  XOR2X1   g07259(.A(new_n7315_), .B(new_n7314_), .Y(new_n7324_));
  AND2X1   g07260(.A(new_n7324_), .B(new_n7323_), .Y(new_n7325_));
  AND2X1   g07261(.A(new_n7041_), .B(new_n7003_), .Y(new_n7326_));
  INVX1    g07262(.A(new_n7326_), .Y(new_n7327_));
  OAI21X1  g07263(.A0(new_n7043_), .A1(new_n7000_), .B0(new_n7327_), .Y(new_n7328_));
  XOR2X1   g07264(.A(new_n7324_), .B(new_n7323_), .Y(new_n7329_));
  AOI21X1  g07265(.A0(new_n7329_), .A1(new_n7328_), .B0(new_n7325_), .Y(new_n7330_));
  OAI21X1  g07266(.A0(new_n7330_), .A1(new_n7320_), .B0(new_n7319_), .Y(new_n7331_));
  AOI21X1  g07267(.A0(new_n7331_), .A1(new_n7303_), .B0(new_n7302_), .Y(new_n7332_));
  XOR2X1   g07268(.A(new_n7279_), .B(new_n7278_), .Y(new_n7333_));
  INVX1    g07269(.A(new_n7333_), .Y(new_n7334_));
  OAI21X1  g07270(.A0(new_n7334_), .A1(new_n7332_), .B0(new_n7281_), .Y(new_n7335_));
  XOR2X1   g07271(.A(new_n7243_), .B(new_n7242_), .Y(new_n7336_));
  AOI21X1  g07272(.A0(new_n7336_), .A1(new_n7335_), .B0(new_n7244_), .Y(new_n7337_));
  OAI21X1  g07273(.A0(new_n7337_), .A1(new_n7229_), .B0(new_n7227_), .Y(new_n7338_));
  AOI21X1  g07274(.A0(new_n7338_), .A1(new_n7163_), .B0(new_n7162_), .Y(new_n7339_));
  OAI21X1  g07275(.A0(new_n7339_), .A1(new_n7123_), .B0(new_n7121_), .Y(new_n7340_));
  NAND3X1  g07276(.A(new_n7340_), .B(new_n7107_), .C(new_n7096_), .Y(new_n7341_));
  NAND3X1  g07277(.A(new_n2874_), .B(new_n2872_), .C(new_n2869_), .Y(new_n7342_));
  AND2X1   g07278(.A(new_n7342_), .B(new_n7341_), .Y(new_n7343_));
  XOR2X1   g07279(.A(new_n7343_), .B(new_n1920_), .Y(new_n7344_));
  OAI22X1  g07280(.A0(new_n161_), .A1(new_n119_), .B0(new_n125_), .B1(new_n106_), .Y(new_n7345_));
  OR4X1    g07281(.A(new_n2920_), .B(new_n7345_), .C(new_n454_), .D(new_n87_), .Y(new_n7346_));
  OR4X1    g07282(.A(new_n292_), .B(new_n399_), .C(new_n757_), .D(new_n291_), .Y(new_n7347_));
  OR4X1    g07283(.A(new_n7347_), .B(new_n488_), .C(new_n218_), .D(new_n202_), .Y(new_n7348_));
  OR4X1    g07284(.A(new_n7348_), .B(new_n1398_), .C(new_n475_), .D(new_n627_), .Y(new_n7349_));
  OR4X1    g07285(.A(new_n7349_), .B(new_n7346_), .C(new_n2127_), .D(new_n1052_), .Y(new_n7350_));
  OR4X1    g07286(.A(new_n483_), .B(new_n329_), .C(new_n243_), .D(new_n159_), .Y(new_n7351_));
  OR2X1    g07287(.A(new_n569_), .B(new_n259_), .Y(new_n7352_));
  OR4X1    g07288(.A(new_n7352_), .B(new_n361_), .C(new_n358_), .D(new_n819_), .Y(new_n7353_));
  OR4X1    g07289(.A(new_n7353_), .B(new_n7351_), .C(new_n657_), .D(new_n552_), .Y(new_n7354_));
  OR4X1    g07290(.A(new_n7354_), .B(new_n830_), .C(new_n751_), .D(new_n669_), .Y(new_n7355_));
  OR2X1    g07291(.A(new_n1772_), .B(new_n866_), .Y(new_n7356_));
  NOR4X1   g07292(.A(new_n7356_), .B(new_n7355_), .C(new_n7350_), .D(new_n1258_), .Y(new_n7357_));
  XOR2X1   g07293(.A(new_n7357_), .B(new_n269_), .Y(new_n7358_));
  XOR2X1   g07294(.A(new_n7358_), .B(new_n7344_), .Y(new_n7359_));
  XOR2X1   g07295(.A(new_n7359_), .B(new_n7054_), .Y(new_n7360_));
  INVX1    g07296(.A(new_n6818_), .Y(new_n7361_));
  OAI21X1  g07297(.A0(new_n6996_), .A1(new_n6819_), .B0(new_n7045_), .Y(new_n7362_));
  OAI21X1  g07298(.A0(new_n7047_), .A1(new_n7361_), .B0(new_n7362_), .Y(new_n7363_));
  XOR2X1   g07299(.A(new_n7329_), .B(new_n7328_), .Y(new_n7364_));
  XOR2X1   g07300(.A(new_n7364_), .B(new_n7044_), .Y(new_n7365_));
  XOR2X1   g07301(.A(new_n7365_), .B(new_n7363_), .Y(new_n7366_));
  INVX1    g07302(.A(new_n7364_), .Y(new_n7367_));
  AOI22X1  g07303(.A0(new_n7044_), .A1(new_n1884_), .B0(new_n6818_), .B1(new_n1890_), .Y(new_n7368_));
  OAI21X1  g07304(.A0(new_n7367_), .A1(new_n3498_), .B0(new_n7368_), .Y(new_n7369_));
  AOI21X1  g07305(.A0(new_n7366_), .A1(new_n407_), .B0(new_n7369_), .Y(new_n7370_));
  XOR2X1   g07306(.A(new_n7370_), .B(new_n7360_), .Y(new_n7371_));
  OAI22X1  g07307(.A0(new_n7054_), .A1(new_n7051_), .B0(new_n7052_), .B1(new_n7050_), .Y(new_n7372_));
  INVX1    g07308(.A(new_n7372_), .Y(new_n7373_));
  OR4X1    g07309(.A(new_n361_), .B(new_n354_), .C(new_n208_), .D(new_n155_), .Y(new_n7374_));
  OR4X1    g07310(.A(new_n7374_), .B(new_n1777_), .C(new_n338_), .D(new_n124_), .Y(new_n7375_));
  OAI22X1  g07311(.A0(new_n117_), .A1(new_n81_), .B0(new_n106_), .B1(new_n78_), .Y(new_n7376_));
  OR4X1    g07312(.A(new_n7376_), .B(new_n2806_), .C(new_n1647_), .D(new_n1493_), .Y(new_n7377_));
  OR4X1    g07313(.A(new_n616_), .B(new_n172_), .C(new_n648_), .D(new_n746_), .Y(new_n7378_));
  OR2X1    g07314(.A(new_n1306_), .B(new_n271_), .Y(new_n7379_));
  OR4X1    g07315(.A(new_n7379_), .B(new_n7378_), .C(new_n7377_), .D(new_n7375_), .Y(new_n7380_));
  OR4X1    g07316(.A(new_n636_), .B(new_n523_), .C(new_n678_), .D(new_n426_), .Y(new_n7381_));
  OR4X1    g07317(.A(new_n7381_), .B(new_n3027_), .C(new_n1627_), .D(new_n1077_), .Y(new_n7382_));
  NOR4X1   g07318(.A(new_n7382_), .B(new_n7380_), .C(new_n1937_), .D(new_n1583_), .Y(new_n7383_));
  NAND3X1  g07319(.A(new_n258_), .B(new_n253_), .C(new_n248_), .Y(new_n7384_));
  NOR3X1   g07320(.A(new_n560_), .B(new_n758_), .C(new_n664_), .Y(new_n7385_));
  NOR4X1   g07321(.A(new_n636_), .B(new_n323_), .C(new_n293_), .D(new_n286_), .Y(new_n7386_));
  NAND3X1  g07322(.A(new_n7386_), .B(new_n7385_), .C(new_n3761_), .Y(new_n7387_));
  OR4X1    g07323(.A(new_n1224_), .B(new_n1100_), .C(new_n417_), .D(new_n1613_), .Y(new_n7388_));
  OR4X1    g07324(.A(new_n598_), .B(new_n191_), .C(new_n181_), .D(new_n175_), .Y(new_n7389_));
  OR4X1    g07325(.A(new_n7389_), .B(new_n7388_), .C(new_n582_), .D(new_n843_), .Y(new_n7390_));
  OR4X1    g07326(.A(new_n7390_), .B(new_n7387_), .C(new_n7384_), .D(new_n122_), .Y(new_n7391_));
  NOR3X1   g07327(.A(new_n7391_), .B(new_n7145_), .C(new_n2821_), .Y(new_n7392_));
  NOR2X1   g07328(.A(new_n7392_), .B(new_n7383_), .Y(new_n7393_));
  NAND3X1  g07329(.A(new_n3230_), .B(new_n3229_), .C(new_n3233_), .Y(new_n7394_));
  AND2X1   g07330(.A(new_n7394_), .B(new_n7341_), .Y(new_n7395_));
  XOR2X1   g07331(.A(new_n7395_), .B(new_n2445_), .Y(new_n7396_));
  XOR2X1   g07332(.A(new_n7392_), .B(new_n7383_), .Y(new_n7397_));
  AOI21X1  g07333(.A0(new_n7397_), .A1(new_n7396_), .B0(new_n7393_), .Y(new_n7398_));
  OR2X1    g07334(.A(new_n7398_), .B(new_n270_), .Y(new_n7399_));
  XOR2X1   g07335(.A(new_n7398_), .B(new_n269_), .Y(new_n7400_));
  NOR2X1   g07336(.A(new_n6996_), .B(new_n6994_), .Y(new_n7401_));
  NOR3X1   g07337(.A(new_n6996_), .B(new_n6995_), .C(new_n6819_), .Y(new_n7402_));
  NOR2X1   g07338(.A(new_n7402_), .B(new_n7401_), .Y(new_n7403_));
  INVX1    g07339(.A(new_n7403_), .Y(new_n7404_));
  AOI22X1  g07340(.A0(new_n6820_), .A1(new_n1890_), .B0(new_n6745_), .B1(new_n1884_), .Y(new_n7405_));
  OAI21X1  g07341(.A0(new_n7361_), .A1(new_n3498_), .B0(new_n7405_), .Y(new_n7406_));
  AOI21X1  g07342(.A0(new_n7404_), .A1(new_n407_), .B0(new_n7406_), .Y(new_n7407_));
  OR2X1    g07343(.A(new_n7407_), .B(new_n7400_), .Y(new_n7408_));
  AND2X1   g07344(.A(new_n7408_), .B(new_n7399_), .Y(new_n7409_));
  NOR2X1   g07345(.A(new_n7409_), .B(new_n7373_), .Y(new_n7410_));
  XOR2X1   g07346(.A(new_n7409_), .B(new_n7373_), .Y(new_n7411_));
  INVX1    g07347(.A(new_n6993_), .Y(new_n7412_));
  AND2X1   g07348(.A(new_n7412_), .B(new_n6992_), .Y(new_n7413_));
  NOR2X1   g07349(.A(new_n6820_), .B(new_n6745_), .Y(new_n7414_));
  NOR3X1   g07350(.A(new_n7414_), .B(new_n6992_), .C(new_n6821_), .Y(new_n7415_));
  NOR2X1   g07351(.A(new_n7415_), .B(new_n7413_), .Y(new_n7416_));
  INVX1    g07352(.A(new_n7416_), .Y(new_n7417_));
  INVX1    g07353(.A(new_n6745_), .Y(new_n7418_));
  AOI22X1  g07354(.A0(new_n6822_), .A1(new_n1890_), .B0(new_n6820_), .B1(new_n1884_), .Y(new_n7419_));
  OAI21X1  g07355(.A0(new_n7418_), .A1(new_n3498_), .B0(new_n7419_), .Y(new_n7420_));
  AOI21X1  g07356(.A0(new_n7417_), .A1(new_n407_), .B0(new_n7420_), .Y(new_n7421_));
  INVX1    g07357(.A(new_n7421_), .Y(new_n7422_));
  XOR2X1   g07358(.A(new_n7397_), .B(new_n7396_), .Y(new_n7423_));
  AND2X1   g07359(.A(new_n7423_), .B(new_n7422_), .Y(new_n7424_));
  OAI22X1  g07360(.A0(new_n88_), .A1(new_n72_), .B0(new_n84_), .B1(new_n81_), .Y(new_n7425_));
  NOR3X1   g07361(.A(new_n7425_), .B(new_n3283_), .C(new_n1105_), .Y(new_n7426_));
  NOR4X1   g07362(.A(new_n475_), .B(new_n299_), .C(new_n273_), .D(new_n194_), .Y(new_n7427_));
  NOR4X1   g07363(.A(new_n493_), .B(new_n229_), .C(new_n217_), .D(new_n116_), .Y(new_n7428_));
  NAND3X1  g07364(.A(new_n7428_), .B(new_n7427_), .C(new_n7426_), .Y(new_n7429_));
  INVX1    g07365(.A(new_n681_), .Y(new_n7430_));
  NOR4X1   g07366(.A(new_n1028_), .B(new_n720_), .C(new_n546_), .D(new_n280_), .Y(new_n7431_));
  NAND3X1  g07367(.A(new_n7431_), .B(new_n7430_), .C(new_n1933_), .Y(new_n7432_));
  OR4X1    g07368(.A(new_n7432_), .B(new_n7429_), .C(new_n3433_), .D(new_n2551_), .Y(new_n7433_));
  NOR4X1   g07369(.A(new_n7433_), .B(new_n998_), .C(new_n478_), .D(new_n147_), .Y(new_n7434_));
  NOR4X1   g07370(.A(new_n1756_), .B(new_n993_), .C(new_n487_), .D(new_n132_), .Y(new_n7435_));
  NOR3X1   g07371(.A(new_n527_), .B(new_n740_), .C(new_n539_), .Y(new_n7436_));
  NOR4X1   g07372(.A(new_n196_), .B(new_n172_), .C(new_n139_), .D(new_n1579_), .Y(new_n7437_));
  NAND3X1  g07373(.A(new_n7437_), .B(new_n7436_), .C(new_n7435_), .Y(new_n7438_));
  NAND3X1  g07374(.A(new_n1130_), .B(new_n320_), .C(new_n762_), .Y(new_n7439_));
  OR4X1    g07375(.A(new_n399_), .B(new_n203_), .C(new_n758_), .D(new_n757_), .Y(new_n7440_));
  OR4X1    g07376(.A(new_n7440_), .B(new_n7439_), .C(new_n1371_), .D(new_n1027_), .Y(new_n7441_));
  OR4X1    g07377(.A(new_n1639_), .B(new_n1224_), .C(new_n433_), .D(new_n340_), .Y(new_n7442_));
  OR2X1    g07378(.A(new_n7442_), .B(new_n3307_), .Y(new_n7443_));
  NOR4X1   g07379(.A(new_n7443_), .B(new_n7441_), .C(new_n7438_), .D(new_n1748_), .Y(new_n7444_));
  AND2X1   g07380(.A(new_n7444_), .B(new_n7434_), .Y(new_n7445_));
  INVX1    g07381(.A(new_n7445_), .Y(new_n7446_));
  AND2X1   g07382(.A(new_n7446_), .B(new_n7383_), .Y(new_n7447_));
  INVX1    g07383(.A(new_n7447_), .Y(new_n7448_));
  OAI22X1  g07384(.A0(new_n148_), .A1(new_n131_), .B0(new_n127_), .B1(new_n115_), .Y(new_n7449_));
  OR2X1    g07385(.A(new_n7449_), .B(new_n2947_), .Y(new_n7450_));
  OAI22X1  g07386(.A0(new_n108_), .A1(new_n84_), .B0(new_n106_), .B1(new_n105_), .Y(new_n7451_));
  OR4X1    g07387(.A(new_n7451_), .B(new_n2561_), .C(new_n1910_), .D(new_n795_), .Y(new_n7452_));
  OR4X1    g07388(.A(new_n869_), .B(new_n421_), .C(new_n681_), .D(new_n263_), .Y(new_n7453_));
  OR4X1    g07389(.A(new_n7453_), .B(new_n7452_), .C(new_n3030_), .D(new_n937_), .Y(new_n7454_));
  NOR4X1   g07390(.A(new_n7454_), .B(new_n7450_), .C(new_n2171_), .D(new_n1729_), .Y(new_n7455_));
  OR4X1    g07391(.A(new_n565_), .B(new_n479_), .C(new_n240_), .D(new_n327_), .Y(new_n7456_));
  OR4X1    g07392(.A(new_n420_), .B(new_n478_), .C(new_n300_), .D(new_n141_), .Y(new_n7457_));
  OR4X1    g07393(.A(new_n7457_), .B(new_n1903_), .C(new_n1105_), .D(new_n561_), .Y(new_n7458_));
  OR4X1    g07394(.A(new_n7458_), .B(new_n7456_), .C(new_n2591_), .D(new_n525_), .Y(new_n7459_));
  OR4X1    g07395(.A(new_n2540_), .B(new_n509_), .C(new_n475_), .D(new_n574_), .Y(new_n7460_));
  OR4X1    g07396(.A(new_n7460_), .B(new_n1300_), .C(new_n2097_), .D(new_n772_), .Y(new_n7461_));
  NOR4X1   g07397(.A(new_n7461_), .B(new_n7459_), .C(new_n3695_), .D(new_n1318_), .Y(new_n7462_));
  NOR2X1   g07398(.A(new_n7462_), .B(new_n7455_), .Y(new_n7463_));
  NAND3X1  g07399(.A(new_n3626_), .B(new_n3623_), .C(new_n3621_), .Y(new_n7464_));
  AND2X1   g07400(.A(new_n7464_), .B(new_n7341_), .Y(new_n7465_));
  XOR2X1   g07401(.A(new_n7465_), .B(new_n2529_), .Y(new_n7466_));
  XOR2X1   g07402(.A(new_n7462_), .B(new_n7455_), .Y(new_n7467_));
  AOI21X1  g07403(.A0(new_n7467_), .A1(new_n7466_), .B0(new_n7463_), .Y(new_n7468_));
  NOR2X1   g07404(.A(new_n7468_), .B(new_n7446_), .Y(new_n7469_));
  XOR2X1   g07405(.A(new_n7468_), .B(new_n7445_), .Y(new_n7470_));
  XOR2X1   g07406(.A(new_n6989_), .B(new_n6988_), .Y(new_n7471_));
  INVX1    g07407(.A(new_n6822_), .Y(new_n7472_));
  AOI22X1  g07408(.A0(new_n6885_), .A1(new_n1890_), .B0(new_n6882_), .B1(new_n1884_), .Y(new_n7473_));
  OAI21X1  g07409(.A0(new_n7472_), .A1(new_n3498_), .B0(new_n7473_), .Y(new_n7474_));
  AOI21X1  g07410(.A0(new_n7471_), .A1(new_n407_), .B0(new_n7474_), .Y(new_n7475_));
  NOR2X1   g07411(.A(new_n7475_), .B(new_n7470_), .Y(new_n7476_));
  XOR2X1   g07412(.A(new_n7446_), .B(new_n7383_), .Y(new_n7477_));
  OAI21X1  g07413(.A0(new_n7476_), .A1(new_n7469_), .B0(new_n7477_), .Y(new_n7478_));
  XOR2X1   g07414(.A(new_n7423_), .B(new_n7421_), .Y(new_n7479_));
  AOI21X1  g07415(.A0(new_n7478_), .A1(new_n7448_), .B0(new_n7479_), .Y(new_n7480_));
  XOR2X1   g07416(.A(new_n7407_), .B(new_n7400_), .Y(new_n7481_));
  OAI21X1  g07417(.A0(new_n7480_), .A1(new_n7424_), .B0(new_n7481_), .Y(new_n7482_));
  NOR2X1   g07418(.A(new_n7480_), .B(new_n7424_), .Y(new_n7483_));
  XOR2X1   g07419(.A(new_n7481_), .B(new_n7483_), .Y(new_n7484_));
  XOR2X1   g07420(.A(new_n7330_), .B(new_n7320_), .Y(new_n7485_));
  OAI22X1  g07421(.A0(new_n7367_), .A1(new_n2431_), .B0(new_n7047_), .B1(new_n2186_), .Y(new_n7486_));
  AOI21X1  g07422(.A0(new_n7485_), .A1(new_n2139_), .B0(new_n7486_), .Y(new_n7487_));
  AND2X1   g07423(.A(new_n7364_), .B(new_n7044_), .Y(new_n7488_));
  AOI21X1  g07424(.A0(new_n7365_), .A1(new_n7363_), .B0(new_n7488_), .Y(new_n7489_));
  AND2X1   g07425(.A(new_n7485_), .B(new_n7364_), .Y(new_n7490_));
  NOR2X1   g07426(.A(new_n7485_), .B(new_n7364_), .Y(new_n7491_));
  NOR3X1   g07427(.A(new_n7491_), .B(new_n7490_), .C(new_n7489_), .Y(new_n7492_));
  NOR2X1   g07428(.A(new_n7492_), .B(new_n7489_), .Y(new_n7493_));
  NOR3X1   g07429(.A(new_n7492_), .B(new_n7491_), .C(new_n7490_), .Y(new_n7494_));
  NOR2X1   g07430(.A(new_n7494_), .B(new_n7493_), .Y(new_n7495_));
  OAI21X1  g07431(.A0(new_n7495_), .A1(new_n2063_), .B0(new_n7487_), .Y(new_n7496_));
  XOR2X1   g07432(.A(new_n7496_), .B(new_n74_), .Y(new_n7497_));
  OAI21X1  g07433(.A0(new_n7497_), .A1(new_n7484_), .B0(new_n7482_), .Y(new_n7498_));
  AOI21X1  g07434(.A0(new_n7498_), .A1(new_n7411_), .B0(new_n7410_), .Y(new_n7499_));
  NOR2X1   g07435(.A(new_n7499_), .B(new_n7371_), .Y(new_n7500_));
  INVX1    g07436(.A(new_n7500_), .Y(new_n7501_));
  XOR2X1   g07437(.A(new_n7499_), .B(new_n7371_), .Y(new_n7502_));
  INVX1    g07438(.A(new_n7502_), .Y(new_n7503_));
  INVX1    g07439(.A(new_n7485_), .Y(new_n7504_));
  INVX1    g07440(.A(new_n7303_), .Y(new_n7505_));
  INVX1    g07441(.A(new_n7320_), .Y(new_n7506_));
  INVX1    g07442(.A(new_n7325_), .Y(new_n7507_));
  INVX1    g07443(.A(new_n2768_), .Y(new_n7508_));
  INVX1    g07444(.A(new_n3104_), .Y(new_n7509_));
  OAI21X1  g07445(.A0(new_n6881_), .A1(new_n6825_), .B0(new_n7509_), .Y(new_n7510_));
  AOI21X1  g07446(.A0(new_n7510_), .A1(new_n2886_), .B0(new_n2884_), .Y(new_n7511_));
  INVX1    g07447(.A(new_n6743_), .Y(new_n7512_));
  OAI21X1  g07448(.A0(new_n7512_), .A1(new_n7511_), .B0(new_n7508_), .Y(new_n7513_));
  AOI21X1  g07449(.A0(new_n7513_), .A1(new_n2702_), .B0(new_n6746_), .Y(new_n7514_));
  INVX1    g07450(.A(new_n6999_), .Y(new_n7515_));
  INVX1    g07451(.A(new_n6817_), .Y(new_n7516_));
  OAI21X1  g07452(.A0(new_n7516_), .A1(new_n7514_), .B0(new_n7515_), .Y(new_n7517_));
  AOI21X1  g07453(.A0(new_n7042_), .A1(new_n7517_), .B0(new_n7326_), .Y(new_n7518_));
  INVX1    g07454(.A(new_n7329_), .Y(new_n7519_));
  OAI21X1  g07455(.A0(new_n7519_), .A1(new_n7518_), .B0(new_n7507_), .Y(new_n7520_));
  AOI21X1  g07456(.A0(new_n7520_), .A1(new_n7506_), .B0(new_n7318_), .Y(new_n7521_));
  XOR2X1   g07457(.A(new_n7521_), .B(new_n7505_), .Y(new_n7522_));
  INVX1    g07458(.A(new_n7522_), .Y(new_n7523_));
  XOR2X1   g07459(.A(new_n7522_), .B(new_n7485_), .Y(new_n7524_));
  OAI21X1  g07460(.A0(new_n7492_), .A1(new_n7490_), .B0(new_n7524_), .Y(new_n7525_));
  OAI21X1  g07461(.A0(new_n7523_), .A1(new_n7504_), .B0(new_n7525_), .Y(new_n7526_));
  INVX1    g07462(.A(new_n7302_), .Y(new_n7527_));
  OAI21X1  g07463(.A0(new_n7521_), .A1(new_n7505_), .B0(new_n7527_), .Y(new_n7528_));
  XOR2X1   g07464(.A(new_n7333_), .B(new_n7528_), .Y(new_n7529_));
  XOR2X1   g07465(.A(new_n7529_), .B(new_n7523_), .Y(new_n7530_));
  AND2X1   g07466(.A(new_n7530_), .B(new_n7526_), .Y(new_n7531_));
  AND2X1   g07467(.A(new_n7529_), .B(new_n7522_), .Y(new_n7532_));
  NOR2X1   g07468(.A(new_n7529_), .B(new_n7522_), .Y(new_n7533_));
  NOR3X1   g07469(.A(new_n7533_), .B(new_n7532_), .C(new_n7526_), .Y(new_n7534_));
  NOR2X1   g07470(.A(new_n7534_), .B(new_n7531_), .Y(new_n7535_));
  INVX1    g07471(.A(new_n7535_), .Y(new_n7536_));
  INVX1    g07472(.A(new_n7529_), .Y(new_n7537_));
  AOI22X1  g07473(.A0(new_n7522_), .A1(new_n2095_), .B0(new_n7485_), .B1(new_n2185_), .Y(new_n7538_));
  OAI21X1  g07474(.A0(new_n7537_), .A1(new_n2140_), .B0(new_n7538_), .Y(new_n7539_));
  AOI21X1  g07475(.A0(new_n7536_), .A1(new_n2062_), .B0(new_n7539_), .Y(new_n7540_));
  XOR2X1   g07476(.A(new_n7540_), .B(\a[29] ), .Y(new_n7541_));
  OAI21X1  g07477(.A0(new_n7541_), .A1(new_n7503_), .B0(new_n7501_), .Y(new_n7542_));
  AND2X1   g07478(.A(new_n7359_), .B(new_n7054_), .Y(new_n7543_));
  INVX1    g07479(.A(new_n7543_), .Y(new_n7544_));
  INVX1    g07480(.A(new_n7360_), .Y(new_n7545_));
  OAI21X1  g07481(.A0(new_n7370_), .A1(new_n7545_), .B0(new_n7544_), .Y(new_n7546_));
  INVX1    g07482(.A(new_n7546_), .Y(new_n7547_));
  INVX1    g07483(.A(new_n7070_), .Y(new_n7548_));
  NOR2X1   g07484(.A(new_n7357_), .B(new_n269_), .Y(new_n7549_));
  AOI21X1  g07485(.A0(new_n7358_), .A1(new_n7344_), .B0(new_n7549_), .Y(new_n7550_));
  XOR2X1   g07486(.A(new_n7550_), .B(new_n7548_), .Y(new_n7551_));
  INVX1    g07487(.A(new_n7495_), .Y(new_n7552_));
  AOI22X1  g07488(.A0(new_n7364_), .A1(new_n1884_), .B0(new_n7044_), .B1(new_n1890_), .Y(new_n7553_));
  OAI21X1  g07489(.A0(new_n7504_), .A1(new_n3498_), .B0(new_n7553_), .Y(new_n7554_));
  AOI21X1  g07490(.A0(new_n7552_), .A1(new_n407_), .B0(new_n7554_), .Y(new_n7555_));
  XOR2X1   g07491(.A(new_n7555_), .B(new_n7551_), .Y(new_n7556_));
  XOR2X1   g07492(.A(new_n7556_), .B(new_n7547_), .Y(new_n7557_));
  XOR2X1   g07493(.A(new_n7336_), .B(new_n7335_), .Y(new_n7558_));
  OAI22X1  g07494(.A0(new_n7537_), .A1(new_n2431_), .B0(new_n7523_), .B1(new_n2186_), .Y(new_n7559_));
  AOI21X1  g07495(.A0(new_n7558_), .A1(new_n2139_), .B0(new_n7559_), .Y(new_n7560_));
  INVX1    g07496(.A(new_n7533_), .Y(new_n7561_));
  AOI21X1  g07497(.A0(new_n7561_), .A1(new_n7526_), .B0(new_n7532_), .Y(new_n7562_));
  XOR2X1   g07498(.A(new_n7558_), .B(new_n7529_), .Y(new_n7563_));
  INVX1    g07499(.A(new_n7563_), .Y(new_n7564_));
  XOR2X1   g07500(.A(new_n7564_), .B(new_n7562_), .Y(new_n7565_));
  INVX1    g07501(.A(new_n7565_), .Y(new_n7566_));
  OAI21X1  g07502(.A0(new_n7566_), .A1(new_n2063_), .B0(new_n7560_), .Y(new_n7567_));
  XOR2X1   g07503(.A(new_n7567_), .B(new_n74_), .Y(new_n7568_));
  XOR2X1   g07504(.A(new_n7568_), .B(new_n7557_), .Y(new_n7569_));
  XOR2X1   g07505(.A(new_n7569_), .B(new_n7542_), .Y(new_n7570_));
  XOR2X1   g07506(.A(new_n7337_), .B(new_n7229_), .Y(new_n7571_));
  INVX1    g07507(.A(new_n7163_), .Y(new_n7572_));
  INVX1    g07508(.A(new_n7244_), .Y(new_n7573_));
  AOI21X1  g07509(.A0(new_n7333_), .A1(new_n7528_), .B0(new_n7280_), .Y(new_n7574_));
  INVX1    g07510(.A(new_n7336_), .Y(new_n7575_));
  OAI21X1  g07511(.A0(new_n7575_), .A1(new_n7574_), .B0(new_n7573_), .Y(new_n7576_));
  AOI21X1  g07512(.A0(new_n7576_), .A1(new_n7228_), .B0(new_n7226_), .Y(new_n7577_));
  XOR2X1   g07513(.A(new_n7577_), .B(new_n7572_), .Y(new_n7578_));
  AND2X1   g07514(.A(new_n7578_), .B(new_n7571_), .Y(new_n7579_));
  AND2X1   g07515(.A(new_n7571_), .B(new_n7558_), .Y(new_n7580_));
  INVX1    g07516(.A(new_n7558_), .Y(new_n7581_));
  OR2X1    g07517(.A(new_n7564_), .B(new_n7562_), .Y(new_n7582_));
  OAI21X1  g07518(.A0(new_n7581_), .A1(new_n7537_), .B0(new_n7582_), .Y(new_n7583_));
  NOR2X1   g07519(.A(new_n7571_), .B(new_n7558_), .Y(new_n7584_));
  INVX1    g07520(.A(new_n7584_), .Y(new_n7585_));
  AOI21X1  g07521(.A0(new_n7585_), .A1(new_n7583_), .B0(new_n7580_), .Y(new_n7586_));
  INVX1    g07522(.A(new_n7586_), .Y(new_n7587_));
  XOR2X1   g07523(.A(new_n7578_), .B(new_n7571_), .Y(new_n7588_));
  AOI21X1  g07524(.A0(new_n7588_), .A1(new_n7587_), .B0(new_n7579_), .Y(new_n7589_));
  XOR2X1   g07525(.A(new_n7339_), .B(new_n7123_), .Y(new_n7590_));
  XOR2X1   g07526(.A(new_n7590_), .B(new_n7578_), .Y(new_n7591_));
  INVX1    g07527(.A(new_n7591_), .Y(new_n7592_));
  XOR2X1   g07528(.A(new_n7592_), .B(new_n7589_), .Y(new_n7593_));
  INVX1    g07529(.A(new_n7590_), .Y(new_n7594_));
  AOI22X1  g07530(.A0(new_n7578_), .A1(new_n2418_), .B0(new_n7571_), .B1(new_n2424_), .Y(new_n7595_));
  OAI21X1  g07531(.A0(new_n7594_), .A1(new_n2626_), .B0(new_n7595_), .Y(new_n7596_));
  AOI21X1  g07532(.A0(new_n7593_), .A1(new_n2301_), .B0(new_n7596_), .Y(new_n7597_));
  XOR2X1   g07533(.A(new_n7597_), .B(\a[26] ), .Y(new_n7598_));
  XOR2X1   g07534(.A(new_n7598_), .B(new_n7570_), .Y(new_n7599_));
  XOR2X1   g07535(.A(new_n7541_), .B(new_n7502_), .Y(new_n7600_));
  XOR2X1   g07536(.A(new_n7588_), .B(new_n7587_), .Y(new_n7601_));
  INVX1    g07537(.A(new_n7578_), .Y(new_n7602_));
  AOI22X1  g07538(.A0(new_n7571_), .A1(new_n2418_), .B0(new_n7558_), .B1(new_n2424_), .Y(new_n7603_));
  OAI21X1  g07539(.A0(new_n7602_), .A1(new_n2626_), .B0(new_n7603_), .Y(new_n7604_));
  AOI21X1  g07540(.A0(new_n7601_), .A1(new_n2301_), .B0(new_n7604_), .Y(new_n7605_));
  XOR2X1   g07541(.A(new_n7605_), .B(\a[26] ), .Y(new_n7606_));
  OR2X1    g07542(.A(new_n7606_), .B(new_n7600_), .Y(new_n7607_));
  XOR2X1   g07543(.A(new_n7606_), .B(new_n7600_), .Y(new_n7608_));
  XOR2X1   g07544(.A(new_n7498_), .B(new_n7411_), .Y(new_n7609_));
  NOR2X1   g07545(.A(new_n7492_), .B(new_n7490_), .Y(new_n7610_));
  XOR2X1   g07546(.A(new_n7524_), .B(new_n7610_), .Y(new_n7611_));
  INVX1    g07547(.A(new_n7611_), .Y(new_n7612_));
  AOI22X1  g07548(.A0(new_n7485_), .A1(new_n2095_), .B0(new_n7364_), .B1(new_n2185_), .Y(new_n7613_));
  OAI21X1  g07549(.A0(new_n7523_), .A1(new_n2140_), .B0(new_n7613_), .Y(new_n7614_));
  AOI21X1  g07550(.A0(new_n7612_), .A1(new_n2062_), .B0(new_n7614_), .Y(new_n7615_));
  XOR2X1   g07551(.A(new_n7615_), .B(\a[29] ), .Y(new_n7616_));
  INVX1    g07552(.A(new_n7616_), .Y(new_n7617_));
  AND2X1   g07553(.A(new_n7617_), .B(new_n7609_), .Y(new_n7618_));
  XOR2X1   g07554(.A(new_n7616_), .B(new_n7609_), .Y(new_n7619_));
  XOR2X1   g07555(.A(new_n7571_), .B(new_n7581_), .Y(new_n7620_));
  AOI22X1  g07556(.A0(new_n7586_), .A1(new_n7585_), .B0(new_n7620_), .B1(new_n7583_), .Y(new_n7621_));
  INVX1    g07557(.A(new_n7621_), .Y(new_n7622_));
  INVX1    g07558(.A(new_n7571_), .Y(new_n7623_));
  AOI22X1  g07559(.A0(new_n7558_), .A1(new_n2418_), .B0(new_n7529_), .B1(new_n2424_), .Y(new_n7624_));
  OAI21X1  g07560(.A0(new_n7623_), .A1(new_n2626_), .B0(new_n7624_), .Y(new_n7625_));
  AOI21X1  g07561(.A0(new_n7622_), .A1(new_n2301_), .B0(new_n7625_), .Y(new_n7626_));
  XOR2X1   g07562(.A(new_n7626_), .B(\a[26] ), .Y(new_n7627_));
  NOR2X1   g07563(.A(new_n7627_), .B(new_n7619_), .Y(new_n7628_));
  OAI21X1  g07564(.A0(new_n7628_), .A1(new_n7618_), .B0(new_n7608_), .Y(new_n7629_));
  AND2X1   g07565(.A(new_n7629_), .B(new_n7607_), .Y(new_n7630_));
  XOR2X1   g07566(.A(new_n7630_), .B(new_n7599_), .Y(new_n7631_));
  INVX1    g07567(.A(new_n7123_), .Y(new_n7632_));
  INVX1    g07568(.A(new_n7162_), .Y(new_n7633_));
  OAI21X1  g07569(.A0(new_n7577_), .A1(new_n7572_), .B0(new_n7633_), .Y(new_n7634_));
  AOI21X1  g07570(.A0(new_n7634_), .A1(new_n7632_), .B0(new_n7120_), .Y(new_n7635_));
  NAND3X1  g07571(.A(new_n7635_), .B(new_n7106_), .C(new_n7095_), .Y(new_n7636_));
  XOR2X1   g07572(.A(new_n7107_), .B(new_n7095_), .Y(new_n7637_));
  NOR2X1   g07573(.A(new_n7637_), .B(new_n7635_), .Y(new_n7638_));
  NOR2X1   g07574(.A(new_n7107_), .B(new_n7095_), .Y(new_n7639_));
  AND2X1   g07575(.A(new_n7107_), .B(new_n7095_), .Y(new_n7640_));
  NOR3X1   g07576(.A(new_n7640_), .B(new_n7639_), .C(new_n7340_), .Y(new_n7641_));
  NOR2X1   g07577(.A(new_n7641_), .B(new_n7638_), .Y(new_n7642_));
  AND2X1   g07578(.A(new_n7636_), .B(new_n7341_), .Y(new_n7643_));
  INVX1    g07579(.A(new_n7643_), .Y(new_n7644_));
  NOR2X1   g07580(.A(new_n7642_), .B(new_n7594_), .Y(new_n7645_));
  NOR3X1   g07581(.A(new_n7641_), .B(new_n7638_), .C(new_n7590_), .Y(new_n7646_));
  INVX1    g07582(.A(new_n7646_), .Y(new_n7647_));
  NAND2X1  g07583(.A(new_n7590_), .B(new_n7578_), .Y(new_n7648_));
  OAI21X1  g07584(.A0(new_n7592_), .A1(new_n7589_), .B0(new_n7648_), .Y(new_n7649_));
  AOI21X1  g07585(.A0(new_n7649_), .A1(new_n7647_), .B0(new_n7645_), .Y(new_n7650_));
  XOR2X1   g07586(.A(new_n7644_), .B(new_n7642_), .Y(new_n7651_));
  INVX1    g07587(.A(new_n7651_), .Y(new_n7652_));
  OR2X1    g07588(.A(new_n7652_), .B(new_n7650_), .Y(new_n7653_));
  OAI21X1  g07589(.A0(new_n7644_), .A1(new_n7642_), .B0(new_n7653_), .Y(new_n7654_));
  XOR2X1   g07590(.A(new_n7654_), .B(new_n7636_), .Y(new_n7655_));
  INVX1    g07591(.A(new_n7655_), .Y(new_n7656_));
  INVX1    g07592(.A(new_n7642_), .Y(new_n7657_));
  AOI22X1  g07593(.A0(new_n7657_), .A1(new_n2657_), .B0(new_n7341_), .B1(new_n2745_), .Y(new_n7658_));
  OAI21X1  g07594(.A0(new_n7644_), .A1(new_n2743_), .B0(new_n7658_), .Y(new_n7659_));
  AOI21X1  g07595(.A0(new_n7656_), .A1(new_n2658_), .B0(new_n7659_), .Y(new_n7660_));
  XOR2X1   g07596(.A(new_n7660_), .B(\a[23] ), .Y(new_n7661_));
  XOR2X1   g07597(.A(new_n7661_), .B(new_n7631_), .Y(new_n7662_));
  XOR2X1   g07598(.A(new_n7627_), .B(new_n7619_), .Y(new_n7663_));
  INVX1    g07599(.A(new_n7663_), .Y(new_n7664_));
  NOR2X1   g07600(.A(new_n7446_), .B(new_n7383_), .Y(new_n7665_));
  OAI22X1  g07601(.A0(new_n7665_), .A1(new_n7447_), .B0(new_n7476_), .B1(new_n7469_), .Y(new_n7666_));
  NOR4X1   g07602(.A(new_n7665_), .B(new_n7476_), .C(new_n7469_), .D(new_n7447_), .Y(new_n7667_));
  INVX1    g07603(.A(new_n7667_), .Y(new_n7668_));
  XOR2X1   g07604(.A(new_n6822_), .B(new_n6820_), .Y(new_n7669_));
  OAI22X1  g07605(.A0(new_n6992_), .A1(new_n6991_), .B0(new_n7669_), .B1(new_n6990_), .Y(new_n7670_));
  INVX1    g07606(.A(new_n6820_), .Y(new_n7671_));
  AOI22X1  g07607(.A0(new_n6882_), .A1(new_n1890_), .B0(new_n6822_), .B1(new_n1884_), .Y(new_n7672_));
  OAI21X1  g07608(.A0(new_n7671_), .A1(new_n3498_), .B0(new_n7672_), .Y(new_n7673_));
  AOI21X1  g07609(.A0(new_n7670_), .A1(new_n407_), .B0(new_n7673_), .Y(new_n7674_));
  AOI21X1  g07610(.A0(new_n7668_), .A1(new_n7666_), .B0(new_n7674_), .Y(new_n7675_));
  INVX1    g07611(.A(new_n7675_), .Y(new_n7676_));
  AND2X1   g07612(.A(new_n7668_), .B(new_n7666_), .Y(new_n7677_));
  INVX1    g07613(.A(new_n7677_), .Y(new_n7678_));
  XOR2X1   g07614(.A(new_n7674_), .B(new_n7678_), .Y(new_n7679_));
  INVX1    g07615(.A(new_n7046_), .Y(new_n7680_));
  OAI22X1  g07616(.A0(new_n7361_), .A1(new_n2431_), .B0(new_n7418_), .B1(new_n2186_), .Y(new_n7681_));
  AOI21X1  g07617(.A0(new_n7044_), .A1(new_n2139_), .B0(new_n7681_), .Y(new_n7682_));
  OAI21X1  g07618(.A0(new_n7680_), .A1(new_n2063_), .B0(new_n7682_), .Y(new_n7683_));
  XOR2X1   g07619(.A(new_n7683_), .B(new_n74_), .Y(new_n7684_));
  OAI21X1  g07620(.A0(new_n7684_), .A1(new_n7679_), .B0(new_n7676_), .Y(new_n7685_));
  AND2X1   g07621(.A(new_n7478_), .B(new_n7448_), .Y(new_n7686_));
  XOR2X1   g07622(.A(new_n7479_), .B(new_n7686_), .Y(new_n7687_));
  AND2X1   g07623(.A(new_n7687_), .B(new_n7685_), .Y(new_n7688_));
  INVX1    g07624(.A(new_n7685_), .Y(new_n7689_));
  XOR2X1   g07625(.A(new_n7687_), .B(new_n7689_), .Y(new_n7690_));
  AOI22X1  g07626(.A0(new_n7044_), .A1(new_n2095_), .B0(new_n6818_), .B1(new_n2185_), .Y(new_n7691_));
  OAI21X1  g07627(.A0(new_n7367_), .A1(new_n2140_), .B0(new_n7691_), .Y(new_n7692_));
  AOI21X1  g07628(.A0(new_n7366_), .A1(new_n2062_), .B0(new_n7692_), .Y(new_n7693_));
  XOR2X1   g07629(.A(new_n7693_), .B(\a[29] ), .Y(new_n7694_));
  NOR2X1   g07630(.A(new_n7694_), .B(new_n7690_), .Y(new_n7695_));
  XOR2X1   g07631(.A(new_n7497_), .B(new_n7484_), .Y(new_n7696_));
  OAI21X1  g07632(.A0(new_n7695_), .A1(new_n7688_), .B0(new_n7696_), .Y(new_n7697_));
  NOR2X1   g07633(.A(new_n7695_), .B(new_n7688_), .Y(new_n7698_));
  XOR2X1   g07634(.A(new_n7696_), .B(new_n7698_), .Y(new_n7699_));
  AOI22X1  g07635(.A0(new_n7529_), .A1(new_n2418_), .B0(new_n7522_), .B1(new_n2424_), .Y(new_n7700_));
  OAI21X1  g07636(.A0(new_n7581_), .A1(new_n2626_), .B0(new_n7700_), .Y(new_n7701_));
  AOI21X1  g07637(.A0(new_n7565_), .A1(new_n2301_), .B0(new_n7701_), .Y(new_n7702_));
  XOR2X1   g07638(.A(new_n7702_), .B(\a[26] ), .Y(new_n7703_));
  OR2X1    g07639(.A(new_n7703_), .B(new_n7699_), .Y(new_n7704_));
  AOI21X1  g07640(.A0(new_n7704_), .A1(new_n7697_), .B0(new_n7664_), .Y(new_n7705_));
  INVX1    g07641(.A(new_n7705_), .Y(new_n7706_));
  AND2X1   g07642(.A(new_n7704_), .B(new_n7697_), .Y(new_n7707_));
  AND2X1   g07643(.A(new_n7707_), .B(new_n7664_), .Y(new_n7708_));
  OAI21X1  g07644(.A0(new_n7646_), .A1(new_n7645_), .B0(new_n7649_), .Y(new_n7709_));
  NAND2X1  g07645(.A(new_n7650_), .B(new_n7647_), .Y(new_n7710_));
  AND2X1   g07646(.A(new_n7710_), .B(new_n7709_), .Y(new_n7711_));
  INVX1    g07647(.A(new_n7711_), .Y(new_n7712_));
  AOI22X1  g07648(.A0(new_n7590_), .A1(new_n2696_), .B0(new_n7578_), .B1(new_n2657_), .Y(new_n7713_));
  OAI21X1  g07649(.A0(new_n7642_), .A1(new_n2753_), .B0(new_n7713_), .Y(new_n7714_));
  AOI21X1  g07650(.A0(new_n7712_), .A1(new_n2658_), .B0(new_n7714_), .Y(new_n7715_));
  XOR2X1   g07651(.A(new_n7715_), .B(\a[23] ), .Y(new_n7716_));
  OAI21X1  g07652(.A0(new_n7716_), .A1(new_n7708_), .B0(new_n7706_), .Y(new_n7717_));
  XOR2X1   g07653(.A(new_n7652_), .B(new_n7650_), .Y(new_n7718_));
  AOI22X1  g07654(.A0(new_n7643_), .A1(new_n2745_), .B0(new_n7590_), .B1(new_n2657_), .Y(new_n7719_));
  OAI21X1  g07655(.A0(new_n7642_), .A1(new_n2743_), .B0(new_n7719_), .Y(new_n7720_));
  AOI21X1  g07656(.A0(new_n7718_), .A1(new_n2658_), .B0(new_n7720_), .Y(new_n7721_));
  XOR2X1   g07657(.A(new_n7721_), .B(\a[23] ), .Y(new_n7722_));
  INVX1    g07658(.A(new_n7722_), .Y(new_n7723_));
  AOI21X1  g07659(.A0(new_n7617_), .A1(new_n7609_), .B0(new_n7628_), .Y(new_n7724_));
  XOR2X1   g07660(.A(new_n7724_), .B(new_n7608_), .Y(new_n7725_));
  XOR2X1   g07661(.A(new_n7722_), .B(new_n7717_), .Y(new_n7726_));
  NOR2X1   g07662(.A(new_n7726_), .B(new_n7725_), .Y(new_n7727_));
  AOI21X1  g07663(.A0(new_n7723_), .A1(new_n7717_), .B0(new_n7727_), .Y(new_n7728_));
  XOR2X1   g07664(.A(new_n7728_), .B(new_n7662_), .Y(new_n7729_));
  INVX1    g07665(.A(new_n7729_), .Y(new_n7730_));
  XOR2X1   g07666(.A(new_n7703_), .B(new_n7699_), .Y(new_n7731_));
  INVX1    g07667(.A(new_n7731_), .Y(new_n7732_));
  XOR2X1   g07668(.A(new_n7694_), .B(new_n7690_), .Y(new_n7733_));
  AOI22X1  g07669(.A0(new_n7522_), .A1(new_n2418_), .B0(new_n7485_), .B1(new_n2424_), .Y(new_n7734_));
  OAI21X1  g07670(.A0(new_n7537_), .A1(new_n2626_), .B0(new_n7734_), .Y(new_n7735_));
  AOI21X1  g07671(.A0(new_n7536_), .A1(new_n2301_), .B0(new_n7735_), .Y(new_n7736_));
  XOR2X1   g07672(.A(new_n7736_), .B(\a[26] ), .Y(new_n7737_));
  INVX1    g07673(.A(new_n7737_), .Y(new_n7738_));
  XOR2X1   g07674(.A(new_n7737_), .B(new_n7733_), .Y(new_n7739_));
  INVX1    g07675(.A(new_n7455_), .Y(new_n7740_));
  OR4X1    g07676(.A(new_n2173_), .B(new_n460_), .C(new_n418_), .D(new_n304_), .Y(new_n7741_));
  AOI21X1  g07677(.A0(new_n131_), .A1(new_n92_), .B0(new_n102_), .Y(new_n7742_));
  AOI21X1  g07678(.A0(new_n161_), .A1(new_n72_), .B0(new_n88_), .Y(new_n7743_));
  OR4X1    g07679(.A(new_n7743_), .B(new_n7742_), .C(new_n348_), .D(new_n201_), .Y(new_n7744_));
  OR4X1    g07680(.A(new_n831_), .B(new_n766_), .C(new_n396_), .D(new_n80_), .Y(new_n7745_));
  OR4X1    g07681(.A(new_n1028_), .B(new_n393_), .C(new_n410_), .D(new_n610_), .Y(new_n7746_));
  OR2X1    g07682(.A(new_n652_), .B(new_n441_), .Y(new_n7747_));
  OR4X1    g07683(.A(new_n7747_), .B(new_n7746_), .C(new_n7745_), .D(new_n7744_), .Y(new_n7748_));
  OR4X1    g07684(.A(new_n7748_), .B(new_n7741_), .C(new_n908_), .D(new_n842_), .Y(new_n7749_));
  OR4X1    g07685(.A(new_n2451_), .B(new_n2572_), .C(new_n1136_), .D(new_n896_), .Y(new_n7750_));
  OR4X1    g07686(.A(new_n1609_), .B(new_n874_), .C(new_n1633_), .D(new_n170_), .Y(new_n7751_));
  OR4X1    g07687(.A(new_n455_), .B(new_n259_), .C(new_n231_), .D(new_n338_), .Y(new_n7752_));
  OR4X1    g07688(.A(new_n7752_), .B(new_n7751_), .C(new_n1963_), .D(new_n1962_), .Y(new_n7753_));
  OR4X1    g07689(.A(new_n296_), .B(new_n191_), .C(new_n327_), .D(new_n1579_), .Y(new_n7754_));
  OR2X1    g07690(.A(new_n823_), .B(new_n552_), .Y(new_n7755_));
  OR4X1    g07691(.A(new_n938_), .B(new_n631_), .C(new_n702_), .D(new_n523_), .Y(new_n7756_));
  OR4X1    g07692(.A(new_n7756_), .B(new_n7755_), .C(new_n7754_), .D(new_n591_), .Y(new_n7757_));
  OR4X1    g07693(.A(new_n7757_), .B(new_n7753_), .C(new_n7750_), .D(new_n2229_), .Y(new_n7758_));
  NOR3X1   g07694(.A(new_n7758_), .B(new_n7749_), .C(new_n1454_), .Y(new_n7759_));
  NOR2X1   g07695(.A(new_n7759_), .B(new_n7740_), .Y(new_n7760_));
  XOR2X1   g07696(.A(new_n6887_), .B(new_n6885_), .Y(new_n7761_));
  OAI22X1  g07697(.A0(new_n6985_), .A1(new_n6984_), .B0(new_n7761_), .B1(new_n6983_), .Y(new_n7762_));
  AOI22X1  g07698(.A0(new_n6890_), .A1(new_n1890_), .B0(new_n6887_), .B1(new_n1884_), .Y(new_n7763_));
  OAI21X1  g07699(.A0(new_n6886_), .A1(new_n3498_), .B0(new_n7763_), .Y(new_n7764_));
  AOI21X1  g07700(.A0(new_n7762_), .A1(new_n407_), .B0(new_n7764_), .Y(new_n7765_));
  XOR2X1   g07701(.A(new_n7759_), .B(new_n7455_), .Y(new_n7766_));
  NOR2X1   g07702(.A(new_n7766_), .B(new_n7765_), .Y(new_n7767_));
  OR2X1    g07703(.A(new_n7767_), .B(new_n7760_), .Y(new_n7768_));
  XOR2X1   g07704(.A(new_n7467_), .B(new_n7466_), .Y(new_n7769_));
  AND2X1   g07705(.A(new_n7769_), .B(new_n7768_), .Y(new_n7770_));
  XOR2X1   g07706(.A(new_n6986_), .B(new_n6985_), .Y(new_n7771_));
  AOI22X1  g07707(.A0(new_n6887_), .A1(new_n1890_), .B0(new_n6885_), .B1(new_n1884_), .Y(new_n7772_));
  OAI21X1  g07708(.A0(new_n6884_), .A1(new_n3498_), .B0(new_n7772_), .Y(new_n7773_));
  AOI21X1  g07709(.A0(new_n7771_), .A1(new_n407_), .B0(new_n7773_), .Y(new_n7774_));
  INVX1    g07710(.A(new_n7774_), .Y(new_n7775_));
  XOR2X1   g07711(.A(new_n7769_), .B(new_n7768_), .Y(new_n7776_));
  AOI21X1  g07712(.A0(new_n7776_), .A1(new_n7775_), .B0(new_n7770_), .Y(new_n7777_));
  INVX1    g07713(.A(new_n7777_), .Y(new_n7778_));
  XOR2X1   g07714(.A(new_n7475_), .B(new_n7470_), .Y(new_n7779_));
  XOR2X1   g07715(.A(new_n7779_), .B(new_n7777_), .Y(new_n7780_));
  OAI22X1  g07716(.A0(new_n7671_), .A1(new_n2186_), .B0(new_n7418_), .B1(new_n2431_), .Y(new_n7781_));
  AOI21X1  g07717(.A0(new_n6818_), .A1(new_n2139_), .B0(new_n7781_), .Y(new_n7782_));
  OAI21X1  g07718(.A0(new_n7403_), .A1(new_n2063_), .B0(new_n7782_), .Y(new_n7783_));
  XOR2X1   g07719(.A(new_n7783_), .B(new_n74_), .Y(new_n7784_));
  NOR2X1   g07720(.A(new_n7784_), .B(new_n7780_), .Y(new_n7785_));
  AOI21X1  g07721(.A0(new_n7779_), .A1(new_n7778_), .B0(new_n7785_), .Y(new_n7786_));
  INVX1    g07722(.A(new_n7786_), .Y(new_n7787_));
  XOR2X1   g07723(.A(new_n7684_), .B(new_n7679_), .Y(new_n7788_));
  AND2X1   g07724(.A(new_n7788_), .B(new_n7787_), .Y(new_n7789_));
  XOR2X1   g07725(.A(new_n7788_), .B(new_n7787_), .Y(new_n7790_));
  AOI22X1  g07726(.A0(new_n7485_), .A1(new_n2418_), .B0(new_n7364_), .B1(new_n2424_), .Y(new_n7791_));
  OAI21X1  g07727(.A0(new_n7523_), .A1(new_n2626_), .B0(new_n7791_), .Y(new_n7792_));
  AOI21X1  g07728(.A0(new_n7612_), .A1(new_n2301_), .B0(new_n7792_), .Y(new_n7793_));
  XOR2X1   g07729(.A(new_n7793_), .B(new_n89_), .Y(new_n7794_));
  AOI21X1  g07730(.A0(new_n7794_), .A1(new_n7790_), .B0(new_n7789_), .Y(new_n7795_));
  NOR2X1   g07731(.A(new_n7795_), .B(new_n7739_), .Y(new_n7796_));
  AOI21X1  g07732(.A0(new_n7738_), .A1(new_n7733_), .B0(new_n7796_), .Y(new_n7797_));
  NOR2X1   g07733(.A(new_n7797_), .B(new_n7732_), .Y(new_n7798_));
  XOR2X1   g07734(.A(new_n7797_), .B(new_n7732_), .Y(new_n7799_));
  AOI22X1  g07735(.A0(new_n7578_), .A1(new_n2696_), .B0(new_n7571_), .B1(new_n2657_), .Y(new_n7800_));
  OAI21X1  g07736(.A0(new_n7594_), .A1(new_n2753_), .B0(new_n7800_), .Y(new_n7801_));
  AOI21X1  g07737(.A0(new_n7593_), .A1(new_n2658_), .B0(new_n7801_), .Y(new_n7802_));
  XOR2X1   g07738(.A(new_n7802_), .B(new_n70_), .Y(new_n7803_));
  AOI21X1  g07739(.A0(new_n7803_), .A1(new_n7799_), .B0(new_n7798_), .Y(new_n7804_));
  MX2X1    g07740(.A(new_n2874_), .B(new_n2873_), .S0(new_n2869_), .Y(new_n7805_));
  AOI22X1  g07741(.A0(new_n7643_), .A1(new_n2875_), .B0(new_n7805_), .B1(new_n7341_), .Y(new_n7806_));
  MX2X1    g07742(.A(new_n7654_), .B(new_n7341_), .S0(new_n7636_), .Y(new_n7807_));
  INVX1    g07743(.A(new_n7807_), .Y(new_n7808_));
  OAI21X1  g07744(.A0(new_n7808_), .A1(new_n3098_), .B0(new_n7806_), .Y(new_n7809_));
  XOR2X1   g07745(.A(new_n7809_), .B(new_n1920_), .Y(new_n7810_));
  NOR2X1   g07746(.A(new_n7810_), .B(new_n7804_), .Y(new_n7811_));
  XOR2X1   g07747(.A(new_n7707_), .B(new_n7664_), .Y(new_n7812_));
  XOR2X1   g07748(.A(new_n7716_), .B(new_n7812_), .Y(new_n7813_));
  INVX1    g07749(.A(new_n7813_), .Y(new_n7814_));
  XOR2X1   g07750(.A(new_n7810_), .B(new_n7804_), .Y(new_n7815_));
  AOI21X1  g07751(.A0(new_n7815_), .A1(new_n7814_), .B0(new_n7811_), .Y(new_n7816_));
  INVX1    g07752(.A(new_n7816_), .Y(new_n7817_));
  XOR2X1   g07753(.A(new_n7726_), .B(new_n7725_), .Y(new_n7818_));
  AND2X1   g07754(.A(new_n7818_), .B(new_n7817_), .Y(new_n7819_));
  XOR2X1   g07755(.A(new_n7815_), .B(new_n7813_), .Y(new_n7820_));
  XOR2X1   g07756(.A(new_n7803_), .B(new_n7799_), .Y(new_n7821_));
  INVX1    g07757(.A(new_n7821_), .Y(new_n7822_));
  XOR2X1   g07758(.A(new_n7795_), .B(new_n7739_), .Y(new_n7823_));
  AOI22X1  g07759(.A0(new_n7571_), .A1(new_n2696_), .B0(new_n7558_), .B1(new_n2657_), .Y(new_n7824_));
  OAI21X1  g07760(.A0(new_n7602_), .A1(new_n2753_), .B0(new_n7824_), .Y(new_n7825_));
  AOI21X1  g07761(.A0(new_n7601_), .A1(new_n2658_), .B0(new_n7825_), .Y(new_n7826_));
  XOR2X1   g07762(.A(new_n7826_), .B(\a[23] ), .Y(new_n7827_));
  INVX1    g07763(.A(new_n7827_), .Y(new_n7828_));
  XOR2X1   g07764(.A(new_n7827_), .B(new_n7823_), .Y(new_n7829_));
  XOR2X1   g07765(.A(new_n7793_), .B(\a[26] ), .Y(new_n7830_));
  XOR2X1   g07766(.A(new_n7830_), .B(new_n7790_), .Y(new_n7831_));
  XOR2X1   g07767(.A(new_n7776_), .B(new_n7774_), .Y(new_n7832_));
  AOI22X1  g07768(.A0(new_n6822_), .A1(new_n2185_), .B0(new_n6820_), .B1(new_n2095_), .Y(new_n7833_));
  OAI21X1  g07769(.A0(new_n7418_), .A1(new_n2140_), .B0(new_n7833_), .Y(new_n7834_));
  AOI21X1  g07770(.A0(new_n7417_), .A1(new_n2062_), .B0(new_n7834_), .Y(new_n7835_));
  XOR2X1   g07771(.A(new_n7835_), .B(\a[29] ), .Y(new_n7836_));
  NOR2X1   g07772(.A(new_n7836_), .B(new_n7832_), .Y(new_n7837_));
  INVX1    g07773(.A(new_n7837_), .Y(new_n7838_));
  XOR2X1   g07774(.A(new_n7836_), .B(new_n7832_), .Y(new_n7839_));
  INVX1    g07775(.A(new_n7839_), .Y(new_n7840_));
  NOR4X1   g07776(.A(new_n7758_), .B(new_n7749_), .C(new_n7455_), .D(new_n1454_), .Y(new_n7841_));
  OAI22X1  g07777(.A0(new_n7768_), .A1(new_n7841_), .B0(new_n7767_), .B1(new_n7765_), .Y(new_n7842_));
  OR4X1    g07778(.A(new_n627_), .B(new_n218_), .C(new_n183_), .D(new_n155_), .Y(new_n7843_));
  OAI22X1  g07779(.A0(new_n152_), .A1(new_n92_), .B0(new_n105_), .B1(new_n75_), .Y(new_n7844_));
  OR4X1    g07780(.A(new_n7844_), .B(new_n2945_), .C(new_n646_), .D(new_n497_), .Y(new_n7845_));
  OR4X1    g07781(.A(new_n1416_), .B(new_n1114_), .C(new_n1090_), .D(new_n164_), .Y(new_n7846_));
  OR4X1    g07782(.A(new_n7846_), .B(new_n7845_), .C(new_n7843_), .D(new_n1336_), .Y(new_n7847_));
  NOR4X1   g07783(.A(new_n400_), .B(new_n177_), .C(new_n327_), .D(new_n581_), .Y(new_n7848_));
  NOR2X1   g07784(.A(new_n1717_), .B(new_n165_), .Y(new_n7849_));
  NOR4X1   g07785(.A(new_n372_), .B(new_n361_), .C(new_n603_), .D(new_n239_), .Y(new_n7850_));
  NAND4X1  g07786(.A(new_n7850_), .B(new_n7849_), .C(new_n7848_), .D(new_n1001_), .Y(new_n7851_));
  OR4X1    g07787(.A(new_n642_), .B(new_n383_), .C(new_n598_), .D(new_n304_), .Y(new_n7852_));
  OR4X1    g07788(.A(new_n7852_), .B(new_n292_), .C(new_n493_), .D(new_n215_), .Y(new_n7853_));
  OR4X1    g07789(.A(new_n7853_), .B(new_n7851_), .C(new_n7134_), .D(new_n1394_), .Y(new_n7854_));
  NOR4X1   g07790(.A(new_n7854_), .B(new_n7847_), .C(new_n3463_), .D(new_n1767_), .Y(new_n7855_));
  OR4X1    g07791(.A(new_n1531_), .B(new_n869_), .C(new_n176_), .D(new_n137_), .Y(new_n7856_));
  OR2X1    g07792(.A(new_n7856_), .B(new_n946_), .Y(new_n7857_));
  NAND3X1  g07793(.A(new_n2168_), .B(new_n1545_), .C(new_n796_), .Y(new_n7858_));
  OR4X1    g07794(.A(new_n1657_), .B(new_n835_), .C(new_n586_), .D(new_n494_), .Y(new_n7859_));
  OR4X1    g07795(.A(new_n1261_), .B(new_n843_), .C(new_n293_), .D(new_n147_), .Y(new_n7860_));
  OR4X1    g07796(.A(new_n7860_), .B(new_n7859_), .C(new_n7858_), .D(new_n216_), .Y(new_n7861_));
  OR4X1    g07797(.A(new_n7861_), .B(new_n7857_), .C(new_n2120_), .D(new_n2113_), .Y(new_n7862_));
  NOR4X1   g07798(.A(new_n7862_), .B(new_n3285_), .C(new_n911_), .D(new_n492_), .Y(new_n7863_));
  NOR2X1   g07799(.A(new_n7863_), .B(new_n7855_), .Y(new_n7864_));
  OR4X1    g07800(.A(new_n4428_), .B(new_n4247_), .C(new_n4080_), .D(new_n4078_), .Y(new_n7865_));
  AND2X1   g07801(.A(new_n7865_), .B(new_n7341_), .Y(new_n7866_));
  XOR2X1   g07802(.A(new_n7866_), .B(new_n2911_), .Y(new_n7867_));
  XOR2X1   g07803(.A(new_n7863_), .B(new_n7855_), .Y(new_n7868_));
  AOI21X1  g07804(.A0(new_n7868_), .A1(new_n7867_), .B0(new_n7864_), .Y(new_n7869_));
  OR2X1    g07805(.A(new_n7869_), .B(new_n7740_), .Y(new_n7870_));
  XOR2X1   g07806(.A(new_n7869_), .B(new_n7455_), .Y(new_n7871_));
  INVX1    g07807(.A(new_n6982_), .Y(new_n7872_));
  AND2X1   g07808(.A(new_n7872_), .B(new_n6981_), .Y(new_n7873_));
  NOR2X1   g07809(.A(new_n6890_), .B(new_n6887_), .Y(new_n7874_));
  NOR3X1   g07810(.A(new_n7874_), .B(new_n6981_), .C(new_n6891_), .Y(new_n7875_));
  NOR2X1   g07811(.A(new_n7875_), .B(new_n7873_), .Y(new_n7876_));
  INVX1    g07812(.A(new_n7876_), .Y(new_n7877_));
  INVX1    g07813(.A(new_n6887_), .Y(new_n7878_));
  AOI22X1  g07814(.A0(new_n6892_), .A1(new_n1890_), .B0(new_n6890_), .B1(new_n1884_), .Y(new_n7879_));
  OAI21X1  g07815(.A0(new_n7878_), .A1(new_n3498_), .B0(new_n7879_), .Y(new_n7880_));
  AOI21X1  g07816(.A0(new_n7877_), .A1(new_n407_), .B0(new_n7880_), .Y(new_n7881_));
  OAI21X1  g07817(.A0(new_n7881_), .A1(new_n7871_), .B0(new_n7870_), .Y(new_n7882_));
  XOR2X1   g07818(.A(new_n7882_), .B(new_n7842_), .Y(new_n7883_));
  XOR2X1   g07819(.A(new_n6980_), .B(new_n6978_), .Y(new_n7884_));
  INVX1    g07820(.A(new_n6890_), .Y(new_n7885_));
  AOI22X1  g07821(.A0(new_n6894_), .A1(new_n1890_), .B0(new_n6892_), .B1(new_n1884_), .Y(new_n7886_));
  OAI21X1  g07822(.A0(new_n7885_), .A1(new_n3498_), .B0(new_n7886_), .Y(new_n7887_));
  AOI21X1  g07823(.A0(new_n7884_), .A1(new_n407_), .B0(new_n7887_), .Y(new_n7888_));
  INVX1    g07824(.A(new_n7888_), .Y(new_n7889_));
  XOR2X1   g07825(.A(new_n7868_), .B(new_n7867_), .Y(new_n7890_));
  AND2X1   g07826(.A(new_n7890_), .B(new_n7889_), .Y(new_n7891_));
  XOR2X1   g07827(.A(new_n7890_), .B(new_n7888_), .Y(new_n7892_));
  INVX1    g07828(.A(new_n7855_), .Y(new_n7893_));
  OR4X1    g07829(.A(new_n509_), .B(new_n263_), .C(new_n1008_), .D(new_n80_), .Y(new_n7894_));
  NOR3X1   g07830(.A(new_n7894_), .B(new_n1061_), .C(new_n1000_), .Y(new_n7895_));
  OR4X1    g07831(.A(new_n812_), .B(new_n226_), .C(new_n197_), .D(new_n175_), .Y(new_n7896_));
  NOR4X1   g07832(.A(new_n7896_), .B(new_n497_), .C(new_n869_), .D(new_n265_), .Y(new_n7897_));
  OR4X1    g07833(.A(new_n2088_), .B(new_n1100_), .C(new_n7149_), .D(new_n1018_), .Y(new_n7898_));
  OR4X1    g07834(.A(new_n571_), .B(new_n323_), .C(new_n162_), .D(new_n124_), .Y(new_n7899_));
  NOR4X1   g07835(.A(new_n7899_), .B(new_n7898_), .C(new_n1702_), .D(new_n430_), .Y(new_n7900_));
  NAND4X1  g07836(.A(new_n7900_), .B(new_n7897_), .C(new_n7895_), .D(new_n1365_), .Y(new_n7901_));
  NOR3X1   g07837(.A(new_n1474_), .B(new_n1623_), .C(new_n641_), .Y(new_n7902_));
  NOR3X1   g07838(.A(new_n372_), .B(new_n280_), .C(new_n144_), .Y(new_n7903_));
  NOR4X1   g07839(.A(new_n246_), .B(new_n231_), .C(new_n229_), .D(new_n974_), .Y(new_n7904_));
  NAND3X1  g07840(.A(new_n7904_), .B(new_n7903_), .C(new_n7902_), .Y(new_n7905_));
  OR4X1    g07841(.A(new_n806_), .B(new_n615_), .C(new_n399_), .D(new_n357_), .Y(new_n7906_));
  OR4X1    g07842(.A(new_n543_), .B(new_n691_), .C(new_n276_), .D(new_n273_), .Y(new_n7907_));
  OR4X1    g07843(.A(new_n7907_), .B(new_n7906_), .C(new_n1234_), .D(new_n435_), .Y(new_n7908_));
  OR4X1    g07844(.A(new_n7908_), .B(new_n7747_), .C(new_n1756_), .D(new_n1989_), .Y(new_n7909_));
  NOR4X1   g07845(.A(new_n7909_), .B(new_n7905_), .C(new_n7901_), .D(new_n2525_), .Y(new_n7910_));
  OR2X1    g07846(.A(new_n7910_), .B(new_n7893_), .Y(new_n7911_));
  OR4X1    g07847(.A(new_n1417_), .B(new_n441_), .C(new_n294_), .D(new_n812_), .Y(new_n7912_));
  OAI22X1  g07848(.A0(new_n148_), .A1(new_n72_), .B0(new_n90_), .B1(new_n79_), .Y(new_n7913_));
  OR4X1    g07849(.A(new_n7913_), .B(new_n1166_), .C(new_n312_), .D(new_n76_), .Y(new_n7914_));
  OR2X1    g07850(.A(new_n2153_), .B(new_n723_), .Y(new_n7915_));
  OR4X1    g07851(.A(new_n1538_), .B(new_n1210_), .C(new_n850_), .D(new_n231_), .Y(new_n7916_));
  OR4X1    g07852(.A(new_n414_), .B(new_n365_), .C(new_n233_), .D(new_n449_), .Y(new_n7917_));
  OAI22X1  g07853(.A0(new_n131_), .A1(new_n115_), .B0(new_n108_), .B1(new_n91_), .Y(new_n7918_));
  OR4X1    g07854(.A(new_n7918_), .B(new_n7917_), .C(new_n7916_), .D(new_n239_), .Y(new_n7919_));
  OR4X1    g07855(.A(new_n7919_), .B(new_n7915_), .C(new_n1876_), .D(new_n189_), .Y(new_n7920_));
  OR4X1    g07856(.A(new_n7920_), .B(new_n7914_), .C(new_n7912_), .D(new_n1944_), .Y(new_n7921_));
  INVX1    g07857(.A(new_n458_), .Y(new_n7922_));
  OAI22X1  g07858(.A0(new_n161_), .A1(new_n106_), .B0(new_n127_), .B1(new_n75_), .Y(new_n7923_));
  NOR4X1   g07859(.A(new_n2101_), .B(new_n7923_), .C(new_n224_), .D(new_n160_), .Y(new_n7924_));
  NOR4X1   g07860(.A(new_n938_), .B(new_n355_), .C(new_n323_), .D(new_n455_), .Y(new_n7925_));
  NAND4X1  g07861(.A(new_n7925_), .B(new_n7924_), .C(new_n7385_), .D(new_n7922_), .Y(new_n7926_));
  OR4X1    g07862(.A(new_n1514_), .B(new_n755_), .C(new_n552_), .D(new_n299_), .Y(new_n7927_));
  OR4X1    g07863(.A(new_n480_), .B(new_n578_), .C(new_n116_), .D(new_n114_), .Y(new_n7928_));
  OR4X1    g07864(.A(new_n7928_), .B(new_n741_), .C(new_n691_), .D(new_n303_), .Y(new_n7929_));
  OR4X1    g07865(.A(new_n7929_), .B(new_n7927_), .C(new_n2459_), .D(new_n1036_), .Y(new_n7930_));
  NOR4X1   g07866(.A(new_n7930_), .B(new_n7926_), .C(new_n7921_), .D(new_n1569_), .Y(new_n7931_));
  NOR4X1   g07867(.A(new_n755_), .B(new_n546_), .C(new_n420_), .D(new_n493_), .Y(new_n7932_));
  NOR2X1   g07868(.A(new_n728_), .B(new_n165_), .Y(new_n7933_));
  NAND4X1  g07869(.A(new_n7933_), .B(new_n7932_), .C(new_n1405_), .D(new_n1250_), .Y(new_n7934_));
  OR4X1    g07870(.A(new_n1082_), .B(new_n527_), .C(new_n1261_), .D(new_n408_), .Y(new_n7935_));
  OR4X1    g07871(.A(new_n276_), .B(new_n265_), .C(new_n381_), .D(new_n449_), .Y(new_n7936_));
  OR4X1    g07872(.A(new_n7936_), .B(new_n7935_), .C(new_n2915_), .D(new_n685_), .Y(new_n7937_));
  OAI22X1  g07873(.A0(new_n131_), .A1(new_n115_), .B0(new_n123_), .B1(new_n72_), .Y(new_n7938_));
  OR2X1    g07874(.A(new_n7938_), .B(new_n455_), .Y(new_n7939_));
  OR4X1    g07875(.A(new_n589_), .B(new_n547_), .C(new_n523_), .D(new_n1008_), .Y(new_n7940_));
  OR2X1    g07876(.A(new_n7940_), .B(new_n7939_), .Y(new_n7941_));
  OR4X1    g07877(.A(new_n1558_), .B(new_n1341_), .C(new_n1255_), .D(new_n440_), .Y(new_n7942_));
  OR4X1    g07878(.A(new_n7942_), .B(new_n7941_), .C(new_n7937_), .D(new_n7934_), .Y(new_n7943_));
  NOR3X1   g07879(.A(new_n7943_), .B(new_n7193_), .C(new_n942_), .Y(new_n7944_));
  NOR2X1   g07880(.A(new_n7944_), .B(new_n7931_), .Y(new_n7945_));
  OR4X1    g07881(.A(new_n5097_), .B(new_n4870_), .C(new_n4637_), .D(new_n4635_), .Y(new_n7946_));
  AND2X1   g07882(.A(new_n7946_), .B(new_n7341_), .Y(new_n7947_));
  XOR2X1   g07883(.A(new_n7947_), .B(new_n2995_), .Y(new_n7948_));
  XOR2X1   g07884(.A(new_n7944_), .B(new_n7931_), .Y(new_n7949_));
  AOI21X1  g07885(.A0(new_n7949_), .A1(new_n7948_), .B0(new_n7945_), .Y(new_n7950_));
  NOR2X1   g07886(.A(new_n7950_), .B(new_n7893_), .Y(new_n7951_));
  XOR2X1   g07887(.A(new_n7950_), .B(new_n7855_), .Y(new_n7952_));
  XOR2X1   g07888(.A(new_n6974_), .B(new_n6973_), .Y(new_n7953_));
  AOI22X1  g07889(.A0(new_n6899_), .A1(new_n1890_), .B0(new_n6897_), .B1(new_n1884_), .Y(new_n7954_));
  OAI21X1  g07890(.A0(new_n6896_), .A1(new_n3498_), .B0(new_n7954_), .Y(new_n7955_));
  AOI21X1  g07891(.A0(new_n7953_), .A1(new_n407_), .B0(new_n7955_), .Y(new_n7956_));
  NOR2X1   g07892(.A(new_n7956_), .B(new_n7952_), .Y(new_n7957_));
  XOR2X1   g07893(.A(new_n7910_), .B(new_n7893_), .Y(new_n7958_));
  OAI21X1  g07894(.A0(new_n7957_), .A1(new_n7951_), .B0(new_n7958_), .Y(new_n7959_));
  AOI21X1  g07895(.A0(new_n7959_), .A1(new_n7911_), .B0(new_n7892_), .Y(new_n7960_));
  XOR2X1   g07896(.A(new_n7881_), .B(new_n7871_), .Y(new_n7961_));
  OAI21X1  g07897(.A0(new_n7960_), .A1(new_n7891_), .B0(new_n7961_), .Y(new_n7962_));
  NOR2X1   g07898(.A(new_n7960_), .B(new_n7891_), .Y(new_n7963_));
  XOR2X1   g07899(.A(new_n7961_), .B(new_n7963_), .Y(new_n7964_));
  INVX1    g07900(.A(new_n7471_), .Y(new_n7965_));
  OAI22X1  g07901(.A0(new_n6886_), .A1(new_n2186_), .B0(new_n6884_), .B1(new_n2431_), .Y(new_n7966_));
  AOI21X1  g07902(.A0(new_n6822_), .A1(new_n2139_), .B0(new_n7966_), .Y(new_n7967_));
  OAI21X1  g07903(.A0(new_n7965_), .A1(new_n2063_), .B0(new_n7967_), .Y(new_n7968_));
  XOR2X1   g07904(.A(new_n7968_), .B(new_n74_), .Y(new_n7969_));
  OAI21X1  g07905(.A0(new_n7969_), .A1(new_n7964_), .B0(new_n7962_), .Y(new_n7970_));
  AND2X1   g07906(.A(new_n7970_), .B(new_n7883_), .Y(new_n7971_));
  AOI21X1  g07907(.A0(new_n7882_), .A1(new_n7842_), .B0(new_n7971_), .Y(new_n7972_));
  OAI21X1  g07908(.A0(new_n7972_), .A1(new_n7840_), .B0(new_n7838_), .Y(new_n7973_));
  XOR2X1   g07909(.A(new_n7784_), .B(new_n7780_), .Y(new_n7974_));
  AND2X1   g07910(.A(new_n7974_), .B(new_n7973_), .Y(new_n7975_));
  XOR2X1   g07911(.A(new_n7974_), .B(new_n7973_), .Y(new_n7976_));
  AOI22X1  g07912(.A0(new_n7364_), .A1(new_n2418_), .B0(new_n7044_), .B1(new_n2424_), .Y(new_n7977_));
  OAI21X1  g07913(.A0(new_n7504_), .A1(new_n2626_), .B0(new_n7977_), .Y(new_n7978_));
  AOI21X1  g07914(.A0(new_n7552_), .A1(new_n2301_), .B0(new_n7978_), .Y(new_n7979_));
  XOR2X1   g07915(.A(new_n7979_), .B(new_n89_), .Y(new_n7980_));
  AOI21X1  g07916(.A0(new_n7980_), .A1(new_n7976_), .B0(new_n7975_), .Y(new_n7981_));
  NOR2X1   g07917(.A(new_n7981_), .B(new_n7831_), .Y(new_n7982_));
  XOR2X1   g07918(.A(new_n7981_), .B(new_n7831_), .Y(new_n7983_));
  AOI22X1  g07919(.A0(new_n7558_), .A1(new_n2696_), .B0(new_n7529_), .B1(new_n2657_), .Y(new_n7984_));
  OAI21X1  g07920(.A0(new_n7623_), .A1(new_n2753_), .B0(new_n7984_), .Y(new_n7985_));
  AOI21X1  g07921(.A0(new_n7622_), .A1(new_n2658_), .B0(new_n7985_), .Y(new_n7986_));
  XOR2X1   g07922(.A(new_n7986_), .B(new_n70_), .Y(new_n7987_));
  AOI21X1  g07923(.A0(new_n7987_), .A1(new_n7983_), .B0(new_n7982_), .Y(new_n7988_));
  NOR2X1   g07924(.A(new_n7988_), .B(new_n7829_), .Y(new_n7989_));
  AOI21X1  g07925(.A0(new_n7828_), .A1(new_n7823_), .B0(new_n7989_), .Y(new_n7990_));
  NOR2X1   g07926(.A(new_n7990_), .B(new_n7822_), .Y(new_n7991_));
  XOR2X1   g07927(.A(new_n7990_), .B(new_n7822_), .Y(new_n7992_));
  AOI22X1  g07928(.A0(new_n7657_), .A1(new_n2875_), .B0(new_n7341_), .B1(new_n3146_), .Y(new_n7993_));
  OAI21X1  g07929(.A0(new_n7644_), .A1(new_n3144_), .B0(new_n7993_), .Y(new_n7994_));
  AOI21X1  g07930(.A0(new_n7656_), .A1(new_n2876_), .B0(new_n7994_), .Y(new_n7995_));
  XOR2X1   g07931(.A(new_n7995_), .B(new_n1920_), .Y(new_n7996_));
  AOI21X1  g07932(.A0(new_n7996_), .A1(new_n7992_), .B0(new_n7991_), .Y(new_n7997_));
  NOR2X1   g07933(.A(new_n7997_), .B(new_n7820_), .Y(new_n7998_));
  INVX1    g07934(.A(new_n7998_), .Y(new_n7999_));
  XOR2X1   g07935(.A(new_n7997_), .B(new_n7820_), .Y(new_n8000_));
  INVX1    g07936(.A(new_n8000_), .Y(new_n8001_));
  XOR2X1   g07937(.A(new_n7996_), .B(new_n7992_), .Y(new_n8002_));
  INVX1    g07938(.A(new_n8002_), .Y(new_n8003_));
  XOR2X1   g07939(.A(new_n7987_), .B(new_n7983_), .Y(new_n8004_));
  INVX1    g07940(.A(new_n8004_), .Y(new_n8005_));
  XOR2X1   g07941(.A(new_n7979_), .B(\a[26] ), .Y(new_n8006_));
  XOR2X1   g07942(.A(new_n8006_), .B(new_n7976_), .Y(new_n8007_));
  XOR2X1   g07943(.A(new_n7972_), .B(new_n7840_), .Y(new_n8008_));
  AOI22X1  g07944(.A0(new_n7044_), .A1(new_n2418_), .B0(new_n6818_), .B1(new_n2424_), .Y(new_n8009_));
  OAI21X1  g07945(.A0(new_n7367_), .A1(new_n2626_), .B0(new_n8009_), .Y(new_n8010_));
  AOI21X1  g07946(.A0(new_n7366_), .A1(new_n2301_), .B0(new_n8010_), .Y(new_n8011_));
  XOR2X1   g07947(.A(new_n8011_), .B(\a[26] ), .Y(new_n8012_));
  INVX1    g07948(.A(new_n8012_), .Y(new_n8013_));
  XOR2X1   g07949(.A(new_n8012_), .B(new_n8008_), .Y(new_n8014_));
  XOR2X1   g07950(.A(new_n7970_), .B(new_n7883_), .Y(new_n8015_));
  AOI22X1  g07951(.A0(new_n6882_), .A1(new_n2185_), .B0(new_n6822_), .B1(new_n2095_), .Y(new_n8016_));
  OAI21X1  g07952(.A0(new_n7671_), .A1(new_n2140_), .B0(new_n8016_), .Y(new_n8017_));
  AOI21X1  g07953(.A0(new_n7670_), .A1(new_n2062_), .B0(new_n8017_), .Y(new_n8018_));
  XOR2X1   g07954(.A(new_n8018_), .B(\a[29] ), .Y(new_n8019_));
  INVX1    g07955(.A(new_n8019_), .Y(new_n8020_));
  XOR2X1   g07956(.A(new_n8019_), .B(new_n8015_), .Y(new_n8021_));
  AOI22X1  g07957(.A0(new_n6818_), .A1(new_n2418_), .B0(new_n6745_), .B1(new_n2424_), .Y(new_n8022_));
  OAI21X1  g07958(.A0(new_n7047_), .A1(new_n2626_), .B0(new_n8022_), .Y(new_n8023_));
  AOI21X1  g07959(.A0(new_n7046_), .A1(new_n2301_), .B0(new_n8023_), .Y(new_n8024_));
  XOR2X1   g07960(.A(new_n8024_), .B(\a[26] ), .Y(new_n8025_));
  NOR2X1   g07961(.A(new_n8025_), .B(new_n8021_), .Y(new_n8026_));
  AOI21X1  g07962(.A0(new_n8020_), .A1(new_n8015_), .B0(new_n8026_), .Y(new_n8027_));
  NOR2X1   g07963(.A(new_n8027_), .B(new_n8014_), .Y(new_n8028_));
  AOI21X1  g07964(.A0(new_n8013_), .A1(new_n8008_), .B0(new_n8028_), .Y(new_n8029_));
  NOR2X1   g07965(.A(new_n8029_), .B(new_n8007_), .Y(new_n8030_));
  XOR2X1   g07966(.A(new_n8029_), .B(new_n8007_), .Y(new_n8031_));
  AOI22X1  g07967(.A0(new_n7529_), .A1(new_n2696_), .B0(new_n7522_), .B1(new_n2657_), .Y(new_n8032_));
  OAI21X1  g07968(.A0(new_n7581_), .A1(new_n2753_), .B0(new_n8032_), .Y(new_n8033_));
  AOI21X1  g07969(.A0(new_n7565_), .A1(new_n2658_), .B0(new_n8033_), .Y(new_n8034_));
  XOR2X1   g07970(.A(new_n8034_), .B(new_n70_), .Y(new_n8035_));
  AOI21X1  g07971(.A0(new_n8035_), .A1(new_n8031_), .B0(new_n8030_), .Y(new_n8036_));
  NOR2X1   g07972(.A(new_n8036_), .B(new_n8005_), .Y(new_n8037_));
  INVX1    g07973(.A(new_n8037_), .Y(new_n8038_));
  XOR2X1   g07974(.A(new_n8036_), .B(new_n8005_), .Y(new_n8039_));
  INVX1    g07975(.A(new_n8039_), .Y(new_n8040_));
  AOI22X1  g07976(.A0(new_n7590_), .A1(new_n3099_), .B0(new_n7578_), .B1(new_n2875_), .Y(new_n8041_));
  OAI21X1  g07977(.A0(new_n7642_), .A1(new_n3152_), .B0(new_n8041_), .Y(new_n8042_));
  AOI21X1  g07978(.A0(new_n7712_), .A1(new_n2876_), .B0(new_n8042_), .Y(new_n8043_));
  XOR2X1   g07979(.A(new_n8043_), .B(\a[20] ), .Y(new_n8044_));
  OAI21X1  g07980(.A0(new_n8044_), .A1(new_n8040_), .B0(new_n8038_), .Y(new_n8045_));
  AOI22X1  g07981(.A0(new_n7643_), .A1(new_n3146_), .B0(new_n7590_), .B1(new_n2875_), .Y(new_n8046_));
  OAI21X1  g07982(.A0(new_n7642_), .A1(new_n3144_), .B0(new_n8046_), .Y(new_n8047_));
  AOI21X1  g07983(.A0(new_n7718_), .A1(new_n2876_), .B0(new_n8047_), .Y(new_n8048_));
  XOR2X1   g07984(.A(new_n8048_), .B(\a[20] ), .Y(new_n8049_));
  INVX1    g07985(.A(new_n8049_), .Y(new_n8050_));
  INVX1    g07986(.A(new_n7829_), .Y(new_n8051_));
  XOR2X1   g07987(.A(new_n7988_), .B(new_n8051_), .Y(new_n8052_));
  XOR2X1   g07988(.A(new_n8049_), .B(new_n8045_), .Y(new_n8053_));
  NOR2X1   g07989(.A(new_n8053_), .B(new_n8052_), .Y(new_n8054_));
  AOI21X1  g07990(.A0(new_n8050_), .A1(new_n8045_), .B0(new_n8054_), .Y(new_n8055_));
  NOR2X1   g07991(.A(new_n8055_), .B(new_n8003_), .Y(new_n8056_));
  XOR2X1   g07992(.A(new_n8055_), .B(new_n8002_), .Y(new_n8057_));
  INVX1    g07993(.A(new_n8057_), .Y(new_n8058_));
  XOR2X1   g07994(.A(new_n8035_), .B(new_n8031_), .Y(new_n8059_));
  INVX1    g07995(.A(new_n8059_), .Y(new_n8060_));
  XOR2X1   g07996(.A(new_n8027_), .B(new_n8014_), .Y(new_n8061_));
  AOI22X1  g07997(.A0(new_n7522_), .A1(new_n2696_), .B0(new_n7485_), .B1(new_n2657_), .Y(new_n8062_));
  OAI21X1  g07998(.A0(new_n7537_), .A1(new_n2753_), .B0(new_n8062_), .Y(new_n8063_));
  AOI21X1  g07999(.A0(new_n7536_), .A1(new_n2658_), .B0(new_n8063_), .Y(new_n8064_));
  XOR2X1   g08000(.A(new_n8064_), .B(\a[23] ), .Y(new_n8065_));
  INVX1    g08001(.A(new_n8065_), .Y(new_n8066_));
  XOR2X1   g08002(.A(new_n8065_), .B(new_n8061_), .Y(new_n8067_));
  XOR2X1   g08003(.A(new_n8025_), .B(new_n8021_), .Y(new_n8068_));
  NAND2X1  g08004(.A(new_n7910_), .B(new_n7893_), .Y(new_n8069_));
  AND2X1   g08005(.A(new_n7959_), .B(new_n7911_), .Y(new_n8070_));
  NOR2X1   g08006(.A(new_n7957_), .B(new_n7951_), .Y(new_n8071_));
  NOR2X1   g08007(.A(new_n7958_), .B(new_n8071_), .Y(new_n8072_));
  AOI21X1  g08008(.A0(new_n8070_), .A1(new_n8069_), .B0(new_n8072_), .Y(new_n8073_));
  XOR2X1   g08009(.A(new_n6977_), .B(new_n6976_), .Y(new_n8074_));
  INVX1    g08010(.A(new_n6892_), .Y(new_n8075_));
  AOI22X1  g08011(.A0(new_n6897_), .A1(new_n1890_), .B0(new_n6894_), .B1(new_n1884_), .Y(new_n8076_));
  OAI21X1  g08012(.A0(new_n8075_), .A1(new_n3498_), .B0(new_n8076_), .Y(new_n8077_));
  AOI21X1  g08013(.A0(new_n8074_), .A1(new_n407_), .B0(new_n8077_), .Y(new_n8078_));
  NOR2X1   g08014(.A(new_n8078_), .B(new_n8073_), .Y(new_n8079_));
  INVX1    g08015(.A(new_n8079_), .Y(new_n8080_));
  INVX1    g08016(.A(new_n8073_), .Y(new_n8081_));
  XOR2X1   g08017(.A(new_n8078_), .B(new_n8081_), .Y(new_n8082_));
  INVX1    g08018(.A(new_n7762_), .Y(new_n8083_));
  OAI22X1  g08019(.A0(new_n7885_), .A1(new_n2186_), .B0(new_n7878_), .B1(new_n2431_), .Y(new_n8084_));
  AOI21X1  g08020(.A0(new_n6885_), .A1(new_n2139_), .B0(new_n8084_), .Y(new_n8085_));
  OAI21X1  g08021(.A0(new_n8083_), .A1(new_n2063_), .B0(new_n8085_), .Y(new_n8086_));
  XOR2X1   g08022(.A(new_n8086_), .B(new_n74_), .Y(new_n8087_));
  OAI21X1  g08023(.A0(new_n8087_), .A1(new_n8082_), .B0(new_n8080_), .Y(new_n8088_));
  XOR2X1   g08024(.A(new_n8070_), .B(new_n7892_), .Y(new_n8089_));
  AND2X1   g08025(.A(new_n8089_), .B(new_n8088_), .Y(new_n8090_));
  INVX1    g08026(.A(new_n8088_), .Y(new_n8091_));
  XOR2X1   g08027(.A(new_n8089_), .B(new_n8091_), .Y(new_n8092_));
  AOI22X1  g08028(.A0(new_n6887_), .A1(new_n2185_), .B0(new_n6885_), .B1(new_n2095_), .Y(new_n8093_));
  OAI21X1  g08029(.A0(new_n6884_), .A1(new_n2140_), .B0(new_n8093_), .Y(new_n8094_));
  AOI21X1  g08030(.A0(new_n7771_), .A1(new_n2062_), .B0(new_n8094_), .Y(new_n8095_));
  XOR2X1   g08031(.A(new_n8095_), .B(\a[29] ), .Y(new_n8096_));
  NOR2X1   g08032(.A(new_n8096_), .B(new_n8092_), .Y(new_n8097_));
  XOR2X1   g08033(.A(new_n7969_), .B(new_n7964_), .Y(new_n8098_));
  OAI21X1  g08034(.A0(new_n8097_), .A1(new_n8090_), .B0(new_n8098_), .Y(new_n8099_));
  NOR2X1   g08035(.A(new_n8097_), .B(new_n8090_), .Y(new_n8100_));
  XOR2X1   g08036(.A(new_n8098_), .B(new_n8100_), .Y(new_n8101_));
  AOI22X1  g08037(.A0(new_n6820_), .A1(new_n2424_), .B0(new_n6745_), .B1(new_n2418_), .Y(new_n8102_));
  OAI21X1  g08038(.A0(new_n7361_), .A1(new_n2626_), .B0(new_n8102_), .Y(new_n8103_));
  AOI21X1  g08039(.A0(new_n7404_), .A1(new_n2301_), .B0(new_n8103_), .Y(new_n8104_));
  XOR2X1   g08040(.A(new_n8104_), .B(\a[26] ), .Y(new_n8105_));
  OAI21X1  g08041(.A0(new_n8105_), .A1(new_n8101_), .B0(new_n8099_), .Y(new_n8106_));
  XOR2X1   g08042(.A(new_n8106_), .B(new_n8068_), .Y(new_n8107_));
  AOI22X1  g08043(.A0(new_n7485_), .A1(new_n2696_), .B0(new_n7364_), .B1(new_n2657_), .Y(new_n8108_));
  OAI21X1  g08044(.A0(new_n7523_), .A1(new_n2753_), .B0(new_n8108_), .Y(new_n8109_));
  AOI21X1  g08045(.A0(new_n7612_), .A1(new_n2658_), .B0(new_n8109_), .Y(new_n8110_));
  XOR2X1   g08046(.A(new_n8110_), .B(new_n70_), .Y(new_n8111_));
  AND2X1   g08047(.A(new_n8111_), .B(new_n8107_), .Y(new_n8112_));
  AOI21X1  g08048(.A0(new_n8106_), .A1(new_n8068_), .B0(new_n8112_), .Y(new_n8113_));
  NOR2X1   g08049(.A(new_n8113_), .B(new_n8067_), .Y(new_n8114_));
  AOI21X1  g08050(.A0(new_n8066_), .A1(new_n8061_), .B0(new_n8114_), .Y(new_n8115_));
  NOR2X1   g08051(.A(new_n8115_), .B(new_n8060_), .Y(new_n8116_));
  XOR2X1   g08052(.A(new_n8115_), .B(new_n8060_), .Y(new_n8117_));
  AOI22X1  g08053(.A0(new_n7578_), .A1(new_n3099_), .B0(new_n7571_), .B1(new_n2875_), .Y(new_n8118_));
  OAI21X1  g08054(.A0(new_n7594_), .A1(new_n3152_), .B0(new_n8118_), .Y(new_n8119_));
  AOI21X1  g08055(.A0(new_n7593_), .A1(new_n2876_), .B0(new_n8119_), .Y(new_n8120_));
  XOR2X1   g08056(.A(new_n8120_), .B(new_n1920_), .Y(new_n8121_));
  AOI21X1  g08057(.A0(new_n8121_), .A1(new_n8117_), .B0(new_n8116_), .Y(new_n8122_));
  MX2X1    g08058(.A(new_n3233_), .B(new_n3228_), .S0(new_n3230_), .Y(new_n8123_));
  AOI22X1  g08059(.A0(new_n7643_), .A1(new_n3232_), .B0(new_n8123_), .B1(new_n7341_), .Y(new_n8124_));
  OAI21X1  g08060(.A0(new_n7808_), .A1(new_n3388_), .B0(new_n8124_), .Y(new_n8125_));
  XOR2X1   g08061(.A(new_n8125_), .B(new_n2445_), .Y(new_n8126_));
  NOR2X1   g08062(.A(new_n8126_), .B(new_n8122_), .Y(new_n8127_));
  XOR2X1   g08063(.A(new_n8044_), .B(new_n8039_), .Y(new_n8128_));
  INVX1    g08064(.A(new_n8128_), .Y(new_n8129_));
  XOR2X1   g08065(.A(new_n8126_), .B(new_n8122_), .Y(new_n8130_));
  AOI21X1  g08066(.A0(new_n8130_), .A1(new_n8129_), .B0(new_n8127_), .Y(new_n8131_));
  INVX1    g08067(.A(new_n8131_), .Y(new_n8132_));
  XOR2X1   g08068(.A(new_n8053_), .B(new_n8052_), .Y(new_n8133_));
  AND2X1   g08069(.A(new_n8133_), .B(new_n8132_), .Y(new_n8134_));
  INVX1    g08070(.A(new_n8134_), .Y(new_n8135_));
  XOR2X1   g08071(.A(new_n8130_), .B(new_n8128_), .Y(new_n8136_));
  XOR2X1   g08072(.A(new_n8121_), .B(new_n8117_), .Y(new_n8137_));
  INVX1    g08073(.A(new_n8137_), .Y(new_n8138_));
  XOR2X1   g08074(.A(new_n8113_), .B(new_n8067_), .Y(new_n8139_));
  AOI22X1  g08075(.A0(new_n7571_), .A1(new_n3099_), .B0(new_n7558_), .B1(new_n2875_), .Y(new_n8140_));
  OAI21X1  g08076(.A0(new_n7602_), .A1(new_n3152_), .B0(new_n8140_), .Y(new_n8141_));
  AOI21X1  g08077(.A0(new_n7601_), .A1(new_n2876_), .B0(new_n8141_), .Y(new_n8142_));
  XOR2X1   g08078(.A(new_n8142_), .B(\a[20] ), .Y(new_n8143_));
  INVX1    g08079(.A(new_n8143_), .Y(new_n8144_));
  XOR2X1   g08080(.A(new_n8143_), .B(new_n8139_), .Y(new_n8145_));
  XOR2X1   g08081(.A(new_n8111_), .B(new_n8107_), .Y(new_n8146_));
  INVX1    g08082(.A(new_n8146_), .Y(new_n8147_));
  XOR2X1   g08083(.A(new_n8105_), .B(new_n8101_), .Y(new_n8148_));
  INVX1    g08084(.A(new_n8148_), .Y(new_n8149_));
  XOR2X1   g08085(.A(new_n8096_), .B(new_n8092_), .Y(new_n8150_));
  AOI22X1  g08086(.A0(new_n6822_), .A1(new_n2424_), .B0(new_n6820_), .B1(new_n2418_), .Y(new_n8151_));
  OAI21X1  g08087(.A0(new_n7418_), .A1(new_n2626_), .B0(new_n8151_), .Y(new_n8152_));
  AOI21X1  g08088(.A0(new_n7417_), .A1(new_n2301_), .B0(new_n8152_), .Y(new_n8153_));
  XOR2X1   g08089(.A(new_n8153_), .B(\a[26] ), .Y(new_n8154_));
  INVX1    g08090(.A(new_n8154_), .Y(new_n8155_));
  AND2X1   g08091(.A(new_n8155_), .B(new_n8150_), .Y(new_n8156_));
  XOR2X1   g08092(.A(new_n8154_), .B(new_n8150_), .Y(new_n8157_));
  INVX1    g08093(.A(new_n8157_), .Y(new_n8158_));
  INVX1    g08094(.A(new_n7931_), .Y(new_n8159_));
  INVX1    g08095(.A(new_n1308_), .Y(new_n8160_));
  NOR4X1   g08096(.A(new_n527_), .B(new_n547_), .C(new_n523_), .D(new_n304_), .Y(new_n8161_));
  NOR4X1   g08097(.A(new_n361_), .B(new_n483_), .C(new_n691_), .D(new_n219_), .Y(new_n8162_));
  NOR4X1   g08098(.A(new_n3012_), .B(new_n945_), .C(new_n229_), .D(new_n194_), .Y(new_n8163_));
  NAND3X1  g08099(.A(new_n8163_), .B(new_n8162_), .C(new_n8161_), .Y(new_n8164_));
  OR4X1    g08100(.A(new_n1751_), .B(new_n1478_), .C(new_n1427_), .D(new_n537_), .Y(new_n8165_));
  OR4X1    g08101(.A(new_n8165_), .B(new_n8164_), .C(new_n2076_), .D(new_n416_), .Y(new_n8166_));
  NOR3X1   g08102(.A(new_n8166_), .B(new_n1377_), .C(new_n8160_), .Y(new_n8167_));
  NOR2X1   g08103(.A(new_n8167_), .B(new_n8159_), .Y(new_n8168_));
  NOR3X1   g08104(.A(\a[2] ), .B(\a[1] ), .C(\a[0] ), .Y(new_n8169_));
  INVX1    g08105(.A(new_n8169_), .Y(new_n8170_));
  AOI21X1  g08106(.A0(new_n8170_), .A1(new_n7341_), .B0(new_n3431_), .Y(new_n8171_));
  NOR3X1   g08107(.A(new_n7635_), .B(new_n7106_), .C(new_n7095_), .Y(new_n8172_));
  NOR3X1   g08108(.A(new_n8169_), .B(new_n8172_), .C(\a[2] ), .Y(new_n8173_));
  NAND3X1  g08109(.A(new_n1151_), .B(new_n2150_), .C(new_n820_), .Y(new_n8174_));
  OR4X1    g08110(.A(new_n286_), .B(new_n850_), .C(new_n246_), .D(new_n147_), .Y(new_n8175_));
  OR4X1    g08111(.A(new_n8175_), .B(new_n570_), .C(new_n292_), .D(new_n138_), .Y(new_n8176_));
  OR4X1    g08112(.A(new_n1275_), .B(new_n7923_), .C(new_n382_), .D(new_n231_), .Y(new_n8177_));
  OR4X1    g08113(.A(new_n8177_), .B(new_n8176_), .C(new_n8174_), .D(new_n2087_), .Y(new_n8178_));
  OR4X1    g08114(.A(new_n7896_), .B(new_n1701_), .C(new_n399_), .D(new_n825_), .Y(new_n8179_));
  OR4X1    g08115(.A(new_n7076_), .B(new_n1502_), .C(new_n1336_), .D(new_n1090_), .Y(new_n8180_));
  OR2X1    g08116(.A(new_n8180_), .B(new_n8179_), .Y(new_n8181_));
  OR4X1    g08117(.A(new_n1950_), .B(new_n2097_), .C(new_n772_), .D(new_n422_), .Y(new_n8182_));
  OR4X1    g08118(.A(new_n8182_), .B(new_n516_), .C(new_n470_), .D(new_n354_), .Y(new_n8183_));
  OR4X1    g08119(.A(new_n8183_), .B(new_n8181_), .C(new_n8178_), .D(new_n136_), .Y(new_n8184_));
  OR4X1    g08120(.A(new_n2209_), .B(new_n490_), .C(new_n447_), .D(new_n313_), .Y(new_n8185_));
  OR4X1    g08121(.A(new_n7352_), .B(new_n357_), .C(new_n146_), .D(new_n585_), .Y(new_n8186_));
  OR4X1    g08122(.A(new_n8186_), .B(new_n8185_), .C(new_n3766_), .D(new_n3468_), .Y(new_n8187_));
  NOR4X1   g08123(.A(new_n8187_), .B(new_n8184_), .C(new_n7851_), .D(new_n6775_), .Y(new_n8188_));
  NOR3X1   g08124(.A(new_n8188_), .B(new_n8173_), .C(new_n8171_), .Y(new_n8189_));
  AND2X1   g08125(.A(new_n8170_), .B(new_n7341_), .Y(new_n8190_));
  XOR2X1   g08126(.A(new_n8190_), .B(new_n3431_), .Y(new_n8191_));
  XOR2X1   g08127(.A(new_n8188_), .B(new_n8191_), .Y(new_n8192_));
  INVX1    g08128(.A(new_n8192_), .Y(new_n8193_));
  NAND3X1  g08129(.A(new_n5371_), .B(new_n5369_), .C(new_n5958_), .Y(new_n8194_));
  AND2X1   g08130(.A(new_n8194_), .B(new_n7341_), .Y(new_n8195_));
  XOR2X1   g08131(.A(new_n8195_), .B(new_n3289_), .Y(new_n8196_));
  AOI21X1  g08132(.A0(new_n8196_), .A1(new_n8193_), .B0(new_n8189_), .Y(new_n8197_));
  OR2X1    g08133(.A(new_n8197_), .B(new_n8159_), .Y(new_n8198_));
  XOR2X1   g08134(.A(new_n8197_), .B(new_n7931_), .Y(new_n8199_));
  INVX1    g08135(.A(new_n6904_), .Y(new_n8200_));
  XOR2X1   g08136(.A(new_n8200_), .B(new_n6902_), .Y(new_n8201_));
  AND2X1   g08137(.A(new_n8201_), .B(new_n6966_), .Y(new_n8202_));
  AOI21X1  g08138(.A0(new_n6968_), .A1(new_n6967_), .B0(new_n8202_), .Y(new_n8203_));
  INVX1    g08139(.A(new_n8203_), .Y(new_n8204_));
  INVX1    g08140(.A(new_n6902_), .Y(new_n8205_));
  AOI22X1  g08141(.A0(new_n6906_), .A1(new_n1890_), .B0(new_n6904_), .B1(new_n1884_), .Y(new_n8206_));
  OAI21X1  g08142(.A0(new_n8205_), .A1(new_n3498_), .B0(new_n8206_), .Y(new_n8207_));
  AOI21X1  g08143(.A0(new_n8204_), .A1(new_n407_), .B0(new_n8207_), .Y(new_n8208_));
  OAI21X1  g08144(.A0(new_n8208_), .A1(new_n8199_), .B0(new_n8198_), .Y(new_n8209_));
  XOR2X1   g08145(.A(new_n8167_), .B(new_n8159_), .Y(new_n8210_));
  AND2X1   g08146(.A(new_n8210_), .B(new_n8209_), .Y(new_n8211_));
  XOR2X1   g08147(.A(new_n7949_), .B(new_n7948_), .Y(new_n8212_));
  OAI21X1  g08148(.A0(new_n8211_), .A1(new_n8168_), .B0(new_n8212_), .Y(new_n8213_));
  XOR2X1   g08149(.A(new_n6899_), .B(new_n6897_), .Y(new_n8214_));
  OAI22X1  g08150(.A0(new_n6973_), .A1(new_n6972_), .B0(new_n8214_), .B1(new_n6971_), .Y(new_n8215_));
  AOI22X1  g08151(.A0(new_n6902_), .A1(new_n1890_), .B0(new_n6899_), .B1(new_n1884_), .Y(new_n8216_));
  OAI21X1  g08152(.A0(new_n6898_), .A1(new_n3498_), .B0(new_n8216_), .Y(new_n8217_));
  AOI21X1  g08153(.A0(new_n8215_), .A1(new_n407_), .B0(new_n8217_), .Y(new_n8218_));
  INVX1    g08154(.A(new_n8218_), .Y(new_n8219_));
  OR2X1    g08155(.A(new_n8211_), .B(new_n8168_), .Y(new_n8220_));
  XOR2X1   g08156(.A(new_n8212_), .B(new_n8220_), .Y(new_n8221_));
  NAND2X1  g08157(.A(new_n8221_), .B(new_n8219_), .Y(new_n8222_));
  AND2X1   g08158(.A(new_n8222_), .B(new_n8213_), .Y(new_n8223_));
  INVX1    g08159(.A(new_n8223_), .Y(new_n8224_));
  XOR2X1   g08160(.A(new_n7956_), .B(new_n7952_), .Y(new_n8225_));
  NAND2X1  g08161(.A(new_n8225_), .B(new_n8224_), .Y(new_n8226_));
  XOR2X1   g08162(.A(new_n8225_), .B(new_n8223_), .Y(new_n8227_));
  OAI22X1  g08163(.A0(new_n8075_), .A1(new_n2186_), .B0(new_n7885_), .B1(new_n2431_), .Y(new_n8228_));
  AOI21X1  g08164(.A0(new_n6887_), .A1(new_n2139_), .B0(new_n8228_), .Y(new_n8229_));
  OAI21X1  g08165(.A0(new_n7876_), .A1(new_n2063_), .B0(new_n8229_), .Y(new_n8230_));
  XOR2X1   g08166(.A(new_n8230_), .B(new_n74_), .Y(new_n8231_));
  OAI21X1  g08167(.A0(new_n8231_), .A1(new_n8227_), .B0(new_n8226_), .Y(new_n8232_));
  XOR2X1   g08168(.A(new_n8087_), .B(new_n8082_), .Y(new_n8233_));
  NAND2X1  g08169(.A(new_n8233_), .B(new_n8232_), .Y(new_n8234_));
  XOR2X1   g08170(.A(new_n8233_), .B(new_n8232_), .Y(new_n8235_));
  INVX1    g08171(.A(new_n8235_), .Y(new_n8236_));
  AOI22X1  g08172(.A0(new_n6882_), .A1(new_n2424_), .B0(new_n6822_), .B1(new_n2418_), .Y(new_n8237_));
  OAI21X1  g08173(.A0(new_n7671_), .A1(new_n2626_), .B0(new_n8237_), .Y(new_n8238_));
  AOI21X1  g08174(.A0(new_n7670_), .A1(new_n2301_), .B0(new_n8238_), .Y(new_n8239_));
  XOR2X1   g08175(.A(new_n8239_), .B(\a[26] ), .Y(new_n8240_));
  OAI21X1  g08176(.A0(new_n8240_), .A1(new_n8236_), .B0(new_n8234_), .Y(new_n8241_));
  AOI21X1  g08177(.A0(new_n8241_), .A1(new_n8158_), .B0(new_n8156_), .Y(new_n8242_));
  NOR2X1   g08178(.A(new_n8242_), .B(new_n8149_), .Y(new_n8243_));
  XOR2X1   g08179(.A(new_n8242_), .B(new_n8149_), .Y(new_n8244_));
  AOI22X1  g08180(.A0(new_n7364_), .A1(new_n2696_), .B0(new_n7044_), .B1(new_n2657_), .Y(new_n8245_));
  OAI21X1  g08181(.A0(new_n7504_), .A1(new_n2753_), .B0(new_n8245_), .Y(new_n8246_));
  AOI21X1  g08182(.A0(new_n7552_), .A1(new_n2658_), .B0(new_n8246_), .Y(new_n8247_));
  XOR2X1   g08183(.A(new_n8247_), .B(new_n70_), .Y(new_n8248_));
  AOI21X1  g08184(.A0(new_n8248_), .A1(new_n8244_), .B0(new_n8243_), .Y(new_n8249_));
  NOR2X1   g08185(.A(new_n8249_), .B(new_n8147_), .Y(new_n8250_));
  XOR2X1   g08186(.A(new_n8249_), .B(new_n8147_), .Y(new_n8251_));
  AOI22X1  g08187(.A0(new_n7558_), .A1(new_n3099_), .B0(new_n7529_), .B1(new_n2875_), .Y(new_n8252_));
  OAI21X1  g08188(.A0(new_n7623_), .A1(new_n3152_), .B0(new_n8252_), .Y(new_n8253_));
  AOI21X1  g08189(.A0(new_n7622_), .A1(new_n2876_), .B0(new_n8253_), .Y(new_n8254_));
  XOR2X1   g08190(.A(new_n8254_), .B(new_n1920_), .Y(new_n8255_));
  AOI21X1  g08191(.A0(new_n8255_), .A1(new_n8251_), .B0(new_n8250_), .Y(new_n8256_));
  NOR2X1   g08192(.A(new_n8256_), .B(new_n8145_), .Y(new_n8257_));
  AOI21X1  g08193(.A0(new_n8144_), .A1(new_n8139_), .B0(new_n8257_), .Y(new_n8258_));
  NOR2X1   g08194(.A(new_n8258_), .B(new_n8138_), .Y(new_n8259_));
  XOR2X1   g08195(.A(new_n8258_), .B(new_n8138_), .Y(new_n8260_));
  AOI22X1  g08196(.A0(new_n7657_), .A1(new_n3232_), .B0(new_n7341_), .B1(new_n3546_), .Y(new_n8261_));
  OAI21X1  g08197(.A0(new_n7644_), .A1(new_n3389_), .B0(new_n8261_), .Y(new_n8262_));
  AOI21X1  g08198(.A0(new_n7656_), .A1(new_n3234_), .B0(new_n8262_), .Y(new_n8263_));
  XOR2X1   g08199(.A(new_n8263_), .B(new_n2445_), .Y(new_n8264_));
  AOI21X1  g08200(.A0(new_n8264_), .A1(new_n8260_), .B0(new_n8259_), .Y(new_n8265_));
  NOR2X1   g08201(.A(new_n8265_), .B(new_n8136_), .Y(new_n8266_));
  XOR2X1   g08202(.A(new_n8265_), .B(new_n8136_), .Y(new_n8267_));
  XOR2X1   g08203(.A(new_n8264_), .B(new_n8260_), .Y(new_n8268_));
  INVX1    g08204(.A(new_n8268_), .Y(new_n8269_));
  XOR2X1   g08205(.A(new_n8255_), .B(new_n8251_), .Y(new_n8270_));
  INVX1    g08206(.A(new_n8270_), .Y(new_n8271_));
  XOR2X1   g08207(.A(new_n8248_), .B(new_n8244_), .Y(new_n8272_));
  XOR2X1   g08208(.A(new_n8241_), .B(new_n8158_), .Y(new_n8273_));
  AOI22X1  g08209(.A0(new_n7044_), .A1(new_n2696_), .B0(new_n6818_), .B1(new_n2657_), .Y(new_n8274_));
  OAI21X1  g08210(.A0(new_n7367_), .A1(new_n2753_), .B0(new_n8274_), .Y(new_n8275_));
  AOI21X1  g08211(.A0(new_n7366_), .A1(new_n2658_), .B0(new_n8275_), .Y(new_n8276_));
  XOR2X1   g08212(.A(new_n8276_), .B(\a[23] ), .Y(new_n8277_));
  INVX1    g08213(.A(new_n8277_), .Y(new_n8278_));
  AND2X1   g08214(.A(new_n8278_), .B(new_n8273_), .Y(new_n8279_));
  XOR2X1   g08215(.A(new_n8277_), .B(new_n8273_), .Y(new_n8280_));
  XOR2X1   g08216(.A(new_n8240_), .B(new_n8235_), .Y(new_n8281_));
  XOR2X1   g08217(.A(new_n8221_), .B(new_n8218_), .Y(new_n8282_));
  AOI22X1  g08218(.A0(new_n6894_), .A1(new_n2185_), .B0(new_n6892_), .B1(new_n2095_), .Y(new_n8283_));
  OAI21X1  g08219(.A0(new_n7885_), .A1(new_n2140_), .B0(new_n8283_), .Y(new_n8284_));
  AOI21X1  g08220(.A0(new_n7884_), .A1(new_n2062_), .B0(new_n8284_), .Y(new_n8285_));
  XOR2X1   g08221(.A(new_n8285_), .B(\a[29] ), .Y(new_n8286_));
  OR2X1    g08222(.A(new_n8286_), .B(new_n8282_), .Y(new_n8287_));
  XOR2X1   g08223(.A(new_n8286_), .B(new_n8282_), .Y(new_n8288_));
  INVX1    g08224(.A(new_n8288_), .Y(new_n8289_));
  INVX1    g08225(.A(new_n8210_), .Y(new_n8290_));
  AOI21X1  g08226(.A0(new_n8167_), .A1(new_n8159_), .B0(new_n8220_), .Y(new_n8291_));
  AOI21X1  g08227(.A0(new_n8290_), .A1(new_n8209_), .B0(new_n8291_), .Y(new_n8292_));
  XOR2X1   g08228(.A(new_n6970_), .B(new_n6968_), .Y(new_n8293_));
  NOR2X1   g08229(.A(new_n8293_), .B(new_n3178_), .Y(new_n8294_));
  INVX1    g08230(.A(new_n6899_), .Y(new_n8295_));
  AOI22X1  g08231(.A0(new_n6904_), .A1(new_n1890_), .B0(new_n6902_), .B1(new_n1884_), .Y(new_n8296_));
  OAI21X1  g08232(.A0(new_n8295_), .A1(new_n3498_), .B0(new_n8296_), .Y(new_n8297_));
  NOR2X1   g08233(.A(new_n8297_), .B(new_n8294_), .Y(new_n8298_));
  NOR2X1   g08234(.A(new_n8298_), .B(new_n8292_), .Y(new_n8299_));
  XOR2X1   g08235(.A(new_n8298_), .B(new_n8292_), .Y(new_n8300_));
  OAI21X1  g08236(.A0(new_n8169_), .A1(new_n8172_), .B0(\a[2] ), .Y(new_n8301_));
  NAND3X1  g08237(.A(new_n8170_), .B(new_n7341_), .C(new_n3431_), .Y(new_n8302_));
  OR4X1    g08238(.A(new_n226_), .B(new_n536_), .C(new_n1008_), .D(new_n307_), .Y(new_n8303_));
  OR2X1    g08239(.A(new_n7345_), .B(new_n76_), .Y(new_n8304_));
  OR4X1    g08240(.A(new_n509_), .B(new_n565_), .C(new_n176_), .D(new_n664_), .Y(new_n8305_));
  OR4X1    g08241(.A(new_n400_), .B(new_n245_), .C(new_n581_), .D(new_n142_), .Y(new_n8306_));
  OR4X1    g08242(.A(new_n8306_), .B(new_n8305_), .C(new_n8304_), .D(new_n8303_), .Y(new_n8307_));
  OR4X1    g08243(.A(new_n8307_), .B(new_n3298_), .C(new_n1746_), .D(new_n958_), .Y(new_n8308_));
  NOR4X1   g08244(.A(new_n8308_), .B(new_n2253_), .C(new_n2225_), .D(new_n801_), .Y(new_n8309_));
  AOI21X1  g08245(.A0(new_n8302_), .A1(new_n8301_), .B0(new_n8309_), .Y(new_n8310_));
  INVX1    g08246(.A(new_n8310_), .Y(new_n8311_));
  NOR3X1   g08247(.A(new_n7425_), .B(new_n659_), .C(new_n460_), .Y(new_n8312_));
  INVX1    g08248(.A(new_n8312_), .Y(new_n8313_));
  OR4X1    g08249(.A(new_n2451_), .B(new_n1385_), .C(new_n1320_), .D(new_n1259_), .Y(new_n8314_));
  OR2X1    g08250(.A(new_n8314_), .B(new_n7067_), .Y(new_n8315_));
  OR4X1    g08251(.A(new_n513_), .B(new_n417_), .C(new_n568_), .D(new_n272_), .Y(new_n8316_));
  OR4X1    g08252(.A(new_n252_), .B(new_n243_), .C(new_n233_), .D(new_n194_), .Y(new_n8317_));
  OR4X1    g08253(.A(new_n8317_), .B(new_n396_), .C(new_n296_), .D(new_n196_), .Y(new_n8318_));
  OR4X1    g08254(.A(new_n8318_), .B(new_n8316_), .C(new_n712_), .D(new_n620_), .Y(new_n8319_));
  NOR4X1   g08255(.A(new_n8319_), .B(new_n8315_), .C(new_n8313_), .D(new_n8184_), .Y(new_n8320_));
  AOI21X1  g08256(.A0(new_n8302_), .A1(new_n8301_), .B0(new_n8320_), .Y(new_n8321_));
  OR4X1    g08257(.A(new_n1540_), .B(new_n451_), .C(new_n423_), .D(new_n681_), .Y(new_n8322_));
  OR4X1    g08258(.A(new_n224_), .B(new_n223_), .C(new_n648_), .D(new_n981_), .Y(new_n8323_));
  OR4X1    g08259(.A(new_n8323_), .B(new_n504_), .C(new_n420_), .D(new_n138_), .Y(new_n8324_));
  OR4X1    g08260(.A(new_n8324_), .B(new_n8322_), .C(new_n6779_), .D(new_n2950_), .Y(new_n8325_));
  OR4X1    g08261(.A(new_n1530_), .B(new_n1173_), .C(new_n116_), .D(new_n307_), .Y(new_n8326_));
  OR4X1    g08262(.A(new_n8326_), .B(new_n497_), .C(new_n383_), .D(new_n358_), .Y(new_n8327_));
  OR2X1    g08263(.A(new_n8327_), .B(new_n1283_), .Y(new_n8328_));
  OR2X1    g08264(.A(new_n8328_), .B(new_n8325_), .Y(new_n8329_));
  OR4X1    g08265(.A(new_n245_), .B(new_n178_), .C(new_n147_), .D(new_n521_), .Y(new_n8330_));
  OR4X1    g08266(.A(new_n8330_), .B(new_n510_), .C(new_n792_), .D(new_n585_), .Y(new_n8331_));
  NOR3X1   g08267(.A(new_n1028_), .B(new_n848_), .C(new_n475_), .Y(new_n8332_));
  NOR4X1   g08268(.A(new_n422_), .B(new_n418_), .C(new_n396_), .D(new_n111_), .Y(new_n8333_));
  NAND3X1  g08269(.A(new_n8333_), .B(new_n8332_), .C(new_n2110_), .Y(new_n8334_));
  OAI22X1  g08270(.A0(new_n152_), .A1(new_n127_), .B0(new_n119_), .B1(new_n90_), .Y(new_n8335_));
  OR2X1    g08271(.A(new_n8335_), .B(new_n546_), .Y(new_n8336_));
  OR4X1    g08272(.A(new_n239_), .B(new_n184_), .C(new_n664_), .D(new_n449_), .Y(new_n8337_));
  OR4X1    g08273(.A(new_n8337_), .B(new_n8336_), .C(new_n7896_), .D(new_n1128_), .Y(new_n8338_));
  OR4X1    g08274(.A(new_n1777_), .B(new_n550_), .C(new_n265_), .D(new_n264_), .Y(new_n8339_));
  NOR4X1   g08275(.A(new_n8339_), .B(new_n8338_), .C(new_n8334_), .D(new_n1291_), .Y(new_n8340_));
  INVX1    g08276(.A(new_n8340_), .Y(new_n8341_));
  NOR4X1   g08277(.A(new_n8341_), .B(new_n8331_), .C(new_n8329_), .D(new_n353_), .Y(new_n8342_));
  INVX1    g08278(.A(new_n8342_), .Y(new_n8343_));
  OAI21X1  g08279(.A0(new_n8173_), .A1(new_n8171_), .B0(new_n8343_), .Y(new_n8344_));
  NOR3X1   g08280(.A(new_n8343_), .B(new_n8173_), .C(new_n8171_), .Y(new_n8345_));
  XOR2X1   g08281(.A(new_n6913_), .B(new_n6911_), .Y(new_n8346_));
  OR2X1    g08282(.A(new_n8346_), .B(new_n6955_), .Y(new_n8347_));
  OAI21X1  g08283(.A0(new_n6957_), .A1(new_n6956_), .B0(new_n8347_), .Y(new_n8348_));
  INVX1    g08284(.A(new_n6911_), .Y(new_n8349_));
  AOI22X1  g08285(.A0(new_n6915_), .A1(new_n1890_), .B0(new_n6913_), .B1(new_n1884_), .Y(new_n8350_));
  OAI21X1  g08286(.A0(new_n8349_), .A1(new_n3498_), .B0(new_n8350_), .Y(new_n8351_));
  AOI21X1  g08287(.A0(new_n8348_), .A1(new_n407_), .B0(new_n8351_), .Y(new_n8352_));
  OAI21X1  g08288(.A0(new_n8352_), .A1(new_n8345_), .B0(new_n8344_), .Y(new_n8353_));
  NAND3X1  g08289(.A(new_n8320_), .B(new_n8302_), .C(new_n8301_), .Y(new_n8354_));
  AOI21X1  g08290(.A0(new_n8354_), .A1(new_n8353_), .B0(new_n8321_), .Y(new_n8355_));
  NAND3X1  g08291(.A(new_n8309_), .B(new_n8302_), .C(new_n8301_), .Y(new_n8356_));
  INVX1    g08292(.A(new_n8356_), .Y(new_n8357_));
  OAI21X1  g08293(.A0(new_n8357_), .A1(new_n8355_), .B0(new_n8311_), .Y(new_n8358_));
  XOR2X1   g08294(.A(new_n8196_), .B(new_n8192_), .Y(new_n8359_));
  XOR2X1   g08295(.A(new_n8359_), .B(new_n8358_), .Y(new_n8360_));
  OR2X1    g08296(.A(new_n6906_), .B(new_n6904_), .Y(new_n8361_));
  INVX1    g08297(.A(new_n6966_), .Y(new_n8362_));
  AOI21X1  g08298(.A0(new_n8361_), .A1(new_n6908_), .B0(new_n6963_), .Y(new_n8363_));
  AOI21X1  g08299(.A0(new_n8362_), .A1(new_n8361_), .B0(new_n8363_), .Y(new_n8364_));
  INVX1    g08300(.A(new_n8364_), .Y(new_n8365_));
  AOI22X1  g08301(.A0(new_n6909_), .A1(new_n1890_), .B0(new_n6906_), .B1(new_n1884_), .Y(new_n8366_));
  OAI21X1  g08302(.A0(new_n8200_), .A1(new_n3498_), .B0(new_n8366_), .Y(new_n8367_));
  AOI21X1  g08303(.A0(new_n8365_), .A1(new_n407_), .B0(new_n8367_), .Y(new_n8368_));
  OR2X1    g08304(.A(new_n8320_), .B(new_n8191_), .Y(new_n8369_));
  AOI21X1  g08305(.A0(new_n8302_), .A1(new_n8301_), .B0(new_n8342_), .Y(new_n8370_));
  NAND3X1  g08306(.A(new_n8342_), .B(new_n8302_), .C(new_n8301_), .Y(new_n8371_));
  INVX1    g08307(.A(new_n8352_), .Y(new_n8372_));
  AOI21X1  g08308(.A0(new_n8372_), .A1(new_n8371_), .B0(new_n8370_), .Y(new_n8373_));
  AND2X1   g08309(.A(new_n8320_), .B(new_n8191_), .Y(new_n8374_));
  OAI21X1  g08310(.A0(new_n8374_), .A1(new_n8373_), .B0(new_n8369_), .Y(new_n8375_));
  AOI21X1  g08311(.A0(new_n8356_), .A1(new_n8375_), .B0(new_n8310_), .Y(new_n8376_));
  OR2X1    g08312(.A(new_n8359_), .B(new_n8376_), .Y(new_n8377_));
  OAI21X1  g08313(.A0(new_n8368_), .A1(new_n8360_), .B0(new_n8377_), .Y(new_n8378_));
  XOR2X1   g08314(.A(new_n8208_), .B(new_n8199_), .Y(new_n8379_));
  NAND2X1  g08315(.A(new_n8379_), .B(new_n8378_), .Y(new_n8380_));
  OR2X1    g08316(.A(new_n8379_), .B(new_n8378_), .Y(new_n8381_));
  NAND2X1  g08317(.A(new_n8381_), .B(new_n8380_), .Y(new_n8382_));
  INVX1    g08318(.A(new_n7953_), .Y(new_n8383_));
  OAI22X1  g08319(.A0(new_n8295_), .A1(new_n2186_), .B0(new_n6898_), .B1(new_n2431_), .Y(new_n8384_));
  AOI21X1  g08320(.A0(new_n6894_), .A1(new_n2139_), .B0(new_n8384_), .Y(new_n8385_));
  OAI21X1  g08321(.A0(new_n8383_), .A1(new_n2063_), .B0(new_n8385_), .Y(new_n8386_));
  XOR2X1   g08322(.A(new_n8386_), .B(new_n74_), .Y(new_n8387_));
  OAI21X1  g08323(.A0(new_n8387_), .A1(new_n8382_), .B0(new_n8380_), .Y(new_n8388_));
  AOI21X1  g08324(.A0(new_n8388_), .A1(new_n8300_), .B0(new_n8299_), .Y(new_n8389_));
  OAI21X1  g08325(.A0(new_n8389_), .A1(new_n8289_), .B0(new_n8287_), .Y(new_n8390_));
  XOR2X1   g08326(.A(new_n8231_), .B(new_n8227_), .Y(new_n8391_));
  NAND2X1  g08327(.A(new_n8391_), .B(new_n8390_), .Y(new_n8392_));
  XOR2X1   g08328(.A(new_n8391_), .B(new_n8390_), .Y(new_n8393_));
  INVX1    g08329(.A(new_n8393_), .Y(new_n8394_));
  AOI22X1  g08330(.A0(new_n6885_), .A1(new_n2424_), .B0(new_n6882_), .B1(new_n2418_), .Y(new_n8395_));
  OAI21X1  g08331(.A0(new_n7472_), .A1(new_n2626_), .B0(new_n8395_), .Y(new_n8396_));
  AOI21X1  g08332(.A0(new_n7471_), .A1(new_n2301_), .B0(new_n8396_), .Y(new_n8397_));
  XOR2X1   g08333(.A(new_n8397_), .B(\a[26] ), .Y(new_n8398_));
  OAI21X1  g08334(.A0(new_n8398_), .A1(new_n8394_), .B0(new_n8392_), .Y(new_n8399_));
  INVX1    g08335(.A(new_n8399_), .Y(new_n8400_));
  OR2X1    g08336(.A(new_n8400_), .B(new_n8281_), .Y(new_n8401_));
  XOR2X1   g08337(.A(new_n8399_), .B(new_n8281_), .Y(new_n8402_));
  AOI22X1  g08338(.A0(new_n6818_), .A1(new_n2696_), .B0(new_n6745_), .B1(new_n2657_), .Y(new_n8403_));
  OAI21X1  g08339(.A0(new_n7047_), .A1(new_n2753_), .B0(new_n8403_), .Y(new_n8404_));
  AOI21X1  g08340(.A0(new_n7046_), .A1(new_n2658_), .B0(new_n8404_), .Y(new_n8405_));
  XOR2X1   g08341(.A(new_n8405_), .B(\a[23] ), .Y(new_n8406_));
  OR2X1    g08342(.A(new_n8406_), .B(new_n8402_), .Y(new_n8407_));
  AND2X1   g08343(.A(new_n8407_), .B(new_n8401_), .Y(new_n8408_));
  NOR2X1   g08344(.A(new_n8408_), .B(new_n8280_), .Y(new_n8409_));
  OAI21X1  g08345(.A0(new_n8409_), .A1(new_n8279_), .B0(new_n8272_), .Y(new_n8410_));
  AOI21X1  g08346(.A0(new_n8278_), .A1(new_n8273_), .B0(new_n8409_), .Y(new_n8411_));
  XOR2X1   g08347(.A(new_n8411_), .B(new_n8272_), .Y(new_n8412_));
  AOI22X1  g08348(.A0(new_n7529_), .A1(new_n3099_), .B0(new_n7522_), .B1(new_n2875_), .Y(new_n8413_));
  OAI21X1  g08349(.A0(new_n7581_), .A1(new_n3152_), .B0(new_n8413_), .Y(new_n8414_));
  AOI21X1  g08350(.A0(new_n7565_), .A1(new_n2876_), .B0(new_n8414_), .Y(new_n8415_));
  XOR2X1   g08351(.A(new_n8415_), .B(\a[20] ), .Y(new_n8416_));
  OR2X1    g08352(.A(new_n8416_), .B(new_n8412_), .Y(new_n8417_));
  AOI21X1  g08353(.A0(new_n8417_), .A1(new_n8410_), .B0(new_n8271_), .Y(new_n8418_));
  INVX1    g08354(.A(new_n8418_), .Y(new_n8419_));
  AND2X1   g08355(.A(new_n8417_), .B(new_n8410_), .Y(new_n8420_));
  AND2X1   g08356(.A(new_n8420_), .B(new_n8271_), .Y(new_n8421_));
  AOI22X1  g08357(.A0(new_n7590_), .A1(new_n3390_), .B0(new_n7578_), .B1(new_n3232_), .Y(new_n8422_));
  OAI21X1  g08358(.A0(new_n7642_), .A1(new_n3545_), .B0(new_n8422_), .Y(new_n8423_));
  AOI21X1  g08359(.A0(new_n7712_), .A1(new_n3234_), .B0(new_n8423_), .Y(new_n8424_));
  XOR2X1   g08360(.A(new_n8424_), .B(\a[17] ), .Y(new_n8425_));
  OAI21X1  g08361(.A0(new_n8425_), .A1(new_n8421_), .B0(new_n8419_), .Y(new_n8426_));
  AOI22X1  g08362(.A0(new_n7643_), .A1(new_n3546_), .B0(new_n7590_), .B1(new_n3232_), .Y(new_n8427_));
  OAI21X1  g08363(.A0(new_n7642_), .A1(new_n3389_), .B0(new_n8427_), .Y(new_n8428_));
  AOI21X1  g08364(.A0(new_n7718_), .A1(new_n3234_), .B0(new_n8428_), .Y(new_n8429_));
  XOR2X1   g08365(.A(new_n8429_), .B(\a[17] ), .Y(new_n8430_));
  INVX1    g08366(.A(new_n8430_), .Y(new_n8431_));
  INVX1    g08367(.A(new_n8145_), .Y(new_n8432_));
  XOR2X1   g08368(.A(new_n8256_), .B(new_n8432_), .Y(new_n8433_));
  XOR2X1   g08369(.A(new_n8430_), .B(new_n8426_), .Y(new_n8434_));
  NOR2X1   g08370(.A(new_n8434_), .B(new_n8433_), .Y(new_n8435_));
  AOI21X1  g08371(.A0(new_n8431_), .A1(new_n8426_), .B0(new_n8435_), .Y(new_n8436_));
  NOR2X1   g08372(.A(new_n8436_), .B(new_n8269_), .Y(new_n8437_));
  INVX1    g08373(.A(new_n8437_), .Y(new_n8438_));
  XOR2X1   g08374(.A(new_n8436_), .B(new_n8268_), .Y(new_n8439_));
  XOR2X1   g08375(.A(new_n8416_), .B(new_n8412_), .Y(new_n8440_));
  INVX1    g08376(.A(new_n8440_), .Y(new_n8441_));
  XOR2X1   g08377(.A(new_n8408_), .B(new_n8280_), .Y(new_n8442_));
  AOI22X1  g08378(.A0(new_n7522_), .A1(new_n3099_), .B0(new_n7485_), .B1(new_n2875_), .Y(new_n8443_));
  OAI21X1  g08379(.A0(new_n7537_), .A1(new_n3152_), .B0(new_n8443_), .Y(new_n8444_));
  AOI21X1  g08380(.A0(new_n7536_), .A1(new_n2876_), .B0(new_n8444_), .Y(new_n8445_));
  XOR2X1   g08381(.A(new_n8445_), .B(\a[20] ), .Y(new_n8446_));
  INVX1    g08382(.A(new_n8446_), .Y(new_n8447_));
  XOR2X1   g08383(.A(new_n8446_), .B(new_n8442_), .Y(new_n8448_));
  INVX1    g08384(.A(new_n8406_), .Y(new_n8449_));
  XOR2X1   g08385(.A(new_n8449_), .B(new_n8402_), .Y(new_n8450_));
  XOR2X1   g08386(.A(new_n8398_), .B(new_n8393_), .Y(new_n8451_));
  XOR2X1   g08387(.A(new_n8389_), .B(new_n8289_), .Y(new_n8452_));
  AOI22X1  g08388(.A0(new_n6887_), .A1(new_n2424_), .B0(new_n6885_), .B1(new_n2418_), .Y(new_n8453_));
  OAI21X1  g08389(.A0(new_n6884_), .A1(new_n2626_), .B0(new_n8453_), .Y(new_n8454_));
  AOI21X1  g08390(.A0(new_n7771_), .A1(new_n2301_), .B0(new_n8454_), .Y(new_n8455_));
  XOR2X1   g08391(.A(new_n8455_), .B(new_n89_), .Y(new_n8456_));
  XOR2X1   g08392(.A(new_n8455_), .B(\a[26] ), .Y(new_n8457_));
  XOR2X1   g08393(.A(new_n8457_), .B(new_n8452_), .Y(new_n8458_));
  INVX1    g08394(.A(new_n8298_), .Y(new_n8459_));
  XOR2X1   g08395(.A(new_n8459_), .B(new_n8292_), .Y(new_n8460_));
  XOR2X1   g08396(.A(new_n8388_), .B(new_n8460_), .Y(new_n8461_));
  AOI22X1  g08397(.A0(new_n6897_), .A1(new_n2185_), .B0(new_n6894_), .B1(new_n2095_), .Y(new_n8462_));
  OAI21X1  g08398(.A0(new_n8075_), .A1(new_n2140_), .B0(new_n8462_), .Y(new_n8463_));
  AOI21X1  g08399(.A0(new_n8074_), .A1(new_n2062_), .B0(new_n8463_), .Y(new_n8464_));
  XOR2X1   g08400(.A(new_n8464_), .B(\a[29] ), .Y(new_n8465_));
  NOR2X1   g08401(.A(new_n8465_), .B(new_n8461_), .Y(new_n8466_));
  XOR2X1   g08402(.A(new_n8465_), .B(new_n8461_), .Y(new_n8467_));
  AOI22X1  g08403(.A0(new_n6890_), .A1(new_n2424_), .B0(new_n6887_), .B1(new_n2418_), .Y(new_n8468_));
  OAI21X1  g08404(.A0(new_n6886_), .A1(new_n2626_), .B0(new_n8468_), .Y(new_n8469_));
  AOI21X1  g08405(.A0(new_n7762_), .A1(new_n2301_), .B0(new_n8469_), .Y(new_n8470_));
  XOR2X1   g08406(.A(new_n8470_), .B(\a[26] ), .Y(new_n8471_));
  INVX1    g08407(.A(new_n8471_), .Y(new_n8472_));
  AOI21X1  g08408(.A0(new_n8472_), .A1(new_n8467_), .B0(new_n8466_), .Y(new_n8473_));
  NOR2X1   g08409(.A(new_n8473_), .B(new_n8458_), .Y(new_n8474_));
  AOI21X1  g08410(.A0(new_n8456_), .A1(new_n8452_), .B0(new_n8474_), .Y(new_n8475_));
  NOR2X1   g08411(.A(new_n8475_), .B(new_n8451_), .Y(new_n8476_));
  XOR2X1   g08412(.A(new_n8475_), .B(new_n8451_), .Y(new_n8477_));
  AOI22X1  g08413(.A0(new_n6820_), .A1(new_n2657_), .B0(new_n6745_), .B1(new_n2696_), .Y(new_n8478_));
  OAI21X1  g08414(.A0(new_n7361_), .A1(new_n2753_), .B0(new_n8478_), .Y(new_n8479_));
  AOI21X1  g08415(.A0(new_n7404_), .A1(new_n2658_), .B0(new_n8479_), .Y(new_n8480_));
  XOR2X1   g08416(.A(new_n8480_), .B(\a[23] ), .Y(new_n8481_));
  INVX1    g08417(.A(new_n8481_), .Y(new_n8482_));
  AOI21X1  g08418(.A0(new_n8482_), .A1(new_n8477_), .B0(new_n8476_), .Y(new_n8483_));
  NOR2X1   g08419(.A(new_n8483_), .B(new_n8450_), .Y(new_n8484_));
  XOR2X1   g08420(.A(new_n8483_), .B(new_n8450_), .Y(new_n8485_));
  AOI22X1  g08421(.A0(new_n7485_), .A1(new_n3099_), .B0(new_n7364_), .B1(new_n2875_), .Y(new_n8486_));
  OAI21X1  g08422(.A0(new_n7523_), .A1(new_n3152_), .B0(new_n8486_), .Y(new_n8487_));
  AOI21X1  g08423(.A0(new_n7612_), .A1(new_n2876_), .B0(new_n8487_), .Y(new_n8488_));
  XOR2X1   g08424(.A(new_n8488_), .B(\a[20] ), .Y(new_n8489_));
  INVX1    g08425(.A(new_n8489_), .Y(new_n8490_));
  AOI21X1  g08426(.A0(new_n8490_), .A1(new_n8485_), .B0(new_n8484_), .Y(new_n8491_));
  NOR2X1   g08427(.A(new_n8491_), .B(new_n8448_), .Y(new_n8492_));
  AOI21X1  g08428(.A0(new_n8447_), .A1(new_n8442_), .B0(new_n8492_), .Y(new_n8493_));
  NOR2X1   g08429(.A(new_n8493_), .B(new_n8441_), .Y(new_n8494_));
  XOR2X1   g08430(.A(new_n8493_), .B(new_n8441_), .Y(new_n8495_));
  AOI22X1  g08431(.A0(new_n7578_), .A1(new_n3390_), .B0(new_n7571_), .B1(new_n3232_), .Y(new_n8496_));
  OAI21X1  g08432(.A0(new_n7594_), .A1(new_n3545_), .B0(new_n8496_), .Y(new_n8497_));
  AOI21X1  g08433(.A0(new_n7593_), .A1(new_n3234_), .B0(new_n8497_), .Y(new_n8498_));
  XOR2X1   g08434(.A(new_n8498_), .B(\a[17] ), .Y(new_n8499_));
  INVX1    g08435(.A(new_n8499_), .Y(new_n8500_));
  AOI21X1  g08436(.A0(new_n8500_), .A1(new_n8495_), .B0(new_n8494_), .Y(new_n8501_));
  MX2X1    g08437(.A(new_n3623_), .B(new_n3625_), .S0(new_n3621_), .Y(new_n8502_));
  AOI22X1  g08438(.A0(new_n7643_), .A1(new_n3628_), .B0(new_n8502_), .B1(new_n7341_), .Y(new_n8503_));
  OAI21X1  g08439(.A0(new_n7808_), .A1(new_n3906_), .B0(new_n8503_), .Y(new_n8504_));
  XOR2X1   g08440(.A(new_n8504_), .B(new_n2529_), .Y(new_n8505_));
  NOR2X1   g08441(.A(new_n8505_), .B(new_n8501_), .Y(new_n8506_));
  XOR2X1   g08442(.A(new_n8420_), .B(new_n8271_), .Y(new_n8507_));
  XOR2X1   g08443(.A(new_n8425_), .B(new_n8507_), .Y(new_n8508_));
  INVX1    g08444(.A(new_n8508_), .Y(new_n8509_));
  XOR2X1   g08445(.A(new_n8505_), .B(new_n8501_), .Y(new_n8510_));
  AOI21X1  g08446(.A0(new_n8510_), .A1(new_n8509_), .B0(new_n8506_), .Y(new_n8511_));
  INVX1    g08447(.A(new_n8511_), .Y(new_n8512_));
  XOR2X1   g08448(.A(new_n8434_), .B(new_n8433_), .Y(new_n8513_));
  AND2X1   g08449(.A(new_n8513_), .B(new_n8512_), .Y(new_n8514_));
  XOR2X1   g08450(.A(new_n8510_), .B(new_n8508_), .Y(new_n8515_));
  XOR2X1   g08451(.A(new_n8499_), .B(new_n8495_), .Y(new_n8516_));
  XOR2X1   g08452(.A(new_n8491_), .B(new_n8448_), .Y(new_n8517_));
  AOI22X1  g08453(.A0(new_n7571_), .A1(new_n3390_), .B0(new_n7558_), .B1(new_n3232_), .Y(new_n8518_));
  OAI21X1  g08454(.A0(new_n7602_), .A1(new_n3545_), .B0(new_n8518_), .Y(new_n8519_));
  AOI21X1  g08455(.A0(new_n7601_), .A1(new_n3234_), .B0(new_n8519_), .Y(new_n8520_));
  XOR2X1   g08456(.A(new_n8520_), .B(\a[17] ), .Y(new_n8521_));
  INVX1    g08457(.A(new_n8521_), .Y(new_n8522_));
  XOR2X1   g08458(.A(new_n8521_), .B(new_n8517_), .Y(new_n8523_));
  XOR2X1   g08459(.A(new_n8489_), .B(new_n8485_), .Y(new_n8524_));
  XOR2X1   g08460(.A(new_n8481_), .B(new_n8477_), .Y(new_n8525_));
  XOR2X1   g08461(.A(new_n8473_), .B(new_n8458_), .Y(new_n8526_));
  AOI22X1  g08462(.A0(new_n6822_), .A1(new_n2657_), .B0(new_n6820_), .B1(new_n2696_), .Y(new_n8527_));
  OAI21X1  g08463(.A0(new_n7418_), .A1(new_n2753_), .B0(new_n8527_), .Y(new_n8528_));
  AOI21X1  g08464(.A0(new_n7417_), .A1(new_n2658_), .B0(new_n8528_), .Y(new_n8529_));
  XOR2X1   g08465(.A(new_n8529_), .B(new_n70_), .Y(new_n8530_));
  XOR2X1   g08466(.A(new_n8529_), .B(\a[23] ), .Y(new_n8531_));
  XOR2X1   g08467(.A(new_n8531_), .B(new_n8526_), .Y(new_n8532_));
  XOR2X1   g08468(.A(new_n8471_), .B(new_n8467_), .Y(new_n8533_));
  XOR2X1   g08469(.A(new_n8309_), .B(new_n8191_), .Y(new_n8534_));
  NOR2X1   g08470(.A(new_n8534_), .B(new_n8355_), .Y(new_n8535_));
  AOI21X1  g08471(.A0(new_n8376_), .A1(new_n8356_), .B0(new_n8535_), .Y(new_n8536_));
  NOR2X1   g08472(.A(new_n6909_), .B(new_n6906_), .Y(new_n8537_));
  INVX1    g08473(.A(new_n6963_), .Y(new_n8538_));
  NAND2X1  g08474(.A(new_n6959_), .B(new_n6912_), .Y(new_n8539_));
  NAND2X1  g08475(.A(new_n6961_), .B(new_n8539_), .Y(new_n8540_));
  OAI21X1  g08476(.A0(new_n8538_), .A1(new_n8537_), .B0(new_n8540_), .Y(new_n8541_));
  AOI22X1  g08477(.A0(new_n6911_), .A1(new_n1890_), .B0(new_n6909_), .B1(new_n1884_), .Y(new_n8542_));
  OAI21X1  g08478(.A0(new_n6964_), .A1(new_n3498_), .B0(new_n8542_), .Y(new_n8543_));
  AOI21X1  g08479(.A0(new_n8541_), .A1(new_n407_), .B0(new_n8543_), .Y(new_n8544_));
  OR2X1    g08480(.A(new_n8544_), .B(new_n8536_), .Y(new_n8545_));
  OAI22X1  g08481(.A0(new_n8358_), .A1(new_n8357_), .B0(new_n8534_), .B1(new_n8355_), .Y(new_n8546_));
  XOR2X1   g08482(.A(new_n8544_), .B(new_n8546_), .Y(new_n8547_));
  XOR2X1   g08483(.A(new_n8190_), .B(\a[2] ), .Y(new_n8548_));
  XOR2X1   g08484(.A(new_n8320_), .B(new_n8548_), .Y(new_n8549_));
  AND2X1   g08485(.A(new_n8549_), .B(new_n8353_), .Y(new_n8550_));
  NOR3X1   g08486(.A(new_n8374_), .B(new_n8353_), .C(new_n8321_), .Y(new_n8551_));
  OR2X1    g08487(.A(new_n8551_), .B(new_n8550_), .Y(new_n8552_));
  XOR2X1   g08488(.A(new_n6958_), .B(new_n6957_), .Y(new_n8553_));
  AOI22X1  g08489(.A0(new_n6913_), .A1(new_n1890_), .B0(new_n6911_), .B1(new_n1884_), .Y(new_n8554_));
  OAI21X1  g08490(.A0(new_n6960_), .A1(new_n3498_), .B0(new_n8554_), .Y(new_n8555_));
  AOI21X1  g08491(.A0(new_n8553_), .A1(new_n407_), .B0(new_n8555_), .Y(new_n8556_));
  INVX1    g08492(.A(new_n8556_), .Y(new_n8557_));
  OAI21X1  g08493(.A0(new_n8551_), .A1(new_n8550_), .B0(new_n8556_), .Y(new_n8558_));
  NAND2X1  g08494(.A(new_n8549_), .B(new_n8353_), .Y(new_n8559_));
  NAND3X1  g08495(.A(new_n8354_), .B(new_n8373_), .C(new_n8369_), .Y(new_n8560_));
  NAND3X1  g08496(.A(new_n8557_), .B(new_n8560_), .C(new_n8559_), .Y(new_n8561_));
  OAI21X1  g08497(.A0(new_n8345_), .A1(new_n8370_), .B0(new_n8372_), .Y(new_n8562_));
  NAND3X1  g08498(.A(new_n8352_), .B(new_n8371_), .C(new_n8344_), .Y(new_n8563_));
  OR4X1    g08499(.A(new_n1778_), .B(new_n1426_), .C(new_n514_), .D(new_n441_), .Y(new_n8564_));
  OR2X1    g08500(.A(new_n8564_), .B(new_n1525_), .Y(new_n8565_));
  INVX1    g08501(.A(new_n547_), .Y(new_n8566_));
  NAND3X1  g08502(.A(new_n8566_), .B(new_n987_), .C(new_n2395_), .Y(new_n8567_));
  OR4X1    g08503(.A(new_n8567_), .B(new_n7249_), .C(new_n578_), .D(new_n173_), .Y(new_n8568_));
  OAI22X1  g08504(.A0(new_n105_), .A1(new_n102_), .B0(new_n92_), .B1(new_n75_), .Y(new_n8569_));
  OR2X1    g08505(.A(new_n8569_), .B(new_n423_), .Y(new_n8570_));
  OR4X1    g08506(.A(new_n234_), .B(new_n200_), .C(new_n184_), .D(new_n120_), .Y(new_n8571_));
  OR4X1    g08507(.A(new_n8571_), .B(new_n8570_), .C(new_n1961_), .D(new_n1743_), .Y(new_n8572_));
  NOR4X1   g08508(.A(new_n8572_), .B(new_n8568_), .C(new_n8565_), .D(new_n7845_), .Y(new_n8573_));
  NAND3X1  g08509(.A(new_n8573_), .B(new_n2820_), .C(new_n644_), .Y(new_n8574_));
  INVX1    g08510(.A(new_n8574_), .Y(new_n8575_));
  INVX1    g08511(.A(new_n6952_), .Y(new_n8576_));
  XOR2X1   g08512(.A(new_n6953_), .B(new_n8576_), .Y(new_n8577_));
  INVX1    g08513(.A(new_n8577_), .Y(new_n8578_));
  INVX1    g08514(.A(new_n6913_), .Y(new_n8579_));
  XOR2X1   g08515(.A(new_n6717_), .B(new_n5670_), .Y(new_n8580_));
  AOI22X1  g08516(.A0(new_n8580_), .A1(new_n1890_), .B0(new_n6915_), .B1(new_n1884_), .Y(new_n8581_));
  OAI21X1  g08517(.A0(new_n8579_), .A1(new_n3498_), .B0(new_n8581_), .Y(new_n8582_));
  AOI21X1  g08518(.A0(new_n8578_), .A1(new_n407_), .B0(new_n8582_), .Y(new_n8583_));
  NOR2X1   g08519(.A(new_n8583_), .B(new_n8575_), .Y(new_n8584_));
  INVX1    g08520(.A(new_n8584_), .Y(new_n8585_));
  OR4X1    g08521(.A(new_n321_), .B(new_n206_), .C(new_n825_), .D(new_n172_), .Y(new_n8586_));
  OR4X1    g08522(.A(new_n399_), .B(new_n479_), .C(new_n226_), .D(new_n521_), .Y(new_n8587_));
  OR4X1    g08523(.A(new_n8587_), .B(new_n8586_), .C(new_n935_), .D(new_n834_), .Y(new_n8588_));
  OR4X1    g08524(.A(new_n1911_), .B(new_n1779_), .C(new_n1724_), .D(new_n1597_), .Y(new_n8589_));
  NOR4X1   g08525(.A(new_n8589_), .B(new_n8588_), .C(new_n7183_), .D(new_n3437_), .Y(new_n8590_));
  NAND3X1  g08526(.A(new_n8590_), .B(new_n859_), .C(new_n593_), .Y(new_n8591_));
  INVX1    g08527(.A(new_n8591_), .Y(new_n8592_));
  NAND2X1  g08528(.A(new_n6918_), .B(new_n6917_), .Y(new_n8593_));
  AOI21X1  g08529(.A0(new_n8593_), .A1(new_n6919_), .B0(new_n6950_), .Y(new_n8594_));
  AOI21X1  g08530(.A0(new_n6918_), .A1(new_n6917_), .B0(new_n6952_), .Y(new_n8595_));
  OAI21X1  g08531(.A0(new_n8595_), .A1(new_n8594_), .B0(new_n407_), .Y(new_n8596_));
  OAI22X1  g08532(.A0(new_n6920_), .A1(new_n2245_), .B0(new_n6918_), .B1(new_n1885_), .Y(new_n8597_));
  AOI21X1  g08533(.A0(new_n6915_), .A1(new_n1889_), .B0(new_n8597_), .Y(new_n8598_));
  AOI21X1  g08534(.A0(new_n8598_), .A1(new_n8596_), .B0(new_n8592_), .Y(new_n8599_));
  INVX1    g08535(.A(new_n8599_), .Y(new_n8600_));
  NOR3X1   g08536(.A(new_n8331_), .B(new_n8328_), .C(new_n8325_), .Y(new_n8601_));
  NAND3X1  g08537(.A(new_n2353_), .B(new_n1175_), .C(new_n145_), .Y(new_n8602_));
  OR4X1    g08538(.A(new_n493_), .B(new_n398_), .C(new_n651_), .D(new_n1579_), .Y(new_n8603_));
  OR4X1    g08539(.A(new_n408_), .B(new_n304_), .C(new_n819_), .D(new_n216_), .Y(new_n8604_));
  OR4X1    g08540(.A(new_n8604_), .B(new_n8603_), .C(new_n1191_), .D(new_n882_), .Y(new_n8605_));
  NOR3X1   g08541(.A(new_n8605_), .B(new_n8602_), .C(new_n1662_), .Y(new_n8606_));
  NAND3X1  g08542(.A(new_n8606_), .B(new_n8601_), .C(new_n1279_), .Y(new_n8607_));
  INVX1    g08543(.A(new_n8607_), .Y(new_n8608_));
  XOR2X1   g08544(.A(new_n6920_), .B(new_n8580_), .Y(new_n8609_));
  AND2X1   g08545(.A(new_n8609_), .B(new_n6948_), .Y(new_n8610_));
  AOI21X1  g08546(.A0(new_n6950_), .A1(new_n6949_), .B0(new_n8610_), .Y(new_n8611_));
  INVX1    g08547(.A(new_n8611_), .Y(new_n8612_));
  AOI22X1  g08548(.A0(new_n6923_), .A1(new_n1890_), .B0(new_n6922_), .B1(new_n1884_), .Y(new_n8613_));
  OAI21X1  g08549(.A0(new_n6918_), .A1(new_n3498_), .B0(new_n8613_), .Y(new_n8614_));
  AOI21X1  g08550(.A0(new_n8612_), .A1(new_n407_), .B0(new_n8614_), .Y(new_n8615_));
  NOR2X1   g08551(.A(new_n8615_), .B(new_n8608_), .Y(new_n8616_));
  INVX1    g08552(.A(new_n8616_), .Y(new_n8617_));
  NOR2X1   g08553(.A(new_n6792_), .B(new_n6788_), .Y(new_n8618_));
  NOR4X1   g08554(.A(new_n496_), .B(new_n224_), .C(new_n206_), .D(new_n303_), .Y(new_n8619_));
  NOR4X1   g08555(.A(new_n717_), .B(new_n746_), .C(new_n379_), .D(new_n118_), .Y(new_n8620_));
  NAND4X1  g08556(.A(new_n8620_), .B(new_n8619_), .C(new_n3781_), .D(new_n1175_), .Y(new_n8621_));
  OR4X1    g08557(.A(new_n1082_), .B(new_n457_), .C(new_n149_), .D(new_n114_), .Y(new_n8622_));
  OR4X1    g08558(.A(new_n8622_), .B(new_n723_), .C(new_n417_), .D(new_n220_), .Y(new_n8623_));
  OR4X1    g08559(.A(new_n8623_), .B(new_n1386_), .C(new_n1211_), .D(new_n1142_), .Y(new_n8624_));
  NOR4X1   g08560(.A(new_n8624_), .B(new_n8621_), .C(new_n2102_), .D(new_n1988_), .Y(new_n8625_));
  NAND3X1  g08561(.A(new_n8625_), .B(new_n8618_), .C(new_n3816_), .Y(new_n8626_));
  INVX1    g08562(.A(new_n8626_), .Y(new_n8627_));
  XOR2X1   g08563(.A(new_n6947_), .B(new_n6946_), .Y(new_n8628_));
  AOI22X1  g08564(.A0(new_n6925_), .A1(new_n1890_), .B0(new_n6923_), .B1(new_n1884_), .Y(new_n8629_));
  OAI21X1  g08565(.A0(new_n6920_), .A1(new_n3498_), .B0(new_n8629_), .Y(new_n8630_));
  AOI21X1  g08566(.A0(new_n8628_), .A1(new_n407_), .B0(new_n8630_), .Y(new_n8631_));
  NOR2X1   g08567(.A(new_n8631_), .B(new_n8627_), .Y(new_n8632_));
  INVX1    g08568(.A(new_n8632_), .Y(new_n8633_));
  OR4X1    g08569(.A(new_n7917_), .B(new_n3782_), .C(new_n2997_), .D(new_n2358_), .Y(new_n8634_));
  OR4X1    g08570(.A(new_n1703_), .B(new_n823_), .C(new_n724_), .D(new_n386_), .Y(new_n8635_));
  OR4X1    g08571(.A(new_n574_), .B(new_n193_), .C(new_n178_), .D(new_n160_), .Y(new_n8636_));
  OR4X1    g08572(.A(new_n8636_), .B(new_n8635_), .C(new_n803_), .D(new_n427_), .Y(new_n8637_));
  NOR3X1   g08573(.A(new_n8637_), .B(new_n8634_), .C(new_n2355_), .Y(new_n8638_));
  OR4X1    g08574(.A(new_n681_), .B(new_n213_), .C(new_n200_), .D(new_n196_), .Y(new_n8639_));
  OR4X1    g08575(.A(new_n8639_), .B(new_n723_), .C(new_n509_), .D(new_n371_), .Y(new_n8640_));
  OR2X1    g08576(.A(new_n88_), .B(new_n81_), .Y(new_n8641_));
  NAND3X1  g08577(.A(new_n214_), .B(new_n380_), .C(new_n8641_), .Y(new_n8642_));
  OR4X1    g08578(.A(new_n8642_), .B(new_n1090_), .C(new_n632_), .D(new_n357_), .Y(new_n8643_));
  OR2X1    g08579(.A(new_n8643_), .B(new_n8640_), .Y(new_n8644_));
  OR4X1    g08580(.A(new_n2451_), .B(new_n1136_), .C(new_n227_), .D(new_n224_), .Y(new_n8645_));
  NOR4X1   g08581(.A(new_n8645_), .B(new_n8644_), .C(new_n3734_), .D(new_n1967_), .Y(new_n8646_));
  OR4X1    g08582(.A(new_n586_), .B(new_n417_), .C(new_n264_), .D(new_n164_), .Y(new_n8647_));
  OR4X1    g08583(.A(new_n420_), .B(new_n300_), .C(new_n299_), .D(new_n292_), .Y(new_n8648_));
  OAI22X1  g08584(.A0(new_n182_), .A1(new_n69_), .B0(new_n81_), .B1(new_n75_), .Y(new_n8649_));
  OR4X1    g08585(.A(new_n8649_), .B(new_n8648_), .C(new_n8647_), .D(new_n222_), .Y(new_n8650_));
  OR2X1    g08586(.A(new_n3685_), .B(new_n1721_), .Y(new_n8651_));
  NOR3X1   g08587(.A(new_n7021_), .B(new_n840_), .C(new_n1046_), .Y(new_n8652_));
  INVX1    g08588(.A(new_n8652_), .Y(new_n8653_));
  OR4X1    g08589(.A(new_n1759_), .B(new_n1002_), .C(new_n280_), .D(new_n928_), .Y(new_n8654_));
  OR2X1    g08590(.A(new_n8654_), .B(new_n8653_), .Y(new_n8655_));
  NOR4X1   g08591(.A(new_n8655_), .B(new_n8651_), .C(new_n8650_), .D(new_n7753_), .Y(new_n8656_));
  NAND3X1  g08592(.A(new_n8656_), .B(new_n8646_), .C(new_n8638_), .Y(new_n8657_));
  INVX1    g08593(.A(new_n8657_), .Y(new_n8658_));
  XOR2X1   g08594(.A(new_n6714_), .B(new_n6859_), .Y(new_n8659_));
  XOR2X1   g08595(.A(new_n6925_), .B(new_n8659_), .Y(new_n8660_));
  AND2X1   g08596(.A(new_n8660_), .B(new_n6944_), .Y(new_n8661_));
  AOI21X1  g08597(.A0(new_n6946_), .A1(new_n6945_), .B0(new_n8661_), .Y(new_n8662_));
  INVX1    g08598(.A(new_n8662_), .Y(new_n8663_));
  AOI22X1  g08599(.A0(new_n6927_), .A1(new_n1890_), .B0(new_n6925_), .B1(new_n1884_), .Y(new_n8664_));
  OAI21X1  g08600(.A0(new_n8659_), .A1(new_n3498_), .B0(new_n8664_), .Y(new_n8665_));
  AOI21X1  g08601(.A0(new_n8663_), .A1(new_n407_), .B0(new_n8665_), .Y(new_n8666_));
  NOR2X1   g08602(.A(new_n8666_), .B(new_n8658_), .Y(new_n8667_));
  INVX1    g08603(.A(new_n8667_), .Y(new_n8668_));
  NOR4X1   g08604(.A(new_n261_), .B(new_n224_), .C(new_n187_), .D(new_n337_), .Y(new_n8669_));
  NAND3X1  g08605(.A(new_n8669_), .B(new_n7187_), .C(new_n7079_), .Y(new_n8670_));
  OR4X1    g08606(.A(new_n659_), .B(new_n652_), .C(new_n490_), .D(new_n272_), .Y(new_n8671_));
  OR4X1    g08607(.A(new_n8671_), .B(new_n1646_), .C(new_n1336_), .D(new_n931_), .Y(new_n8672_));
  NOR4X1   g08608(.A(new_n8672_), .B(new_n8670_), .C(new_n7934_), .D(new_n997_), .Y(new_n8673_));
  INVX1    g08609(.A(new_n8673_), .Y(new_n8674_));
  OR4X1    g08610(.A(new_n1416_), .B(new_n873_), .C(new_n716_), .D(new_n188_), .Y(new_n8675_));
  OAI22X1  g08611(.A0(new_n152_), .A1(new_n99_), .B0(new_n125_), .B1(new_n119_), .Y(new_n8676_));
  OR2X1    g08612(.A(new_n8676_), .B(new_n408_), .Y(new_n8677_));
  OR4X1    g08613(.A(new_n296_), .B(new_n398_), .C(new_n141_), .D(new_n1008_), .Y(new_n8678_));
  OR4X1    g08614(.A(new_n8678_), .B(new_n8677_), .C(new_n8675_), .D(new_n1315_), .Y(new_n8679_));
  NOR4X1   g08615(.A(new_n8679_), .B(new_n8674_), .C(new_n7087_), .D(new_n7074_), .Y(new_n8680_));
  XOR2X1   g08616(.A(new_n6927_), .B(new_n6925_), .Y(new_n8681_));
  OAI22X1  g08617(.A0(new_n6944_), .A1(new_n6943_), .B0(new_n8681_), .B1(new_n6942_), .Y(new_n8682_));
  INVX1    g08618(.A(new_n6925_), .Y(new_n8683_));
  AOI22X1  g08619(.A0(new_n6932_), .A1(new_n1890_), .B0(new_n6927_), .B1(new_n1884_), .Y(new_n8684_));
  OAI21X1  g08620(.A0(new_n8683_), .A1(new_n3498_), .B0(new_n8684_), .Y(new_n8685_));
  AOI21X1  g08621(.A0(new_n8682_), .A1(new_n407_), .B0(new_n8685_), .Y(new_n8686_));
  NOR2X1   g08622(.A(new_n8686_), .B(new_n8680_), .Y(new_n8687_));
  INVX1    g08623(.A(new_n8687_), .Y(new_n8688_));
  OR4X1    g08624(.A(new_n396_), .B(new_n747_), .C(new_n717_), .D(new_n240_), .Y(new_n8689_));
  OR4X1    g08625(.A(new_n494_), .B(new_n327_), .C(new_n648_), .D(new_n158_), .Y(new_n8690_));
  OR4X1    g08626(.A(new_n8690_), .B(new_n8689_), .C(new_n188_), .D(new_n187_), .Y(new_n8691_));
  OR4X1    g08627(.A(new_n7376_), .B(new_n356_), .C(new_n199_), .D(new_n100_), .Y(new_n8692_));
  OR4X1    g08628(.A(new_n8692_), .B(new_n857_), .C(new_n743_), .D(new_n537_), .Y(new_n8693_));
  OR4X1    g08629(.A(new_n3283_), .B(new_n259_), .C(new_n616_), .D(new_n147_), .Y(new_n8694_));
  OR4X1    g08630(.A(new_n8694_), .B(new_n527_), .C(new_n348_), .D(new_n400_), .Y(new_n8695_));
  NOR4X1   g08631(.A(new_n8695_), .B(new_n8693_), .C(new_n8691_), .D(new_n7905_), .Y(new_n8696_));
  INVX1    g08632(.A(new_n8696_), .Y(new_n8697_));
  OAI22X1  g08633(.A0(new_n123_), .A1(new_n94_), .B0(new_n115_), .B1(new_n81_), .Y(new_n8698_));
  OR4X1    g08634(.A(new_n468_), .B(new_n819_), .C(new_n651_), .D(new_n1284_), .Y(new_n8699_));
  OR4X1    g08635(.A(new_n8699_), .B(new_n8698_), .C(new_n724_), .D(new_n363_), .Y(new_n8700_));
  OR4X1    g08636(.A(new_n1514_), .B(new_n1096_), .C(new_n612_), .D(new_n191_), .Y(new_n8701_));
  OR4X1    g08637(.A(new_n8701_), .B(new_n8700_), .C(new_n2786_), .D(new_n549_), .Y(new_n8702_));
  NOR4X1   g08638(.A(new_n8702_), .B(new_n8697_), .C(new_n1544_), .D(new_n7015_), .Y(new_n8703_));
  XOR2X1   g08639(.A(new_n6930_), .B(new_n6927_), .Y(new_n8704_));
  XOR2X1   g08640(.A(new_n8704_), .B(new_n6940_), .Y(new_n8705_));
  INVX1    g08641(.A(new_n8705_), .Y(new_n8706_));
  AOI22X1  g08642(.A0(new_n6933_), .A1(new_n1890_), .B0(new_n6932_), .B1(new_n1884_), .Y(new_n8707_));
  OAI21X1  g08643(.A0(new_n6929_), .A1(new_n3498_), .B0(new_n8707_), .Y(new_n8708_));
  AOI21X1  g08644(.A0(new_n8706_), .A1(new_n407_), .B0(new_n8708_), .Y(new_n8709_));
  NOR2X1   g08645(.A(new_n8709_), .B(new_n8703_), .Y(new_n8710_));
  OR4X1    g08646(.A(new_n2315_), .B(new_n686_), .C(new_n815_), .D(new_n274_), .Y(new_n8711_));
  OR4X1    g08647(.A(new_n589_), .B(new_n196_), .C(new_n156_), .D(new_n155_), .Y(new_n8712_));
  OR4X1    g08648(.A(new_n594_), .B(new_n395_), .C(new_n321_), .D(new_n535_), .Y(new_n8713_));
  OR4X1    g08649(.A(new_n8713_), .B(new_n8712_), .C(new_n1974_), .D(new_n1473_), .Y(new_n8714_));
  OR4X1    g08650(.A(new_n8714_), .B(new_n8711_), .C(new_n3703_), .D(new_n3045_), .Y(new_n8715_));
  NOR4X1   g08651(.A(new_n8715_), .B(new_n7173_), .C(new_n7144_), .D(new_n1958_), .Y(new_n8716_));
  XOR2X1   g08652(.A(new_n6939_), .B(new_n6938_), .Y(new_n8717_));
  AOI22X1  g08653(.A0(new_n6935_), .A1(new_n1890_), .B0(new_n6933_), .B1(new_n1884_), .Y(new_n8718_));
  OAI21X1  g08654(.A0(new_n6930_), .A1(new_n3498_), .B0(new_n8718_), .Y(new_n8719_));
  AOI21X1  g08655(.A0(new_n8717_), .A1(new_n407_), .B0(new_n8719_), .Y(new_n8720_));
  NOR2X1   g08656(.A(new_n8720_), .B(new_n8716_), .Y(new_n8721_));
  NOR4X1   g08657(.A(new_n1158_), .B(new_n1118_), .C(new_n904_), .D(new_n827_), .Y(new_n8722_));
  OR4X1    g08658(.A(new_n293_), .B(new_n239_), .C(new_n202_), .D(new_n521_), .Y(new_n8723_));
  NOR4X1   g08659(.A(new_n8723_), .B(new_n631_), .C(new_n184_), .D(new_n181_), .Y(new_n8724_));
  NOR4X1   g08660(.A(new_n739_), .B(new_n395_), .C(new_n307_), .D(new_n86_), .Y(new_n8725_));
  NAND3X1  g08661(.A(new_n8725_), .B(new_n8724_), .C(new_n8722_), .Y(new_n8726_));
  AOI21X1  g08662(.A0(new_n108_), .A1(new_n99_), .B0(new_n119_), .Y(new_n8727_));
  OR2X1    g08663(.A(new_n8727_), .B(new_n1044_), .Y(new_n8728_));
  OR4X1    g08664(.A(new_n8728_), .B(new_n7058_), .C(new_n2950_), .D(new_n1875_), .Y(new_n8729_));
  NOR3X1   g08665(.A(new_n2101_), .B(new_n1005_), .C(new_n638_), .Y(new_n8730_));
  NOR4X1   g08666(.A(new_n478_), .B(new_n321_), .C(new_n180_), .D(new_n173_), .Y(new_n8731_));
  NOR4X1   g08667(.A(new_n354_), .B(new_n218_), .C(new_n581_), .D(new_n149_), .Y(new_n8732_));
  NAND3X1  g08668(.A(new_n8732_), .B(new_n8731_), .C(new_n8730_), .Y(new_n8733_));
  OR4X1    g08669(.A(new_n8733_), .B(new_n8729_), .C(new_n8726_), .D(new_n8334_), .Y(new_n8734_));
  OR2X1    g08670(.A(new_n8734_), .B(new_n7901_), .Y(new_n8735_));
  NOR3X1   g08671(.A(new_n500_), .B(new_n206_), .C(new_n202_), .Y(new_n8736_));
  NOR3X1   g08672(.A(new_n720_), .B(new_n421_), .C(new_n365_), .Y(new_n8737_));
  NOR3X1   g08673(.A(new_n1515_), .B(new_n196_), .C(new_n410_), .Y(new_n8738_));
  NAND3X1  g08674(.A(new_n8738_), .B(new_n8737_), .C(new_n8736_), .Y(new_n8739_));
  OR4X1    g08675(.A(new_n1402_), .B(new_n743_), .C(new_n498_), .D(new_n154_), .Y(new_n8740_));
  OR4X1    g08676(.A(new_n679_), .B(new_n387_), .C(new_n474_), .D(new_n1046_), .Y(new_n8741_));
  OR4X1    g08677(.A(new_n8741_), .B(new_n8740_), .C(new_n8739_), .D(new_n1921_), .Y(new_n8742_));
  OR4X1    g08678(.A(new_n8742_), .B(new_n8623_), .C(new_n7200_), .D(new_n2310_), .Y(new_n8743_));
  OAI22X1  g08679(.A0(new_n161_), .A1(new_n123_), .B0(new_n152_), .B1(new_n129_), .Y(new_n8744_));
  OR4X1    g08680(.A(new_n8744_), .B(new_n1540_), .C(new_n1223_), .D(new_n1118_), .Y(new_n8745_));
  NOR4X1   g08681(.A(new_n8745_), .B(new_n1044_), .C(new_n396_), .D(new_n356_), .Y(new_n8746_));
  OR4X1    g08682(.A(new_n2272_), .B(new_n1478_), .C(new_n441_), .D(new_n539_), .Y(new_n8747_));
  NOR4X1   g08683(.A(new_n8747_), .B(new_n1458_), .C(new_n1457_), .D(new_n1442_), .Y(new_n8748_));
  NAND3X1  g08684(.A(new_n8748_), .B(new_n8746_), .C(new_n3757_), .Y(new_n8749_));
  NOR4X1   g08685(.A(new_n8749_), .B(new_n8743_), .C(new_n1604_), .D(new_n1603_), .Y(new_n8750_));
  XOR2X1   g08686(.A(new_n6937_), .B(new_n6935_), .Y(new_n8751_));
  INVX1    g08687(.A(new_n6935_), .Y(new_n8752_));
  OAI22X1  g08688(.A0(new_n6936_), .A1(new_n1885_), .B0(new_n8752_), .B1(new_n3498_), .Y(new_n8753_));
  AOI21X1  g08689(.A0(new_n8751_), .A1(new_n407_), .B0(new_n8753_), .Y(new_n8754_));
  NOR2X1   g08690(.A(new_n8754_), .B(new_n8750_), .Y(new_n8755_));
  AND2X1   g08691(.A(new_n8755_), .B(new_n8735_), .Y(new_n8756_));
  XOR2X1   g08692(.A(new_n6854_), .B(new_n6704_), .Y(new_n8757_));
  AND2X1   g08693(.A(new_n6936_), .B(new_n6935_), .Y(new_n8758_));
  XOR2X1   g08694(.A(new_n8758_), .B(new_n8757_), .Y(new_n8759_));
  OAI22X1  g08695(.A0(new_n6936_), .A1(new_n2245_), .B0(new_n8752_), .B1(new_n1885_), .Y(new_n8760_));
  AOI21X1  g08696(.A0(new_n6933_), .A1(new_n1889_), .B0(new_n8760_), .Y(new_n8761_));
  OAI21X1  g08697(.A0(new_n8759_), .A1(new_n3178_), .B0(new_n8761_), .Y(new_n8762_));
  XOR2X1   g08698(.A(new_n8755_), .B(new_n8735_), .Y(new_n8763_));
  AOI21X1  g08699(.A0(new_n8763_), .A1(new_n8762_), .B0(new_n8756_), .Y(new_n8764_));
  INVX1    g08700(.A(new_n8716_), .Y(new_n8765_));
  XOR2X1   g08701(.A(new_n8720_), .B(new_n8765_), .Y(new_n8766_));
  NOR2X1   g08702(.A(new_n8766_), .B(new_n8764_), .Y(new_n8767_));
  NOR2X1   g08703(.A(new_n8767_), .B(new_n8721_), .Y(new_n8768_));
  INVX1    g08704(.A(new_n8768_), .Y(new_n8769_));
  XOR2X1   g08705(.A(new_n8709_), .B(new_n8703_), .Y(new_n8770_));
  AOI21X1  g08706(.A0(new_n8770_), .A1(new_n8769_), .B0(new_n8710_), .Y(new_n8771_));
  XOR2X1   g08707(.A(new_n8686_), .B(new_n8680_), .Y(new_n8772_));
  INVX1    g08708(.A(new_n8772_), .Y(new_n8773_));
  OAI21X1  g08709(.A0(new_n8773_), .A1(new_n8771_), .B0(new_n8688_), .Y(new_n8774_));
  INVX1    g08710(.A(new_n8774_), .Y(new_n8775_));
  XOR2X1   g08711(.A(new_n8666_), .B(new_n8657_), .Y(new_n8776_));
  OAI21X1  g08712(.A0(new_n8776_), .A1(new_n8775_), .B0(new_n8668_), .Y(new_n8777_));
  INVX1    g08713(.A(new_n8777_), .Y(new_n8778_));
  XOR2X1   g08714(.A(new_n8631_), .B(new_n8626_), .Y(new_n8779_));
  OAI21X1  g08715(.A0(new_n8779_), .A1(new_n8778_), .B0(new_n8633_), .Y(new_n8780_));
  INVX1    g08716(.A(new_n8780_), .Y(new_n8781_));
  XOR2X1   g08717(.A(new_n8615_), .B(new_n8607_), .Y(new_n8782_));
  OAI21X1  g08718(.A0(new_n8782_), .A1(new_n8781_), .B0(new_n8617_), .Y(new_n8783_));
  INVX1    g08719(.A(new_n8783_), .Y(new_n8784_));
  AND2X1   g08720(.A(new_n8598_), .B(new_n8596_), .Y(new_n8785_));
  XOR2X1   g08721(.A(new_n8785_), .B(new_n8591_), .Y(new_n8786_));
  OAI21X1  g08722(.A0(new_n8786_), .A1(new_n8784_), .B0(new_n8600_), .Y(new_n8787_));
  INVX1    g08723(.A(new_n8787_), .Y(new_n8788_));
  XOR2X1   g08724(.A(new_n8583_), .B(new_n8574_), .Y(new_n8789_));
  OAI21X1  g08725(.A0(new_n8789_), .A1(new_n8788_), .B0(new_n8585_), .Y(new_n8790_));
  INVX1    g08726(.A(new_n8790_), .Y(new_n8791_));
  AOI21X1  g08727(.A0(new_n8563_), .A1(new_n8562_), .B0(new_n8791_), .Y(new_n8792_));
  NAND3X1  g08728(.A(new_n8791_), .B(new_n8563_), .C(new_n8562_), .Y(new_n8793_));
  OAI22X1  g08729(.A0(new_n6960_), .A1(new_n2186_), .B0(new_n6964_), .B1(new_n2431_), .Y(new_n8794_));
  AOI21X1  g08730(.A0(new_n6904_), .A1(new_n2139_), .B0(new_n8794_), .Y(new_n8795_));
  OAI21X1  g08731(.A0(new_n8364_), .A1(new_n2063_), .B0(new_n8795_), .Y(new_n8796_));
  XOR2X1   g08732(.A(new_n8796_), .B(new_n74_), .Y(new_n8797_));
  INVX1    g08733(.A(new_n8797_), .Y(new_n8798_));
  AOI21X1  g08734(.A0(new_n8798_), .A1(new_n8793_), .B0(new_n8792_), .Y(new_n8799_));
  AOI21X1  g08735(.A0(new_n8561_), .A1(new_n8558_), .B0(new_n8799_), .Y(new_n8800_));
  AOI21X1  g08736(.A0(new_n8557_), .A1(new_n8552_), .B0(new_n8800_), .Y(new_n8801_));
  OAI21X1  g08737(.A0(new_n8801_), .A1(new_n8547_), .B0(new_n8545_), .Y(new_n8802_));
  XOR2X1   g08738(.A(new_n8368_), .B(new_n8360_), .Y(new_n8803_));
  AND2X1   g08739(.A(new_n8803_), .B(new_n8802_), .Y(new_n8804_));
  XOR2X1   g08740(.A(new_n8803_), .B(new_n8802_), .Y(new_n8805_));
  AOI22X1  g08741(.A0(new_n6902_), .A1(new_n2185_), .B0(new_n6899_), .B1(new_n2095_), .Y(new_n8806_));
  OAI21X1  g08742(.A0(new_n6898_), .A1(new_n2140_), .B0(new_n8806_), .Y(new_n8807_));
  AOI21X1  g08743(.A0(new_n8215_), .A1(new_n2062_), .B0(new_n8807_), .Y(new_n8808_));
  XOR2X1   g08744(.A(new_n8808_), .B(\a[29] ), .Y(new_n8809_));
  INVX1    g08745(.A(new_n8809_), .Y(new_n8810_));
  AOI21X1  g08746(.A0(new_n8810_), .A1(new_n8805_), .B0(new_n8804_), .Y(new_n8811_));
  INVX1    g08747(.A(new_n8811_), .Y(new_n8812_));
  XOR2X1   g08748(.A(new_n8387_), .B(new_n8382_), .Y(new_n8813_));
  XOR2X1   g08749(.A(new_n8813_), .B(new_n8811_), .Y(new_n8814_));
  AOI22X1  g08750(.A0(new_n6892_), .A1(new_n2424_), .B0(new_n6890_), .B1(new_n2418_), .Y(new_n8815_));
  OAI21X1  g08751(.A0(new_n7878_), .A1(new_n2626_), .B0(new_n8815_), .Y(new_n8816_));
  AOI21X1  g08752(.A0(new_n7877_), .A1(new_n2301_), .B0(new_n8816_), .Y(new_n8817_));
  XOR2X1   g08753(.A(new_n8817_), .B(\a[26] ), .Y(new_n8818_));
  NOR2X1   g08754(.A(new_n8818_), .B(new_n8814_), .Y(new_n8819_));
  AOI21X1  g08755(.A0(new_n8813_), .A1(new_n8812_), .B0(new_n8819_), .Y(new_n8820_));
  NOR2X1   g08756(.A(new_n8820_), .B(new_n8533_), .Y(new_n8821_));
  XOR2X1   g08757(.A(new_n8820_), .B(new_n8533_), .Y(new_n8822_));
  AOI22X1  g08758(.A0(new_n6882_), .A1(new_n2657_), .B0(new_n6822_), .B1(new_n2696_), .Y(new_n8823_));
  OAI21X1  g08759(.A0(new_n7671_), .A1(new_n2753_), .B0(new_n8823_), .Y(new_n8824_));
  AOI21X1  g08760(.A0(new_n7670_), .A1(new_n2658_), .B0(new_n8824_), .Y(new_n8825_));
  XOR2X1   g08761(.A(new_n8825_), .B(\a[23] ), .Y(new_n8826_));
  INVX1    g08762(.A(new_n8826_), .Y(new_n8827_));
  AOI21X1  g08763(.A0(new_n8827_), .A1(new_n8822_), .B0(new_n8821_), .Y(new_n8828_));
  NOR2X1   g08764(.A(new_n8828_), .B(new_n8532_), .Y(new_n8829_));
  AOI21X1  g08765(.A0(new_n8530_), .A1(new_n8526_), .B0(new_n8829_), .Y(new_n8830_));
  NOR2X1   g08766(.A(new_n8830_), .B(new_n8525_), .Y(new_n8831_));
  XOR2X1   g08767(.A(new_n8830_), .B(new_n8525_), .Y(new_n8832_));
  AOI22X1  g08768(.A0(new_n7364_), .A1(new_n3099_), .B0(new_n7044_), .B1(new_n2875_), .Y(new_n8833_));
  OAI21X1  g08769(.A0(new_n7504_), .A1(new_n3152_), .B0(new_n8833_), .Y(new_n8834_));
  AOI21X1  g08770(.A0(new_n7552_), .A1(new_n2876_), .B0(new_n8834_), .Y(new_n8835_));
  XOR2X1   g08771(.A(new_n8835_), .B(\a[20] ), .Y(new_n8836_));
  INVX1    g08772(.A(new_n8836_), .Y(new_n8837_));
  AOI21X1  g08773(.A0(new_n8837_), .A1(new_n8832_), .B0(new_n8831_), .Y(new_n8838_));
  NOR2X1   g08774(.A(new_n8838_), .B(new_n8524_), .Y(new_n8839_));
  XOR2X1   g08775(.A(new_n8838_), .B(new_n8524_), .Y(new_n8840_));
  AOI22X1  g08776(.A0(new_n7558_), .A1(new_n3390_), .B0(new_n7529_), .B1(new_n3232_), .Y(new_n8841_));
  OAI21X1  g08777(.A0(new_n7623_), .A1(new_n3545_), .B0(new_n8841_), .Y(new_n8842_));
  AOI21X1  g08778(.A0(new_n7622_), .A1(new_n3234_), .B0(new_n8842_), .Y(new_n8843_));
  XOR2X1   g08779(.A(new_n8843_), .B(\a[17] ), .Y(new_n8844_));
  INVX1    g08780(.A(new_n8844_), .Y(new_n8845_));
  AOI21X1  g08781(.A0(new_n8845_), .A1(new_n8840_), .B0(new_n8839_), .Y(new_n8846_));
  NOR2X1   g08782(.A(new_n8846_), .B(new_n8523_), .Y(new_n8847_));
  AOI21X1  g08783(.A0(new_n8522_), .A1(new_n8517_), .B0(new_n8847_), .Y(new_n8848_));
  NOR2X1   g08784(.A(new_n8848_), .B(new_n8516_), .Y(new_n8849_));
  XOR2X1   g08785(.A(new_n8848_), .B(new_n8516_), .Y(new_n8850_));
  AOI22X1  g08786(.A0(new_n7657_), .A1(new_n3628_), .B0(new_n7341_), .B1(new_n3984_), .Y(new_n8851_));
  OAI21X1  g08787(.A0(new_n7644_), .A1(new_n3907_), .B0(new_n8851_), .Y(new_n8852_));
  AOI21X1  g08788(.A0(new_n7656_), .A1(new_n3624_), .B0(new_n8852_), .Y(new_n8853_));
  XOR2X1   g08789(.A(new_n8853_), .B(\a[14] ), .Y(new_n8854_));
  INVX1    g08790(.A(new_n8854_), .Y(new_n8855_));
  AOI21X1  g08791(.A0(new_n8855_), .A1(new_n8850_), .B0(new_n8849_), .Y(new_n8856_));
  NOR2X1   g08792(.A(new_n8856_), .B(new_n8515_), .Y(new_n8857_));
  INVX1    g08793(.A(new_n8857_), .Y(new_n8858_));
  XOR2X1   g08794(.A(new_n8856_), .B(new_n8515_), .Y(new_n8859_));
  INVX1    g08795(.A(new_n8859_), .Y(new_n8860_));
  XOR2X1   g08796(.A(new_n8854_), .B(new_n8850_), .Y(new_n8861_));
  XOR2X1   g08797(.A(new_n8844_), .B(new_n8840_), .Y(new_n8862_));
  XOR2X1   g08798(.A(new_n8836_), .B(new_n8832_), .Y(new_n8863_));
  XOR2X1   g08799(.A(new_n8828_), .B(new_n8532_), .Y(new_n8864_));
  AOI22X1  g08800(.A0(new_n7044_), .A1(new_n3099_), .B0(new_n6818_), .B1(new_n2875_), .Y(new_n8865_));
  OAI21X1  g08801(.A0(new_n7367_), .A1(new_n3152_), .B0(new_n8865_), .Y(new_n8866_));
  AOI21X1  g08802(.A0(new_n7366_), .A1(new_n2876_), .B0(new_n8866_), .Y(new_n8867_));
  XOR2X1   g08803(.A(new_n8867_), .B(new_n1920_), .Y(new_n8868_));
  XOR2X1   g08804(.A(new_n8867_), .B(\a[20] ), .Y(new_n8869_));
  XOR2X1   g08805(.A(new_n8869_), .B(new_n8864_), .Y(new_n8870_));
  XOR2X1   g08806(.A(new_n8826_), .B(new_n8822_), .Y(new_n8871_));
  INVX1    g08807(.A(new_n8818_), .Y(new_n8872_));
  XOR2X1   g08808(.A(new_n8872_), .B(new_n8814_), .Y(new_n8873_));
  XOR2X1   g08809(.A(new_n8809_), .B(new_n8805_), .Y(new_n8874_));
  AOI22X1  g08810(.A0(new_n6894_), .A1(new_n2424_), .B0(new_n6892_), .B1(new_n2418_), .Y(new_n8875_));
  OAI21X1  g08811(.A0(new_n7885_), .A1(new_n2626_), .B0(new_n8875_), .Y(new_n8876_));
  AOI21X1  g08812(.A0(new_n7884_), .A1(new_n2301_), .B0(new_n8876_), .Y(new_n8877_));
  XOR2X1   g08813(.A(new_n8877_), .B(\a[26] ), .Y(new_n8878_));
  NOR2X1   g08814(.A(new_n8878_), .B(new_n8874_), .Y(new_n8879_));
  XOR2X1   g08815(.A(new_n8878_), .B(new_n8874_), .Y(new_n8880_));
  XOR2X1   g08816(.A(new_n8544_), .B(new_n8536_), .Y(new_n8881_));
  XOR2X1   g08817(.A(new_n8801_), .B(new_n8881_), .Y(new_n8882_));
  INVX1    g08818(.A(new_n8293_), .Y(new_n8883_));
  AOI22X1  g08819(.A0(new_n6904_), .A1(new_n2185_), .B0(new_n6902_), .B1(new_n2095_), .Y(new_n8884_));
  OAI21X1  g08820(.A0(new_n8295_), .A1(new_n2140_), .B0(new_n8884_), .Y(new_n8885_));
  AOI21X1  g08821(.A0(new_n8883_), .A1(new_n2062_), .B0(new_n8885_), .Y(new_n8886_));
  XOR2X1   g08822(.A(new_n8886_), .B(\a[29] ), .Y(new_n8887_));
  OR2X1    g08823(.A(new_n8887_), .B(new_n8882_), .Y(new_n8888_));
  XOR2X1   g08824(.A(new_n8801_), .B(new_n8547_), .Y(new_n8889_));
  XOR2X1   g08825(.A(new_n8887_), .B(new_n8889_), .Y(new_n8890_));
  AOI22X1  g08826(.A0(new_n6897_), .A1(new_n2424_), .B0(new_n6894_), .B1(new_n2418_), .Y(new_n8891_));
  OAI21X1  g08827(.A0(new_n8075_), .A1(new_n2626_), .B0(new_n8891_), .Y(new_n8892_));
  AOI21X1  g08828(.A0(new_n8074_), .A1(new_n2301_), .B0(new_n8892_), .Y(new_n8893_));
  XOR2X1   g08829(.A(new_n8893_), .B(\a[26] ), .Y(new_n8894_));
  OAI21X1  g08830(.A0(new_n8894_), .A1(new_n8890_), .B0(new_n8888_), .Y(new_n8895_));
  AOI21X1  g08831(.A0(new_n8895_), .A1(new_n8880_), .B0(new_n8879_), .Y(new_n8896_));
  NOR2X1   g08832(.A(new_n8896_), .B(new_n8873_), .Y(new_n8897_));
  XOR2X1   g08833(.A(new_n8896_), .B(new_n8873_), .Y(new_n8898_));
  AOI22X1  g08834(.A0(new_n6885_), .A1(new_n2657_), .B0(new_n6882_), .B1(new_n2696_), .Y(new_n8899_));
  OAI21X1  g08835(.A0(new_n7472_), .A1(new_n2753_), .B0(new_n8899_), .Y(new_n8900_));
  AOI21X1  g08836(.A0(new_n7471_), .A1(new_n2658_), .B0(new_n8900_), .Y(new_n8901_));
  XOR2X1   g08837(.A(new_n8901_), .B(\a[23] ), .Y(new_n8902_));
  INVX1    g08838(.A(new_n8902_), .Y(new_n8903_));
  AOI21X1  g08839(.A0(new_n8903_), .A1(new_n8898_), .B0(new_n8897_), .Y(new_n8904_));
  NOR2X1   g08840(.A(new_n8904_), .B(new_n8871_), .Y(new_n8905_));
  XOR2X1   g08841(.A(new_n8904_), .B(new_n8871_), .Y(new_n8906_));
  AOI22X1  g08842(.A0(new_n6818_), .A1(new_n3099_), .B0(new_n6745_), .B1(new_n2875_), .Y(new_n8907_));
  OAI21X1  g08843(.A0(new_n7047_), .A1(new_n3152_), .B0(new_n8907_), .Y(new_n8908_));
  AOI21X1  g08844(.A0(new_n7046_), .A1(new_n2876_), .B0(new_n8908_), .Y(new_n8909_));
  XOR2X1   g08845(.A(new_n8909_), .B(\a[20] ), .Y(new_n8910_));
  INVX1    g08846(.A(new_n8910_), .Y(new_n8911_));
  AOI21X1  g08847(.A0(new_n8911_), .A1(new_n8906_), .B0(new_n8905_), .Y(new_n8912_));
  NOR2X1   g08848(.A(new_n8912_), .B(new_n8870_), .Y(new_n8913_));
  AOI21X1  g08849(.A0(new_n8868_), .A1(new_n8864_), .B0(new_n8913_), .Y(new_n8914_));
  NOR2X1   g08850(.A(new_n8914_), .B(new_n8863_), .Y(new_n8915_));
  XOR2X1   g08851(.A(new_n8914_), .B(new_n8863_), .Y(new_n8916_));
  AOI22X1  g08852(.A0(new_n7529_), .A1(new_n3390_), .B0(new_n7522_), .B1(new_n3232_), .Y(new_n8917_));
  OAI21X1  g08853(.A0(new_n7581_), .A1(new_n3545_), .B0(new_n8917_), .Y(new_n8918_));
  AOI21X1  g08854(.A0(new_n7565_), .A1(new_n3234_), .B0(new_n8918_), .Y(new_n8919_));
  XOR2X1   g08855(.A(new_n8919_), .B(\a[17] ), .Y(new_n8920_));
  INVX1    g08856(.A(new_n8920_), .Y(new_n8921_));
  AOI21X1  g08857(.A0(new_n8921_), .A1(new_n8916_), .B0(new_n8915_), .Y(new_n8922_));
  NOR2X1   g08858(.A(new_n8922_), .B(new_n8862_), .Y(new_n8923_));
  INVX1    g08859(.A(new_n8923_), .Y(new_n8924_));
  XOR2X1   g08860(.A(new_n8922_), .B(new_n8862_), .Y(new_n8925_));
  INVX1    g08861(.A(new_n8925_), .Y(new_n8926_));
  AOI22X1  g08862(.A0(new_n7590_), .A1(new_n3908_), .B0(new_n7578_), .B1(new_n3628_), .Y(new_n8927_));
  OAI21X1  g08863(.A0(new_n7642_), .A1(new_n3983_), .B0(new_n8927_), .Y(new_n8928_));
  AOI21X1  g08864(.A0(new_n7712_), .A1(new_n3624_), .B0(new_n8928_), .Y(new_n8929_));
  XOR2X1   g08865(.A(new_n8929_), .B(\a[14] ), .Y(new_n8930_));
  OR2X1    g08866(.A(new_n8930_), .B(new_n8926_), .Y(new_n8931_));
  AOI22X1  g08867(.A0(new_n7643_), .A1(new_n3984_), .B0(new_n7590_), .B1(new_n3628_), .Y(new_n8932_));
  OAI21X1  g08868(.A0(new_n7642_), .A1(new_n3907_), .B0(new_n8932_), .Y(new_n8933_));
  AOI21X1  g08869(.A0(new_n7718_), .A1(new_n3624_), .B0(new_n8933_), .Y(new_n8934_));
  XOR2X1   g08870(.A(new_n8934_), .B(\a[14] ), .Y(new_n8935_));
  AOI21X1  g08871(.A0(new_n8931_), .A1(new_n8924_), .B0(new_n8935_), .Y(new_n8936_));
  INVX1    g08872(.A(new_n8523_), .Y(new_n8937_));
  XOR2X1   g08873(.A(new_n8846_), .B(new_n8937_), .Y(new_n8938_));
  OAI21X1  g08874(.A0(new_n8930_), .A1(new_n8926_), .B0(new_n8924_), .Y(new_n8939_));
  XOR2X1   g08875(.A(new_n8935_), .B(new_n8939_), .Y(new_n8940_));
  NOR2X1   g08876(.A(new_n8940_), .B(new_n8938_), .Y(new_n8941_));
  NOR2X1   g08877(.A(new_n8941_), .B(new_n8936_), .Y(new_n8942_));
  NOR2X1   g08878(.A(new_n8942_), .B(new_n8861_), .Y(new_n8943_));
  XOR2X1   g08879(.A(new_n8942_), .B(new_n8861_), .Y(new_n8944_));
  XOR2X1   g08880(.A(new_n8920_), .B(new_n8916_), .Y(new_n8945_));
  XOR2X1   g08881(.A(new_n8912_), .B(new_n8870_), .Y(new_n8946_));
  AOI22X1  g08882(.A0(new_n7522_), .A1(new_n3390_), .B0(new_n7485_), .B1(new_n3232_), .Y(new_n8947_));
  OAI21X1  g08883(.A0(new_n7537_), .A1(new_n3545_), .B0(new_n8947_), .Y(new_n8948_));
  AOI21X1  g08884(.A0(new_n7536_), .A1(new_n3234_), .B0(new_n8948_), .Y(new_n8949_));
  XOR2X1   g08885(.A(new_n8949_), .B(new_n2445_), .Y(new_n8950_));
  XOR2X1   g08886(.A(new_n8949_), .B(\a[17] ), .Y(new_n8951_));
  XOR2X1   g08887(.A(new_n8951_), .B(new_n8946_), .Y(new_n8952_));
  XOR2X1   g08888(.A(new_n8910_), .B(new_n8906_), .Y(new_n8953_));
  XOR2X1   g08889(.A(new_n8902_), .B(new_n8898_), .Y(new_n8954_));
  OR2X1    g08890(.A(new_n8894_), .B(new_n8890_), .Y(new_n8955_));
  AND2X1   g08891(.A(new_n8955_), .B(new_n8888_), .Y(new_n8956_));
  XOR2X1   g08892(.A(new_n8956_), .B(new_n8880_), .Y(new_n8957_));
  AOI22X1  g08893(.A0(new_n6887_), .A1(new_n2657_), .B0(new_n6885_), .B1(new_n2696_), .Y(new_n8958_));
  OAI21X1  g08894(.A0(new_n6884_), .A1(new_n2753_), .B0(new_n8958_), .Y(new_n8959_));
  AOI21X1  g08895(.A0(new_n7771_), .A1(new_n2658_), .B0(new_n8959_), .Y(new_n8960_));
  XOR2X1   g08896(.A(new_n8960_), .B(\a[23] ), .Y(new_n8961_));
  NOR2X1   g08897(.A(new_n8961_), .B(new_n8957_), .Y(new_n8962_));
  XOR2X1   g08898(.A(new_n8961_), .B(new_n8957_), .Y(new_n8963_));
  XOR2X1   g08899(.A(new_n8887_), .B(new_n8882_), .Y(new_n8964_));
  XOR2X1   g08900(.A(new_n8894_), .B(new_n8964_), .Y(new_n8965_));
  AOI21X1  g08901(.A0(new_n8560_), .A1(new_n8559_), .B0(new_n8557_), .Y(new_n8966_));
  NOR3X1   g08902(.A(new_n8556_), .B(new_n8551_), .C(new_n8550_), .Y(new_n8967_));
  AOI21X1  g08903(.A0(new_n8371_), .A1(new_n8344_), .B0(new_n8352_), .Y(new_n8968_));
  NOR3X1   g08904(.A(new_n8372_), .B(new_n8345_), .C(new_n8370_), .Y(new_n8969_));
  OAI21X1  g08905(.A0(new_n8969_), .A1(new_n8968_), .B0(new_n8790_), .Y(new_n8970_));
  NOR3X1   g08906(.A(new_n8790_), .B(new_n8969_), .C(new_n8968_), .Y(new_n8971_));
  OAI21X1  g08907(.A0(new_n8797_), .A1(new_n8971_), .B0(new_n8970_), .Y(new_n8972_));
  OAI21X1  g08908(.A0(new_n8967_), .A1(new_n8966_), .B0(new_n8972_), .Y(new_n8973_));
  NAND3X1  g08909(.A(new_n8799_), .B(new_n8561_), .C(new_n8558_), .Y(new_n8974_));
  AOI22X1  g08910(.A0(new_n6906_), .A1(new_n2185_), .B0(new_n6904_), .B1(new_n2095_), .Y(new_n8975_));
  OAI21X1  g08911(.A0(new_n8205_), .A1(new_n2140_), .B0(new_n8975_), .Y(new_n8976_));
  AOI21X1  g08912(.A0(new_n8204_), .A1(new_n2062_), .B0(new_n8976_), .Y(new_n8977_));
  XOR2X1   g08913(.A(new_n8977_), .B(\a[29] ), .Y(new_n8978_));
  INVX1    g08914(.A(new_n8978_), .Y(new_n8979_));
  NAND3X1  g08915(.A(new_n8979_), .B(new_n8974_), .C(new_n8973_), .Y(new_n8980_));
  NOR3X1   g08916(.A(new_n8972_), .B(new_n8967_), .C(new_n8966_), .Y(new_n8981_));
  NOR3X1   g08917(.A(new_n8979_), .B(new_n8981_), .C(new_n8800_), .Y(new_n8982_));
  AOI21X1  g08918(.A0(new_n8974_), .A1(new_n8973_), .B0(new_n8978_), .Y(new_n8983_));
  AOI22X1  g08919(.A0(new_n6899_), .A1(new_n2424_), .B0(new_n6897_), .B1(new_n2418_), .Y(new_n8984_));
  OAI21X1  g08920(.A0(new_n6896_), .A1(new_n2626_), .B0(new_n8984_), .Y(new_n8985_));
  AOI21X1  g08921(.A0(new_n7953_), .A1(new_n2301_), .B0(new_n8985_), .Y(new_n8986_));
  XOR2X1   g08922(.A(new_n8986_), .B(\a[26] ), .Y(new_n8987_));
  INVX1    g08923(.A(new_n8987_), .Y(new_n8988_));
  OAI21X1  g08924(.A0(new_n8983_), .A1(new_n8982_), .B0(new_n8988_), .Y(new_n8989_));
  AND2X1   g08925(.A(new_n8989_), .B(new_n8980_), .Y(new_n8990_));
  OR2X1    g08926(.A(new_n8990_), .B(new_n8965_), .Y(new_n8991_));
  XOR2X1   g08927(.A(new_n8894_), .B(new_n8890_), .Y(new_n8992_));
  XOR2X1   g08928(.A(new_n8990_), .B(new_n8992_), .Y(new_n8993_));
  AOI22X1  g08929(.A0(new_n6890_), .A1(new_n2657_), .B0(new_n6887_), .B1(new_n2696_), .Y(new_n8994_));
  OAI21X1  g08930(.A0(new_n6886_), .A1(new_n2753_), .B0(new_n8994_), .Y(new_n8995_));
  AOI21X1  g08931(.A0(new_n7762_), .A1(new_n2658_), .B0(new_n8995_), .Y(new_n8996_));
  XOR2X1   g08932(.A(new_n8996_), .B(\a[23] ), .Y(new_n8997_));
  OAI21X1  g08933(.A0(new_n8997_), .A1(new_n8993_), .B0(new_n8991_), .Y(new_n8998_));
  AOI21X1  g08934(.A0(new_n8998_), .A1(new_n8963_), .B0(new_n8962_), .Y(new_n8999_));
  NOR2X1   g08935(.A(new_n8999_), .B(new_n8954_), .Y(new_n9000_));
  XOR2X1   g08936(.A(new_n8999_), .B(new_n8954_), .Y(new_n9001_));
  AOI22X1  g08937(.A0(new_n6820_), .A1(new_n2875_), .B0(new_n6745_), .B1(new_n3099_), .Y(new_n9002_));
  OAI21X1  g08938(.A0(new_n7361_), .A1(new_n3152_), .B0(new_n9002_), .Y(new_n9003_));
  AOI21X1  g08939(.A0(new_n7404_), .A1(new_n2876_), .B0(new_n9003_), .Y(new_n9004_));
  XOR2X1   g08940(.A(new_n9004_), .B(\a[20] ), .Y(new_n9005_));
  INVX1    g08941(.A(new_n9005_), .Y(new_n9006_));
  AOI21X1  g08942(.A0(new_n9006_), .A1(new_n9001_), .B0(new_n9000_), .Y(new_n9007_));
  NOR2X1   g08943(.A(new_n9007_), .B(new_n8953_), .Y(new_n9008_));
  XOR2X1   g08944(.A(new_n9007_), .B(new_n8953_), .Y(new_n9009_));
  AOI22X1  g08945(.A0(new_n7485_), .A1(new_n3390_), .B0(new_n7364_), .B1(new_n3232_), .Y(new_n9010_));
  OAI21X1  g08946(.A0(new_n7523_), .A1(new_n3545_), .B0(new_n9010_), .Y(new_n9011_));
  AOI21X1  g08947(.A0(new_n7612_), .A1(new_n3234_), .B0(new_n9011_), .Y(new_n9012_));
  XOR2X1   g08948(.A(new_n9012_), .B(\a[17] ), .Y(new_n9013_));
  INVX1    g08949(.A(new_n9013_), .Y(new_n9014_));
  AOI21X1  g08950(.A0(new_n9014_), .A1(new_n9009_), .B0(new_n9008_), .Y(new_n9015_));
  NOR2X1   g08951(.A(new_n9015_), .B(new_n8952_), .Y(new_n9016_));
  AOI21X1  g08952(.A0(new_n8950_), .A1(new_n8946_), .B0(new_n9016_), .Y(new_n9017_));
  NOR2X1   g08953(.A(new_n9017_), .B(new_n8945_), .Y(new_n9018_));
  XOR2X1   g08954(.A(new_n9017_), .B(new_n8945_), .Y(new_n9019_));
  AOI22X1  g08955(.A0(new_n7578_), .A1(new_n3908_), .B0(new_n7571_), .B1(new_n3628_), .Y(new_n9020_));
  OAI21X1  g08956(.A0(new_n7594_), .A1(new_n3983_), .B0(new_n9020_), .Y(new_n9021_));
  AOI21X1  g08957(.A0(new_n7593_), .A1(new_n3624_), .B0(new_n9021_), .Y(new_n9022_));
  XOR2X1   g08958(.A(new_n9022_), .B(\a[14] ), .Y(new_n9023_));
  INVX1    g08959(.A(new_n9023_), .Y(new_n9024_));
  AOI21X1  g08960(.A0(new_n9024_), .A1(new_n9019_), .B0(new_n9018_), .Y(new_n9025_));
  NAND2X1  g08961(.A(new_n4427_), .B(new_n4246_), .Y(new_n9026_));
  AOI22X1  g08962(.A0(new_n9026_), .A1(new_n7341_), .B0(new_n7643_), .B1(new_n4078_), .Y(new_n9027_));
  OAI21X1  g08963(.A0(new_n7808_), .A1(new_n4245_), .B0(new_n9027_), .Y(new_n9028_));
  XOR2X1   g08964(.A(new_n9028_), .B(new_n2911_), .Y(new_n9029_));
  NOR2X1   g08965(.A(new_n9029_), .B(new_n9025_), .Y(new_n9030_));
  XOR2X1   g08966(.A(new_n8930_), .B(new_n8925_), .Y(new_n9031_));
  INVX1    g08967(.A(new_n9031_), .Y(new_n9032_));
  XOR2X1   g08968(.A(new_n9029_), .B(new_n9025_), .Y(new_n9033_));
  AOI21X1  g08969(.A0(new_n9033_), .A1(new_n9032_), .B0(new_n9030_), .Y(new_n9034_));
  INVX1    g08970(.A(new_n9034_), .Y(new_n9035_));
  XOR2X1   g08971(.A(new_n8940_), .B(new_n8938_), .Y(new_n9036_));
  AND2X1   g08972(.A(new_n9036_), .B(new_n9035_), .Y(new_n9037_));
  INVX1    g08973(.A(new_n9037_), .Y(new_n9038_));
  XOR2X1   g08974(.A(new_n9033_), .B(new_n9031_), .Y(new_n9039_));
  XOR2X1   g08975(.A(new_n9023_), .B(new_n9019_), .Y(new_n9040_));
  XOR2X1   g08976(.A(new_n9015_), .B(new_n8952_), .Y(new_n9041_));
  INVX1    g08977(.A(new_n9041_), .Y(new_n9042_));
  AOI22X1  g08978(.A0(new_n7571_), .A1(new_n3908_), .B0(new_n7558_), .B1(new_n3628_), .Y(new_n9043_));
  OAI21X1  g08979(.A0(new_n7602_), .A1(new_n3983_), .B0(new_n9043_), .Y(new_n9044_));
  AOI21X1  g08980(.A0(new_n7601_), .A1(new_n3624_), .B0(new_n9044_), .Y(new_n9045_));
  XOR2X1   g08981(.A(new_n9045_), .B(\a[14] ), .Y(new_n9046_));
  NOR2X1   g08982(.A(new_n9046_), .B(new_n9042_), .Y(new_n9047_));
  XOR2X1   g08983(.A(new_n9046_), .B(new_n9041_), .Y(new_n9048_));
  INVX1    g08984(.A(new_n9048_), .Y(new_n9049_));
  XOR2X1   g08985(.A(new_n9013_), .B(new_n9009_), .Y(new_n9050_));
  XOR2X1   g08986(.A(new_n9005_), .B(new_n9001_), .Y(new_n9051_));
  OR2X1    g08987(.A(new_n8997_), .B(new_n8993_), .Y(new_n9052_));
  AND2X1   g08988(.A(new_n9052_), .B(new_n8991_), .Y(new_n9053_));
  XOR2X1   g08989(.A(new_n9053_), .B(new_n8963_), .Y(new_n9054_));
  AOI22X1  g08990(.A0(new_n6822_), .A1(new_n2875_), .B0(new_n6820_), .B1(new_n3099_), .Y(new_n9055_));
  OAI21X1  g08991(.A0(new_n7418_), .A1(new_n3152_), .B0(new_n9055_), .Y(new_n9056_));
  AOI21X1  g08992(.A0(new_n7417_), .A1(new_n2876_), .B0(new_n9056_), .Y(new_n9057_));
  XOR2X1   g08993(.A(new_n9057_), .B(\a[20] ), .Y(new_n9058_));
  NOR2X1   g08994(.A(new_n9058_), .B(new_n9054_), .Y(new_n9059_));
  XOR2X1   g08995(.A(new_n9058_), .B(new_n9054_), .Y(new_n9060_));
  XOR2X1   g08996(.A(new_n8990_), .B(new_n8965_), .Y(new_n9061_));
  XOR2X1   g08997(.A(new_n8997_), .B(new_n9061_), .Y(new_n9062_));
  OAI21X1  g08998(.A0(new_n8983_), .A1(new_n8982_), .B0(new_n8987_), .Y(new_n9063_));
  NAND3X1  g08999(.A(new_n8978_), .B(new_n8974_), .C(new_n8973_), .Y(new_n9064_));
  OAI21X1  g09000(.A0(new_n8981_), .A1(new_n8800_), .B0(new_n8979_), .Y(new_n9065_));
  NAND3X1  g09001(.A(new_n8988_), .B(new_n9065_), .C(new_n9064_), .Y(new_n9066_));
  NOR3X1   g09002(.A(new_n8797_), .B(new_n8971_), .C(new_n8792_), .Y(new_n9067_));
  XOR2X1   g09003(.A(new_n8789_), .B(new_n8787_), .Y(new_n9068_));
  AOI22X1  g09004(.A0(new_n6911_), .A1(new_n2185_), .B0(new_n6909_), .B1(new_n2095_), .Y(new_n9069_));
  OAI21X1  g09005(.A0(new_n6964_), .A1(new_n2140_), .B0(new_n9069_), .Y(new_n9070_));
  AOI21X1  g09006(.A0(new_n8541_), .A1(new_n2062_), .B0(new_n9070_), .Y(new_n9071_));
  XOR2X1   g09007(.A(new_n9071_), .B(\a[29] ), .Y(new_n9072_));
  NOR2X1   g09008(.A(new_n9072_), .B(new_n9068_), .Y(new_n9073_));
  XOR2X1   g09009(.A(new_n8786_), .B(new_n8783_), .Y(new_n9074_));
  INVX1    g09010(.A(new_n8553_), .Y(new_n9075_));
  OAI22X1  g09011(.A0(new_n8579_), .A1(new_n2186_), .B0(new_n8349_), .B1(new_n2431_), .Y(new_n9076_));
  AOI21X1  g09012(.A0(new_n6909_), .A1(new_n2139_), .B0(new_n9076_), .Y(new_n9077_));
  OAI21X1  g09013(.A0(new_n9075_), .A1(new_n2063_), .B0(new_n9077_), .Y(new_n9078_));
  XOR2X1   g09014(.A(new_n9078_), .B(new_n74_), .Y(new_n9079_));
  NOR2X1   g09015(.A(new_n9079_), .B(new_n9074_), .Y(new_n9080_));
  XOR2X1   g09016(.A(new_n8782_), .B(new_n8780_), .Y(new_n9081_));
  INVX1    g09017(.A(new_n8348_), .Y(new_n9082_));
  OAI22X1  g09018(.A0(new_n6917_), .A1(new_n2186_), .B0(new_n8579_), .B1(new_n2431_), .Y(new_n9083_));
  AOI21X1  g09019(.A0(new_n6911_), .A1(new_n2139_), .B0(new_n9083_), .Y(new_n9084_));
  OAI21X1  g09020(.A0(new_n9082_), .A1(new_n2063_), .B0(new_n9084_), .Y(new_n9085_));
  XOR2X1   g09021(.A(new_n9085_), .B(new_n74_), .Y(new_n9086_));
  XOR2X1   g09022(.A(new_n8779_), .B(new_n8777_), .Y(new_n9087_));
  OAI22X1  g09023(.A0(new_n6918_), .A1(new_n2186_), .B0(new_n6917_), .B1(new_n2431_), .Y(new_n9088_));
  AOI21X1  g09024(.A0(new_n6913_), .A1(new_n2139_), .B0(new_n9088_), .Y(new_n9089_));
  OAI21X1  g09025(.A0(new_n8577_), .A1(new_n2063_), .B0(new_n9089_), .Y(new_n9090_));
  XOR2X1   g09026(.A(new_n9090_), .B(new_n74_), .Y(new_n9091_));
  XOR2X1   g09027(.A(new_n8776_), .B(new_n8774_), .Y(new_n9092_));
  NOR2X1   g09028(.A(new_n8595_), .B(new_n8594_), .Y(new_n9093_));
  OAI22X1  g09029(.A0(new_n6920_), .A1(new_n2186_), .B0(new_n6918_), .B1(new_n2431_), .Y(new_n9094_));
  AOI21X1  g09030(.A0(new_n6915_), .A1(new_n2139_), .B0(new_n9094_), .Y(new_n9095_));
  OAI21X1  g09031(.A0(new_n9093_), .A1(new_n2063_), .B0(new_n9095_), .Y(new_n9096_));
  XOR2X1   g09032(.A(new_n9096_), .B(new_n74_), .Y(new_n9097_));
  AOI22X1  g09033(.A0(new_n6923_), .A1(new_n2185_), .B0(new_n6922_), .B1(new_n2095_), .Y(new_n9098_));
  OAI21X1  g09034(.A0(new_n6918_), .A1(new_n2140_), .B0(new_n9098_), .Y(new_n9099_));
  AOI21X1  g09035(.A0(new_n8612_), .A1(new_n2062_), .B0(new_n9099_), .Y(new_n9100_));
  XOR2X1   g09036(.A(new_n9100_), .B(\a[29] ), .Y(new_n9101_));
  XOR2X1   g09037(.A(new_n8772_), .B(new_n8771_), .Y(new_n9102_));
  NOR2X1   g09038(.A(new_n9102_), .B(new_n9101_), .Y(new_n9103_));
  INVX1    g09039(.A(new_n9103_), .Y(new_n9104_));
  INVX1    g09040(.A(new_n9102_), .Y(new_n9105_));
  XOR2X1   g09041(.A(new_n9105_), .B(new_n9101_), .Y(new_n9106_));
  AOI22X1  g09042(.A0(new_n6925_), .A1(new_n2185_), .B0(new_n6923_), .B1(new_n2095_), .Y(new_n9107_));
  OAI21X1  g09043(.A0(new_n6920_), .A1(new_n2140_), .B0(new_n9107_), .Y(new_n9108_));
  AOI21X1  g09044(.A0(new_n8628_), .A1(new_n2062_), .B0(new_n9108_), .Y(new_n9109_));
  XOR2X1   g09045(.A(new_n9109_), .B(\a[29] ), .Y(new_n9110_));
  XOR2X1   g09046(.A(new_n8770_), .B(new_n8768_), .Y(new_n9111_));
  NOR2X1   g09047(.A(new_n9111_), .B(new_n9110_), .Y(new_n9112_));
  XOR2X1   g09048(.A(new_n9111_), .B(new_n9110_), .Y(new_n9113_));
  AOI22X1  g09049(.A0(new_n6927_), .A1(new_n2185_), .B0(new_n6925_), .B1(new_n2095_), .Y(new_n9114_));
  OAI21X1  g09050(.A0(new_n8659_), .A1(new_n2140_), .B0(new_n9114_), .Y(new_n9115_));
  AOI21X1  g09051(.A0(new_n8663_), .A1(new_n2062_), .B0(new_n9115_), .Y(new_n9116_));
  XOR2X1   g09052(.A(new_n9116_), .B(\a[29] ), .Y(new_n9117_));
  XOR2X1   g09053(.A(new_n8720_), .B(new_n8716_), .Y(new_n9118_));
  XOR2X1   g09054(.A(new_n9118_), .B(new_n8764_), .Y(new_n9119_));
  OR2X1    g09055(.A(new_n9119_), .B(new_n9117_), .Y(new_n9120_));
  XOR2X1   g09056(.A(new_n9119_), .B(new_n9117_), .Y(new_n9121_));
  INVX1    g09057(.A(new_n9121_), .Y(new_n9122_));
  AOI22X1  g09058(.A0(new_n6932_), .A1(new_n2185_), .B0(new_n6927_), .B1(new_n2095_), .Y(new_n9123_));
  OAI21X1  g09059(.A0(new_n8683_), .A1(new_n2140_), .B0(new_n9123_), .Y(new_n9124_));
  AOI21X1  g09060(.A0(new_n8682_), .A1(new_n2062_), .B0(new_n9124_), .Y(new_n9125_));
  XOR2X1   g09061(.A(new_n9125_), .B(\a[29] ), .Y(new_n9126_));
  INVX1    g09062(.A(new_n8762_), .Y(new_n9127_));
  XOR2X1   g09063(.A(new_n8763_), .B(new_n9127_), .Y(new_n9128_));
  NOR2X1   g09064(.A(new_n9128_), .B(new_n9126_), .Y(new_n9129_));
  XOR2X1   g09065(.A(new_n9128_), .B(new_n9126_), .Y(new_n9130_));
  AOI22X1  g09066(.A0(new_n6933_), .A1(new_n2185_), .B0(new_n6932_), .B1(new_n2095_), .Y(new_n9131_));
  OAI21X1  g09067(.A0(new_n6929_), .A1(new_n2140_), .B0(new_n9131_), .Y(new_n9132_));
  AOI21X1  g09068(.A0(new_n8706_), .A1(new_n2062_), .B0(new_n9132_), .Y(new_n9133_));
  XOR2X1   g09069(.A(new_n9133_), .B(\a[29] ), .Y(new_n9134_));
  INVX1    g09070(.A(new_n8750_), .Y(new_n9135_));
  XOR2X1   g09071(.A(new_n8754_), .B(new_n9135_), .Y(new_n9136_));
  OR2X1    g09072(.A(new_n9136_), .B(new_n9134_), .Y(new_n9137_));
  XOR2X1   g09073(.A(new_n9136_), .B(new_n9134_), .Y(new_n9138_));
  INVX1    g09074(.A(new_n9138_), .Y(new_n9139_));
  NOR2X1   g09075(.A(new_n6936_), .B(new_n4171_), .Y(new_n9140_));
  OAI22X1  g09076(.A0(new_n6936_), .A1(new_n2431_), .B0(new_n8752_), .B1(new_n2140_), .Y(new_n9141_));
  AOI21X1  g09077(.A0(new_n8751_), .A1(new_n2062_), .B0(new_n9141_), .Y(new_n9142_));
  XOR2X1   g09078(.A(new_n9142_), .B(\a[29] ), .Y(new_n9143_));
  NOR2X1   g09079(.A(new_n6936_), .B(new_n2061_), .Y(new_n9144_));
  OAI22X1  g09080(.A0(new_n6936_), .A1(new_n2186_), .B0(new_n8752_), .B1(new_n2431_), .Y(new_n9145_));
  AOI21X1  g09081(.A0(new_n6933_), .A1(new_n2139_), .B0(new_n9145_), .Y(new_n9146_));
  OAI21X1  g09082(.A0(new_n8759_), .A1(new_n2063_), .B0(new_n9146_), .Y(new_n9147_));
  NOR4X1   g09083(.A(new_n9147_), .B(new_n9144_), .C(new_n9143_), .D(new_n74_), .Y(new_n9148_));
  AOI22X1  g09084(.A0(new_n6935_), .A1(new_n2185_), .B0(new_n6933_), .B1(new_n2095_), .Y(new_n9149_));
  OAI21X1  g09085(.A0(new_n6930_), .A1(new_n2140_), .B0(new_n9149_), .Y(new_n9150_));
  AOI21X1  g09086(.A0(new_n8717_), .A1(new_n2062_), .B0(new_n9150_), .Y(new_n9151_));
  XOR2X1   g09087(.A(new_n9151_), .B(\a[29] ), .Y(new_n9152_));
  INVX1    g09088(.A(new_n9140_), .Y(new_n9153_));
  XOR2X1   g09089(.A(new_n9148_), .B(new_n9153_), .Y(new_n9154_));
  NOR2X1   g09090(.A(new_n9154_), .B(new_n9152_), .Y(new_n9155_));
  AOI21X1  g09091(.A0(new_n9148_), .A1(new_n9140_), .B0(new_n9155_), .Y(new_n9156_));
  OAI21X1  g09092(.A0(new_n9156_), .A1(new_n9139_), .B0(new_n9137_), .Y(new_n9157_));
  AOI21X1  g09093(.A0(new_n9157_), .A1(new_n9130_), .B0(new_n9129_), .Y(new_n9158_));
  OAI21X1  g09094(.A0(new_n9158_), .A1(new_n9122_), .B0(new_n9120_), .Y(new_n9159_));
  AOI21X1  g09095(.A0(new_n9159_), .A1(new_n9113_), .B0(new_n9112_), .Y(new_n9160_));
  OAI21X1  g09096(.A0(new_n9160_), .A1(new_n9106_), .B0(new_n9104_), .Y(new_n9161_));
  XOR2X1   g09097(.A(new_n9097_), .B(new_n9092_), .Y(new_n9162_));
  NAND2X1  g09098(.A(new_n9162_), .B(new_n9161_), .Y(new_n9163_));
  OAI21X1  g09099(.A0(new_n9097_), .A1(new_n9092_), .B0(new_n9163_), .Y(new_n9164_));
  XOR2X1   g09100(.A(new_n9091_), .B(new_n9087_), .Y(new_n9165_));
  NAND2X1  g09101(.A(new_n9165_), .B(new_n9164_), .Y(new_n9166_));
  OAI21X1  g09102(.A0(new_n9091_), .A1(new_n9087_), .B0(new_n9166_), .Y(new_n9167_));
  XOR2X1   g09103(.A(new_n9086_), .B(new_n9081_), .Y(new_n9168_));
  NAND2X1  g09104(.A(new_n9168_), .B(new_n9167_), .Y(new_n9169_));
  OAI21X1  g09105(.A0(new_n9086_), .A1(new_n9081_), .B0(new_n9169_), .Y(new_n9170_));
  XOR2X1   g09106(.A(new_n9079_), .B(new_n9074_), .Y(new_n9171_));
  AOI21X1  g09107(.A0(new_n9171_), .A1(new_n9170_), .B0(new_n9080_), .Y(new_n9172_));
  INVX1    g09108(.A(new_n9172_), .Y(new_n9173_));
  XOR2X1   g09109(.A(new_n9072_), .B(new_n9068_), .Y(new_n9174_));
  AOI21X1  g09110(.A0(new_n9174_), .A1(new_n9173_), .B0(new_n9073_), .Y(new_n9175_));
  AOI21X1  g09111(.A0(new_n8793_), .A1(new_n8970_), .B0(new_n8798_), .Y(new_n9176_));
  NOR3X1   g09112(.A(new_n9176_), .B(new_n9175_), .C(new_n9067_), .Y(new_n9177_));
  OAI21X1  g09113(.A0(new_n9176_), .A1(new_n9067_), .B0(new_n9175_), .Y(new_n9178_));
  AOI22X1  g09114(.A0(new_n6902_), .A1(new_n2424_), .B0(new_n6899_), .B1(new_n2418_), .Y(new_n9179_));
  OAI21X1  g09115(.A0(new_n6898_), .A1(new_n2626_), .B0(new_n9179_), .Y(new_n9180_));
  AOI21X1  g09116(.A0(new_n8215_), .A1(new_n2301_), .B0(new_n9180_), .Y(new_n9181_));
  XOR2X1   g09117(.A(new_n9181_), .B(\a[26] ), .Y(new_n9182_));
  INVX1    g09118(.A(new_n9182_), .Y(new_n9183_));
  AOI21X1  g09119(.A0(new_n9183_), .A1(new_n9178_), .B0(new_n9177_), .Y(new_n9184_));
  AOI21X1  g09120(.A0(new_n9066_), .A1(new_n9063_), .B0(new_n9184_), .Y(new_n9185_));
  NAND3X1  g09121(.A(new_n9184_), .B(new_n9066_), .C(new_n9063_), .Y(new_n9186_));
  AOI22X1  g09122(.A0(new_n6892_), .A1(new_n2657_), .B0(new_n6890_), .B1(new_n2696_), .Y(new_n9187_));
  OAI21X1  g09123(.A0(new_n7878_), .A1(new_n2753_), .B0(new_n9187_), .Y(new_n9188_));
  AOI21X1  g09124(.A0(new_n7877_), .A1(new_n2658_), .B0(new_n9188_), .Y(new_n9189_));
  XOR2X1   g09125(.A(new_n9189_), .B(\a[23] ), .Y(new_n9190_));
  INVX1    g09126(.A(new_n9190_), .Y(new_n9191_));
  AOI21X1  g09127(.A0(new_n9191_), .A1(new_n9186_), .B0(new_n9185_), .Y(new_n9192_));
  OR2X1    g09128(.A(new_n9192_), .B(new_n9062_), .Y(new_n9193_));
  XOR2X1   g09129(.A(new_n8997_), .B(new_n8993_), .Y(new_n9194_));
  XOR2X1   g09130(.A(new_n9192_), .B(new_n9194_), .Y(new_n9195_));
  AOI22X1  g09131(.A0(new_n6882_), .A1(new_n2875_), .B0(new_n6822_), .B1(new_n3099_), .Y(new_n9196_));
  OAI21X1  g09132(.A0(new_n7671_), .A1(new_n3152_), .B0(new_n9196_), .Y(new_n9197_));
  AOI21X1  g09133(.A0(new_n7670_), .A1(new_n2876_), .B0(new_n9197_), .Y(new_n9198_));
  XOR2X1   g09134(.A(new_n9198_), .B(\a[20] ), .Y(new_n9199_));
  OAI21X1  g09135(.A0(new_n9199_), .A1(new_n9195_), .B0(new_n9193_), .Y(new_n9200_));
  AOI21X1  g09136(.A0(new_n9200_), .A1(new_n9060_), .B0(new_n9059_), .Y(new_n9201_));
  NOR2X1   g09137(.A(new_n9201_), .B(new_n9051_), .Y(new_n9202_));
  XOR2X1   g09138(.A(new_n9201_), .B(new_n9051_), .Y(new_n9203_));
  AOI22X1  g09139(.A0(new_n7364_), .A1(new_n3390_), .B0(new_n7044_), .B1(new_n3232_), .Y(new_n9204_));
  OAI21X1  g09140(.A0(new_n7504_), .A1(new_n3545_), .B0(new_n9204_), .Y(new_n9205_));
  AOI21X1  g09141(.A0(new_n7552_), .A1(new_n3234_), .B0(new_n9205_), .Y(new_n9206_));
  XOR2X1   g09142(.A(new_n9206_), .B(\a[17] ), .Y(new_n9207_));
  INVX1    g09143(.A(new_n9207_), .Y(new_n9208_));
  AOI21X1  g09144(.A0(new_n9208_), .A1(new_n9203_), .B0(new_n9202_), .Y(new_n9209_));
  OR2X1    g09145(.A(new_n9209_), .B(new_n9050_), .Y(new_n9210_));
  XOR2X1   g09146(.A(new_n9014_), .B(new_n9009_), .Y(new_n9211_));
  XOR2X1   g09147(.A(new_n9209_), .B(new_n9211_), .Y(new_n9212_));
  AOI22X1  g09148(.A0(new_n7558_), .A1(new_n3908_), .B0(new_n7529_), .B1(new_n3628_), .Y(new_n9213_));
  OAI21X1  g09149(.A0(new_n7623_), .A1(new_n3983_), .B0(new_n9213_), .Y(new_n9214_));
  AOI21X1  g09150(.A0(new_n7622_), .A1(new_n3624_), .B0(new_n9214_), .Y(new_n9215_));
  XOR2X1   g09151(.A(new_n9215_), .B(\a[14] ), .Y(new_n9216_));
  OAI21X1  g09152(.A0(new_n9216_), .A1(new_n9212_), .B0(new_n9210_), .Y(new_n9217_));
  AOI21X1  g09153(.A0(new_n9217_), .A1(new_n9049_), .B0(new_n9047_), .Y(new_n9218_));
  NOR2X1   g09154(.A(new_n9218_), .B(new_n9040_), .Y(new_n9219_));
  XOR2X1   g09155(.A(new_n9218_), .B(new_n9040_), .Y(new_n9220_));
  AOI22X1  g09156(.A0(new_n7657_), .A1(new_n4078_), .B0(new_n7341_), .B1(new_n4428_), .Y(new_n9221_));
  OAI21X1  g09157(.A0(new_n7644_), .A1(new_n4246_), .B0(new_n9221_), .Y(new_n9222_));
  AOI21X1  g09158(.A0(new_n7656_), .A1(new_n4080_), .B0(new_n9222_), .Y(new_n9223_));
  XOR2X1   g09159(.A(new_n9223_), .B(\a[11] ), .Y(new_n9224_));
  INVX1    g09160(.A(new_n9224_), .Y(new_n9225_));
  AOI21X1  g09161(.A0(new_n9225_), .A1(new_n9220_), .B0(new_n9219_), .Y(new_n9226_));
  NOR2X1   g09162(.A(new_n9226_), .B(new_n9039_), .Y(new_n9227_));
  XOR2X1   g09163(.A(new_n9226_), .B(new_n9039_), .Y(new_n9228_));
  XOR2X1   g09164(.A(new_n9224_), .B(new_n9220_), .Y(new_n9229_));
  XOR2X1   g09165(.A(new_n9209_), .B(new_n9050_), .Y(new_n9230_));
  XOR2X1   g09166(.A(new_n9216_), .B(new_n9230_), .Y(new_n9231_));
  XOR2X1   g09167(.A(new_n9207_), .B(new_n9203_), .Y(new_n9232_));
  OR2X1    g09168(.A(new_n9199_), .B(new_n9195_), .Y(new_n9233_));
  AND2X1   g09169(.A(new_n9233_), .B(new_n9193_), .Y(new_n9234_));
  XOR2X1   g09170(.A(new_n9234_), .B(new_n9060_), .Y(new_n9235_));
  AOI22X1  g09171(.A0(new_n7044_), .A1(new_n3390_), .B0(new_n6818_), .B1(new_n3232_), .Y(new_n9236_));
  OAI21X1  g09172(.A0(new_n7367_), .A1(new_n3545_), .B0(new_n9236_), .Y(new_n9237_));
  AOI21X1  g09173(.A0(new_n7366_), .A1(new_n3234_), .B0(new_n9237_), .Y(new_n9238_));
  XOR2X1   g09174(.A(new_n9238_), .B(\a[17] ), .Y(new_n9239_));
  NOR2X1   g09175(.A(new_n9239_), .B(new_n9235_), .Y(new_n9240_));
  XOR2X1   g09176(.A(new_n9239_), .B(new_n9235_), .Y(new_n9241_));
  XOR2X1   g09177(.A(new_n9192_), .B(new_n9062_), .Y(new_n9242_));
  XOR2X1   g09178(.A(new_n9199_), .B(new_n9242_), .Y(new_n9243_));
  AOI21X1  g09179(.A0(new_n9065_), .A1(new_n9064_), .B0(new_n8988_), .Y(new_n9244_));
  NOR3X1   g09180(.A(new_n8987_), .B(new_n8983_), .C(new_n8982_), .Y(new_n9245_));
  NAND3X1  g09181(.A(new_n8798_), .B(new_n8793_), .C(new_n8970_), .Y(new_n9246_));
  INVX1    g09182(.A(new_n9175_), .Y(new_n9247_));
  OAI21X1  g09183(.A0(new_n8971_), .A1(new_n8792_), .B0(new_n8797_), .Y(new_n9248_));
  NAND3X1  g09184(.A(new_n9248_), .B(new_n9247_), .C(new_n9246_), .Y(new_n9249_));
  AOI21X1  g09185(.A0(new_n9248_), .A1(new_n9246_), .B0(new_n9247_), .Y(new_n9250_));
  OAI21X1  g09186(.A0(new_n9182_), .A1(new_n9250_), .B0(new_n9249_), .Y(new_n9251_));
  OAI21X1  g09187(.A0(new_n9245_), .A1(new_n9244_), .B0(new_n9251_), .Y(new_n9252_));
  NAND3X1  g09188(.A(new_n9190_), .B(new_n9186_), .C(new_n9252_), .Y(new_n9253_));
  NOR3X1   g09189(.A(new_n9251_), .B(new_n9245_), .C(new_n9244_), .Y(new_n9254_));
  OAI21X1  g09190(.A0(new_n9254_), .A1(new_n9185_), .B0(new_n9191_), .Y(new_n9255_));
  NAND3X1  g09191(.A(new_n9182_), .B(new_n9178_), .C(new_n9249_), .Y(new_n9256_));
  OAI21X1  g09192(.A0(new_n9250_), .A1(new_n9177_), .B0(new_n9183_), .Y(new_n9257_));
  XOR2X1   g09193(.A(new_n9174_), .B(new_n9172_), .Y(new_n9258_));
  OAI22X1  g09194(.A0(new_n8200_), .A1(new_n2666_), .B0(new_n8205_), .B1(new_n2419_), .Y(new_n9259_));
  AOI21X1  g09195(.A0(new_n6899_), .A1(new_n2423_), .B0(new_n9259_), .Y(new_n9260_));
  OAI21X1  g09196(.A0(new_n8293_), .A1(new_n2665_), .B0(new_n9260_), .Y(new_n9261_));
  XOR2X1   g09197(.A(new_n9261_), .B(new_n89_), .Y(new_n9262_));
  NOR2X1   g09198(.A(new_n9262_), .B(new_n9258_), .Y(new_n9263_));
  XOR2X1   g09199(.A(new_n9171_), .B(new_n9170_), .Y(new_n9264_));
  OAI22X1  g09200(.A0(new_n6964_), .A1(new_n2666_), .B0(new_n8200_), .B1(new_n2419_), .Y(new_n9265_));
  AOI21X1  g09201(.A0(new_n6902_), .A1(new_n2423_), .B0(new_n9265_), .Y(new_n9266_));
  OAI21X1  g09202(.A0(new_n8203_), .A1(new_n2665_), .B0(new_n9266_), .Y(new_n9267_));
  XOR2X1   g09203(.A(new_n9267_), .B(new_n89_), .Y(new_n9268_));
  INVX1    g09204(.A(new_n9268_), .Y(new_n9269_));
  NAND2X1  g09205(.A(new_n9269_), .B(new_n9264_), .Y(new_n9270_));
  XOR2X1   g09206(.A(new_n9168_), .B(new_n9167_), .Y(new_n9271_));
  OAI22X1  g09207(.A0(new_n6960_), .A1(new_n2666_), .B0(new_n6964_), .B1(new_n2419_), .Y(new_n9272_));
  AOI21X1  g09208(.A0(new_n6904_), .A1(new_n2423_), .B0(new_n9272_), .Y(new_n9273_));
  OAI21X1  g09209(.A0(new_n8364_), .A1(new_n2665_), .B0(new_n9273_), .Y(new_n9274_));
  XOR2X1   g09210(.A(new_n9274_), .B(new_n89_), .Y(new_n9275_));
  INVX1    g09211(.A(new_n9275_), .Y(new_n9276_));
  AND2X1   g09212(.A(new_n9276_), .B(new_n9271_), .Y(new_n9277_));
  INVX1    g09213(.A(new_n9277_), .Y(new_n9278_));
  XOR2X1   g09214(.A(new_n9165_), .B(new_n9164_), .Y(new_n9279_));
  INVX1    g09215(.A(new_n8541_), .Y(new_n9280_));
  OAI22X1  g09216(.A0(new_n8349_), .A1(new_n2666_), .B0(new_n6960_), .B1(new_n2419_), .Y(new_n9281_));
  AOI21X1  g09217(.A0(new_n6906_), .A1(new_n2423_), .B0(new_n9281_), .Y(new_n9282_));
  OAI21X1  g09218(.A0(new_n9280_), .A1(new_n2665_), .B0(new_n9282_), .Y(new_n9283_));
  XOR2X1   g09219(.A(new_n9283_), .B(new_n89_), .Y(new_n9284_));
  INVX1    g09220(.A(new_n9284_), .Y(new_n9285_));
  AND2X1   g09221(.A(new_n9285_), .B(new_n9279_), .Y(new_n9286_));
  INVX1    g09222(.A(new_n9286_), .Y(new_n9287_));
  XOR2X1   g09223(.A(new_n9162_), .B(new_n9161_), .Y(new_n9288_));
  OAI22X1  g09224(.A0(new_n8579_), .A1(new_n2666_), .B0(new_n8349_), .B1(new_n2419_), .Y(new_n9289_));
  AOI21X1  g09225(.A0(new_n6909_), .A1(new_n2423_), .B0(new_n9289_), .Y(new_n9290_));
  OAI21X1  g09226(.A0(new_n9075_), .A1(new_n2665_), .B0(new_n9290_), .Y(new_n9291_));
  XOR2X1   g09227(.A(new_n9291_), .B(\a[26] ), .Y(new_n9292_));
  AND2X1   g09228(.A(new_n9292_), .B(new_n9288_), .Y(new_n9293_));
  INVX1    g09229(.A(new_n9293_), .Y(new_n9294_));
  XOR2X1   g09230(.A(new_n9160_), .B(new_n9106_), .Y(new_n9295_));
  OAI22X1  g09231(.A0(new_n6917_), .A1(new_n2666_), .B0(new_n8579_), .B1(new_n2419_), .Y(new_n9296_));
  AOI21X1  g09232(.A0(new_n6911_), .A1(new_n2423_), .B0(new_n9296_), .Y(new_n9297_));
  OAI21X1  g09233(.A0(new_n9082_), .A1(new_n2665_), .B0(new_n9297_), .Y(new_n9298_));
  XOR2X1   g09234(.A(new_n9298_), .B(new_n89_), .Y(new_n9299_));
  INVX1    g09235(.A(new_n9299_), .Y(new_n9300_));
  AND2X1   g09236(.A(new_n9300_), .B(new_n9295_), .Y(new_n9301_));
  INVX1    g09237(.A(new_n9301_), .Y(new_n9302_));
  XOR2X1   g09238(.A(new_n9159_), .B(new_n9113_), .Y(new_n9303_));
  OAI22X1  g09239(.A0(new_n6918_), .A1(new_n2666_), .B0(new_n6917_), .B1(new_n2419_), .Y(new_n9304_));
  AOI21X1  g09240(.A0(new_n6913_), .A1(new_n2423_), .B0(new_n9304_), .Y(new_n9305_));
  OAI21X1  g09241(.A0(new_n8577_), .A1(new_n2665_), .B0(new_n9305_), .Y(new_n9306_));
  XOR2X1   g09242(.A(new_n9306_), .B(\a[26] ), .Y(new_n9307_));
  AND2X1   g09243(.A(new_n9307_), .B(new_n9303_), .Y(new_n9308_));
  INVX1    g09244(.A(new_n9308_), .Y(new_n9309_));
  XOR2X1   g09245(.A(new_n9158_), .B(new_n9122_), .Y(new_n9310_));
  OAI22X1  g09246(.A0(new_n6920_), .A1(new_n2666_), .B0(new_n6918_), .B1(new_n2419_), .Y(new_n9311_));
  AOI21X1  g09247(.A0(new_n6915_), .A1(new_n2423_), .B0(new_n9311_), .Y(new_n9312_));
  OAI21X1  g09248(.A0(new_n9093_), .A1(new_n2665_), .B0(new_n9312_), .Y(new_n9313_));
  XOR2X1   g09249(.A(new_n9313_), .B(\a[26] ), .Y(new_n9314_));
  AND2X1   g09250(.A(new_n9314_), .B(new_n9310_), .Y(new_n9315_));
  INVX1    g09251(.A(new_n9315_), .Y(new_n9316_));
  XOR2X1   g09252(.A(new_n9157_), .B(new_n9130_), .Y(new_n9317_));
  OAI22X1  g09253(.A0(new_n8659_), .A1(new_n2666_), .B0(new_n6920_), .B1(new_n2419_), .Y(new_n9318_));
  AOI21X1  g09254(.A0(new_n8580_), .A1(new_n2423_), .B0(new_n9318_), .Y(new_n9319_));
  OAI21X1  g09255(.A0(new_n8611_), .A1(new_n2665_), .B0(new_n9319_), .Y(new_n9320_));
  XOR2X1   g09256(.A(new_n9320_), .B(\a[26] ), .Y(new_n9321_));
  AND2X1   g09257(.A(new_n9321_), .B(new_n9317_), .Y(new_n9322_));
  INVX1    g09258(.A(new_n9322_), .Y(new_n9323_));
  XOR2X1   g09259(.A(new_n9156_), .B(new_n9138_), .Y(new_n9324_));
  AOI22X1  g09260(.A0(new_n6925_), .A1(new_n2424_), .B0(new_n6923_), .B1(new_n2418_), .Y(new_n9325_));
  OAI21X1  g09261(.A0(new_n6920_), .A1(new_n2626_), .B0(new_n9325_), .Y(new_n9326_));
  AOI21X1  g09262(.A0(new_n8628_), .A1(new_n2301_), .B0(new_n9326_), .Y(new_n9327_));
  XOR2X1   g09263(.A(new_n9327_), .B(\a[26] ), .Y(new_n9328_));
  NOR2X1   g09264(.A(new_n9328_), .B(new_n9324_), .Y(new_n9329_));
  INVX1    g09265(.A(new_n9329_), .Y(new_n9330_));
  AOI22X1  g09266(.A0(new_n6927_), .A1(new_n2424_), .B0(new_n6925_), .B1(new_n2418_), .Y(new_n9331_));
  OAI21X1  g09267(.A0(new_n8659_), .A1(new_n2626_), .B0(new_n9331_), .Y(new_n9332_));
  AOI21X1  g09268(.A0(new_n8663_), .A1(new_n2301_), .B0(new_n9332_), .Y(new_n9333_));
  XOR2X1   g09269(.A(new_n9333_), .B(\a[26] ), .Y(new_n9334_));
  INVX1    g09270(.A(new_n9334_), .Y(new_n9335_));
  XOR2X1   g09271(.A(new_n9154_), .B(new_n9152_), .Y(new_n9336_));
  XOR2X1   g09272(.A(new_n9336_), .B(new_n9334_), .Y(new_n9337_));
  AOI22X1  g09273(.A0(new_n6932_), .A1(new_n2424_), .B0(new_n6927_), .B1(new_n2418_), .Y(new_n9338_));
  OAI21X1  g09274(.A0(new_n8683_), .A1(new_n2626_), .B0(new_n9338_), .Y(new_n9339_));
  AOI21X1  g09275(.A0(new_n8682_), .A1(new_n2301_), .B0(new_n9339_), .Y(new_n9340_));
  XOR2X1   g09276(.A(new_n9340_), .B(\a[26] ), .Y(new_n9341_));
  INVX1    g09277(.A(new_n9341_), .Y(new_n9342_));
  NOR3X1   g09278(.A(new_n9144_), .B(new_n9143_), .C(new_n74_), .Y(new_n9343_));
  XOR2X1   g09279(.A(new_n9147_), .B(\a[29] ), .Y(new_n9344_));
  XOR2X1   g09280(.A(new_n9344_), .B(new_n9343_), .Y(new_n9345_));
  XOR2X1   g09281(.A(new_n9345_), .B(new_n9341_), .Y(new_n9346_));
  NOR2X1   g09282(.A(new_n9144_), .B(new_n74_), .Y(new_n9347_));
  XOR2X1   g09283(.A(new_n9347_), .B(new_n9143_), .Y(new_n9348_));
  OAI22X1  g09284(.A0(new_n8757_), .A1(new_n2666_), .B0(new_n6930_), .B1(new_n2419_), .Y(new_n9349_));
  AOI21X1  g09285(.A0(new_n6927_), .A1(new_n2423_), .B0(new_n9349_), .Y(new_n9350_));
  OAI21X1  g09286(.A0(new_n8705_), .A1(new_n2665_), .B0(new_n9350_), .Y(new_n9351_));
  XOR2X1   g09287(.A(new_n9351_), .B(new_n89_), .Y(new_n9352_));
  NOR2X1   g09288(.A(new_n9352_), .B(new_n9348_), .Y(new_n9353_));
  OAI22X1  g09289(.A0(new_n6936_), .A1(new_n2419_), .B0(new_n8752_), .B1(new_n2626_), .Y(new_n9354_));
  AOI21X1  g09290(.A0(new_n8751_), .A1(new_n2301_), .B0(new_n9354_), .Y(new_n9355_));
  XOR2X1   g09291(.A(new_n9355_), .B(\a[26] ), .Y(new_n9356_));
  NOR2X1   g09292(.A(new_n6936_), .B(new_n2299_), .Y(new_n9357_));
  OAI22X1  g09293(.A0(new_n6936_), .A1(new_n2666_), .B0(new_n8752_), .B1(new_n2419_), .Y(new_n9358_));
  AOI21X1  g09294(.A0(new_n6933_), .A1(new_n2423_), .B0(new_n9358_), .Y(new_n9359_));
  OAI21X1  g09295(.A0(new_n8759_), .A1(new_n2665_), .B0(new_n9359_), .Y(new_n9360_));
  NOR4X1   g09296(.A(new_n9360_), .B(new_n9357_), .C(new_n9356_), .D(new_n89_), .Y(new_n9361_));
  NAND2X1  g09297(.A(new_n9361_), .B(new_n9144_), .Y(new_n9362_));
  XOR2X1   g09298(.A(new_n9361_), .B(new_n9144_), .Y(new_n9363_));
  INVX1    g09299(.A(new_n9363_), .Y(new_n9364_));
  AOI22X1  g09300(.A0(new_n6935_), .A1(new_n2424_), .B0(new_n6933_), .B1(new_n2418_), .Y(new_n9365_));
  OAI21X1  g09301(.A0(new_n6930_), .A1(new_n2626_), .B0(new_n9365_), .Y(new_n9366_));
  AOI21X1  g09302(.A0(new_n8717_), .A1(new_n2301_), .B0(new_n9366_), .Y(new_n9367_));
  XOR2X1   g09303(.A(new_n9367_), .B(\a[26] ), .Y(new_n9368_));
  OAI21X1  g09304(.A0(new_n9368_), .A1(new_n9364_), .B0(new_n9362_), .Y(new_n9369_));
  XOR2X1   g09305(.A(new_n9352_), .B(new_n9348_), .Y(new_n9370_));
  AOI21X1  g09306(.A0(new_n9370_), .A1(new_n9369_), .B0(new_n9353_), .Y(new_n9371_));
  NOR2X1   g09307(.A(new_n9371_), .B(new_n9346_), .Y(new_n9372_));
  AOI21X1  g09308(.A0(new_n9345_), .A1(new_n9342_), .B0(new_n9372_), .Y(new_n9373_));
  NOR2X1   g09309(.A(new_n9373_), .B(new_n9337_), .Y(new_n9374_));
  AOI21X1  g09310(.A0(new_n9336_), .A1(new_n9335_), .B0(new_n9374_), .Y(new_n9375_));
  XOR2X1   g09311(.A(new_n9328_), .B(new_n9324_), .Y(new_n9376_));
  INVX1    g09312(.A(new_n9376_), .Y(new_n9377_));
  OAI21X1  g09313(.A0(new_n9377_), .A1(new_n9375_), .B0(new_n9330_), .Y(new_n9378_));
  INVX1    g09314(.A(new_n9378_), .Y(new_n9379_));
  XOR2X1   g09315(.A(new_n9320_), .B(new_n89_), .Y(new_n9380_));
  XOR2X1   g09316(.A(new_n9380_), .B(new_n9317_), .Y(new_n9381_));
  OAI21X1  g09317(.A0(new_n9381_), .A1(new_n9379_), .B0(new_n9323_), .Y(new_n9382_));
  INVX1    g09318(.A(new_n9382_), .Y(new_n9383_));
  XOR2X1   g09319(.A(new_n9313_), .B(new_n89_), .Y(new_n9384_));
  XOR2X1   g09320(.A(new_n9384_), .B(new_n9310_), .Y(new_n9385_));
  OAI21X1  g09321(.A0(new_n9385_), .A1(new_n9383_), .B0(new_n9316_), .Y(new_n9386_));
  INVX1    g09322(.A(new_n9386_), .Y(new_n9387_));
  XOR2X1   g09323(.A(new_n9306_), .B(new_n89_), .Y(new_n9388_));
  XOR2X1   g09324(.A(new_n9388_), .B(new_n9303_), .Y(new_n9389_));
  OAI21X1  g09325(.A0(new_n9389_), .A1(new_n9387_), .B0(new_n9309_), .Y(new_n9390_));
  INVX1    g09326(.A(new_n9390_), .Y(new_n9391_));
  XOR2X1   g09327(.A(new_n9299_), .B(new_n9295_), .Y(new_n9392_));
  OAI21X1  g09328(.A0(new_n9392_), .A1(new_n9391_), .B0(new_n9302_), .Y(new_n9393_));
  INVX1    g09329(.A(new_n9393_), .Y(new_n9394_));
  XOR2X1   g09330(.A(new_n9291_), .B(new_n89_), .Y(new_n9395_));
  XOR2X1   g09331(.A(new_n9395_), .B(new_n9288_), .Y(new_n9396_));
  OAI21X1  g09332(.A0(new_n9396_), .A1(new_n9394_), .B0(new_n9294_), .Y(new_n9397_));
  INVX1    g09333(.A(new_n9397_), .Y(new_n9398_));
  XOR2X1   g09334(.A(new_n9284_), .B(new_n9279_), .Y(new_n9399_));
  OAI21X1  g09335(.A0(new_n9399_), .A1(new_n9398_), .B0(new_n9287_), .Y(new_n9400_));
  INVX1    g09336(.A(new_n9400_), .Y(new_n9401_));
  XOR2X1   g09337(.A(new_n9275_), .B(new_n9271_), .Y(new_n9402_));
  OAI21X1  g09338(.A0(new_n9402_), .A1(new_n9401_), .B0(new_n9278_), .Y(new_n9403_));
  INVX1    g09339(.A(new_n9403_), .Y(new_n9404_));
  XOR2X1   g09340(.A(new_n9268_), .B(new_n9264_), .Y(new_n9405_));
  OAI21X1  g09341(.A0(new_n9405_), .A1(new_n9404_), .B0(new_n9270_), .Y(new_n9406_));
  XOR2X1   g09342(.A(new_n9262_), .B(new_n9258_), .Y(new_n9407_));
  AOI21X1  g09343(.A0(new_n9407_), .A1(new_n9406_), .B0(new_n9263_), .Y(new_n9408_));
  AOI21X1  g09344(.A0(new_n9257_), .A1(new_n9256_), .B0(new_n9408_), .Y(new_n9409_));
  NAND3X1  g09345(.A(new_n9408_), .B(new_n9257_), .C(new_n9256_), .Y(new_n9410_));
  AOI22X1  g09346(.A0(new_n6894_), .A1(new_n2657_), .B0(new_n6892_), .B1(new_n2696_), .Y(new_n9411_));
  OAI21X1  g09347(.A0(new_n7885_), .A1(new_n2753_), .B0(new_n9411_), .Y(new_n9412_));
  AOI21X1  g09348(.A0(new_n7884_), .A1(new_n2658_), .B0(new_n9412_), .Y(new_n9413_));
  XOR2X1   g09349(.A(new_n9413_), .B(\a[23] ), .Y(new_n9414_));
  INVX1    g09350(.A(new_n9414_), .Y(new_n9415_));
  AOI21X1  g09351(.A0(new_n9415_), .A1(new_n9410_), .B0(new_n9409_), .Y(new_n9416_));
  AOI21X1  g09352(.A0(new_n9255_), .A1(new_n9253_), .B0(new_n9416_), .Y(new_n9417_));
  NAND3X1  g09353(.A(new_n9416_), .B(new_n9255_), .C(new_n9253_), .Y(new_n9418_));
  AOI22X1  g09354(.A0(new_n6885_), .A1(new_n2875_), .B0(new_n6882_), .B1(new_n3099_), .Y(new_n9419_));
  OAI21X1  g09355(.A0(new_n7472_), .A1(new_n3152_), .B0(new_n9419_), .Y(new_n9420_));
  AOI21X1  g09356(.A0(new_n7471_), .A1(new_n2876_), .B0(new_n9420_), .Y(new_n9421_));
  XOR2X1   g09357(.A(new_n9421_), .B(\a[20] ), .Y(new_n9422_));
  INVX1    g09358(.A(new_n9422_), .Y(new_n9423_));
  AOI21X1  g09359(.A0(new_n9423_), .A1(new_n9418_), .B0(new_n9417_), .Y(new_n9424_));
  OR2X1    g09360(.A(new_n9424_), .B(new_n9243_), .Y(new_n9425_));
  XOR2X1   g09361(.A(new_n9199_), .B(new_n9195_), .Y(new_n9426_));
  XOR2X1   g09362(.A(new_n9424_), .B(new_n9426_), .Y(new_n9427_));
  AOI22X1  g09363(.A0(new_n6818_), .A1(new_n3390_), .B0(new_n6745_), .B1(new_n3232_), .Y(new_n9428_));
  OAI21X1  g09364(.A0(new_n7047_), .A1(new_n3545_), .B0(new_n9428_), .Y(new_n9429_));
  AOI21X1  g09365(.A0(new_n7046_), .A1(new_n3234_), .B0(new_n9429_), .Y(new_n9430_));
  XOR2X1   g09366(.A(new_n9430_), .B(\a[17] ), .Y(new_n9431_));
  OAI21X1  g09367(.A0(new_n9431_), .A1(new_n9427_), .B0(new_n9425_), .Y(new_n9432_));
  AOI21X1  g09368(.A0(new_n9432_), .A1(new_n9241_), .B0(new_n9240_), .Y(new_n9433_));
  NOR2X1   g09369(.A(new_n9433_), .B(new_n9232_), .Y(new_n9434_));
  XOR2X1   g09370(.A(new_n9433_), .B(new_n9232_), .Y(new_n9435_));
  AOI22X1  g09371(.A0(new_n7529_), .A1(new_n3908_), .B0(new_n7522_), .B1(new_n3628_), .Y(new_n9436_));
  OAI21X1  g09372(.A0(new_n7581_), .A1(new_n3983_), .B0(new_n9436_), .Y(new_n9437_));
  AOI21X1  g09373(.A0(new_n7565_), .A1(new_n3624_), .B0(new_n9437_), .Y(new_n9438_));
  XOR2X1   g09374(.A(new_n9438_), .B(\a[14] ), .Y(new_n9439_));
  INVX1    g09375(.A(new_n9439_), .Y(new_n9440_));
  AOI21X1  g09376(.A0(new_n9440_), .A1(new_n9435_), .B0(new_n9434_), .Y(new_n9441_));
  OR2X1    g09377(.A(new_n9441_), .B(new_n9231_), .Y(new_n9442_));
  XOR2X1   g09378(.A(new_n9216_), .B(new_n9212_), .Y(new_n9443_));
  XOR2X1   g09379(.A(new_n9441_), .B(new_n9443_), .Y(new_n9444_));
  AOI22X1  g09380(.A0(new_n7590_), .A1(new_n4247_), .B0(new_n7578_), .B1(new_n4078_), .Y(new_n9445_));
  OAI21X1  g09381(.A0(new_n7642_), .A1(new_n4427_), .B0(new_n9445_), .Y(new_n9446_));
  AOI21X1  g09382(.A0(new_n7712_), .A1(new_n4080_), .B0(new_n9446_), .Y(new_n9447_));
  XOR2X1   g09383(.A(new_n9447_), .B(\a[11] ), .Y(new_n9448_));
  OAI21X1  g09384(.A0(new_n9448_), .A1(new_n9444_), .B0(new_n9442_), .Y(new_n9449_));
  AOI22X1  g09385(.A0(new_n7643_), .A1(new_n4428_), .B0(new_n7590_), .B1(new_n4078_), .Y(new_n9450_));
  OAI21X1  g09386(.A0(new_n7642_), .A1(new_n4246_), .B0(new_n9450_), .Y(new_n9451_));
  AOI21X1  g09387(.A0(new_n7718_), .A1(new_n4080_), .B0(new_n9451_), .Y(new_n9452_));
  XOR2X1   g09388(.A(new_n9452_), .B(\a[11] ), .Y(new_n9453_));
  INVX1    g09389(.A(new_n9453_), .Y(new_n9454_));
  XOR2X1   g09390(.A(new_n9217_), .B(new_n9048_), .Y(new_n9455_));
  XOR2X1   g09391(.A(new_n9453_), .B(new_n9449_), .Y(new_n9456_));
  NOR2X1   g09392(.A(new_n9456_), .B(new_n9455_), .Y(new_n9457_));
  AOI21X1  g09393(.A0(new_n9454_), .A1(new_n9449_), .B0(new_n9457_), .Y(new_n9458_));
  OR2X1    g09394(.A(new_n9458_), .B(new_n9229_), .Y(new_n9459_));
  XOR2X1   g09395(.A(new_n9225_), .B(new_n9220_), .Y(new_n9460_));
  XOR2X1   g09396(.A(new_n9458_), .B(new_n9460_), .Y(new_n9461_));
  XOR2X1   g09397(.A(new_n9439_), .B(new_n9435_), .Y(new_n9462_));
  OR2X1    g09398(.A(new_n9431_), .B(new_n9427_), .Y(new_n9463_));
  AND2X1   g09399(.A(new_n9463_), .B(new_n9425_), .Y(new_n9464_));
  XOR2X1   g09400(.A(new_n9464_), .B(new_n9241_), .Y(new_n9465_));
  AOI22X1  g09401(.A0(new_n7522_), .A1(new_n3908_), .B0(new_n7485_), .B1(new_n3628_), .Y(new_n9466_));
  OAI21X1  g09402(.A0(new_n7537_), .A1(new_n3983_), .B0(new_n9466_), .Y(new_n9467_));
  AOI21X1  g09403(.A0(new_n7536_), .A1(new_n3624_), .B0(new_n9467_), .Y(new_n9468_));
  XOR2X1   g09404(.A(new_n9468_), .B(\a[14] ), .Y(new_n9469_));
  NOR2X1   g09405(.A(new_n9469_), .B(new_n9465_), .Y(new_n9470_));
  XOR2X1   g09406(.A(new_n9469_), .B(new_n9465_), .Y(new_n9471_));
  XOR2X1   g09407(.A(new_n9424_), .B(new_n9243_), .Y(new_n9472_));
  XOR2X1   g09408(.A(new_n9431_), .B(new_n9472_), .Y(new_n9473_));
  NOR3X1   g09409(.A(new_n9191_), .B(new_n9254_), .C(new_n9185_), .Y(new_n9474_));
  AOI21X1  g09410(.A0(new_n9186_), .A1(new_n9252_), .B0(new_n9190_), .Y(new_n9475_));
  NOR3X1   g09411(.A(new_n9183_), .B(new_n9250_), .C(new_n9177_), .Y(new_n9476_));
  AOI21X1  g09412(.A0(new_n9178_), .A1(new_n9249_), .B0(new_n9182_), .Y(new_n9477_));
  INVX1    g09413(.A(new_n9408_), .Y(new_n9478_));
  OAI21X1  g09414(.A0(new_n9477_), .A1(new_n9476_), .B0(new_n9478_), .Y(new_n9479_));
  NOR3X1   g09415(.A(new_n9478_), .B(new_n9477_), .C(new_n9476_), .Y(new_n9480_));
  OAI21X1  g09416(.A0(new_n9414_), .A1(new_n9480_), .B0(new_n9479_), .Y(new_n9481_));
  OAI21X1  g09417(.A0(new_n9475_), .A1(new_n9474_), .B0(new_n9481_), .Y(new_n9482_));
  NAND3X1  g09418(.A(new_n9422_), .B(new_n9418_), .C(new_n9482_), .Y(new_n9483_));
  NOR3X1   g09419(.A(new_n9481_), .B(new_n9475_), .C(new_n9474_), .Y(new_n9484_));
  OAI21X1  g09420(.A0(new_n9484_), .A1(new_n9417_), .B0(new_n9423_), .Y(new_n9485_));
  NAND3X1  g09421(.A(new_n9414_), .B(new_n9410_), .C(new_n9479_), .Y(new_n9486_));
  OAI21X1  g09422(.A0(new_n9480_), .A1(new_n9409_), .B0(new_n9415_), .Y(new_n9487_));
  AOI22X1  g09423(.A0(new_n6897_), .A1(new_n2657_), .B0(new_n6894_), .B1(new_n2696_), .Y(new_n9488_));
  OAI21X1  g09424(.A0(new_n8075_), .A1(new_n2753_), .B0(new_n9488_), .Y(new_n9489_));
  AOI21X1  g09425(.A0(new_n8074_), .A1(new_n2658_), .B0(new_n9489_), .Y(new_n9490_));
  XOR2X1   g09426(.A(new_n9490_), .B(\a[23] ), .Y(new_n9491_));
  INVX1    g09427(.A(new_n9491_), .Y(new_n9492_));
  XOR2X1   g09428(.A(new_n9407_), .B(new_n9406_), .Y(new_n9493_));
  AND2X1   g09429(.A(new_n9493_), .B(new_n9492_), .Y(new_n9494_));
  XOR2X1   g09430(.A(new_n9493_), .B(new_n9491_), .Y(new_n9495_));
  AOI22X1  g09431(.A0(new_n6899_), .A1(new_n2657_), .B0(new_n6897_), .B1(new_n2696_), .Y(new_n9496_));
  OAI21X1  g09432(.A0(new_n6896_), .A1(new_n2753_), .B0(new_n9496_), .Y(new_n9497_));
  AOI21X1  g09433(.A0(new_n7953_), .A1(new_n2658_), .B0(new_n9497_), .Y(new_n9498_));
  XOR2X1   g09434(.A(new_n9498_), .B(\a[23] ), .Y(new_n9499_));
  XOR2X1   g09435(.A(new_n9405_), .B(new_n9403_), .Y(new_n9500_));
  OR2X1    g09436(.A(new_n9500_), .B(new_n9499_), .Y(new_n9501_));
  XOR2X1   g09437(.A(new_n9500_), .B(new_n9499_), .Y(new_n9502_));
  INVX1    g09438(.A(new_n9502_), .Y(new_n9503_));
  AOI22X1  g09439(.A0(new_n6902_), .A1(new_n2657_), .B0(new_n6899_), .B1(new_n2696_), .Y(new_n9504_));
  OAI21X1  g09440(.A0(new_n6898_), .A1(new_n2753_), .B0(new_n9504_), .Y(new_n9505_));
  AOI21X1  g09441(.A0(new_n8215_), .A1(new_n2658_), .B0(new_n9505_), .Y(new_n9506_));
  XOR2X1   g09442(.A(new_n9506_), .B(\a[23] ), .Y(new_n9507_));
  XOR2X1   g09443(.A(new_n9402_), .B(new_n9400_), .Y(new_n9508_));
  NOR2X1   g09444(.A(new_n9508_), .B(new_n9507_), .Y(new_n9509_));
  XOR2X1   g09445(.A(new_n9508_), .B(new_n9507_), .Y(new_n9510_));
  AOI22X1  g09446(.A0(new_n6904_), .A1(new_n2657_), .B0(new_n6902_), .B1(new_n2696_), .Y(new_n9511_));
  OAI21X1  g09447(.A0(new_n8295_), .A1(new_n2753_), .B0(new_n9511_), .Y(new_n9512_));
  AOI21X1  g09448(.A0(new_n8883_), .A1(new_n2658_), .B0(new_n9512_), .Y(new_n9513_));
  XOR2X1   g09449(.A(new_n9513_), .B(\a[23] ), .Y(new_n9514_));
  XOR2X1   g09450(.A(new_n9399_), .B(new_n9397_), .Y(new_n9515_));
  OR2X1    g09451(.A(new_n9515_), .B(new_n9514_), .Y(new_n9516_));
  XOR2X1   g09452(.A(new_n9515_), .B(new_n9514_), .Y(new_n9517_));
  INVX1    g09453(.A(new_n9517_), .Y(new_n9518_));
  AOI22X1  g09454(.A0(new_n6906_), .A1(new_n2657_), .B0(new_n6904_), .B1(new_n2696_), .Y(new_n9519_));
  OAI21X1  g09455(.A0(new_n8205_), .A1(new_n2753_), .B0(new_n9519_), .Y(new_n9520_));
  AOI21X1  g09456(.A0(new_n8204_), .A1(new_n2658_), .B0(new_n9520_), .Y(new_n9521_));
  XOR2X1   g09457(.A(new_n9521_), .B(\a[23] ), .Y(new_n9522_));
  XOR2X1   g09458(.A(new_n9396_), .B(new_n9393_), .Y(new_n9523_));
  NOR2X1   g09459(.A(new_n9523_), .B(new_n9522_), .Y(new_n9524_));
  XOR2X1   g09460(.A(new_n9523_), .B(new_n9522_), .Y(new_n9525_));
  AOI22X1  g09461(.A0(new_n6909_), .A1(new_n2657_), .B0(new_n6906_), .B1(new_n2696_), .Y(new_n9526_));
  OAI21X1  g09462(.A0(new_n8200_), .A1(new_n2753_), .B0(new_n9526_), .Y(new_n9527_));
  AOI21X1  g09463(.A0(new_n8365_), .A1(new_n2658_), .B0(new_n9527_), .Y(new_n9528_));
  XOR2X1   g09464(.A(new_n9528_), .B(\a[23] ), .Y(new_n9529_));
  XOR2X1   g09465(.A(new_n9392_), .B(new_n9390_), .Y(new_n9530_));
  OR2X1    g09466(.A(new_n9530_), .B(new_n9529_), .Y(new_n9531_));
  XOR2X1   g09467(.A(new_n9530_), .B(new_n9529_), .Y(new_n9532_));
  INVX1    g09468(.A(new_n9532_), .Y(new_n9533_));
  AOI22X1  g09469(.A0(new_n6911_), .A1(new_n2657_), .B0(new_n6909_), .B1(new_n2696_), .Y(new_n9534_));
  OAI21X1  g09470(.A0(new_n6964_), .A1(new_n2753_), .B0(new_n9534_), .Y(new_n9535_));
  AOI21X1  g09471(.A0(new_n8541_), .A1(new_n2658_), .B0(new_n9535_), .Y(new_n9536_));
  XOR2X1   g09472(.A(new_n9536_), .B(\a[23] ), .Y(new_n9537_));
  XOR2X1   g09473(.A(new_n9389_), .B(new_n9386_), .Y(new_n9538_));
  NOR2X1   g09474(.A(new_n9538_), .B(new_n9537_), .Y(new_n9539_));
  XOR2X1   g09475(.A(new_n9538_), .B(new_n9537_), .Y(new_n9540_));
  AOI22X1  g09476(.A0(new_n6913_), .A1(new_n2657_), .B0(new_n6911_), .B1(new_n2696_), .Y(new_n9541_));
  OAI21X1  g09477(.A0(new_n6960_), .A1(new_n2753_), .B0(new_n9541_), .Y(new_n9542_));
  AOI21X1  g09478(.A0(new_n8553_), .A1(new_n2658_), .B0(new_n9542_), .Y(new_n9543_));
  XOR2X1   g09479(.A(new_n9543_), .B(\a[23] ), .Y(new_n9544_));
  XOR2X1   g09480(.A(new_n9385_), .B(new_n9382_), .Y(new_n9545_));
  OR2X1    g09481(.A(new_n9545_), .B(new_n9544_), .Y(new_n9546_));
  XOR2X1   g09482(.A(new_n9545_), .B(new_n9544_), .Y(new_n9547_));
  INVX1    g09483(.A(new_n9547_), .Y(new_n9548_));
  AOI22X1  g09484(.A0(new_n6915_), .A1(new_n2657_), .B0(new_n6913_), .B1(new_n2696_), .Y(new_n9549_));
  OAI21X1  g09485(.A0(new_n8349_), .A1(new_n2753_), .B0(new_n9549_), .Y(new_n9550_));
  AOI21X1  g09486(.A0(new_n8348_), .A1(new_n2658_), .B0(new_n9550_), .Y(new_n9551_));
  XOR2X1   g09487(.A(new_n9551_), .B(\a[23] ), .Y(new_n9552_));
  XOR2X1   g09488(.A(new_n9381_), .B(new_n9378_), .Y(new_n9553_));
  NOR2X1   g09489(.A(new_n9553_), .B(new_n9552_), .Y(new_n9554_));
  XOR2X1   g09490(.A(new_n9553_), .B(new_n9552_), .Y(new_n9555_));
  AOI22X1  g09491(.A0(new_n8580_), .A1(new_n2657_), .B0(new_n6915_), .B1(new_n2696_), .Y(new_n9556_));
  OAI21X1  g09492(.A0(new_n8579_), .A1(new_n2753_), .B0(new_n9556_), .Y(new_n9557_));
  AOI21X1  g09493(.A0(new_n8578_), .A1(new_n2658_), .B0(new_n9557_), .Y(new_n9558_));
  XOR2X1   g09494(.A(new_n9558_), .B(\a[23] ), .Y(new_n9559_));
  XOR2X1   g09495(.A(new_n9376_), .B(new_n9375_), .Y(new_n9560_));
  OR2X1    g09496(.A(new_n9560_), .B(new_n9559_), .Y(new_n9561_));
  XOR2X1   g09497(.A(new_n9560_), .B(new_n9559_), .Y(new_n9562_));
  INVX1    g09498(.A(new_n9562_), .Y(new_n9563_));
  INVX1    g09499(.A(new_n9337_), .Y(new_n9564_));
  XOR2X1   g09500(.A(new_n9373_), .B(new_n9564_), .Y(new_n9565_));
  OAI22X1  g09501(.A0(new_n6920_), .A1(new_n4016_), .B0(new_n6918_), .B1(new_n2743_), .Y(new_n9566_));
  AOI21X1  g09502(.A0(new_n6915_), .A1(new_n2745_), .B0(new_n9566_), .Y(new_n9567_));
  OAI21X1  g09503(.A0(new_n9093_), .A1(new_n2692_), .B0(new_n9567_), .Y(new_n9568_));
  XOR2X1   g09504(.A(new_n9568_), .B(new_n70_), .Y(new_n9569_));
  NOR2X1   g09505(.A(new_n9569_), .B(new_n9565_), .Y(new_n9570_));
  XOR2X1   g09506(.A(new_n9371_), .B(new_n9346_), .Y(new_n9571_));
  INVX1    g09507(.A(new_n9571_), .Y(new_n9572_));
  OAI22X1  g09508(.A0(new_n8659_), .A1(new_n4016_), .B0(new_n6920_), .B1(new_n2743_), .Y(new_n9573_));
  AOI21X1  g09509(.A0(new_n8580_), .A1(new_n2745_), .B0(new_n9573_), .Y(new_n9574_));
  OAI21X1  g09510(.A0(new_n8611_), .A1(new_n2692_), .B0(new_n9574_), .Y(new_n9575_));
  XOR2X1   g09511(.A(new_n9575_), .B(new_n70_), .Y(new_n9576_));
  OR2X1    g09512(.A(new_n9576_), .B(new_n9572_), .Y(new_n9577_));
  AOI22X1  g09513(.A0(new_n6925_), .A1(new_n2657_), .B0(new_n6923_), .B1(new_n2696_), .Y(new_n9578_));
  OAI21X1  g09514(.A0(new_n6920_), .A1(new_n2753_), .B0(new_n9578_), .Y(new_n9579_));
  AOI21X1  g09515(.A0(new_n8628_), .A1(new_n2658_), .B0(new_n9579_), .Y(new_n9580_));
  XOR2X1   g09516(.A(new_n9580_), .B(\a[23] ), .Y(new_n9581_));
  INVX1    g09517(.A(new_n9581_), .Y(new_n9582_));
  XOR2X1   g09518(.A(new_n9370_), .B(new_n9369_), .Y(new_n9583_));
  AND2X1   g09519(.A(new_n9583_), .B(new_n9582_), .Y(new_n9584_));
  INVX1    g09520(.A(new_n9584_), .Y(new_n9585_));
  XOR2X1   g09521(.A(new_n9583_), .B(new_n9581_), .Y(new_n9586_));
  XOR2X1   g09522(.A(new_n9368_), .B(new_n9363_), .Y(new_n9587_));
  OAI22X1  g09523(.A0(new_n6929_), .A1(new_n4016_), .B0(new_n8683_), .B1(new_n2743_), .Y(new_n9588_));
  AOI21X1  g09524(.A0(new_n6923_), .A1(new_n2745_), .B0(new_n9588_), .Y(new_n9589_));
  OAI21X1  g09525(.A0(new_n8662_), .A1(new_n2692_), .B0(new_n9589_), .Y(new_n9590_));
  XOR2X1   g09526(.A(new_n9590_), .B(new_n70_), .Y(new_n9591_));
  NOR2X1   g09527(.A(new_n9591_), .B(new_n9587_), .Y(new_n9592_));
  AOI22X1  g09528(.A0(new_n6932_), .A1(new_n2657_), .B0(new_n6927_), .B1(new_n2696_), .Y(new_n9593_));
  OAI21X1  g09529(.A0(new_n8683_), .A1(new_n2753_), .B0(new_n9593_), .Y(new_n9594_));
  AOI21X1  g09530(.A0(new_n8682_), .A1(new_n2658_), .B0(new_n9594_), .Y(new_n9595_));
  XOR2X1   g09531(.A(new_n9595_), .B(\a[23] ), .Y(new_n9596_));
  NOR3X1   g09532(.A(new_n9357_), .B(new_n9356_), .C(new_n89_), .Y(new_n9597_));
  XOR2X1   g09533(.A(new_n9360_), .B(\a[26] ), .Y(new_n9598_));
  NOR2X1   g09534(.A(new_n9598_), .B(new_n9597_), .Y(new_n9599_));
  NOR3X1   g09535(.A(new_n9599_), .B(new_n9596_), .C(new_n9361_), .Y(new_n9600_));
  XOR2X1   g09536(.A(new_n9598_), .B(new_n9597_), .Y(new_n9601_));
  XOR2X1   g09537(.A(new_n9601_), .B(new_n9596_), .Y(new_n9602_));
  NOR2X1   g09538(.A(new_n9357_), .B(new_n89_), .Y(new_n9603_));
  XOR2X1   g09539(.A(new_n9603_), .B(new_n9356_), .Y(new_n9604_));
  OAI22X1  g09540(.A0(new_n8757_), .A1(new_n4016_), .B0(new_n6930_), .B1(new_n2743_), .Y(new_n9605_));
  AOI21X1  g09541(.A0(new_n6927_), .A1(new_n2745_), .B0(new_n9605_), .Y(new_n9606_));
  OAI21X1  g09542(.A0(new_n8705_), .A1(new_n2692_), .B0(new_n9606_), .Y(new_n9607_));
  XOR2X1   g09543(.A(new_n9607_), .B(new_n70_), .Y(new_n9608_));
  NOR2X1   g09544(.A(new_n9608_), .B(new_n9604_), .Y(new_n9609_));
  OAI22X1  g09545(.A0(new_n6936_), .A1(new_n2743_), .B0(new_n8752_), .B1(new_n2753_), .Y(new_n9610_));
  AOI21X1  g09546(.A0(new_n8751_), .A1(new_n2658_), .B0(new_n9610_), .Y(new_n9611_));
  XOR2X1   g09547(.A(new_n9611_), .B(\a[23] ), .Y(new_n9612_));
  NOR2X1   g09548(.A(new_n6936_), .B(new_n2655_), .Y(new_n9613_));
  OAI22X1  g09549(.A0(new_n6936_), .A1(new_n4016_), .B0(new_n8752_), .B1(new_n2743_), .Y(new_n9614_));
  AOI21X1  g09550(.A0(new_n6933_), .A1(new_n2745_), .B0(new_n9614_), .Y(new_n9615_));
  OAI21X1  g09551(.A0(new_n8759_), .A1(new_n2692_), .B0(new_n9615_), .Y(new_n9616_));
  NOR4X1   g09552(.A(new_n9616_), .B(new_n9613_), .C(new_n9612_), .D(new_n70_), .Y(new_n9617_));
  NAND2X1  g09553(.A(new_n9617_), .B(new_n9357_), .Y(new_n9618_));
  XOR2X1   g09554(.A(new_n9617_), .B(new_n9357_), .Y(new_n9619_));
  INVX1    g09555(.A(new_n9619_), .Y(new_n9620_));
  AOI22X1  g09556(.A0(new_n6935_), .A1(new_n2657_), .B0(new_n6933_), .B1(new_n2696_), .Y(new_n9621_));
  OAI21X1  g09557(.A0(new_n6930_), .A1(new_n2753_), .B0(new_n9621_), .Y(new_n9622_));
  AOI21X1  g09558(.A0(new_n8717_), .A1(new_n2658_), .B0(new_n9622_), .Y(new_n9623_));
  XOR2X1   g09559(.A(new_n9623_), .B(\a[23] ), .Y(new_n9624_));
  OAI21X1  g09560(.A0(new_n9624_), .A1(new_n9620_), .B0(new_n9618_), .Y(new_n9625_));
  XOR2X1   g09561(.A(new_n9608_), .B(new_n9604_), .Y(new_n9626_));
  AOI21X1  g09562(.A0(new_n9626_), .A1(new_n9625_), .B0(new_n9609_), .Y(new_n9627_));
  NOR2X1   g09563(.A(new_n9627_), .B(new_n9602_), .Y(new_n9628_));
  OR2X1    g09564(.A(new_n9628_), .B(new_n9600_), .Y(new_n9629_));
  XOR2X1   g09565(.A(new_n9591_), .B(new_n9587_), .Y(new_n9630_));
  AOI21X1  g09566(.A0(new_n9630_), .A1(new_n9629_), .B0(new_n9592_), .Y(new_n9631_));
  OAI21X1  g09567(.A0(new_n9631_), .A1(new_n9586_), .B0(new_n9585_), .Y(new_n9632_));
  INVX1    g09568(.A(new_n9632_), .Y(new_n9633_));
  XOR2X1   g09569(.A(new_n9576_), .B(new_n9571_), .Y(new_n9634_));
  OAI21X1  g09570(.A0(new_n9634_), .A1(new_n9633_), .B0(new_n9577_), .Y(new_n9635_));
  XOR2X1   g09571(.A(new_n9569_), .B(new_n9565_), .Y(new_n9636_));
  AOI21X1  g09572(.A0(new_n9636_), .A1(new_n9635_), .B0(new_n9570_), .Y(new_n9637_));
  OAI21X1  g09573(.A0(new_n9637_), .A1(new_n9563_), .B0(new_n9561_), .Y(new_n9638_));
  AOI21X1  g09574(.A0(new_n9638_), .A1(new_n9555_), .B0(new_n9554_), .Y(new_n9639_));
  OAI21X1  g09575(.A0(new_n9639_), .A1(new_n9548_), .B0(new_n9546_), .Y(new_n9640_));
  AOI21X1  g09576(.A0(new_n9640_), .A1(new_n9540_), .B0(new_n9539_), .Y(new_n9641_));
  OAI21X1  g09577(.A0(new_n9641_), .A1(new_n9533_), .B0(new_n9531_), .Y(new_n9642_));
  AOI21X1  g09578(.A0(new_n9642_), .A1(new_n9525_), .B0(new_n9524_), .Y(new_n9643_));
  OAI21X1  g09579(.A0(new_n9643_), .A1(new_n9518_), .B0(new_n9516_), .Y(new_n9644_));
  AOI21X1  g09580(.A0(new_n9644_), .A1(new_n9510_), .B0(new_n9509_), .Y(new_n9645_));
  OR2X1    g09581(.A(new_n9645_), .B(new_n9503_), .Y(new_n9646_));
  AOI21X1  g09582(.A0(new_n9646_), .A1(new_n9501_), .B0(new_n9495_), .Y(new_n9647_));
  NOR2X1   g09583(.A(new_n9647_), .B(new_n9494_), .Y(new_n9648_));
  AOI21X1  g09584(.A0(new_n9487_), .A1(new_n9486_), .B0(new_n9648_), .Y(new_n9649_));
  NAND3X1  g09585(.A(new_n9648_), .B(new_n9487_), .C(new_n9486_), .Y(new_n9650_));
  AOI22X1  g09586(.A0(new_n6887_), .A1(new_n2875_), .B0(new_n6885_), .B1(new_n3099_), .Y(new_n9651_));
  OAI21X1  g09587(.A0(new_n6884_), .A1(new_n3152_), .B0(new_n9651_), .Y(new_n9652_));
  AOI21X1  g09588(.A0(new_n7771_), .A1(new_n2876_), .B0(new_n9652_), .Y(new_n9653_));
  XOR2X1   g09589(.A(new_n9653_), .B(\a[20] ), .Y(new_n9654_));
  INVX1    g09590(.A(new_n9654_), .Y(new_n9655_));
  AOI21X1  g09591(.A0(new_n9655_), .A1(new_n9650_), .B0(new_n9649_), .Y(new_n9656_));
  AOI21X1  g09592(.A0(new_n9485_), .A1(new_n9483_), .B0(new_n9656_), .Y(new_n9657_));
  NAND3X1  g09593(.A(new_n9656_), .B(new_n9485_), .C(new_n9483_), .Y(new_n9658_));
  AOI22X1  g09594(.A0(new_n6820_), .A1(new_n3232_), .B0(new_n6745_), .B1(new_n3390_), .Y(new_n9659_));
  OAI21X1  g09595(.A0(new_n7361_), .A1(new_n3545_), .B0(new_n9659_), .Y(new_n9660_));
  AOI21X1  g09596(.A0(new_n7404_), .A1(new_n3234_), .B0(new_n9660_), .Y(new_n9661_));
  XOR2X1   g09597(.A(new_n9661_), .B(\a[17] ), .Y(new_n9662_));
  INVX1    g09598(.A(new_n9662_), .Y(new_n9663_));
  AOI21X1  g09599(.A0(new_n9663_), .A1(new_n9658_), .B0(new_n9657_), .Y(new_n9664_));
  OR2X1    g09600(.A(new_n9664_), .B(new_n9473_), .Y(new_n9665_));
  XOR2X1   g09601(.A(new_n9431_), .B(new_n9427_), .Y(new_n9666_));
  XOR2X1   g09602(.A(new_n9664_), .B(new_n9666_), .Y(new_n9667_));
  AOI22X1  g09603(.A0(new_n7485_), .A1(new_n3908_), .B0(new_n7364_), .B1(new_n3628_), .Y(new_n9668_));
  OAI21X1  g09604(.A0(new_n7523_), .A1(new_n3983_), .B0(new_n9668_), .Y(new_n9669_));
  AOI21X1  g09605(.A0(new_n7612_), .A1(new_n3624_), .B0(new_n9669_), .Y(new_n9670_));
  XOR2X1   g09606(.A(new_n9670_), .B(\a[14] ), .Y(new_n9671_));
  OAI21X1  g09607(.A0(new_n9671_), .A1(new_n9667_), .B0(new_n9665_), .Y(new_n9672_));
  AOI21X1  g09608(.A0(new_n9672_), .A1(new_n9471_), .B0(new_n9470_), .Y(new_n9673_));
  NOR2X1   g09609(.A(new_n9673_), .B(new_n9462_), .Y(new_n9674_));
  XOR2X1   g09610(.A(new_n9673_), .B(new_n9462_), .Y(new_n9675_));
  AOI22X1  g09611(.A0(new_n7578_), .A1(new_n4247_), .B0(new_n7571_), .B1(new_n4078_), .Y(new_n9676_));
  OAI21X1  g09612(.A0(new_n7594_), .A1(new_n4427_), .B0(new_n9676_), .Y(new_n9677_));
  AOI21X1  g09613(.A0(new_n7593_), .A1(new_n4080_), .B0(new_n9677_), .Y(new_n9678_));
  XOR2X1   g09614(.A(new_n9678_), .B(new_n2911_), .Y(new_n9679_));
  AOI21X1  g09615(.A0(new_n9679_), .A1(new_n9675_), .B0(new_n9674_), .Y(new_n9680_));
  NAND2X1  g09616(.A(new_n5096_), .B(new_n4869_), .Y(new_n9681_));
  AOI22X1  g09617(.A0(new_n9681_), .A1(new_n7341_), .B0(new_n7643_), .B1(new_n4635_), .Y(new_n9682_));
  OAI21X1  g09618(.A0(new_n7808_), .A1(new_n4868_), .B0(new_n9682_), .Y(new_n9683_));
  XOR2X1   g09619(.A(new_n9683_), .B(new_n2995_), .Y(new_n9684_));
  OR2X1    g09620(.A(new_n9684_), .B(new_n9680_), .Y(new_n9685_));
  XOR2X1   g09621(.A(new_n9448_), .B(new_n9444_), .Y(new_n9686_));
  XOR2X1   g09622(.A(new_n9684_), .B(new_n9680_), .Y(new_n9687_));
  NAND2X1  g09623(.A(new_n9687_), .B(new_n9686_), .Y(new_n9688_));
  NAND2X1  g09624(.A(new_n9688_), .B(new_n9685_), .Y(new_n9689_));
  XOR2X1   g09625(.A(new_n9456_), .B(new_n9455_), .Y(new_n9690_));
  AND2X1   g09626(.A(new_n9690_), .B(new_n9689_), .Y(new_n9691_));
  XOR2X1   g09627(.A(new_n9441_), .B(new_n9231_), .Y(new_n9692_));
  XOR2X1   g09628(.A(new_n9448_), .B(new_n9692_), .Y(new_n9693_));
  XOR2X1   g09629(.A(new_n9687_), .B(new_n9693_), .Y(new_n9694_));
  XOR2X1   g09630(.A(new_n9679_), .B(new_n9675_), .Y(new_n9695_));
  OR2X1    g09631(.A(new_n9671_), .B(new_n9667_), .Y(new_n9696_));
  AND2X1   g09632(.A(new_n9696_), .B(new_n9665_), .Y(new_n9697_));
  XOR2X1   g09633(.A(new_n9697_), .B(new_n9471_), .Y(new_n9698_));
  AOI22X1  g09634(.A0(new_n7571_), .A1(new_n4247_), .B0(new_n7558_), .B1(new_n4078_), .Y(new_n9699_));
  OAI21X1  g09635(.A0(new_n7602_), .A1(new_n4427_), .B0(new_n9699_), .Y(new_n9700_));
  AOI21X1  g09636(.A0(new_n7601_), .A1(new_n4080_), .B0(new_n9700_), .Y(new_n9701_));
  XOR2X1   g09637(.A(new_n9701_), .B(\a[11] ), .Y(new_n9702_));
  NOR2X1   g09638(.A(new_n9702_), .B(new_n9698_), .Y(new_n9703_));
  INVX1    g09639(.A(new_n9702_), .Y(new_n9704_));
  XOR2X1   g09640(.A(new_n9704_), .B(new_n9698_), .Y(new_n9705_));
  XOR2X1   g09641(.A(new_n9664_), .B(new_n9473_), .Y(new_n9706_));
  XOR2X1   g09642(.A(new_n9671_), .B(new_n9706_), .Y(new_n9707_));
  NOR3X1   g09643(.A(new_n9423_), .B(new_n9484_), .C(new_n9417_), .Y(new_n9708_));
  AOI21X1  g09644(.A0(new_n9418_), .A1(new_n9482_), .B0(new_n9422_), .Y(new_n9709_));
  NOR3X1   g09645(.A(new_n9415_), .B(new_n9480_), .C(new_n9409_), .Y(new_n9710_));
  AOI21X1  g09646(.A0(new_n9410_), .A1(new_n9479_), .B0(new_n9414_), .Y(new_n9711_));
  INVX1    g09647(.A(new_n9648_), .Y(new_n9712_));
  OAI21X1  g09648(.A0(new_n9711_), .A1(new_n9710_), .B0(new_n9712_), .Y(new_n9713_));
  NOR3X1   g09649(.A(new_n9712_), .B(new_n9711_), .C(new_n9710_), .Y(new_n9714_));
  OAI21X1  g09650(.A0(new_n9654_), .A1(new_n9714_), .B0(new_n9713_), .Y(new_n9715_));
  OAI21X1  g09651(.A0(new_n9709_), .A1(new_n9708_), .B0(new_n9715_), .Y(new_n9716_));
  NAND3X1  g09652(.A(new_n9662_), .B(new_n9658_), .C(new_n9716_), .Y(new_n9717_));
  NOR3X1   g09653(.A(new_n9715_), .B(new_n9709_), .C(new_n9708_), .Y(new_n9718_));
  OAI21X1  g09654(.A0(new_n9718_), .A1(new_n9657_), .B0(new_n9663_), .Y(new_n9719_));
  NAND3X1  g09655(.A(new_n9654_), .B(new_n9650_), .C(new_n9713_), .Y(new_n9720_));
  OAI21X1  g09656(.A0(new_n9714_), .A1(new_n9649_), .B0(new_n9655_), .Y(new_n9721_));
  AND2X1   g09657(.A(new_n9646_), .B(new_n9501_), .Y(new_n9722_));
  XOR2X1   g09658(.A(new_n9722_), .B(new_n9495_), .Y(new_n9723_));
  INVX1    g09659(.A(new_n9723_), .Y(new_n9724_));
  OAI22X1  g09660(.A0(new_n7885_), .A1(new_n3250_), .B0(new_n7878_), .B1(new_n3144_), .Y(new_n9725_));
  AOI21X1  g09661(.A0(new_n6885_), .A1(new_n3146_), .B0(new_n9725_), .Y(new_n9726_));
  OAI21X1  g09662(.A0(new_n8083_), .A1(new_n3098_), .B0(new_n9726_), .Y(new_n9727_));
  XOR2X1   g09663(.A(new_n9727_), .B(new_n1920_), .Y(new_n9728_));
  NOR2X1   g09664(.A(new_n9728_), .B(new_n9724_), .Y(new_n9729_));
  XOR2X1   g09665(.A(new_n9645_), .B(new_n9503_), .Y(new_n9730_));
  OAI22X1  g09666(.A0(new_n8075_), .A1(new_n3250_), .B0(new_n7885_), .B1(new_n3144_), .Y(new_n9731_));
  AOI21X1  g09667(.A0(new_n6887_), .A1(new_n3146_), .B0(new_n9731_), .Y(new_n9732_));
  OAI21X1  g09668(.A0(new_n7876_), .A1(new_n3098_), .B0(new_n9732_), .Y(new_n9733_));
  XOR2X1   g09669(.A(new_n9733_), .B(new_n1920_), .Y(new_n9734_));
  INVX1    g09670(.A(new_n9734_), .Y(new_n9735_));
  NAND2X1  g09671(.A(new_n9735_), .B(new_n9730_), .Y(new_n9736_));
  XOR2X1   g09672(.A(new_n9644_), .B(new_n9510_), .Y(new_n9737_));
  INVX1    g09673(.A(new_n7884_), .Y(new_n9738_));
  OAI22X1  g09674(.A0(new_n6896_), .A1(new_n3250_), .B0(new_n8075_), .B1(new_n3144_), .Y(new_n9739_));
  AOI21X1  g09675(.A0(new_n6890_), .A1(new_n3146_), .B0(new_n9739_), .Y(new_n9740_));
  OAI21X1  g09676(.A0(new_n9738_), .A1(new_n3098_), .B0(new_n9740_), .Y(new_n9741_));
  XOR2X1   g09677(.A(new_n9741_), .B(\a[20] ), .Y(new_n9742_));
  XOR2X1   g09678(.A(new_n9643_), .B(new_n9518_), .Y(new_n9743_));
  INVX1    g09679(.A(new_n8074_), .Y(new_n9744_));
  OAI22X1  g09680(.A0(new_n6898_), .A1(new_n3250_), .B0(new_n6896_), .B1(new_n3144_), .Y(new_n9745_));
  AOI21X1  g09681(.A0(new_n6892_), .A1(new_n3146_), .B0(new_n9745_), .Y(new_n9746_));
  OAI21X1  g09682(.A0(new_n9744_), .A1(new_n3098_), .B0(new_n9746_), .Y(new_n9747_));
  XOR2X1   g09683(.A(new_n9747_), .B(\a[20] ), .Y(new_n9748_));
  AND2X1   g09684(.A(new_n9748_), .B(new_n9743_), .Y(new_n9749_));
  XOR2X1   g09685(.A(new_n9642_), .B(new_n9525_), .Y(new_n9750_));
  OAI22X1  g09686(.A0(new_n8295_), .A1(new_n3250_), .B0(new_n6898_), .B1(new_n3144_), .Y(new_n9751_));
  AOI21X1  g09687(.A0(new_n6894_), .A1(new_n3146_), .B0(new_n9751_), .Y(new_n9752_));
  OAI21X1  g09688(.A0(new_n8383_), .A1(new_n3098_), .B0(new_n9752_), .Y(new_n9753_));
  XOR2X1   g09689(.A(new_n9753_), .B(\a[20] ), .Y(new_n9754_));
  AND2X1   g09690(.A(new_n9754_), .B(new_n9750_), .Y(new_n9755_));
  INVX1    g09691(.A(new_n9755_), .Y(new_n9756_));
  XOR2X1   g09692(.A(new_n9641_), .B(new_n9533_), .Y(new_n9757_));
  AOI22X1  g09693(.A0(new_n6902_), .A1(new_n2875_), .B0(new_n6899_), .B1(new_n3099_), .Y(new_n9758_));
  OAI21X1  g09694(.A0(new_n6898_), .A1(new_n3152_), .B0(new_n9758_), .Y(new_n9759_));
  AOI21X1  g09695(.A0(new_n8215_), .A1(new_n2876_), .B0(new_n9759_), .Y(new_n9760_));
  XOR2X1   g09696(.A(new_n9760_), .B(new_n1920_), .Y(new_n9761_));
  AND2X1   g09697(.A(new_n9761_), .B(new_n9757_), .Y(new_n9762_));
  INVX1    g09698(.A(new_n9762_), .Y(new_n9763_));
  XOR2X1   g09699(.A(new_n9640_), .B(new_n9540_), .Y(new_n9764_));
  OAI22X1  g09700(.A0(new_n8200_), .A1(new_n3250_), .B0(new_n8205_), .B1(new_n3144_), .Y(new_n9765_));
  AOI21X1  g09701(.A0(new_n6899_), .A1(new_n3146_), .B0(new_n9765_), .Y(new_n9766_));
  OAI21X1  g09702(.A0(new_n8293_), .A1(new_n3098_), .B0(new_n9766_), .Y(new_n9767_));
  XOR2X1   g09703(.A(new_n9767_), .B(\a[20] ), .Y(new_n9768_));
  AND2X1   g09704(.A(new_n9768_), .B(new_n9764_), .Y(new_n9769_));
  INVX1    g09705(.A(new_n9769_), .Y(new_n9770_));
  XOR2X1   g09706(.A(new_n9639_), .B(new_n9548_), .Y(new_n9771_));
  OAI22X1  g09707(.A0(new_n6964_), .A1(new_n3250_), .B0(new_n8200_), .B1(new_n3144_), .Y(new_n9772_));
  AOI21X1  g09708(.A0(new_n6902_), .A1(new_n3146_), .B0(new_n9772_), .Y(new_n9773_));
  OAI21X1  g09709(.A0(new_n8203_), .A1(new_n3098_), .B0(new_n9773_), .Y(new_n9774_));
  XOR2X1   g09710(.A(new_n9774_), .B(\a[20] ), .Y(new_n9775_));
  AND2X1   g09711(.A(new_n9775_), .B(new_n9771_), .Y(new_n9776_));
  INVX1    g09712(.A(new_n9776_), .Y(new_n9777_));
  XOR2X1   g09713(.A(new_n9638_), .B(new_n9555_), .Y(new_n9778_));
  INVX1    g09714(.A(new_n9778_), .Y(new_n9779_));
  OAI22X1  g09715(.A0(new_n6960_), .A1(new_n3250_), .B0(new_n6964_), .B1(new_n3144_), .Y(new_n9780_));
  AOI21X1  g09716(.A0(new_n6904_), .A1(new_n3146_), .B0(new_n9780_), .Y(new_n9781_));
  OAI21X1  g09717(.A0(new_n8364_), .A1(new_n3098_), .B0(new_n9781_), .Y(new_n9782_));
  XOR2X1   g09718(.A(new_n9782_), .B(new_n1920_), .Y(new_n9783_));
  NOR2X1   g09719(.A(new_n9783_), .B(new_n9779_), .Y(new_n9784_));
  INVX1    g09720(.A(new_n9784_), .Y(new_n9785_));
  XOR2X1   g09721(.A(new_n9637_), .B(new_n9563_), .Y(new_n9786_));
  INVX1    g09722(.A(new_n9786_), .Y(new_n9787_));
  AOI22X1  g09723(.A0(new_n6911_), .A1(new_n2875_), .B0(new_n6909_), .B1(new_n3099_), .Y(new_n9788_));
  OAI21X1  g09724(.A0(new_n6964_), .A1(new_n3152_), .B0(new_n9788_), .Y(new_n9789_));
  AOI21X1  g09725(.A0(new_n8541_), .A1(new_n2876_), .B0(new_n9789_), .Y(new_n9790_));
  XOR2X1   g09726(.A(new_n9790_), .B(\a[20] ), .Y(new_n9791_));
  NOR2X1   g09727(.A(new_n9791_), .B(new_n9787_), .Y(new_n9792_));
  INVX1    g09728(.A(new_n9792_), .Y(new_n9793_));
  AOI22X1  g09729(.A0(new_n6913_), .A1(new_n2875_), .B0(new_n6911_), .B1(new_n3099_), .Y(new_n9794_));
  OAI21X1  g09730(.A0(new_n6960_), .A1(new_n3152_), .B0(new_n9794_), .Y(new_n9795_));
  AOI21X1  g09731(.A0(new_n8553_), .A1(new_n2876_), .B0(new_n9795_), .Y(new_n9796_));
  XOR2X1   g09732(.A(new_n9796_), .B(\a[20] ), .Y(new_n9797_));
  INVX1    g09733(.A(new_n9797_), .Y(new_n9798_));
  XOR2X1   g09734(.A(new_n9636_), .B(new_n9635_), .Y(new_n9799_));
  AND2X1   g09735(.A(new_n9799_), .B(new_n9798_), .Y(new_n9800_));
  XOR2X1   g09736(.A(new_n9799_), .B(new_n9797_), .Y(new_n9801_));
  INVX1    g09737(.A(new_n9801_), .Y(new_n9802_));
  AOI22X1  g09738(.A0(new_n6915_), .A1(new_n2875_), .B0(new_n6913_), .B1(new_n3099_), .Y(new_n9803_));
  OAI21X1  g09739(.A0(new_n8349_), .A1(new_n3152_), .B0(new_n9803_), .Y(new_n9804_));
  AOI21X1  g09740(.A0(new_n8348_), .A1(new_n2876_), .B0(new_n9804_), .Y(new_n9805_));
  XOR2X1   g09741(.A(new_n9805_), .B(\a[20] ), .Y(new_n9806_));
  XOR2X1   g09742(.A(new_n9634_), .B(new_n9632_), .Y(new_n9807_));
  OR2X1    g09743(.A(new_n9807_), .B(new_n9806_), .Y(new_n9808_));
  XOR2X1   g09744(.A(new_n9807_), .B(new_n9806_), .Y(new_n9809_));
  INVX1    g09745(.A(new_n9809_), .Y(new_n9810_));
  INVX1    g09746(.A(new_n9586_), .Y(new_n9811_));
  XOR2X1   g09747(.A(new_n9631_), .B(new_n9811_), .Y(new_n9812_));
  OAI22X1  g09748(.A0(new_n6918_), .A1(new_n3250_), .B0(new_n6917_), .B1(new_n3144_), .Y(new_n9813_));
  AOI21X1  g09749(.A0(new_n6913_), .A1(new_n3146_), .B0(new_n9813_), .Y(new_n9814_));
  OAI21X1  g09750(.A0(new_n8577_), .A1(new_n3098_), .B0(new_n9814_), .Y(new_n9815_));
  XOR2X1   g09751(.A(new_n9815_), .B(new_n1920_), .Y(new_n9816_));
  NOR2X1   g09752(.A(new_n9816_), .B(new_n9812_), .Y(new_n9817_));
  XOR2X1   g09753(.A(new_n9630_), .B(new_n9629_), .Y(new_n9818_));
  INVX1    g09754(.A(new_n9818_), .Y(new_n9819_));
  OAI22X1  g09755(.A0(new_n6920_), .A1(new_n3250_), .B0(new_n6918_), .B1(new_n3144_), .Y(new_n9820_));
  AOI21X1  g09756(.A0(new_n6915_), .A1(new_n3146_), .B0(new_n9820_), .Y(new_n9821_));
  OAI21X1  g09757(.A0(new_n9093_), .A1(new_n3098_), .B0(new_n9821_), .Y(new_n9822_));
  XOR2X1   g09758(.A(new_n9822_), .B(new_n1920_), .Y(new_n9823_));
  OR2X1    g09759(.A(new_n9823_), .B(new_n9819_), .Y(new_n9824_));
  XOR2X1   g09760(.A(new_n9627_), .B(new_n9602_), .Y(new_n9825_));
  INVX1    g09761(.A(new_n9825_), .Y(new_n9826_));
  OAI22X1  g09762(.A0(new_n8659_), .A1(new_n3250_), .B0(new_n6920_), .B1(new_n3144_), .Y(new_n9827_));
  AOI21X1  g09763(.A0(new_n8580_), .A1(new_n3146_), .B0(new_n9827_), .Y(new_n9828_));
  OAI21X1  g09764(.A0(new_n8611_), .A1(new_n3098_), .B0(new_n9828_), .Y(new_n9829_));
  XOR2X1   g09765(.A(new_n9829_), .B(new_n1920_), .Y(new_n9830_));
  NOR2X1   g09766(.A(new_n9830_), .B(new_n9826_), .Y(new_n9831_));
  INVX1    g09767(.A(new_n9831_), .Y(new_n9832_));
  AOI22X1  g09768(.A0(new_n6925_), .A1(new_n2875_), .B0(new_n6923_), .B1(new_n3099_), .Y(new_n9833_));
  OAI21X1  g09769(.A0(new_n6920_), .A1(new_n3152_), .B0(new_n9833_), .Y(new_n9834_));
  AOI21X1  g09770(.A0(new_n8628_), .A1(new_n2876_), .B0(new_n9834_), .Y(new_n9835_));
  XOR2X1   g09771(.A(new_n9835_), .B(\a[20] ), .Y(new_n9836_));
  INVX1    g09772(.A(new_n9836_), .Y(new_n9837_));
  XOR2X1   g09773(.A(new_n9626_), .B(new_n9625_), .Y(new_n9838_));
  AND2X1   g09774(.A(new_n9838_), .B(new_n9837_), .Y(new_n9839_));
  INVX1    g09775(.A(new_n9839_), .Y(new_n9840_));
  XOR2X1   g09776(.A(new_n9838_), .B(new_n9836_), .Y(new_n9841_));
  XOR2X1   g09777(.A(new_n9624_), .B(new_n9619_), .Y(new_n9842_));
  OAI22X1  g09778(.A0(new_n6929_), .A1(new_n3250_), .B0(new_n8683_), .B1(new_n3144_), .Y(new_n9843_));
  AOI21X1  g09779(.A0(new_n6923_), .A1(new_n3146_), .B0(new_n9843_), .Y(new_n9844_));
  OAI21X1  g09780(.A0(new_n8662_), .A1(new_n3098_), .B0(new_n9844_), .Y(new_n9845_));
  XOR2X1   g09781(.A(new_n9845_), .B(new_n1920_), .Y(new_n9846_));
  NOR2X1   g09782(.A(new_n9846_), .B(new_n9842_), .Y(new_n9847_));
  AOI22X1  g09783(.A0(new_n6932_), .A1(new_n2875_), .B0(new_n6927_), .B1(new_n3099_), .Y(new_n9848_));
  OAI21X1  g09784(.A0(new_n8683_), .A1(new_n3152_), .B0(new_n9848_), .Y(new_n9849_));
  AOI21X1  g09785(.A0(new_n8682_), .A1(new_n2876_), .B0(new_n9849_), .Y(new_n9850_));
  XOR2X1   g09786(.A(new_n9850_), .B(\a[20] ), .Y(new_n9851_));
  NOR3X1   g09787(.A(new_n9613_), .B(new_n9612_), .C(new_n70_), .Y(new_n9852_));
  XOR2X1   g09788(.A(new_n9616_), .B(\a[23] ), .Y(new_n9853_));
  NOR2X1   g09789(.A(new_n9853_), .B(new_n9852_), .Y(new_n9854_));
  NOR3X1   g09790(.A(new_n9854_), .B(new_n9851_), .C(new_n9617_), .Y(new_n9855_));
  XOR2X1   g09791(.A(new_n9853_), .B(new_n9852_), .Y(new_n9856_));
  XOR2X1   g09792(.A(new_n9856_), .B(new_n9851_), .Y(new_n9857_));
  NOR2X1   g09793(.A(new_n9613_), .B(new_n70_), .Y(new_n9858_));
  XOR2X1   g09794(.A(new_n9858_), .B(new_n9612_), .Y(new_n9859_));
  OAI22X1  g09795(.A0(new_n8757_), .A1(new_n3250_), .B0(new_n6930_), .B1(new_n3144_), .Y(new_n9860_));
  AOI21X1  g09796(.A0(new_n6927_), .A1(new_n3146_), .B0(new_n9860_), .Y(new_n9861_));
  OAI21X1  g09797(.A0(new_n8705_), .A1(new_n3098_), .B0(new_n9861_), .Y(new_n9862_));
  XOR2X1   g09798(.A(new_n9862_), .B(new_n1920_), .Y(new_n9863_));
  NOR2X1   g09799(.A(new_n9863_), .B(new_n9859_), .Y(new_n9864_));
  OAI22X1  g09800(.A0(new_n6936_), .A1(new_n3144_), .B0(new_n8752_), .B1(new_n3152_), .Y(new_n9865_));
  AOI21X1  g09801(.A0(new_n8751_), .A1(new_n2876_), .B0(new_n9865_), .Y(new_n9866_));
  NOR2X1   g09802(.A(new_n6936_), .B(new_n2869_), .Y(new_n9867_));
  INVX1    g09803(.A(new_n9867_), .Y(new_n9868_));
  NAND3X1  g09804(.A(new_n9868_), .B(new_n9866_), .C(\a[20] ), .Y(new_n9869_));
  OAI22X1  g09805(.A0(new_n6936_), .A1(new_n3250_), .B0(new_n8752_), .B1(new_n3144_), .Y(new_n9870_));
  AOI21X1  g09806(.A0(new_n6933_), .A1(new_n3146_), .B0(new_n9870_), .Y(new_n9871_));
  OAI21X1  g09807(.A0(new_n8759_), .A1(new_n3098_), .B0(new_n9871_), .Y(new_n9872_));
  XOR2X1   g09808(.A(new_n9872_), .B(new_n1920_), .Y(new_n9873_));
  OR4X1    g09809(.A(new_n9873_), .B(new_n9869_), .C(new_n6936_), .D(new_n2655_), .Y(new_n9874_));
  XOR2X1   g09810(.A(new_n9866_), .B(\a[20] ), .Y(new_n9875_));
  OR4X1    g09811(.A(new_n9872_), .B(new_n9867_), .C(new_n9875_), .D(new_n1920_), .Y(new_n9876_));
  XOR2X1   g09812(.A(new_n9876_), .B(new_n9613_), .Y(new_n9877_));
  AOI22X1  g09813(.A0(new_n6935_), .A1(new_n2875_), .B0(new_n6933_), .B1(new_n3099_), .Y(new_n9878_));
  OAI21X1  g09814(.A0(new_n6930_), .A1(new_n3152_), .B0(new_n9878_), .Y(new_n9879_));
  AOI21X1  g09815(.A0(new_n8717_), .A1(new_n2876_), .B0(new_n9879_), .Y(new_n9880_));
  XOR2X1   g09816(.A(new_n9880_), .B(\a[20] ), .Y(new_n9881_));
  OAI21X1  g09817(.A0(new_n9881_), .A1(new_n9877_), .B0(new_n9874_), .Y(new_n9882_));
  XOR2X1   g09818(.A(new_n9863_), .B(new_n9859_), .Y(new_n9883_));
  AOI21X1  g09819(.A0(new_n9883_), .A1(new_n9882_), .B0(new_n9864_), .Y(new_n9884_));
  NOR2X1   g09820(.A(new_n9884_), .B(new_n9857_), .Y(new_n9885_));
  OR2X1    g09821(.A(new_n9885_), .B(new_n9855_), .Y(new_n9886_));
  XOR2X1   g09822(.A(new_n9846_), .B(new_n9842_), .Y(new_n9887_));
  AOI21X1  g09823(.A0(new_n9887_), .A1(new_n9886_), .B0(new_n9847_), .Y(new_n9888_));
  OAI21X1  g09824(.A0(new_n9888_), .A1(new_n9841_), .B0(new_n9840_), .Y(new_n9889_));
  INVX1    g09825(.A(new_n9889_), .Y(new_n9890_));
  XOR2X1   g09826(.A(new_n9830_), .B(new_n9825_), .Y(new_n9891_));
  OAI21X1  g09827(.A0(new_n9891_), .A1(new_n9890_), .B0(new_n9832_), .Y(new_n9892_));
  INVX1    g09828(.A(new_n9892_), .Y(new_n9893_));
  XOR2X1   g09829(.A(new_n9823_), .B(new_n9818_), .Y(new_n9894_));
  OAI21X1  g09830(.A0(new_n9894_), .A1(new_n9893_), .B0(new_n9824_), .Y(new_n9895_));
  XOR2X1   g09831(.A(new_n9816_), .B(new_n9812_), .Y(new_n9896_));
  AOI21X1  g09832(.A0(new_n9896_), .A1(new_n9895_), .B0(new_n9817_), .Y(new_n9897_));
  OAI21X1  g09833(.A0(new_n9897_), .A1(new_n9810_), .B0(new_n9808_), .Y(new_n9898_));
  AOI21X1  g09834(.A0(new_n9898_), .A1(new_n9802_), .B0(new_n9800_), .Y(new_n9899_));
  XOR2X1   g09835(.A(new_n9791_), .B(new_n9786_), .Y(new_n9900_));
  OAI21X1  g09836(.A0(new_n9900_), .A1(new_n9899_), .B0(new_n9793_), .Y(new_n9901_));
  INVX1    g09837(.A(new_n9901_), .Y(new_n9902_));
  XOR2X1   g09838(.A(new_n9783_), .B(new_n9778_), .Y(new_n9903_));
  OAI21X1  g09839(.A0(new_n9903_), .A1(new_n9902_), .B0(new_n9785_), .Y(new_n9904_));
  INVX1    g09840(.A(new_n9904_), .Y(new_n9905_));
  XOR2X1   g09841(.A(new_n9774_), .B(new_n1920_), .Y(new_n9906_));
  XOR2X1   g09842(.A(new_n9906_), .B(new_n9771_), .Y(new_n9907_));
  OAI21X1  g09843(.A0(new_n9907_), .A1(new_n9905_), .B0(new_n9777_), .Y(new_n9908_));
  INVX1    g09844(.A(new_n9908_), .Y(new_n9909_));
  XOR2X1   g09845(.A(new_n9767_), .B(new_n1920_), .Y(new_n9910_));
  XOR2X1   g09846(.A(new_n9910_), .B(new_n9764_), .Y(new_n9911_));
  OAI21X1  g09847(.A0(new_n9911_), .A1(new_n9909_), .B0(new_n9770_), .Y(new_n9912_));
  INVX1    g09848(.A(new_n9912_), .Y(new_n9913_));
  XOR2X1   g09849(.A(new_n9760_), .B(\a[20] ), .Y(new_n9914_));
  XOR2X1   g09850(.A(new_n9914_), .B(new_n9757_), .Y(new_n9915_));
  OAI21X1  g09851(.A0(new_n9915_), .A1(new_n9913_), .B0(new_n9763_), .Y(new_n9916_));
  INVX1    g09852(.A(new_n9916_), .Y(new_n9917_));
  XOR2X1   g09853(.A(new_n9753_), .B(new_n1920_), .Y(new_n9918_));
  XOR2X1   g09854(.A(new_n9918_), .B(new_n9750_), .Y(new_n9919_));
  OAI21X1  g09855(.A0(new_n9919_), .A1(new_n9917_), .B0(new_n9756_), .Y(new_n9920_));
  XOR2X1   g09856(.A(new_n9747_), .B(new_n1920_), .Y(new_n9921_));
  XOR2X1   g09857(.A(new_n9921_), .B(new_n9743_), .Y(new_n9922_));
  INVX1    g09858(.A(new_n9922_), .Y(new_n9923_));
  AOI21X1  g09859(.A0(new_n9923_), .A1(new_n9920_), .B0(new_n9749_), .Y(new_n9924_));
  XOR2X1   g09860(.A(new_n9741_), .B(new_n1920_), .Y(new_n9925_));
  XOR2X1   g09861(.A(new_n9925_), .B(new_n9737_), .Y(new_n9926_));
  NOR2X1   g09862(.A(new_n9926_), .B(new_n9924_), .Y(new_n9927_));
  AOI21X1  g09863(.A0(new_n9742_), .A1(new_n9737_), .B0(new_n9927_), .Y(new_n9928_));
  XOR2X1   g09864(.A(new_n9734_), .B(new_n9730_), .Y(new_n9929_));
  OAI21X1  g09865(.A0(new_n9929_), .A1(new_n9928_), .B0(new_n9736_), .Y(new_n9930_));
  XOR2X1   g09866(.A(new_n9728_), .B(new_n9724_), .Y(new_n9931_));
  AOI21X1  g09867(.A0(new_n9931_), .A1(new_n9930_), .B0(new_n9729_), .Y(new_n9932_));
  AOI21X1  g09868(.A0(new_n9721_), .A1(new_n9720_), .B0(new_n9932_), .Y(new_n9933_));
  NAND3X1  g09869(.A(new_n9932_), .B(new_n9721_), .C(new_n9720_), .Y(new_n9934_));
  AOI22X1  g09870(.A0(new_n6822_), .A1(new_n3232_), .B0(new_n6820_), .B1(new_n3390_), .Y(new_n9935_));
  OAI21X1  g09871(.A0(new_n7418_), .A1(new_n3545_), .B0(new_n9935_), .Y(new_n9936_));
  AOI21X1  g09872(.A0(new_n7417_), .A1(new_n3234_), .B0(new_n9936_), .Y(new_n9937_));
  XOR2X1   g09873(.A(new_n9937_), .B(\a[17] ), .Y(new_n9938_));
  INVX1    g09874(.A(new_n9938_), .Y(new_n9939_));
  AOI21X1  g09875(.A0(new_n9939_), .A1(new_n9934_), .B0(new_n9933_), .Y(new_n9940_));
  AOI21X1  g09876(.A0(new_n9719_), .A1(new_n9717_), .B0(new_n9940_), .Y(new_n9941_));
  NAND3X1  g09877(.A(new_n9940_), .B(new_n9719_), .C(new_n9717_), .Y(new_n9942_));
  AOI22X1  g09878(.A0(new_n7364_), .A1(new_n3908_), .B0(new_n7044_), .B1(new_n3628_), .Y(new_n9943_));
  OAI21X1  g09879(.A0(new_n7504_), .A1(new_n3983_), .B0(new_n9943_), .Y(new_n9944_));
  AOI21X1  g09880(.A0(new_n7552_), .A1(new_n3624_), .B0(new_n9944_), .Y(new_n9945_));
  XOR2X1   g09881(.A(new_n9945_), .B(\a[14] ), .Y(new_n9946_));
  INVX1    g09882(.A(new_n9946_), .Y(new_n9947_));
  AOI21X1  g09883(.A0(new_n9947_), .A1(new_n9942_), .B0(new_n9941_), .Y(new_n9948_));
  NOR2X1   g09884(.A(new_n9948_), .B(new_n9707_), .Y(new_n9949_));
  XOR2X1   g09885(.A(new_n9948_), .B(new_n9707_), .Y(new_n9950_));
  AOI22X1  g09886(.A0(new_n7558_), .A1(new_n4247_), .B0(new_n7529_), .B1(new_n4078_), .Y(new_n9951_));
  OAI21X1  g09887(.A0(new_n7623_), .A1(new_n4427_), .B0(new_n9951_), .Y(new_n9952_));
  AOI21X1  g09888(.A0(new_n7622_), .A1(new_n4080_), .B0(new_n9952_), .Y(new_n9953_));
  XOR2X1   g09889(.A(new_n9953_), .B(new_n2911_), .Y(new_n9954_));
  AOI21X1  g09890(.A0(new_n9954_), .A1(new_n9950_), .B0(new_n9949_), .Y(new_n9955_));
  NOR2X1   g09891(.A(new_n9955_), .B(new_n9705_), .Y(new_n9956_));
  OR2X1    g09892(.A(new_n9956_), .B(new_n9703_), .Y(new_n9957_));
  NOR2X1   g09893(.A(new_n9956_), .B(new_n9703_), .Y(new_n9958_));
  XOR2X1   g09894(.A(new_n9958_), .B(new_n9695_), .Y(new_n9959_));
  AOI22X1  g09895(.A0(new_n7657_), .A1(new_n4635_), .B0(new_n7341_), .B1(new_n5097_), .Y(new_n9960_));
  OAI21X1  g09896(.A0(new_n7644_), .A1(new_n4869_), .B0(new_n9960_), .Y(new_n9961_));
  AOI21X1  g09897(.A0(new_n7656_), .A1(new_n4637_), .B0(new_n9961_), .Y(new_n9962_));
  XOR2X1   g09898(.A(new_n9962_), .B(\a[8] ), .Y(new_n9963_));
  NOR2X1   g09899(.A(new_n9963_), .B(new_n9959_), .Y(new_n9964_));
  AOI21X1  g09900(.A0(new_n9957_), .A1(new_n9695_), .B0(new_n9964_), .Y(new_n9965_));
  OR2X1    g09901(.A(new_n9965_), .B(new_n9694_), .Y(new_n9966_));
  XOR2X1   g09902(.A(new_n9687_), .B(new_n9686_), .Y(new_n9967_));
  XOR2X1   g09903(.A(new_n9965_), .B(new_n9967_), .Y(new_n9968_));
  XOR2X1   g09904(.A(new_n9957_), .B(new_n9695_), .Y(new_n9969_));
  XOR2X1   g09905(.A(new_n9963_), .B(new_n9969_), .Y(new_n9970_));
  XOR2X1   g09906(.A(new_n9953_), .B(\a[11] ), .Y(new_n9971_));
  XOR2X1   g09907(.A(new_n9971_), .B(new_n9950_), .Y(new_n9972_));
  NOR3X1   g09908(.A(new_n9663_), .B(new_n9718_), .C(new_n9657_), .Y(new_n9973_));
  AOI21X1  g09909(.A0(new_n9658_), .A1(new_n9716_), .B0(new_n9662_), .Y(new_n9974_));
  NOR3X1   g09910(.A(new_n9655_), .B(new_n9714_), .C(new_n9649_), .Y(new_n9975_));
  AOI21X1  g09911(.A0(new_n9650_), .A1(new_n9713_), .B0(new_n9654_), .Y(new_n9976_));
  INVX1    g09912(.A(new_n9932_), .Y(new_n9977_));
  OAI21X1  g09913(.A0(new_n9976_), .A1(new_n9975_), .B0(new_n9977_), .Y(new_n9978_));
  NOR3X1   g09914(.A(new_n9977_), .B(new_n9976_), .C(new_n9975_), .Y(new_n9979_));
  OAI21X1  g09915(.A0(new_n9938_), .A1(new_n9979_), .B0(new_n9978_), .Y(new_n9980_));
  OAI21X1  g09916(.A0(new_n9974_), .A1(new_n9973_), .B0(new_n9980_), .Y(new_n9981_));
  NAND3X1  g09917(.A(new_n9946_), .B(new_n9942_), .C(new_n9981_), .Y(new_n9982_));
  NOR3X1   g09918(.A(new_n9980_), .B(new_n9974_), .C(new_n9973_), .Y(new_n9983_));
  OAI21X1  g09919(.A0(new_n9983_), .A1(new_n9941_), .B0(new_n9947_), .Y(new_n9984_));
  NAND3X1  g09920(.A(new_n9938_), .B(new_n9934_), .C(new_n9978_), .Y(new_n9985_));
  OAI21X1  g09921(.A0(new_n9979_), .A1(new_n9933_), .B0(new_n9939_), .Y(new_n9986_));
  AOI22X1  g09922(.A0(new_n6882_), .A1(new_n3232_), .B0(new_n6822_), .B1(new_n3390_), .Y(new_n9987_));
  OAI21X1  g09923(.A0(new_n7671_), .A1(new_n3545_), .B0(new_n9987_), .Y(new_n9988_));
  AOI21X1  g09924(.A0(new_n7670_), .A1(new_n3234_), .B0(new_n9988_), .Y(new_n9989_));
  XOR2X1   g09925(.A(new_n9989_), .B(\a[17] ), .Y(new_n9990_));
  INVX1    g09926(.A(new_n9990_), .Y(new_n9991_));
  XOR2X1   g09927(.A(new_n9931_), .B(new_n9930_), .Y(new_n9992_));
  AND2X1   g09928(.A(new_n9992_), .B(new_n9991_), .Y(new_n9993_));
  XOR2X1   g09929(.A(new_n9992_), .B(new_n9991_), .Y(new_n9994_));
  AOI22X1  g09930(.A0(new_n6885_), .A1(new_n3232_), .B0(new_n6882_), .B1(new_n3390_), .Y(new_n9995_));
  OAI21X1  g09931(.A0(new_n7472_), .A1(new_n3545_), .B0(new_n9995_), .Y(new_n9996_));
  AOI21X1  g09932(.A0(new_n7471_), .A1(new_n3234_), .B0(new_n9996_), .Y(new_n9997_));
  XOR2X1   g09933(.A(new_n9997_), .B(\a[17] ), .Y(new_n9998_));
  INVX1    g09934(.A(new_n9929_), .Y(new_n9999_));
  XOR2X1   g09935(.A(new_n9999_), .B(new_n9928_), .Y(new_n10000_));
  OR2X1    g09936(.A(new_n10000_), .B(new_n9998_), .Y(new_n10001_));
  XOR2X1   g09937(.A(new_n10000_), .B(new_n9998_), .Y(new_n10002_));
  AOI22X1  g09938(.A0(new_n6887_), .A1(new_n3232_), .B0(new_n6885_), .B1(new_n3390_), .Y(new_n10003_));
  OAI21X1  g09939(.A0(new_n6884_), .A1(new_n3545_), .B0(new_n10003_), .Y(new_n10004_));
  AOI21X1  g09940(.A0(new_n7771_), .A1(new_n3234_), .B0(new_n10004_), .Y(new_n10005_));
  XOR2X1   g09941(.A(new_n10005_), .B(\a[17] ), .Y(new_n10006_));
  INVX1    g09942(.A(new_n9926_), .Y(new_n10007_));
  XOR2X1   g09943(.A(new_n10007_), .B(new_n9924_), .Y(new_n10008_));
  NOR2X1   g09944(.A(new_n10008_), .B(new_n10006_), .Y(new_n10009_));
  XOR2X1   g09945(.A(new_n10008_), .B(new_n10006_), .Y(new_n10010_));
  INVX1    g09946(.A(new_n10010_), .Y(new_n10011_));
  AOI22X1  g09947(.A0(new_n6890_), .A1(new_n3232_), .B0(new_n6887_), .B1(new_n3390_), .Y(new_n10012_));
  OAI21X1  g09948(.A0(new_n6886_), .A1(new_n3545_), .B0(new_n10012_), .Y(new_n10013_));
  AOI21X1  g09949(.A0(new_n7762_), .A1(new_n3234_), .B0(new_n10013_), .Y(new_n10014_));
  XOR2X1   g09950(.A(new_n10014_), .B(\a[17] ), .Y(new_n10015_));
  XOR2X1   g09951(.A(new_n9922_), .B(new_n9920_), .Y(new_n10016_));
  NOR2X1   g09952(.A(new_n10016_), .B(new_n10015_), .Y(new_n10017_));
  XOR2X1   g09953(.A(new_n10016_), .B(new_n10015_), .Y(new_n10018_));
  AOI22X1  g09954(.A0(new_n6892_), .A1(new_n3232_), .B0(new_n6890_), .B1(new_n3390_), .Y(new_n10019_));
  OAI21X1  g09955(.A0(new_n7878_), .A1(new_n3545_), .B0(new_n10019_), .Y(new_n10020_));
  AOI21X1  g09956(.A0(new_n7877_), .A1(new_n3234_), .B0(new_n10020_), .Y(new_n10021_));
  XOR2X1   g09957(.A(new_n10021_), .B(\a[17] ), .Y(new_n10022_));
  XOR2X1   g09958(.A(new_n9919_), .B(new_n9916_), .Y(new_n10023_));
  NOR2X1   g09959(.A(new_n10023_), .B(new_n10022_), .Y(new_n10024_));
  XOR2X1   g09960(.A(new_n10023_), .B(new_n10022_), .Y(new_n10025_));
  AOI22X1  g09961(.A0(new_n6894_), .A1(new_n3232_), .B0(new_n6892_), .B1(new_n3390_), .Y(new_n10026_));
  OAI21X1  g09962(.A0(new_n7885_), .A1(new_n3545_), .B0(new_n10026_), .Y(new_n10027_));
  AOI21X1  g09963(.A0(new_n7884_), .A1(new_n3234_), .B0(new_n10027_), .Y(new_n10028_));
  XOR2X1   g09964(.A(new_n10028_), .B(\a[17] ), .Y(new_n10029_));
  XOR2X1   g09965(.A(new_n9915_), .B(new_n9912_), .Y(new_n10030_));
  NOR2X1   g09966(.A(new_n10030_), .B(new_n10029_), .Y(new_n10031_));
  XOR2X1   g09967(.A(new_n10030_), .B(new_n10029_), .Y(new_n10032_));
  AOI22X1  g09968(.A0(new_n6897_), .A1(new_n3232_), .B0(new_n6894_), .B1(new_n3390_), .Y(new_n10033_));
  OAI21X1  g09969(.A0(new_n8075_), .A1(new_n3545_), .B0(new_n10033_), .Y(new_n10034_));
  AOI21X1  g09970(.A0(new_n8074_), .A1(new_n3234_), .B0(new_n10034_), .Y(new_n10035_));
  XOR2X1   g09971(.A(new_n10035_), .B(\a[17] ), .Y(new_n10036_));
  XOR2X1   g09972(.A(new_n9911_), .B(new_n9908_), .Y(new_n10037_));
  NOR2X1   g09973(.A(new_n10037_), .B(new_n10036_), .Y(new_n10038_));
  XOR2X1   g09974(.A(new_n10037_), .B(new_n10036_), .Y(new_n10039_));
  AOI22X1  g09975(.A0(new_n6899_), .A1(new_n3232_), .B0(new_n6897_), .B1(new_n3390_), .Y(new_n10040_));
  OAI21X1  g09976(.A0(new_n6896_), .A1(new_n3545_), .B0(new_n10040_), .Y(new_n10041_));
  AOI21X1  g09977(.A0(new_n7953_), .A1(new_n3234_), .B0(new_n10041_), .Y(new_n10042_));
  XOR2X1   g09978(.A(new_n10042_), .B(\a[17] ), .Y(new_n10043_));
  XOR2X1   g09979(.A(new_n9907_), .B(new_n9904_), .Y(new_n10044_));
  NOR2X1   g09980(.A(new_n10044_), .B(new_n10043_), .Y(new_n10045_));
  XOR2X1   g09981(.A(new_n10044_), .B(new_n10043_), .Y(new_n10046_));
  AOI22X1  g09982(.A0(new_n6902_), .A1(new_n3232_), .B0(new_n6899_), .B1(new_n3390_), .Y(new_n10047_));
  OAI21X1  g09983(.A0(new_n6898_), .A1(new_n3545_), .B0(new_n10047_), .Y(new_n10048_));
  AOI21X1  g09984(.A0(new_n8215_), .A1(new_n3234_), .B0(new_n10048_), .Y(new_n10049_));
  XOR2X1   g09985(.A(new_n10049_), .B(\a[17] ), .Y(new_n10050_));
  XOR2X1   g09986(.A(new_n9903_), .B(new_n9901_), .Y(new_n10051_));
  NOR2X1   g09987(.A(new_n10051_), .B(new_n10050_), .Y(new_n10052_));
  XOR2X1   g09988(.A(new_n10051_), .B(new_n10050_), .Y(new_n10053_));
  INVX1    g09989(.A(new_n10053_), .Y(new_n10054_));
  AOI22X1  g09990(.A0(new_n6904_), .A1(new_n3232_), .B0(new_n6902_), .B1(new_n3390_), .Y(new_n10055_));
  OAI21X1  g09991(.A0(new_n8295_), .A1(new_n3545_), .B0(new_n10055_), .Y(new_n10056_));
  AOI21X1  g09992(.A0(new_n8883_), .A1(new_n3234_), .B0(new_n10056_), .Y(new_n10057_));
  XOR2X1   g09993(.A(new_n10057_), .B(\a[17] ), .Y(new_n10058_));
  INVX1    g09994(.A(new_n9900_), .Y(new_n10059_));
  XOR2X1   g09995(.A(new_n10059_), .B(new_n9899_), .Y(new_n10060_));
  OR2X1    g09996(.A(new_n10060_), .B(new_n10058_), .Y(new_n10061_));
  XOR2X1   g09997(.A(new_n10060_), .B(new_n10058_), .Y(new_n10062_));
  INVX1    g09998(.A(new_n10062_), .Y(new_n10063_));
  XOR2X1   g09999(.A(new_n9898_), .B(new_n9801_), .Y(new_n10064_));
  OAI22X1  g10000(.A0(new_n6964_), .A1(new_n3231_), .B0(new_n8200_), .B1(new_n3389_), .Y(new_n10065_));
  AOI21X1  g10001(.A0(new_n6902_), .A1(new_n3546_), .B0(new_n10065_), .Y(new_n10066_));
  OAI21X1  g10002(.A0(new_n8203_), .A1(new_n3388_), .B0(new_n10066_), .Y(new_n10067_));
  XOR2X1   g10003(.A(new_n10067_), .B(new_n2445_), .Y(new_n10068_));
  NOR2X1   g10004(.A(new_n10068_), .B(new_n10064_), .Y(new_n10069_));
  XOR2X1   g10005(.A(new_n9897_), .B(new_n9810_), .Y(new_n10070_));
  INVX1    g10006(.A(new_n10070_), .Y(new_n10071_));
  OAI22X1  g10007(.A0(new_n6960_), .A1(new_n3231_), .B0(new_n6964_), .B1(new_n3389_), .Y(new_n10072_));
  AOI21X1  g10008(.A0(new_n6904_), .A1(new_n3546_), .B0(new_n10072_), .Y(new_n10073_));
  OAI21X1  g10009(.A0(new_n8364_), .A1(new_n3388_), .B0(new_n10073_), .Y(new_n10074_));
  XOR2X1   g10010(.A(new_n10074_), .B(new_n2445_), .Y(new_n10075_));
  OR2X1    g10011(.A(new_n10075_), .B(new_n10071_), .Y(new_n10076_));
  AOI22X1  g10012(.A0(new_n6911_), .A1(new_n3232_), .B0(new_n6909_), .B1(new_n3390_), .Y(new_n10077_));
  OAI21X1  g10013(.A0(new_n6964_), .A1(new_n3545_), .B0(new_n10077_), .Y(new_n10078_));
  AOI21X1  g10014(.A0(new_n8541_), .A1(new_n3234_), .B0(new_n10078_), .Y(new_n10079_));
  XOR2X1   g10015(.A(new_n10079_), .B(\a[17] ), .Y(new_n10080_));
  INVX1    g10016(.A(new_n10080_), .Y(new_n10081_));
  XOR2X1   g10017(.A(new_n9896_), .B(new_n9895_), .Y(new_n10082_));
  AND2X1   g10018(.A(new_n10082_), .B(new_n10081_), .Y(new_n10083_));
  XOR2X1   g10019(.A(new_n10082_), .B(new_n10080_), .Y(new_n10084_));
  AOI22X1  g10020(.A0(new_n6913_), .A1(new_n3232_), .B0(new_n6911_), .B1(new_n3390_), .Y(new_n10085_));
  OAI21X1  g10021(.A0(new_n6960_), .A1(new_n3545_), .B0(new_n10085_), .Y(new_n10086_));
  AOI21X1  g10022(.A0(new_n8553_), .A1(new_n3234_), .B0(new_n10086_), .Y(new_n10087_));
  XOR2X1   g10023(.A(new_n10087_), .B(\a[17] ), .Y(new_n10088_));
  XOR2X1   g10024(.A(new_n9894_), .B(new_n9892_), .Y(new_n10089_));
  NOR2X1   g10025(.A(new_n10089_), .B(new_n10088_), .Y(new_n10090_));
  XOR2X1   g10026(.A(new_n10089_), .B(new_n10088_), .Y(new_n10091_));
  AOI22X1  g10027(.A0(new_n6915_), .A1(new_n3232_), .B0(new_n6913_), .B1(new_n3390_), .Y(new_n10092_));
  OAI21X1  g10028(.A0(new_n8349_), .A1(new_n3545_), .B0(new_n10092_), .Y(new_n10093_));
  AOI21X1  g10029(.A0(new_n8348_), .A1(new_n3234_), .B0(new_n10093_), .Y(new_n10094_));
  XOR2X1   g10030(.A(new_n10094_), .B(\a[17] ), .Y(new_n10095_));
  XOR2X1   g10031(.A(new_n9891_), .B(new_n9889_), .Y(new_n10096_));
  OR2X1    g10032(.A(new_n10096_), .B(new_n10095_), .Y(new_n10097_));
  XOR2X1   g10033(.A(new_n10096_), .B(new_n10095_), .Y(new_n10098_));
  INVX1    g10034(.A(new_n10098_), .Y(new_n10099_));
  INVX1    g10035(.A(new_n9841_), .Y(new_n10100_));
  XOR2X1   g10036(.A(new_n9888_), .B(new_n10100_), .Y(new_n10101_));
  OAI22X1  g10037(.A0(new_n6918_), .A1(new_n3231_), .B0(new_n6917_), .B1(new_n3389_), .Y(new_n10102_));
  AOI21X1  g10038(.A0(new_n6913_), .A1(new_n3546_), .B0(new_n10102_), .Y(new_n10103_));
  OAI21X1  g10039(.A0(new_n8577_), .A1(new_n3388_), .B0(new_n10103_), .Y(new_n10104_));
  XOR2X1   g10040(.A(new_n10104_), .B(new_n2445_), .Y(new_n10105_));
  NOR2X1   g10041(.A(new_n10105_), .B(new_n10101_), .Y(new_n10106_));
  XOR2X1   g10042(.A(new_n9887_), .B(new_n9886_), .Y(new_n10107_));
  INVX1    g10043(.A(new_n10107_), .Y(new_n10108_));
  OAI22X1  g10044(.A0(new_n6920_), .A1(new_n3231_), .B0(new_n6918_), .B1(new_n3389_), .Y(new_n10109_));
  AOI21X1  g10045(.A0(new_n6915_), .A1(new_n3546_), .B0(new_n10109_), .Y(new_n10110_));
  OAI21X1  g10046(.A0(new_n9093_), .A1(new_n3388_), .B0(new_n10110_), .Y(new_n10111_));
  XOR2X1   g10047(.A(new_n10111_), .B(new_n2445_), .Y(new_n10112_));
  OR2X1    g10048(.A(new_n10112_), .B(new_n10108_), .Y(new_n10113_));
  XOR2X1   g10049(.A(new_n9884_), .B(new_n9857_), .Y(new_n10114_));
  INVX1    g10050(.A(new_n10114_), .Y(new_n10115_));
  OAI22X1  g10051(.A0(new_n8659_), .A1(new_n3231_), .B0(new_n6920_), .B1(new_n3389_), .Y(new_n10116_));
  AOI21X1  g10052(.A0(new_n8580_), .A1(new_n3546_), .B0(new_n10116_), .Y(new_n10117_));
  OAI21X1  g10053(.A0(new_n8611_), .A1(new_n3388_), .B0(new_n10117_), .Y(new_n10118_));
  XOR2X1   g10054(.A(new_n10118_), .B(new_n2445_), .Y(new_n10119_));
  NOR2X1   g10055(.A(new_n10119_), .B(new_n10115_), .Y(new_n10120_));
  INVX1    g10056(.A(new_n10120_), .Y(new_n10121_));
  AOI22X1  g10057(.A0(new_n6925_), .A1(new_n3232_), .B0(new_n6923_), .B1(new_n3390_), .Y(new_n10122_));
  OAI21X1  g10058(.A0(new_n6920_), .A1(new_n3545_), .B0(new_n10122_), .Y(new_n10123_));
  AOI21X1  g10059(.A0(new_n8628_), .A1(new_n3234_), .B0(new_n10123_), .Y(new_n10124_));
  XOR2X1   g10060(.A(new_n10124_), .B(\a[17] ), .Y(new_n10125_));
  INVX1    g10061(.A(new_n10125_), .Y(new_n10126_));
  XOR2X1   g10062(.A(new_n9883_), .B(new_n9882_), .Y(new_n10127_));
  AND2X1   g10063(.A(new_n10127_), .B(new_n10126_), .Y(new_n10128_));
  INVX1    g10064(.A(new_n10128_), .Y(new_n10129_));
  XOR2X1   g10065(.A(new_n10127_), .B(new_n10125_), .Y(new_n10130_));
  XOR2X1   g10066(.A(new_n9880_), .B(new_n1920_), .Y(new_n10131_));
  XOR2X1   g10067(.A(new_n10131_), .B(new_n9877_), .Y(new_n10132_));
  OAI22X1  g10068(.A0(new_n6929_), .A1(new_n3231_), .B0(new_n8683_), .B1(new_n3389_), .Y(new_n10133_));
  AOI21X1  g10069(.A0(new_n6923_), .A1(new_n3546_), .B0(new_n10133_), .Y(new_n10134_));
  OAI21X1  g10070(.A0(new_n8662_), .A1(new_n3388_), .B0(new_n10134_), .Y(new_n10135_));
  XOR2X1   g10071(.A(new_n10135_), .B(new_n2445_), .Y(new_n10136_));
  NOR2X1   g10072(.A(new_n10136_), .B(new_n10132_), .Y(new_n10137_));
  AOI22X1  g10073(.A0(new_n6932_), .A1(new_n3232_), .B0(new_n6927_), .B1(new_n3390_), .Y(new_n10138_));
  OAI21X1  g10074(.A0(new_n8683_), .A1(new_n3545_), .B0(new_n10138_), .Y(new_n10139_));
  AOI21X1  g10075(.A0(new_n8682_), .A1(new_n3234_), .B0(new_n10139_), .Y(new_n10140_));
  XOR2X1   g10076(.A(new_n10140_), .B(\a[17] ), .Y(new_n10141_));
  INVX1    g10077(.A(new_n10141_), .Y(new_n10142_));
  XOR2X1   g10078(.A(new_n9873_), .B(new_n9869_), .Y(new_n10143_));
  AND2X1   g10079(.A(new_n10143_), .B(new_n10142_), .Y(new_n10144_));
  XOR2X1   g10080(.A(new_n10143_), .B(new_n10141_), .Y(new_n10145_));
  NOR2X1   g10081(.A(new_n9867_), .B(new_n1920_), .Y(new_n10146_));
  XOR2X1   g10082(.A(new_n10146_), .B(new_n9875_), .Y(new_n10147_));
  OAI22X1  g10083(.A0(new_n8757_), .A1(new_n3231_), .B0(new_n6930_), .B1(new_n3389_), .Y(new_n10148_));
  AOI21X1  g10084(.A0(new_n6927_), .A1(new_n3546_), .B0(new_n10148_), .Y(new_n10149_));
  OAI21X1  g10085(.A0(new_n8705_), .A1(new_n3388_), .B0(new_n10149_), .Y(new_n10150_));
  XOR2X1   g10086(.A(new_n10150_), .B(new_n2445_), .Y(new_n10151_));
  NOR2X1   g10087(.A(new_n10151_), .B(new_n10147_), .Y(new_n10152_));
  OAI22X1  g10088(.A0(new_n6936_), .A1(new_n3389_), .B0(new_n8752_), .B1(new_n3545_), .Y(new_n10153_));
  AOI21X1  g10089(.A0(new_n8751_), .A1(new_n3234_), .B0(new_n10153_), .Y(new_n10154_));
  XOR2X1   g10090(.A(new_n10154_), .B(\a[17] ), .Y(new_n10155_));
  NOR2X1   g10091(.A(new_n6936_), .B(new_n3230_), .Y(new_n10156_));
  OAI22X1  g10092(.A0(new_n6936_), .A1(new_n3231_), .B0(new_n8752_), .B1(new_n3389_), .Y(new_n10157_));
  AOI21X1  g10093(.A0(new_n6933_), .A1(new_n3546_), .B0(new_n10157_), .Y(new_n10158_));
  OAI21X1  g10094(.A0(new_n8759_), .A1(new_n3388_), .B0(new_n10158_), .Y(new_n10159_));
  OR4X1    g10095(.A(new_n10159_), .B(new_n10156_), .C(new_n10155_), .D(new_n2445_), .Y(new_n10160_));
  OR2X1    g10096(.A(new_n10160_), .B(new_n9868_), .Y(new_n10161_));
  XOR2X1   g10097(.A(new_n10160_), .B(new_n9867_), .Y(new_n10162_));
  AOI22X1  g10098(.A0(new_n6935_), .A1(new_n3232_), .B0(new_n6933_), .B1(new_n3390_), .Y(new_n10163_));
  OAI21X1  g10099(.A0(new_n6930_), .A1(new_n3545_), .B0(new_n10163_), .Y(new_n10164_));
  AOI21X1  g10100(.A0(new_n8717_), .A1(new_n3234_), .B0(new_n10164_), .Y(new_n10165_));
  XOR2X1   g10101(.A(new_n10165_), .B(\a[17] ), .Y(new_n10166_));
  OAI21X1  g10102(.A0(new_n10166_), .A1(new_n10162_), .B0(new_n10161_), .Y(new_n10167_));
  XOR2X1   g10103(.A(new_n10151_), .B(new_n10147_), .Y(new_n10168_));
  AOI21X1  g10104(.A0(new_n10168_), .A1(new_n10167_), .B0(new_n10152_), .Y(new_n10169_));
  NOR2X1   g10105(.A(new_n10169_), .B(new_n10145_), .Y(new_n10170_));
  OR2X1    g10106(.A(new_n10170_), .B(new_n10144_), .Y(new_n10171_));
  XOR2X1   g10107(.A(new_n10136_), .B(new_n10132_), .Y(new_n10172_));
  AOI21X1  g10108(.A0(new_n10172_), .A1(new_n10171_), .B0(new_n10137_), .Y(new_n10173_));
  OAI21X1  g10109(.A0(new_n10173_), .A1(new_n10130_), .B0(new_n10129_), .Y(new_n10174_));
  INVX1    g10110(.A(new_n10174_), .Y(new_n10175_));
  XOR2X1   g10111(.A(new_n10119_), .B(new_n10114_), .Y(new_n10176_));
  OAI21X1  g10112(.A0(new_n10176_), .A1(new_n10175_), .B0(new_n10121_), .Y(new_n10177_));
  INVX1    g10113(.A(new_n10177_), .Y(new_n10178_));
  XOR2X1   g10114(.A(new_n10112_), .B(new_n10107_), .Y(new_n10179_));
  OAI21X1  g10115(.A0(new_n10179_), .A1(new_n10178_), .B0(new_n10113_), .Y(new_n10180_));
  XOR2X1   g10116(.A(new_n10105_), .B(new_n10101_), .Y(new_n10181_));
  AOI21X1  g10117(.A0(new_n10181_), .A1(new_n10180_), .B0(new_n10106_), .Y(new_n10182_));
  OAI21X1  g10118(.A0(new_n10182_), .A1(new_n10099_), .B0(new_n10097_), .Y(new_n10183_));
  AOI21X1  g10119(.A0(new_n10183_), .A1(new_n10091_), .B0(new_n10090_), .Y(new_n10184_));
  NOR2X1   g10120(.A(new_n10184_), .B(new_n10084_), .Y(new_n10185_));
  NOR2X1   g10121(.A(new_n10185_), .B(new_n10083_), .Y(new_n10186_));
  XOR2X1   g10122(.A(new_n10075_), .B(new_n10070_), .Y(new_n10187_));
  OAI21X1  g10123(.A0(new_n10187_), .A1(new_n10186_), .B0(new_n10076_), .Y(new_n10188_));
  XOR2X1   g10124(.A(new_n10068_), .B(new_n10064_), .Y(new_n10189_));
  AOI21X1  g10125(.A0(new_n10189_), .A1(new_n10188_), .B0(new_n10069_), .Y(new_n10190_));
  OR2X1    g10126(.A(new_n10190_), .B(new_n10063_), .Y(new_n10191_));
  AOI21X1  g10127(.A0(new_n10191_), .A1(new_n10061_), .B0(new_n10054_), .Y(new_n10192_));
  NOR2X1   g10128(.A(new_n10192_), .B(new_n10052_), .Y(new_n10193_));
  INVX1    g10129(.A(new_n10193_), .Y(new_n10194_));
  AOI21X1  g10130(.A0(new_n10194_), .A1(new_n10046_), .B0(new_n10045_), .Y(new_n10195_));
  INVX1    g10131(.A(new_n10195_), .Y(new_n10196_));
  AOI21X1  g10132(.A0(new_n10196_), .A1(new_n10039_), .B0(new_n10038_), .Y(new_n10197_));
  INVX1    g10133(.A(new_n10197_), .Y(new_n10198_));
  AOI21X1  g10134(.A0(new_n10198_), .A1(new_n10032_), .B0(new_n10031_), .Y(new_n10199_));
  INVX1    g10135(.A(new_n10199_), .Y(new_n10200_));
  AOI21X1  g10136(.A0(new_n10200_), .A1(new_n10025_), .B0(new_n10024_), .Y(new_n10201_));
  INVX1    g10137(.A(new_n10201_), .Y(new_n10202_));
  AOI21X1  g10138(.A0(new_n10202_), .A1(new_n10018_), .B0(new_n10017_), .Y(new_n10203_));
  NOR2X1   g10139(.A(new_n10203_), .B(new_n10011_), .Y(new_n10204_));
  OAI21X1  g10140(.A0(new_n10204_), .A1(new_n10009_), .B0(new_n10002_), .Y(new_n10205_));
  AND2X1   g10141(.A(new_n10205_), .B(new_n10001_), .Y(new_n10206_));
  INVX1    g10142(.A(new_n10206_), .Y(new_n10207_));
  AOI21X1  g10143(.A0(new_n10207_), .A1(new_n9994_), .B0(new_n9993_), .Y(new_n10208_));
  AOI21X1  g10144(.A0(new_n9986_), .A1(new_n9985_), .B0(new_n10208_), .Y(new_n10209_));
  NAND3X1  g10145(.A(new_n10208_), .B(new_n9986_), .C(new_n9985_), .Y(new_n10210_));
  AOI22X1  g10146(.A0(new_n7044_), .A1(new_n3908_), .B0(new_n6818_), .B1(new_n3628_), .Y(new_n10211_));
  OAI21X1  g10147(.A0(new_n7367_), .A1(new_n3983_), .B0(new_n10211_), .Y(new_n10212_));
  AOI21X1  g10148(.A0(new_n7366_), .A1(new_n3624_), .B0(new_n10212_), .Y(new_n10213_));
  XOR2X1   g10149(.A(new_n10213_), .B(\a[14] ), .Y(new_n10214_));
  INVX1    g10150(.A(new_n10214_), .Y(new_n10215_));
  AOI21X1  g10151(.A0(new_n10215_), .A1(new_n10210_), .B0(new_n10209_), .Y(new_n10216_));
  AOI21X1  g10152(.A0(new_n9984_), .A1(new_n9982_), .B0(new_n10216_), .Y(new_n10217_));
  NAND3X1  g10153(.A(new_n10216_), .B(new_n9984_), .C(new_n9982_), .Y(new_n10218_));
  AOI22X1  g10154(.A0(new_n7529_), .A1(new_n4247_), .B0(new_n7522_), .B1(new_n4078_), .Y(new_n10219_));
  OAI21X1  g10155(.A0(new_n7581_), .A1(new_n4427_), .B0(new_n10219_), .Y(new_n10220_));
  AOI21X1  g10156(.A0(new_n7565_), .A1(new_n4080_), .B0(new_n10220_), .Y(new_n10221_));
  XOR2X1   g10157(.A(new_n10221_), .B(\a[11] ), .Y(new_n10222_));
  INVX1    g10158(.A(new_n10222_), .Y(new_n10223_));
  AOI21X1  g10159(.A0(new_n10223_), .A1(new_n10218_), .B0(new_n10217_), .Y(new_n10224_));
  NOR2X1   g10160(.A(new_n10224_), .B(new_n9972_), .Y(new_n10225_));
  XOR2X1   g10161(.A(new_n10224_), .B(new_n9972_), .Y(new_n10226_));
  AOI22X1  g10162(.A0(new_n7590_), .A1(new_n4870_), .B0(new_n7578_), .B1(new_n4635_), .Y(new_n10227_));
  OAI21X1  g10163(.A0(new_n7642_), .A1(new_n5096_), .B0(new_n10227_), .Y(new_n10228_));
  AOI21X1  g10164(.A0(new_n7712_), .A1(new_n4637_), .B0(new_n10228_), .Y(new_n10229_));
  XOR2X1   g10165(.A(new_n10229_), .B(\a[8] ), .Y(new_n10230_));
  INVX1    g10166(.A(new_n10230_), .Y(new_n10231_));
  AOI21X1  g10167(.A0(new_n10231_), .A1(new_n10226_), .B0(new_n10225_), .Y(new_n10232_));
  AOI22X1  g10168(.A0(new_n7643_), .A1(new_n5097_), .B0(new_n7590_), .B1(new_n4635_), .Y(new_n10233_));
  OAI21X1  g10169(.A0(new_n7642_), .A1(new_n4869_), .B0(new_n10233_), .Y(new_n10234_));
  AOI21X1  g10170(.A0(new_n7718_), .A1(new_n4637_), .B0(new_n10234_), .Y(new_n10235_));
  XOR2X1   g10171(.A(new_n10235_), .B(\a[8] ), .Y(new_n10236_));
  NOR2X1   g10172(.A(new_n10236_), .B(new_n10232_), .Y(new_n10237_));
  XOR2X1   g10173(.A(new_n10236_), .B(new_n10232_), .Y(new_n10238_));
  XOR2X1   g10174(.A(new_n9955_), .B(new_n9705_), .Y(new_n10239_));
  AOI21X1  g10175(.A0(new_n10239_), .A1(new_n10238_), .B0(new_n10237_), .Y(new_n10240_));
  NOR2X1   g10176(.A(new_n10240_), .B(new_n9970_), .Y(new_n10241_));
  XOR2X1   g10177(.A(new_n10240_), .B(new_n9970_), .Y(new_n10242_));
  NOR3X1   g10178(.A(new_n9947_), .B(new_n9983_), .C(new_n9941_), .Y(new_n10243_));
  AOI21X1  g10179(.A0(new_n9942_), .A1(new_n9981_), .B0(new_n9946_), .Y(new_n10244_));
  NOR3X1   g10180(.A(new_n9939_), .B(new_n9979_), .C(new_n9933_), .Y(new_n10245_));
  AOI21X1  g10181(.A0(new_n9934_), .A1(new_n9978_), .B0(new_n9938_), .Y(new_n10246_));
  INVX1    g10182(.A(new_n10208_), .Y(new_n10247_));
  OAI21X1  g10183(.A0(new_n10246_), .A1(new_n10245_), .B0(new_n10247_), .Y(new_n10248_));
  NOR3X1   g10184(.A(new_n10247_), .B(new_n10246_), .C(new_n10245_), .Y(new_n10249_));
  OAI21X1  g10185(.A0(new_n10214_), .A1(new_n10249_), .B0(new_n10248_), .Y(new_n10250_));
  OAI21X1  g10186(.A0(new_n10244_), .A1(new_n10243_), .B0(new_n10250_), .Y(new_n10251_));
  NAND3X1  g10187(.A(new_n10222_), .B(new_n10218_), .C(new_n10251_), .Y(new_n10252_));
  NOR3X1   g10188(.A(new_n10250_), .B(new_n10244_), .C(new_n10243_), .Y(new_n10253_));
  OAI21X1  g10189(.A0(new_n10253_), .A1(new_n10217_), .B0(new_n10223_), .Y(new_n10254_));
  NAND3X1  g10190(.A(new_n10214_), .B(new_n10210_), .C(new_n10248_), .Y(new_n10255_));
  OAI21X1  g10191(.A0(new_n10249_), .A1(new_n10209_), .B0(new_n10215_), .Y(new_n10256_));
  XOR2X1   g10192(.A(new_n10206_), .B(new_n9994_), .Y(new_n10257_));
  OAI22X1  g10193(.A0(new_n7361_), .A1(new_n3907_), .B0(new_n7418_), .B1(new_n3627_), .Y(new_n10258_));
  AOI21X1  g10194(.A0(new_n7044_), .A1(new_n3984_), .B0(new_n10258_), .Y(new_n10259_));
  OAI21X1  g10195(.A0(new_n7680_), .A1(new_n3906_), .B0(new_n10259_), .Y(new_n10260_));
  XOR2X1   g10196(.A(new_n10260_), .B(new_n2529_), .Y(new_n10261_));
  NOR2X1   g10197(.A(new_n10261_), .B(new_n10257_), .Y(new_n10262_));
  INVX1    g10198(.A(new_n10002_), .Y(new_n10263_));
  NOR2X1   g10199(.A(new_n10204_), .B(new_n10009_), .Y(new_n10264_));
  XOR2X1   g10200(.A(new_n10264_), .B(new_n10263_), .Y(new_n10265_));
  OAI22X1  g10201(.A0(new_n7671_), .A1(new_n3627_), .B0(new_n7418_), .B1(new_n3907_), .Y(new_n10266_));
  AOI21X1  g10202(.A0(new_n6818_), .A1(new_n3984_), .B0(new_n10266_), .Y(new_n10267_));
  OAI21X1  g10203(.A0(new_n7403_), .A1(new_n3906_), .B0(new_n10267_), .Y(new_n10268_));
  XOR2X1   g10204(.A(new_n10268_), .B(new_n2529_), .Y(new_n10269_));
  INVX1    g10205(.A(new_n10269_), .Y(new_n10270_));
  NAND2X1  g10206(.A(new_n10270_), .B(new_n10265_), .Y(new_n10271_));
  XOR2X1   g10207(.A(new_n10203_), .B(new_n10011_), .Y(new_n10272_));
  OAI22X1  g10208(.A0(new_n7472_), .A1(new_n3627_), .B0(new_n7671_), .B1(new_n3907_), .Y(new_n10273_));
  AOI21X1  g10209(.A0(new_n6745_), .A1(new_n3984_), .B0(new_n10273_), .Y(new_n10274_));
  OAI21X1  g10210(.A0(new_n7416_), .A1(new_n3906_), .B0(new_n10274_), .Y(new_n10275_));
  XOR2X1   g10211(.A(new_n10275_), .B(\a[14] ), .Y(new_n10276_));
  AND2X1   g10212(.A(new_n10276_), .B(new_n10272_), .Y(new_n10277_));
  INVX1    g10213(.A(new_n10277_), .Y(new_n10278_));
  XOR2X1   g10214(.A(new_n10202_), .B(new_n10018_), .Y(new_n10279_));
  INVX1    g10215(.A(new_n7670_), .Y(new_n10280_));
  OAI22X1  g10216(.A0(new_n6884_), .A1(new_n3627_), .B0(new_n7472_), .B1(new_n3907_), .Y(new_n10281_));
  AOI21X1  g10217(.A0(new_n6820_), .A1(new_n3984_), .B0(new_n10281_), .Y(new_n10282_));
  OAI21X1  g10218(.A0(new_n10280_), .A1(new_n3906_), .B0(new_n10282_), .Y(new_n10283_));
  XOR2X1   g10219(.A(new_n10283_), .B(\a[14] ), .Y(new_n10284_));
  AND2X1   g10220(.A(new_n10284_), .B(new_n10279_), .Y(new_n10285_));
  XOR2X1   g10221(.A(new_n10200_), .B(new_n10025_), .Y(new_n10286_));
  INVX1    g10222(.A(new_n10286_), .Y(new_n10287_));
  OAI22X1  g10223(.A0(new_n6886_), .A1(new_n3627_), .B0(new_n6884_), .B1(new_n3907_), .Y(new_n10288_));
  AOI21X1  g10224(.A0(new_n6822_), .A1(new_n3984_), .B0(new_n10288_), .Y(new_n10289_));
  OAI21X1  g10225(.A0(new_n7965_), .A1(new_n3906_), .B0(new_n10289_), .Y(new_n10290_));
  XOR2X1   g10226(.A(new_n10290_), .B(new_n2529_), .Y(new_n10291_));
  XOR2X1   g10227(.A(new_n10198_), .B(new_n10032_), .Y(new_n10292_));
  AOI22X1  g10228(.A0(new_n6887_), .A1(new_n3628_), .B0(new_n6885_), .B1(new_n3908_), .Y(new_n10293_));
  OAI21X1  g10229(.A0(new_n6884_), .A1(new_n3983_), .B0(new_n10293_), .Y(new_n10294_));
  AOI21X1  g10230(.A0(new_n7771_), .A1(new_n3624_), .B0(new_n10294_), .Y(new_n10295_));
  XOR2X1   g10231(.A(new_n10295_), .B(new_n2529_), .Y(new_n10296_));
  XOR2X1   g10232(.A(new_n10196_), .B(new_n10039_), .Y(new_n10297_));
  OAI22X1  g10233(.A0(new_n7885_), .A1(new_n3627_), .B0(new_n7878_), .B1(new_n3907_), .Y(new_n10298_));
  AOI21X1  g10234(.A0(new_n6885_), .A1(new_n3984_), .B0(new_n10298_), .Y(new_n10299_));
  OAI21X1  g10235(.A0(new_n8083_), .A1(new_n3906_), .B0(new_n10299_), .Y(new_n10300_));
  XOR2X1   g10236(.A(new_n10300_), .B(\a[14] ), .Y(new_n10301_));
  AND2X1   g10237(.A(new_n10301_), .B(new_n10297_), .Y(new_n10302_));
  INVX1    g10238(.A(new_n10302_), .Y(new_n10303_));
  XOR2X1   g10239(.A(new_n10193_), .B(new_n10046_), .Y(new_n10304_));
  OAI22X1  g10240(.A0(new_n8075_), .A1(new_n3627_), .B0(new_n7885_), .B1(new_n3907_), .Y(new_n10305_));
  AOI21X1  g10241(.A0(new_n6887_), .A1(new_n3984_), .B0(new_n10305_), .Y(new_n10306_));
  OAI21X1  g10242(.A0(new_n7876_), .A1(new_n3906_), .B0(new_n10306_), .Y(new_n10307_));
  XOR2X1   g10243(.A(new_n10307_), .B(new_n2529_), .Y(new_n10308_));
  NOR2X1   g10244(.A(new_n10308_), .B(new_n10304_), .Y(new_n10309_));
  AND2X1   g10245(.A(new_n10191_), .B(new_n10061_), .Y(new_n10310_));
  XOR2X1   g10246(.A(new_n10310_), .B(new_n10054_), .Y(new_n10311_));
  OAI22X1  g10247(.A0(new_n6896_), .A1(new_n3627_), .B0(new_n8075_), .B1(new_n3907_), .Y(new_n10312_));
  AOI21X1  g10248(.A0(new_n6890_), .A1(new_n3984_), .B0(new_n10312_), .Y(new_n10313_));
  OAI21X1  g10249(.A0(new_n9738_), .A1(new_n3906_), .B0(new_n10313_), .Y(new_n10314_));
  XOR2X1   g10250(.A(new_n10314_), .B(\a[14] ), .Y(new_n10315_));
  AND2X1   g10251(.A(new_n10315_), .B(new_n10311_), .Y(new_n10316_));
  XOR2X1   g10252(.A(new_n10190_), .B(new_n10063_), .Y(new_n10317_));
  OAI22X1  g10253(.A0(new_n6898_), .A1(new_n3627_), .B0(new_n6896_), .B1(new_n3907_), .Y(new_n10318_));
  AOI21X1  g10254(.A0(new_n6892_), .A1(new_n3984_), .B0(new_n10318_), .Y(new_n10319_));
  OAI21X1  g10255(.A0(new_n9744_), .A1(new_n3906_), .B0(new_n10319_), .Y(new_n10320_));
  XOR2X1   g10256(.A(new_n10320_), .B(\a[14] ), .Y(new_n10321_));
  AOI22X1  g10257(.A0(new_n6899_), .A1(new_n3628_), .B0(new_n6897_), .B1(new_n3908_), .Y(new_n10322_));
  OAI21X1  g10258(.A0(new_n6896_), .A1(new_n3983_), .B0(new_n10322_), .Y(new_n10323_));
  AOI21X1  g10259(.A0(new_n7953_), .A1(new_n3624_), .B0(new_n10323_), .Y(new_n10324_));
  XOR2X1   g10260(.A(new_n10324_), .B(\a[14] ), .Y(new_n10325_));
  INVX1    g10261(.A(new_n10325_), .Y(new_n10326_));
  XOR2X1   g10262(.A(new_n10189_), .B(new_n10188_), .Y(new_n10327_));
  XOR2X1   g10263(.A(new_n10327_), .B(new_n10325_), .Y(new_n10328_));
  AOI22X1  g10264(.A0(new_n6902_), .A1(new_n3628_), .B0(new_n6899_), .B1(new_n3908_), .Y(new_n10329_));
  OAI21X1  g10265(.A0(new_n6898_), .A1(new_n3983_), .B0(new_n10329_), .Y(new_n10330_));
  AOI21X1  g10266(.A0(new_n8215_), .A1(new_n3624_), .B0(new_n10330_), .Y(new_n10331_));
  XOR2X1   g10267(.A(new_n10331_), .B(\a[14] ), .Y(new_n10332_));
  XOR2X1   g10268(.A(new_n10075_), .B(new_n10071_), .Y(new_n10333_));
  XOR2X1   g10269(.A(new_n10333_), .B(new_n10186_), .Y(new_n10334_));
  NOR2X1   g10270(.A(new_n10334_), .B(new_n10332_), .Y(new_n10335_));
  INVX1    g10271(.A(new_n10335_), .Y(new_n10336_));
  XOR2X1   g10272(.A(new_n10334_), .B(new_n10332_), .Y(new_n10337_));
  INVX1    g10273(.A(new_n10337_), .Y(new_n10338_));
  INVX1    g10274(.A(new_n10084_), .Y(new_n10339_));
  XOR2X1   g10275(.A(new_n10184_), .B(new_n10339_), .Y(new_n10340_));
  OAI22X1  g10276(.A0(new_n8200_), .A1(new_n3627_), .B0(new_n8205_), .B1(new_n3907_), .Y(new_n10341_));
  AOI21X1  g10277(.A0(new_n6899_), .A1(new_n3984_), .B0(new_n10341_), .Y(new_n10342_));
  OAI21X1  g10278(.A0(new_n8293_), .A1(new_n3906_), .B0(new_n10342_), .Y(new_n10343_));
  XOR2X1   g10279(.A(new_n10343_), .B(new_n2529_), .Y(new_n10344_));
  NOR2X1   g10280(.A(new_n10344_), .B(new_n10340_), .Y(new_n10345_));
  XOR2X1   g10281(.A(new_n10183_), .B(new_n10091_), .Y(new_n10346_));
  OAI22X1  g10282(.A0(new_n6964_), .A1(new_n3627_), .B0(new_n8200_), .B1(new_n3907_), .Y(new_n10347_));
  AOI21X1  g10283(.A0(new_n6902_), .A1(new_n3984_), .B0(new_n10347_), .Y(new_n10348_));
  OAI21X1  g10284(.A0(new_n8203_), .A1(new_n3906_), .B0(new_n10348_), .Y(new_n10349_));
  XOR2X1   g10285(.A(new_n10349_), .B(\a[14] ), .Y(new_n10350_));
  NAND2X1  g10286(.A(new_n10350_), .B(new_n10346_), .Y(new_n10351_));
  XOR2X1   g10287(.A(new_n10182_), .B(new_n10099_), .Y(new_n10352_));
  INVX1    g10288(.A(new_n10352_), .Y(new_n10353_));
  OAI22X1  g10289(.A0(new_n6960_), .A1(new_n3627_), .B0(new_n6964_), .B1(new_n3907_), .Y(new_n10354_));
  AOI21X1  g10290(.A0(new_n6904_), .A1(new_n3984_), .B0(new_n10354_), .Y(new_n10355_));
  OAI21X1  g10291(.A0(new_n8364_), .A1(new_n3906_), .B0(new_n10355_), .Y(new_n10356_));
  XOR2X1   g10292(.A(new_n10356_), .B(new_n2529_), .Y(new_n10357_));
  NOR2X1   g10293(.A(new_n10357_), .B(new_n10353_), .Y(new_n10358_));
  INVX1    g10294(.A(new_n10358_), .Y(new_n10359_));
  AOI22X1  g10295(.A0(new_n6911_), .A1(new_n3628_), .B0(new_n6909_), .B1(new_n3908_), .Y(new_n10360_));
  OAI21X1  g10296(.A0(new_n6964_), .A1(new_n3983_), .B0(new_n10360_), .Y(new_n10361_));
  AOI21X1  g10297(.A0(new_n8541_), .A1(new_n3624_), .B0(new_n10361_), .Y(new_n10362_));
  XOR2X1   g10298(.A(new_n10362_), .B(\a[14] ), .Y(new_n10363_));
  INVX1    g10299(.A(new_n10363_), .Y(new_n10364_));
  XOR2X1   g10300(.A(new_n10181_), .B(new_n10180_), .Y(new_n10365_));
  XOR2X1   g10301(.A(new_n10365_), .B(new_n10363_), .Y(new_n10366_));
  AOI22X1  g10302(.A0(new_n6913_), .A1(new_n3628_), .B0(new_n6911_), .B1(new_n3908_), .Y(new_n10367_));
  OAI21X1  g10303(.A0(new_n6960_), .A1(new_n3983_), .B0(new_n10367_), .Y(new_n10368_));
  AOI21X1  g10304(.A0(new_n8553_), .A1(new_n3624_), .B0(new_n10368_), .Y(new_n10369_));
  XOR2X1   g10305(.A(new_n10369_), .B(\a[14] ), .Y(new_n10370_));
  XOR2X1   g10306(.A(new_n10179_), .B(new_n10177_), .Y(new_n10371_));
  NOR2X1   g10307(.A(new_n10371_), .B(new_n10370_), .Y(new_n10372_));
  XOR2X1   g10308(.A(new_n10371_), .B(new_n10370_), .Y(new_n10373_));
  AOI22X1  g10309(.A0(new_n6915_), .A1(new_n3628_), .B0(new_n6913_), .B1(new_n3908_), .Y(new_n10374_));
  OAI21X1  g10310(.A0(new_n8349_), .A1(new_n3983_), .B0(new_n10374_), .Y(new_n10375_));
  AOI21X1  g10311(.A0(new_n8348_), .A1(new_n3624_), .B0(new_n10375_), .Y(new_n10376_));
  XOR2X1   g10312(.A(new_n10376_), .B(\a[14] ), .Y(new_n10377_));
  XOR2X1   g10313(.A(new_n10176_), .B(new_n10174_), .Y(new_n10378_));
  OR2X1    g10314(.A(new_n10378_), .B(new_n10377_), .Y(new_n10379_));
  XOR2X1   g10315(.A(new_n10378_), .B(new_n10377_), .Y(new_n10380_));
  INVX1    g10316(.A(new_n10380_), .Y(new_n10381_));
  INVX1    g10317(.A(new_n10130_), .Y(new_n10382_));
  XOR2X1   g10318(.A(new_n10173_), .B(new_n10382_), .Y(new_n10383_));
  OAI22X1  g10319(.A0(new_n6918_), .A1(new_n3627_), .B0(new_n6917_), .B1(new_n3907_), .Y(new_n10384_));
  AOI21X1  g10320(.A0(new_n6913_), .A1(new_n3984_), .B0(new_n10384_), .Y(new_n10385_));
  OAI21X1  g10321(.A0(new_n8577_), .A1(new_n3906_), .B0(new_n10385_), .Y(new_n10386_));
  XOR2X1   g10322(.A(new_n10386_), .B(new_n2529_), .Y(new_n10387_));
  NOR2X1   g10323(.A(new_n10387_), .B(new_n10383_), .Y(new_n10388_));
  XOR2X1   g10324(.A(new_n10172_), .B(new_n10171_), .Y(new_n10389_));
  INVX1    g10325(.A(new_n10389_), .Y(new_n10390_));
  OAI22X1  g10326(.A0(new_n6920_), .A1(new_n3627_), .B0(new_n6918_), .B1(new_n3907_), .Y(new_n10391_));
  AOI21X1  g10327(.A0(new_n6915_), .A1(new_n3984_), .B0(new_n10391_), .Y(new_n10392_));
  OAI21X1  g10328(.A0(new_n9093_), .A1(new_n3906_), .B0(new_n10392_), .Y(new_n10393_));
  XOR2X1   g10329(.A(new_n10393_), .B(new_n2529_), .Y(new_n10394_));
  OR2X1    g10330(.A(new_n10394_), .B(new_n10390_), .Y(new_n10395_));
  XOR2X1   g10331(.A(new_n10169_), .B(new_n10145_), .Y(new_n10396_));
  INVX1    g10332(.A(new_n10396_), .Y(new_n10397_));
  OAI22X1  g10333(.A0(new_n8659_), .A1(new_n3627_), .B0(new_n6920_), .B1(new_n3907_), .Y(new_n10398_));
  AOI21X1  g10334(.A0(new_n8580_), .A1(new_n3984_), .B0(new_n10398_), .Y(new_n10399_));
  OAI21X1  g10335(.A0(new_n8611_), .A1(new_n3906_), .B0(new_n10399_), .Y(new_n10400_));
  XOR2X1   g10336(.A(new_n10400_), .B(new_n2529_), .Y(new_n10401_));
  NOR2X1   g10337(.A(new_n10401_), .B(new_n10397_), .Y(new_n10402_));
  INVX1    g10338(.A(new_n10402_), .Y(new_n10403_));
  AOI22X1  g10339(.A0(new_n6925_), .A1(new_n3628_), .B0(new_n6923_), .B1(new_n3908_), .Y(new_n10404_));
  OAI21X1  g10340(.A0(new_n6920_), .A1(new_n3983_), .B0(new_n10404_), .Y(new_n10405_));
  AOI21X1  g10341(.A0(new_n8628_), .A1(new_n3624_), .B0(new_n10405_), .Y(new_n10406_));
  XOR2X1   g10342(.A(new_n10406_), .B(\a[14] ), .Y(new_n10407_));
  INVX1    g10343(.A(new_n10407_), .Y(new_n10408_));
  XOR2X1   g10344(.A(new_n10168_), .B(new_n10167_), .Y(new_n10409_));
  AND2X1   g10345(.A(new_n10409_), .B(new_n10408_), .Y(new_n10410_));
  INVX1    g10346(.A(new_n10410_), .Y(new_n10411_));
  XOR2X1   g10347(.A(new_n10409_), .B(new_n10407_), .Y(new_n10412_));
  XOR2X1   g10348(.A(new_n10165_), .B(new_n2445_), .Y(new_n10413_));
  XOR2X1   g10349(.A(new_n10413_), .B(new_n10162_), .Y(new_n10414_));
  OAI22X1  g10350(.A0(new_n6929_), .A1(new_n3627_), .B0(new_n8683_), .B1(new_n3907_), .Y(new_n10415_));
  AOI21X1  g10351(.A0(new_n6923_), .A1(new_n3984_), .B0(new_n10415_), .Y(new_n10416_));
  OAI21X1  g10352(.A0(new_n8662_), .A1(new_n3906_), .B0(new_n10416_), .Y(new_n10417_));
  XOR2X1   g10353(.A(new_n10417_), .B(new_n2529_), .Y(new_n10418_));
  NOR2X1   g10354(.A(new_n10418_), .B(new_n10414_), .Y(new_n10419_));
  AOI22X1  g10355(.A0(new_n6932_), .A1(new_n3628_), .B0(new_n6927_), .B1(new_n3908_), .Y(new_n10420_));
  OAI21X1  g10356(.A0(new_n8683_), .A1(new_n3983_), .B0(new_n10420_), .Y(new_n10421_));
  AOI21X1  g10357(.A0(new_n8682_), .A1(new_n3624_), .B0(new_n10421_), .Y(new_n10422_));
  XOR2X1   g10358(.A(new_n10422_), .B(\a[14] ), .Y(new_n10423_));
  INVX1    g10359(.A(new_n10423_), .Y(new_n10424_));
  NOR3X1   g10360(.A(new_n10156_), .B(new_n10155_), .C(new_n2445_), .Y(new_n10425_));
  XOR2X1   g10361(.A(new_n10159_), .B(\a[17] ), .Y(new_n10426_));
  XOR2X1   g10362(.A(new_n10426_), .B(new_n10425_), .Y(new_n10427_));
  AND2X1   g10363(.A(new_n10427_), .B(new_n10424_), .Y(new_n10428_));
  XOR2X1   g10364(.A(new_n10427_), .B(new_n10423_), .Y(new_n10429_));
  NOR2X1   g10365(.A(new_n10156_), .B(new_n2445_), .Y(new_n10430_));
  XOR2X1   g10366(.A(new_n10430_), .B(new_n10155_), .Y(new_n10431_));
  OAI22X1  g10367(.A0(new_n8757_), .A1(new_n3627_), .B0(new_n6930_), .B1(new_n3907_), .Y(new_n10432_));
  AOI21X1  g10368(.A0(new_n6927_), .A1(new_n3984_), .B0(new_n10432_), .Y(new_n10433_));
  OAI21X1  g10369(.A0(new_n8705_), .A1(new_n3906_), .B0(new_n10433_), .Y(new_n10434_));
  XOR2X1   g10370(.A(new_n10434_), .B(new_n2529_), .Y(new_n10435_));
  NOR2X1   g10371(.A(new_n10435_), .B(new_n10431_), .Y(new_n10436_));
  OAI22X1  g10372(.A0(new_n6936_), .A1(new_n3907_), .B0(new_n8752_), .B1(new_n3983_), .Y(new_n10437_));
  AOI21X1  g10373(.A0(new_n8751_), .A1(new_n3624_), .B0(new_n10437_), .Y(new_n10438_));
  NOR2X1   g10374(.A(new_n6936_), .B(new_n3621_), .Y(new_n10439_));
  INVX1    g10375(.A(new_n10439_), .Y(new_n10440_));
  NAND3X1  g10376(.A(new_n10440_), .B(new_n10438_), .C(\a[14] ), .Y(new_n10441_));
  OAI22X1  g10377(.A0(new_n6936_), .A1(new_n3627_), .B0(new_n8752_), .B1(new_n3907_), .Y(new_n10442_));
  AOI21X1  g10378(.A0(new_n6933_), .A1(new_n3984_), .B0(new_n10442_), .Y(new_n10443_));
  OAI21X1  g10379(.A0(new_n8759_), .A1(new_n3906_), .B0(new_n10443_), .Y(new_n10444_));
  XOR2X1   g10380(.A(new_n10444_), .B(new_n2529_), .Y(new_n10445_));
  OR4X1    g10381(.A(new_n10445_), .B(new_n10441_), .C(new_n6936_), .D(new_n3230_), .Y(new_n10446_));
  XOR2X1   g10382(.A(new_n10438_), .B(\a[14] ), .Y(new_n10447_));
  OR4X1    g10383(.A(new_n10444_), .B(new_n10439_), .C(new_n10447_), .D(new_n2529_), .Y(new_n10448_));
  XOR2X1   g10384(.A(new_n10448_), .B(new_n10156_), .Y(new_n10449_));
  AOI22X1  g10385(.A0(new_n6935_), .A1(new_n3628_), .B0(new_n6933_), .B1(new_n3908_), .Y(new_n10450_));
  OAI21X1  g10386(.A0(new_n6930_), .A1(new_n3983_), .B0(new_n10450_), .Y(new_n10451_));
  AOI21X1  g10387(.A0(new_n8717_), .A1(new_n3624_), .B0(new_n10451_), .Y(new_n10452_));
  XOR2X1   g10388(.A(new_n10452_), .B(\a[14] ), .Y(new_n10453_));
  OAI21X1  g10389(.A0(new_n10453_), .A1(new_n10449_), .B0(new_n10446_), .Y(new_n10454_));
  XOR2X1   g10390(.A(new_n10435_), .B(new_n10431_), .Y(new_n10455_));
  AOI21X1  g10391(.A0(new_n10455_), .A1(new_n10454_), .B0(new_n10436_), .Y(new_n10456_));
  NOR2X1   g10392(.A(new_n10456_), .B(new_n10429_), .Y(new_n10457_));
  OR2X1    g10393(.A(new_n10457_), .B(new_n10428_), .Y(new_n10458_));
  XOR2X1   g10394(.A(new_n10418_), .B(new_n10414_), .Y(new_n10459_));
  AOI21X1  g10395(.A0(new_n10459_), .A1(new_n10458_), .B0(new_n10419_), .Y(new_n10460_));
  OAI21X1  g10396(.A0(new_n10460_), .A1(new_n10412_), .B0(new_n10411_), .Y(new_n10461_));
  INVX1    g10397(.A(new_n10461_), .Y(new_n10462_));
  XOR2X1   g10398(.A(new_n10401_), .B(new_n10396_), .Y(new_n10463_));
  OAI21X1  g10399(.A0(new_n10463_), .A1(new_n10462_), .B0(new_n10403_), .Y(new_n10464_));
  INVX1    g10400(.A(new_n10464_), .Y(new_n10465_));
  XOR2X1   g10401(.A(new_n10394_), .B(new_n10389_), .Y(new_n10466_));
  OAI21X1  g10402(.A0(new_n10466_), .A1(new_n10465_), .B0(new_n10395_), .Y(new_n10467_));
  XOR2X1   g10403(.A(new_n10387_), .B(new_n10383_), .Y(new_n10468_));
  AOI21X1  g10404(.A0(new_n10468_), .A1(new_n10467_), .B0(new_n10388_), .Y(new_n10469_));
  OAI21X1  g10405(.A0(new_n10469_), .A1(new_n10381_), .B0(new_n10379_), .Y(new_n10470_));
  AOI21X1  g10406(.A0(new_n10470_), .A1(new_n10373_), .B0(new_n10372_), .Y(new_n10471_));
  NOR2X1   g10407(.A(new_n10471_), .B(new_n10366_), .Y(new_n10472_));
  AOI21X1  g10408(.A0(new_n10365_), .A1(new_n10364_), .B0(new_n10472_), .Y(new_n10473_));
  XOR2X1   g10409(.A(new_n10357_), .B(new_n10352_), .Y(new_n10474_));
  OAI21X1  g10410(.A0(new_n10474_), .A1(new_n10473_), .B0(new_n10359_), .Y(new_n10475_));
  INVX1    g10411(.A(new_n10475_), .Y(new_n10476_));
  XOR2X1   g10412(.A(new_n10349_), .B(new_n2529_), .Y(new_n10477_));
  XOR2X1   g10413(.A(new_n10477_), .B(new_n10346_), .Y(new_n10478_));
  OAI21X1  g10414(.A0(new_n10478_), .A1(new_n10476_), .B0(new_n10351_), .Y(new_n10479_));
  XOR2X1   g10415(.A(new_n10344_), .B(new_n10340_), .Y(new_n10480_));
  AOI21X1  g10416(.A0(new_n10480_), .A1(new_n10479_), .B0(new_n10345_), .Y(new_n10481_));
  OR2X1    g10417(.A(new_n10481_), .B(new_n10338_), .Y(new_n10482_));
  AOI21X1  g10418(.A0(new_n10482_), .A1(new_n10336_), .B0(new_n10328_), .Y(new_n10483_));
  AOI21X1  g10419(.A0(new_n10327_), .A1(new_n10326_), .B0(new_n10483_), .Y(new_n10484_));
  XOR2X1   g10420(.A(new_n10320_), .B(new_n2529_), .Y(new_n10485_));
  XOR2X1   g10421(.A(new_n10485_), .B(new_n10317_), .Y(new_n10486_));
  NOR2X1   g10422(.A(new_n10486_), .B(new_n10484_), .Y(new_n10487_));
  AOI21X1  g10423(.A0(new_n10321_), .A1(new_n10317_), .B0(new_n10487_), .Y(new_n10488_));
  XOR2X1   g10424(.A(new_n10314_), .B(new_n2529_), .Y(new_n10489_));
  XOR2X1   g10425(.A(new_n10489_), .B(new_n10311_), .Y(new_n10490_));
  NOR2X1   g10426(.A(new_n10490_), .B(new_n10488_), .Y(new_n10491_));
  NOR2X1   g10427(.A(new_n10491_), .B(new_n10316_), .Y(new_n10492_));
  INVX1    g10428(.A(new_n10492_), .Y(new_n10493_));
  XOR2X1   g10429(.A(new_n10308_), .B(new_n10304_), .Y(new_n10494_));
  AOI21X1  g10430(.A0(new_n10494_), .A1(new_n10493_), .B0(new_n10309_), .Y(new_n10495_));
  XOR2X1   g10431(.A(new_n10300_), .B(new_n2529_), .Y(new_n10496_));
  XOR2X1   g10432(.A(new_n10496_), .B(new_n10297_), .Y(new_n10497_));
  OR2X1    g10433(.A(new_n10497_), .B(new_n10495_), .Y(new_n10498_));
  XOR2X1   g10434(.A(new_n10295_), .B(\a[14] ), .Y(new_n10499_));
  XOR2X1   g10435(.A(new_n10499_), .B(new_n10292_), .Y(new_n10500_));
  AOI21X1  g10436(.A0(new_n10498_), .A1(new_n10303_), .B0(new_n10500_), .Y(new_n10501_));
  AOI21X1  g10437(.A0(new_n10296_), .A1(new_n10292_), .B0(new_n10501_), .Y(new_n10502_));
  XOR2X1   g10438(.A(new_n10291_), .B(new_n10286_), .Y(new_n10503_));
  OR2X1    g10439(.A(new_n10503_), .B(new_n10502_), .Y(new_n10504_));
  OAI21X1  g10440(.A0(new_n10291_), .A1(new_n10287_), .B0(new_n10504_), .Y(new_n10505_));
  XOR2X1   g10441(.A(new_n10283_), .B(new_n2529_), .Y(new_n10506_));
  XOR2X1   g10442(.A(new_n10506_), .B(new_n10279_), .Y(new_n10507_));
  INVX1    g10443(.A(new_n10507_), .Y(new_n10508_));
  AOI21X1  g10444(.A0(new_n10508_), .A1(new_n10505_), .B0(new_n10285_), .Y(new_n10509_));
  XOR2X1   g10445(.A(new_n10275_), .B(new_n2529_), .Y(new_n10510_));
  XOR2X1   g10446(.A(new_n10510_), .B(new_n10272_), .Y(new_n10511_));
  OAI21X1  g10447(.A0(new_n10511_), .A1(new_n10509_), .B0(new_n10278_), .Y(new_n10512_));
  INVX1    g10448(.A(new_n10512_), .Y(new_n10513_));
  XOR2X1   g10449(.A(new_n10269_), .B(new_n10265_), .Y(new_n10514_));
  OAI21X1  g10450(.A0(new_n10514_), .A1(new_n10513_), .B0(new_n10271_), .Y(new_n10515_));
  XOR2X1   g10451(.A(new_n10261_), .B(new_n10257_), .Y(new_n10516_));
  AOI21X1  g10452(.A0(new_n10516_), .A1(new_n10515_), .B0(new_n10262_), .Y(new_n10517_));
  AOI21X1  g10453(.A0(new_n10256_), .A1(new_n10255_), .B0(new_n10517_), .Y(new_n10518_));
  NAND3X1  g10454(.A(new_n10517_), .B(new_n10256_), .C(new_n10255_), .Y(new_n10519_));
  AOI22X1  g10455(.A0(new_n7522_), .A1(new_n4247_), .B0(new_n7485_), .B1(new_n4078_), .Y(new_n10520_));
  OAI21X1  g10456(.A0(new_n7537_), .A1(new_n4427_), .B0(new_n10520_), .Y(new_n10521_));
  AOI21X1  g10457(.A0(new_n7536_), .A1(new_n4080_), .B0(new_n10521_), .Y(new_n10522_));
  XOR2X1   g10458(.A(new_n10522_), .B(\a[11] ), .Y(new_n10523_));
  INVX1    g10459(.A(new_n10523_), .Y(new_n10524_));
  AOI21X1  g10460(.A0(new_n10524_), .A1(new_n10519_), .B0(new_n10518_), .Y(new_n10525_));
  AOI21X1  g10461(.A0(new_n10254_), .A1(new_n10252_), .B0(new_n10525_), .Y(new_n10526_));
  NAND3X1  g10462(.A(new_n10525_), .B(new_n10254_), .C(new_n10252_), .Y(new_n10527_));
  AOI22X1  g10463(.A0(new_n7578_), .A1(new_n4870_), .B0(new_n7571_), .B1(new_n4635_), .Y(new_n10528_));
  OAI21X1  g10464(.A0(new_n7594_), .A1(new_n5096_), .B0(new_n10528_), .Y(new_n10529_));
  AOI21X1  g10465(.A0(new_n7593_), .A1(new_n4637_), .B0(new_n10529_), .Y(new_n10530_));
  XOR2X1   g10466(.A(new_n10530_), .B(\a[8] ), .Y(new_n10531_));
  INVX1    g10467(.A(new_n10531_), .Y(new_n10532_));
  AOI21X1  g10468(.A0(new_n10532_), .A1(new_n10527_), .B0(new_n10526_), .Y(new_n10533_));
  MX2X1    g10469(.A(new_n5370_), .B(new_n5958_), .S0(new_n66_), .Y(new_n10534_));
  AOI22X1  g10470(.A0(new_n10534_), .A1(new_n7341_), .B0(new_n7643_), .B1(new_n5373_), .Y(new_n10535_));
  OAI21X1  g10471(.A0(new_n7808_), .A1(new_n5657_), .B0(new_n10535_), .Y(new_n10536_));
  XOR2X1   g10472(.A(new_n10536_), .B(new_n3289_), .Y(new_n10537_));
  OR2X1    g10473(.A(new_n10537_), .B(new_n10533_), .Y(new_n10538_));
  XOR2X1   g10474(.A(new_n10231_), .B(new_n10226_), .Y(new_n10539_));
  XOR2X1   g10475(.A(new_n10537_), .B(new_n10533_), .Y(new_n10540_));
  NAND2X1  g10476(.A(new_n10540_), .B(new_n10539_), .Y(new_n10541_));
  NAND2X1  g10477(.A(new_n10541_), .B(new_n10538_), .Y(new_n10542_));
  XOR2X1   g10478(.A(new_n10239_), .B(new_n10238_), .Y(new_n10543_));
  NAND2X1  g10479(.A(new_n10543_), .B(new_n10542_), .Y(new_n10544_));
  XOR2X1   g10480(.A(new_n10230_), .B(new_n10226_), .Y(new_n10545_));
  XOR2X1   g10481(.A(new_n10540_), .B(new_n10545_), .Y(new_n10546_));
  NOR3X1   g10482(.A(new_n10223_), .B(new_n10253_), .C(new_n10217_), .Y(new_n10547_));
  AOI21X1  g10483(.A0(new_n10218_), .A1(new_n10251_), .B0(new_n10222_), .Y(new_n10548_));
  NOR3X1   g10484(.A(new_n10215_), .B(new_n10249_), .C(new_n10209_), .Y(new_n10549_));
  AOI21X1  g10485(.A0(new_n10210_), .A1(new_n10248_), .B0(new_n10214_), .Y(new_n10550_));
  INVX1    g10486(.A(new_n10517_), .Y(new_n10551_));
  OAI21X1  g10487(.A0(new_n10550_), .A1(new_n10549_), .B0(new_n10551_), .Y(new_n10552_));
  NOR3X1   g10488(.A(new_n10551_), .B(new_n10550_), .C(new_n10549_), .Y(new_n10553_));
  OAI21X1  g10489(.A0(new_n10523_), .A1(new_n10553_), .B0(new_n10552_), .Y(new_n10554_));
  OAI21X1  g10490(.A0(new_n10548_), .A1(new_n10547_), .B0(new_n10554_), .Y(new_n10555_));
  NAND3X1  g10491(.A(new_n10531_), .B(new_n10527_), .C(new_n10555_), .Y(new_n10556_));
  NOR3X1   g10492(.A(new_n10554_), .B(new_n10548_), .C(new_n10547_), .Y(new_n10557_));
  OAI21X1  g10493(.A0(new_n10557_), .A1(new_n10526_), .B0(new_n10532_), .Y(new_n10558_));
  NAND3X1  g10494(.A(new_n10523_), .B(new_n10519_), .C(new_n10552_), .Y(new_n10559_));
  OAI21X1  g10495(.A0(new_n10553_), .A1(new_n10518_), .B0(new_n10524_), .Y(new_n10560_));
  AOI22X1  g10496(.A0(new_n7485_), .A1(new_n4247_), .B0(new_n7364_), .B1(new_n4078_), .Y(new_n10561_));
  OAI21X1  g10497(.A0(new_n7523_), .A1(new_n4427_), .B0(new_n10561_), .Y(new_n10562_));
  AOI21X1  g10498(.A0(new_n7612_), .A1(new_n4080_), .B0(new_n10562_), .Y(new_n10563_));
  XOR2X1   g10499(.A(new_n10563_), .B(\a[11] ), .Y(new_n10564_));
  INVX1    g10500(.A(new_n10564_), .Y(new_n10565_));
  XOR2X1   g10501(.A(new_n10516_), .B(new_n10515_), .Y(new_n10566_));
  AND2X1   g10502(.A(new_n10566_), .B(new_n10565_), .Y(new_n10567_));
  XOR2X1   g10503(.A(new_n10566_), .B(new_n10565_), .Y(new_n10568_));
  AOI22X1  g10504(.A0(new_n7364_), .A1(new_n4247_), .B0(new_n7044_), .B1(new_n4078_), .Y(new_n10569_));
  OAI21X1  g10505(.A0(new_n7504_), .A1(new_n4427_), .B0(new_n10569_), .Y(new_n10570_));
  AOI21X1  g10506(.A0(new_n7552_), .A1(new_n4080_), .B0(new_n10570_), .Y(new_n10571_));
  XOR2X1   g10507(.A(new_n10571_), .B(\a[11] ), .Y(new_n10572_));
  XOR2X1   g10508(.A(new_n10514_), .B(new_n10512_), .Y(new_n10573_));
  NOR2X1   g10509(.A(new_n10573_), .B(new_n10572_), .Y(new_n10574_));
  XOR2X1   g10510(.A(new_n10573_), .B(new_n10572_), .Y(new_n10575_));
  AOI22X1  g10511(.A0(new_n7044_), .A1(new_n4247_), .B0(new_n6818_), .B1(new_n4078_), .Y(new_n10576_));
  OAI21X1  g10512(.A0(new_n7367_), .A1(new_n4427_), .B0(new_n10576_), .Y(new_n10577_));
  AOI21X1  g10513(.A0(new_n7366_), .A1(new_n4080_), .B0(new_n10577_), .Y(new_n10578_));
  XOR2X1   g10514(.A(new_n10578_), .B(\a[11] ), .Y(new_n10579_));
  INVX1    g10515(.A(new_n10511_), .Y(new_n10580_));
  XOR2X1   g10516(.A(new_n10580_), .B(new_n10509_), .Y(new_n10581_));
  XOR2X1   g10517(.A(new_n10581_), .B(new_n10579_), .Y(new_n10582_));
  INVX1    g10518(.A(new_n10582_), .Y(new_n10583_));
  AOI22X1  g10519(.A0(new_n6818_), .A1(new_n4247_), .B0(new_n6745_), .B1(new_n4078_), .Y(new_n10584_));
  OAI21X1  g10520(.A0(new_n7047_), .A1(new_n4427_), .B0(new_n10584_), .Y(new_n10585_));
  AOI21X1  g10521(.A0(new_n7046_), .A1(new_n4080_), .B0(new_n10585_), .Y(new_n10586_));
  XOR2X1   g10522(.A(new_n10586_), .B(\a[11] ), .Y(new_n10587_));
  XOR2X1   g10523(.A(new_n10507_), .B(new_n10505_), .Y(new_n10588_));
  NOR2X1   g10524(.A(new_n10588_), .B(new_n10587_), .Y(new_n10589_));
  XOR2X1   g10525(.A(new_n10588_), .B(new_n10587_), .Y(new_n10590_));
  AOI22X1  g10526(.A0(new_n6820_), .A1(new_n4078_), .B0(new_n6745_), .B1(new_n4247_), .Y(new_n10591_));
  OAI21X1  g10527(.A0(new_n7361_), .A1(new_n4427_), .B0(new_n10591_), .Y(new_n10592_));
  AOI21X1  g10528(.A0(new_n7404_), .A1(new_n4080_), .B0(new_n10592_), .Y(new_n10593_));
  XOR2X1   g10529(.A(new_n10593_), .B(\a[11] ), .Y(new_n10594_));
  INVX1    g10530(.A(new_n10503_), .Y(new_n10595_));
  XOR2X1   g10531(.A(new_n10595_), .B(new_n10502_), .Y(new_n10596_));
  XOR2X1   g10532(.A(new_n10596_), .B(new_n10594_), .Y(new_n10597_));
  INVX1    g10533(.A(new_n10597_), .Y(new_n10598_));
  AOI22X1  g10534(.A0(new_n6822_), .A1(new_n4078_), .B0(new_n6820_), .B1(new_n4247_), .Y(new_n10599_));
  OAI21X1  g10535(.A0(new_n7418_), .A1(new_n4427_), .B0(new_n10599_), .Y(new_n10600_));
  AOI21X1  g10536(.A0(new_n7417_), .A1(new_n4080_), .B0(new_n10600_), .Y(new_n10601_));
  XOR2X1   g10537(.A(new_n10601_), .B(\a[11] ), .Y(new_n10602_));
  AND2X1   g10538(.A(new_n10498_), .B(new_n10303_), .Y(new_n10603_));
  INVX1    g10539(.A(new_n10500_), .Y(new_n10604_));
  XOR2X1   g10540(.A(new_n10604_), .B(new_n10603_), .Y(new_n10605_));
  NOR2X1   g10541(.A(new_n10605_), .B(new_n10602_), .Y(new_n10606_));
  XOR2X1   g10542(.A(new_n10605_), .B(new_n10602_), .Y(new_n10607_));
  AOI22X1  g10543(.A0(new_n6882_), .A1(new_n4078_), .B0(new_n6822_), .B1(new_n4247_), .Y(new_n10608_));
  OAI21X1  g10544(.A0(new_n7671_), .A1(new_n4427_), .B0(new_n10608_), .Y(new_n10609_));
  AOI21X1  g10545(.A0(new_n7670_), .A1(new_n4080_), .B0(new_n10609_), .Y(new_n10610_));
  XOR2X1   g10546(.A(new_n10610_), .B(\a[11] ), .Y(new_n10611_));
  INVX1    g10547(.A(new_n10497_), .Y(new_n10612_));
  XOR2X1   g10548(.A(new_n10612_), .B(new_n10495_), .Y(new_n10613_));
  NOR2X1   g10549(.A(new_n10613_), .B(new_n10611_), .Y(new_n10614_));
  XOR2X1   g10550(.A(new_n10613_), .B(new_n10611_), .Y(new_n10615_));
  AOI22X1  g10551(.A0(new_n6885_), .A1(new_n4078_), .B0(new_n6882_), .B1(new_n4247_), .Y(new_n10616_));
  OAI21X1  g10552(.A0(new_n7472_), .A1(new_n4427_), .B0(new_n10616_), .Y(new_n10617_));
  AOI21X1  g10553(.A0(new_n7471_), .A1(new_n4080_), .B0(new_n10617_), .Y(new_n10618_));
  XOR2X1   g10554(.A(new_n10618_), .B(\a[11] ), .Y(new_n10619_));
  XOR2X1   g10555(.A(new_n10494_), .B(new_n10492_), .Y(new_n10620_));
  NOR2X1   g10556(.A(new_n10620_), .B(new_n10619_), .Y(new_n10621_));
  XOR2X1   g10557(.A(new_n10620_), .B(new_n10619_), .Y(new_n10622_));
  AOI22X1  g10558(.A0(new_n6887_), .A1(new_n4078_), .B0(new_n6885_), .B1(new_n4247_), .Y(new_n10623_));
  OAI21X1  g10559(.A0(new_n6884_), .A1(new_n4427_), .B0(new_n10623_), .Y(new_n10624_));
  AOI21X1  g10560(.A0(new_n7771_), .A1(new_n4080_), .B0(new_n10624_), .Y(new_n10625_));
  XOR2X1   g10561(.A(new_n10625_), .B(\a[11] ), .Y(new_n10626_));
  INVX1    g10562(.A(new_n10490_), .Y(new_n10627_));
  XOR2X1   g10563(.A(new_n10627_), .B(new_n10488_), .Y(new_n10628_));
  NOR2X1   g10564(.A(new_n10628_), .B(new_n10626_), .Y(new_n10629_));
  XOR2X1   g10565(.A(new_n10628_), .B(new_n10626_), .Y(new_n10630_));
  INVX1    g10566(.A(new_n10630_), .Y(new_n10631_));
  AOI22X1  g10567(.A0(new_n6890_), .A1(new_n4078_), .B0(new_n6887_), .B1(new_n4247_), .Y(new_n10632_));
  OAI21X1  g10568(.A0(new_n6886_), .A1(new_n4427_), .B0(new_n10632_), .Y(new_n10633_));
  AOI21X1  g10569(.A0(new_n7762_), .A1(new_n4080_), .B0(new_n10633_), .Y(new_n10634_));
  XOR2X1   g10570(.A(new_n10634_), .B(\a[11] ), .Y(new_n10635_));
  INVX1    g10571(.A(new_n10486_), .Y(new_n10636_));
  XOR2X1   g10572(.A(new_n10636_), .B(new_n10484_), .Y(new_n10637_));
  NOR2X1   g10573(.A(new_n10637_), .B(new_n10635_), .Y(new_n10638_));
  INVX1    g10574(.A(new_n10638_), .Y(new_n10639_));
  XOR2X1   g10575(.A(new_n10637_), .B(new_n10635_), .Y(new_n10640_));
  INVX1    g10576(.A(new_n10640_), .Y(new_n10641_));
  AND2X1   g10577(.A(new_n10482_), .B(new_n10336_), .Y(new_n10642_));
  XOR2X1   g10578(.A(new_n10642_), .B(new_n10328_), .Y(new_n10643_));
  INVX1    g10579(.A(new_n10643_), .Y(new_n10644_));
  OAI22X1  g10580(.A0(new_n8075_), .A1(new_n4077_), .B0(new_n7885_), .B1(new_n4246_), .Y(new_n10645_));
  AOI21X1  g10581(.A0(new_n6887_), .A1(new_n4428_), .B0(new_n10645_), .Y(new_n10646_));
  OAI21X1  g10582(.A0(new_n7876_), .A1(new_n4245_), .B0(new_n10646_), .Y(new_n10647_));
  XOR2X1   g10583(.A(new_n10647_), .B(new_n2911_), .Y(new_n10648_));
  NOR2X1   g10584(.A(new_n10648_), .B(new_n10644_), .Y(new_n10649_));
  XOR2X1   g10585(.A(new_n10481_), .B(new_n10338_), .Y(new_n10650_));
  OAI22X1  g10586(.A0(new_n6896_), .A1(new_n4077_), .B0(new_n8075_), .B1(new_n4246_), .Y(new_n10651_));
  AOI21X1  g10587(.A0(new_n6890_), .A1(new_n4428_), .B0(new_n10651_), .Y(new_n10652_));
  OAI21X1  g10588(.A0(new_n9738_), .A1(new_n4245_), .B0(new_n10652_), .Y(new_n10653_));
  XOR2X1   g10589(.A(new_n10653_), .B(\a[11] ), .Y(new_n10654_));
  AOI22X1  g10590(.A0(new_n6897_), .A1(new_n4078_), .B0(new_n6894_), .B1(new_n4247_), .Y(new_n10655_));
  OAI21X1  g10591(.A0(new_n8075_), .A1(new_n4427_), .B0(new_n10655_), .Y(new_n10656_));
  AOI21X1  g10592(.A0(new_n8074_), .A1(new_n4080_), .B0(new_n10656_), .Y(new_n10657_));
  XOR2X1   g10593(.A(new_n10657_), .B(\a[11] ), .Y(new_n10658_));
  INVX1    g10594(.A(new_n10658_), .Y(new_n10659_));
  XOR2X1   g10595(.A(new_n10480_), .B(new_n10479_), .Y(new_n10660_));
  XOR2X1   g10596(.A(new_n10660_), .B(new_n10658_), .Y(new_n10661_));
  AOI22X1  g10597(.A0(new_n6899_), .A1(new_n4078_), .B0(new_n6897_), .B1(new_n4247_), .Y(new_n10662_));
  OAI21X1  g10598(.A0(new_n6896_), .A1(new_n4427_), .B0(new_n10662_), .Y(new_n10663_));
  AOI21X1  g10599(.A0(new_n7953_), .A1(new_n4080_), .B0(new_n10663_), .Y(new_n10664_));
  XOR2X1   g10600(.A(new_n10664_), .B(\a[11] ), .Y(new_n10665_));
  XOR2X1   g10601(.A(new_n10478_), .B(new_n10475_), .Y(new_n10666_));
  OR2X1    g10602(.A(new_n10666_), .B(new_n10665_), .Y(new_n10667_));
  XOR2X1   g10603(.A(new_n10666_), .B(new_n10665_), .Y(new_n10668_));
  INVX1    g10604(.A(new_n10668_), .Y(new_n10669_));
  AOI22X1  g10605(.A0(new_n6902_), .A1(new_n4078_), .B0(new_n6899_), .B1(new_n4247_), .Y(new_n10670_));
  OAI21X1  g10606(.A0(new_n6898_), .A1(new_n4427_), .B0(new_n10670_), .Y(new_n10671_));
  AOI21X1  g10607(.A0(new_n8215_), .A1(new_n4080_), .B0(new_n10671_), .Y(new_n10672_));
  XOR2X1   g10608(.A(new_n10672_), .B(\a[11] ), .Y(new_n10673_));
  INVX1    g10609(.A(new_n10474_), .Y(new_n10674_));
  XOR2X1   g10610(.A(new_n10674_), .B(new_n10473_), .Y(new_n10675_));
  NOR2X1   g10611(.A(new_n10675_), .B(new_n10673_), .Y(new_n10676_));
  XOR2X1   g10612(.A(new_n10675_), .B(new_n10673_), .Y(new_n10677_));
  XOR2X1   g10613(.A(new_n10471_), .B(new_n10366_), .Y(new_n10678_));
  INVX1    g10614(.A(new_n10678_), .Y(new_n10679_));
  OAI22X1  g10615(.A0(new_n8200_), .A1(new_n4077_), .B0(new_n8205_), .B1(new_n4246_), .Y(new_n10680_));
  AOI21X1  g10616(.A0(new_n6899_), .A1(new_n4428_), .B0(new_n10680_), .Y(new_n10681_));
  OAI21X1  g10617(.A0(new_n8293_), .A1(new_n4245_), .B0(new_n10681_), .Y(new_n10682_));
  XOR2X1   g10618(.A(new_n10682_), .B(new_n2911_), .Y(new_n10683_));
  NOR2X1   g10619(.A(new_n10683_), .B(new_n10679_), .Y(new_n10684_));
  XOR2X1   g10620(.A(new_n10470_), .B(new_n10373_), .Y(new_n10685_));
  OAI22X1  g10621(.A0(new_n6964_), .A1(new_n4077_), .B0(new_n8200_), .B1(new_n4246_), .Y(new_n10686_));
  AOI21X1  g10622(.A0(new_n6902_), .A1(new_n4428_), .B0(new_n10686_), .Y(new_n10687_));
  OAI21X1  g10623(.A0(new_n8203_), .A1(new_n4245_), .B0(new_n10687_), .Y(new_n10688_));
  XOR2X1   g10624(.A(new_n10688_), .B(\a[11] ), .Y(new_n10689_));
  NAND2X1  g10625(.A(new_n10689_), .B(new_n10685_), .Y(new_n10690_));
  XOR2X1   g10626(.A(new_n10469_), .B(new_n10381_), .Y(new_n10691_));
  INVX1    g10627(.A(new_n10691_), .Y(new_n10692_));
  OAI22X1  g10628(.A0(new_n6960_), .A1(new_n4077_), .B0(new_n6964_), .B1(new_n4246_), .Y(new_n10693_));
  AOI21X1  g10629(.A0(new_n6904_), .A1(new_n4428_), .B0(new_n10693_), .Y(new_n10694_));
  OAI21X1  g10630(.A0(new_n8364_), .A1(new_n4245_), .B0(new_n10694_), .Y(new_n10695_));
  XOR2X1   g10631(.A(new_n10695_), .B(new_n2911_), .Y(new_n10696_));
  NOR2X1   g10632(.A(new_n10696_), .B(new_n10692_), .Y(new_n10697_));
  AOI22X1  g10633(.A0(new_n6911_), .A1(new_n4078_), .B0(new_n6909_), .B1(new_n4247_), .Y(new_n10698_));
  OAI21X1  g10634(.A0(new_n6964_), .A1(new_n4427_), .B0(new_n10698_), .Y(new_n10699_));
  AOI21X1  g10635(.A0(new_n8541_), .A1(new_n4080_), .B0(new_n10699_), .Y(new_n10700_));
  XOR2X1   g10636(.A(new_n10700_), .B(\a[11] ), .Y(new_n10701_));
  INVX1    g10637(.A(new_n10701_), .Y(new_n10702_));
  XOR2X1   g10638(.A(new_n10468_), .B(new_n10467_), .Y(new_n10703_));
  NAND2X1  g10639(.A(new_n10703_), .B(new_n10702_), .Y(new_n10704_));
  XOR2X1   g10640(.A(new_n10703_), .B(new_n10701_), .Y(new_n10705_));
  AOI22X1  g10641(.A0(new_n6913_), .A1(new_n4078_), .B0(new_n6911_), .B1(new_n4247_), .Y(new_n10706_));
  OAI21X1  g10642(.A0(new_n6960_), .A1(new_n4427_), .B0(new_n10706_), .Y(new_n10707_));
  AOI21X1  g10643(.A0(new_n8553_), .A1(new_n4080_), .B0(new_n10707_), .Y(new_n10708_));
  XOR2X1   g10644(.A(new_n10708_), .B(\a[11] ), .Y(new_n10709_));
  XOR2X1   g10645(.A(new_n10466_), .B(new_n10464_), .Y(new_n10710_));
  NOR2X1   g10646(.A(new_n10710_), .B(new_n10709_), .Y(new_n10711_));
  XOR2X1   g10647(.A(new_n10710_), .B(new_n10709_), .Y(new_n10712_));
  AOI22X1  g10648(.A0(new_n6915_), .A1(new_n4078_), .B0(new_n6913_), .B1(new_n4247_), .Y(new_n10713_));
  OAI21X1  g10649(.A0(new_n8349_), .A1(new_n4427_), .B0(new_n10713_), .Y(new_n10714_));
  AOI21X1  g10650(.A0(new_n8348_), .A1(new_n4080_), .B0(new_n10714_), .Y(new_n10715_));
  XOR2X1   g10651(.A(new_n10715_), .B(\a[11] ), .Y(new_n10716_));
  XOR2X1   g10652(.A(new_n10463_), .B(new_n10461_), .Y(new_n10717_));
  OR2X1    g10653(.A(new_n10717_), .B(new_n10716_), .Y(new_n10718_));
  XOR2X1   g10654(.A(new_n10717_), .B(new_n10716_), .Y(new_n10719_));
  INVX1    g10655(.A(new_n10719_), .Y(new_n10720_));
  INVX1    g10656(.A(new_n10412_), .Y(new_n10721_));
  XOR2X1   g10657(.A(new_n10460_), .B(new_n10721_), .Y(new_n10722_));
  OAI22X1  g10658(.A0(new_n6918_), .A1(new_n4077_), .B0(new_n6917_), .B1(new_n4246_), .Y(new_n10723_));
  AOI21X1  g10659(.A0(new_n6913_), .A1(new_n4428_), .B0(new_n10723_), .Y(new_n10724_));
  OAI21X1  g10660(.A0(new_n8577_), .A1(new_n4245_), .B0(new_n10724_), .Y(new_n10725_));
  XOR2X1   g10661(.A(new_n10725_), .B(new_n2911_), .Y(new_n10726_));
  NOR2X1   g10662(.A(new_n10726_), .B(new_n10722_), .Y(new_n10727_));
  XOR2X1   g10663(.A(new_n10459_), .B(new_n10458_), .Y(new_n10728_));
  INVX1    g10664(.A(new_n10728_), .Y(new_n10729_));
  OAI22X1  g10665(.A0(new_n6920_), .A1(new_n4077_), .B0(new_n6918_), .B1(new_n4246_), .Y(new_n10730_));
  AOI21X1  g10666(.A0(new_n6915_), .A1(new_n4428_), .B0(new_n10730_), .Y(new_n10731_));
  OAI21X1  g10667(.A0(new_n9093_), .A1(new_n4245_), .B0(new_n10731_), .Y(new_n10732_));
  XOR2X1   g10668(.A(new_n10732_), .B(new_n2911_), .Y(new_n10733_));
  OR2X1    g10669(.A(new_n10733_), .B(new_n10729_), .Y(new_n10734_));
  XOR2X1   g10670(.A(new_n10456_), .B(new_n10429_), .Y(new_n10735_));
  INVX1    g10671(.A(new_n10735_), .Y(new_n10736_));
  OAI22X1  g10672(.A0(new_n8659_), .A1(new_n4077_), .B0(new_n6920_), .B1(new_n4246_), .Y(new_n10737_));
  AOI21X1  g10673(.A0(new_n8580_), .A1(new_n4428_), .B0(new_n10737_), .Y(new_n10738_));
  OAI21X1  g10674(.A0(new_n8611_), .A1(new_n4245_), .B0(new_n10738_), .Y(new_n10739_));
  XOR2X1   g10675(.A(new_n10739_), .B(new_n2911_), .Y(new_n10740_));
  NOR2X1   g10676(.A(new_n10740_), .B(new_n10736_), .Y(new_n10741_));
  INVX1    g10677(.A(new_n10741_), .Y(new_n10742_));
  AOI22X1  g10678(.A0(new_n6925_), .A1(new_n4078_), .B0(new_n6923_), .B1(new_n4247_), .Y(new_n10743_));
  OAI21X1  g10679(.A0(new_n6920_), .A1(new_n4427_), .B0(new_n10743_), .Y(new_n10744_));
  AOI21X1  g10680(.A0(new_n8628_), .A1(new_n4080_), .B0(new_n10744_), .Y(new_n10745_));
  XOR2X1   g10681(.A(new_n10745_), .B(\a[11] ), .Y(new_n10746_));
  INVX1    g10682(.A(new_n10746_), .Y(new_n10747_));
  XOR2X1   g10683(.A(new_n10455_), .B(new_n10454_), .Y(new_n10748_));
  AND2X1   g10684(.A(new_n10748_), .B(new_n10747_), .Y(new_n10749_));
  INVX1    g10685(.A(new_n10749_), .Y(new_n10750_));
  XOR2X1   g10686(.A(new_n10748_), .B(new_n10746_), .Y(new_n10751_));
  XOR2X1   g10687(.A(new_n10452_), .B(new_n2529_), .Y(new_n10752_));
  XOR2X1   g10688(.A(new_n10752_), .B(new_n10449_), .Y(new_n10753_));
  OAI22X1  g10689(.A0(new_n6929_), .A1(new_n4077_), .B0(new_n8683_), .B1(new_n4246_), .Y(new_n10754_));
  AOI21X1  g10690(.A0(new_n6923_), .A1(new_n4428_), .B0(new_n10754_), .Y(new_n10755_));
  OAI21X1  g10691(.A0(new_n8662_), .A1(new_n4245_), .B0(new_n10755_), .Y(new_n10756_));
  XOR2X1   g10692(.A(new_n10756_), .B(new_n2911_), .Y(new_n10757_));
  NOR2X1   g10693(.A(new_n10757_), .B(new_n10753_), .Y(new_n10758_));
  AOI22X1  g10694(.A0(new_n6932_), .A1(new_n4078_), .B0(new_n6927_), .B1(new_n4247_), .Y(new_n10759_));
  OAI21X1  g10695(.A0(new_n8683_), .A1(new_n4427_), .B0(new_n10759_), .Y(new_n10760_));
  AOI21X1  g10696(.A0(new_n8682_), .A1(new_n4080_), .B0(new_n10760_), .Y(new_n10761_));
  XOR2X1   g10697(.A(new_n10761_), .B(\a[11] ), .Y(new_n10762_));
  INVX1    g10698(.A(new_n10762_), .Y(new_n10763_));
  XOR2X1   g10699(.A(new_n10445_), .B(new_n10441_), .Y(new_n10764_));
  AND2X1   g10700(.A(new_n10764_), .B(new_n10763_), .Y(new_n10765_));
  XOR2X1   g10701(.A(new_n10764_), .B(new_n10762_), .Y(new_n10766_));
  NOR2X1   g10702(.A(new_n10439_), .B(new_n2529_), .Y(new_n10767_));
  XOR2X1   g10703(.A(new_n10767_), .B(new_n10447_), .Y(new_n10768_));
  OAI22X1  g10704(.A0(new_n8757_), .A1(new_n4077_), .B0(new_n6930_), .B1(new_n4246_), .Y(new_n10769_));
  AOI21X1  g10705(.A0(new_n6927_), .A1(new_n4428_), .B0(new_n10769_), .Y(new_n10770_));
  OAI21X1  g10706(.A0(new_n8705_), .A1(new_n4245_), .B0(new_n10770_), .Y(new_n10771_));
  XOR2X1   g10707(.A(new_n10771_), .B(new_n2911_), .Y(new_n10772_));
  NOR2X1   g10708(.A(new_n10772_), .B(new_n10768_), .Y(new_n10773_));
  OAI22X1  g10709(.A0(new_n6936_), .A1(new_n4246_), .B0(new_n8752_), .B1(new_n4427_), .Y(new_n10774_));
  AOI21X1  g10710(.A0(new_n8751_), .A1(new_n4080_), .B0(new_n10774_), .Y(new_n10775_));
  XOR2X1   g10711(.A(new_n10775_), .B(\a[11] ), .Y(new_n10776_));
  NOR2X1   g10712(.A(new_n6936_), .B(new_n4073_), .Y(new_n10777_));
  OAI22X1  g10713(.A0(new_n6936_), .A1(new_n4077_), .B0(new_n8752_), .B1(new_n4246_), .Y(new_n10778_));
  AOI21X1  g10714(.A0(new_n6933_), .A1(new_n4428_), .B0(new_n10778_), .Y(new_n10779_));
  OAI21X1  g10715(.A0(new_n8759_), .A1(new_n4245_), .B0(new_n10779_), .Y(new_n10780_));
  OR4X1    g10716(.A(new_n10780_), .B(new_n10777_), .C(new_n10776_), .D(new_n2911_), .Y(new_n10781_));
  OR2X1    g10717(.A(new_n10781_), .B(new_n10440_), .Y(new_n10782_));
  XOR2X1   g10718(.A(new_n10781_), .B(new_n10439_), .Y(new_n10783_));
  AOI22X1  g10719(.A0(new_n6935_), .A1(new_n4078_), .B0(new_n6933_), .B1(new_n4247_), .Y(new_n10784_));
  OAI21X1  g10720(.A0(new_n6930_), .A1(new_n4427_), .B0(new_n10784_), .Y(new_n10785_));
  AOI21X1  g10721(.A0(new_n8717_), .A1(new_n4080_), .B0(new_n10785_), .Y(new_n10786_));
  XOR2X1   g10722(.A(new_n10786_), .B(\a[11] ), .Y(new_n10787_));
  OAI21X1  g10723(.A0(new_n10787_), .A1(new_n10783_), .B0(new_n10782_), .Y(new_n10788_));
  XOR2X1   g10724(.A(new_n10772_), .B(new_n10768_), .Y(new_n10789_));
  AOI21X1  g10725(.A0(new_n10789_), .A1(new_n10788_), .B0(new_n10773_), .Y(new_n10790_));
  NOR2X1   g10726(.A(new_n10790_), .B(new_n10766_), .Y(new_n10791_));
  OR2X1    g10727(.A(new_n10791_), .B(new_n10765_), .Y(new_n10792_));
  XOR2X1   g10728(.A(new_n10757_), .B(new_n10753_), .Y(new_n10793_));
  AOI21X1  g10729(.A0(new_n10793_), .A1(new_n10792_), .B0(new_n10758_), .Y(new_n10794_));
  OAI21X1  g10730(.A0(new_n10794_), .A1(new_n10751_), .B0(new_n10750_), .Y(new_n10795_));
  INVX1    g10731(.A(new_n10795_), .Y(new_n10796_));
  XOR2X1   g10732(.A(new_n10740_), .B(new_n10735_), .Y(new_n10797_));
  OAI21X1  g10733(.A0(new_n10797_), .A1(new_n10796_), .B0(new_n10742_), .Y(new_n10798_));
  INVX1    g10734(.A(new_n10798_), .Y(new_n10799_));
  XOR2X1   g10735(.A(new_n10733_), .B(new_n10728_), .Y(new_n10800_));
  OAI21X1  g10736(.A0(new_n10800_), .A1(new_n10799_), .B0(new_n10734_), .Y(new_n10801_));
  XOR2X1   g10737(.A(new_n10726_), .B(new_n10722_), .Y(new_n10802_));
  AOI21X1  g10738(.A0(new_n10802_), .A1(new_n10801_), .B0(new_n10727_), .Y(new_n10803_));
  OAI21X1  g10739(.A0(new_n10803_), .A1(new_n10720_), .B0(new_n10718_), .Y(new_n10804_));
  AOI21X1  g10740(.A0(new_n10804_), .A1(new_n10712_), .B0(new_n10711_), .Y(new_n10805_));
  OAI21X1  g10741(.A0(new_n10805_), .A1(new_n10705_), .B0(new_n10704_), .Y(new_n10806_));
  XOR2X1   g10742(.A(new_n10696_), .B(new_n10691_), .Y(new_n10807_));
  INVX1    g10743(.A(new_n10807_), .Y(new_n10808_));
  AOI21X1  g10744(.A0(new_n10808_), .A1(new_n10806_), .B0(new_n10697_), .Y(new_n10809_));
  XOR2X1   g10745(.A(new_n10688_), .B(new_n2911_), .Y(new_n10810_));
  XOR2X1   g10746(.A(new_n10810_), .B(new_n10685_), .Y(new_n10811_));
  OAI21X1  g10747(.A0(new_n10811_), .A1(new_n10809_), .B0(new_n10690_), .Y(new_n10812_));
  XOR2X1   g10748(.A(new_n10683_), .B(new_n10679_), .Y(new_n10813_));
  AOI21X1  g10749(.A0(new_n10813_), .A1(new_n10812_), .B0(new_n10684_), .Y(new_n10814_));
  INVX1    g10750(.A(new_n10814_), .Y(new_n10815_));
  AOI21X1  g10751(.A0(new_n10815_), .A1(new_n10677_), .B0(new_n10676_), .Y(new_n10816_));
  OR2X1    g10752(.A(new_n10816_), .B(new_n10669_), .Y(new_n10817_));
  AOI21X1  g10753(.A0(new_n10817_), .A1(new_n10667_), .B0(new_n10661_), .Y(new_n10818_));
  AOI21X1  g10754(.A0(new_n10660_), .A1(new_n10659_), .B0(new_n10818_), .Y(new_n10819_));
  XOR2X1   g10755(.A(new_n10653_), .B(new_n2911_), .Y(new_n10820_));
  XOR2X1   g10756(.A(new_n10820_), .B(new_n10650_), .Y(new_n10821_));
  NOR2X1   g10757(.A(new_n10821_), .B(new_n10819_), .Y(new_n10822_));
  AOI21X1  g10758(.A0(new_n10654_), .A1(new_n10650_), .B0(new_n10822_), .Y(new_n10823_));
  INVX1    g10759(.A(new_n10823_), .Y(new_n10824_));
  XOR2X1   g10760(.A(new_n10648_), .B(new_n10644_), .Y(new_n10825_));
  AOI21X1  g10761(.A0(new_n10825_), .A1(new_n10824_), .B0(new_n10649_), .Y(new_n10826_));
  OR2X1    g10762(.A(new_n10826_), .B(new_n10641_), .Y(new_n10827_));
  AOI21X1  g10763(.A0(new_n10827_), .A1(new_n10639_), .B0(new_n10631_), .Y(new_n10828_));
  NOR2X1   g10764(.A(new_n10828_), .B(new_n10629_), .Y(new_n10829_));
  INVX1    g10765(.A(new_n10829_), .Y(new_n10830_));
  AOI21X1  g10766(.A0(new_n10830_), .A1(new_n10622_), .B0(new_n10621_), .Y(new_n10831_));
  INVX1    g10767(.A(new_n10831_), .Y(new_n10832_));
  AOI21X1  g10768(.A0(new_n10832_), .A1(new_n10615_), .B0(new_n10614_), .Y(new_n10833_));
  INVX1    g10769(.A(new_n10833_), .Y(new_n10834_));
  AOI21X1  g10770(.A0(new_n10834_), .A1(new_n10607_), .B0(new_n10606_), .Y(new_n10835_));
  OR2X1    g10771(.A(new_n10835_), .B(new_n10598_), .Y(new_n10836_));
  OAI21X1  g10772(.A0(new_n10596_), .A1(new_n10594_), .B0(new_n10836_), .Y(new_n10837_));
  AOI21X1  g10773(.A0(new_n10837_), .A1(new_n10590_), .B0(new_n10589_), .Y(new_n10838_));
  OR2X1    g10774(.A(new_n10838_), .B(new_n10583_), .Y(new_n10839_));
  OAI21X1  g10775(.A0(new_n10581_), .A1(new_n10579_), .B0(new_n10839_), .Y(new_n10840_));
  AOI21X1  g10776(.A0(new_n10840_), .A1(new_n10575_), .B0(new_n10574_), .Y(new_n10841_));
  INVX1    g10777(.A(new_n10841_), .Y(new_n10842_));
  AOI21X1  g10778(.A0(new_n10842_), .A1(new_n10568_), .B0(new_n10567_), .Y(new_n10843_));
  AOI21X1  g10779(.A0(new_n10560_), .A1(new_n10559_), .B0(new_n10843_), .Y(new_n10844_));
  NAND3X1  g10780(.A(new_n10843_), .B(new_n10560_), .C(new_n10559_), .Y(new_n10845_));
  AOI22X1  g10781(.A0(new_n7571_), .A1(new_n4870_), .B0(new_n7558_), .B1(new_n4635_), .Y(new_n10846_));
  OAI21X1  g10782(.A0(new_n7602_), .A1(new_n5096_), .B0(new_n10846_), .Y(new_n10847_));
  AOI21X1  g10783(.A0(new_n7601_), .A1(new_n4637_), .B0(new_n10847_), .Y(new_n10848_));
  XOR2X1   g10784(.A(new_n10848_), .B(\a[8] ), .Y(new_n10849_));
  INVX1    g10785(.A(new_n10849_), .Y(new_n10850_));
  AOI21X1  g10786(.A0(new_n10850_), .A1(new_n10845_), .B0(new_n10844_), .Y(new_n10851_));
  AOI21X1  g10787(.A0(new_n10558_), .A1(new_n10556_), .B0(new_n10851_), .Y(new_n10852_));
  NAND3X1  g10788(.A(new_n10851_), .B(new_n10558_), .C(new_n10556_), .Y(new_n10853_));
  AOI22X1  g10789(.A0(new_n7657_), .A1(new_n5373_), .B0(new_n7341_), .B1(new_n5960_), .Y(new_n10854_));
  OAI21X1  g10790(.A0(new_n7644_), .A1(new_n5658_), .B0(new_n10854_), .Y(new_n10855_));
  AOI21X1  g10791(.A0(new_n7656_), .A1(new_n67_), .B0(new_n10855_), .Y(new_n10856_));
  XOR2X1   g10792(.A(new_n10856_), .B(\a[5] ), .Y(new_n10857_));
  INVX1    g10793(.A(new_n10857_), .Y(new_n10858_));
  AOI21X1  g10794(.A0(new_n10858_), .A1(new_n10853_), .B0(new_n10852_), .Y(new_n10859_));
  NOR2X1   g10795(.A(new_n10859_), .B(new_n10546_), .Y(new_n10860_));
  XOR2X1   g10796(.A(new_n10859_), .B(new_n10546_), .Y(new_n10861_));
  NOR3X1   g10797(.A(new_n10532_), .B(new_n10557_), .C(new_n10526_), .Y(new_n10862_));
  AOI21X1  g10798(.A0(new_n10527_), .A1(new_n10555_), .B0(new_n10531_), .Y(new_n10863_));
  NOR3X1   g10799(.A(new_n10524_), .B(new_n10553_), .C(new_n10518_), .Y(new_n10864_));
  AOI21X1  g10800(.A0(new_n10519_), .A1(new_n10552_), .B0(new_n10523_), .Y(new_n10865_));
  INVX1    g10801(.A(new_n10843_), .Y(new_n10866_));
  OAI21X1  g10802(.A0(new_n10865_), .A1(new_n10864_), .B0(new_n10866_), .Y(new_n10867_));
  NOR3X1   g10803(.A(new_n10866_), .B(new_n10865_), .C(new_n10864_), .Y(new_n10868_));
  OAI21X1  g10804(.A0(new_n10849_), .A1(new_n10868_), .B0(new_n10867_), .Y(new_n10869_));
  NOR3X1   g10805(.A(new_n10869_), .B(new_n10863_), .C(new_n10862_), .Y(new_n10870_));
  NOR3X1   g10806(.A(new_n10858_), .B(new_n10870_), .C(new_n10852_), .Y(new_n10871_));
  OAI21X1  g10807(.A0(new_n10863_), .A1(new_n10862_), .B0(new_n10869_), .Y(new_n10872_));
  AOI21X1  g10808(.A0(new_n10853_), .A1(new_n10872_), .B0(new_n10857_), .Y(new_n10873_));
  NOR3X1   g10809(.A(new_n10850_), .B(new_n10868_), .C(new_n10844_), .Y(new_n10874_));
  AOI21X1  g10810(.A0(new_n10845_), .A1(new_n10867_), .B0(new_n10849_), .Y(new_n10875_));
  XOR2X1   g10811(.A(new_n10841_), .B(new_n10568_), .Y(new_n10876_));
  OAI22X1  g10812(.A0(new_n7581_), .A1(new_n4869_), .B0(new_n7537_), .B1(new_n4634_), .Y(new_n10877_));
  AOI21X1  g10813(.A0(new_n7571_), .A1(new_n5097_), .B0(new_n10877_), .Y(new_n10878_));
  OAI21X1  g10814(.A0(new_n7621_), .A1(new_n4868_), .B0(new_n10878_), .Y(new_n10879_));
  XOR2X1   g10815(.A(new_n10879_), .B(new_n2995_), .Y(new_n10880_));
  NOR2X1   g10816(.A(new_n10880_), .B(new_n10876_), .Y(new_n10881_));
  XOR2X1   g10817(.A(new_n10840_), .B(new_n10575_), .Y(new_n10882_));
  OAI22X1  g10818(.A0(new_n7537_), .A1(new_n4869_), .B0(new_n7523_), .B1(new_n4634_), .Y(new_n10883_));
  AOI21X1  g10819(.A0(new_n7558_), .A1(new_n5097_), .B0(new_n10883_), .Y(new_n10884_));
  OAI21X1  g10820(.A0(new_n7566_), .A1(new_n4868_), .B0(new_n10884_), .Y(new_n10885_));
  XOR2X1   g10821(.A(new_n10885_), .B(new_n2995_), .Y(new_n10886_));
  INVX1    g10822(.A(new_n10886_), .Y(new_n10887_));
  NAND2X1  g10823(.A(new_n10887_), .B(new_n10882_), .Y(new_n10888_));
  XOR2X1   g10824(.A(new_n10838_), .B(new_n10582_), .Y(new_n10889_));
  OAI22X1  g10825(.A0(new_n7523_), .A1(new_n4869_), .B0(new_n7504_), .B1(new_n4634_), .Y(new_n10890_));
  AOI21X1  g10826(.A0(new_n7529_), .A1(new_n5097_), .B0(new_n10890_), .Y(new_n10891_));
  OAI21X1  g10827(.A0(new_n7535_), .A1(new_n4868_), .B0(new_n10891_), .Y(new_n10892_));
  XOR2X1   g10828(.A(new_n10892_), .B(new_n2995_), .Y(new_n10893_));
  OR2X1    g10829(.A(new_n10893_), .B(new_n10889_), .Y(new_n10894_));
  INVX1    g10830(.A(new_n10590_), .Y(new_n10895_));
  XOR2X1   g10831(.A(new_n10837_), .B(new_n10895_), .Y(new_n10896_));
  OAI22X1  g10832(.A0(new_n7504_), .A1(new_n4869_), .B0(new_n7367_), .B1(new_n4634_), .Y(new_n10897_));
  AOI21X1  g10833(.A0(new_n7522_), .A1(new_n5097_), .B0(new_n10897_), .Y(new_n10898_));
  OAI21X1  g10834(.A0(new_n7611_), .A1(new_n4868_), .B0(new_n10898_), .Y(new_n10899_));
  XOR2X1   g10835(.A(new_n10899_), .B(new_n2995_), .Y(new_n10900_));
  NOR2X1   g10836(.A(new_n10900_), .B(new_n10896_), .Y(new_n10901_));
  XOR2X1   g10837(.A(new_n10835_), .B(new_n10597_), .Y(new_n10902_));
  OAI22X1  g10838(.A0(new_n7367_), .A1(new_n4869_), .B0(new_n7047_), .B1(new_n4634_), .Y(new_n10903_));
  AOI21X1  g10839(.A0(new_n7485_), .A1(new_n5097_), .B0(new_n10903_), .Y(new_n10904_));
  OAI21X1  g10840(.A0(new_n7495_), .A1(new_n4868_), .B0(new_n10904_), .Y(new_n10905_));
  XOR2X1   g10841(.A(new_n10905_), .B(new_n2995_), .Y(new_n10906_));
  OR2X1    g10842(.A(new_n10906_), .B(new_n10902_), .Y(new_n10907_));
  XOR2X1   g10843(.A(new_n10833_), .B(new_n10607_), .Y(new_n10908_));
  AOI22X1  g10844(.A0(new_n7044_), .A1(new_n4870_), .B0(new_n6818_), .B1(new_n4635_), .Y(new_n10909_));
  OAI21X1  g10845(.A0(new_n7367_), .A1(new_n5096_), .B0(new_n10909_), .Y(new_n10910_));
  AOI21X1  g10846(.A0(new_n7366_), .A1(new_n4637_), .B0(new_n10910_), .Y(new_n10911_));
  XOR2X1   g10847(.A(new_n10911_), .B(\a[8] ), .Y(new_n10912_));
  NOR2X1   g10848(.A(new_n10912_), .B(new_n10908_), .Y(new_n10913_));
  XOR2X1   g10849(.A(new_n10832_), .B(new_n10615_), .Y(new_n10914_));
  OAI22X1  g10850(.A0(new_n7361_), .A1(new_n4869_), .B0(new_n7418_), .B1(new_n4634_), .Y(new_n10915_));
  AOI21X1  g10851(.A0(new_n7044_), .A1(new_n5097_), .B0(new_n10915_), .Y(new_n10916_));
  OAI21X1  g10852(.A0(new_n7680_), .A1(new_n4868_), .B0(new_n10916_), .Y(new_n10917_));
  XOR2X1   g10853(.A(new_n10917_), .B(\a[8] ), .Y(new_n10918_));
  NAND2X1  g10854(.A(new_n10918_), .B(new_n10914_), .Y(new_n10919_));
  XOR2X1   g10855(.A(new_n10829_), .B(new_n10622_), .Y(new_n10920_));
  OAI22X1  g10856(.A0(new_n7671_), .A1(new_n4634_), .B0(new_n7418_), .B1(new_n4869_), .Y(new_n10921_));
  AOI21X1  g10857(.A0(new_n6818_), .A1(new_n5097_), .B0(new_n10921_), .Y(new_n10922_));
  OAI21X1  g10858(.A0(new_n7403_), .A1(new_n4868_), .B0(new_n10922_), .Y(new_n10923_));
  XOR2X1   g10859(.A(new_n10923_), .B(new_n2995_), .Y(new_n10924_));
  NOR2X1   g10860(.A(new_n10924_), .B(new_n10920_), .Y(new_n10925_));
  INVX1    g10861(.A(new_n10925_), .Y(new_n10926_));
  AND2X1   g10862(.A(new_n10827_), .B(new_n10639_), .Y(new_n10927_));
  XOR2X1   g10863(.A(new_n10927_), .B(new_n10631_), .Y(new_n10928_));
  OAI22X1  g10864(.A0(new_n7472_), .A1(new_n4634_), .B0(new_n7671_), .B1(new_n4869_), .Y(new_n10929_));
  AOI21X1  g10865(.A0(new_n6745_), .A1(new_n5097_), .B0(new_n10929_), .Y(new_n10930_));
  OAI21X1  g10866(.A0(new_n7416_), .A1(new_n4868_), .B0(new_n10930_), .Y(new_n10931_));
  XOR2X1   g10867(.A(new_n10931_), .B(\a[8] ), .Y(new_n10932_));
  AND2X1   g10868(.A(new_n10932_), .B(new_n10928_), .Y(new_n10933_));
  XOR2X1   g10869(.A(new_n10826_), .B(new_n10641_), .Y(new_n10934_));
  INVX1    g10870(.A(new_n10934_), .Y(new_n10935_));
  OAI22X1  g10871(.A0(new_n6884_), .A1(new_n4634_), .B0(new_n7472_), .B1(new_n4869_), .Y(new_n10936_));
  AOI21X1  g10872(.A0(new_n6820_), .A1(new_n5097_), .B0(new_n10936_), .Y(new_n10937_));
  OAI21X1  g10873(.A0(new_n10280_), .A1(new_n4868_), .B0(new_n10937_), .Y(new_n10938_));
  XOR2X1   g10874(.A(new_n10938_), .B(new_n2995_), .Y(new_n10939_));
  AOI22X1  g10875(.A0(new_n6885_), .A1(new_n4635_), .B0(new_n6882_), .B1(new_n4870_), .Y(new_n10940_));
  OAI21X1  g10876(.A0(new_n7472_), .A1(new_n5096_), .B0(new_n10940_), .Y(new_n10941_));
  AOI21X1  g10877(.A0(new_n7471_), .A1(new_n4637_), .B0(new_n10941_), .Y(new_n10942_));
  XOR2X1   g10878(.A(new_n10942_), .B(\a[8] ), .Y(new_n10943_));
  XOR2X1   g10879(.A(new_n10825_), .B(new_n10823_), .Y(new_n10944_));
  NOR2X1   g10880(.A(new_n10944_), .B(new_n10943_), .Y(new_n10945_));
  INVX1    g10881(.A(new_n10943_), .Y(new_n10946_));
  XOR2X1   g10882(.A(new_n10944_), .B(new_n10946_), .Y(new_n10947_));
  AOI22X1  g10883(.A0(new_n6887_), .A1(new_n4635_), .B0(new_n6885_), .B1(new_n4870_), .Y(new_n10948_));
  OAI21X1  g10884(.A0(new_n6884_), .A1(new_n5096_), .B0(new_n10948_), .Y(new_n10949_));
  AOI21X1  g10885(.A0(new_n7771_), .A1(new_n4637_), .B0(new_n10949_), .Y(new_n10950_));
  XOR2X1   g10886(.A(new_n10950_), .B(\a[8] ), .Y(new_n10951_));
  INVX1    g10887(.A(new_n10821_), .Y(new_n10952_));
  XOR2X1   g10888(.A(new_n10952_), .B(new_n10819_), .Y(new_n10953_));
  NOR2X1   g10889(.A(new_n10953_), .B(new_n10951_), .Y(new_n10954_));
  INVX1    g10890(.A(new_n10954_), .Y(new_n10955_));
  XOR2X1   g10891(.A(new_n10953_), .B(new_n10951_), .Y(new_n10956_));
  INVX1    g10892(.A(new_n10956_), .Y(new_n10957_));
  AND2X1   g10893(.A(new_n10817_), .B(new_n10667_), .Y(new_n10958_));
  XOR2X1   g10894(.A(new_n10958_), .B(new_n10661_), .Y(new_n10959_));
  INVX1    g10895(.A(new_n10959_), .Y(new_n10960_));
  OAI22X1  g10896(.A0(new_n7885_), .A1(new_n4634_), .B0(new_n7878_), .B1(new_n4869_), .Y(new_n10961_));
  AOI21X1  g10897(.A0(new_n6885_), .A1(new_n5097_), .B0(new_n10961_), .Y(new_n10962_));
  OAI21X1  g10898(.A0(new_n8083_), .A1(new_n4868_), .B0(new_n10962_), .Y(new_n10963_));
  XOR2X1   g10899(.A(new_n10963_), .B(new_n2995_), .Y(new_n10964_));
  NOR2X1   g10900(.A(new_n10964_), .B(new_n10960_), .Y(new_n10965_));
  XOR2X1   g10901(.A(new_n10816_), .B(new_n10669_), .Y(new_n10966_));
  OAI22X1  g10902(.A0(new_n8075_), .A1(new_n4634_), .B0(new_n7885_), .B1(new_n4869_), .Y(new_n10967_));
  AOI21X1  g10903(.A0(new_n6887_), .A1(new_n5097_), .B0(new_n10967_), .Y(new_n10968_));
  OAI21X1  g10904(.A0(new_n7876_), .A1(new_n4868_), .B0(new_n10968_), .Y(new_n10969_));
  XOR2X1   g10905(.A(new_n10969_), .B(\a[8] ), .Y(new_n10970_));
  XOR2X1   g10906(.A(new_n10815_), .B(new_n10677_), .Y(new_n10971_));
  OAI22X1  g10907(.A0(new_n6896_), .A1(new_n4634_), .B0(new_n8075_), .B1(new_n4869_), .Y(new_n10972_));
  AOI21X1  g10908(.A0(new_n6890_), .A1(new_n5097_), .B0(new_n10972_), .Y(new_n10973_));
  OAI21X1  g10909(.A0(new_n9738_), .A1(new_n4868_), .B0(new_n10973_), .Y(new_n10974_));
  XOR2X1   g10910(.A(new_n10974_), .B(\a[8] ), .Y(new_n10975_));
  AND2X1   g10911(.A(new_n10975_), .B(new_n10971_), .Y(new_n10976_));
  AOI22X1  g10912(.A0(new_n6897_), .A1(new_n4635_), .B0(new_n6894_), .B1(new_n4870_), .Y(new_n10977_));
  OAI21X1  g10913(.A0(new_n8075_), .A1(new_n5096_), .B0(new_n10977_), .Y(new_n10978_));
  AOI21X1  g10914(.A0(new_n8074_), .A1(new_n4637_), .B0(new_n10978_), .Y(new_n10979_));
  XOR2X1   g10915(.A(new_n10979_), .B(\a[8] ), .Y(new_n10980_));
  XOR2X1   g10916(.A(new_n10813_), .B(new_n10812_), .Y(new_n10981_));
  INVX1    g10917(.A(new_n10981_), .Y(new_n10982_));
  OR2X1    g10918(.A(new_n10982_), .B(new_n10980_), .Y(new_n10983_));
  XOR2X1   g10919(.A(new_n10981_), .B(new_n10980_), .Y(new_n10984_));
  AOI22X1  g10920(.A0(new_n6899_), .A1(new_n4635_), .B0(new_n6897_), .B1(new_n4870_), .Y(new_n10985_));
  OAI21X1  g10921(.A0(new_n6896_), .A1(new_n5096_), .B0(new_n10985_), .Y(new_n10986_));
  AOI21X1  g10922(.A0(new_n7953_), .A1(new_n4637_), .B0(new_n10986_), .Y(new_n10987_));
  XOR2X1   g10923(.A(new_n10987_), .B(\a[8] ), .Y(new_n10988_));
  INVX1    g10924(.A(new_n10811_), .Y(new_n10989_));
  XOR2X1   g10925(.A(new_n10989_), .B(new_n10809_), .Y(new_n10990_));
  OR2X1    g10926(.A(new_n10990_), .B(new_n10988_), .Y(new_n10991_));
  XOR2X1   g10927(.A(new_n10990_), .B(new_n10988_), .Y(new_n10992_));
  INVX1    g10928(.A(new_n10992_), .Y(new_n10993_));
  AOI22X1  g10929(.A0(new_n6902_), .A1(new_n4635_), .B0(new_n6899_), .B1(new_n4870_), .Y(new_n10994_));
  OAI21X1  g10930(.A0(new_n6898_), .A1(new_n5096_), .B0(new_n10994_), .Y(new_n10995_));
  AOI21X1  g10931(.A0(new_n8215_), .A1(new_n4637_), .B0(new_n10995_), .Y(new_n10996_));
  XOR2X1   g10932(.A(new_n10996_), .B(\a[8] ), .Y(new_n10997_));
  XOR2X1   g10933(.A(new_n10807_), .B(new_n10806_), .Y(new_n10998_));
  NOR2X1   g10934(.A(new_n10998_), .B(new_n10997_), .Y(new_n10999_));
  XOR2X1   g10935(.A(new_n10998_), .B(new_n10997_), .Y(new_n11000_));
  INVX1    g10936(.A(new_n10705_), .Y(new_n11001_));
  XOR2X1   g10937(.A(new_n10805_), .B(new_n11001_), .Y(new_n11002_));
  OAI22X1  g10938(.A0(new_n8200_), .A1(new_n4634_), .B0(new_n8205_), .B1(new_n4869_), .Y(new_n11003_));
  AOI21X1  g10939(.A0(new_n6899_), .A1(new_n5097_), .B0(new_n11003_), .Y(new_n11004_));
  OAI21X1  g10940(.A0(new_n8293_), .A1(new_n4868_), .B0(new_n11004_), .Y(new_n11005_));
  XOR2X1   g10941(.A(new_n11005_), .B(new_n2995_), .Y(new_n11006_));
  NOR2X1   g10942(.A(new_n11006_), .B(new_n11002_), .Y(new_n11007_));
  XOR2X1   g10943(.A(new_n10804_), .B(new_n10712_), .Y(new_n11008_));
  OAI22X1  g10944(.A0(new_n6964_), .A1(new_n4634_), .B0(new_n8200_), .B1(new_n4869_), .Y(new_n11009_));
  AOI21X1  g10945(.A0(new_n6902_), .A1(new_n5097_), .B0(new_n11009_), .Y(new_n11010_));
  OAI21X1  g10946(.A0(new_n8203_), .A1(new_n4868_), .B0(new_n11010_), .Y(new_n11011_));
  XOR2X1   g10947(.A(new_n11011_), .B(new_n2995_), .Y(new_n11012_));
  INVX1    g10948(.A(new_n11012_), .Y(new_n11013_));
  NAND2X1  g10949(.A(new_n11013_), .B(new_n11008_), .Y(new_n11014_));
  XOR2X1   g10950(.A(new_n10803_), .B(new_n10720_), .Y(new_n11015_));
  INVX1    g10951(.A(new_n11015_), .Y(new_n11016_));
  OAI22X1  g10952(.A0(new_n6960_), .A1(new_n4634_), .B0(new_n6964_), .B1(new_n4869_), .Y(new_n11017_));
  AOI21X1  g10953(.A0(new_n6904_), .A1(new_n5097_), .B0(new_n11017_), .Y(new_n11018_));
  OAI21X1  g10954(.A0(new_n8364_), .A1(new_n4868_), .B0(new_n11018_), .Y(new_n11019_));
  XOR2X1   g10955(.A(new_n11019_), .B(new_n2995_), .Y(new_n11020_));
  NOR2X1   g10956(.A(new_n11020_), .B(new_n11016_), .Y(new_n11021_));
  AOI22X1  g10957(.A0(new_n6911_), .A1(new_n4635_), .B0(new_n6909_), .B1(new_n4870_), .Y(new_n11022_));
  OAI21X1  g10958(.A0(new_n6964_), .A1(new_n5096_), .B0(new_n11022_), .Y(new_n11023_));
  AOI21X1  g10959(.A0(new_n8541_), .A1(new_n4637_), .B0(new_n11023_), .Y(new_n11024_));
  XOR2X1   g10960(.A(new_n11024_), .B(\a[8] ), .Y(new_n11025_));
  INVX1    g10961(.A(new_n11025_), .Y(new_n11026_));
  XOR2X1   g10962(.A(new_n10802_), .B(new_n10801_), .Y(new_n11027_));
  NAND2X1  g10963(.A(new_n11027_), .B(new_n11026_), .Y(new_n11028_));
  XOR2X1   g10964(.A(new_n11027_), .B(new_n11025_), .Y(new_n11029_));
  AOI22X1  g10965(.A0(new_n6913_), .A1(new_n4635_), .B0(new_n6911_), .B1(new_n4870_), .Y(new_n11030_));
  OAI21X1  g10966(.A0(new_n6960_), .A1(new_n5096_), .B0(new_n11030_), .Y(new_n11031_));
  AOI21X1  g10967(.A0(new_n8553_), .A1(new_n4637_), .B0(new_n11031_), .Y(new_n11032_));
  XOR2X1   g10968(.A(new_n11032_), .B(\a[8] ), .Y(new_n11033_));
  XOR2X1   g10969(.A(new_n10800_), .B(new_n10798_), .Y(new_n11034_));
  NOR2X1   g10970(.A(new_n11034_), .B(new_n11033_), .Y(new_n11035_));
  XOR2X1   g10971(.A(new_n11034_), .B(new_n11033_), .Y(new_n11036_));
  AOI22X1  g10972(.A0(new_n6915_), .A1(new_n4635_), .B0(new_n6913_), .B1(new_n4870_), .Y(new_n11037_));
  OAI21X1  g10973(.A0(new_n8349_), .A1(new_n5096_), .B0(new_n11037_), .Y(new_n11038_));
  AOI21X1  g10974(.A0(new_n8348_), .A1(new_n4637_), .B0(new_n11038_), .Y(new_n11039_));
  XOR2X1   g10975(.A(new_n11039_), .B(\a[8] ), .Y(new_n11040_));
  XOR2X1   g10976(.A(new_n10797_), .B(new_n10795_), .Y(new_n11041_));
  XOR2X1   g10977(.A(new_n11041_), .B(new_n11040_), .Y(new_n11042_));
  INVX1    g10978(.A(new_n11042_), .Y(new_n11043_));
  INVX1    g10979(.A(new_n10751_), .Y(new_n11044_));
  XOR2X1   g10980(.A(new_n10794_), .B(new_n11044_), .Y(new_n11045_));
  OAI22X1  g10981(.A0(new_n6918_), .A1(new_n4634_), .B0(new_n6917_), .B1(new_n4869_), .Y(new_n11046_));
  AOI21X1  g10982(.A0(new_n6913_), .A1(new_n5097_), .B0(new_n11046_), .Y(new_n11047_));
  OAI21X1  g10983(.A0(new_n8577_), .A1(new_n4868_), .B0(new_n11047_), .Y(new_n11048_));
  XOR2X1   g10984(.A(new_n11048_), .B(new_n2995_), .Y(new_n11049_));
  NOR2X1   g10985(.A(new_n11049_), .B(new_n11045_), .Y(new_n11050_));
  XOR2X1   g10986(.A(new_n10793_), .B(new_n10792_), .Y(new_n11051_));
  INVX1    g10987(.A(new_n11051_), .Y(new_n11052_));
  OAI22X1  g10988(.A0(new_n6920_), .A1(new_n4634_), .B0(new_n6918_), .B1(new_n4869_), .Y(new_n11053_));
  AOI21X1  g10989(.A0(new_n6915_), .A1(new_n5097_), .B0(new_n11053_), .Y(new_n11054_));
  OAI21X1  g10990(.A0(new_n9093_), .A1(new_n4868_), .B0(new_n11054_), .Y(new_n11055_));
  XOR2X1   g10991(.A(new_n11055_), .B(new_n2995_), .Y(new_n11056_));
  OR2X1    g10992(.A(new_n11056_), .B(new_n11052_), .Y(new_n11057_));
  XOR2X1   g10993(.A(new_n10790_), .B(new_n10766_), .Y(new_n11058_));
  INVX1    g10994(.A(new_n11058_), .Y(new_n11059_));
  OAI22X1  g10995(.A0(new_n8659_), .A1(new_n4634_), .B0(new_n6920_), .B1(new_n4869_), .Y(new_n11060_));
  AOI21X1  g10996(.A0(new_n8580_), .A1(new_n5097_), .B0(new_n11060_), .Y(new_n11061_));
  OAI21X1  g10997(.A0(new_n8611_), .A1(new_n4868_), .B0(new_n11061_), .Y(new_n11062_));
  XOR2X1   g10998(.A(new_n11062_), .B(new_n2995_), .Y(new_n11063_));
  NOR2X1   g10999(.A(new_n11063_), .B(new_n11059_), .Y(new_n11064_));
  INVX1    g11000(.A(new_n11064_), .Y(new_n11065_));
  AOI22X1  g11001(.A0(new_n6925_), .A1(new_n4635_), .B0(new_n6923_), .B1(new_n4870_), .Y(new_n11066_));
  OAI21X1  g11002(.A0(new_n6920_), .A1(new_n5096_), .B0(new_n11066_), .Y(new_n11067_));
  AOI21X1  g11003(.A0(new_n8628_), .A1(new_n4637_), .B0(new_n11067_), .Y(new_n11068_));
  XOR2X1   g11004(.A(new_n11068_), .B(\a[8] ), .Y(new_n11069_));
  INVX1    g11005(.A(new_n11069_), .Y(new_n11070_));
  XOR2X1   g11006(.A(new_n10789_), .B(new_n10788_), .Y(new_n11071_));
  AND2X1   g11007(.A(new_n11071_), .B(new_n11070_), .Y(new_n11072_));
  INVX1    g11008(.A(new_n11072_), .Y(new_n11073_));
  XOR2X1   g11009(.A(new_n11071_), .B(new_n11069_), .Y(new_n11074_));
  XOR2X1   g11010(.A(new_n10786_), .B(new_n2911_), .Y(new_n11075_));
  XOR2X1   g11011(.A(new_n11075_), .B(new_n10783_), .Y(new_n11076_));
  OAI22X1  g11012(.A0(new_n6929_), .A1(new_n4634_), .B0(new_n8683_), .B1(new_n4869_), .Y(new_n11077_));
  AOI21X1  g11013(.A0(new_n6923_), .A1(new_n5097_), .B0(new_n11077_), .Y(new_n11078_));
  OAI21X1  g11014(.A0(new_n8662_), .A1(new_n4868_), .B0(new_n11078_), .Y(new_n11079_));
  XOR2X1   g11015(.A(new_n11079_), .B(new_n2995_), .Y(new_n11080_));
  NOR2X1   g11016(.A(new_n11080_), .B(new_n11076_), .Y(new_n11081_));
  AOI22X1  g11017(.A0(new_n6932_), .A1(new_n4635_), .B0(new_n6927_), .B1(new_n4870_), .Y(new_n11082_));
  OAI21X1  g11018(.A0(new_n8683_), .A1(new_n5096_), .B0(new_n11082_), .Y(new_n11083_));
  AOI21X1  g11019(.A0(new_n8682_), .A1(new_n4637_), .B0(new_n11083_), .Y(new_n11084_));
  XOR2X1   g11020(.A(new_n11084_), .B(\a[8] ), .Y(new_n11085_));
  INVX1    g11021(.A(new_n11085_), .Y(new_n11086_));
  NOR3X1   g11022(.A(new_n10777_), .B(new_n10776_), .C(new_n2911_), .Y(new_n11087_));
  XOR2X1   g11023(.A(new_n10780_), .B(\a[11] ), .Y(new_n11088_));
  XOR2X1   g11024(.A(new_n11088_), .B(new_n11087_), .Y(new_n11089_));
  AND2X1   g11025(.A(new_n11089_), .B(new_n11086_), .Y(new_n11090_));
  INVX1    g11026(.A(new_n11090_), .Y(new_n11091_));
  XOR2X1   g11027(.A(new_n11089_), .B(new_n11085_), .Y(new_n11092_));
  NOR2X1   g11028(.A(new_n10777_), .B(new_n2911_), .Y(new_n11093_));
  XOR2X1   g11029(.A(new_n11093_), .B(new_n10776_), .Y(new_n11094_));
  OAI22X1  g11030(.A0(new_n8757_), .A1(new_n4634_), .B0(new_n6930_), .B1(new_n4869_), .Y(new_n11095_));
  AOI21X1  g11031(.A0(new_n6927_), .A1(new_n5097_), .B0(new_n11095_), .Y(new_n11096_));
  OAI21X1  g11032(.A0(new_n8705_), .A1(new_n4868_), .B0(new_n11096_), .Y(new_n11097_));
  XOR2X1   g11033(.A(new_n11097_), .B(new_n2995_), .Y(new_n11098_));
  NOR2X1   g11034(.A(new_n11098_), .B(new_n11094_), .Y(new_n11099_));
  OAI22X1  g11035(.A0(new_n6936_), .A1(new_n4869_), .B0(new_n8752_), .B1(new_n5096_), .Y(new_n11100_));
  AOI21X1  g11036(.A0(new_n8751_), .A1(new_n4637_), .B0(new_n11100_), .Y(new_n11101_));
  NOR2X1   g11037(.A(new_n6936_), .B(new_n4630_), .Y(new_n11102_));
  INVX1    g11038(.A(new_n11102_), .Y(new_n11103_));
  NAND3X1  g11039(.A(new_n11103_), .B(new_n11101_), .C(\a[8] ), .Y(new_n11104_));
  OAI22X1  g11040(.A0(new_n6936_), .A1(new_n4634_), .B0(new_n8752_), .B1(new_n4869_), .Y(new_n11105_));
  AOI21X1  g11041(.A0(new_n6933_), .A1(new_n5097_), .B0(new_n11105_), .Y(new_n11106_));
  OAI21X1  g11042(.A0(new_n8759_), .A1(new_n4868_), .B0(new_n11106_), .Y(new_n11107_));
  XOR2X1   g11043(.A(new_n11107_), .B(new_n2995_), .Y(new_n11108_));
  OR4X1    g11044(.A(new_n11108_), .B(new_n11104_), .C(new_n6936_), .D(new_n4073_), .Y(new_n11109_));
  XOR2X1   g11045(.A(new_n11101_), .B(\a[8] ), .Y(new_n11110_));
  OR4X1    g11046(.A(new_n11107_), .B(new_n11102_), .C(new_n11110_), .D(new_n2995_), .Y(new_n11111_));
  XOR2X1   g11047(.A(new_n11111_), .B(new_n10777_), .Y(new_n11112_));
  AOI22X1  g11048(.A0(new_n6935_), .A1(new_n4635_), .B0(new_n6933_), .B1(new_n4870_), .Y(new_n11113_));
  OAI21X1  g11049(.A0(new_n6930_), .A1(new_n5096_), .B0(new_n11113_), .Y(new_n11114_));
  AOI21X1  g11050(.A0(new_n8717_), .A1(new_n4637_), .B0(new_n11114_), .Y(new_n11115_));
  XOR2X1   g11051(.A(new_n11115_), .B(\a[8] ), .Y(new_n11116_));
  OAI21X1  g11052(.A0(new_n11116_), .A1(new_n11112_), .B0(new_n11109_), .Y(new_n11117_));
  XOR2X1   g11053(.A(new_n11098_), .B(new_n11094_), .Y(new_n11118_));
  AOI21X1  g11054(.A0(new_n11118_), .A1(new_n11117_), .B0(new_n11099_), .Y(new_n11119_));
  OR2X1    g11055(.A(new_n11119_), .B(new_n11092_), .Y(new_n11120_));
  AND2X1   g11056(.A(new_n11120_), .B(new_n11091_), .Y(new_n11121_));
  INVX1    g11057(.A(new_n11121_), .Y(new_n11122_));
  XOR2X1   g11058(.A(new_n11080_), .B(new_n11076_), .Y(new_n11123_));
  AOI21X1  g11059(.A0(new_n11123_), .A1(new_n11122_), .B0(new_n11081_), .Y(new_n11124_));
  OAI21X1  g11060(.A0(new_n11124_), .A1(new_n11074_), .B0(new_n11073_), .Y(new_n11125_));
  INVX1    g11061(.A(new_n11125_), .Y(new_n11126_));
  XOR2X1   g11062(.A(new_n11063_), .B(new_n11058_), .Y(new_n11127_));
  OAI21X1  g11063(.A0(new_n11127_), .A1(new_n11126_), .B0(new_n11065_), .Y(new_n11128_));
  INVX1    g11064(.A(new_n11128_), .Y(new_n11129_));
  XOR2X1   g11065(.A(new_n11056_), .B(new_n11051_), .Y(new_n11130_));
  OAI21X1  g11066(.A0(new_n11130_), .A1(new_n11129_), .B0(new_n11057_), .Y(new_n11131_));
  XOR2X1   g11067(.A(new_n11049_), .B(new_n11045_), .Y(new_n11132_));
  AOI21X1  g11068(.A0(new_n11132_), .A1(new_n11131_), .B0(new_n11050_), .Y(new_n11133_));
  OR2X1    g11069(.A(new_n11133_), .B(new_n11043_), .Y(new_n11134_));
  OAI21X1  g11070(.A0(new_n11041_), .A1(new_n11040_), .B0(new_n11134_), .Y(new_n11135_));
  AOI21X1  g11071(.A0(new_n11135_), .A1(new_n11036_), .B0(new_n11035_), .Y(new_n11136_));
  OAI21X1  g11072(.A0(new_n11136_), .A1(new_n11029_), .B0(new_n11028_), .Y(new_n11137_));
  XOR2X1   g11073(.A(new_n11020_), .B(new_n11015_), .Y(new_n11138_));
  INVX1    g11074(.A(new_n11138_), .Y(new_n11139_));
  AOI21X1  g11075(.A0(new_n11139_), .A1(new_n11137_), .B0(new_n11021_), .Y(new_n11140_));
  XOR2X1   g11076(.A(new_n11012_), .B(new_n11008_), .Y(new_n11141_));
  OAI21X1  g11077(.A0(new_n11141_), .A1(new_n11140_), .B0(new_n11014_), .Y(new_n11142_));
  XOR2X1   g11078(.A(new_n11006_), .B(new_n11002_), .Y(new_n11143_));
  AOI21X1  g11079(.A0(new_n11143_), .A1(new_n11142_), .B0(new_n11007_), .Y(new_n11144_));
  INVX1    g11080(.A(new_n11144_), .Y(new_n11145_));
  AOI21X1  g11081(.A0(new_n11145_), .A1(new_n11000_), .B0(new_n10999_), .Y(new_n11146_));
  OR2X1    g11082(.A(new_n11146_), .B(new_n10993_), .Y(new_n11147_));
  AND2X1   g11083(.A(new_n11147_), .B(new_n10991_), .Y(new_n11148_));
  OAI21X1  g11084(.A0(new_n11148_), .A1(new_n10984_), .B0(new_n10983_), .Y(new_n11149_));
  XOR2X1   g11085(.A(new_n10974_), .B(new_n2995_), .Y(new_n11150_));
  XOR2X1   g11086(.A(new_n11150_), .B(new_n10971_), .Y(new_n11151_));
  INVX1    g11087(.A(new_n11151_), .Y(new_n11152_));
  AOI21X1  g11088(.A0(new_n11152_), .A1(new_n11149_), .B0(new_n10976_), .Y(new_n11153_));
  XOR2X1   g11089(.A(new_n10969_), .B(new_n2995_), .Y(new_n11154_));
  XOR2X1   g11090(.A(new_n11154_), .B(new_n10966_), .Y(new_n11155_));
  NOR2X1   g11091(.A(new_n11155_), .B(new_n11153_), .Y(new_n11156_));
  AOI21X1  g11092(.A0(new_n10970_), .A1(new_n10966_), .B0(new_n11156_), .Y(new_n11157_));
  INVX1    g11093(.A(new_n11157_), .Y(new_n11158_));
  XOR2X1   g11094(.A(new_n10964_), .B(new_n10960_), .Y(new_n11159_));
  AOI21X1  g11095(.A0(new_n11159_), .A1(new_n11158_), .B0(new_n10965_), .Y(new_n11160_));
  OR2X1    g11096(.A(new_n11160_), .B(new_n10957_), .Y(new_n11161_));
  AOI21X1  g11097(.A0(new_n11161_), .A1(new_n10955_), .B0(new_n10947_), .Y(new_n11162_));
  XOR2X1   g11098(.A(new_n10939_), .B(new_n10934_), .Y(new_n11163_));
  INVX1    g11099(.A(new_n11163_), .Y(new_n11164_));
  OAI21X1  g11100(.A0(new_n11162_), .A1(new_n10945_), .B0(new_n11164_), .Y(new_n11165_));
  OAI21X1  g11101(.A0(new_n10939_), .A1(new_n10935_), .B0(new_n11165_), .Y(new_n11166_));
  XOR2X1   g11102(.A(new_n10931_), .B(new_n2995_), .Y(new_n11167_));
  XOR2X1   g11103(.A(new_n11167_), .B(new_n10928_), .Y(new_n11168_));
  INVX1    g11104(.A(new_n11168_), .Y(new_n11169_));
  AOI21X1  g11105(.A0(new_n11169_), .A1(new_n11166_), .B0(new_n10933_), .Y(new_n11170_));
  XOR2X1   g11106(.A(new_n10924_), .B(new_n10920_), .Y(new_n11171_));
  INVX1    g11107(.A(new_n11171_), .Y(new_n11172_));
  OAI21X1  g11108(.A0(new_n11172_), .A1(new_n11170_), .B0(new_n10926_), .Y(new_n11173_));
  INVX1    g11109(.A(new_n11173_), .Y(new_n11174_));
  XOR2X1   g11110(.A(new_n10917_), .B(new_n2995_), .Y(new_n11175_));
  XOR2X1   g11111(.A(new_n11175_), .B(new_n10914_), .Y(new_n11176_));
  OAI21X1  g11112(.A0(new_n11176_), .A1(new_n11174_), .B0(new_n10919_), .Y(new_n11177_));
  XOR2X1   g11113(.A(new_n10912_), .B(new_n10908_), .Y(new_n11178_));
  AOI21X1  g11114(.A0(new_n11178_), .A1(new_n11177_), .B0(new_n10913_), .Y(new_n11179_));
  XOR2X1   g11115(.A(new_n10835_), .B(new_n10598_), .Y(new_n11180_));
  XOR2X1   g11116(.A(new_n10906_), .B(new_n11180_), .Y(new_n11181_));
  OAI21X1  g11117(.A0(new_n11181_), .A1(new_n11179_), .B0(new_n10907_), .Y(new_n11182_));
  XOR2X1   g11118(.A(new_n10900_), .B(new_n10896_), .Y(new_n11183_));
  AOI21X1  g11119(.A0(new_n11183_), .A1(new_n11182_), .B0(new_n10901_), .Y(new_n11184_));
  XOR2X1   g11120(.A(new_n10838_), .B(new_n10583_), .Y(new_n11185_));
  XOR2X1   g11121(.A(new_n10893_), .B(new_n11185_), .Y(new_n11186_));
  OR2X1    g11122(.A(new_n11186_), .B(new_n11184_), .Y(new_n11187_));
  AND2X1   g11123(.A(new_n11187_), .B(new_n10894_), .Y(new_n11188_));
  XOR2X1   g11124(.A(new_n10886_), .B(new_n10882_), .Y(new_n11189_));
  OAI21X1  g11125(.A0(new_n11189_), .A1(new_n11188_), .B0(new_n10888_), .Y(new_n11190_));
  XOR2X1   g11126(.A(new_n10880_), .B(new_n10876_), .Y(new_n11191_));
  AOI21X1  g11127(.A0(new_n11191_), .A1(new_n11190_), .B0(new_n10881_), .Y(new_n11192_));
  INVX1    g11128(.A(new_n11192_), .Y(new_n11193_));
  OAI21X1  g11129(.A0(new_n10875_), .A1(new_n10874_), .B0(new_n11193_), .Y(new_n11194_));
  NOR3X1   g11130(.A(new_n11193_), .B(new_n10875_), .C(new_n10874_), .Y(new_n11195_));
  AOI22X1  g11131(.A0(new_n7643_), .A1(new_n5960_), .B0(new_n7590_), .B1(new_n5373_), .Y(new_n11196_));
  OAI21X1  g11132(.A0(new_n7642_), .A1(new_n5658_), .B0(new_n11196_), .Y(new_n11197_));
  AOI21X1  g11133(.A0(new_n7718_), .A1(new_n67_), .B0(new_n11197_), .Y(new_n11198_));
  XOR2X1   g11134(.A(new_n11198_), .B(\a[5] ), .Y(new_n11199_));
  OAI21X1  g11135(.A0(new_n11199_), .A1(new_n11195_), .B0(new_n11194_), .Y(new_n11200_));
  OAI21X1  g11136(.A0(new_n10873_), .A1(new_n10871_), .B0(new_n11200_), .Y(new_n11201_));
  NOR3X1   g11137(.A(new_n11200_), .B(new_n10873_), .C(new_n10871_), .Y(new_n11202_));
  NAND3X1  g11138(.A(new_n10849_), .B(new_n10845_), .C(new_n10867_), .Y(new_n11203_));
  OAI21X1  g11139(.A0(new_n10868_), .A1(new_n10844_), .B0(new_n10850_), .Y(new_n11204_));
  NAND3X1  g11140(.A(new_n11192_), .B(new_n11204_), .C(new_n11203_), .Y(new_n11205_));
  NAND3X1  g11141(.A(new_n11199_), .B(new_n11205_), .C(new_n11194_), .Y(new_n11206_));
  AOI21X1  g11142(.A0(new_n11204_), .A1(new_n11203_), .B0(new_n11192_), .Y(new_n11207_));
  INVX1    g11143(.A(new_n11199_), .Y(new_n11208_));
  OAI21X1  g11144(.A0(new_n11195_), .A1(new_n11207_), .B0(new_n11208_), .Y(new_n11209_));
  AOI22X1  g11145(.A0(new_n7590_), .A1(new_n5659_), .B0(new_n7578_), .B1(new_n5373_), .Y(new_n11210_));
  OAI21X1  g11146(.A0(new_n7642_), .A1(new_n5959_), .B0(new_n11210_), .Y(new_n11211_));
  AOI21X1  g11147(.A0(new_n7712_), .A1(new_n67_), .B0(new_n11211_), .Y(new_n11212_));
  XOR2X1   g11148(.A(new_n11212_), .B(\a[5] ), .Y(new_n11213_));
  INVX1    g11149(.A(new_n11213_), .Y(new_n11214_));
  XOR2X1   g11150(.A(new_n11191_), .B(new_n11190_), .Y(new_n11215_));
  AND2X1   g11151(.A(new_n11215_), .B(new_n11214_), .Y(new_n11216_));
  INVX1    g11152(.A(new_n11216_), .Y(new_n11217_));
  XOR2X1   g11153(.A(new_n11215_), .B(new_n11213_), .Y(new_n11218_));
  OR2X1    g11154(.A(new_n6308_), .B(new_n6300_), .Y(new_n11219_));
  AOI22X1  g11155(.A0(new_n11219_), .A1(new_n7341_), .B0(new_n7643_), .B1(new_n5970_), .Y(new_n11220_));
  OAI21X1  g11156(.A0(new_n7808_), .A1(new_n6298_), .B0(new_n11220_), .Y(new_n11221_));
  XOR2X1   g11157(.A(new_n11221_), .B(new_n3431_), .Y(new_n11222_));
  OR2X1    g11158(.A(new_n11222_), .B(new_n11218_), .Y(new_n11223_));
  AND2X1   g11159(.A(new_n11223_), .B(new_n11217_), .Y(new_n11224_));
  AOI21X1  g11160(.A0(new_n11209_), .A1(new_n11206_), .B0(new_n11224_), .Y(new_n11225_));
  NAND3X1  g11161(.A(new_n11224_), .B(new_n11209_), .C(new_n11206_), .Y(new_n11226_));
  XOR2X1   g11162(.A(new_n11215_), .B(new_n11214_), .Y(new_n11227_));
  XOR2X1   g11163(.A(new_n11222_), .B(new_n11227_), .Y(new_n11228_));
  AOI22X1  g11164(.A0(new_n7578_), .A1(new_n5659_), .B0(new_n7571_), .B1(new_n5373_), .Y(new_n11229_));
  OAI21X1  g11165(.A0(new_n7594_), .A1(new_n5959_), .B0(new_n11229_), .Y(new_n11230_));
  AOI21X1  g11166(.A0(new_n7593_), .A1(new_n67_), .B0(new_n11230_), .Y(new_n11231_));
  XOR2X1   g11167(.A(new_n11231_), .B(\a[5] ), .Y(new_n11232_));
  OAI21X1  g11168(.A0(new_n11186_), .A1(new_n11184_), .B0(new_n10894_), .Y(new_n11233_));
  XOR2X1   g11169(.A(new_n11189_), .B(new_n11233_), .Y(new_n11234_));
  NOR2X1   g11170(.A(new_n11234_), .B(new_n11232_), .Y(new_n11235_));
  XOR2X1   g11171(.A(new_n11234_), .B(new_n11232_), .Y(new_n11236_));
  AOI22X1  g11172(.A0(new_n7571_), .A1(new_n5659_), .B0(new_n7558_), .B1(new_n5373_), .Y(new_n11237_));
  OAI21X1  g11173(.A0(new_n7602_), .A1(new_n5959_), .B0(new_n11237_), .Y(new_n11238_));
  AOI21X1  g11174(.A0(new_n7601_), .A1(new_n67_), .B0(new_n11238_), .Y(new_n11239_));
  XOR2X1   g11175(.A(new_n11239_), .B(\a[5] ), .Y(new_n11240_));
  XOR2X1   g11176(.A(new_n10893_), .B(new_n10889_), .Y(new_n11241_));
  XOR2X1   g11177(.A(new_n11241_), .B(new_n11184_), .Y(new_n11242_));
  NOR2X1   g11178(.A(new_n11242_), .B(new_n11240_), .Y(new_n11243_));
  XOR2X1   g11179(.A(new_n11242_), .B(new_n11240_), .Y(new_n11244_));
  AOI22X1  g11180(.A0(new_n7558_), .A1(new_n5659_), .B0(new_n7529_), .B1(new_n5373_), .Y(new_n11245_));
  OAI21X1  g11181(.A0(new_n7623_), .A1(new_n5959_), .B0(new_n11245_), .Y(new_n11246_));
  AOI21X1  g11182(.A0(new_n7622_), .A1(new_n67_), .B0(new_n11246_), .Y(new_n11247_));
  XOR2X1   g11183(.A(new_n11247_), .B(\a[5] ), .Y(new_n11248_));
  XOR2X1   g11184(.A(new_n10837_), .B(new_n10590_), .Y(new_n11249_));
  XOR2X1   g11185(.A(new_n10900_), .B(new_n11249_), .Y(new_n11250_));
  XOR2X1   g11186(.A(new_n11250_), .B(new_n11182_), .Y(new_n11251_));
  OR2X1    g11187(.A(new_n11251_), .B(new_n11248_), .Y(new_n11252_));
  INVX1    g11188(.A(new_n11248_), .Y(new_n11253_));
  XOR2X1   g11189(.A(new_n11251_), .B(new_n11253_), .Y(new_n11254_));
  AOI22X1  g11190(.A0(new_n7529_), .A1(new_n5659_), .B0(new_n7522_), .B1(new_n5373_), .Y(new_n11255_));
  OAI21X1  g11191(.A0(new_n7581_), .A1(new_n5959_), .B0(new_n11255_), .Y(new_n11256_));
  AOI21X1  g11192(.A0(new_n7565_), .A1(new_n67_), .B0(new_n11256_), .Y(new_n11257_));
  XOR2X1   g11193(.A(new_n11257_), .B(\a[5] ), .Y(new_n11258_));
  INVX1    g11194(.A(new_n11181_), .Y(new_n11259_));
  XOR2X1   g11195(.A(new_n11259_), .B(new_n11179_), .Y(new_n11260_));
  NOR2X1   g11196(.A(new_n11260_), .B(new_n11258_), .Y(new_n11261_));
  XOR2X1   g11197(.A(new_n11260_), .B(new_n11258_), .Y(new_n11262_));
  AOI22X1  g11198(.A0(new_n7522_), .A1(new_n5659_), .B0(new_n7485_), .B1(new_n5373_), .Y(new_n11263_));
  OAI21X1  g11199(.A0(new_n7537_), .A1(new_n5959_), .B0(new_n11263_), .Y(new_n11264_));
  AOI21X1  g11200(.A0(new_n7536_), .A1(new_n67_), .B0(new_n11264_), .Y(new_n11265_));
  XOR2X1   g11201(.A(new_n11265_), .B(\a[5] ), .Y(new_n11266_));
  INVX1    g11202(.A(new_n11178_), .Y(new_n11267_));
  XOR2X1   g11203(.A(new_n11267_), .B(new_n11177_), .Y(new_n11268_));
  OR2X1    g11204(.A(new_n11268_), .B(new_n11266_), .Y(new_n11269_));
  INVX1    g11205(.A(new_n11266_), .Y(new_n11270_));
  XOR2X1   g11206(.A(new_n11268_), .B(new_n11270_), .Y(new_n11271_));
  AOI22X1  g11207(.A0(new_n7485_), .A1(new_n5659_), .B0(new_n7364_), .B1(new_n5373_), .Y(new_n11272_));
  OAI21X1  g11208(.A0(new_n7523_), .A1(new_n5959_), .B0(new_n11272_), .Y(new_n11273_));
  AOI21X1  g11209(.A0(new_n7612_), .A1(new_n67_), .B0(new_n11273_), .Y(new_n11274_));
  XOR2X1   g11210(.A(new_n11274_), .B(\a[5] ), .Y(new_n11275_));
  XOR2X1   g11211(.A(new_n11176_), .B(new_n11173_), .Y(new_n11276_));
  NOR2X1   g11212(.A(new_n11276_), .B(new_n11275_), .Y(new_n11277_));
  XOR2X1   g11213(.A(new_n11276_), .B(new_n11275_), .Y(new_n11278_));
  AOI22X1  g11214(.A0(new_n7364_), .A1(new_n5659_), .B0(new_n7044_), .B1(new_n5373_), .Y(new_n11279_));
  OAI21X1  g11215(.A0(new_n7504_), .A1(new_n5959_), .B0(new_n11279_), .Y(new_n11280_));
  AOI21X1  g11216(.A0(new_n7552_), .A1(new_n67_), .B0(new_n11280_), .Y(new_n11281_));
  XOR2X1   g11217(.A(new_n11281_), .B(\a[5] ), .Y(new_n11282_));
  XOR2X1   g11218(.A(new_n11171_), .B(new_n11170_), .Y(new_n11283_));
  NOR2X1   g11219(.A(new_n11283_), .B(new_n11282_), .Y(new_n11284_));
  INVX1    g11220(.A(new_n11284_), .Y(new_n11285_));
  XOR2X1   g11221(.A(new_n11283_), .B(new_n11282_), .Y(new_n11286_));
  INVX1    g11222(.A(new_n11286_), .Y(new_n11287_));
  AOI22X1  g11223(.A0(new_n7044_), .A1(new_n5659_), .B0(new_n6818_), .B1(new_n5373_), .Y(new_n11288_));
  OAI21X1  g11224(.A0(new_n7367_), .A1(new_n5959_), .B0(new_n11288_), .Y(new_n11289_));
  AOI21X1  g11225(.A0(new_n7366_), .A1(new_n67_), .B0(new_n11289_), .Y(new_n11290_));
  XOR2X1   g11226(.A(new_n11290_), .B(\a[5] ), .Y(new_n11291_));
  XOR2X1   g11227(.A(new_n11168_), .B(new_n11166_), .Y(new_n11292_));
  NOR2X1   g11228(.A(new_n11292_), .B(new_n11291_), .Y(new_n11293_));
  XOR2X1   g11229(.A(new_n11292_), .B(new_n11291_), .Y(new_n11294_));
  AOI22X1  g11230(.A0(new_n6818_), .A1(new_n5659_), .B0(new_n6745_), .B1(new_n5373_), .Y(new_n11295_));
  OAI21X1  g11231(.A0(new_n7047_), .A1(new_n5959_), .B0(new_n11295_), .Y(new_n11296_));
  AOI21X1  g11232(.A0(new_n7046_), .A1(new_n67_), .B0(new_n11296_), .Y(new_n11297_));
  XOR2X1   g11233(.A(new_n11297_), .B(\a[5] ), .Y(new_n11298_));
  NOR2X1   g11234(.A(new_n11162_), .B(new_n10945_), .Y(new_n11299_));
  XOR2X1   g11235(.A(new_n11164_), .B(new_n11299_), .Y(new_n11300_));
  NOR2X1   g11236(.A(new_n11300_), .B(new_n11298_), .Y(new_n11301_));
  INVX1    g11237(.A(new_n11301_), .Y(new_n11302_));
  XOR2X1   g11238(.A(new_n11300_), .B(new_n11298_), .Y(new_n11303_));
  INVX1    g11239(.A(new_n11303_), .Y(new_n11304_));
  AND2X1   g11240(.A(new_n11161_), .B(new_n10955_), .Y(new_n11305_));
  XOR2X1   g11241(.A(new_n11305_), .B(new_n10947_), .Y(new_n11306_));
  OAI22X1  g11242(.A0(new_n7671_), .A1(new_n5372_), .B0(new_n7418_), .B1(new_n5658_), .Y(new_n11307_));
  AOI21X1  g11243(.A0(new_n6818_), .A1(new_n5960_), .B0(new_n11307_), .Y(new_n11308_));
  OAI21X1  g11244(.A0(new_n7403_), .A1(new_n5657_), .B0(new_n11308_), .Y(new_n11309_));
  XOR2X1   g11245(.A(new_n11309_), .B(\a[5] ), .Y(new_n11310_));
  AND2X1   g11246(.A(new_n11310_), .B(new_n11306_), .Y(new_n11311_));
  XOR2X1   g11247(.A(new_n11160_), .B(new_n10957_), .Y(new_n11312_));
  INVX1    g11248(.A(new_n11312_), .Y(new_n11313_));
  OAI22X1  g11249(.A0(new_n7472_), .A1(new_n5372_), .B0(new_n7671_), .B1(new_n5658_), .Y(new_n11314_));
  AOI21X1  g11250(.A0(new_n6745_), .A1(new_n5960_), .B0(new_n11314_), .Y(new_n11315_));
  OAI21X1  g11251(.A0(new_n7416_), .A1(new_n5657_), .B0(new_n11315_), .Y(new_n11316_));
  XOR2X1   g11252(.A(new_n11316_), .B(new_n3289_), .Y(new_n11317_));
  AOI22X1  g11253(.A0(new_n6882_), .A1(new_n5373_), .B0(new_n6822_), .B1(new_n5659_), .Y(new_n11318_));
  OAI21X1  g11254(.A0(new_n7671_), .A1(new_n5959_), .B0(new_n11318_), .Y(new_n11319_));
  AOI21X1  g11255(.A0(new_n7670_), .A1(new_n67_), .B0(new_n11319_), .Y(new_n11320_));
  XOR2X1   g11256(.A(new_n11320_), .B(\a[5] ), .Y(new_n11321_));
  XOR2X1   g11257(.A(new_n11159_), .B(new_n11157_), .Y(new_n11322_));
  NOR2X1   g11258(.A(new_n11322_), .B(new_n11321_), .Y(new_n11323_));
  INVX1    g11259(.A(new_n11321_), .Y(new_n11324_));
  XOR2X1   g11260(.A(new_n11322_), .B(new_n11324_), .Y(new_n11325_));
  AOI22X1  g11261(.A0(new_n6885_), .A1(new_n5373_), .B0(new_n6882_), .B1(new_n5659_), .Y(new_n11326_));
  OAI21X1  g11262(.A0(new_n7472_), .A1(new_n5959_), .B0(new_n11326_), .Y(new_n11327_));
  AOI21X1  g11263(.A0(new_n7471_), .A1(new_n67_), .B0(new_n11327_), .Y(new_n11328_));
  XOR2X1   g11264(.A(new_n11328_), .B(\a[5] ), .Y(new_n11329_));
  INVX1    g11265(.A(new_n11155_), .Y(new_n11330_));
  XOR2X1   g11266(.A(new_n11330_), .B(new_n11153_), .Y(new_n11331_));
  NOR2X1   g11267(.A(new_n11331_), .B(new_n11329_), .Y(new_n11332_));
  XOR2X1   g11268(.A(new_n11331_), .B(new_n11329_), .Y(new_n11333_));
  AOI22X1  g11269(.A0(new_n6887_), .A1(new_n5373_), .B0(new_n6885_), .B1(new_n5659_), .Y(new_n11334_));
  OAI21X1  g11270(.A0(new_n6884_), .A1(new_n5959_), .B0(new_n11334_), .Y(new_n11335_));
  AOI21X1  g11271(.A0(new_n7771_), .A1(new_n67_), .B0(new_n11335_), .Y(new_n11336_));
  XOR2X1   g11272(.A(new_n11336_), .B(\a[5] ), .Y(new_n11337_));
  XOR2X1   g11273(.A(new_n11151_), .B(new_n11149_), .Y(new_n11338_));
  NOR2X1   g11274(.A(new_n11338_), .B(new_n11337_), .Y(new_n11339_));
  INVX1    g11275(.A(new_n11339_), .Y(new_n11340_));
  XOR2X1   g11276(.A(new_n11338_), .B(new_n11337_), .Y(new_n11341_));
  INVX1    g11277(.A(new_n11341_), .Y(new_n11342_));
  XOR2X1   g11278(.A(new_n11148_), .B(new_n10984_), .Y(new_n11343_));
  INVX1    g11279(.A(new_n11343_), .Y(new_n11344_));
  OAI22X1  g11280(.A0(new_n7885_), .A1(new_n5372_), .B0(new_n7878_), .B1(new_n5658_), .Y(new_n11345_));
  AOI21X1  g11281(.A0(new_n6885_), .A1(new_n5960_), .B0(new_n11345_), .Y(new_n11346_));
  OAI21X1  g11282(.A0(new_n8083_), .A1(new_n5657_), .B0(new_n11346_), .Y(new_n11347_));
  XOR2X1   g11283(.A(new_n11347_), .B(new_n3289_), .Y(new_n11348_));
  NOR2X1   g11284(.A(new_n11348_), .B(new_n11344_), .Y(new_n11349_));
  XOR2X1   g11285(.A(new_n11146_), .B(new_n10993_), .Y(new_n11350_));
  OAI22X1  g11286(.A0(new_n8075_), .A1(new_n5372_), .B0(new_n7885_), .B1(new_n5658_), .Y(new_n11351_));
  AOI21X1  g11287(.A0(new_n6887_), .A1(new_n5960_), .B0(new_n11351_), .Y(new_n11352_));
  OAI21X1  g11288(.A0(new_n7876_), .A1(new_n5657_), .B0(new_n11352_), .Y(new_n11353_));
  XOR2X1   g11289(.A(new_n11353_), .B(\a[5] ), .Y(new_n11354_));
  AND2X1   g11290(.A(new_n11354_), .B(new_n11350_), .Y(new_n11355_));
  XOR2X1   g11291(.A(new_n11145_), .B(new_n11000_), .Y(new_n11356_));
  OAI22X1  g11292(.A0(new_n6896_), .A1(new_n5372_), .B0(new_n8075_), .B1(new_n5658_), .Y(new_n11357_));
  AOI21X1  g11293(.A0(new_n6890_), .A1(new_n5960_), .B0(new_n11357_), .Y(new_n11358_));
  OAI21X1  g11294(.A0(new_n9738_), .A1(new_n5657_), .B0(new_n11358_), .Y(new_n11359_));
  XOR2X1   g11295(.A(new_n11359_), .B(\a[5] ), .Y(new_n11360_));
  AND2X1   g11296(.A(new_n11360_), .B(new_n11356_), .Y(new_n11361_));
  INVX1    g11297(.A(new_n11361_), .Y(new_n11362_));
  AOI22X1  g11298(.A0(new_n6897_), .A1(new_n5373_), .B0(new_n6894_), .B1(new_n5659_), .Y(new_n11363_));
  OAI21X1  g11299(.A0(new_n8075_), .A1(new_n5959_), .B0(new_n11363_), .Y(new_n11364_));
  AOI21X1  g11300(.A0(new_n8074_), .A1(new_n67_), .B0(new_n11364_), .Y(new_n11365_));
  XOR2X1   g11301(.A(new_n11365_), .B(\a[5] ), .Y(new_n11366_));
  INVX1    g11302(.A(new_n11366_), .Y(new_n11367_));
  XOR2X1   g11303(.A(new_n11143_), .B(new_n11142_), .Y(new_n11368_));
  AND2X1   g11304(.A(new_n11368_), .B(new_n11367_), .Y(new_n11369_));
  INVX1    g11305(.A(new_n11369_), .Y(new_n11370_));
  XOR2X1   g11306(.A(new_n11368_), .B(new_n11366_), .Y(new_n11371_));
  AOI22X1  g11307(.A0(new_n6899_), .A1(new_n5373_), .B0(new_n6897_), .B1(new_n5659_), .Y(new_n11372_));
  OAI21X1  g11308(.A0(new_n6896_), .A1(new_n5959_), .B0(new_n11372_), .Y(new_n11373_));
  AOI21X1  g11309(.A0(new_n7953_), .A1(new_n67_), .B0(new_n11373_), .Y(new_n11374_));
  XOR2X1   g11310(.A(new_n11374_), .B(\a[5] ), .Y(new_n11375_));
  INVX1    g11311(.A(new_n11141_), .Y(new_n11376_));
  XOR2X1   g11312(.A(new_n11376_), .B(new_n11140_), .Y(new_n11377_));
  NOR2X1   g11313(.A(new_n11377_), .B(new_n11375_), .Y(new_n11378_));
  XOR2X1   g11314(.A(new_n11377_), .B(new_n11375_), .Y(new_n11379_));
  AOI22X1  g11315(.A0(new_n6902_), .A1(new_n5373_), .B0(new_n6899_), .B1(new_n5659_), .Y(new_n11380_));
  OAI21X1  g11316(.A0(new_n6898_), .A1(new_n5959_), .B0(new_n11380_), .Y(new_n11381_));
  AOI21X1  g11317(.A0(new_n8215_), .A1(new_n67_), .B0(new_n11381_), .Y(new_n11382_));
  XOR2X1   g11318(.A(new_n11382_), .B(\a[5] ), .Y(new_n11383_));
  XOR2X1   g11319(.A(new_n11138_), .B(new_n11137_), .Y(new_n11384_));
  XOR2X1   g11320(.A(new_n11384_), .B(new_n11383_), .Y(new_n11385_));
  INVX1    g11321(.A(new_n11385_), .Y(new_n11386_));
  XOR2X1   g11322(.A(new_n11136_), .B(new_n11029_), .Y(new_n11387_));
  INVX1    g11323(.A(new_n11387_), .Y(new_n11388_));
  OAI22X1  g11324(.A0(new_n8200_), .A1(new_n5372_), .B0(new_n8205_), .B1(new_n5658_), .Y(new_n11389_));
  AOI21X1  g11325(.A0(new_n6899_), .A1(new_n5960_), .B0(new_n11389_), .Y(new_n11390_));
  OAI21X1  g11326(.A0(new_n8293_), .A1(new_n5657_), .B0(new_n11390_), .Y(new_n11391_));
  XOR2X1   g11327(.A(new_n11391_), .B(new_n3289_), .Y(new_n11392_));
  NOR2X1   g11328(.A(new_n11392_), .B(new_n11388_), .Y(new_n11393_));
  XOR2X1   g11329(.A(new_n11135_), .B(new_n11036_), .Y(new_n11394_));
  OAI22X1  g11330(.A0(new_n6964_), .A1(new_n5372_), .B0(new_n8200_), .B1(new_n5658_), .Y(new_n11395_));
  AOI21X1  g11331(.A0(new_n6902_), .A1(new_n5960_), .B0(new_n11395_), .Y(new_n11396_));
  OAI21X1  g11332(.A0(new_n8203_), .A1(new_n5657_), .B0(new_n11396_), .Y(new_n11397_));
  XOR2X1   g11333(.A(new_n11397_), .B(\a[5] ), .Y(new_n11398_));
  AND2X1   g11334(.A(new_n11398_), .B(new_n11394_), .Y(new_n11399_));
  XOR2X1   g11335(.A(new_n11133_), .B(new_n11043_), .Y(new_n11400_));
  OAI22X1  g11336(.A0(new_n6960_), .A1(new_n5372_), .B0(new_n6964_), .B1(new_n5658_), .Y(new_n11401_));
  AOI21X1  g11337(.A0(new_n6904_), .A1(new_n5960_), .B0(new_n11401_), .Y(new_n11402_));
  OAI21X1  g11338(.A0(new_n8364_), .A1(new_n5657_), .B0(new_n11402_), .Y(new_n11403_));
  XOR2X1   g11339(.A(new_n11403_), .B(\a[5] ), .Y(new_n11404_));
  NAND2X1  g11340(.A(new_n11404_), .B(new_n11400_), .Y(new_n11405_));
  AOI22X1  g11341(.A0(new_n6911_), .A1(new_n5373_), .B0(new_n6909_), .B1(new_n5659_), .Y(new_n11406_));
  OAI21X1  g11342(.A0(new_n6964_), .A1(new_n5959_), .B0(new_n11406_), .Y(new_n11407_));
  AOI21X1  g11343(.A0(new_n8541_), .A1(new_n67_), .B0(new_n11407_), .Y(new_n11408_));
  XOR2X1   g11344(.A(new_n11408_), .B(\a[5] ), .Y(new_n11409_));
  INVX1    g11345(.A(new_n11409_), .Y(new_n11410_));
  XOR2X1   g11346(.A(new_n11132_), .B(new_n11131_), .Y(new_n11411_));
  NAND2X1  g11347(.A(new_n11411_), .B(new_n11410_), .Y(new_n11412_));
  XOR2X1   g11348(.A(new_n11411_), .B(new_n11409_), .Y(new_n11413_));
  AOI22X1  g11349(.A0(new_n6913_), .A1(new_n5373_), .B0(new_n6911_), .B1(new_n5659_), .Y(new_n11414_));
  OAI21X1  g11350(.A0(new_n6960_), .A1(new_n5959_), .B0(new_n11414_), .Y(new_n11415_));
  AOI21X1  g11351(.A0(new_n8553_), .A1(new_n67_), .B0(new_n11415_), .Y(new_n11416_));
  XOR2X1   g11352(.A(new_n11416_), .B(\a[5] ), .Y(new_n11417_));
  XOR2X1   g11353(.A(new_n11130_), .B(new_n11128_), .Y(new_n11418_));
  NOR2X1   g11354(.A(new_n11418_), .B(new_n11417_), .Y(new_n11419_));
  XOR2X1   g11355(.A(new_n11418_), .B(new_n11417_), .Y(new_n11420_));
  AOI22X1  g11356(.A0(new_n6915_), .A1(new_n5373_), .B0(new_n6913_), .B1(new_n5659_), .Y(new_n11421_));
  OAI21X1  g11357(.A0(new_n8349_), .A1(new_n5959_), .B0(new_n11421_), .Y(new_n11422_));
  AOI21X1  g11358(.A0(new_n8348_), .A1(new_n67_), .B0(new_n11422_), .Y(new_n11423_));
  XOR2X1   g11359(.A(new_n11423_), .B(\a[5] ), .Y(new_n11424_));
  XOR2X1   g11360(.A(new_n11127_), .B(new_n11125_), .Y(new_n11425_));
  NOR2X1   g11361(.A(new_n11425_), .B(new_n11424_), .Y(new_n11426_));
  INVX1    g11362(.A(new_n11426_), .Y(new_n11427_));
  XOR2X1   g11363(.A(new_n11425_), .B(new_n11424_), .Y(new_n11428_));
  INVX1    g11364(.A(new_n11428_), .Y(new_n11429_));
  XOR2X1   g11365(.A(new_n11124_), .B(new_n11074_), .Y(new_n11430_));
  INVX1    g11366(.A(new_n11430_), .Y(new_n11431_));
  OAI22X1  g11367(.A0(new_n6918_), .A1(new_n5372_), .B0(new_n6917_), .B1(new_n5658_), .Y(new_n11432_));
  AOI21X1  g11368(.A0(new_n6913_), .A1(new_n5960_), .B0(new_n11432_), .Y(new_n11433_));
  OAI21X1  g11369(.A0(new_n8577_), .A1(new_n5657_), .B0(new_n11433_), .Y(new_n11434_));
  XOR2X1   g11370(.A(new_n11434_), .B(new_n3289_), .Y(new_n11435_));
  NOR2X1   g11371(.A(new_n11435_), .B(new_n11431_), .Y(new_n11436_));
  XOR2X1   g11372(.A(new_n11123_), .B(new_n11122_), .Y(new_n11437_));
  OAI22X1  g11373(.A0(new_n6920_), .A1(new_n5372_), .B0(new_n6918_), .B1(new_n5658_), .Y(new_n11438_));
  AOI21X1  g11374(.A0(new_n6915_), .A1(new_n5960_), .B0(new_n11438_), .Y(new_n11439_));
  OAI21X1  g11375(.A0(new_n9093_), .A1(new_n5657_), .B0(new_n11439_), .Y(new_n11440_));
  XOR2X1   g11376(.A(new_n11440_), .B(\a[5] ), .Y(new_n11441_));
  NAND2X1  g11377(.A(new_n11441_), .B(new_n11437_), .Y(new_n11442_));
  INVX1    g11378(.A(new_n11092_), .Y(new_n11443_));
  XOR2X1   g11379(.A(new_n11119_), .B(new_n11443_), .Y(new_n11444_));
  OAI22X1  g11380(.A0(new_n8659_), .A1(new_n5372_), .B0(new_n6920_), .B1(new_n5658_), .Y(new_n11445_));
  AOI21X1  g11381(.A0(new_n8580_), .A1(new_n5960_), .B0(new_n11445_), .Y(new_n11446_));
  OAI21X1  g11382(.A0(new_n8611_), .A1(new_n5657_), .B0(new_n11446_), .Y(new_n11447_));
  XOR2X1   g11383(.A(new_n11447_), .B(new_n3289_), .Y(new_n11448_));
  OR2X1    g11384(.A(new_n11448_), .B(new_n11444_), .Y(new_n11449_));
  AOI22X1  g11385(.A0(new_n6925_), .A1(new_n5373_), .B0(new_n6923_), .B1(new_n5659_), .Y(new_n11450_));
  OAI21X1  g11386(.A0(new_n6920_), .A1(new_n5959_), .B0(new_n11450_), .Y(new_n11451_));
  AOI21X1  g11387(.A0(new_n8628_), .A1(new_n67_), .B0(new_n11451_), .Y(new_n11452_));
  XOR2X1   g11388(.A(new_n11452_), .B(\a[5] ), .Y(new_n11453_));
  INVX1    g11389(.A(new_n11453_), .Y(new_n11454_));
  XOR2X1   g11390(.A(new_n11118_), .B(new_n11117_), .Y(new_n11455_));
  NAND2X1  g11391(.A(new_n11455_), .B(new_n11454_), .Y(new_n11456_));
  XOR2X1   g11392(.A(new_n11455_), .B(new_n11453_), .Y(new_n11457_));
  XOR2X1   g11393(.A(new_n11116_), .B(new_n11112_), .Y(new_n11458_));
  INVX1    g11394(.A(new_n11458_), .Y(new_n11459_));
  OAI22X1  g11395(.A0(new_n6929_), .A1(new_n5372_), .B0(new_n8683_), .B1(new_n5658_), .Y(new_n11460_));
  AOI21X1  g11396(.A0(new_n6923_), .A1(new_n5960_), .B0(new_n11460_), .Y(new_n11461_));
  OAI21X1  g11397(.A0(new_n8662_), .A1(new_n5657_), .B0(new_n11461_), .Y(new_n11462_));
  XOR2X1   g11398(.A(new_n11462_), .B(new_n3289_), .Y(new_n11463_));
  NOR2X1   g11399(.A(new_n11463_), .B(new_n11459_), .Y(new_n11464_));
  AOI22X1  g11400(.A0(new_n6932_), .A1(new_n5373_), .B0(new_n6927_), .B1(new_n5659_), .Y(new_n11465_));
  OAI21X1  g11401(.A0(new_n8683_), .A1(new_n5959_), .B0(new_n11465_), .Y(new_n11466_));
  AOI21X1  g11402(.A0(new_n8682_), .A1(new_n67_), .B0(new_n11466_), .Y(new_n11467_));
  XOR2X1   g11403(.A(new_n11467_), .B(\a[5] ), .Y(new_n11468_));
  INVX1    g11404(.A(new_n11468_), .Y(new_n11469_));
  XOR2X1   g11405(.A(new_n11108_), .B(new_n11104_), .Y(new_n11470_));
  NAND2X1  g11406(.A(new_n11470_), .B(new_n11469_), .Y(new_n11471_));
  XOR2X1   g11407(.A(new_n11470_), .B(new_n11468_), .Y(new_n11472_));
  NOR2X1   g11408(.A(new_n11102_), .B(new_n2995_), .Y(new_n11473_));
  XOR2X1   g11409(.A(new_n11473_), .B(new_n11110_), .Y(new_n11474_));
  OAI22X1  g11410(.A0(new_n8757_), .A1(new_n5372_), .B0(new_n6930_), .B1(new_n5658_), .Y(new_n11475_));
  AOI21X1  g11411(.A0(new_n6927_), .A1(new_n5960_), .B0(new_n11475_), .Y(new_n11476_));
  OAI21X1  g11412(.A0(new_n8705_), .A1(new_n5657_), .B0(new_n11476_), .Y(new_n11477_));
  XOR2X1   g11413(.A(new_n11477_), .B(new_n3289_), .Y(new_n11478_));
  NOR2X1   g11414(.A(new_n11478_), .B(new_n11474_), .Y(new_n11479_));
  OAI22X1  g11415(.A0(new_n6936_), .A1(new_n5658_), .B0(new_n8752_), .B1(new_n5959_), .Y(new_n11480_));
  AOI21X1  g11416(.A0(new_n8751_), .A1(new_n67_), .B0(new_n11480_), .Y(new_n11481_));
  XOR2X1   g11417(.A(new_n11481_), .B(\a[5] ), .Y(new_n11482_));
  NOR2X1   g11418(.A(new_n6936_), .B(new_n5369_), .Y(new_n11483_));
  OAI22X1  g11419(.A0(new_n6936_), .A1(new_n5372_), .B0(new_n8752_), .B1(new_n5658_), .Y(new_n11484_));
  AOI21X1  g11420(.A0(new_n6933_), .A1(new_n5960_), .B0(new_n11484_), .Y(new_n11485_));
  OAI21X1  g11421(.A0(new_n8759_), .A1(new_n5657_), .B0(new_n11485_), .Y(new_n11486_));
  NOR4X1   g11422(.A(new_n11486_), .B(new_n11483_), .C(new_n11482_), .D(new_n3289_), .Y(new_n11487_));
  NAND2X1  g11423(.A(new_n11487_), .B(new_n11102_), .Y(new_n11488_));
  XOR2X1   g11424(.A(new_n11487_), .B(new_n11103_), .Y(new_n11489_));
  AOI22X1  g11425(.A0(new_n6935_), .A1(new_n5373_), .B0(new_n6933_), .B1(new_n5659_), .Y(new_n11490_));
  OAI21X1  g11426(.A0(new_n6930_), .A1(new_n5959_), .B0(new_n11490_), .Y(new_n11491_));
  AOI21X1  g11427(.A0(new_n8717_), .A1(new_n67_), .B0(new_n11491_), .Y(new_n11492_));
  XOR2X1   g11428(.A(new_n11492_), .B(\a[5] ), .Y(new_n11493_));
  OAI21X1  g11429(.A0(new_n11493_), .A1(new_n11489_), .B0(new_n11488_), .Y(new_n11494_));
  XOR2X1   g11430(.A(new_n11478_), .B(new_n11474_), .Y(new_n11495_));
  AOI21X1  g11431(.A0(new_n11495_), .A1(new_n11494_), .B0(new_n11479_), .Y(new_n11496_));
  OAI21X1  g11432(.A0(new_n11496_), .A1(new_n11472_), .B0(new_n11471_), .Y(new_n11497_));
  XOR2X1   g11433(.A(new_n11463_), .B(new_n11459_), .Y(new_n11498_));
  AOI21X1  g11434(.A0(new_n11498_), .A1(new_n11497_), .B0(new_n11464_), .Y(new_n11499_));
  OAI21X1  g11435(.A0(new_n11499_), .A1(new_n11457_), .B0(new_n11456_), .Y(new_n11500_));
  XOR2X1   g11436(.A(new_n11448_), .B(new_n11444_), .Y(new_n11501_));
  NAND2X1  g11437(.A(new_n11501_), .B(new_n11500_), .Y(new_n11502_));
  AND2X1   g11438(.A(new_n11502_), .B(new_n11449_), .Y(new_n11503_));
  XOR2X1   g11439(.A(new_n11440_), .B(new_n3289_), .Y(new_n11504_));
  XOR2X1   g11440(.A(new_n11504_), .B(new_n11437_), .Y(new_n11505_));
  OAI21X1  g11441(.A0(new_n11505_), .A1(new_n11503_), .B0(new_n11442_), .Y(new_n11506_));
  XOR2X1   g11442(.A(new_n11435_), .B(new_n11430_), .Y(new_n11507_));
  INVX1    g11443(.A(new_n11507_), .Y(new_n11508_));
  AOI21X1  g11444(.A0(new_n11508_), .A1(new_n11506_), .B0(new_n11436_), .Y(new_n11509_));
  OAI21X1  g11445(.A0(new_n11509_), .A1(new_n11429_), .B0(new_n11427_), .Y(new_n11510_));
  AOI21X1  g11446(.A0(new_n11510_), .A1(new_n11420_), .B0(new_n11419_), .Y(new_n11511_));
  OAI21X1  g11447(.A0(new_n11511_), .A1(new_n11413_), .B0(new_n11412_), .Y(new_n11512_));
  INVX1    g11448(.A(new_n11512_), .Y(new_n11513_));
  XOR2X1   g11449(.A(new_n11403_), .B(new_n3289_), .Y(new_n11514_));
  XOR2X1   g11450(.A(new_n11514_), .B(new_n11400_), .Y(new_n11515_));
  OAI21X1  g11451(.A0(new_n11515_), .A1(new_n11513_), .B0(new_n11405_), .Y(new_n11516_));
  XOR2X1   g11452(.A(new_n11397_), .B(new_n3289_), .Y(new_n11517_));
  XOR2X1   g11453(.A(new_n11517_), .B(new_n11394_), .Y(new_n11518_));
  INVX1    g11454(.A(new_n11518_), .Y(new_n11519_));
  AND2X1   g11455(.A(new_n11519_), .B(new_n11516_), .Y(new_n11520_));
  OR2X1    g11456(.A(new_n11520_), .B(new_n11399_), .Y(new_n11521_));
  XOR2X1   g11457(.A(new_n11392_), .B(new_n11388_), .Y(new_n11522_));
  AOI21X1  g11458(.A0(new_n11522_), .A1(new_n11521_), .B0(new_n11393_), .Y(new_n11523_));
  OR2X1    g11459(.A(new_n11523_), .B(new_n11386_), .Y(new_n11524_));
  OAI21X1  g11460(.A0(new_n11384_), .A1(new_n11383_), .B0(new_n11524_), .Y(new_n11525_));
  AOI21X1  g11461(.A0(new_n11525_), .A1(new_n11379_), .B0(new_n11378_), .Y(new_n11526_));
  OAI21X1  g11462(.A0(new_n11526_), .A1(new_n11371_), .B0(new_n11370_), .Y(new_n11527_));
  INVX1    g11463(.A(new_n11527_), .Y(new_n11528_));
  XOR2X1   g11464(.A(new_n11359_), .B(new_n3289_), .Y(new_n11529_));
  XOR2X1   g11465(.A(new_n11529_), .B(new_n11356_), .Y(new_n11530_));
  OAI21X1  g11466(.A0(new_n11530_), .A1(new_n11528_), .B0(new_n11362_), .Y(new_n11531_));
  XOR2X1   g11467(.A(new_n11353_), .B(new_n3289_), .Y(new_n11532_));
  XOR2X1   g11468(.A(new_n11532_), .B(new_n11350_), .Y(new_n11533_));
  INVX1    g11469(.A(new_n11533_), .Y(new_n11534_));
  AOI21X1  g11470(.A0(new_n11534_), .A1(new_n11531_), .B0(new_n11355_), .Y(new_n11535_));
  INVX1    g11471(.A(new_n11535_), .Y(new_n11536_));
  XOR2X1   g11472(.A(new_n11348_), .B(new_n11344_), .Y(new_n11537_));
  AOI21X1  g11473(.A0(new_n11537_), .A1(new_n11536_), .B0(new_n11349_), .Y(new_n11538_));
  OAI21X1  g11474(.A0(new_n11538_), .A1(new_n11342_), .B0(new_n11340_), .Y(new_n11539_));
  AOI21X1  g11475(.A0(new_n11539_), .A1(new_n11333_), .B0(new_n11332_), .Y(new_n11540_));
  NOR2X1   g11476(.A(new_n11540_), .B(new_n11325_), .Y(new_n11541_));
  NOR2X1   g11477(.A(new_n11541_), .B(new_n11323_), .Y(new_n11542_));
  XOR2X1   g11478(.A(new_n11317_), .B(new_n11312_), .Y(new_n11543_));
  OR2X1    g11479(.A(new_n11543_), .B(new_n11542_), .Y(new_n11544_));
  OAI21X1  g11480(.A0(new_n11317_), .A1(new_n11313_), .B0(new_n11544_), .Y(new_n11545_));
  XOR2X1   g11481(.A(new_n11309_), .B(new_n3289_), .Y(new_n11546_));
  XOR2X1   g11482(.A(new_n11546_), .B(new_n11306_), .Y(new_n11547_));
  INVX1    g11483(.A(new_n11547_), .Y(new_n11548_));
  AOI21X1  g11484(.A0(new_n11548_), .A1(new_n11545_), .B0(new_n11311_), .Y(new_n11549_));
  OAI21X1  g11485(.A0(new_n11549_), .A1(new_n11304_), .B0(new_n11302_), .Y(new_n11550_));
  AOI21X1  g11486(.A0(new_n11550_), .A1(new_n11294_), .B0(new_n11293_), .Y(new_n11551_));
  OAI21X1  g11487(.A0(new_n11551_), .A1(new_n11287_), .B0(new_n11285_), .Y(new_n11552_));
  AOI21X1  g11488(.A0(new_n11552_), .A1(new_n11278_), .B0(new_n11277_), .Y(new_n11553_));
  OAI21X1  g11489(.A0(new_n11553_), .A1(new_n11271_), .B0(new_n11269_), .Y(new_n11554_));
  AOI21X1  g11490(.A0(new_n11554_), .A1(new_n11262_), .B0(new_n11261_), .Y(new_n11555_));
  OAI21X1  g11491(.A0(new_n11555_), .A1(new_n11254_), .B0(new_n11252_), .Y(new_n11556_));
  AOI21X1  g11492(.A0(new_n11556_), .A1(new_n11244_), .B0(new_n11243_), .Y(new_n11557_));
  INVX1    g11493(.A(new_n11557_), .Y(new_n11558_));
  AOI21X1  g11494(.A0(new_n11558_), .A1(new_n11236_), .B0(new_n11235_), .Y(new_n11559_));
  NOR2X1   g11495(.A(new_n11559_), .B(new_n11228_), .Y(new_n11560_));
  XOR2X1   g11496(.A(new_n11222_), .B(new_n11218_), .Y(new_n11561_));
  XOR2X1   g11497(.A(new_n11559_), .B(new_n11561_), .Y(new_n11562_));
  XOR2X1   g11498(.A(new_n11557_), .B(new_n11236_), .Y(new_n11563_));
  OAI22X1  g11499(.A0(new_n7642_), .A1(new_n6325_), .B0(new_n8172_), .B1(new_n6309_), .Y(new_n11564_));
  AOI21X1  g11500(.A0(new_n7643_), .A1(new_n6300_), .B0(new_n11564_), .Y(new_n11565_));
  OAI21X1  g11501(.A0(new_n7655_), .A1(new_n6298_), .B0(new_n11565_), .Y(new_n11566_));
  XOR2X1   g11502(.A(new_n11566_), .B(new_n3431_), .Y(new_n11567_));
  OR2X1    g11503(.A(new_n11567_), .B(new_n11563_), .Y(new_n11568_));
  XOR2X1   g11504(.A(new_n11556_), .B(new_n11244_), .Y(new_n11569_));
  AOI22X1  g11505(.A0(new_n7643_), .A1(new_n6308_), .B0(new_n7590_), .B1(new_n5970_), .Y(new_n11570_));
  OAI21X1  g11506(.A0(new_n7642_), .A1(new_n6307_), .B0(new_n11570_), .Y(new_n11571_));
  AOI21X1  g11507(.A0(new_n7718_), .A1(new_n5972_), .B0(new_n11571_), .Y(new_n11572_));
  XOR2X1   g11508(.A(new_n11572_), .B(new_n3431_), .Y(new_n11573_));
  AND2X1   g11509(.A(new_n11573_), .B(new_n11569_), .Y(new_n11574_));
  XOR2X1   g11510(.A(new_n11251_), .B(new_n11248_), .Y(new_n11575_));
  XOR2X1   g11511(.A(new_n11555_), .B(new_n11575_), .Y(new_n11576_));
  OAI22X1  g11512(.A0(new_n7594_), .A1(new_n6307_), .B0(new_n7602_), .B1(new_n6325_), .Y(new_n11577_));
  AOI21X1  g11513(.A0(new_n7657_), .A1(new_n6308_), .B0(new_n11577_), .Y(new_n11578_));
  OAI21X1  g11514(.A0(new_n7711_), .A1(new_n6298_), .B0(new_n11578_), .Y(new_n11579_));
  XOR2X1   g11515(.A(new_n11579_), .B(new_n3431_), .Y(new_n11580_));
  OR2X1    g11516(.A(new_n11580_), .B(new_n11576_), .Y(new_n11581_));
  XOR2X1   g11517(.A(new_n11554_), .B(new_n11262_), .Y(new_n11582_));
  INVX1    g11518(.A(new_n7593_), .Y(new_n11583_));
  OAI22X1  g11519(.A0(new_n7602_), .A1(new_n6307_), .B0(new_n7623_), .B1(new_n6325_), .Y(new_n11584_));
  AOI21X1  g11520(.A0(new_n7590_), .A1(new_n6308_), .B0(new_n11584_), .Y(new_n11585_));
  OAI21X1  g11521(.A0(new_n11583_), .A1(new_n6298_), .B0(new_n11585_), .Y(new_n11586_));
  XOR2X1   g11522(.A(new_n11586_), .B(\a[2] ), .Y(new_n11587_));
  AND2X1   g11523(.A(new_n11587_), .B(new_n11582_), .Y(new_n11588_));
  XOR2X1   g11524(.A(new_n11268_), .B(new_n11266_), .Y(new_n11589_));
  XOR2X1   g11525(.A(new_n11553_), .B(new_n11589_), .Y(new_n11590_));
  AOI22X1  g11526(.A0(new_n7571_), .A1(new_n6300_), .B0(new_n7558_), .B1(new_n5970_), .Y(new_n11591_));
  OAI21X1  g11527(.A0(new_n7602_), .A1(new_n6309_), .B0(new_n11591_), .Y(new_n11592_));
  AOI21X1  g11528(.A0(new_n7601_), .A1(new_n5972_), .B0(new_n11592_), .Y(new_n11593_));
  XOR2X1   g11529(.A(new_n11593_), .B(\a[2] ), .Y(new_n11594_));
  OR2X1    g11530(.A(new_n11594_), .B(new_n11590_), .Y(new_n11595_));
  XOR2X1   g11531(.A(new_n11552_), .B(new_n11278_), .Y(new_n11596_));
  OAI22X1  g11532(.A0(new_n7581_), .A1(new_n6307_), .B0(new_n7537_), .B1(new_n6325_), .Y(new_n11597_));
  AOI21X1  g11533(.A0(new_n7571_), .A1(new_n6308_), .B0(new_n11597_), .Y(new_n11598_));
  OAI21X1  g11534(.A0(new_n7621_), .A1(new_n6298_), .B0(new_n11598_), .Y(new_n11599_));
  XOR2X1   g11535(.A(new_n11599_), .B(\a[2] ), .Y(new_n11600_));
  AND2X1   g11536(.A(new_n11600_), .B(new_n11596_), .Y(new_n11601_));
  XOR2X1   g11537(.A(new_n11551_), .B(new_n11286_), .Y(new_n11602_));
  OAI22X1  g11538(.A0(new_n7537_), .A1(new_n6307_), .B0(new_n7523_), .B1(new_n6325_), .Y(new_n11603_));
  AOI21X1  g11539(.A0(new_n7558_), .A1(new_n6308_), .B0(new_n11603_), .Y(new_n11604_));
  OAI21X1  g11540(.A0(new_n7566_), .A1(new_n6298_), .B0(new_n11604_), .Y(new_n11605_));
  XOR2X1   g11541(.A(new_n11605_), .B(new_n3431_), .Y(new_n11606_));
  NOR2X1   g11542(.A(new_n11606_), .B(new_n11602_), .Y(new_n11607_));
  INVX1    g11543(.A(new_n11607_), .Y(new_n11608_));
  XOR2X1   g11544(.A(new_n11550_), .B(new_n11294_), .Y(new_n11609_));
  OAI22X1  g11545(.A0(new_n7523_), .A1(new_n6307_), .B0(new_n7504_), .B1(new_n6325_), .Y(new_n11610_));
  AOI21X1  g11546(.A0(new_n7529_), .A1(new_n6308_), .B0(new_n11610_), .Y(new_n11611_));
  OAI21X1  g11547(.A0(new_n7535_), .A1(new_n6298_), .B0(new_n11611_), .Y(new_n11612_));
  XOR2X1   g11548(.A(new_n11612_), .B(\a[2] ), .Y(new_n11613_));
  AND2X1   g11549(.A(new_n11613_), .B(new_n11609_), .Y(new_n11614_));
  XOR2X1   g11550(.A(new_n11549_), .B(new_n11303_), .Y(new_n11615_));
  OAI22X1  g11551(.A0(new_n7504_), .A1(new_n6307_), .B0(new_n7367_), .B1(new_n6325_), .Y(new_n11616_));
  AOI21X1  g11552(.A0(new_n7522_), .A1(new_n6308_), .B0(new_n11616_), .Y(new_n11617_));
  OAI21X1  g11553(.A0(new_n7611_), .A1(new_n6298_), .B0(new_n11617_), .Y(new_n11618_));
  XOR2X1   g11554(.A(new_n11618_), .B(new_n3431_), .Y(new_n11619_));
  NOR2X1   g11555(.A(new_n11619_), .B(new_n11615_), .Y(new_n11620_));
  INVX1    g11556(.A(new_n11620_), .Y(new_n11621_));
  XOR2X1   g11557(.A(new_n11548_), .B(new_n11545_), .Y(new_n11622_));
  XOR2X1   g11558(.A(new_n11537_), .B(new_n11535_), .Y(new_n11623_));
  INVX1    g11559(.A(new_n11623_), .Y(new_n11624_));
  AOI21X1  g11560(.A0(new_n11519_), .A1(new_n11516_), .B0(new_n11399_), .Y(new_n11625_));
  XOR2X1   g11561(.A(new_n11522_), .B(new_n11625_), .Y(new_n11626_));
  XOR2X1   g11562(.A(new_n11507_), .B(new_n11506_), .Y(new_n11627_));
  INVX1    g11563(.A(new_n11627_), .Y(new_n11628_));
  XOR2X1   g11564(.A(new_n11495_), .B(new_n11494_), .Y(new_n11629_));
  INVX1    g11565(.A(new_n11629_), .Y(new_n11630_));
  OAI21X1  g11566(.A0(new_n6936_), .A1(new_n5369_), .B0(\a[5] ), .Y(new_n11631_));
  NOR2X1   g11567(.A(new_n11631_), .B(new_n11482_), .Y(new_n11632_));
  XOR2X1   g11568(.A(new_n11486_), .B(new_n3289_), .Y(new_n11633_));
  XOR2X1   g11569(.A(new_n11633_), .B(new_n11632_), .Y(new_n11634_));
  INVX1    g11570(.A(new_n11634_), .Y(new_n11635_));
  AOI22X1  g11571(.A0(new_n6937_), .A1(new_n5970_), .B0(new_n6935_), .B1(new_n6300_), .Y(new_n11636_));
  OAI21X1  g11572(.A0(new_n8757_), .A1(new_n6309_), .B0(new_n11636_), .Y(new_n11637_));
  AND2X1   g11573(.A(new_n11637_), .B(\a[2] ), .Y(new_n11638_));
  NOR2X1   g11574(.A(new_n8759_), .B(new_n6351_), .Y(new_n11639_));
  AND2X1   g11575(.A(new_n8751_), .B(new_n6350_), .Y(new_n11640_));
  OAI21X1  g11576(.A0(new_n6936_), .A1(new_n6357_), .B0(\a[2] ), .Y(new_n11641_));
  AOI21X1  g11577(.A0(new_n6937_), .A1(new_n6360_), .B0(new_n11641_), .Y(new_n11642_));
  OAI21X1  g11578(.A0(new_n8752_), .A1(new_n6362_), .B0(new_n11642_), .Y(new_n11643_));
  NOR4X1   g11579(.A(new_n11643_), .B(new_n11640_), .C(new_n11639_), .D(new_n11638_), .Y(new_n11644_));
  AND2X1   g11580(.A(new_n11644_), .B(new_n11483_), .Y(new_n11645_));
  OR2X1    g11581(.A(new_n11644_), .B(new_n11483_), .Y(new_n11646_));
  AOI22X1  g11582(.A0(new_n6935_), .A1(new_n5970_), .B0(new_n6933_), .B1(new_n6300_), .Y(new_n11647_));
  OAI21X1  g11583(.A0(new_n6930_), .A1(new_n6309_), .B0(new_n11647_), .Y(new_n11648_));
  AOI21X1  g11584(.A0(new_n8717_), .A1(new_n5972_), .B0(new_n11648_), .Y(new_n11649_));
  XOR2X1   g11585(.A(new_n11649_), .B(new_n3431_), .Y(new_n11650_));
  AOI21X1  g11586(.A0(new_n11650_), .A1(new_n11646_), .B0(new_n11645_), .Y(new_n11651_));
  OAI22X1  g11587(.A0(new_n8757_), .A1(new_n6325_), .B0(new_n6930_), .B1(new_n6307_), .Y(new_n11652_));
  AOI21X1  g11588(.A0(new_n6927_), .A1(new_n6308_), .B0(new_n11652_), .Y(new_n11653_));
  OAI21X1  g11589(.A0(new_n8705_), .A1(new_n6298_), .B0(new_n11653_), .Y(new_n11654_));
  XOR2X1   g11590(.A(new_n11654_), .B(new_n3431_), .Y(new_n11655_));
  XOR2X1   g11591(.A(new_n11631_), .B(new_n11482_), .Y(new_n11656_));
  INVX1    g11592(.A(new_n11656_), .Y(new_n11657_));
  AOI21X1  g11593(.A0(new_n11655_), .A1(new_n11651_), .B0(new_n11657_), .Y(new_n11658_));
  NAND2X1  g11594(.A(new_n11644_), .B(new_n11483_), .Y(new_n11659_));
  NOR2X1   g11595(.A(new_n11644_), .B(new_n11483_), .Y(new_n11660_));
  XOR2X1   g11596(.A(new_n11649_), .B(\a[2] ), .Y(new_n11661_));
  OAI21X1  g11597(.A0(new_n11661_), .A1(new_n11660_), .B0(new_n11659_), .Y(new_n11662_));
  XOR2X1   g11598(.A(new_n11654_), .B(\a[2] ), .Y(new_n11663_));
  AND2X1   g11599(.A(new_n11663_), .B(new_n11662_), .Y(new_n11664_));
  OAI21X1  g11600(.A0(new_n11664_), .A1(new_n11658_), .B0(new_n11635_), .Y(new_n11665_));
  NOR3X1   g11601(.A(new_n11664_), .B(new_n11658_), .C(new_n11635_), .Y(new_n11666_));
  AOI22X1  g11602(.A0(new_n6932_), .A1(new_n5970_), .B0(new_n6927_), .B1(new_n6300_), .Y(new_n11667_));
  OAI21X1  g11603(.A0(new_n8683_), .A1(new_n6309_), .B0(new_n11667_), .Y(new_n11668_));
  AOI21X1  g11604(.A0(new_n8682_), .A1(new_n5972_), .B0(new_n11668_), .Y(new_n11669_));
  XOR2X1   g11605(.A(new_n11669_), .B(\a[2] ), .Y(new_n11670_));
  OAI21X1  g11606(.A0(new_n11670_), .A1(new_n11666_), .B0(new_n11665_), .Y(new_n11671_));
  OAI22X1  g11607(.A0(new_n6929_), .A1(new_n6325_), .B0(new_n8683_), .B1(new_n6307_), .Y(new_n11672_));
  AOI21X1  g11608(.A0(new_n6923_), .A1(new_n6308_), .B0(new_n11672_), .Y(new_n11673_));
  OAI21X1  g11609(.A0(new_n8662_), .A1(new_n6298_), .B0(new_n11673_), .Y(new_n11674_));
  XOR2X1   g11610(.A(new_n11674_), .B(\a[2] ), .Y(new_n11675_));
  NAND2X1  g11611(.A(new_n11675_), .B(new_n11671_), .Y(new_n11676_));
  XOR2X1   g11612(.A(new_n11493_), .B(new_n11489_), .Y(new_n11677_));
  OAI21X1  g11613(.A0(new_n11675_), .A1(new_n11671_), .B0(new_n11677_), .Y(new_n11678_));
  AOI21X1  g11614(.A0(new_n11678_), .A1(new_n11676_), .B0(new_n11630_), .Y(new_n11679_));
  NAND3X1  g11615(.A(new_n11678_), .B(new_n11676_), .C(new_n11630_), .Y(new_n11680_));
  AOI22X1  g11616(.A0(new_n6925_), .A1(new_n5970_), .B0(new_n6923_), .B1(new_n6300_), .Y(new_n11681_));
  OAI21X1  g11617(.A0(new_n6920_), .A1(new_n6309_), .B0(new_n11681_), .Y(new_n11682_));
  AOI21X1  g11618(.A0(new_n8628_), .A1(new_n5972_), .B0(new_n11682_), .Y(new_n11683_));
  XOR2X1   g11619(.A(new_n11683_), .B(\a[2] ), .Y(new_n11684_));
  INVX1    g11620(.A(new_n11684_), .Y(new_n11685_));
  AOI21X1  g11621(.A0(new_n11685_), .A1(new_n11680_), .B0(new_n11679_), .Y(new_n11686_));
  OAI22X1  g11622(.A0(new_n8659_), .A1(new_n6325_), .B0(new_n6920_), .B1(new_n6307_), .Y(new_n11687_));
  AOI21X1  g11623(.A0(new_n8580_), .A1(new_n6308_), .B0(new_n11687_), .Y(new_n11688_));
  OAI21X1  g11624(.A0(new_n8611_), .A1(new_n6298_), .B0(new_n11688_), .Y(new_n11689_));
  XOR2X1   g11625(.A(new_n11689_), .B(new_n3431_), .Y(new_n11690_));
  XOR2X1   g11626(.A(new_n11496_), .B(new_n11472_), .Y(new_n11691_));
  INVX1    g11627(.A(new_n11691_), .Y(new_n11692_));
  AOI21X1  g11628(.A0(new_n11690_), .A1(new_n11686_), .B0(new_n11692_), .Y(new_n11693_));
  NOR2X1   g11629(.A(new_n11690_), .B(new_n11686_), .Y(new_n11694_));
  OAI22X1  g11630(.A0(new_n6920_), .A1(new_n6325_), .B0(new_n6918_), .B1(new_n6307_), .Y(new_n11695_));
  AOI21X1  g11631(.A0(new_n6915_), .A1(new_n6308_), .B0(new_n11695_), .Y(new_n11696_));
  OAI21X1  g11632(.A0(new_n9093_), .A1(new_n6298_), .B0(new_n11696_), .Y(new_n11697_));
  XOR2X1   g11633(.A(new_n11697_), .B(\a[2] ), .Y(new_n11698_));
  NOR3X1   g11634(.A(new_n11698_), .B(new_n11694_), .C(new_n11693_), .Y(new_n11699_));
  XOR2X1   g11635(.A(new_n11498_), .B(new_n11497_), .Y(new_n11700_));
  INVX1    g11636(.A(new_n11700_), .Y(new_n11701_));
  OAI21X1  g11637(.A0(new_n11694_), .A1(new_n11693_), .B0(new_n11698_), .Y(new_n11702_));
  OAI21X1  g11638(.A0(new_n11701_), .A1(new_n11699_), .B0(new_n11702_), .Y(new_n11703_));
  OAI22X1  g11639(.A0(new_n6918_), .A1(new_n6325_), .B0(new_n6917_), .B1(new_n6307_), .Y(new_n11704_));
  AOI21X1  g11640(.A0(new_n6913_), .A1(new_n6308_), .B0(new_n11704_), .Y(new_n11705_));
  OAI21X1  g11641(.A0(new_n8577_), .A1(new_n6298_), .B0(new_n11705_), .Y(new_n11706_));
  XOR2X1   g11642(.A(new_n11706_), .B(new_n3431_), .Y(new_n11707_));
  INVX1    g11643(.A(new_n11707_), .Y(new_n11708_));
  XOR2X1   g11644(.A(new_n11499_), .B(new_n11457_), .Y(new_n11709_));
  OAI21X1  g11645(.A0(new_n11708_), .A1(new_n11703_), .B0(new_n11709_), .Y(new_n11710_));
  NAND2X1  g11646(.A(new_n11708_), .B(new_n11703_), .Y(new_n11711_));
  XOR2X1   g11647(.A(new_n11501_), .B(new_n11500_), .Y(new_n11712_));
  INVX1    g11648(.A(new_n11712_), .Y(new_n11713_));
  AOI21X1  g11649(.A0(new_n11711_), .A1(new_n11710_), .B0(new_n11713_), .Y(new_n11714_));
  NAND3X1  g11650(.A(new_n11713_), .B(new_n11711_), .C(new_n11710_), .Y(new_n11715_));
  AOI22X1  g11651(.A0(new_n6915_), .A1(new_n5970_), .B0(new_n6913_), .B1(new_n6300_), .Y(new_n11716_));
  OAI21X1  g11652(.A0(new_n8349_), .A1(new_n6309_), .B0(new_n11716_), .Y(new_n11717_));
  AOI21X1  g11653(.A0(new_n8348_), .A1(new_n5972_), .B0(new_n11717_), .Y(new_n11718_));
  XOR2X1   g11654(.A(new_n11718_), .B(\a[2] ), .Y(new_n11719_));
  INVX1    g11655(.A(new_n11719_), .Y(new_n11720_));
  AOI21X1  g11656(.A0(new_n11720_), .A1(new_n11715_), .B0(new_n11714_), .Y(new_n11721_));
  XOR2X1   g11657(.A(new_n11505_), .B(new_n11503_), .Y(new_n11722_));
  INVX1    g11658(.A(new_n11722_), .Y(new_n11723_));
  NOR2X1   g11659(.A(new_n11723_), .B(new_n11721_), .Y(new_n11724_));
  AOI22X1  g11660(.A0(new_n6913_), .A1(new_n5970_), .B0(new_n6911_), .B1(new_n6300_), .Y(new_n11725_));
  OAI21X1  g11661(.A0(new_n6960_), .A1(new_n6309_), .B0(new_n11725_), .Y(new_n11726_));
  AOI21X1  g11662(.A0(new_n8553_), .A1(new_n5972_), .B0(new_n11726_), .Y(new_n11727_));
  XOR2X1   g11663(.A(new_n11727_), .B(\a[2] ), .Y(new_n11728_));
  AOI21X1  g11664(.A0(new_n11723_), .A1(new_n11721_), .B0(new_n11728_), .Y(new_n11729_));
  OAI21X1  g11665(.A0(new_n11729_), .A1(new_n11724_), .B0(new_n11628_), .Y(new_n11730_));
  NOR3X1   g11666(.A(new_n11729_), .B(new_n11724_), .C(new_n11628_), .Y(new_n11731_));
  AOI22X1  g11667(.A0(new_n6911_), .A1(new_n5970_), .B0(new_n6909_), .B1(new_n6300_), .Y(new_n11732_));
  OAI21X1  g11668(.A0(new_n6964_), .A1(new_n6309_), .B0(new_n11732_), .Y(new_n11733_));
  AOI21X1  g11669(.A0(new_n8541_), .A1(new_n5972_), .B0(new_n11733_), .Y(new_n11734_));
  XOR2X1   g11670(.A(new_n11734_), .B(\a[2] ), .Y(new_n11735_));
  OAI21X1  g11671(.A0(new_n11735_), .A1(new_n11731_), .B0(new_n11730_), .Y(new_n11736_));
  OAI22X1  g11672(.A0(new_n6960_), .A1(new_n6325_), .B0(new_n6964_), .B1(new_n6307_), .Y(new_n11737_));
  AOI21X1  g11673(.A0(new_n6904_), .A1(new_n6308_), .B0(new_n11737_), .Y(new_n11738_));
  OAI21X1  g11674(.A0(new_n8364_), .A1(new_n6298_), .B0(new_n11738_), .Y(new_n11739_));
  XOR2X1   g11675(.A(new_n11739_), .B(\a[2] ), .Y(new_n11740_));
  XOR2X1   g11676(.A(new_n11509_), .B(new_n11429_), .Y(new_n11741_));
  OAI21X1  g11677(.A0(new_n11740_), .A1(new_n11736_), .B0(new_n11741_), .Y(new_n11742_));
  NAND2X1  g11678(.A(new_n11740_), .B(new_n11736_), .Y(new_n11743_));
  OAI22X1  g11679(.A0(new_n6964_), .A1(new_n6325_), .B0(new_n8200_), .B1(new_n6307_), .Y(new_n11744_));
  AOI21X1  g11680(.A0(new_n6902_), .A1(new_n6308_), .B0(new_n11744_), .Y(new_n11745_));
  OAI21X1  g11681(.A0(new_n8203_), .A1(new_n6298_), .B0(new_n11745_), .Y(new_n11746_));
  XOR2X1   g11682(.A(new_n11746_), .B(new_n3431_), .Y(new_n11747_));
  NAND3X1  g11683(.A(new_n11747_), .B(new_n11743_), .C(new_n11742_), .Y(new_n11748_));
  XOR2X1   g11684(.A(new_n11510_), .B(new_n11420_), .Y(new_n11749_));
  AOI21X1  g11685(.A0(new_n11743_), .A1(new_n11742_), .B0(new_n11747_), .Y(new_n11750_));
  AOI21X1  g11686(.A0(new_n11749_), .A1(new_n11748_), .B0(new_n11750_), .Y(new_n11751_));
  OAI22X1  g11687(.A0(new_n8200_), .A1(new_n6325_), .B0(new_n8205_), .B1(new_n6307_), .Y(new_n11752_));
  AOI21X1  g11688(.A0(new_n6899_), .A1(new_n6308_), .B0(new_n11752_), .Y(new_n11753_));
  OAI21X1  g11689(.A0(new_n8293_), .A1(new_n6298_), .B0(new_n11753_), .Y(new_n11754_));
  XOR2X1   g11690(.A(new_n11754_), .B(new_n3431_), .Y(new_n11755_));
  XOR2X1   g11691(.A(new_n11511_), .B(new_n11413_), .Y(new_n11756_));
  INVX1    g11692(.A(new_n11756_), .Y(new_n11757_));
  AOI21X1  g11693(.A0(new_n11755_), .A1(new_n11751_), .B0(new_n11757_), .Y(new_n11758_));
  NOR2X1   g11694(.A(new_n11755_), .B(new_n11751_), .Y(new_n11759_));
  XOR2X1   g11695(.A(new_n11515_), .B(new_n11512_), .Y(new_n11760_));
  INVX1    g11696(.A(new_n11760_), .Y(new_n11761_));
  OAI21X1  g11697(.A0(new_n11759_), .A1(new_n11758_), .B0(new_n11761_), .Y(new_n11762_));
  NOR3X1   g11698(.A(new_n11761_), .B(new_n11759_), .C(new_n11758_), .Y(new_n11763_));
  AOI22X1  g11699(.A0(new_n6902_), .A1(new_n5970_), .B0(new_n6899_), .B1(new_n6300_), .Y(new_n11764_));
  OAI21X1  g11700(.A0(new_n6898_), .A1(new_n6309_), .B0(new_n11764_), .Y(new_n11765_));
  AOI21X1  g11701(.A0(new_n8215_), .A1(new_n5972_), .B0(new_n11765_), .Y(new_n11766_));
  XOR2X1   g11702(.A(new_n11766_), .B(\a[2] ), .Y(new_n11767_));
  OAI21X1  g11703(.A0(new_n11767_), .A1(new_n11763_), .B0(new_n11762_), .Y(new_n11768_));
  XOR2X1   g11704(.A(new_n11518_), .B(new_n11516_), .Y(new_n11769_));
  INVX1    g11705(.A(new_n11769_), .Y(new_n11770_));
  NAND2X1  g11706(.A(new_n11770_), .B(new_n11768_), .Y(new_n11771_));
  AOI22X1  g11707(.A0(new_n6899_), .A1(new_n5970_), .B0(new_n6897_), .B1(new_n6300_), .Y(new_n11772_));
  OAI21X1  g11708(.A0(new_n6896_), .A1(new_n6309_), .B0(new_n11772_), .Y(new_n11773_));
  AOI21X1  g11709(.A0(new_n7953_), .A1(new_n5972_), .B0(new_n11773_), .Y(new_n11774_));
  XOR2X1   g11710(.A(new_n11774_), .B(\a[2] ), .Y(new_n11775_));
  INVX1    g11711(.A(new_n11775_), .Y(new_n11776_));
  OAI21X1  g11712(.A0(new_n11770_), .A1(new_n11768_), .B0(new_n11776_), .Y(new_n11777_));
  AOI21X1  g11713(.A0(new_n11777_), .A1(new_n11771_), .B0(new_n11626_), .Y(new_n11778_));
  NAND3X1  g11714(.A(new_n11777_), .B(new_n11771_), .C(new_n11626_), .Y(new_n11779_));
  AOI22X1  g11715(.A0(new_n6897_), .A1(new_n5970_), .B0(new_n6894_), .B1(new_n6300_), .Y(new_n11780_));
  OAI21X1  g11716(.A0(new_n8075_), .A1(new_n6309_), .B0(new_n11780_), .Y(new_n11781_));
  AOI21X1  g11717(.A0(new_n8074_), .A1(new_n5972_), .B0(new_n11781_), .Y(new_n11782_));
  XOR2X1   g11718(.A(new_n11782_), .B(\a[2] ), .Y(new_n11783_));
  INVX1    g11719(.A(new_n11783_), .Y(new_n11784_));
  AOI21X1  g11720(.A0(new_n11784_), .A1(new_n11779_), .B0(new_n11778_), .Y(new_n11785_));
  OAI22X1  g11721(.A0(new_n6896_), .A1(new_n6325_), .B0(new_n8075_), .B1(new_n6307_), .Y(new_n11786_));
  AOI21X1  g11722(.A0(new_n6890_), .A1(new_n6308_), .B0(new_n11786_), .Y(new_n11787_));
  OAI21X1  g11723(.A0(new_n9738_), .A1(new_n6298_), .B0(new_n11787_), .Y(new_n11788_));
  XOR2X1   g11724(.A(new_n11788_), .B(new_n3431_), .Y(new_n11789_));
  XOR2X1   g11725(.A(new_n11523_), .B(new_n11385_), .Y(new_n11790_));
  AOI21X1  g11726(.A0(new_n11789_), .A1(new_n11785_), .B0(new_n11790_), .Y(new_n11791_));
  NOR2X1   g11727(.A(new_n11789_), .B(new_n11785_), .Y(new_n11792_));
  OAI22X1  g11728(.A0(new_n8075_), .A1(new_n6325_), .B0(new_n7885_), .B1(new_n6307_), .Y(new_n11793_));
  AOI21X1  g11729(.A0(new_n6887_), .A1(new_n6308_), .B0(new_n11793_), .Y(new_n11794_));
  OAI21X1  g11730(.A0(new_n7876_), .A1(new_n6298_), .B0(new_n11794_), .Y(new_n11795_));
  XOR2X1   g11731(.A(new_n11795_), .B(new_n3431_), .Y(new_n11796_));
  INVX1    g11732(.A(new_n11796_), .Y(new_n11797_));
  NOR3X1   g11733(.A(new_n11797_), .B(new_n11792_), .C(new_n11791_), .Y(new_n11798_));
  XOR2X1   g11734(.A(new_n11525_), .B(new_n11379_), .Y(new_n11799_));
  INVX1    g11735(.A(new_n11799_), .Y(new_n11800_));
  OAI21X1  g11736(.A0(new_n11792_), .A1(new_n11791_), .B0(new_n11797_), .Y(new_n11801_));
  OAI21X1  g11737(.A0(new_n11800_), .A1(new_n11798_), .B0(new_n11801_), .Y(new_n11802_));
  OAI22X1  g11738(.A0(new_n7885_), .A1(new_n6325_), .B0(new_n7878_), .B1(new_n6307_), .Y(new_n11803_));
  AOI21X1  g11739(.A0(new_n6885_), .A1(new_n6308_), .B0(new_n11803_), .Y(new_n11804_));
  OAI21X1  g11740(.A0(new_n8083_), .A1(new_n6298_), .B0(new_n11804_), .Y(new_n11805_));
  XOR2X1   g11741(.A(new_n11805_), .B(new_n3431_), .Y(new_n11806_));
  INVX1    g11742(.A(new_n11806_), .Y(new_n11807_));
  XOR2X1   g11743(.A(new_n11526_), .B(new_n11371_), .Y(new_n11808_));
  OAI21X1  g11744(.A0(new_n11807_), .A1(new_n11802_), .B0(new_n11808_), .Y(new_n11809_));
  NAND2X1  g11745(.A(new_n11807_), .B(new_n11802_), .Y(new_n11810_));
  XOR2X1   g11746(.A(new_n11530_), .B(new_n11527_), .Y(new_n11811_));
  AOI21X1  g11747(.A0(new_n11810_), .A1(new_n11809_), .B0(new_n11811_), .Y(new_n11812_));
  NAND3X1  g11748(.A(new_n11811_), .B(new_n11810_), .C(new_n11809_), .Y(new_n11813_));
  AOI22X1  g11749(.A0(new_n6887_), .A1(new_n5970_), .B0(new_n6885_), .B1(new_n6300_), .Y(new_n11814_));
  OAI21X1  g11750(.A0(new_n6884_), .A1(new_n6309_), .B0(new_n11814_), .Y(new_n11815_));
  AOI21X1  g11751(.A0(new_n7771_), .A1(new_n5972_), .B0(new_n11815_), .Y(new_n11816_));
  XOR2X1   g11752(.A(new_n11816_), .B(\a[2] ), .Y(new_n11817_));
  INVX1    g11753(.A(new_n11817_), .Y(new_n11818_));
  AOI21X1  g11754(.A0(new_n11818_), .A1(new_n11813_), .B0(new_n11812_), .Y(new_n11819_));
  XOR2X1   g11755(.A(new_n11534_), .B(new_n11531_), .Y(new_n11820_));
  INVX1    g11756(.A(new_n11820_), .Y(new_n11821_));
  NOR2X1   g11757(.A(new_n11821_), .B(new_n11819_), .Y(new_n11822_));
  AOI22X1  g11758(.A0(new_n6885_), .A1(new_n5970_), .B0(new_n6882_), .B1(new_n6300_), .Y(new_n11823_));
  OAI21X1  g11759(.A0(new_n7472_), .A1(new_n6309_), .B0(new_n11823_), .Y(new_n11824_));
  AOI21X1  g11760(.A0(new_n7471_), .A1(new_n5972_), .B0(new_n11824_), .Y(new_n11825_));
  XOR2X1   g11761(.A(new_n11825_), .B(\a[2] ), .Y(new_n11826_));
  AOI21X1  g11762(.A0(new_n11821_), .A1(new_n11819_), .B0(new_n11826_), .Y(new_n11827_));
  OAI21X1  g11763(.A0(new_n11827_), .A1(new_n11822_), .B0(new_n11624_), .Y(new_n11828_));
  NOR3X1   g11764(.A(new_n11827_), .B(new_n11822_), .C(new_n11624_), .Y(new_n11829_));
  AOI22X1  g11765(.A0(new_n6882_), .A1(new_n5970_), .B0(new_n6822_), .B1(new_n6300_), .Y(new_n11830_));
  OAI21X1  g11766(.A0(new_n7671_), .A1(new_n6309_), .B0(new_n11830_), .Y(new_n11831_));
  AOI21X1  g11767(.A0(new_n7670_), .A1(new_n5972_), .B0(new_n11831_), .Y(new_n11832_));
  XOR2X1   g11768(.A(new_n11832_), .B(\a[2] ), .Y(new_n11833_));
  OAI21X1  g11769(.A0(new_n11833_), .A1(new_n11829_), .B0(new_n11828_), .Y(new_n11834_));
  OAI22X1  g11770(.A0(new_n7472_), .A1(new_n6325_), .B0(new_n7671_), .B1(new_n6307_), .Y(new_n11835_));
  AOI21X1  g11771(.A0(new_n6745_), .A1(new_n6308_), .B0(new_n11835_), .Y(new_n11836_));
  OAI21X1  g11772(.A0(new_n7416_), .A1(new_n6298_), .B0(new_n11836_), .Y(new_n11837_));
  XOR2X1   g11773(.A(new_n11837_), .B(new_n3431_), .Y(new_n11838_));
  INVX1    g11774(.A(new_n11838_), .Y(new_n11839_));
  XOR2X1   g11775(.A(new_n11538_), .B(new_n11342_), .Y(new_n11840_));
  OAI21X1  g11776(.A0(new_n11839_), .A1(new_n11834_), .B0(new_n11840_), .Y(new_n11841_));
  NAND2X1  g11777(.A(new_n11839_), .B(new_n11834_), .Y(new_n11842_));
  OAI22X1  g11778(.A0(new_n7671_), .A1(new_n6325_), .B0(new_n7418_), .B1(new_n6307_), .Y(new_n11843_));
  AOI21X1  g11779(.A0(new_n6818_), .A1(new_n6308_), .B0(new_n11843_), .Y(new_n11844_));
  OAI21X1  g11780(.A0(new_n7403_), .A1(new_n6298_), .B0(new_n11844_), .Y(new_n11845_));
  XOR2X1   g11781(.A(new_n11845_), .B(new_n3431_), .Y(new_n11846_));
  NAND3X1  g11782(.A(new_n11846_), .B(new_n11842_), .C(new_n11841_), .Y(new_n11847_));
  XOR2X1   g11783(.A(new_n11539_), .B(new_n11333_), .Y(new_n11848_));
  AOI21X1  g11784(.A0(new_n11842_), .A1(new_n11841_), .B0(new_n11846_), .Y(new_n11849_));
  AOI21X1  g11785(.A0(new_n11848_), .A1(new_n11847_), .B0(new_n11849_), .Y(new_n11850_));
  OAI22X1  g11786(.A0(new_n7361_), .A1(new_n6307_), .B0(new_n7418_), .B1(new_n6325_), .Y(new_n11851_));
  AOI21X1  g11787(.A0(new_n7044_), .A1(new_n6308_), .B0(new_n11851_), .Y(new_n11852_));
  OAI21X1  g11788(.A0(new_n7680_), .A1(new_n6298_), .B0(new_n11852_), .Y(new_n11853_));
  XOR2X1   g11789(.A(new_n11853_), .B(new_n3431_), .Y(new_n11854_));
  XOR2X1   g11790(.A(new_n11540_), .B(new_n11325_), .Y(new_n11855_));
  INVX1    g11791(.A(new_n11855_), .Y(new_n11856_));
  AOI21X1  g11792(.A0(new_n11854_), .A1(new_n11850_), .B0(new_n11856_), .Y(new_n11857_));
  NOR2X1   g11793(.A(new_n11854_), .B(new_n11850_), .Y(new_n11858_));
  XOR2X1   g11794(.A(new_n11543_), .B(new_n11542_), .Y(new_n11859_));
  OAI21X1  g11795(.A0(new_n11858_), .A1(new_n11857_), .B0(new_n11859_), .Y(new_n11860_));
  NOR3X1   g11796(.A(new_n11859_), .B(new_n11858_), .C(new_n11857_), .Y(new_n11861_));
  AOI22X1  g11797(.A0(new_n7044_), .A1(new_n6300_), .B0(new_n6818_), .B1(new_n5970_), .Y(new_n11862_));
  OAI21X1  g11798(.A0(new_n7367_), .A1(new_n6309_), .B0(new_n11862_), .Y(new_n11863_));
  AOI21X1  g11799(.A0(new_n7366_), .A1(new_n5972_), .B0(new_n11863_), .Y(new_n11864_));
  XOR2X1   g11800(.A(new_n11864_), .B(\a[2] ), .Y(new_n11865_));
  OAI21X1  g11801(.A0(new_n11865_), .A1(new_n11861_), .B0(new_n11860_), .Y(new_n11866_));
  AND2X1   g11802(.A(new_n11866_), .B(new_n11622_), .Y(new_n11867_));
  INVX1    g11803(.A(new_n11622_), .Y(new_n11868_));
  OR2X1    g11804(.A(new_n11821_), .B(new_n11819_), .Y(new_n11869_));
  XOR2X1   g11805(.A(new_n11522_), .B(new_n11521_), .Y(new_n11870_));
  AND2X1   g11806(.A(new_n11770_), .B(new_n11768_), .Y(new_n11871_));
  OR2X1    g11807(.A(new_n11723_), .B(new_n11721_), .Y(new_n11872_));
  AND2X1   g11808(.A(new_n11675_), .B(new_n11671_), .Y(new_n11873_));
  OAI21X1  g11809(.A0(new_n11663_), .A1(new_n11662_), .B0(new_n11656_), .Y(new_n11874_));
  OR2X1    g11810(.A(new_n11655_), .B(new_n11651_), .Y(new_n11875_));
  AOI21X1  g11811(.A0(new_n11875_), .A1(new_n11874_), .B0(new_n11634_), .Y(new_n11876_));
  NAND3X1  g11812(.A(new_n11875_), .B(new_n11874_), .C(new_n11634_), .Y(new_n11877_));
  XOR2X1   g11813(.A(new_n11669_), .B(new_n3431_), .Y(new_n11878_));
  AOI21X1  g11814(.A0(new_n11878_), .A1(new_n11877_), .B0(new_n11876_), .Y(new_n11879_));
  XOR2X1   g11815(.A(new_n11674_), .B(new_n3431_), .Y(new_n11880_));
  INVX1    g11816(.A(new_n11677_), .Y(new_n11881_));
  AOI21X1  g11817(.A0(new_n11880_), .A1(new_n11879_), .B0(new_n11881_), .Y(new_n11882_));
  OAI21X1  g11818(.A0(new_n11882_), .A1(new_n11873_), .B0(new_n11629_), .Y(new_n11883_));
  NOR3X1   g11819(.A(new_n11882_), .B(new_n11873_), .C(new_n11629_), .Y(new_n11884_));
  OAI21X1  g11820(.A0(new_n11684_), .A1(new_n11884_), .B0(new_n11883_), .Y(new_n11885_));
  XOR2X1   g11821(.A(new_n11689_), .B(\a[2] ), .Y(new_n11886_));
  OAI21X1  g11822(.A0(new_n11886_), .A1(new_n11885_), .B0(new_n11691_), .Y(new_n11887_));
  OR2X1    g11823(.A(new_n11690_), .B(new_n11686_), .Y(new_n11888_));
  XOR2X1   g11824(.A(new_n11697_), .B(new_n3431_), .Y(new_n11889_));
  NAND3X1  g11825(.A(new_n11889_), .B(new_n11888_), .C(new_n11887_), .Y(new_n11890_));
  AOI21X1  g11826(.A0(new_n11888_), .A1(new_n11887_), .B0(new_n11889_), .Y(new_n11891_));
  AOI21X1  g11827(.A0(new_n11700_), .A1(new_n11890_), .B0(new_n11891_), .Y(new_n11892_));
  INVX1    g11828(.A(new_n11709_), .Y(new_n11893_));
  AOI21X1  g11829(.A0(new_n11707_), .A1(new_n11892_), .B0(new_n11893_), .Y(new_n11894_));
  AND2X1   g11830(.A(new_n11708_), .B(new_n11703_), .Y(new_n11895_));
  OAI21X1  g11831(.A0(new_n11895_), .A1(new_n11894_), .B0(new_n11712_), .Y(new_n11896_));
  NOR3X1   g11832(.A(new_n11712_), .B(new_n11895_), .C(new_n11894_), .Y(new_n11897_));
  OAI21X1  g11833(.A0(new_n11719_), .A1(new_n11897_), .B0(new_n11896_), .Y(new_n11898_));
  INVX1    g11834(.A(new_n11728_), .Y(new_n11899_));
  OAI21X1  g11835(.A0(new_n11722_), .A1(new_n11898_), .B0(new_n11899_), .Y(new_n11900_));
  AOI21X1  g11836(.A0(new_n11900_), .A1(new_n11872_), .B0(new_n11627_), .Y(new_n11901_));
  NAND3X1  g11837(.A(new_n11900_), .B(new_n11872_), .C(new_n11627_), .Y(new_n11902_));
  XOR2X1   g11838(.A(new_n11734_), .B(new_n3431_), .Y(new_n11903_));
  AOI21X1  g11839(.A0(new_n11903_), .A1(new_n11902_), .B0(new_n11901_), .Y(new_n11904_));
  XOR2X1   g11840(.A(new_n11739_), .B(new_n3431_), .Y(new_n11905_));
  INVX1    g11841(.A(new_n11741_), .Y(new_n11906_));
  AOI21X1  g11842(.A0(new_n11905_), .A1(new_n11904_), .B0(new_n11906_), .Y(new_n11907_));
  AND2X1   g11843(.A(new_n11740_), .B(new_n11736_), .Y(new_n11908_));
  INVX1    g11844(.A(new_n11747_), .Y(new_n11909_));
  NOR3X1   g11845(.A(new_n11909_), .B(new_n11908_), .C(new_n11907_), .Y(new_n11910_));
  INVX1    g11846(.A(new_n11749_), .Y(new_n11911_));
  OAI21X1  g11847(.A0(new_n11908_), .A1(new_n11907_), .B0(new_n11909_), .Y(new_n11912_));
  OAI21X1  g11848(.A0(new_n11911_), .A1(new_n11910_), .B0(new_n11912_), .Y(new_n11913_));
  INVX1    g11849(.A(new_n11755_), .Y(new_n11914_));
  OAI21X1  g11850(.A0(new_n11914_), .A1(new_n11913_), .B0(new_n11756_), .Y(new_n11915_));
  OR2X1    g11851(.A(new_n11755_), .B(new_n11751_), .Y(new_n11916_));
  AOI21X1  g11852(.A0(new_n11916_), .A1(new_n11915_), .B0(new_n11760_), .Y(new_n11917_));
  NAND3X1  g11853(.A(new_n11760_), .B(new_n11916_), .C(new_n11915_), .Y(new_n11918_));
  INVX1    g11854(.A(new_n11767_), .Y(new_n11919_));
  AOI21X1  g11855(.A0(new_n11919_), .A1(new_n11918_), .B0(new_n11917_), .Y(new_n11920_));
  AOI21X1  g11856(.A0(new_n11769_), .A1(new_n11920_), .B0(new_n11775_), .Y(new_n11921_));
  OAI21X1  g11857(.A0(new_n11921_), .A1(new_n11871_), .B0(new_n11870_), .Y(new_n11922_));
  NOR3X1   g11858(.A(new_n11921_), .B(new_n11871_), .C(new_n11870_), .Y(new_n11923_));
  OAI21X1  g11859(.A0(new_n11783_), .A1(new_n11923_), .B0(new_n11922_), .Y(new_n11924_));
  INVX1    g11860(.A(new_n11789_), .Y(new_n11925_));
  XOR2X1   g11861(.A(new_n11523_), .B(new_n11386_), .Y(new_n11926_));
  OAI21X1  g11862(.A0(new_n11925_), .A1(new_n11924_), .B0(new_n11926_), .Y(new_n11927_));
  OR2X1    g11863(.A(new_n11789_), .B(new_n11785_), .Y(new_n11928_));
  NAND3X1  g11864(.A(new_n11796_), .B(new_n11928_), .C(new_n11927_), .Y(new_n11929_));
  AOI21X1  g11865(.A0(new_n11928_), .A1(new_n11927_), .B0(new_n11796_), .Y(new_n11930_));
  AOI21X1  g11866(.A0(new_n11799_), .A1(new_n11929_), .B0(new_n11930_), .Y(new_n11931_));
  INVX1    g11867(.A(new_n11808_), .Y(new_n11932_));
  AOI21X1  g11868(.A0(new_n11806_), .A1(new_n11931_), .B0(new_n11932_), .Y(new_n11933_));
  AND2X1   g11869(.A(new_n11807_), .B(new_n11802_), .Y(new_n11934_));
  INVX1    g11870(.A(new_n11811_), .Y(new_n11935_));
  OAI21X1  g11871(.A0(new_n11934_), .A1(new_n11933_), .B0(new_n11935_), .Y(new_n11936_));
  NOR3X1   g11872(.A(new_n11935_), .B(new_n11934_), .C(new_n11933_), .Y(new_n11937_));
  OAI21X1  g11873(.A0(new_n11817_), .A1(new_n11937_), .B0(new_n11936_), .Y(new_n11938_));
  INVX1    g11874(.A(new_n11826_), .Y(new_n11939_));
  OAI21X1  g11875(.A0(new_n11820_), .A1(new_n11938_), .B0(new_n11939_), .Y(new_n11940_));
  AOI21X1  g11876(.A0(new_n11940_), .A1(new_n11869_), .B0(new_n11623_), .Y(new_n11941_));
  NAND3X1  g11877(.A(new_n11940_), .B(new_n11869_), .C(new_n11623_), .Y(new_n11942_));
  INVX1    g11878(.A(new_n11833_), .Y(new_n11943_));
  AOI21X1  g11879(.A0(new_n11943_), .A1(new_n11942_), .B0(new_n11941_), .Y(new_n11944_));
  INVX1    g11880(.A(new_n11840_), .Y(new_n11945_));
  AOI21X1  g11881(.A0(new_n11838_), .A1(new_n11944_), .B0(new_n11945_), .Y(new_n11946_));
  AND2X1   g11882(.A(new_n11839_), .B(new_n11834_), .Y(new_n11947_));
  INVX1    g11883(.A(new_n11846_), .Y(new_n11948_));
  NOR3X1   g11884(.A(new_n11948_), .B(new_n11947_), .C(new_n11946_), .Y(new_n11949_));
  INVX1    g11885(.A(new_n11848_), .Y(new_n11950_));
  OAI21X1  g11886(.A0(new_n11947_), .A1(new_n11946_), .B0(new_n11948_), .Y(new_n11951_));
  OAI21X1  g11887(.A0(new_n11950_), .A1(new_n11949_), .B0(new_n11951_), .Y(new_n11952_));
  INVX1    g11888(.A(new_n11854_), .Y(new_n11953_));
  OAI21X1  g11889(.A0(new_n11953_), .A1(new_n11952_), .B0(new_n11855_), .Y(new_n11954_));
  OR2X1    g11890(.A(new_n11854_), .B(new_n11850_), .Y(new_n11955_));
  INVX1    g11891(.A(new_n11859_), .Y(new_n11956_));
  AOI21X1  g11892(.A0(new_n11955_), .A1(new_n11954_), .B0(new_n11956_), .Y(new_n11957_));
  NAND3X1  g11893(.A(new_n11956_), .B(new_n11955_), .C(new_n11954_), .Y(new_n11958_));
  INVX1    g11894(.A(new_n11865_), .Y(new_n11959_));
  AOI21X1  g11895(.A0(new_n11959_), .A1(new_n11958_), .B0(new_n11957_), .Y(new_n11960_));
  AOI22X1  g11896(.A0(new_n7364_), .A1(new_n6300_), .B0(new_n7044_), .B1(new_n5970_), .Y(new_n11961_));
  OAI21X1  g11897(.A0(new_n7504_), .A1(new_n6309_), .B0(new_n11961_), .Y(new_n11962_));
  AOI21X1  g11898(.A0(new_n7552_), .A1(new_n5972_), .B0(new_n11962_), .Y(new_n11963_));
  XOR2X1   g11899(.A(new_n11963_), .B(\a[2] ), .Y(new_n11964_));
  AOI21X1  g11900(.A0(new_n11960_), .A1(new_n11868_), .B0(new_n11964_), .Y(new_n11965_));
  XOR2X1   g11901(.A(new_n11619_), .B(new_n11615_), .Y(new_n11966_));
  OAI21X1  g11902(.A0(new_n11965_), .A1(new_n11867_), .B0(new_n11966_), .Y(new_n11967_));
  XOR2X1   g11903(.A(new_n11612_), .B(new_n3431_), .Y(new_n11968_));
  XOR2X1   g11904(.A(new_n11968_), .B(new_n11609_), .Y(new_n11969_));
  AOI21X1  g11905(.A0(new_n11967_), .A1(new_n11621_), .B0(new_n11969_), .Y(new_n11970_));
  XOR2X1   g11906(.A(new_n11606_), .B(new_n11602_), .Y(new_n11971_));
  OAI21X1  g11907(.A0(new_n11970_), .A1(new_n11614_), .B0(new_n11971_), .Y(new_n11972_));
  XOR2X1   g11908(.A(new_n11599_), .B(new_n3431_), .Y(new_n11973_));
  XOR2X1   g11909(.A(new_n11973_), .B(new_n11596_), .Y(new_n11974_));
  AOI21X1  g11910(.A0(new_n11972_), .A1(new_n11608_), .B0(new_n11974_), .Y(new_n11975_));
  XOR2X1   g11911(.A(new_n11594_), .B(new_n11590_), .Y(new_n11976_));
  OAI21X1  g11912(.A0(new_n11975_), .A1(new_n11601_), .B0(new_n11976_), .Y(new_n11977_));
  XOR2X1   g11913(.A(new_n11586_), .B(new_n3431_), .Y(new_n11978_));
  XOR2X1   g11914(.A(new_n11978_), .B(new_n11582_), .Y(new_n11979_));
  AOI21X1  g11915(.A0(new_n11977_), .A1(new_n11595_), .B0(new_n11979_), .Y(new_n11980_));
  XOR2X1   g11916(.A(new_n11580_), .B(new_n11576_), .Y(new_n11981_));
  OAI21X1  g11917(.A0(new_n11980_), .A1(new_n11588_), .B0(new_n11981_), .Y(new_n11982_));
  XOR2X1   g11918(.A(new_n11572_), .B(\a[2] ), .Y(new_n11983_));
  XOR2X1   g11919(.A(new_n11983_), .B(new_n11569_), .Y(new_n11984_));
  AOI21X1  g11920(.A0(new_n11982_), .A1(new_n11581_), .B0(new_n11984_), .Y(new_n11985_));
  XOR2X1   g11921(.A(new_n11567_), .B(new_n11563_), .Y(new_n11986_));
  OAI21X1  g11922(.A0(new_n11985_), .A1(new_n11574_), .B0(new_n11986_), .Y(new_n11987_));
  AOI21X1  g11923(.A0(new_n11987_), .A1(new_n11568_), .B0(new_n11562_), .Y(new_n11988_));
  OR2X1    g11924(.A(new_n11988_), .B(new_n11560_), .Y(new_n11989_));
  AOI21X1  g11925(.A0(new_n11989_), .A1(new_n11226_), .B0(new_n11225_), .Y(new_n11990_));
  OAI21X1  g11926(.A0(new_n11990_), .A1(new_n11202_), .B0(new_n11201_), .Y(new_n11991_));
  AOI21X1  g11927(.A0(new_n11991_), .A1(new_n10861_), .B0(new_n10860_), .Y(new_n11992_));
  AND2X1   g11928(.A(new_n10541_), .B(new_n10538_), .Y(new_n11993_));
  XOR2X1   g11929(.A(new_n10543_), .B(new_n11993_), .Y(new_n11994_));
  OAI21X1  g11930(.A0(new_n11994_), .A1(new_n11992_), .B0(new_n10544_), .Y(new_n11995_));
  AOI21X1  g11931(.A0(new_n11995_), .A1(new_n10242_), .B0(new_n10241_), .Y(new_n11996_));
  OAI21X1  g11932(.A0(new_n11996_), .A1(new_n9968_), .B0(new_n9966_), .Y(new_n11997_));
  XOR2X1   g11933(.A(new_n9690_), .B(new_n9689_), .Y(new_n11998_));
  AOI21X1  g11934(.A0(new_n11998_), .A1(new_n11997_), .B0(new_n9691_), .Y(new_n11999_));
  OAI21X1  g11935(.A0(new_n11999_), .A1(new_n9461_), .B0(new_n9459_), .Y(new_n12000_));
  AOI21X1  g11936(.A0(new_n12000_), .A1(new_n9228_), .B0(new_n9227_), .Y(new_n12001_));
  XOR2X1   g11937(.A(new_n9036_), .B(new_n9035_), .Y(new_n12002_));
  INVX1    g11938(.A(new_n12002_), .Y(new_n12003_));
  OAI21X1  g11939(.A0(new_n12003_), .A1(new_n12001_), .B0(new_n9038_), .Y(new_n12004_));
  AOI21X1  g11940(.A0(new_n12004_), .A1(new_n8944_), .B0(new_n8943_), .Y(new_n12005_));
  OAI21X1  g11941(.A0(new_n12005_), .A1(new_n8860_), .B0(new_n8858_), .Y(new_n12006_));
  XOR2X1   g11942(.A(new_n8513_), .B(new_n8512_), .Y(new_n12007_));
  AOI21X1  g11943(.A0(new_n12007_), .A1(new_n12006_), .B0(new_n8514_), .Y(new_n12008_));
  OAI21X1  g11944(.A0(new_n12008_), .A1(new_n8439_), .B0(new_n8438_), .Y(new_n12009_));
  AOI21X1  g11945(.A0(new_n12009_), .A1(new_n8267_), .B0(new_n8266_), .Y(new_n12010_));
  XOR2X1   g11946(.A(new_n8133_), .B(new_n8132_), .Y(new_n12011_));
  INVX1    g11947(.A(new_n12011_), .Y(new_n12012_));
  OAI21X1  g11948(.A0(new_n12012_), .A1(new_n12010_), .B0(new_n8135_), .Y(new_n12013_));
  AOI21X1  g11949(.A0(new_n12013_), .A1(new_n8058_), .B0(new_n8056_), .Y(new_n12014_));
  OAI21X1  g11950(.A0(new_n12014_), .A1(new_n8001_), .B0(new_n7999_), .Y(new_n12015_));
  XOR2X1   g11951(.A(new_n7818_), .B(new_n7817_), .Y(new_n12016_));
  AOI21X1  g11952(.A0(new_n12016_), .A1(new_n12015_), .B0(new_n7819_), .Y(new_n12017_));
  XOR2X1   g11953(.A(new_n12017_), .B(new_n7730_), .Y(new_n12018_));
  AND2X1   g11954(.A(new_n7556_), .B(new_n7546_), .Y(new_n12019_));
  INVX1    g11955(.A(new_n12019_), .Y(new_n12020_));
  OAI21X1  g11956(.A0(new_n7568_), .A1(new_n7557_), .B0(new_n12020_), .Y(new_n12021_));
  NOR2X1   g11957(.A(new_n7550_), .B(new_n7070_), .Y(new_n12022_));
  NOR2X1   g11958(.A(new_n7555_), .B(new_n7551_), .Y(new_n12023_));
  NOR2X1   g11959(.A(new_n12023_), .B(new_n12022_), .Y(new_n12024_));
  INVX1    g11960(.A(new_n2811_), .Y(new_n12025_));
  OR4X1    g11961(.A(new_n2089_), .B(new_n874_), .C(new_n460_), .D(new_n358_), .Y(new_n12026_));
  OR4X1    g11962(.A(new_n938_), .B(new_n505_), .C(new_n869_), .D(new_n678_), .Y(new_n12027_));
  OR4X1    g11963(.A(new_n12027_), .B(new_n513_), .C(new_n137_), .D(new_n928_), .Y(new_n12028_));
  NOR4X1   g11964(.A(new_n12028_), .B(new_n12026_), .C(new_n12025_), .D(new_n2275_), .Y(new_n12029_));
  INVX1    g11965(.A(new_n12029_), .Y(new_n12030_));
  OR4X1    g11966(.A(new_n2302_), .B(new_n1415_), .C(new_n480_), .D(new_n133_), .Y(new_n12031_));
  NAND3X1  g11967(.A(new_n719_), .B(new_n862_), .C(new_n469_), .Y(new_n12032_));
  OR4X1    g11968(.A(new_n12032_), .B(new_n12031_), .C(new_n785_), .D(new_n128_), .Y(new_n12033_));
  OR4X1    g11969(.A(new_n12033_), .B(new_n6767_), .C(new_n3282_), .D(new_n2118_), .Y(new_n12034_));
  NOR4X1   g11970(.A(new_n12034_), .B(new_n12030_), .C(new_n2539_), .D(new_n212_), .Y(new_n12035_));
  XOR2X1   g11971(.A(new_n12035_), .B(new_n7070_), .Y(new_n12036_));
  NOR2X1   g11972(.A(new_n12036_), .B(new_n12024_), .Y(new_n12037_));
  AND2X1   g11973(.A(new_n12035_), .B(new_n7070_), .Y(new_n12038_));
  NOR2X1   g11974(.A(new_n12035_), .B(new_n7070_), .Y(new_n12039_));
  NOR4X1   g11975(.A(new_n12039_), .B(new_n12038_), .C(new_n12023_), .D(new_n12022_), .Y(new_n12040_));
  NOR2X1   g11976(.A(new_n12040_), .B(new_n12037_), .Y(new_n12041_));
  AOI22X1  g11977(.A0(new_n7485_), .A1(new_n1884_), .B0(new_n7364_), .B1(new_n1890_), .Y(new_n12042_));
  OAI21X1  g11978(.A0(new_n7523_), .A1(new_n3498_), .B0(new_n12042_), .Y(new_n12043_));
  AOI21X1  g11979(.A0(new_n7612_), .A1(new_n407_), .B0(new_n12043_), .Y(new_n12044_));
  XOR2X1   g11980(.A(new_n12044_), .B(new_n12041_), .Y(new_n12045_));
  OAI22X1  g11981(.A0(new_n7581_), .A1(new_n2431_), .B0(new_n7537_), .B1(new_n2186_), .Y(new_n12046_));
  AOI21X1  g11982(.A0(new_n7571_), .A1(new_n2139_), .B0(new_n12046_), .Y(new_n12047_));
  OAI21X1  g11983(.A0(new_n7621_), .A1(new_n2063_), .B0(new_n12047_), .Y(new_n12048_));
  XOR2X1   g11984(.A(new_n12048_), .B(new_n74_), .Y(new_n12049_));
  INVX1    g11985(.A(new_n12049_), .Y(new_n12050_));
  XOR2X1   g11986(.A(new_n12050_), .B(new_n12045_), .Y(new_n12051_));
  XOR2X1   g11987(.A(new_n12051_), .B(new_n12021_), .Y(new_n12052_));
  AOI22X1  g11988(.A0(new_n7590_), .A1(new_n2418_), .B0(new_n7578_), .B1(new_n2424_), .Y(new_n12053_));
  OAI21X1  g11989(.A0(new_n7642_), .A1(new_n2626_), .B0(new_n12053_), .Y(new_n12054_));
  AOI21X1  g11990(.A0(new_n7712_), .A1(new_n2301_), .B0(new_n12054_), .Y(new_n12055_));
  XOR2X1   g11991(.A(new_n12055_), .B(\a[26] ), .Y(new_n12056_));
  XOR2X1   g11992(.A(new_n12056_), .B(new_n12052_), .Y(new_n12057_));
  AND2X1   g11993(.A(new_n7569_), .B(new_n7542_), .Y(new_n12058_));
  INVX1    g11994(.A(new_n7598_), .Y(new_n12059_));
  AOI21X1  g11995(.A0(new_n12059_), .A1(new_n7570_), .B0(new_n12058_), .Y(new_n12060_));
  MX2X1    g11996(.A(new_n2653_), .B(new_n2654_), .S0(new_n2655_), .Y(new_n12061_));
  AOI22X1  g11997(.A0(new_n12061_), .A1(new_n7341_), .B0(new_n7643_), .B1(new_n2657_), .Y(new_n12062_));
  OAI21X1  g11998(.A0(new_n7808_), .A1(new_n2692_), .B0(new_n12062_), .Y(new_n12063_));
  XOR2X1   g11999(.A(new_n12063_), .B(new_n70_), .Y(new_n12064_));
  XOR2X1   g12000(.A(new_n12064_), .B(new_n12060_), .Y(new_n12065_));
  XOR2X1   g12001(.A(new_n12065_), .B(new_n12057_), .Y(new_n12066_));
  NOR2X1   g12002(.A(new_n7630_), .B(new_n7599_), .Y(new_n12067_));
  INVX1    g12003(.A(new_n7661_), .Y(new_n12068_));
  AOI21X1  g12004(.A0(new_n12068_), .A1(new_n7631_), .B0(new_n12067_), .Y(new_n12069_));
  XOR2X1   g12005(.A(new_n12069_), .B(new_n12066_), .Y(new_n12070_));
  NOR2X1   g12006(.A(new_n7728_), .B(new_n7662_), .Y(new_n12071_));
  INVX1    g12007(.A(new_n12071_), .Y(new_n12072_));
  OAI21X1  g12008(.A0(new_n12017_), .A1(new_n7730_), .B0(new_n12072_), .Y(new_n12073_));
  XOR2X1   g12009(.A(new_n12073_), .B(new_n12070_), .Y(new_n12074_));
  AND2X1   g12010(.A(new_n12074_), .B(new_n12018_), .Y(new_n12075_));
  XOR2X1   g12011(.A(new_n12016_), .B(new_n12015_), .Y(new_n12076_));
  AND2X1   g12012(.A(new_n12076_), .B(new_n12018_), .Y(new_n12077_));
  INVX1    g12013(.A(new_n12077_), .Y(new_n12078_));
  XOR2X1   g12014(.A(new_n12014_), .B(new_n8001_), .Y(new_n12079_));
  AND2X1   g12015(.A(new_n12079_), .B(new_n12076_), .Y(new_n12080_));
  XOR2X1   g12016(.A(new_n12013_), .B(new_n8058_), .Y(new_n12081_));
  NAND2X1  g12017(.A(new_n12081_), .B(new_n12079_), .Y(new_n12082_));
  XOR2X1   g12018(.A(new_n12012_), .B(new_n12010_), .Y(new_n12083_));
  AND2X1   g12019(.A(new_n12083_), .B(new_n12081_), .Y(new_n12084_));
  XOR2X1   g12020(.A(new_n12009_), .B(new_n8267_), .Y(new_n12085_));
  AND2X1   g12021(.A(new_n12085_), .B(new_n12083_), .Y(new_n12086_));
  INVX1    g12022(.A(new_n12086_), .Y(new_n12087_));
  XOR2X1   g12023(.A(new_n12008_), .B(new_n8439_), .Y(new_n12088_));
  AND2X1   g12024(.A(new_n12088_), .B(new_n12085_), .Y(new_n12089_));
  XOR2X1   g12025(.A(new_n12007_), .B(new_n12006_), .Y(new_n12090_));
  AND2X1   g12026(.A(new_n12090_), .B(new_n12088_), .Y(new_n12091_));
  INVX1    g12027(.A(new_n12091_), .Y(new_n12092_));
  XOR2X1   g12028(.A(new_n12005_), .B(new_n8860_), .Y(new_n12093_));
  AND2X1   g12029(.A(new_n12093_), .B(new_n12090_), .Y(new_n12094_));
  XOR2X1   g12030(.A(new_n12004_), .B(new_n8944_), .Y(new_n12095_));
  NAND2X1  g12031(.A(new_n12095_), .B(new_n12093_), .Y(new_n12096_));
  XOR2X1   g12032(.A(new_n12003_), .B(new_n12001_), .Y(new_n12097_));
  AND2X1   g12033(.A(new_n12097_), .B(new_n12095_), .Y(new_n12098_));
  XOR2X1   g12034(.A(new_n12000_), .B(new_n9228_), .Y(new_n12099_));
  AND2X1   g12035(.A(new_n12099_), .B(new_n12097_), .Y(new_n12100_));
  INVX1    g12036(.A(new_n12100_), .Y(new_n12101_));
  XOR2X1   g12037(.A(new_n11999_), .B(new_n9461_), .Y(new_n12102_));
  AND2X1   g12038(.A(new_n12102_), .B(new_n12099_), .Y(new_n12103_));
  XOR2X1   g12039(.A(new_n11998_), .B(new_n11997_), .Y(new_n12104_));
  AND2X1   g12040(.A(new_n12104_), .B(new_n12102_), .Y(new_n12105_));
  INVX1    g12041(.A(new_n12105_), .Y(new_n12106_));
  XOR2X1   g12042(.A(new_n11996_), .B(new_n9968_), .Y(new_n12107_));
  AND2X1   g12043(.A(new_n12107_), .B(new_n12104_), .Y(new_n12108_));
  INVX1    g12044(.A(new_n12107_), .Y(new_n12109_));
  INVX1    g12045(.A(new_n11995_), .Y(new_n12110_));
  XOR2X1   g12046(.A(new_n12110_), .B(new_n10242_), .Y(new_n12111_));
  INVX1    g12047(.A(new_n11992_), .Y(new_n12112_));
  XOR2X1   g12048(.A(new_n11994_), .B(new_n12112_), .Y(new_n12113_));
  NOR2X1   g12049(.A(new_n12113_), .B(new_n12111_), .Y(new_n12114_));
  INVX1    g12050(.A(new_n12114_), .Y(new_n12115_));
  INVX1    g12051(.A(new_n11991_), .Y(new_n12116_));
  XOR2X1   g12052(.A(new_n12116_), .B(new_n10861_), .Y(new_n12117_));
  NOR2X1   g12053(.A(new_n12117_), .B(new_n12113_), .Y(new_n12118_));
  NAND3X1  g12054(.A(new_n10857_), .B(new_n10853_), .C(new_n10872_), .Y(new_n12119_));
  OAI21X1  g12055(.A0(new_n10870_), .A1(new_n10852_), .B0(new_n10858_), .Y(new_n12120_));
  INVX1    g12056(.A(new_n11200_), .Y(new_n12121_));
  NAND3X1  g12057(.A(new_n12121_), .B(new_n12120_), .C(new_n12119_), .Y(new_n12122_));
  NOR3X1   g12058(.A(new_n11208_), .B(new_n11195_), .C(new_n11207_), .Y(new_n12123_));
  AOI21X1  g12059(.A0(new_n11205_), .A1(new_n11194_), .B0(new_n11199_), .Y(new_n12124_));
  NAND2X1  g12060(.A(new_n11223_), .B(new_n11217_), .Y(new_n12125_));
  OAI21X1  g12061(.A0(new_n12124_), .A1(new_n12123_), .B0(new_n12125_), .Y(new_n12126_));
  NOR3X1   g12062(.A(new_n12125_), .B(new_n12124_), .C(new_n12123_), .Y(new_n12127_));
  NOR2X1   g12063(.A(new_n11988_), .B(new_n11560_), .Y(new_n12128_));
  OAI21X1  g12064(.A0(new_n12128_), .A1(new_n12127_), .B0(new_n12126_), .Y(new_n12129_));
  NAND3X1  g12065(.A(new_n12129_), .B(new_n12122_), .C(new_n11201_), .Y(new_n12130_));
  AOI21X1  g12066(.A0(new_n12120_), .A1(new_n12119_), .B0(new_n12121_), .Y(new_n12131_));
  OAI21X1  g12067(.A0(new_n11202_), .A1(new_n12131_), .B0(new_n11990_), .Y(new_n12132_));
  AND2X1   g12068(.A(new_n12132_), .B(new_n12130_), .Y(new_n12133_));
  INVX1    g12069(.A(new_n12133_), .Y(new_n12134_));
  OR2X1    g12070(.A(new_n12134_), .B(new_n12117_), .Y(new_n12135_));
  NAND3X1  g12071(.A(new_n11989_), .B(new_n11226_), .C(new_n12126_), .Y(new_n12136_));
  OAI21X1  g12072(.A0(new_n12127_), .A1(new_n11225_), .B0(new_n12128_), .Y(new_n12137_));
  AND2X1   g12073(.A(new_n12137_), .B(new_n12136_), .Y(new_n12138_));
  AND2X1   g12074(.A(new_n12138_), .B(new_n12133_), .Y(new_n12139_));
  AND2X1   g12075(.A(new_n11987_), .B(new_n11568_), .Y(new_n12140_));
  XOR2X1   g12076(.A(new_n12140_), .B(new_n11562_), .Y(new_n12141_));
  NAND3X1  g12077(.A(new_n12141_), .B(new_n12137_), .C(new_n12136_), .Y(new_n12142_));
  OR2X1    g12078(.A(new_n11985_), .B(new_n11574_), .Y(new_n12143_));
  XOR2X1   g12079(.A(new_n11986_), .B(new_n12143_), .Y(new_n12144_));
  AND2X1   g12080(.A(new_n12144_), .B(new_n12141_), .Y(new_n12145_));
  NAND2X1  g12081(.A(new_n11982_), .B(new_n11581_), .Y(new_n12146_));
  INVX1    g12082(.A(new_n11984_), .Y(new_n12147_));
  XOR2X1   g12083(.A(new_n12147_), .B(new_n12146_), .Y(new_n12148_));
  NAND2X1  g12084(.A(new_n12148_), .B(new_n12144_), .Y(new_n12149_));
  OR2X1    g12085(.A(new_n11980_), .B(new_n11588_), .Y(new_n12150_));
  XOR2X1   g12086(.A(new_n11981_), .B(new_n12150_), .Y(new_n12151_));
  AND2X1   g12087(.A(new_n12151_), .B(new_n12148_), .Y(new_n12152_));
  NAND2X1  g12088(.A(new_n11977_), .B(new_n11595_), .Y(new_n12153_));
  INVX1    g12089(.A(new_n11979_), .Y(new_n12154_));
  XOR2X1   g12090(.A(new_n12154_), .B(new_n12153_), .Y(new_n12155_));
  NAND2X1  g12091(.A(new_n12155_), .B(new_n12151_), .Y(new_n12156_));
  OR2X1    g12092(.A(new_n11975_), .B(new_n11601_), .Y(new_n12157_));
  XOR2X1   g12093(.A(new_n11976_), .B(new_n12157_), .Y(new_n12158_));
  AND2X1   g12094(.A(new_n12158_), .B(new_n12155_), .Y(new_n12159_));
  NAND2X1  g12095(.A(new_n11972_), .B(new_n11608_), .Y(new_n12160_));
  INVX1    g12096(.A(new_n11974_), .Y(new_n12161_));
  XOR2X1   g12097(.A(new_n12161_), .B(new_n12160_), .Y(new_n12162_));
  NAND2X1  g12098(.A(new_n12162_), .B(new_n12158_), .Y(new_n12163_));
  OR2X1    g12099(.A(new_n11970_), .B(new_n11614_), .Y(new_n12164_));
  XOR2X1   g12100(.A(new_n11971_), .B(new_n12164_), .Y(new_n12165_));
  AND2X1   g12101(.A(new_n12165_), .B(new_n12162_), .Y(new_n12166_));
  NOR2X1   g12102(.A(new_n11970_), .B(new_n11614_), .Y(new_n12167_));
  XOR2X1   g12103(.A(new_n11971_), .B(new_n12167_), .Y(new_n12168_));
  NAND2X1  g12104(.A(new_n11967_), .B(new_n11621_), .Y(new_n12169_));
  XOR2X1   g12105(.A(new_n11969_), .B(new_n12169_), .Y(new_n12170_));
  OAI21X1  g12106(.A0(new_n11965_), .A1(new_n11867_), .B0(new_n11967_), .Y(new_n12171_));
  NAND2X1  g12107(.A(new_n11866_), .B(new_n11622_), .Y(new_n12172_));
  INVX1    g12108(.A(new_n11964_), .Y(new_n12173_));
  OAI21X1  g12109(.A0(new_n11866_), .A1(new_n11622_), .B0(new_n12173_), .Y(new_n12174_));
  NAND3X1  g12110(.A(new_n11966_), .B(new_n12174_), .C(new_n12172_), .Y(new_n12175_));
  AND2X1   g12111(.A(new_n12175_), .B(new_n12171_), .Y(new_n12176_));
  AOI21X1  g12112(.A0(new_n12176_), .A1(new_n12168_), .B0(new_n12170_), .Y(new_n12177_));
  XOR2X1   g12113(.A(new_n12165_), .B(new_n12162_), .Y(new_n12178_));
  AOI21X1  g12114(.A0(new_n12178_), .A1(new_n12177_), .B0(new_n12166_), .Y(new_n12179_));
  NOR2X1   g12115(.A(new_n12162_), .B(new_n12158_), .Y(new_n12180_));
  OAI21X1  g12116(.A0(new_n12180_), .A1(new_n12179_), .B0(new_n12163_), .Y(new_n12181_));
  XOR2X1   g12117(.A(new_n12158_), .B(new_n12155_), .Y(new_n12182_));
  AND2X1   g12118(.A(new_n12182_), .B(new_n12181_), .Y(new_n12183_));
  XOR2X1   g12119(.A(new_n12155_), .B(new_n12151_), .Y(new_n12184_));
  OAI21X1  g12120(.A0(new_n12183_), .A1(new_n12159_), .B0(new_n12184_), .Y(new_n12185_));
  XOR2X1   g12121(.A(new_n11984_), .B(new_n12146_), .Y(new_n12186_));
  XOR2X1   g12122(.A(new_n12151_), .B(new_n12186_), .Y(new_n12187_));
  AOI21X1  g12123(.A0(new_n12185_), .A1(new_n12156_), .B0(new_n12187_), .Y(new_n12188_));
  XOR2X1   g12124(.A(new_n12148_), .B(new_n12144_), .Y(new_n12189_));
  OAI21X1  g12125(.A0(new_n12188_), .A1(new_n12152_), .B0(new_n12189_), .Y(new_n12190_));
  NOR2X1   g12126(.A(new_n11985_), .B(new_n11574_), .Y(new_n12191_));
  XOR2X1   g12127(.A(new_n11986_), .B(new_n12191_), .Y(new_n12192_));
  XOR2X1   g12128(.A(new_n12192_), .B(new_n12141_), .Y(new_n12193_));
  AOI21X1  g12129(.A0(new_n12190_), .A1(new_n12149_), .B0(new_n12193_), .Y(new_n12194_));
  NOR2X1   g12130(.A(new_n12194_), .B(new_n12145_), .Y(new_n12195_));
  AOI21X1  g12131(.A0(new_n12137_), .A1(new_n12136_), .B0(new_n12141_), .Y(new_n12196_));
  OAI21X1  g12132(.A0(new_n12196_), .A1(new_n12195_), .B0(new_n12142_), .Y(new_n12197_));
  XOR2X1   g12133(.A(new_n12138_), .B(new_n12133_), .Y(new_n12198_));
  AND2X1   g12134(.A(new_n12198_), .B(new_n12197_), .Y(new_n12199_));
  XOR2X1   g12135(.A(new_n12134_), .B(new_n12117_), .Y(new_n12200_));
  OAI21X1  g12136(.A0(new_n12199_), .A1(new_n12139_), .B0(new_n12200_), .Y(new_n12201_));
  NAND2X1  g12137(.A(new_n12201_), .B(new_n12135_), .Y(new_n12202_));
  AND2X1   g12138(.A(new_n12117_), .B(new_n12113_), .Y(new_n12203_));
  INVX1    g12139(.A(new_n12203_), .Y(new_n12204_));
  AOI21X1  g12140(.A0(new_n12204_), .A1(new_n12202_), .B0(new_n12118_), .Y(new_n12205_));
  AND2X1   g12141(.A(new_n12113_), .B(new_n12111_), .Y(new_n12206_));
  OAI21X1  g12142(.A0(new_n12206_), .A1(new_n12205_), .B0(new_n12115_), .Y(new_n12207_));
  INVX1    g12143(.A(new_n12111_), .Y(new_n12208_));
  XOR2X1   g12144(.A(new_n12208_), .B(new_n12107_), .Y(new_n12209_));
  NAND2X1  g12145(.A(new_n12209_), .B(new_n12207_), .Y(new_n12210_));
  OAI21X1  g12146(.A0(new_n12111_), .A1(new_n12109_), .B0(new_n12210_), .Y(new_n12211_));
  NOR2X1   g12147(.A(new_n12107_), .B(new_n12104_), .Y(new_n12212_));
  INVX1    g12148(.A(new_n12212_), .Y(new_n12213_));
  AOI21X1  g12149(.A0(new_n12213_), .A1(new_n12211_), .B0(new_n12108_), .Y(new_n12214_));
  NOR2X1   g12150(.A(new_n12104_), .B(new_n12102_), .Y(new_n12215_));
  OAI21X1  g12151(.A0(new_n12215_), .A1(new_n12214_), .B0(new_n12106_), .Y(new_n12216_));
  XOR2X1   g12152(.A(new_n12102_), .B(new_n12099_), .Y(new_n12217_));
  AOI21X1  g12153(.A0(new_n12217_), .A1(new_n12216_), .B0(new_n12103_), .Y(new_n12218_));
  NOR2X1   g12154(.A(new_n12099_), .B(new_n12097_), .Y(new_n12219_));
  OAI21X1  g12155(.A0(new_n12219_), .A1(new_n12218_), .B0(new_n12101_), .Y(new_n12220_));
  OR2X1    g12156(.A(new_n12097_), .B(new_n12095_), .Y(new_n12221_));
  AOI21X1  g12157(.A0(new_n12221_), .A1(new_n12220_), .B0(new_n12098_), .Y(new_n12222_));
  XOR2X1   g12158(.A(new_n12095_), .B(new_n12093_), .Y(new_n12223_));
  INVX1    g12159(.A(new_n12223_), .Y(new_n12224_));
  OAI21X1  g12160(.A0(new_n12224_), .A1(new_n12222_), .B0(new_n12096_), .Y(new_n12225_));
  OR2X1    g12161(.A(new_n12093_), .B(new_n12090_), .Y(new_n12226_));
  AOI21X1  g12162(.A0(new_n12226_), .A1(new_n12225_), .B0(new_n12094_), .Y(new_n12227_));
  NOR2X1   g12163(.A(new_n12090_), .B(new_n12088_), .Y(new_n12228_));
  OAI21X1  g12164(.A0(new_n12228_), .A1(new_n12227_), .B0(new_n12092_), .Y(new_n12229_));
  XOR2X1   g12165(.A(new_n12088_), .B(new_n12085_), .Y(new_n12230_));
  AOI21X1  g12166(.A0(new_n12230_), .A1(new_n12229_), .B0(new_n12089_), .Y(new_n12231_));
  NOR2X1   g12167(.A(new_n12085_), .B(new_n12083_), .Y(new_n12232_));
  OAI21X1  g12168(.A0(new_n12232_), .A1(new_n12231_), .B0(new_n12087_), .Y(new_n12233_));
  XOR2X1   g12169(.A(new_n12083_), .B(new_n12081_), .Y(new_n12234_));
  AOI21X1  g12170(.A0(new_n12234_), .A1(new_n12233_), .B0(new_n12084_), .Y(new_n12235_));
  NOR2X1   g12171(.A(new_n12081_), .B(new_n12079_), .Y(new_n12236_));
  OAI21X1  g12172(.A0(new_n12236_), .A1(new_n12235_), .B0(new_n12082_), .Y(new_n12237_));
  XOR2X1   g12173(.A(new_n12079_), .B(new_n12076_), .Y(new_n12238_));
  AOI21X1  g12174(.A0(new_n12238_), .A1(new_n12237_), .B0(new_n12080_), .Y(new_n12239_));
  NOR2X1   g12175(.A(new_n12076_), .B(new_n12018_), .Y(new_n12240_));
  OAI21X1  g12176(.A0(new_n12240_), .A1(new_n12239_), .B0(new_n12078_), .Y(new_n12241_));
  XOR2X1   g12177(.A(new_n12074_), .B(new_n12018_), .Y(new_n12242_));
  AOI21X1  g12178(.A0(new_n12242_), .A1(new_n12241_), .B0(new_n12075_), .Y(new_n12243_));
  NOR2X1   g12179(.A(new_n12069_), .B(new_n12066_), .Y(new_n12244_));
  AOI21X1  g12180(.A0(new_n12073_), .A1(new_n12070_), .B0(new_n12244_), .Y(new_n12245_));
  INVX1    g12181(.A(new_n12057_), .Y(new_n12246_));
  NOR2X1   g12182(.A(new_n12064_), .B(new_n12060_), .Y(new_n12247_));
  AOI21X1  g12183(.A0(new_n12065_), .A1(new_n12246_), .B0(new_n12247_), .Y(new_n12248_));
  AND2X1   g12184(.A(new_n12051_), .B(new_n12021_), .Y(new_n12249_));
  INVX1    g12185(.A(new_n12056_), .Y(new_n12250_));
  AOI21X1  g12186(.A0(new_n12250_), .A1(new_n12052_), .B0(new_n12249_), .Y(new_n12251_));
  AOI22X1  g12187(.A0(new_n7643_), .A1(new_n2423_), .B0(new_n7590_), .B1(new_n2424_), .Y(new_n12252_));
  OAI21X1  g12188(.A0(new_n7642_), .A1(new_n2419_), .B0(new_n12252_), .Y(new_n12253_));
  AOI21X1  g12189(.A0(new_n7718_), .A1(new_n2301_), .B0(new_n12253_), .Y(new_n12254_));
  XOR2X1   g12190(.A(new_n12254_), .B(\a[26] ), .Y(new_n12255_));
  XOR2X1   g12191(.A(new_n12255_), .B(new_n12251_), .Y(new_n12256_));
  INVX1    g12192(.A(new_n12038_), .Y(new_n12257_));
  OAI21X1  g12193(.A0(new_n12039_), .A1(new_n12024_), .B0(new_n12257_), .Y(new_n12258_));
  OR4X1    g12194(.A(new_n2745_), .B(new_n2696_), .C(new_n2658_), .D(new_n2657_), .Y(new_n12259_));
  AND2X1   g12195(.A(new_n12259_), .B(new_n7341_), .Y(new_n12260_));
  XOR2X1   g12196(.A(new_n12260_), .B(new_n70_), .Y(new_n12261_));
  OR4X1    g12197(.A(new_n480_), .B(new_n282_), .C(new_n175_), .D(new_n338_), .Y(new_n12262_));
  OR4X1    g12198(.A(new_n12262_), .B(new_n3765_), .C(new_n3709_), .D(new_n508_), .Y(new_n12263_));
  OR4X1    g12199(.A(new_n1911_), .B(new_n1000_), .C(new_n766_), .D(new_n537_), .Y(new_n12264_));
  OR4X1    g12200(.A(new_n12264_), .B(new_n12263_), .C(new_n2789_), .D(new_n2261_), .Y(new_n12265_));
  NOR4X1   g12201(.A(new_n12265_), .B(new_n8726_), .C(new_n7926_), .D(new_n7433_), .Y(new_n12266_));
  XOR2X1   g12202(.A(new_n12266_), .B(new_n12035_), .Y(new_n12267_));
  XOR2X1   g12203(.A(new_n12267_), .B(new_n12261_), .Y(new_n12268_));
  XOR2X1   g12204(.A(new_n12268_), .B(new_n12258_), .Y(new_n12269_));
  AOI22X1  g12205(.A0(new_n7522_), .A1(new_n1884_), .B0(new_n7485_), .B1(new_n1890_), .Y(new_n12270_));
  OAI21X1  g12206(.A0(new_n7537_), .A1(new_n3498_), .B0(new_n12270_), .Y(new_n12271_));
  AOI21X1  g12207(.A0(new_n7536_), .A1(new_n407_), .B0(new_n12271_), .Y(new_n12272_));
  XOR2X1   g12208(.A(new_n12272_), .B(new_n12269_), .Y(new_n12273_));
  NOR2X1   g12209(.A(new_n12044_), .B(new_n12041_), .Y(new_n12274_));
  AOI21X1  g12210(.A0(new_n12050_), .A1(new_n12045_), .B0(new_n12274_), .Y(new_n12275_));
  XOR2X1   g12211(.A(new_n12275_), .B(new_n12273_), .Y(new_n12276_));
  AOI22X1  g12212(.A0(new_n7571_), .A1(new_n2095_), .B0(new_n7558_), .B1(new_n2185_), .Y(new_n12277_));
  OAI21X1  g12213(.A0(new_n7602_), .A1(new_n2140_), .B0(new_n12277_), .Y(new_n12278_));
  AOI21X1  g12214(.A0(new_n7601_), .A1(new_n2062_), .B0(new_n12278_), .Y(new_n12279_));
  XOR2X1   g12215(.A(new_n12279_), .B(\a[29] ), .Y(new_n12280_));
  XOR2X1   g12216(.A(new_n12280_), .B(new_n12276_), .Y(new_n12281_));
  XOR2X1   g12217(.A(new_n12281_), .B(new_n12256_), .Y(new_n12282_));
  XOR2X1   g12218(.A(new_n12282_), .B(new_n12248_), .Y(new_n12283_));
  INVX1    g12219(.A(new_n12283_), .Y(new_n12284_));
  XOR2X1   g12220(.A(new_n12284_), .B(new_n12245_), .Y(new_n12285_));
  NOR2X1   g12221(.A(new_n12285_), .B(new_n12074_), .Y(new_n12286_));
  XOR2X1   g12222(.A(new_n12285_), .B(new_n12074_), .Y(new_n12287_));
  AND2X1   g12223(.A(new_n12285_), .B(new_n12074_), .Y(new_n12288_));
  INVX1    g12224(.A(new_n12288_), .Y(new_n12289_));
  OAI21X1  g12225(.A0(new_n12286_), .A1(new_n12243_), .B0(new_n12289_), .Y(new_n12290_));
  OAI22X1  g12226(.A0(new_n12290_), .A1(new_n12286_), .B0(new_n12287_), .B1(new_n12243_), .Y(new_n12291_));
  INVX1    g12227(.A(new_n12285_), .Y(new_n12292_));
  AOI22X1  g12228(.A0(new_n12074_), .A1(new_n5659_), .B0(new_n12018_), .B1(new_n5373_), .Y(new_n12293_));
  OAI21X1  g12229(.A0(new_n12292_), .A1(new_n5959_), .B0(new_n12293_), .Y(new_n12294_));
  AOI21X1  g12230(.A0(new_n12291_), .A1(new_n67_), .B0(new_n12294_), .Y(new_n12295_));
  XOR2X1   g12231(.A(new_n12295_), .B(\a[5] ), .Y(new_n12296_));
  XOR2X1   g12232(.A(new_n12230_), .B(new_n12229_), .Y(new_n12297_));
  INVX1    g12233(.A(new_n12085_), .Y(new_n12298_));
  AOI22X1  g12234(.A0(new_n12090_), .A1(new_n4078_), .B0(new_n12088_), .B1(new_n4247_), .Y(new_n12299_));
  OAI21X1  g12235(.A0(new_n12298_), .A1(new_n4427_), .B0(new_n12299_), .Y(new_n12300_));
  AOI21X1  g12236(.A0(new_n12297_), .A1(new_n4080_), .B0(new_n12300_), .Y(new_n12301_));
  XOR2X1   g12237(.A(new_n12301_), .B(\a[11] ), .Y(new_n12302_));
  XOR2X1   g12238(.A(new_n12104_), .B(new_n12102_), .Y(new_n12303_));
  OR2X1    g12239(.A(new_n12303_), .B(new_n12214_), .Y(new_n12304_));
  OAI21X1  g12240(.A0(new_n12216_), .A1(new_n12215_), .B0(new_n12304_), .Y(new_n12305_));
  INVX1    g12241(.A(new_n12102_), .Y(new_n12306_));
  AOI22X1  g12242(.A0(new_n12107_), .A1(new_n3232_), .B0(new_n12104_), .B1(new_n3390_), .Y(new_n12307_));
  OAI21X1  g12243(.A0(new_n12306_), .A1(new_n3545_), .B0(new_n12307_), .Y(new_n12308_));
  AOI21X1  g12244(.A0(new_n12305_), .A1(new_n3234_), .B0(new_n12308_), .Y(new_n12309_));
  XOR2X1   g12245(.A(new_n12309_), .B(\a[17] ), .Y(new_n12310_));
  OR2X1    g12246(.A(new_n12194_), .B(new_n12145_), .Y(new_n12311_));
  XOR2X1   g12247(.A(new_n12141_), .B(new_n12138_), .Y(new_n12312_));
  XOR2X1   g12248(.A(new_n12312_), .B(new_n12311_), .Y(new_n12313_));
  INVX1    g12249(.A(new_n12138_), .Y(new_n12314_));
  AOI22X1  g12250(.A0(new_n12144_), .A1(new_n2657_), .B0(new_n12141_), .B1(new_n2696_), .Y(new_n12315_));
  OAI21X1  g12251(.A0(new_n12314_), .A1(new_n2753_), .B0(new_n12315_), .Y(new_n12316_));
  AOI21X1  g12252(.A0(new_n12313_), .A1(new_n2658_), .B0(new_n12316_), .Y(new_n12317_));
  XOR2X1   g12253(.A(new_n12317_), .B(\a[23] ), .Y(new_n12318_));
  AOI21X1  g12254(.A0(new_n12182_), .A1(new_n12181_), .B0(new_n12159_), .Y(new_n12319_));
  XOR2X1   g12255(.A(new_n12184_), .B(new_n12319_), .Y(new_n12320_));
  INVX1    g12256(.A(new_n12320_), .Y(new_n12321_));
  INVX1    g12257(.A(new_n12151_), .Y(new_n12322_));
  AOI22X1  g12258(.A0(new_n12158_), .A1(new_n2424_), .B0(new_n12155_), .B1(new_n2418_), .Y(new_n12323_));
  OAI21X1  g12259(.A0(new_n12322_), .A1(new_n2626_), .B0(new_n12323_), .Y(new_n12324_));
  AOI21X1  g12260(.A0(new_n12321_), .A1(new_n2301_), .B0(new_n12324_), .Y(new_n12325_));
  XOR2X1   g12261(.A(new_n12325_), .B(\a[26] ), .Y(new_n12326_));
  INVX1    g12262(.A(new_n12326_), .Y(new_n12327_));
  XOR2X1   g12263(.A(new_n12178_), .B(new_n12177_), .Y(new_n12328_));
  XOR2X1   g12264(.A(new_n11974_), .B(new_n12160_), .Y(new_n12329_));
  INVX1    g12265(.A(new_n11969_), .Y(new_n12330_));
  XOR2X1   g12266(.A(new_n12330_), .B(new_n12169_), .Y(new_n12331_));
  AOI22X1  g12267(.A0(new_n12331_), .A1(new_n2185_), .B0(new_n12165_), .B1(new_n2095_), .Y(new_n12332_));
  OAI21X1  g12268(.A0(new_n12329_), .A1(new_n2140_), .B0(new_n12332_), .Y(new_n12333_));
  AOI21X1  g12269(.A0(new_n12328_), .A1(new_n2062_), .B0(new_n12333_), .Y(new_n12334_));
  XOR2X1   g12270(.A(new_n12334_), .B(\a[29] ), .Y(new_n12335_));
  AOI21X1  g12271(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n2061_), .Y(new_n12336_));
  XOR2X1   g12272(.A(new_n12176_), .B(new_n12170_), .Y(new_n12337_));
  OAI22X1  g12273(.A0(new_n12176_), .A1(new_n2431_), .B0(new_n12170_), .B1(new_n2140_), .Y(new_n12338_));
  AOI21X1  g12274(.A0(new_n12337_), .A1(new_n2062_), .B0(new_n12338_), .Y(new_n12339_));
  XOR2X1   g12275(.A(new_n12339_), .B(\a[29] ), .Y(new_n12340_));
  OAI22X1  g12276(.A0(new_n12176_), .A1(new_n2186_), .B0(new_n12170_), .B1(new_n2431_), .Y(new_n12341_));
  AOI21X1  g12277(.A0(new_n12165_), .A1(new_n2139_), .B0(new_n12341_), .Y(new_n12342_));
  NAND2X1  g12278(.A(new_n12176_), .B(new_n12331_), .Y(new_n12343_));
  XOR2X1   g12279(.A(new_n12343_), .B(new_n12165_), .Y(new_n12344_));
  OAI21X1  g12280(.A0(new_n12344_), .A1(new_n2063_), .B0(new_n12342_), .Y(new_n12345_));
  NOR4X1   g12281(.A(new_n12345_), .B(new_n12340_), .C(new_n12336_), .D(new_n74_), .Y(new_n12346_));
  AOI21X1  g12282(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n4171_), .Y(new_n12347_));
  INVX1    g12283(.A(new_n12347_), .Y(new_n12348_));
  XOR2X1   g12284(.A(new_n12348_), .B(new_n12346_), .Y(new_n12349_));
  XOR2X1   g12285(.A(new_n12349_), .B(new_n12335_), .Y(new_n12350_));
  XOR2X1   g12286(.A(new_n12350_), .B(new_n12326_), .Y(new_n12351_));
  XOR2X1   g12287(.A(new_n12182_), .B(new_n12181_), .Y(new_n12352_));
  INVX1    g12288(.A(new_n12155_), .Y(new_n12353_));
  AOI22X1  g12289(.A0(new_n12162_), .A1(new_n2424_), .B0(new_n12158_), .B1(new_n2418_), .Y(new_n12354_));
  OAI21X1  g12290(.A0(new_n12353_), .A1(new_n2626_), .B0(new_n12354_), .Y(new_n12355_));
  AOI21X1  g12291(.A0(new_n12352_), .A1(new_n2301_), .B0(new_n12355_), .Y(new_n12356_));
  XOR2X1   g12292(.A(new_n12356_), .B(\a[26] ), .Y(new_n12357_));
  INVX1    g12293(.A(new_n12357_), .Y(new_n12358_));
  NOR3X1   g12294(.A(new_n12340_), .B(new_n12336_), .C(new_n74_), .Y(new_n12359_));
  XOR2X1   g12295(.A(new_n12345_), .B(\a[29] ), .Y(new_n12360_));
  XOR2X1   g12296(.A(new_n12360_), .B(new_n12359_), .Y(new_n12361_));
  XOR2X1   g12297(.A(new_n12361_), .B(new_n12357_), .Y(new_n12362_));
  NOR2X1   g12298(.A(new_n12336_), .B(new_n74_), .Y(new_n12363_));
  XOR2X1   g12299(.A(new_n12340_), .B(new_n12363_), .Y(new_n12364_));
  OAI22X1  g12300(.A0(new_n12168_), .A1(new_n2666_), .B0(new_n12329_), .B1(new_n2419_), .Y(new_n12365_));
  AOI21X1  g12301(.A0(new_n12158_), .A1(new_n2423_), .B0(new_n12365_), .Y(new_n12366_));
  XOR2X1   g12302(.A(new_n12162_), .B(new_n12158_), .Y(new_n12367_));
  XOR2X1   g12303(.A(new_n12367_), .B(new_n12179_), .Y(new_n12368_));
  OAI21X1  g12304(.A0(new_n12368_), .A1(new_n2665_), .B0(new_n12366_), .Y(new_n12369_));
  XOR2X1   g12305(.A(new_n12369_), .B(new_n89_), .Y(new_n12370_));
  NOR2X1   g12306(.A(new_n12370_), .B(new_n12364_), .Y(new_n12371_));
  AOI21X1  g12307(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n2299_), .Y(new_n12372_));
  OAI22X1  g12308(.A0(new_n12176_), .A1(new_n2419_), .B0(new_n12170_), .B1(new_n2626_), .Y(new_n12373_));
  AOI21X1  g12309(.A0(new_n12337_), .A1(new_n2301_), .B0(new_n12373_), .Y(new_n12374_));
  XOR2X1   g12310(.A(new_n12374_), .B(\a[26] ), .Y(new_n12375_));
  OAI22X1  g12311(.A0(new_n12176_), .A1(new_n2666_), .B0(new_n12170_), .B1(new_n2419_), .Y(new_n12376_));
  AOI21X1  g12312(.A0(new_n12165_), .A1(new_n2423_), .B0(new_n12376_), .Y(new_n12377_));
  OAI21X1  g12313(.A0(new_n12344_), .A1(new_n2665_), .B0(new_n12377_), .Y(new_n12378_));
  NOR4X1   g12314(.A(new_n12378_), .B(new_n12375_), .C(new_n12372_), .D(new_n89_), .Y(new_n12379_));
  NAND2X1  g12315(.A(new_n12379_), .B(new_n12336_), .Y(new_n12380_));
  XOR2X1   g12316(.A(new_n12379_), .B(new_n12336_), .Y(new_n12381_));
  INVX1    g12317(.A(new_n12381_), .Y(new_n12382_));
  AOI22X1  g12318(.A0(new_n12331_), .A1(new_n2424_), .B0(new_n12165_), .B1(new_n2418_), .Y(new_n12383_));
  OAI21X1  g12319(.A0(new_n12329_), .A1(new_n2626_), .B0(new_n12383_), .Y(new_n12384_));
  AOI21X1  g12320(.A0(new_n12328_), .A1(new_n2301_), .B0(new_n12384_), .Y(new_n12385_));
  XOR2X1   g12321(.A(new_n12385_), .B(\a[26] ), .Y(new_n12386_));
  OAI21X1  g12322(.A0(new_n12386_), .A1(new_n12382_), .B0(new_n12380_), .Y(new_n12387_));
  XOR2X1   g12323(.A(new_n12370_), .B(new_n12364_), .Y(new_n12388_));
  AOI21X1  g12324(.A0(new_n12388_), .A1(new_n12387_), .B0(new_n12371_), .Y(new_n12389_));
  NOR2X1   g12325(.A(new_n12389_), .B(new_n12362_), .Y(new_n12390_));
  AOI21X1  g12326(.A0(new_n12361_), .A1(new_n12358_), .B0(new_n12390_), .Y(new_n12391_));
  NOR2X1   g12327(.A(new_n12391_), .B(new_n12351_), .Y(new_n12392_));
  AOI21X1  g12328(.A0(new_n12350_), .A1(new_n12327_), .B0(new_n12392_), .Y(new_n12393_));
  XOR2X1   g12329(.A(new_n12329_), .B(new_n12158_), .Y(new_n12394_));
  XOR2X1   g12330(.A(new_n12394_), .B(new_n12179_), .Y(new_n12395_));
  INVX1    g12331(.A(new_n12158_), .Y(new_n12396_));
  AOI22X1  g12332(.A0(new_n12165_), .A1(new_n2185_), .B0(new_n12162_), .B1(new_n2095_), .Y(new_n12397_));
  OAI21X1  g12333(.A0(new_n12396_), .A1(new_n2140_), .B0(new_n12397_), .Y(new_n12398_));
  AOI21X1  g12334(.A0(new_n12395_), .A1(new_n2062_), .B0(new_n12398_), .Y(new_n12399_));
  XOR2X1   g12335(.A(new_n12399_), .B(\a[29] ), .Y(new_n12400_));
  INVX1    g12336(.A(new_n8646_), .Y(new_n12401_));
  NAND3X1  g12337(.A(new_n930_), .B(new_n2996_), .C(new_n349_), .Y(new_n12402_));
  OR4X1    g12338(.A(new_n423_), .B(new_n479_), .C(new_n757_), .D(new_n187_), .Y(new_n12403_));
  OR4X1    g12339(.A(new_n12403_), .B(new_n12402_), .C(new_n530_), .D(new_n464_), .Y(new_n12404_));
  OR4X1    g12340(.A(new_n12404_), .B(new_n1426_), .C(new_n1114_), .D(new_n786_), .Y(new_n12405_));
  OR4X1    g12341(.A(new_n426_), .B(new_n85_), .C(new_n1579_), .D(new_n1284_), .Y(new_n12406_));
  OR4X1    g12342(.A(new_n1452_), .B(new_n455_), .C(new_n265_), .D(new_n223_), .Y(new_n12407_));
  OR4X1    g12343(.A(new_n12407_), .B(new_n12406_), .C(new_n1467_), .D(new_n340_), .Y(new_n12408_));
  OR4X1    g12344(.A(new_n1000_), .B(new_n1094_), .C(new_n728_), .D(new_n701_), .Y(new_n12409_));
  OR4X1    g12345(.A(new_n12409_), .B(new_n12408_), .C(new_n8692_), .D(new_n883_), .Y(new_n12410_));
  NOR4X1   g12346(.A(new_n382_), .B(new_n372_), .C(new_n207_), .D(new_n307_), .Y(new_n12411_));
  NAND3X1  g12347(.A(new_n12411_), .B(new_n2448_), .C(new_n2401_), .Y(new_n12412_));
  OR4X1    g12348(.A(new_n1984_), .B(new_n1962_), .C(new_n1777_), .D(new_n1780_), .Y(new_n12413_));
  OR4X1    g12349(.A(new_n750_), .B(new_n659_), .C(new_n566_), .D(new_n559_), .Y(new_n12414_));
  OR4X1    g12350(.A(new_n12414_), .B(new_n12413_), .C(new_n12412_), .D(new_n7744_), .Y(new_n12415_));
  NOR4X1   g12351(.A(new_n12415_), .B(new_n12410_), .C(new_n12405_), .D(new_n12401_), .Y(new_n12416_));
  INVX1    g12352(.A(new_n12416_), .Y(new_n12417_));
  OAI22X1  g12353(.A0(new_n12176_), .A1(new_n1885_), .B0(new_n12170_), .B1(new_n3498_), .Y(new_n12418_));
  AOI21X1  g12354(.A0(new_n12337_), .A1(new_n407_), .B0(new_n12418_), .Y(new_n12419_));
  XOR2X1   g12355(.A(new_n12419_), .B(new_n12417_), .Y(new_n12420_));
  XOR2X1   g12356(.A(new_n12420_), .B(new_n12400_), .Y(new_n12421_));
  OR2X1    g12357(.A(new_n12349_), .B(new_n12335_), .Y(new_n12422_));
  NAND2X1  g12358(.A(new_n12347_), .B(new_n12346_), .Y(new_n12423_));
  AND2X1   g12359(.A(new_n12423_), .B(new_n12422_), .Y(new_n12424_));
  XOR2X1   g12360(.A(new_n12424_), .B(new_n12421_), .Y(new_n12425_));
  AOI22X1  g12361(.A0(new_n12155_), .A1(new_n2424_), .B0(new_n12151_), .B1(new_n2418_), .Y(new_n12426_));
  OAI21X1  g12362(.A0(new_n12186_), .A1(new_n2626_), .B0(new_n12426_), .Y(new_n12427_));
  NAND2X1  g12363(.A(new_n12185_), .B(new_n12156_), .Y(new_n12428_));
  INVX1    g12364(.A(new_n12187_), .Y(new_n12429_));
  XOR2X1   g12365(.A(new_n12429_), .B(new_n12428_), .Y(new_n12430_));
  AOI21X1  g12366(.A0(new_n12430_), .A1(new_n2301_), .B0(new_n12427_), .Y(new_n12431_));
  XOR2X1   g12367(.A(new_n12431_), .B(\a[26] ), .Y(new_n12432_));
  XOR2X1   g12368(.A(new_n12432_), .B(new_n12425_), .Y(new_n12433_));
  XOR2X1   g12369(.A(new_n12433_), .B(new_n12393_), .Y(new_n12434_));
  XOR2X1   g12370(.A(new_n12434_), .B(new_n12318_), .Y(new_n12435_));
  INVX1    g12371(.A(new_n12435_), .Y(new_n12436_));
  INVX1    g12372(.A(new_n12351_), .Y(new_n12437_));
  XOR2X1   g12373(.A(new_n12391_), .B(new_n12437_), .Y(new_n12438_));
  OAI22X1  g12374(.A0(new_n12186_), .A1(new_n4016_), .B0(new_n12192_), .B1(new_n2743_), .Y(new_n12439_));
  AOI21X1  g12375(.A0(new_n12141_), .A1(new_n2745_), .B0(new_n12439_), .Y(new_n12440_));
  NAND2X1  g12376(.A(new_n12190_), .B(new_n12149_), .Y(new_n12441_));
  NOR2X1   g12377(.A(new_n12144_), .B(new_n12141_), .Y(new_n12442_));
  NOR3X1   g12378(.A(new_n12442_), .B(new_n12441_), .C(new_n12145_), .Y(new_n12443_));
  AOI21X1  g12379(.A0(new_n12193_), .A1(new_n12441_), .B0(new_n12443_), .Y(new_n12444_));
  OAI21X1  g12380(.A0(new_n12444_), .A1(new_n2692_), .B0(new_n12440_), .Y(new_n12445_));
  XOR2X1   g12381(.A(new_n12445_), .B(new_n70_), .Y(new_n12446_));
  NOR2X1   g12382(.A(new_n12446_), .B(new_n12438_), .Y(new_n12447_));
  XOR2X1   g12383(.A(new_n12389_), .B(new_n12362_), .Y(new_n12448_));
  INVX1    g12384(.A(new_n12448_), .Y(new_n12449_));
  OAI22X1  g12385(.A0(new_n12322_), .A1(new_n4016_), .B0(new_n12186_), .B1(new_n2743_), .Y(new_n12450_));
  AOI21X1  g12386(.A0(new_n12144_), .A1(new_n2745_), .B0(new_n12450_), .Y(new_n12451_));
  NOR2X1   g12387(.A(new_n12188_), .B(new_n12152_), .Y(new_n12452_));
  XOR2X1   g12388(.A(new_n12189_), .B(new_n12452_), .Y(new_n12453_));
  OAI21X1  g12389(.A0(new_n12453_), .A1(new_n2692_), .B0(new_n12451_), .Y(new_n12454_));
  XOR2X1   g12390(.A(new_n12454_), .B(new_n70_), .Y(new_n12455_));
  OR2X1    g12391(.A(new_n12455_), .B(new_n12449_), .Y(new_n12456_));
  AOI22X1  g12392(.A0(new_n12155_), .A1(new_n2657_), .B0(new_n12151_), .B1(new_n2696_), .Y(new_n12457_));
  OAI21X1  g12393(.A0(new_n12186_), .A1(new_n2753_), .B0(new_n12457_), .Y(new_n12458_));
  AOI21X1  g12394(.A0(new_n12430_), .A1(new_n2658_), .B0(new_n12458_), .Y(new_n12459_));
  XOR2X1   g12395(.A(new_n12459_), .B(\a[23] ), .Y(new_n12460_));
  INVX1    g12396(.A(new_n12460_), .Y(new_n12461_));
  XOR2X1   g12397(.A(new_n12388_), .B(new_n12387_), .Y(new_n12462_));
  XOR2X1   g12398(.A(new_n12462_), .B(new_n12460_), .Y(new_n12463_));
  XOR2X1   g12399(.A(new_n12386_), .B(new_n12381_), .Y(new_n12464_));
  AOI22X1  g12400(.A0(new_n12158_), .A1(new_n2657_), .B0(new_n12155_), .B1(new_n2696_), .Y(new_n12465_));
  OAI21X1  g12401(.A0(new_n12322_), .A1(new_n2753_), .B0(new_n12465_), .Y(new_n12466_));
  AOI21X1  g12402(.A0(new_n12321_), .A1(new_n2658_), .B0(new_n12466_), .Y(new_n12467_));
  XOR2X1   g12403(.A(new_n12467_), .B(\a[23] ), .Y(new_n12468_));
  NOR2X1   g12404(.A(new_n12468_), .B(new_n12464_), .Y(new_n12469_));
  AOI22X1  g12405(.A0(new_n12162_), .A1(new_n2657_), .B0(new_n12158_), .B1(new_n2696_), .Y(new_n12470_));
  OAI21X1  g12406(.A0(new_n12353_), .A1(new_n2753_), .B0(new_n12470_), .Y(new_n12471_));
  AOI21X1  g12407(.A0(new_n12352_), .A1(new_n2658_), .B0(new_n12471_), .Y(new_n12472_));
  XOR2X1   g12408(.A(new_n12472_), .B(\a[23] ), .Y(new_n12473_));
  INVX1    g12409(.A(new_n12473_), .Y(new_n12474_));
  NOR3X1   g12410(.A(new_n12375_), .B(new_n12372_), .C(new_n89_), .Y(new_n12475_));
  XOR2X1   g12411(.A(new_n12378_), .B(\a[26] ), .Y(new_n12476_));
  XOR2X1   g12412(.A(new_n12476_), .B(new_n12475_), .Y(new_n12477_));
  XOR2X1   g12413(.A(new_n12477_), .B(new_n12473_), .Y(new_n12478_));
  NOR2X1   g12414(.A(new_n12372_), .B(new_n89_), .Y(new_n12479_));
  XOR2X1   g12415(.A(new_n12375_), .B(new_n12479_), .Y(new_n12480_));
  OAI22X1  g12416(.A0(new_n12168_), .A1(new_n4016_), .B0(new_n12329_), .B1(new_n2743_), .Y(new_n12481_));
  AOI21X1  g12417(.A0(new_n12158_), .A1(new_n2745_), .B0(new_n12481_), .Y(new_n12482_));
  OAI21X1  g12418(.A0(new_n12368_), .A1(new_n2692_), .B0(new_n12482_), .Y(new_n12483_));
  XOR2X1   g12419(.A(new_n12483_), .B(new_n70_), .Y(new_n12484_));
  NOR2X1   g12420(.A(new_n12484_), .B(new_n12480_), .Y(new_n12485_));
  AOI21X1  g12421(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n2655_), .Y(new_n12486_));
  OAI22X1  g12422(.A0(new_n12176_), .A1(new_n2743_), .B0(new_n12170_), .B1(new_n2753_), .Y(new_n12487_));
  AOI21X1  g12423(.A0(new_n12337_), .A1(new_n2658_), .B0(new_n12487_), .Y(new_n12488_));
  XOR2X1   g12424(.A(new_n12488_), .B(\a[23] ), .Y(new_n12489_));
  OAI22X1  g12425(.A0(new_n12176_), .A1(new_n4016_), .B0(new_n12170_), .B1(new_n2743_), .Y(new_n12490_));
  AOI21X1  g12426(.A0(new_n12165_), .A1(new_n2745_), .B0(new_n12490_), .Y(new_n12491_));
  OAI21X1  g12427(.A0(new_n12344_), .A1(new_n2692_), .B0(new_n12491_), .Y(new_n12492_));
  NOR4X1   g12428(.A(new_n12492_), .B(new_n12489_), .C(new_n12486_), .D(new_n70_), .Y(new_n12493_));
  NAND2X1  g12429(.A(new_n12493_), .B(new_n12372_), .Y(new_n12494_));
  XOR2X1   g12430(.A(new_n12493_), .B(new_n12372_), .Y(new_n12495_));
  INVX1    g12431(.A(new_n12495_), .Y(new_n12496_));
  AOI22X1  g12432(.A0(new_n12331_), .A1(new_n2657_), .B0(new_n12165_), .B1(new_n2696_), .Y(new_n12497_));
  OAI21X1  g12433(.A0(new_n12329_), .A1(new_n2753_), .B0(new_n12497_), .Y(new_n12498_));
  AOI21X1  g12434(.A0(new_n12328_), .A1(new_n2658_), .B0(new_n12498_), .Y(new_n12499_));
  XOR2X1   g12435(.A(new_n12499_), .B(\a[23] ), .Y(new_n12500_));
  OAI21X1  g12436(.A0(new_n12500_), .A1(new_n12496_), .B0(new_n12494_), .Y(new_n12501_));
  XOR2X1   g12437(.A(new_n12484_), .B(new_n12480_), .Y(new_n12502_));
  AOI21X1  g12438(.A0(new_n12502_), .A1(new_n12501_), .B0(new_n12485_), .Y(new_n12503_));
  NOR2X1   g12439(.A(new_n12503_), .B(new_n12478_), .Y(new_n12504_));
  AOI21X1  g12440(.A0(new_n12477_), .A1(new_n12474_), .B0(new_n12504_), .Y(new_n12505_));
  INVX1    g12441(.A(new_n12505_), .Y(new_n12506_));
  XOR2X1   g12442(.A(new_n12468_), .B(new_n12464_), .Y(new_n12507_));
  AOI21X1  g12443(.A0(new_n12507_), .A1(new_n12506_), .B0(new_n12469_), .Y(new_n12508_));
  NOR2X1   g12444(.A(new_n12508_), .B(new_n12463_), .Y(new_n12509_));
  AOI21X1  g12445(.A0(new_n12462_), .A1(new_n12461_), .B0(new_n12509_), .Y(new_n12510_));
  XOR2X1   g12446(.A(new_n12455_), .B(new_n12448_), .Y(new_n12511_));
  OAI21X1  g12447(.A0(new_n12511_), .A1(new_n12510_), .B0(new_n12456_), .Y(new_n12512_));
  XOR2X1   g12448(.A(new_n12446_), .B(new_n12438_), .Y(new_n12513_));
  AOI21X1  g12449(.A0(new_n12513_), .A1(new_n12512_), .B0(new_n12447_), .Y(new_n12514_));
  XOR2X1   g12450(.A(new_n12514_), .B(new_n12436_), .Y(new_n12515_));
  INVX1    g12451(.A(new_n12113_), .Y(new_n12516_));
  OAI22X1  g12452(.A0(new_n12134_), .A1(new_n3250_), .B0(new_n12117_), .B1(new_n3144_), .Y(new_n12517_));
  AOI21X1  g12453(.A0(new_n12516_), .A1(new_n3146_), .B0(new_n12517_), .Y(new_n12518_));
  XOR2X1   g12454(.A(new_n12117_), .B(new_n12113_), .Y(new_n12519_));
  AOI21X1  g12455(.A0(new_n12201_), .A1(new_n12135_), .B0(new_n12519_), .Y(new_n12520_));
  NOR3X1   g12456(.A(new_n12203_), .B(new_n12202_), .C(new_n12118_), .Y(new_n12521_));
  NOR2X1   g12457(.A(new_n12521_), .B(new_n12520_), .Y(new_n12522_));
  OAI21X1  g12458(.A0(new_n12522_), .A1(new_n3098_), .B0(new_n12518_), .Y(new_n12523_));
  XOR2X1   g12459(.A(new_n12523_), .B(\a[20] ), .Y(new_n12524_));
  OR2X1    g12460(.A(new_n12199_), .B(new_n12139_), .Y(new_n12525_));
  XOR2X1   g12461(.A(new_n12200_), .B(new_n12525_), .Y(new_n12526_));
  AOI22X1  g12462(.A0(new_n12138_), .A1(new_n2875_), .B0(new_n12133_), .B1(new_n3099_), .Y(new_n12527_));
  OAI21X1  g12463(.A0(new_n12117_), .A1(new_n3152_), .B0(new_n12527_), .Y(new_n12528_));
  AOI21X1  g12464(.A0(new_n12526_), .A1(new_n2876_), .B0(new_n12528_), .Y(new_n12529_));
  XOR2X1   g12465(.A(new_n12529_), .B(\a[20] ), .Y(new_n12530_));
  INVX1    g12466(.A(new_n12530_), .Y(new_n12531_));
  XOR2X1   g12467(.A(new_n12513_), .B(new_n12512_), .Y(new_n12532_));
  AND2X1   g12468(.A(new_n12532_), .B(new_n12531_), .Y(new_n12533_));
  XOR2X1   g12469(.A(new_n12532_), .B(new_n12530_), .Y(new_n12534_));
  INVX1    g12470(.A(new_n12534_), .Y(new_n12535_));
  XOR2X1   g12471(.A(new_n12198_), .B(new_n12197_), .Y(new_n12536_));
  AOI22X1  g12472(.A0(new_n12141_), .A1(new_n2875_), .B0(new_n12138_), .B1(new_n3099_), .Y(new_n12537_));
  OAI21X1  g12473(.A0(new_n12134_), .A1(new_n3152_), .B0(new_n12537_), .Y(new_n12538_));
  AOI21X1  g12474(.A0(new_n12536_), .A1(new_n2876_), .B0(new_n12538_), .Y(new_n12539_));
  XOR2X1   g12475(.A(new_n12539_), .B(\a[20] ), .Y(new_n12540_));
  INVX1    g12476(.A(new_n12511_), .Y(new_n12541_));
  XOR2X1   g12477(.A(new_n12541_), .B(new_n12510_), .Y(new_n12542_));
  OR2X1    g12478(.A(new_n12542_), .B(new_n12540_), .Y(new_n12543_));
  XOR2X1   g12479(.A(new_n12542_), .B(new_n12540_), .Y(new_n12544_));
  INVX1    g12480(.A(new_n12544_), .Y(new_n12545_));
  INVX1    g12481(.A(new_n12463_), .Y(new_n12546_));
  XOR2X1   g12482(.A(new_n12508_), .B(new_n12546_), .Y(new_n12547_));
  AOI22X1  g12483(.A0(new_n12144_), .A1(new_n2875_), .B0(new_n12141_), .B1(new_n3099_), .Y(new_n12548_));
  OAI21X1  g12484(.A0(new_n12314_), .A1(new_n3152_), .B0(new_n12548_), .Y(new_n12549_));
  AOI21X1  g12485(.A0(new_n12313_), .A1(new_n2876_), .B0(new_n12549_), .Y(new_n12550_));
  XOR2X1   g12486(.A(new_n12550_), .B(\a[20] ), .Y(new_n12551_));
  NOR2X1   g12487(.A(new_n12551_), .B(new_n12547_), .Y(new_n12552_));
  XOR2X1   g12488(.A(new_n12507_), .B(new_n12506_), .Y(new_n12553_));
  INVX1    g12489(.A(new_n12553_), .Y(new_n12554_));
  OAI22X1  g12490(.A0(new_n12186_), .A1(new_n3250_), .B0(new_n12192_), .B1(new_n3144_), .Y(new_n12555_));
  AOI21X1  g12491(.A0(new_n12141_), .A1(new_n3146_), .B0(new_n12555_), .Y(new_n12556_));
  OAI21X1  g12492(.A0(new_n12444_), .A1(new_n3098_), .B0(new_n12556_), .Y(new_n12557_));
  XOR2X1   g12493(.A(new_n12557_), .B(new_n1920_), .Y(new_n12558_));
  OR2X1    g12494(.A(new_n12558_), .B(new_n12554_), .Y(new_n12559_));
  XOR2X1   g12495(.A(new_n12503_), .B(new_n12478_), .Y(new_n12560_));
  INVX1    g12496(.A(new_n12560_), .Y(new_n12561_));
  OAI22X1  g12497(.A0(new_n12322_), .A1(new_n3250_), .B0(new_n12186_), .B1(new_n3144_), .Y(new_n12562_));
  AOI21X1  g12498(.A0(new_n12144_), .A1(new_n3146_), .B0(new_n12562_), .Y(new_n12563_));
  OAI21X1  g12499(.A0(new_n12453_), .A1(new_n3098_), .B0(new_n12563_), .Y(new_n12564_));
  XOR2X1   g12500(.A(new_n12564_), .B(new_n1920_), .Y(new_n12565_));
  NOR2X1   g12501(.A(new_n12565_), .B(new_n12561_), .Y(new_n12566_));
  AOI22X1  g12502(.A0(new_n12155_), .A1(new_n2875_), .B0(new_n12151_), .B1(new_n3099_), .Y(new_n12567_));
  OAI21X1  g12503(.A0(new_n12186_), .A1(new_n3152_), .B0(new_n12567_), .Y(new_n12568_));
  AOI21X1  g12504(.A0(new_n12430_), .A1(new_n2876_), .B0(new_n12568_), .Y(new_n12569_));
  XOR2X1   g12505(.A(new_n12569_), .B(\a[20] ), .Y(new_n12570_));
  INVX1    g12506(.A(new_n12570_), .Y(new_n12571_));
  XOR2X1   g12507(.A(new_n12502_), .B(new_n12501_), .Y(new_n12572_));
  NAND2X1  g12508(.A(new_n12572_), .B(new_n12571_), .Y(new_n12573_));
  XOR2X1   g12509(.A(new_n12572_), .B(new_n12570_), .Y(new_n12574_));
  XOR2X1   g12510(.A(new_n12500_), .B(new_n12495_), .Y(new_n12575_));
  AOI22X1  g12511(.A0(new_n12158_), .A1(new_n2875_), .B0(new_n12155_), .B1(new_n3099_), .Y(new_n12576_));
  OAI21X1  g12512(.A0(new_n12322_), .A1(new_n3152_), .B0(new_n12576_), .Y(new_n12577_));
  AOI21X1  g12513(.A0(new_n12321_), .A1(new_n2876_), .B0(new_n12577_), .Y(new_n12578_));
  XOR2X1   g12514(.A(new_n12578_), .B(\a[20] ), .Y(new_n12579_));
  NOR2X1   g12515(.A(new_n12579_), .B(new_n12575_), .Y(new_n12580_));
  AOI22X1  g12516(.A0(new_n12162_), .A1(new_n2875_), .B0(new_n12158_), .B1(new_n3099_), .Y(new_n12581_));
  OAI21X1  g12517(.A0(new_n12353_), .A1(new_n3152_), .B0(new_n12581_), .Y(new_n12582_));
  AOI21X1  g12518(.A0(new_n12352_), .A1(new_n2876_), .B0(new_n12582_), .Y(new_n12583_));
  XOR2X1   g12519(.A(new_n12583_), .B(\a[20] ), .Y(new_n12584_));
  NOR3X1   g12520(.A(new_n12489_), .B(new_n12486_), .C(new_n70_), .Y(new_n12585_));
  XOR2X1   g12521(.A(new_n12492_), .B(\a[23] ), .Y(new_n12586_));
  NOR2X1   g12522(.A(new_n12586_), .B(new_n12585_), .Y(new_n12587_));
  NOR3X1   g12523(.A(new_n12587_), .B(new_n12584_), .C(new_n12493_), .Y(new_n12588_));
  XOR2X1   g12524(.A(new_n12586_), .B(new_n12585_), .Y(new_n12589_));
  XOR2X1   g12525(.A(new_n12589_), .B(new_n12584_), .Y(new_n12590_));
  NOR2X1   g12526(.A(new_n12486_), .B(new_n70_), .Y(new_n12591_));
  XOR2X1   g12527(.A(new_n12489_), .B(new_n12591_), .Y(new_n12592_));
  OAI22X1  g12528(.A0(new_n12168_), .A1(new_n3250_), .B0(new_n12329_), .B1(new_n3144_), .Y(new_n12593_));
  AOI21X1  g12529(.A0(new_n12158_), .A1(new_n3146_), .B0(new_n12593_), .Y(new_n12594_));
  OAI21X1  g12530(.A0(new_n12368_), .A1(new_n3098_), .B0(new_n12594_), .Y(new_n12595_));
  XOR2X1   g12531(.A(new_n12595_), .B(new_n1920_), .Y(new_n12596_));
  NOR2X1   g12532(.A(new_n12596_), .B(new_n12592_), .Y(new_n12597_));
  OAI22X1  g12533(.A0(new_n12176_), .A1(new_n3144_), .B0(new_n12170_), .B1(new_n3152_), .Y(new_n12598_));
  AOI21X1  g12534(.A0(new_n12337_), .A1(new_n2876_), .B0(new_n12598_), .Y(new_n12599_));
  XOR2X1   g12535(.A(new_n12599_), .B(\a[20] ), .Y(new_n12600_));
  AOI21X1  g12536(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n2869_), .Y(new_n12601_));
  OAI22X1  g12537(.A0(new_n12176_), .A1(new_n3250_), .B0(new_n12170_), .B1(new_n3144_), .Y(new_n12602_));
  AOI21X1  g12538(.A0(new_n12165_), .A1(new_n3146_), .B0(new_n12602_), .Y(new_n12603_));
  OAI21X1  g12539(.A0(new_n12344_), .A1(new_n3098_), .B0(new_n12603_), .Y(new_n12604_));
  NOR4X1   g12540(.A(new_n12604_), .B(new_n12601_), .C(new_n12600_), .D(new_n1920_), .Y(new_n12605_));
  NAND2X1  g12541(.A(new_n12605_), .B(new_n12486_), .Y(new_n12606_));
  INVX1    g12542(.A(new_n12605_), .Y(new_n12607_));
  XOR2X1   g12543(.A(new_n12607_), .B(new_n12486_), .Y(new_n12608_));
  AOI22X1  g12544(.A0(new_n12331_), .A1(new_n2875_), .B0(new_n12165_), .B1(new_n3099_), .Y(new_n12609_));
  OAI21X1  g12545(.A0(new_n12329_), .A1(new_n3152_), .B0(new_n12609_), .Y(new_n12610_));
  AOI21X1  g12546(.A0(new_n12328_), .A1(new_n2876_), .B0(new_n12610_), .Y(new_n12611_));
  XOR2X1   g12547(.A(new_n12611_), .B(\a[20] ), .Y(new_n12612_));
  OAI21X1  g12548(.A0(new_n12612_), .A1(new_n12608_), .B0(new_n12606_), .Y(new_n12613_));
  XOR2X1   g12549(.A(new_n12596_), .B(new_n12592_), .Y(new_n12614_));
  AOI21X1  g12550(.A0(new_n12614_), .A1(new_n12613_), .B0(new_n12597_), .Y(new_n12615_));
  NOR2X1   g12551(.A(new_n12615_), .B(new_n12590_), .Y(new_n12616_));
  OR2X1    g12552(.A(new_n12616_), .B(new_n12588_), .Y(new_n12617_));
  XOR2X1   g12553(.A(new_n12579_), .B(new_n12575_), .Y(new_n12618_));
  AOI21X1  g12554(.A0(new_n12618_), .A1(new_n12617_), .B0(new_n12580_), .Y(new_n12619_));
  OR2X1    g12555(.A(new_n12619_), .B(new_n12574_), .Y(new_n12620_));
  XOR2X1   g12556(.A(new_n12565_), .B(new_n12560_), .Y(new_n12621_));
  AOI21X1  g12557(.A0(new_n12620_), .A1(new_n12573_), .B0(new_n12621_), .Y(new_n12622_));
  NOR2X1   g12558(.A(new_n12622_), .B(new_n12566_), .Y(new_n12623_));
  XOR2X1   g12559(.A(new_n12558_), .B(new_n12553_), .Y(new_n12624_));
  OAI21X1  g12560(.A0(new_n12624_), .A1(new_n12623_), .B0(new_n12559_), .Y(new_n12625_));
  XOR2X1   g12561(.A(new_n12551_), .B(new_n12547_), .Y(new_n12626_));
  AOI21X1  g12562(.A0(new_n12626_), .A1(new_n12625_), .B0(new_n12552_), .Y(new_n12627_));
  OAI21X1  g12563(.A0(new_n12627_), .A1(new_n12545_), .B0(new_n12543_), .Y(new_n12628_));
  AOI21X1  g12564(.A0(new_n12628_), .A1(new_n12535_), .B0(new_n12533_), .Y(new_n12629_));
  XOR2X1   g12565(.A(new_n12523_), .B(new_n1920_), .Y(new_n12630_));
  XOR2X1   g12566(.A(new_n12630_), .B(new_n12515_), .Y(new_n12631_));
  NOR2X1   g12567(.A(new_n12631_), .B(new_n12629_), .Y(new_n12632_));
  AOI21X1  g12568(.A0(new_n12524_), .A1(new_n12515_), .B0(new_n12632_), .Y(new_n12633_));
  AOI22X1  g12569(.A0(new_n12141_), .A1(new_n2657_), .B0(new_n12138_), .B1(new_n2696_), .Y(new_n12634_));
  OAI21X1  g12570(.A0(new_n12134_), .A1(new_n2753_), .B0(new_n12634_), .Y(new_n12635_));
  AOI21X1  g12571(.A0(new_n12536_), .A1(new_n2658_), .B0(new_n12635_), .Y(new_n12636_));
  XOR2X1   g12572(.A(new_n12636_), .B(\a[23] ), .Y(new_n12637_));
  NOR2X1   g12573(.A(new_n12432_), .B(new_n12425_), .Y(new_n12638_));
  INVX1    g12574(.A(new_n12638_), .Y(new_n12639_));
  INVX1    g12575(.A(new_n12433_), .Y(new_n12640_));
  OAI21X1  g12576(.A0(new_n12640_), .A1(new_n12393_), .B0(new_n12639_), .Y(new_n12641_));
  AOI22X1  g12577(.A0(new_n12162_), .A1(new_n2185_), .B0(new_n12158_), .B1(new_n2095_), .Y(new_n12642_));
  OAI21X1  g12578(.A0(new_n12353_), .A1(new_n2140_), .B0(new_n12642_), .Y(new_n12643_));
  AOI21X1  g12579(.A0(new_n12352_), .A1(new_n2062_), .B0(new_n12643_), .Y(new_n12644_));
  XOR2X1   g12580(.A(new_n12644_), .B(\a[29] ), .Y(new_n12645_));
  OAI22X1  g12581(.A0(new_n12176_), .A1(new_n2245_), .B0(new_n12170_), .B1(new_n1885_), .Y(new_n12646_));
  AOI21X1  g12582(.A0(new_n12165_), .A1(new_n1889_), .B0(new_n12646_), .Y(new_n12647_));
  OAI21X1  g12583(.A0(new_n12344_), .A1(new_n3178_), .B0(new_n12647_), .Y(new_n12648_));
  INVX1    g12584(.A(new_n12648_), .Y(new_n12649_));
  OR2X1    g12585(.A(new_n12419_), .B(new_n12416_), .Y(new_n12650_));
  INVX1    g12586(.A(new_n3742_), .Y(new_n12651_));
  OR4X1    g12587(.A(new_n7425_), .B(new_n1910_), .C(new_n888_), .D(new_n700_), .Y(new_n12652_));
  OR2X1    g12588(.A(new_n6768_), .B(new_n2015_), .Y(new_n12653_));
  OR4X1    g12589(.A(new_n479_), .B(new_n536_), .C(new_n522_), .D(new_n160_), .Y(new_n12654_));
  OR4X1    g12590(.A(new_n293_), .B(new_n239_), .C(new_n218_), .D(new_n202_), .Y(new_n12655_));
  OAI22X1  g12591(.A0(new_n143_), .A1(new_n79_), .B0(new_n108_), .B1(new_n96_), .Y(new_n12656_));
  OR2X1    g12592(.A(new_n12656_), .B(new_n370_), .Y(new_n12657_));
  OR4X1    g12593(.A(new_n740_), .B(new_n383_), .C(new_n350_), .D(new_n203_), .Y(new_n12658_));
  OR4X1    g12594(.A(new_n12658_), .B(new_n12657_), .C(new_n12655_), .D(new_n12654_), .Y(new_n12659_));
  OR4X1    g12595(.A(new_n12659_), .B(new_n12653_), .C(new_n12652_), .D(new_n402_), .Y(new_n12660_));
  NOR3X1   g12596(.A(new_n12660_), .B(new_n12401_), .C(new_n12651_), .Y(new_n12661_));
  XOR2X1   g12597(.A(new_n12661_), .B(new_n12650_), .Y(new_n12662_));
  XOR2X1   g12598(.A(new_n12662_), .B(new_n12649_), .Y(new_n12663_));
  XOR2X1   g12599(.A(new_n12663_), .B(new_n12645_), .Y(new_n12664_));
  INVX1    g12600(.A(new_n12664_), .Y(new_n12665_));
  NOR2X1   g12601(.A(new_n12420_), .B(new_n12400_), .Y(new_n12666_));
  INVX1    g12602(.A(new_n12424_), .Y(new_n12667_));
  AOI21X1  g12603(.A0(new_n12667_), .A1(new_n12421_), .B0(new_n12666_), .Y(new_n12668_));
  XOR2X1   g12604(.A(new_n12668_), .B(new_n12665_), .Y(new_n12669_));
  OAI22X1  g12605(.A0(new_n12322_), .A1(new_n2666_), .B0(new_n12186_), .B1(new_n2419_), .Y(new_n12670_));
  AOI21X1  g12606(.A0(new_n12144_), .A1(new_n2423_), .B0(new_n12670_), .Y(new_n12671_));
  OAI21X1  g12607(.A0(new_n12453_), .A1(new_n2665_), .B0(new_n12671_), .Y(new_n12672_));
  XOR2X1   g12608(.A(new_n12672_), .B(new_n89_), .Y(new_n12673_));
  XOR2X1   g12609(.A(new_n12673_), .B(new_n12669_), .Y(new_n12674_));
  XOR2X1   g12610(.A(new_n12674_), .B(new_n12641_), .Y(new_n12675_));
  XOR2X1   g12611(.A(new_n12675_), .B(new_n12637_), .Y(new_n12676_));
  OR2X1    g12612(.A(new_n12434_), .B(new_n12318_), .Y(new_n12677_));
  OAI21X1  g12613(.A0(new_n12514_), .A1(new_n12436_), .B0(new_n12677_), .Y(new_n12678_));
  XOR2X1   g12614(.A(new_n12678_), .B(new_n12676_), .Y(new_n12679_));
  OAI22X1  g12615(.A0(new_n12117_), .A1(new_n3250_), .B0(new_n12113_), .B1(new_n3144_), .Y(new_n12680_));
  AOI21X1  g12616(.A0(new_n12208_), .A1(new_n3146_), .B0(new_n12680_), .Y(new_n12681_));
  INVX1    g12617(.A(new_n12206_), .Y(new_n12682_));
  INVX1    g12618(.A(new_n12207_), .Y(new_n12683_));
  AOI21X1  g12619(.A0(new_n12682_), .A1(new_n12115_), .B0(new_n12205_), .Y(new_n12684_));
  AOI21X1  g12620(.A0(new_n12683_), .A1(new_n12682_), .B0(new_n12684_), .Y(new_n12685_));
  OAI21X1  g12621(.A0(new_n12685_), .A1(new_n3098_), .B0(new_n12681_), .Y(new_n12686_));
  XOR2X1   g12622(.A(new_n12686_), .B(new_n1920_), .Y(new_n12687_));
  XOR2X1   g12623(.A(new_n12687_), .B(new_n12679_), .Y(new_n12688_));
  INVX1    g12624(.A(new_n12688_), .Y(new_n12689_));
  XOR2X1   g12625(.A(new_n12689_), .B(new_n12633_), .Y(new_n12690_));
  XOR2X1   g12626(.A(new_n12690_), .B(new_n12310_), .Y(new_n12691_));
  XOR2X1   g12627(.A(new_n12109_), .B(new_n12104_), .Y(new_n12692_));
  AOI22X1  g12628(.A0(new_n12214_), .A1(new_n12213_), .B0(new_n12692_), .B1(new_n12211_), .Y(new_n12693_));
  INVX1    g12629(.A(new_n12693_), .Y(new_n12694_));
  INVX1    g12630(.A(new_n12104_), .Y(new_n12695_));
  AOI22X1  g12631(.A0(new_n12208_), .A1(new_n3232_), .B0(new_n12107_), .B1(new_n3390_), .Y(new_n12696_));
  OAI21X1  g12632(.A0(new_n12695_), .A1(new_n3545_), .B0(new_n12696_), .Y(new_n12697_));
  AOI21X1  g12633(.A0(new_n12694_), .A1(new_n3234_), .B0(new_n12697_), .Y(new_n12698_));
  XOR2X1   g12634(.A(new_n12698_), .B(\a[17] ), .Y(new_n12699_));
  INVX1    g12635(.A(new_n12631_), .Y(new_n12700_));
  XOR2X1   g12636(.A(new_n12700_), .B(new_n12629_), .Y(new_n12701_));
  OR2X1    g12637(.A(new_n12701_), .B(new_n12699_), .Y(new_n12702_));
  XOR2X1   g12638(.A(new_n12701_), .B(new_n12699_), .Y(new_n12703_));
  INVX1    g12639(.A(new_n12703_), .Y(new_n12704_));
  XOR2X1   g12640(.A(new_n12628_), .B(new_n12534_), .Y(new_n12705_));
  OAI22X1  g12641(.A0(new_n12113_), .A1(new_n3231_), .B0(new_n12111_), .B1(new_n3389_), .Y(new_n12706_));
  AOI21X1  g12642(.A0(new_n12107_), .A1(new_n3546_), .B0(new_n12706_), .Y(new_n12707_));
  XOR2X1   g12643(.A(new_n12209_), .B(new_n12683_), .Y(new_n12708_));
  OAI21X1  g12644(.A0(new_n12708_), .A1(new_n3388_), .B0(new_n12707_), .Y(new_n12709_));
  XOR2X1   g12645(.A(new_n12709_), .B(new_n2445_), .Y(new_n12710_));
  NOR2X1   g12646(.A(new_n12710_), .B(new_n12705_), .Y(new_n12711_));
  XOR2X1   g12647(.A(new_n12627_), .B(new_n12545_), .Y(new_n12712_));
  INVX1    g12648(.A(new_n12712_), .Y(new_n12713_));
  OAI22X1  g12649(.A0(new_n12117_), .A1(new_n3231_), .B0(new_n12113_), .B1(new_n3389_), .Y(new_n12714_));
  AOI21X1  g12650(.A0(new_n12208_), .A1(new_n3546_), .B0(new_n12714_), .Y(new_n12715_));
  OAI21X1  g12651(.A0(new_n12685_), .A1(new_n3388_), .B0(new_n12715_), .Y(new_n12716_));
  XOR2X1   g12652(.A(new_n12716_), .B(new_n2445_), .Y(new_n12717_));
  OR2X1    g12653(.A(new_n12717_), .B(new_n12713_), .Y(new_n12718_));
  INVX1    g12654(.A(new_n12522_), .Y(new_n12719_));
  INVX1    g12655(.A(new_n12117_), .Y(new_n12720_));
  AOI22X1  g12656(.A0(new_n12133_), .A1(new_n3232_), .B0(new_n12720_), .B1(new_n3390_), .Y(new_n12721_));
  OAI21X1  g12657(.A0(new_n12113_), .A1(new_n3545_), .B0(new_n12721_), .Y(new_n12722_));
  AOI21X1  g12658(.A0(new_n12719_), .A1(new_n3234_), .B0(new_n12722_), .Y(new_n12723_));
  XOR2X1   g12659(.A(new_n12723_), .B(\a[17] ), .Y(new_n12724_));
  INVX1    g12660(.A(new_n12724_), .Y(new_n12725_));
  XOR2X1   g12661(.A(new_n12626_), .B(new_n12625_), .Y(new_n12726_));
  XOR2X1   g12662(.A(new_n12726_), .B(new_n12724_), .Y(new_n12727_));
  AOI22X1  g12663(.A0(new_n12138_), .A1(new_n3232_), .B0(new_n12133_), .B1(new_n3390_), .Y(new_n12728_));
  OAI21X1  g12664(.A0(new_n12117_), .A1(new_n3545_), .B0(new_n12728_), .Y(new_n12729_));
  AOI21X1  g12665(.A0(new_n12526_), .A1(new_n3234_), .B0(new_n12729_), .Y(new_n12730_));
  XOR2X1   g12666(.A(new_n12730_), .B(\a[17] ), .Y(new_n12731_));
  INVX1    g12667(.A(new_n12624_), .Y(new_n12732_));
  XOR2X1   g12668(.A(new_n12732_), .B(new_n12623_), .Y(new_n12733_));
  NOR2X1   g12669(.A(new_n12733_), .B(new_n12731_), .Y(new_n12734_));
  XOR2X1   g12670(.A(new_n12733_), .B(new_n12731_), .Y(new_n12735_));
  AOI22X1  g12671(.A0(new_n12141_), .A1(new_n3232_), .B0(new_n12138_), .B1(new_n3390_), .Y(new_n12736_));
  OAI21X1  g12672(.A0(new_n12134_), .A1(new_n3545_), .B0(new_n12736_), .Y(new_n12737_));
  AOI21X1  g12673(.A0(new_n12536_), .A1(new_n3234_), .B0(new_n12737_), .Y(new_n12738_));
  XOR2X1   g12674(.A(new_n12738_), .B(\a[17] ), .Y(new_n12739_));
  AND2X1   g12675(.A(new_n12620_), .B(new_n12573_), .Y(new_n12740_));
  INVX1    g12676(.A(new_n12621_), .Y(new_n12741_));
  XOR2X1   g12677(.A(new_n12741_), .B(new_n12740_), .Y(new_n12742_));
  OR2X1    g12678(.A(new_n12742_), .B(new_n12739_), .Y(new_n12743_));
  XOR2X1   g12679(.A(new_n12742_), .B(new_n12739_), .Y(new_n12744_));
  INVX1    g12680(.A(new_n12744_), .Y(new_n12745_));
  INVX1    g12681(.A(new_n12574_), .Y(new_n12746_));
  XOR2X1   g12682(.A(new_n12619_), .B(new_n12746_), .Y(new_n12747_));
  AOI22X1  g12683(.A0(new_n12144_), .A1(new_n3232_), .B0(new_n12141_), .B1(new_n3390_), .Y(new_n12748_));
  OAI21X1  g12684(.A0(new_n12314_), .A1(new_n3545_), .B0(new_n12748_), .Y(new_n12749_));
  AOI21X1  g12685(.A0(new_n12313_), .A1(new_n3234_), .B0(new_n12749_), .Y(new_n12750_));
  XOR2X1   g12686(.A(new_n12750_), .B(\a[17] ), .Y(new_n12751_));
  NOR2X1   g12687(.A(new_n12751_), .B(new_n12747_), .Y(new_n12752_));
  XOR2X1   g12688(.A(new_n12618_), .B(new_n12617_), .Y(new_n12753_));
  INVX1    g12689(.A(new_n12753_), .Y(new_n12754_));
  OAI22X1  g12690(.A0(new_n12186_), .A1(new_n3231_), .B0(new_n12192_), .B1(new_n3389_), .Y(new_n12755_));
  AOI21X1  g12691(.A0(new_n12141_), .A1(new_n3546_), .B0(new_n12755_), .Y(new_n12756_));
  OAI21X1  g12692(.A0(new_n12444_), .A1(new_n3388_), .B0(new_n12756_), .Y(new_n12757_));
  XOR2X1   g12693(.A(new_n12757_), .B(new_n2445_), .Y(new_n12758_));
  OR2X1    g12694(.A(new_n12758_), .B(new_n12754_), .Y(new_n12759_));
  XOR2X1   g12695(.A(new_n12615_), .B(new_n12590_), .Y(new_n12760_));
  INVX1    g12696(.A(new_n12760_), .Y(new_n12761_));
  OAI22X1  g12697(.A0(new_n12322_), .A1(new_n3231_), .B0(new_n12186_), .B1(new_n3389_), .Y(new_n12762_));
  AOI21X1  g12698(.A0(new_n12144_), .A1(new_n3546_), .B0(new_n12762_), .Y(new_n12763_));
  OAI21X1  g12699(.A0(new_n12453_), .A1(new_n3388_), .B0(new_n12763_), .Y(new_n12764_));
  XOR2X1   g12700(.A(new_n12764_), .B(new_n2445_), .Y(new_n12765_));
  NOR2X1   g12701(.A(new_n12765_), .B(new_n12761_), .Y(new_n12766_));
  AOI22X1  g12702(.A0(new_n12155_), .A1(new_n3232_), .B0(new_n12151_), .B1(new_n3390_), .Y(new_n12767_));
  OAI21X1  g12703(.A0(new_n12186_), .A1(new_n3545_), .B0(new_n12767_), .Y(new_n12768_));
  AOI21X1  g12704(.A0(new_n12430_), .A1(new_n3234_), .B0(new_n12768_), .Y(new_n12769_));
  XOR2X1   g12705(.A(new_n12769_), .B(\a[17] ), .Y(new_n12770_));
  INVX1    g12706(.A(new_n12770_), .Y(new_n12771_));
  XOR2X1   g12707(.A(new_n12614_), .B(new_n12613_), .Y(new_n12772_));
  NAND2X1  g12708(.A(new_n12772_), .B(new_n12771_), .Y(new_n12773_));
  XOR2X1   g12709(.A(new_n12772_), .B(new_n12770_), .Y(new_n12774_));
  XOR2X1   g12710(.A(new_n12611_), .B(new_n1920_), .Y(new_n12775_));
  XOR2X1   g12711(.A(new_n12775_), .B(new_n12608_), .Y(new_n12776_));
  AOI22X1  g12712(.A0(new_n12158_), .A1(new_n3232_), .B0(new_n12155_), .B1(new_n3390_), .Y(new_n12777_));
  OAI21X1  g12713(.A0(new_n12322_), .A1(new_n3545_), .B0(new_n12777_), .Y(new_n12778_));
  AOI21X1  g12714(.A0(new_n12321_), .A1(new_n3234_), .B0(new_n12778_), .Y(new_n12779_));
  XOR2X1   g12715(.A(new_n12779_), .B(\a[17] ), .Y(new_n12780_));
  NOR2X1   g12716(.A(new_n12780_), .B(new_n12776_), .Y(new_n12781_));
  AOI22X1  g12717(.A0(new_n12162_), .A1(new_n3232_), .B0(new_n12158_), .B1(new_n3390_), .Y(new_n12782_));
  OAI21X1  g12718(.A0(new_n12353_), .A1(new_n3545_), .B0(new_n12782_), .Y(new_n12783_));
  AOI21X1  g12719(.A0(new_n12352_), .A1(new_n3234_), .B0(new_n12783_), .Y(new_n12784_));
  XOR2X1   g12720(.A(new_n12784_), .B(\a[17] ), .Y(new_n12785_));
  NOR3X1   g12721(.A(new_n12601_), .B(new_n12600_), .C(new_n1920_), .Y(new_n12786_));
  XOR2X1   g12722(.A(new_n12604_), .B(\a[20] ), .Y(new_n12787_));
  NOR2X1   g12723(.A(new_n12787_), .B(new_n12786_), .Y(new_n12788_));
  NOR3X1   g12724(.A(new_n12788_), .B(new_n12785_), .C(new_n12605_), .Y(new_n12789_));
  XOR2X1   g12725(.A(new_n12787_), .B(new_n12786_), .Y(new_n12790_));
  XOR2X1   g12726(.A(new_n12790_), .B(new_n12785_), .Y(new_n12791_));
  NOR2X1   g12727(.A(new_n12601_), .B(new_n1920_), .Y(new_n12792_));
  XOR2X1   g12728(.A(new_n12792_), .B(new_n12600_), .Y(new_n12793_));
  OAI22X1  g12729(.A0(new_n12168_), .A1(new_n3231_), .B0(new_n12329_), .B1(new_n3389_), .Y(new_n12794_));
  AOI21X1  g12730(.A0(new_n12158_), .A1(new_n3546_), .B0(new_n12794_), .Y(new_n12795_));
  OAI21X1  g12731(.A0(new_n12368_), .A1(new_n3388_), .B0(new_n12795_), .Y(new_n12796_));
  XOR2X1   g12732(.A(new_n12796_), .B(new_n2445_), .Y(new_n12797_));
  NOR2X1   g12733(.A(new_n12797_), .B(new_n12793_), .Y(new_n12798_));
  OAI22X1  g12734(.A0(new_n12176_), .A1(new_n3389_), .B0(new_n12170_), .B1(new_n3545_), .Y(new_n12799_));
  AOI21X1  g12735(.A0(new_n12337_), .A1(new_n3234_), .B0(new_n12799_), .Y(new_n12800_));
  XOR2X1   g12736(.A(new_n12800_), .B(\a[17] ), .Y(new_n12801_));
  AOI21X1  g12737(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n3230_), .Y(new_n12802_));
  OAI22X1  g12738(.A0(new_n12176_), .A1(new_n3231_), .B0(new_n12170_), .B1(new_n3389_), .Y(new_n12803_));
  AOI21X1  g12739(.A0(new_n12165_), .A1(new_n3546_), .B0(new_n12803_), .Y(new_n12804_));
  OAI21X1  g12740(.A0(new_n12344_), .A1(new_n3388_), .B0(new_n12804_), .Y(new_n12805_));
  NOR4X1   g12741(.A(new_n12805_), .B(new_n12802_), .C(new_n12801_), .D(new_n2445_), .Y(new_n12806_));
  NAND2X1  g12742(.A(new_n12806_), .B(new_n12601_), .Y(new_n12807_));
  INVX1    g12743(.A(new_n12806_), .Y(new_n12808_));
  XOR2X1   g12744(.A(new_n12808_), .B(new_n12601_), .Y(new_n12809_));
  AOI22X1  g12745(.A0(new_n12331_), .A1(new_n3232_), .B0(new_n12165_), .B1(new_n3390_), .Y(new_n12810_));
  OAI21X1  g12746(.A0(new_n12329_), .A1(new_n3545_), .B0(new_n12810_), .Y(new_n12811_));
  AOI21X1  g12747(.A0(new_n12328_), .A1(new_n3234_), .B0(new_n12811_), .Y(new_n12812_));
  XOR2X1   g12748(.A(new_n12812_), .B(\a[17] ), .Y(new_n12813_));
  OAI21X1  g12749(.A0(new_n12813_), .A1(new_n12809_), .B0(new_n12807_), .Y(new_n12814_));
  XOR2X1   g12750(.A(new_n12797_), .B(new_n12793_), .Y(new_n12815_));
  AOI21X1  g12751(.A0(new_n12815_), .A1(new_n12814_), .B0(new_n12798_), .Y(new_n12816_));
  NOR2X1   g12752(.A(new_n12816_), .B(new_n12791_), .Y(new_n12817_));
  OR2X1    g12753(.A(new_n12817_), .B(new_n12789_), .Y(new_n12818_));
  XOR2X1   g12754(.A(new_n12780_), .B(new_n12776_), .Y(new_n12819_));
  AOI21X1  g12755(.A0(new_n12819_), .A1(new_n12818_), .B0(new_n12781_), .Y(new_n12820_));
  OR2X1    g12756(.A(new_n12820_), .B(new_n12774_), .Y(new_n12821_));
  XOR2X1   g12757(.A(new_n12765_), .B(new_n12760_), .Y(new_n12822_));
  AOI21X1  g12758(.A0(new_n12821_), .A1(new_n12773_), .B0(new_n12822_), .Y(new_n12823_));
  NOR2X1   g12759(.A(new_n12823_), .B(new_n12766_), .Y(new_n12824_));
  XOR2X1   g12760(.A(new_n12758_), .B(new_n12753_), .Y(new_n12825_));
  OAI21X1  g12761(.A0(new_n12825_), .A1(new_n12824_), .B0(new_n12759_), .Y(new_n12826_));
  XOR2X1   g12762(.A(new_n12751_), .B(new_n12747_), .Y(new_n12827_));
  AOI21X1  g12763(.A0(new_n12827_), .A1(new_n12826_), .B0(new_n12752_), .Y(new_n12828_));
  OAI21X1  g12764(.A0(new_n12828_), .A1(new_n12745_), .B0(new_n12743_), .Y(new_n12829_));
  AOI21X1  g12765(.A0(new_n12829_), .A1(new_n12735_), .B0(new_n12734_), .Y(new_n12830_));
  NOR2X1   g12766(.A(new_n12830_), .B(new_n12727_), .Y(new_n12831_));
  AOI21X1  g12767(.A0(new_n12726_), .A1(new_n12725_), .B0(new_n12831_), .Y(new_n12832_));
  XOR2X1   g12768(.A(new_n12717_), .B(new_n12712_), .Y(new_n12833_));
  OAI21X1  g12769(.A0(new_n12833_), .A1(new_n12832_), .B0(new_n12718_), .Y(new_n12834_));
  XOR2X1   g12770(.A(new_n12710_), .B(new_n12705_), .Y(new_n12835_));
  AOI21X1  g12771(.A0(new_n12835_), .A1(new_n12834_), .B0(new_n12711_), .Y(new_n12836_));
  OAI21X1  g12772(.A0(new_n12836_), .A1(new_n12704_), .B0(new_n12702_), .Y(new_n12837_));
  XOR2X1   g12773(.A(new_n12837_), .B(new_n12691_), .Y(new_n12838_));
  INVX1    g12774(.A(new_n12097_), .Y(new_n12839_));
  INVX1    g12775(.A(new_n12099_), .Y(new_n12840_));
  OAI22X1  g12776(.A0(new_n12840_), .A1(new_n3627_), .B0(new_n12839_), .B1(new_n3907_), .Y(new_n12841_));
  AOI21X1  g12777(.A0(new_n12095_), .A1(new_n3984_), .B0(new_n12841_), .Y(new_n12842_));
  XOR2X1   g12778(.A(new_n12097_), .B(new_n12095_), .Y(new_n12843_));
  INVX1    g12779(.A(new_n12843_), .Y(new_n12844_));
  AND2X1   g12780(.A(new_n12844_), .B(new_n12220_), .Y(new_n12845_));
  AOI21X1  g12781(.A0(new_n12222_), .A1(new_n12221_), .B0(new_n12845_), .Y(new_n12846_));
  OAI21X1  g12782(.A0(new_n12846_), .A1(new_n3906_), .B0(new_n12842_), .Y(new_n12847_));
  XOR2X1   g12783(.A(new_n12847_), .B(\a[14] ), .Y(new_n12848_));
  AND2X1   g12784(.A(new_n12848_), .B(new_n12838_), .Y(new_n12849_));
  XOR2X1   g12785(.A(new_n12836_), .B(new_n12704_), .Y(new_n12850_));
  OAI22X1  g12786(.A0(new_n12306_), .A1(new_n3627_), .B0(new_n12840_), .B1(new_n3907_), .Y(new_n12851_));
  AOI21X1  g12787(.A0(new_n12097_), .A1(new_n3984_), .B0(new_n12851_), .Y(new_n12852_));
  XOR2X1   g12788(.A(new_n12099_), .B(new_n12097_), .Y(new_n12853_));
  OR2X1    g12789(.A(new_n12853_), .B(new_n12218_), .Y(new_n12854_));
  OAI21X1  g12790(.A0(new_n12220_), .A1(new_n12219_), .B0(new_n12854_), .Y(new_n12855_));
  INVX1    g12791(.A(new_n12855_), .Y(new_n12856_));
  OAI21X1  g12792(.A0(new_n12856_), .A1(new_n3906_), .B0(new_n12852_), .Y(new_n12857_));
  XOR2X1   g12793(.A(new_n12857_), .B(\a[14] ), .Y(new_n12858_));
  XOR2X1   g12794(.A(new_n12217_), .B(new_n12216_), .Y(new_n12859_));
  AOI22X1  g12795(.A0(new_n12104_), .A1(new_n3628_), .B0(new_n12102_), .B1(new_n3908_), .Y(new_n12860_));
  OAI21X1  g12796(.A0(new_n12840_), .A1(new_n3983_), .B0(new_n12860_), .Y(new_n12861_));
  AOI21X1  g12797(.A0(new_n12859_), .A1(new_n3624_), .B0(new_n12861_), .Y(new_n12862_));
  XOR2X1   g12798(.A(new_n12862_), .B(\a[14] ), .Y(new_n12863_));
  INVX1    g12799(.A(new_n12863_), .Y(new_n12864_));
  XOR2X1   g12800(.A(new_n12835_), .B(new_n12834_), .Y(new_n12865_));
  AND2X1   g12801(.A(new_n12865_), .B(new_n12864_), .Y(new_n12866_));
  XOR2X1   g12802(.A(new_n12865_), .B(new_n12863_), .Y(new_n12867_));
  INVX1    g12803(.A(new_n12867_), .Y(new_n12868_));
  AOI22X1  g12804(.A0(new_n12107_), .A1(new_n3628_), .B0(new_n12104_), .B1(new_n3908_), .Y(new_n12869_));
  OAI21X1  g12805(.A0(new_n12306_), .A1(new_n3983_), .B0(new_n12869_), .Y(new_n12870_));
  AOI21X1  g12806(.A0(new_n12305_), .A1(new_n3624_), .B0(new_n12870_), .Y(new_n12871_));
  XOR2X1   g12807(.A(new_n12871_), .B(\a[14] ), .Y(new_n12872_));
  INVX1    g12808(.A(new_n12833_), .Y(new_n12873_));
  XOR2X1   g12809(.A(new_n12873_), .B(new_n12832_), .Y(new_n12874_));
  OR2X1    g12810(.A(new_n12874_), .B(new_n12872_), .Y(new_n12875_));
  XOR2X1   g12811(.A(new_n12874_), .B(new_n12872_), .Y(new_n12876_));
  INVX1    g12812(.A(new_n12876_), .Y(new_n12877_));
  INVX1    g12813(.A(new_n12727_), .Y(new_n12878_));
  XOR2X1   g12814(.A(new_n12830_), .B(new_n12878_), .Y(new_n12879_));
  OAI22X1  g12815(.A0(new_n12111_), .A1(new_n3627_), .B0(new_n12109_), .B1(new_n3907_), .Y(new_n12880_));
  AOI21X1  g12816(.A0(new_n12104_), .A1(new_n3984_), .B0(new_n12880_), .Y(new_n12881_));
  OAI21X1  g12817(.A0(new_n12693_), .A1(new_n3906_), .B0(new_n12881_), .Y(new_n12882_));
  XOR2X1   g12818(.A(new_n12882_), .B(new_n2529_), .Y(new_n12883_));
  NOR2X1   g12819(.A(new_n12883_), .B(new_n12879_), .Y(new_n12884_));
  XOR2X1   g12820(.A(new_n12829_), .B(new_n12735_), .Y(new_n12885_));
  INVX1    g12821(.A(new_n12885_), .Y(new_n12886_));
  OAI22X1  g12822(.A0(new_n12113_), .A1(new_n3627_), .B0(new_n12111_), .B1(new_n3907_), .Y(new_n12887_));
  AOI21X1  g12823(.A0(new_n12107_), .A1(new_n3984_), .B0(new_n12887_), .Y(new_n12888_));
  OAI21X1  g12824(.A0(new_n12708_), .A1(new_n3906_), .B0(new_n12888_), .Y(new_n12889_));
  XOR2X1   g12825(.A(new_n12889_), .B(new_n2529_), .Y(new_n12890_));
  OR2X1    g12826(.A(new_n12890_), .B(new_n12886_), .Y(new_n12891_));
  XOR2X1   g12827(.A(new_n12828_), .B(new_n12745_), .Y(new_n12892_));
  OAI22X1  g12828(.A0(new_n12117_), .A1(new_n3627_), .B0(new_n12113_), .B1(new_n3907_), .Y(new_n12893_));
  AOI21X1  g12829(.A0(new_n12208_), .A1(new_n3984_), .B0(new_n12893_), .Y(new_n12894_));
  OAI21X1  g12830(.A0(new_n12685_), .A1(new_n3906_), .B0(new_n12894_), .Y(new_n12895_));
  XOR2X1   g12831(.A(new_n12895_), .B(\a[14] ), .Y(new_n12896_));
  AOI22X1  g12832(.A0(new_n12133_), .A1(new_n3628_), .B0(new_n12720_), .B1(new_n3908_), .Y(new_n12897_));
  OAI21X1  g12833(.A0(new_n12113_), .A1(new_n3983_), .B0(new_n12897_), .Y(new_n12898_));
  AOI21X1  g12834(.A0(new_n12719_), .A1(new_n3624_), .B0(new_n12898_), .Y(new_n12899_));
  XOR2X1   g12835(.A(new_n12899_), .B(\a[14] ), .Y(new_n12900_));
  INVX1    g12836(.A(new_n12900_), .Y(new_n12901_));
  XOR2X1   g12837(.A(new_n12827_), .B(new_n12826_), .Y(new_n12902_));
  XOR2X1   g12838(.A(new_n12902_), .B(new_n12900_), .Y(new_n12903_));
  AOI22X1  g12839(.A0(new_n12138_), .A1(new_n3628_), .B0(new_n12133_), .B1(new_n3908_), .Y(new_n12904_));
  OAI21X1  g12840(.A0(new_n12117_), .A1(new_n3983_), .B0(new_n12904_), .Y(new_n12905_));
  AOI21X1  g12841(.A0(new_n12526_), .A1(new_n3624_), .B0(new_n12905_), .Y(new_n12906_));
  XOR2X1   g12842(.A(new_n12906_), .B(\a[14] ), .Y(new_n12907_));
  INVX1    g12843(.A(new_n12825_), .Y(new_n12908_));
  XOR2X1   g12844(.A(new_n12908_), .B(new_n12824_), .Y(new_n12909_));
  NOR2X1   g12845(.A(new_n12909_), .B(new_n12907_), .Y(new_n12910_));
  XOR2X1   g12846(.A(new_n12909_), .B(new_n12907_), .Y(new_n12911_));
  AOI22X1  g12847(.A0(new_n12141_), .A1(new_n3628_), .B0(new_n12138_), .B1(new_n3908_), .Y(new_n12912_));
  OAI21X1  g12848(.A0(new_n12134_), .A1(new_n3983_), .B0(new_n12912_), .Y(new_n12913_));
  AOI21X1  g12849(.A0(new_n12536_), .A1(new_n3624_), .B0(new_n12913_), .Y(new_n12914_));
  XOR2X1   g12850(.A(new_n12914_), .B(\a[14] ), .Y(new_n12915_));
  AND2X1   g12851(.A(new_n12821_), .B(new_n12773_), .Y(new_n12916_));
  INVX1    g12852(.A(new_n12822_), .Y(new_n12917_));
  XOR2X1   g12853(.A(new_n12917_), .B(new_n12916_), .Y(new_n12918_));
  OR2X1    g12854(.A(new_n12918_), .B(new_n12915_), .Y(new_n12919_));
  XOR2X1   g12855(.A(new_n12918_), .B(new_n12915_), .Y(new_n12920_));
  INVX1    g12856(.A(new_n12920_), .Y(new_n12921_));
  INVX1    g12857(.A(new_n12774_), .Y(new_n12922_));
  XOR2X1   g12858(.A(new_n12820_), .B(new_n12922_), .Y(new_n12923_));
  AOI22X1  g12859(.A0(new_n12144_), .A1(new_n3628_), .B0(new_n12141_), .B1(new_n3908_), .Y(new_n12924_));
  OAI21X1  g12860(.A0(new_n12314_), .A1(new_n3983_), .B0(new_n12924_), .Y(new_n12925_));
  AOI21X1  g12861(.A0(new_n12313_), .A1(new_n3624_), .B0(new_n12925_), .Y(new_n12926_));
  XOR2X1   g12862(.A(new_n12926_), .B(\a[14] ), .Y(new_n12927_));
  NOR2X1   g12863(.A(new_n12927_), .B(new_n12923_), .Y(new_n12928_));
  XOR2X1   g12864(.A(new_n12819_), .B(new_n12818_), .Y(new_n12929_));
  INVX1    g12865(.A(new_n12929_), .Y(new_n12930_));
  OAI22X1  g12866(.A0(new_n12186_), .A1(new_n3627_), .B0(new_n12192_), .B1(new_n3907_), .Y(new_n12931_));
  AOI21X1  g12867(.A0(new_n12141_), .A1(new_n3984_), .B0(new_n12931_), .Y(new_n12932_));
  OAI21X1  g12868(.A0(new_n12444_), .A1(new_n3906_), .B0(new_n12932_), .Y(new_n12933_));
  XOR2X1   g12869(.A(new_n12933_), .B(new_n2529_), .Y(new_n12934_));
  OR2X1    g12870(.A(new_n12934_), .B(new_n12930_), .Y(new_n12935_));
  XOR2X1   g12871(.A(new_n12816_), .B(new_n12791_), .Y(new_n12936_));
  INVX1    g12872(.A(new_n12936_), .Y(new_n12937_));
  OAI22X1  g12873(.A0(new_n12322_), .A1(new_n3627_), .B0(new_n12186_), .B1(new_n3907_), .Y(new_n12938_));
  AOI21X1  g12874(.A0(new_n12144_), .A1(new_n3984_), .B0(new_n12938_), .Y(new_n12939_));
  OAI21X1  g12875(.A0(new_n12453_), .A1(new_n3906_), .B0(new_n12939_), .Y(new_n12940_));
  XOR2X1   g12876(.A(new_n12940_), .B(new_n2529_), .Y(new_n12941_));
  NOR2X1   g12877(.A(new_n12941_), .B(new_n12937_), .Y(new_n12942_));
  AOI22X1  g12878(.A0(new_n12155_), .A1(new_n3628_), .B0(new_n12151_), .B1(new_n3908_), .Y(new_n12943_));
  OAI21X1  g12879(.A0(new_n12186_), .A1(new_n3983_), .B0(new_n12943_), .Y(new_n12944_));
  AOI21X1  g12880(.A0(new_n12430_), .A1(new_n3624_), .B0(new_n12944_), .Y(new_n12945_));
  XOR2X1   g12881(.A(new_n12945_), .B(\a[14] ), .Y(new_n12946_));
  INVX1    g12882(.A(new_n12946_), .Y(new_n12947_));
  XOR2X1   g12883(.A(new_n12815_), .B(new_n12814_), .Y(new_n12948_));
  NAND2X1  g12884(.A(new_n12948_), .B(new_n12947_), .Y(new_n12949_));
  XOR2X1   g12885(.A(new_n12948_), .B(new_n12946_), .Y(new_n12950_));
  XOR2X1   g12886(.A(new_n12812_), .B(new_n2445_), .Y(new_n12951_));
  XOR2X1   g12887(.A(new_n12951_), .B(new_n12809_), .Y(new_n12952_));
  AOI22X1  g12888(.A0(new_n12158_), .A1(new_n3628_), .B0(new_n12155_), .B1(new_n3908_), .Y(new_n12953_));
  OAI21X1  g12889(.A0(new_n12322_), .A1(new_n3983_), .B0(new_n12953_), .Y(new_n12954_));
  AOI21X1  g12890(.A0(new_n12321_), .A1(new_n3624_), .B0(new_n12954_), .Y(new_n12955_));
  XOR2X1   g12891(.A(new_n12955_), .B(\a[14] ), .Y(new_n12956_));
  NOR2X1   g12892(.A(new_n12956_), .B(new_n12952_), .Y(new_n12957_));
  AOI22X1  g12893(.A0(new_n12162_), .A1(new_n3628_), .B0(new_n12158_), .B1(new_n3908_), .Y(new_n12958_));
  OAI21X1  g12894(.A0(new_n12353_), .A1(new_n3983_), .B0(new_n12958_), .Y(new_n12959_));
  AOI21X1  g12895(.A0(new_n12352_), .A1(new_n3624_), .B0(new_n12959_), .Y(new_n12960_));
  XOR2X1   g12896(.A(new_n12960_), .B(\a[14] ), .Y(new_n12961_));
  NOR3X1   g12897(.A(new_n12802_), .B(new_n12801_), .C(new_n2445_), .Y(new_n12962_));
  XOR2X1   g12898(.A(new_n12805_), .B(\a[17] ), .Y(new_n12963_));
  NOR2X1   g12899(.A(new_n12963_), .B(new_n12962_), .Y(new_n12964_));
  NOR3X1   g12900(.A(new_n12964_), .B(new_n12961_), .C(new_n12806_), .Y(new_n12965_));
  XOR2X1   g12901(.A(new_n12963_), .B(new_n12962_), .Y(new_n12966_));
  XOR2X1   g12902(.A(new_n12966_), .B(new_n12961_), .Y(new_n12967_));
  NOR2X1   g12903(.A(new_n12802_), .B(new_n2445_), .Y(new_n12968_));
  XOR2X1   g12904(.A(new_n12968_), .B(new_n12801_), .Y(new_n12969_));
  OAI22X1  g12905(.A0(new_n12168_), .A1(new_n3627_), .B0(new_n12329_), .B1(new_n3907_), .Y(new_n12970_));
  AOI21X1  g12906(.A0(new_n12158_), .A1(new_n3984_), .B0(new_n12970_), .Y(new_n12971_));
  OAI21X1  g12907(.A0(new_n12368_), .A1(new_n3906_), .B0(new_n12971_), .Y(new_n12972_));
  XOR2X1   g12908(.A(new_n12972_), .B(new_n2529_), .Y(new_n12973_));
  NOR2X1   g12909(.A(new_n12973_), .B(new_n12969_), .Y(new_n12974_));
  OAI22X1  g12910(.A0(new_n12176_), .A1(new_n3907_), .B0(new_n12170_), .B1(new_n3983_), .Y(new_n12975_));
  AOI21X1  g12911(.A0(new_n12337_), .A1(new_n3624_), .B0(new_n12975_), .Y(new_n12976_));
  XOR2X1   g12912(.A(new_n12976_), .B(\a[14] ), .Y(new_n12977_));
  AOI21X1  g12913(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n3621_), .Y(new_n12978_));
  OAI22X1  g12914(.A0(new_n12176_), .A1(new_n3627_), .B0(new_n12170_), .B1(new_n3907_), .Y(new_n12979_));
  AOI21X1  g12915(.A0(new_n12165_), .A1(new_n3984_), .B0(new_n12979_), .Y(new_n12980_));
  OAI21X1  g12916(.A0(new_n12344_), .A1(new_n3906_), .B0(new_n12980_), .Y(new_n12981_));
  NOR4X1   g12917(.A(new_n12981_), .B(new_n12978_), .C(new_n12977_), .D(new_n2529_), .Y(new_n12982_));
  NAND2X1  g12918(.A(new_n12982_), .B(new_n12802_), .Y(new_n12983_));
  INVX1    g12919(.A(new_n12982_), .Y(new_n12984_));
  XOR2X1   g12920(.A(new_n12984_), .B(new_n12802_), .Y(new_n12985_));
  AOI22X1  g12921(.A0(new_n12331_), .A1(new_n3628_), .B0(new_n12165_), .B1(new_n3908_), .Y(new_n12986_));
  OAI21X1  g12922(.A0(new_n12329_), .A1(new_n3983_), .B0(new_n12986_), .Y(new_n12987_));
  AOI21X1  g12923(.A0(new_n12328_), .A1(new_n3624_), .B0(new_n12987_), .Y(new_n12988_));
  XOR2X1   g12924(.A(new_n12988_), .B(\a[14] ), .Y(new_n12989_));
  OAI21X1  g12925(.A0(new_n12989_), .A1(new_n12985_), .B0(new_n12983_), .Y(new_n12990_));
  XOR2X1   g12926(.A(new_n12973_), .B(new_n12969_), .Y(new_n12991_));
  AOI21X1  g12927(.A0(new_n12991_), .A1(new_n12990_), .B0(new_n12974_), .Y(new_n12992_));
  NOR2X1   g12928(.A(new_n12992_), .B(new_n12967_), .Y(new_n12993_));
  OR2X1    g12929(.A(new_n12993_), .B(new_n12965_), .Y(new_n12994_));
  XOR2X1   g12930(.A(new_n12956_), .B(new_n12952_), .Y(new_n12995_));
  AOI21X1  g12931(.A0(new_n12995_), .A1(new_n12994_), .B0(new_n12957_), .Y(new_n12996_));
  OR2X1    g12932(.A(new_n12996_), .B(new_n12950_), .Y(new_n12997_));
  XOR2X1   g12933(.A(new_n12941_), .B(new_n12936_), .Y(new_n12998_));
  AOI21X1  g12934(.A0(new_n12997_), .A1(new_n12949_), .B0(new_n12998_), .Y(new_n12999_));
  NOR2X1   g12935(.A(new_n12999_), .B(new_n12942_), .Y(new_n13000_));
  XOR2X1   g12936(.A(new_n12934_), .B(new_n12929_), .Y(new_n13001_));
  OAI21X1  g12937(.A0(new_n13001_), .A1(new_n13000_), .B0(new_n12935_), .Y(new_n13002_));
  XOR2X1   g12938(.A(new_n12927_), .B(new_n12923_), .Y(new_n13003_));
  AOI21X1  g12939(.A0(new_n13003_), .A1(new_n13002_), .B0(new_n12928_), .Y(new_n13004_));
  OAI21X1  g12940(.A0(new_n13004_), .A1(new_n12921_), .B0(new_n12919_), .Y(new_n13005_));
  AOI21X1  g12941(.A0(new_n13005_), .A1(new_n12911_), .B0(new_n12910_), .Y(new_n13006_));
  NOR2X1   g12942(.A(new_n13006_), .B(new_n12903_), .Y(new_n13007_));
  AOI21X1  g12943(.A0(new_n12902_), .A1(new_n12901_), .B0(new_n13007_), .Y(new_n13008_));
  XOR2X1   g12944(.A(new_n12895_), .B(new_n2529_), .Y(new_n13009_));
  XOR2X1   g12945(.A(new_n13009_), .B(new_n12892_), .Y(new_n13010_));
  NOR2X1   g12946(.A(new_n13010_), .B(new_n13008_), .Y(new_n13011_));
  AOI21X1  g12947(.A0(new_n12896_), .A1(new_n12892_), .B0(new_n13011_), .Y(new_n13012_));
  XOR2X1   g12948(.A(new_n12890_), .B(new_n12885_), .Y(new_n13013_));
  OAI21X1  g12949(.A0(new_n13013_), .A1(new_n13012_), .B0(new_n12891_), .Y(new_n13014_));
  XOR2X1   g12950(.A(new_n12883_), .B(new_n12879_), .Y(new_n13015_));
  AOI21X1  g12951(.A0(new_n13015_), .A1(new_n13014_), .B0(new_n12884_), .Y(new_n13016_));
  OAI21X1  g12952(.A0(new_n13016_), .A1(new_n12877_), .B0(new_n12875_), .Y(new_n13017_));
  AOI21X1  g12953(.A0(new_n13017_), .A1(new_n12868_), .B0(new_n12866_), .Y(new_n13018_));
  XOR2X1   g12954(.A(new_n12857_), .B(new_n2529_), .Y(new_n13019_));
  XOR2X1   g12955(.A(new_n13019_), .B(new_n12850_), .Y(new_n13020_));
  NOR2X1   g12956(.A(new_n13020_), .B(new_n13018_), .Y(new_n13021_));
  AOI21X1  g12957(.A0(new_n12858_), .A1(new_n12850_), .B0(new_n13021_), .Y(new_n13022_));
  XOR2X1   g12958(.A(new_n12847_), .B(new_n2529_), .Y(new_n13023_));
  XOR2X1   g12959(.A(new_n13023_), .B(new_n12838_), .Y(new_n13024_));
  NOR2X1   g12960(.A(new_n13024_), .B(new_n13022_), .Y(new_n13025_));
  NOR2X1   g12961(.A(new_n13025_), .B(new_n12849_), .Y(new_n13026_));
  AOI22X1  g12962(.A0(new_n12104_), .A1(new_n3232_), .B0(new_n12102_), .B1(new_n3390_), .Y(new_n13027_));
  OAI21X1  g12963(.A0(new_n12840_), .A1(new_n3545_), .B0(new_n13027_), .Y(new_n13028_));
  AOI21X1  g12964(.A0(new_n12859_), .A1(new_n3234_), .B0(new_n13028_), .Y(new_n13029_));
  XOR2X1   g12965(.A(new_n13029_), .B(\a[17] ), .Y(new_n13030_));
  XOR2X1   g12966(.A(new_n12686_), .B(\a[20] ), .Y(new_n13031_));
  NOR2X1   g12967(.A(new_n12688_), .B(new_n12633_), .Y(new_n13032_));
  AOI21X1  g12968(.A0(new_n13031_), .A1(new_n12679_), .B0(new_n13032_), .Y(new_n13033_));
  AOI22X1  g12969(.A0(new_n12138_), .A1(new_n2657_), .B0(new_n12133_), .B1(new_n2696_), .Y(new_n13034_));
  OAI21X1  g12970(.A0(new_n12117_), .A1(new_n2753_), .B0(new_n13034_), .Y(new_n13035_));
  AOI21X1  g12971(.A0(new_n12526_), .A1(new_n2658_), .B0(new_n13035_), .Y(new_n13036_));
  XOR2X1   g12972(.A(new_n13036_), .B(\a[23] ), .Y(new_n13037_));
  INVX1    g12973(.A(new_n12641_), .Y(new_n13038_));
  INVX1    g12974(.A(new_n12669_), .Y(new_n13039_));
  NOR2X1   g12975(.A(new_n12673_), .B(new_n13039_), .Y(new_n13040_));
  INVX1    g12976(.A(new_n13040_), .Y(new_n13041_));
  OAI21X1  g12977(.A0(new_n12674_), .A1(new_n13038_), .B0(new_n13041_), .Y(new_n13042_));
  AOI22X1  g12978(.A0(new_n12158_), .A1(new_n2185_), .B0(new_n12155_), .B1(new_n2095_), .Y(new_n13043_));
  OAI21X1  g12979(.A0(new_n12322_), .A1(new_n2140_), .B0(new_n13043_), .Y(new_n13044_));
  AOI21X1  g12980(.A0(new_n12321_), .A1(new_n2062_), .B0(new_n13044_), .Y(new_n13045_));
  XOR2X1   g12981(.A(new_n13045_), .B(\a[29] ), .Y(new_n13046_));
  NOR3X1   g12982(.A(new_n12661_), .B(new_n12419_), .C(new_n12416_), .Y(new_n13047_));
  AOI21X1  g12983(.A0(new_n12662_), .A1(new_n12648_), .B0(new_n13047_), .Y(new_n13048_));
  INVX1    g12984(.A(new_n13048_), .Y(new_n13049_));
  NOR4X1   g12985(.A(new_n1142_), .B(new_n582_), .C(new_n537_), .D(new_n515_), .Y(new_n13050_));
  NOR3X1   g12986(.A(new_n465_), .B(new_n274_), .C(new_n118_), .Y(new_n13051_));
  NOR4X1   g12987(.A(new_n885_), .B(new_n187_), .C(new_n449_), .D(new_n114_), .Y(new_n13052_));
  NAND3X1  g12988(.A(new_n13052_), .B(new_n13051_), .C(new_n13050_), .Y(new_n13053_));
  OR4X1    g12989(.A(new_n2920_), .B(new_n2506_), .C(new_n1540_), .D(new_n1203_), .Y(new_n13054_));
  OR4X1    g12990(.A(new_n13054_), .B(new_n13053_), .C(new_n3042_), .D(new_n2003_), .Y(new_n13055_));
  NOR4X1   g12991(.A(new_n13055_), .B(new_n1360_), .C(new_n810_), .D(new_n438_), .Y(new_n13056_));
  INVX1    g12992(.A(new_n13056_), .Y(new_n13057_));
  AOI22X1  g12993(.A0(new_n12331_), .A1(new_n1890_), .B0(new_n12165_), .B1(new_n1884_), .Y(new_n13058_));
  OAI21X1  g12994(.A0(new_n12329_), .A1(new_n3498_), .B0(new_n13058_), .Y(new_n13059_));
  AOI21X1  g12995(.A0(new_n12328_), .A1(new_n407_), .B0(new_n13059_), .Y(new_n13060_));
  XOR2X1   g12996(.A(new_n13060_), .B(new_n13057_), .Y(new_n13061_));
  XOR2X1   g12997(.A(new_n13061_), .B(new_n13049_), .Y(new_n13062_));
  XOR2X1   g12998(.A(new_n13062_), .B(new_n13046_), .Y(new_n13063_));
  OR2X1    g12999(.A(new_n12663_), .B(new_n12645_), .Y(new_n13064_));
  OAI21X1  g13000(.A0(new_n12668_), .A1(new_n12665_), .B0(new_n13064_), .Y(new_n13065_));
  XOR2X1   g13001(.A(new_n13065_), .B(new_n13063_), .Y(new_n13066_));
  OAI22X1  g13002(.A0(new_n12186_), .A1(new_n2666_), .B0(new_n12192_), .B1(new_n2419_), .Y(new_n13067_));
  AOI21X1  g13003(.A0(new_n12141_), .A1(new_n2423_), .B0(new_n13067_), .Y(new_n13068_));
  OAI21X1  g13004(.A0(new_n12444_), .A1(new_n2665_), .B0(new_n13068_), .Y(new_n13069_));
  XOR2X1   g13005(.A(new_n13069_), .B(new_n89_), .Y(new_n13070_));
  XOR2X1   g13006(.A(new_n13070_), .B(new_n13066_), .Y(new_n13071_));
  XOR2X1   g13007(.A(new_n13071_), .B(new_n13042_), .Y(new_n13072_));
  XOR2X1   g13008(.A(new_n13072_), .B(new_n13037_), .Y(new_n13073_));
  INVX1    g13009(.A(new_n13073_), .Y(new_n13074_));
  NOR2X1   g13010(.A(new_n12675_), .B(new_n12637_), .Y(new_n13075_));
  AOI21X1  g13011(.A0(new_n12678_), .A1(new_n12676_), .B0(new_n13075_), .Y(new_n13076_));
  XOR2X1   g13012(.A(new_n13076_), .B(new_n13074_), .Y(new_n13077_));
  OAI22X1  g13013(.A0(new_n12113_), .A1(new_n3250_), .B0(new_n12111_), .B1(new_n3144_), .Y(new_n13078_));
  AOI21X1  g13014(.A0(new_n12107_), .A1(new_n3146_), .B0(new_n13078_), .Y(new_n13079_));
  OAI21X1  g13015(.A0(new_n12708_), .A1(new_n3098_), .B0(new_n13079_), .Y(new_n13080_));
  XOR2X1   g13016(.A(new_n13080_), .B(new_n1920_), .Y(new_n13081_));
  XOR2X1   g13017(.A(new_n13081_), .B(new_n13077_), .Y(new_n13082_));
  INVX1    g13018(.A(new_n13082_), .Y(new_n13083_));
  XOR2X1   g13019(.A(new_n13083_), .B(new_n13033_), .Y(new_n13084_));
  XOR2X1   g13020(.A(new_n13084_), .B(new_n13030_), .Y(new_n13085_));
  INVX1    g13021(.A(new_n13085_), .Y(new_n13086_));
  NOR2X1   g13022(.A(new_n12690_), .B(new_n12310_), .Y(new_n13087_));
  AOI21X1  g13023(.A0(new_n12837_), .A1(new_n12691_), .B0(new_n13087_), .Y(new_n13088_));
  XOR2X1   g13024(.A(new_n13088_), .B(new_n13086_), .Y(new_n13089_));
  INVX1    g13025(.A(new_n12095_), .Y(new_n13090_));
  OAI22X1  g13026(.A0(new_n12839_), .A1(new_n3627_), .B0(new_n13090_), .B1(new_n3907_), .Y(new_n13091_));
  AOI21X1  g13027(.A0(new_n12093_), .A1(new_n3984_), .B0(new_n13091_), .Y(new_n13092_));
  XOR2X1   g13028(.A(new_n12224_), .B(new_n12222_), .Y(new_n13093_));
  INVX1    g13029(.A(new_n13093_), .Y(new_n13094_));
  OAI21X1  g13030(.A0(new_n13094_), .A1(new_n3906_), .B0(new_n13092_), .Y(new_n13095_));
  XOR2X1   g13031(.A(new_n13095_), .B(new_n2529_), .Y(new_n13096_));
  XOR2X1   g13032(.A(new_n13096_), .B(new_n13089_), .Y(new_n13097_));
  INVX1    g13033(.A(new_n13097_), .Y(new_n13098_));
  XOR2X1   g13034(.A(new_n13098_), .B(new_n13026_), .Y(new_n13099_));
  XOR2X1   g13035(.A(new_n13099_), .B(new_n12302_), .Y(new_n13100_));
  XOR2X1   g13036(.A(new_n12090_), .B(new_n12088_), .Y(new_n13101_));
  OR2X1    g13037(.A(new_n13101_), .B(new_n12227_), .Y(new_n13102_));
  OAI21X1  g13038(.A0(new_n12229_), .A1(new_n12228_), .B0(new_n13102_), .Y(new_n13103_));
  INVX1    g13039(.A(new_n12088_), .Y(new_n13104_));
  AOI22X1  g13040(.A0(new_n12093_), .A1(new_n4078_), .B0(new_n12090_), .B1(new_n4247_), .Y(new_n13105_));
  OAI21X1  g13041(.A0(new_n13104_), .A1(new_n4427_), .B0(new_n13105_), .Y(new_n13106_));
  AOI21X1  g13042(.A0(new_n13103_), .A1(new_n4080_), .B0(new_n13106_), .Y(new_n13107_));
  XOR2X1   g13043(.A(new_n13107_), .B(\a[11] ), .Y(new_n13108_));
  INVX1    g13044(.A(new_n13024_), .Y(new_n13109_));
  XOR2X1   g13045(.A(new_n13109_), .B(new_n13022_), .Y(new_n13110_));
  NOR2X1   g13046(.A(new_n13110_), .B(new_n13108_), .Y(new_n13111_));
  XOR2X1   g13047(.A(new_n13110_), .B(new_n13108_), .Y(new_n13112_));
  XOR2X1   g13048(.A(new_n12093_), .B(new_n12090_), .Y(new_n13113_));
  INVX1    g13049(.A(new_n13113_), .Y(new_n13114_));
  AND2X1   g13050(.A(new_n13114_), .B(new_n12225_), .Y(new_n13115_));
  AOI21X1  g13051(.A0(new_n12227_), .A1(new_n12226_), .B0(new_n13115_), .Y(new_n13116_));
  INVX1    g13052(.A(new_n13116_), .Y(new_n13117_));
  INVX1    g13053(.A(new_n12090_), .Y(new_n13118_));
  AOI22X1  g13054(.A0(new_n12095_), .A1(new_n4078_), .B0(new_n12093_), .B1(new_n4247_), .Y(new_n13119_));
  OAI21X1  g13055(.A0(new_n13118_), .A1(new_n4427_), .B0(new_n13119_), .Y(new_n13120_));
  AOI21X1  g13056(.A0(new_n13117_), .A1(new_n4080_), .B0(new_n13120_), .Y(new_n13121_));
  XOR2X1   g13057(.A(new_n13121_), .B(\a[11] ), .Y(new_n13122_));
  INVX1    g13058(.A(new_n13020_), .Y(new_n13123_));
  XOR2X1   g13059(.A(new_n13123_), .B(new_n13018_), .Y(new_n13124_));
  NOR2X1   g13060(.A(new_n13124_), .B(new_n13122_), .Y(new_n13125_));
  INVX1    g13061(.A(new_n13125_), .Y(new_n13126_));
  XOR2X1   g13062(.A(new_n13124_), .B(new_n13122_), .Y(new_n13127_));
  INVX1    g13063(.A(new_n13127_), .Y(new_n13128_));
  XOR2X1   g13064(.A(new_n13017_), .B(new_n12867_), .Y(new_n13129_));
  OAI22X1  g13065(.A0(new_n12839_), .A1(new_n4077_), .B0(new_n13090_), .B1(new_n4246_), .Y(new_n13130_));
  AOI21X1  g13066(.A0(new_n12093_), .A1(new_n4428_), .B0(new_n13130_), .Y(new_n13131_));
  OAI21X1  g13067(.A0(new_n13094_), .A1(new_n4245_), .B0(new_n13131_), .Y(new_n13132_));
  XOR2X1   g13068(.A(new_n13132_), .B(new_n2911_), .Y(new_n13133_));
  NOR2X1   g13069(.A(new_n13133_), .B(new_n13129_), .Y(new_n13134_));
  XOR2X1   g13070(.A(new_n13016_), .B(new_n12877_), .Y(new_n13135_));
  OAI22X1  g13071(.A0(new_n12840_), .A1(new_n4077_), .B0(new_n12839_), .B1(new_n4246_), .Y(new_n13136_));
  AOI21X1  g13072(.A0(new_n12095_), .A1(new_n4428_), .B0(new_n13136_), .Y(new_n13137_));
  OAI21X1  g13073(.A0(new_n12846_), .A1(new_n4245_), .B0(new_n13137_), .Y(new_n13138_));
  XOR2X1   g13074(.A(new_n13138_), .B(\a[11] ), .Y(new_n13139_));
  NAND2X1  g13075(.A(new_n13139_), .B(new_n13135_), .Y(new_n13140_));
  AOI22X1  g13076(.A0(new_n12102_), .A1(new_n4078_), .B0(new_n12099_), .B1(new_n4247_), .Y(new_n13141_));
  OAI21X1  g13077(.A0(new_n12839_), .A1(new_n4427_), .B0(new_n13141_), .Y(new_n13142_));
  AOI21X1  g13078(.A0(new_n12855_), .A1(new_n4080_), .B0(new_n13142_), .Y(new_n13143_));
  XOR2X1   g13079(.A(new_n13143_), .B(\a[11] ), .Y(new_n13144_));
  INVX1    g13080(.A(new_n13144_), .Y(new_n13145_));
  XOR2X1   g13081(.A(new_n13015_), .B(new_n13014_), .Y(new_n13146_));
  XOR2X1   g13082(.A(new_n13146_), .B(new_n13144_), .Y(new_n13147_));
  AOI22X1  g13083(.A0(new_n12104_), .A1(new_n4078_), .B0(new_n12102_), .B1(new_n4247_), .Y(new_n13148_));
  OAI21X1  g13084(.A0(new_n12840_), .A1(new_n4427_), .B0(new_n13148_), .Y(new_n13149_));
  AOI21X1  g13085(.A0(new_n12859_), .A1(new_n4080_), .B0(new_n13149_), .Y(new_n13150_));
  XOR2X1   g13086(.A(new_n13150_), .B(\a[11] ), .Y(new_n13151_));
  INVX1    g13087(.A(new_n13013_), .Y(new_n13152_));
  XOR2X1   g13088(.A(new_n13152_), .B(new_n13012_), .Y(new_n13153_));
  NOR2X1   g13089(.A(new_n13153_), .B(new_n13151_), .Y(new_n13154_));
  XOR2X1   g13090(.A(new_n13153_), .B(new_n13151_), .Y(new_n13155_));
  INVX1    g13091(.A(new_n13155_), .Y(new_n13156_));
  AOI22X1  g13092(.A0(new_n12107_), .A1(new_n4078_), .B0(new_n12104_), .B1(new_n4247_), .Y(new_n13157_));
  OAI21X1  g13093(.A0(new_n12306_), .A1(new_n4427_), .B0(new_n13157_), .Y(new_n13158_));
  AOI21X1  g13094(.A0(new_n12305_), .A1(new_n4080_), .B0(new_n13158_), .Y(new_n13159_));
  XOR2X1   g13095(.A(new_n13159_), .B(\a[11] ), .Y(new_n13160_));
  INVX1    g13096(.A(new_n13010_), .Y(new_n13161_));
  XOR2X1   g13097(.A(new_n13161_), .B(new_n13008_), .Y(new_n13162_));
  OR2X1    g13098(.A(new_n13162_), .B(new_n13160_), .Y(new_n13163_));
  XOR2X1   g13099(.A(new_n13162_), .B(new_n13160_), .Y(new_n13164_));
  INVX1    g13100(.A(new_n13164_), .Y(new_n13165_));
  INVX1    g13101(.A(new_n12903_), .Y(new_n13166_));
  XOR2X1   g13102(.A(new_n13006_), .B(new_n13166_), .Y(new_n13167_));
  OAI22X1  g13103(.A0(new_n12111_), .A1(new_n4077_), .B0(new_n12109_), .B1(new_n4246_), .Y(new_n13168_));
  AOI21X1  g13104(.A0(new_n12104_), .A1(new_n4428_), .B0(new_n13168_), .Y(new_n13169_));
  OAI21X1  g13105(.A0(new_n12693_), .A1(new_n4245_), .B0(new_n13169_), .Y(new_n13170_));
  XOR2X1   g13106(.A(new_n13170_), .B(new_n2911_), .Y(new_n13171_));
  NOR2X1   g13107(.A(new_n13171_), .B(new_n13167_), .Y(new_n13172_));
  XOR2X1   g13108(.A(new_n13005_), .B(new_n12911_), .Y(new_n13173_));
  INVX1    g13109(.A(new_n13173_), .Y(new_n13174_));
  OAI22X1  g13110(.A0(new_n12113_), .A1(new_n4077_), .B0(new_n12111_), .B1(new_n4246_), .Y(new_n13175_));
  AOI21X1  g13111(.A0(new_n12107_), .A1(new_n4428_), .B0(new_n13175_), .Y(new_n13176_));
  OAI21X1  g13112(.A0(new_n12708_), .A1(new_n4245_), .B0(new_n13176_), .Y(new_n13177_));
  XOR2X1   g13113(.A(new_n13177_), .B(new_n2911_), .Y(new_n13178_));
  OR2X1    g13114(.A(new_n13178_), .B(new_n13174_), .Y(new_n13179_));
  XOR2X1   g13115(.A(new_n13004_), .B(new_n12921_), .Y(new_n13180_));
  OAI22X1  g13116(.A0(new_n12117_), .A1(new_n4077_), .B0(new_n12113_), .B1(new_n4246_), .Y(new_n13181_));
  AOI21X1  g13117(.A0(new_n12208_), .A1(new_n4428_), .B0(new_n13181_), .Y(new_n13182_));
  OAI21X1  g13118(.A0(new_n12685_), .A1(new_n4245_), .B0(new_n13182_), .Y(new_n13183_));
  XOR2X1   g13119(.A(new_n13183_), .B(\a[11] ), .Y(new_n13184_));
  AOI22X1  g13120(.A0(new_n12133_), .A1(new_n4078_), .B0(new_n12720_), .B1(new_n4247_), .Y(new_n13185_));
  OAI21X1  g13121(.A0(new_n12113_), .A1(new_n4427_), .B0(new_n13185_), .Y(new_n13186_));
  AOI21X1  g13122(.A0(new_n12719_), .A1(new_n4080_), .B0(new_n13186_), .Y(new_n13187_));
  XOR2X1   g13123(.A(new_n13187_), .B(\a[11] ), .Y(new_n13188_));
  INVX1    g13124(.A(new_n13188_), .Y(new_n13189_));
  XOR2X1   g13125(.A(new_n13003_), .B(new_n13002_), .Y(new_n13190_));
  XOR2X1   g13126(.A(new_n13190_), .B(new_n13188_), .Y(new_n13191_));
  AOI22X1  g13127(.A0(new_n12138_), .A1(new_n4078_), .B0(new_n12133_), .B1(new_n4247_), .Y(new_n13192_));
  OAI21X1  g13128(.A0(new_n12117_), .A1(new_n4427_), .B0(new_n13192_), .Y(new_n13193_));
  AOI21X1  g13129(.A0(new_n12526_), .A1(new_n4080_), .B0(new_n13193_), .Y(new_n13194_));
  XOR2X1   g13130(.A(new_n13194_), .B(\a[11] ), .Y(new_n13195_));
  INVX1    g13131(.A(new_n13001_), .Y(new_n13196_));
  XOR2X1   g13132(.A(new_n13196_), .B(new_n13000_), .Y(new_n13197_));
  NOR2X1   g13133(.A(new_n13197_), .B(new_n13195_), .Y(new_n13198_));
  XOR2X1   g13134(.A(new_n13197_), .B(new_n13195_), .Y(new_n13199_));
  AOI22X1  g13135(.A0(new_n12141_), .A1(new_n4078_), .B0(new_n12138_), .B1(new_n4247_), .Y(new_n13200_));
  OAI21X1  g13136(.A0(new_n12134_), .A1(new_n4427_), .B0(new_n13200_), .Y(new_n13201_));
  AOI21X1  g13137(.A0(new_n12536_), .A1(new_n4080_), .B0(new_n13201_), .Y(new_n13202_));
  XOR2X1   g13138(.A(new_n13202_), .B(\a[11] ), .Y(new_n13203_));
  AND2X1   g13139(.A(new_n12997_), .B(new_n12949_), .Y(new_n13204_));
  INVX1    g13140(.A(new_n12998_), .Y(new_n13205_));
  XOR2X1   g13141(.A(new_n13205_), .B(new_n13204_), .Y(new_n13206_));
  OR2X1    g13142(.A(new_n13206_), .B(new_n13203_), .Y(new_n13207_));
  XOR2X1   g13143(.A(new_n13206_), .B(new_n13203_), .Y(new_n13208_));
  INVX1    g13144(.A(new_n13208_), .Y(new_n13209_));
  INVX1    g13145(.A(new_n12950_), .Y(new_n13210_));
  XOR2X1   g13146(.A(new_n12996_), .B(new_n13210_), .Y(new_n13211_));
  AOI22X1  g13147(.A0(new_n12144_), .A1(new_n4078_), .B0(new_n12141_), .B1(new_n4247_), .Y(new_n13212_));
  OAI21X1  g13148(.A0(new_n12314_), .A1(new_n4427_), .B0(new_n13212_), .Y(new_n13213_));
  AOI21X1  g13149(.A0(new_n12313_), .A1(new_n4080_), .B0(new_n13213_), .Y(new_n13214_));
  XOR2X1   g13150(.A(new_n13214_), .B(\a[11] ), .Y(new_n13215_));
  NOR2X1   g13151(.A(new_n13215_), .B(new_n13211_), .Y(new_n13216_));
  XOR2X1   g13152(.A(new_n12995_), .B(new_n12994_), .Y(new_n13217_));
  INVX1    g13153(.A(new_n13217_), .Y(new_n13218_));
  OAI22X1  g13154(.A0(new_n12186_), .A1(new_n4077_), .B0(new_n12192_), .B1(new_n4246_), .Y(new_n13219_));
  AOI21X1  g13155(.A0(new_n12141_), .A1(new_n4428_), .B0(new_n13219_), .Y(new_n13220_));
  OAI21X1  g13156(.A0(new_n12444_), .A1(new_n4245_), .B0(new_n13220_), .Y(new_n13221_));
  XOR2X1   g13157(.A(new_n13221_), .B(new_n2911_), .Y(new_n13222_));
  OR2X1    g13158(.A(new_n13222_), .B(new_n13218_), .Y(new_n13223_));
  XOR2X1   g13159(.A(new_n12992_), .B(new_n12967_), .Y(new_n13224_));
  INVX1    g13160(.A(new_n13224_), .Y(new_n13225_));
  OAI22X1  g13161(.A0(new_n12322_), .A1(new_n4077_), .B0(new_n12186_), .B1(new_n4246_), .Y(new_n13226_));
  AOI21X1  g13162(.A0(new_n12144_), .A1(new_n4428_), .B0(new_n13226_), .Y(new_n13227_));
  OAI21X1  g13163(.A0(new_n12453_), .A1(new_n4245_), .B0(new_n13227_), .Y(new_n13228_));
  XOR2X1   g13164(.A(new_n13228_), .B(new_n2911_), .Y(new_n13229_));
  NOR2X1   g13165(.A(new_n13229_), .B(new_n13225_), .Y(new_n13230_));
  AOI22X1  g13166(.A0(new_n12155_), .A1(new_n4078_), .B0(new_n12151_), .B1(new_n4247_), .Y(new_n13231_));
  OAI21X1  g13167(.A0(new_n12186_), .A1(new_n4427_), .B0(new_n13231_), .Y(new_n13232_));
  AOI21X1  g13168(.A0(new_n12430_), .A1(new_n4080_), .B0(new_n13232_), .Y(new_n13233_));
  XOR2X1   g13169(.A(new_n13233_), .B(\a[11] ), .Y(new_n13234_));
  INVX1    g13170(.A(new_n13234_), .Y(new_n13235_));
  XOR2X1   g13171(.A(new_n12991_), .B(new_n12990_), .Y(new_n13236_));
  NAND2X1  g13172(.A(new_n13236_), .B(new_n13235_), .Y(new_n13237_));
  XOR2X1   g13173(.A(new_n13236_), .B(new_n13234_), .Y(new_n13238_));
  XOR2X1   g13174(.A(new_n12988_), .B(new_n2529_), .Y(new_n13239_));
  XOR2X1   g13175(.A(new_n13239_), .B(new_n12985_), .Y(new_n13240_));
  AOI22X1  g13176(.A0(new_n12158_), .A1(new_n4078_), .B0(new_n12155_), .B1(new_n4247_), .Y(new_n13241_));
  OAI21X1  g13177(.A0(new_n12322_), .A1(new_n4427_), .B0(new_n13241_), .Y(new_n13242_));
  AOI21X1  g13178(.A0(new_n12321_), .A1(new_n4080_), .B0(new_n13242_), .Y(new_n13243_));
  XOR2X1   g13179(.A(new_n13243_), .B(\a[11] ), .Y(new_n13244_));
  NOR2X1   g13180(.A(new_n13244_), .B(new_n13240_), .Y(new_n13245_));
  AOI22X1  g13181(.A0(new_n12162_), .A1(new_n4078_), .B0(new_n12158_), .B1(new_n4247_), .Y(new_n13246_));
  OAI21X1  g13182(.A0(new_n12353_), .A1(new_n4427_), .B0(new_n13246_), .Y(new_n13247_));
  AOI21X1  g13183(.A0(new_n12352_), .A1(new_n4080_), .B0(new_n13247_), .Y(new_n13248_));
  XOR2X1   g13184(.A(new_n13248_), .B(\a[11] ), .Y(new_n13249_));
  NOR3X1   g13185(.A(new_n12978_), .B(new_n12977_), .C(new_n2529_), .Y(new_n13250_));
  XOR2X1   g13186(.A(new_n12981_), .B(\a[14] ), .Y(new_n13251_));
  NOR2X1   g13187(.A(new_n13251_), .B(new_n13250_), .Y(new_n13252_));
  NOR3X1   g13188(.A(new_n13252_), .B(new_n13249_), .C(new_n12982_), .Y(new_n13253_));
  XOR2X1   g13189(.A(new_n13251_), .B(new_n13250_), .Y(new_n13254_));
  XOR2X1   g13190(.A(new_n13254_), .B(new_n13249_), .Y(new_n13255_));
  NOR2X1   g13191(.A(new_n12978_), .B(new_n2529_), .Y(new_n13256_));
  XOR2X1   g13192(.A(new_n13256_), .B(new_n12977_), .Y(new_n13257_));
  OAI22X1  g13193(.A0(new_n12168_), .A1(new_n4077_), .B0(new_n12329_), .B1(new_n4246_), .Y(new_n13258_));
  AOI21X1  g13194(.A0(new_n12158_), .A1(new_n4428_), .B0(new_n13258_), .Y(new_n13259_));
  OAI21X1  g13195(.A0(new_n12368_), .A1(new_n4245_), .B0(new_n13259_), .Y(new_n13260_));
  XOR2X1   g13196(.A(new_n13260_), .B(new_n2911_), .Y(new_n13261_));
  NOR2X1   g13197(.A(new_n13261_), .B(new_n13257_), .Y(new_n13262_));
  OAI22X1  g13198(.A0(new_n12176_), .A1(new_n4246_), .B0(new_n12170_), .B1(new_n4427_), .Y(new_n13263_));
  AOI21X1  g13199(.A0(new_n12337_), .A1(new_n4080_), .B0(new_n13263_), .Y(new_n13264_));
  XOR2X1   g13200(.A(new_n13264_), .B(\a[11] ), .Y(new_n13265_));
  AOI21X1  g13201(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n4073_), .Y(new_n13266_));
  OAI22X1  g13202(.A0(new_n12176_), .A1(new_n4077_), .B0(new_n12170_), .B1(new_n4246_), .Y(new_n13267_));
  AOI21X1  g13203(.A0(new_n12165_), .A1(new_n4428_), .B0(new_n13267_), .Y(new_n13268_));
  OAI21X1  g13204(.A0(new_n12344_), .A1(new_n4245_), .B0(new_n13268_), .Y(new_n13269_));
  NOR4X1   g13205(.A(new_n13269_), .B(new_n13266_), .C(new_n13265_), .D(new_n2911_), .Y(new_n13270_));
  NAND2X1  g13206(.A(new_n13270_), .B(new_n12978_), .Y(new_n13271_));
  INVX1    g13207(.A(new_n13270_), .Y(new_n13272_));
  XOR2X1   g13208(.A(new_n13272_), .B(new_n12978_), .Y(new_n13273_));
  AOI22X1  g13209(.A0(new_n12331_), .A1(new_n4078_), .B0(new_n12165_), .B1(new_n4247_), .Y(new_n13274_));
  OAI21X1  g13210(.A0(new_n12329_), .A1(new_n4427_), .B0(new_n13274_), .Y(new_n13275_));
  AOI21X1  g13211(.A0(new_n12328_), .A1(new_n4080_), .B0(new_n13275_), .Y(new_n13276_));
  XOR2X1   g13212(.A(new_n13276_), .B(\a[11] ), .Y(new_n13277_));
  OAI21X1  g13213(.A0(new_n13277_), .A1(new_n13273_), .B0(new_n13271_), .Y(new_n13278_));
  XOR2X1   g13214(.A(new_n13261_), .B(new_n13257_), .Y(new_n13279_));
  AOI21X1  g13215(.A0(new_n13279_), .A1(new_n13278_), .B0(new_n13262_), .Y(new_n13280_));
  NOR2X1   g13216(.A(new_n13280_), .B(new_n13255_), .Y(new_n13281_));
  OR2X1    g13217(.A(new_n13281_), .B(new_n13253_), .Y(new_n13282_));
  XOR2X1   g13218(.A(new_n13244_), .B(new_n13240_), .Y(new_n13283_));
  AOI21X1  g13219(.A0(new_n13283_), .A1(new_n13282_), .B0(new_n13245_), .Y(new_n13284_));
  OR2X1    g13220(.A(new_n13284_), .B(new_n13238_), .Y(new_n13285_));
  XOR2X1   g13221(.A(new_n13229_), .B(new_n13224_), .Y(new_n13286_));
  AOI21X1  g13222(.A0(new_n13285_), .A1(new_n13237_), .B0(new_n13286_), .Y(new_n13287_));
  NOR2X1   g13223(.A(new_n13287_), .B(new_n13230_), .Y(new_n13288_));
  XOR2X1   g13224(.A(new_n13222_), .B(new_n13217_), .Y(new_n13289_));
  OAI21X1  g13225(.A0(new_n13289_), .A1(new_n13288_), .B0(new_n13223_), .Y(new_n13290_));
  XOR2X1   g13226(.A(new_n13215_), .B(new_n13211_), .Y(new_n13291_));
  AOI21X1  g13227(.A0(new_n13291_), .A1(new_n13290_), .B0(new_n13216_), .Y(new_n13292_));
  OAI21X1  g13228(.A0(new_n13292_), .A1(new_n13209_), .B0(new_n13207_), .Y(new_n13293_));
  AOI21X1  g13229(.A0(new_n13293_), .A1(new_n13199_), .B0(new_n13198_), .Y(new_n13294_));
  NOR2X1   g13230(.A(new_n13294_), .B(new_n13191_), .Y(new_n13295_));
  AOI21X1  g13231(.A0(new_n13190_), .A1(new_n13189_), .B0(new_n13295_), .Y(new_n13296_));
  XOR2X1   g13232(.A(new_n13183_), .B(new_n2911_), .Y(new_n13297_));
  XOR2X1   g13233(.A(new_n13297_), .B(new_n13180_), .Y(new_n13298_));
  NOR2X1   g13234(.A(new_n13298_), .B(new_n13296_), .Y(new_n13299_));
  AOI21X1  g13235(.A0(new_n13184_), .A1(new_n13180_), .B0(new_n13299_), .Y(new_n13300_));
  XOR2X1   g13236(.A(new_n13178_), .B(new_n13173_), .Y(new_n13301_));
  OAI21X1  g13237(.A0(new_n13301_), .A1(new_n13300_), .B0(new_n13179_), .Y(new_n13302_));
  XOR2X1   g13238(.A(new_n13171_), .B(new_n13167_), .Y(new_n13303_));
  AOI21X1  g13239(.A0(new_n13303_), .A1(new_n13302_), .B0(new_n13172_), .Y(new_n13304_));
  OR2X1    g13240(.A(new_n13304_), .B(new_n13165_), .Y(new_n13305_));
  AOI21X1  g13241(.A0(new_n13305_), .A1(new_n13163_), .B0(new_n13156_), .Y(new_n13306_));
  NOR2X1   g13242(.A(new_n13306_), .B(new_n13154_), .Y(new_n13307_));
  NOR2X1   g13243(.A(new_n13307_), .B(new_n13147_), .Y(new_n13308_));
  AOI21X1  g13244(.A0(new_n13146_), .A1(new_n13145_), .B0(new_n13308_), .Y(new_n13309_));
  XOR2X1   g13245(.A(new_n13138_), .B(new_n2911_), .Y(new_n13310_));
  XOR2X1   g13246(.A(new_n13310_), .B(new_n13135_), .Y(new_n13311_));
  OAI21X1  g13247(.A0(new_n13311_), .A1(new_n13309_), .B0(new_n13140_), .Y(new_n13312_));
  XOR2X1   g13248(.A(new_n13133_), .B(new_n13129_), .Y(new_n13313_));
  AOI21X1  g13249(.A0(new_n13313_), .A1(new_n13312_), .B0(new_n13134_), .Y(new_n13314_));
  OAI21X1  g13250(.A0(new_n13314_), .A1(new_n13128_), .B0(new_n13126_), .Y(new_n13315_));
  AOI21X1  g13251(.A0(new_n13315_), .A1(new_n13112_), .B0(new_n13111_), .Y(new_n13316_));
  INVX1    g13252(.A(new_n13316_), .Y(new_n13317_));
  XOR2X1   g13253(.A(new_n13317_), .B(new_n13100_), .Y(new_n13318_));
  INVX1    g13254(.A(new_n13318_), .Y(new_n13319_));
  INVX1    g13255(.A(new_n12081_), .Y(new_n13320_));
  INVX1    g13256(.A(new_n12083_), .Y(new_n13321_));
  OAI22X1  g13257(.A0(new_n13321_), .A1(new_n4634_), .B0(new_n13320_), .B1(new_n4869_), .Y(new_n13322_));
  AOI21X1  g13258(.A0(new_n12079_), .A1(new_n5097_), .B0(new_n13322_), .Y(new_n13323_));
  XOR2X1   g13259(.A(new_n12081_), .B(new_n12079_), .Y(new_n13324_));
  XOR2X1   g13260(.A(new_n13324_), .B(new_n12235_), .Y(new_n13325_));
  OAI21X1  g13261(.A0(new_n13325_), .A1(new_n4868_), .B0(new_n13323_), .Y(new_n13326_));
  XOR2X1   g13262(.A(new_n13326_), .B(new_n2995_), .Y(new_n13327_));
  XOR2X1   g13263(.A(new_n13315_), .B(new_n13112_), .Y(new_n13328_));
  OAI22X1  g13264(.A0(new_n12298_), .A1(new_n4634_), .B0(new_n13321_), .B1(new_n4869_), .Y(new_n13329_));
  AOI21X1  g13265(.A0(new_n12081_), .A1(new_n5097_), .B0(new_n13329_), .Y(new_n13330_));
  NOR2X1   g13266(.A(new_n12083_), .B(new_n12081_), .Y(new_n13331_));
  OAI21X1  g13267(.A0(new_n13331_), .A1(new_n12084_), .B0(new_n12233_), .Y(new_n13332_));
  NOR3X1   g13268(.A(new_n13331_), .B(new_n12233_), .C(new_n12084_), .Y(new_n13333_));
  INVX1    g13269(.A(new_n13333_), .Y(new_n13334_));
  AND2X1   g13270(.A(new_n13334_), .B(new_n13332_), .Y(new_n13335_));
  OAI21X1  g13271(.A0(new_n13335_), .A1(new_n4868_), .B0(new_n13330_), .Y(new_n13336_));
  XOR2X1   g13272(.A(new_n13336_), .B(\a[8] ), .Y(new_n13337_));
  AND2X1   g13273(.A(new_n13337_), .B(new_n13328_), .Y(new_n13338_));
  XOR2X1   g13274(.A(new_n13314_), .B(new_n13128_), .Y(new_n13339_));
  INVX1    g13275(.A(new_n13339_), .Y(new_n13340_));
  OAI22X1  g13276(.A0(new_n13104_), .A1(new_n4634_), .B0(new_n12298_), .B1(new_n4869_), .Y(new_n13341_));
  AOI21X1  g13277(.A0(new_n12083_), .A1(new_n5097_), .B0(new_n13341_), .Y(new_n13342_));
  XOR2X1   g13278(.A(new_n12085_), .B(new_n12083_), .Y(new_n13343_));
  OAI22X1  g13279(.A0(new_n12233_), .A1(new_n12232_), .B0(new_n13343_), .B1(new_n12231_), .Y(new_n13344_));
  INVX1    g13280(.A(new_n13344_), .Y(new_n13345_));
  OAI21X1  g13281(.A0(new_n13345_), .A1(new_n4868_), .B0(new_n13342_), .Y(new_n13346_));
  XOR2X1   g13282(.A(new_n13346_), .B(new_n2995_), .Y(new_n13347_));
  AOI22X1  g13283(.A0(new_n12090_), .A1(new_n4635_), .B0(new_n12088_), .B1(new_n4870_), .Y(new_n13348_));
  OAI21X1  g13284(.A0(new_n12298_), .A1(new_n5096_), .B0(new_n13348_), .Y(new_n13349_));
  AOI21X1  g13285(.A0(new_n12297_), .A1(new_n4637_), .B0(new_n13349_), .Y(new_n13350_));
  XOR2X1   g13286(.A(new_n13350_), .B(\a[8] ), .Y(new_n13351_));
  INVX1    g13287(.A(new_n13351_), .Y(new_n13352_));
  XOR2X1   g13288(.A(new_n13313_), .B(new_n13312_), .Y(new_n13353_));
  XOR2X1   g13289(.A(new_n13353_), .B(new_n13351_), .Y(new_n13354_));
  AOI22X1  g13290(.A0(new_n12093_), .A1(new_n4635_), .B0(new_n12090_), .B1(new_n4870_), .Y(new_n13355_));
  OAI21X1  g13291(.A0(new_n13104_), .A1(new_n5096_), .B0(new_n13355_), .Y(new_n13356_));
  AOI21X1  g13292(.A0(new_n13103_), .A1(new_n4637_), .B0(new_n13356_), .Y(new_n13357_));
  XOR2X1   g13293(.A(new_n13357_), .B(\a[8] ), .Y(new_n13358_));
  INVX1    g13294(.A(new_n13311_), .Y(new_n13359_));
  XOR2X1   g13295(.A(new_n13359_), .B(new_n13309_), .Y(new_n13360_));
  OR2X1    g13296(.A(new_n13360_), .B(new_n13358_), .Y(new_n13361_));
  XOR2X1   g13297(.A(new_n13360_), .B(new_n13358_), .Y(new_n13362_));
  INVX1    g13298(.A(new_n13362_), .Y(new_n13363_));
  XOR2X1   g13299(.A(new_n13307_), .B(new_n13147_), .Y(new_n13364_));
  INVX1    g13300(.A(new_n13364_), .Y(new_n13365_));
  INVX1    g13301(.A(new_n12093_), .Y(new_n13366_));
  OAI22X1  g13302(.A0(new_n13090_), .A1(new_n4634_), .B0(new_n13366_), .B1(new_n4869_), .Y(new_n13367_));
  AOI21X1  g13303(.A0(new_n12090_), .A1(new_n5097_), .B0(new_n13367_), .Y(new_n13368_));
  OAI21X1  g13304(.A0(new_n13116_), .A1(new_n4868_), .B0(new_n13368_), .Y(new_n13369_));
  XOR2X1   g13305(.A(new_n13369_), .B(new_n2995_), .Y(new_n13370_));
  NOR2X1   g13306(.A(new_n13370_), .B(new_n13365_), .Y(new_n13371_));
  AND2X1   g13307(.A(new_n13305_), .B(new_n13163_), .Y(new_n13372_));
  XOR2X1   g13308(.A(new_n13372_), .B(new_n13156_), .Y(new_n13373_));
  OAI22X1  g13309(.A0(new_n12839_), .A1(new_n4634_), .B0(new_n13090_), .B1(new_n4869_), .Y(new_n13374_));
  AOI21X1  g13310(.A0(new_n12093_), .A1(new_n5097_), .B0(new_n13374_), .Y(new_n13375_));
  OAI21X1  g13311(.A0(new_n13094_), .A1(new_n4868_), .B0(new_n13375_), .Y(new_n13376_));
  XOR2X1   g13312(.A(new_n13376_), .B(\a[8] ), .Y(new_n13377_));
  AND2X1   g13313(.A(new_n13377_), .B(new_n13373_), .Y(new_n13378_));
  XOR2X1   g13314(.A(new_n13304_), .B(new_n13165_), .Y(new_n13379_));
  OAI22X1  g13315(.A0(new_n12840_), .A1(new_n4634_), .B0(new_n12839_), .B1(new_n4869_), .Y(new_n13380_));
  AOI21X1  g13316(.A0(new_n12095_), .A1(new_n5097_), .B0(new_n13380_), .Y(new_n13381_));
  OAI21X1  g13317(.A0(new_n12846_), .A1(new_n4868_), .B0(new_n13381_), .Y(new_n13382_));
  XOR2X1   g13318(.A(new_n13382_), .B(new_n2995_), .Y(new_n13383_));
  INVX1    g13319(.A(new_n13383_), .Y(new_n13384_));
  NAND2X1  g13320(.A(new_n13384_), .B(new_n13379_), .Y(new_n13385_));
  AOI22X1  g13321(.A0(new_n12102_), .A1(new_n4635_), .B0(new_n12099_), .B1(new_n4870_), .Y(new_n13386_));
  OAI21X1  g13322(.A0(new_n12839_), .A1(new_n5096_), .B0(new_n13386_), .Y(new_n13387_));
  AOI21X1  g13323(.A0(new_n12855_), .A1(new_n4637_), .B0(new_n13387_), .Y(new_n13388_));
  XOR2X1   g13324(.A(new_n13388_), .B(\a[8] ), .Y(new_n13389_));
  INVX1    g13325(.A(new_n13389_), .Y(new_n13390_));
  XOR2X1   g13326(.A(new_n13303_), .B(new_n13302_), .Y(new_n13391_));
  XOR2X1   g13327(.A(new_n13391_), .B(new_n13389_), .Y(new_n13392_));
  AOI22X1  g13328(.A0(new_n12104_), .A1(new_n4635_), .B0(new_n12102_), .B1(new_n4870_), .Y(new_n13393_));
  OAI21X1  g13329(.A0(new_n12840_), .A1(new_n5096_), .B0(new_n13393_), .Y(new_n13394_));
  AOI21X1  g13330(.A0(new_n12859_), .A1(new_n4637_), .B0(new_n13394_), .Y(new_n13395_));
  XOR2X1   g13331(.A(new_n13395_), .B(\a[8] ), .Y(new_n13396_));
  INVX1    g13332(.A(new_n13301_), .Y(new_n13397_));
  XOR2X1   g13333(.A(new_n13397_), .B(new_n13300_), .Y(new_n13398_));
  NOR2X1   g13334(.A(new_n13398_), .B(new_n13396_), .Y(new_n13399_));
  XOR2X1   g13335(.A(new_n13398_), .B(new_n13396_), .Y(new_n13400_));
  INVX1    g13336(.A(new_n13400_), .Y(new_n13401_));
  AOI22X1  g13337(.A0(new_n12107_), .A1(new_n4635_), .B0(new_n12104_), .B1(new_n4870_), .Y(new_n13402_));
  OAI21X1  g13338(.A0(new_n12306_), .A1(new_n5096_), .B0(new_n13402_), .Y(new_n13403_));
  AOI21X1  g13339(.A0(new_n12305_), .A1(new_n4637_), .B0(new_n13403_), .Y(new_n13404_));
  XOR2X1   g13340(.A(new_n13404_), .B(\a[8] ), .Y(new_n13405_));
  INVX1    g13341(.A(new_n13298_), .Y(new_n13406_));
  XOR2X1   g13342(.A(new_n13406_), .B(new_n13296_), .Y(new_n13407_));
  OR2X1    g13343(.A(new_n13407_), .B(new_n13405_), .Y(new_n13408_));
  XOR2X1   g13344(.A(new_n13407_), .B(new_n13405_), .Y(new_n13409_));
  INVX1    g13345(.A(new_n13409_), .Y(new_n13410_));
  XOR2X1   g13346(.A(new_n13294_), .B(new_n13191_), .Y(new_n13411_));
  INVX1    g13347(.A(new_n13411_), .Y(new_n13412_));
  OAI22X1  g13348(.A0(new_n12111_), .A1(new_n4634_), .B0(new_n12109_), .B1(new_n4869_), .Y(new_n13413_));
  AOI21X1  g13349(.A0(new_n12104_), .A1(new_n5097_), .B0(new_n13413_), .Y(new_n13414_));
  OAI21X1  g13350(.A0(new_n12693_), .A1(new_n4868_), .B0(new_n13414_), .Y(new_n13415_));
  XOR2X1   g13351(.A(new_n13415_), .B(new_n2995_), .Y(new_n13416_));
  NOR2X1   g13352(.A(new_n13416_), .B(new_n13412_), .Y(new_n13417_));
  XOR2X1   g13353(.A(new_n13293_), .B(new_n13199_), .Y(new_n13418_));
  OAI22X1  g13354(.A0(new_n12113_), .A1(new_n4634_), .B0(new_n12111_), .B1(new_n4869_), .Y(new_n13419_));
  AOI21X1  g13355(.A0(new_n12107_), .A1(new_n5097_), .B0(new_n13419_), .Y(new_n13420_));
  OAI21X1  g13356(.A0(new_n12708_), .A1(new_n4868_), .B0(new_n13420_), .Y(new_n13421_));
  XOR2X1   g13357(.A(new_n13421_), .B(\a[8] ), .Y(new_n13422_));
  XOR2X1   g13358(.A(new_n13292_), .B(new_n13209_), .Y(new_n13423_));
  INVX1    g13359(.A(new_n13423_), .Y(new_n13424_));
  OAI22X1  g13360(.A0(new_n12117_), .A1(new_n4634_), .B0(new_n12113_), .B1(new_n4869_), .Y(new_n13425_));
  AOI21X1  g13361(.A0(new_n12208_), .A1(new_n5097_), .B0(new_n13425_), .Y(new_n13426_));
  OAI21X1  g13362(.A0(new_n12685_), .A1(new_n4868_), .B0(new_n13426_), .Y(new_n13427_));
  XOR2X1   g13363(.A(new_n13427_), .B(new_n2995_), .Y(new_n13428_));
  OR2X1    g13364(.A(new_n13428_), .B(new_n13424_), .Y(new_n13429_));
  AOI22X1  g13365(.A0(new_n12133_), .A1(new_n4635_), .B0(new_n12720_), .B1(new_n4870_), .Y(new_n13430_));
  OAI21X1  g13366(.A0(new_n12113_), .A1(new_n5096_), .B0(new_n13430_), .Y(new_n13431_));
  AOI21X1  g13367(.A0(new_n12719_), .A1(new_n4637_), .B0(new_n13431_), .Y(new_n13432_));
  XOR2X1   g13368(.A(new_n13432_), .B(\a[8] ), .Y(new_n13433_));
  INVX1    g13369(.A(new_n13433_), .Y(new_n13434_));
  XOR2X1   g13370(.A(new_n13291_), .B(new_n13290_), .Y(new_n13435_));
  XOR2X1   g13371(.A(new_n13435_), .B(new_n13433_), .Y(new_n13436_));
  AOI22X1  g13372(.A0(new_n12138_), .A1(new_n4635_), .B0(new_n12133_), .B1(new_n4870_), .Y(new_n13437_));
  OAI21X1  g13373(.A0(new_n12117_), .A1(new_n5096_), .B0(new_n13437_), .Y(new_n13438_));
  AOI21X1  g13374(.A0(new_n12526_), .A1(new_n4637_), .B0(new_n13438_), .Y(new_n13439_));
  XOR2X1   g13375(.A(new_n13439_), .B(\a[8] ), .Y(new_n13440_));
  INVX1    g13376(.A(new_n13289_), .Y(new_n13441_));
  XOR2X1   g13377(.A(new_n13441_), .B(new_n13288_), .Y(new_n13442_));
  OR2X1    g13378(.A(new_n13442_), .B(new_n13440_), .Y(new_n13443_));
  XOR2X1   g13379(.A(new_n13442_), .B(new_n13440_), .Y(new_n13444_));
  INVX1    g13380(.A(new_n13444_), .Y(new_n13445_));
  AOI22X1  g13381(.A0(new_n12141_), .A1(new_n4635_), .B0(new_n12138_), .B1(new_n4870_), .Y(new_n13446_));
  OAI21X1  g13382(.A0(new_n12134_), .A1(new_n5096_), .B0(new_n13446_), .Y(new_n13447_));
  AOI21X1  g13383(.A0(new_n12536_), .A1(new_n4637_), .B0(new_n13447_), .Y(new_n13448_));
  XOR2X1   g13384(.A(new_n13448_), .B(\a[8] ), .Y(new_n13449_));
  AND2X1   g13385(.A(new_n13285_), .B(new_n13237_), .Y(new_n13450_));
  INVX1    g13386(.A(new_n13286_), .Y(new_n13451_));
  XOR2X1   g13387(.A(new_n13451_), .B(new_n13450_), .Y(new_n13452_));
  OR2X1    g13388(.A(new_n13452_), .B(new_n13449_), .Y(new_n13453_));
  XOR2X1   g13389(.A(new_n13452_), .B(new_n13449_), .Y(new_n13454_));
  INVX1    g13390(.A(new_n13454_), .Y(new_n13455_));
  INVX1    g13391(.A(new_n13238_), .Y(new_n13456_));
  XOR2X1   g13392(.A(new_n13284_), .B(new_n13456_), .Y(new_n13457_));
  AOI22X1  g13393(.A0(new_n12144_), .A1(new_n4635_), .B0(new_n12141_), .B1(new_n4870_), .Y(new_n13458_));
  OAI21X1  g13394(.A0(new_n12314_), .A1(new_n5096_), .B0(new_n13458_), .Y(new_n13459_));
  AOI21X1  g13395(.A0(new_n12313_), .A1(new_n4637_), .B0(new_n13459_), .Y(new_n13460_));
  XOR2X1   g13396(.A(new_n13460_), .B(\a[8] ), .Y(new_n13461_));
  NOR2X1   g13397(.A(new_n13461_), .B(new_n13457_), .Y(new_n13462_));
  XOR2X1   g13398(.A(new_n13283_), .B(new_n13282_), .Y(new_n13463_));
  INVX1    g13399(.A(new_n13463_), .Y(new_n13464_));
  OAI22X1  g13400(.A0(new_n12186_), .A1(new_n4634_), .B0(new_n12192_), .B1(new_n4869_), .Y(new_n13465_));
  AOI21X1  g13401(.A0(new_n12141_), .A1(new_n5097_), .B0(new_n13465_), .Y(new_n13466_));
  OAI21X1  g13402(.A0(new_n12444_), .A1(new_n4868_), .B0(new_n13466_), .Y(new_n13467_));
  XOR2X1   g13403(.A(new_n13467_), .B(new_n2995_), .Y(new_n13468_));
  OR2X1    g13404(.A(new_n13468_), .B(new_n13464_), .Y(new_n13469_));
  XOR2X1   g13405(.A(new_n13280_), .B(new_n13255_), .Y(new_n13470_));
  INVX1    g13406(.A(new_n13470_), .Y(new_n13471_));
  OAI22X1  g13407(.A0(new_n12322_), .A1(new_n4634_), .B0(new_n12186_), .B1(new_n4869_), .Y(new_n13472_));
  AOI21X1  g13408(.A0(new_n12144_), .A1(new_n5097_), .B0(new_n13472_), .Y(new_n13473_));
  OAI21X1  g13409(.A0(new_n12453_), .A1(new_n4868_), .B0(new_n13473_), .Y(new_n13474_));
  XOR2X1   g13410(.A(new_n13474_), .B(new_n2995_), .Y(new_n13475_));
  NOR2X1   g13411(.A(new_n13475_), .B(new_n13471_), .Y(new_n13476_));
  AOI22X1  g13412(.A0(new_n12155_), .A1(new_n4635_), .B0(new_n12151_), .B1(new_n4870_), .Y(new_n13477_));
  OAI21X1  g13413(.A0(new_n12186_), .A1(new_n5096_), .B0(new_n13477_), .Y(new_n13478_));
  AOI21X1  g13414(.A0(new_n12430_), .A1(new_n4637_), .B0(new_n13478_), .Y(new_n13479_));
  XOR2X1   g13415(.A(new_n13479_), .B(\a[8] ), .Y(new_n13480_));
  INVX1    g13416(.A(new_n13480_), .Y(new_n13481_));
  XOR2X1   g13417(.A(new_n13279_), .B(new_n13278_), .Y(new_n13482_));
  NAND2X1  g13418(.A(new_n13482_), .B(new_n13481_), .Y(new_n13483_));
  XOR2X1   g13419(.A(new_n13482_), .B(new_n13480_), .Y(new_n13484_));
  XOR2X1   g13420(.A(new_n13276_), .B(new_n2911_), .Y(new_n13485_));
  XOR2X1   g13421(.A(new_n13485_), .B(new_n13273_), .Y(new_n13486_));
  AOI22X1  g13422(.A0(new_n12158_), .A1(new_n4635_), .B0(new_n12155_), .B1(new_n4870_), .Y(new_n13487_));
  OAI21X1  g13423(.A0(new_n12322_), .A1(new_n5096_), .B0(new_n13487_), .Y(new_n13488_));
  AOI21X1  g13424(.A0(new_n12321_), .A1(new_n4637_), .B0(new_n13488_), .Y(new_n13489_));
  XOR2X1   g13425(.A(new_n13489_), .B(\a[8] ), .Y(new_n13490_));
  NOR2X1   g13426(.A(new_n13490_), .B(new_n13486_), .Y(new_n13491_));
  AOI22X1  g13427(.A0(new_n12162_), .A1(new_n4635_), .B0(new_n12158_), .B1(new_n4870_), .Y(new_n13492_));
  OAI21X1  g13428(.A0(new_n12353_), .A1(new_n5096_), .B0(new_n13492_), .Y(new_n13493_));
  AOI21X1  g13429(.A0(new_n12352_), .A1(new_n4637_), .B0(new_n13493_), .Y(new_n13494_));
  XOR2X1   g13430(.A(new_n13494_), .B(\a[8] ), .Y(new_n13495_));
  INVX1    g13431(.A(new_n13495_), .Y(new_n13496_));
  NOR3X1   g13432(.A(new_n13266_), .B(new_n13265_), .C(new_n2911_), .Y(new_n13497_));
  XOR2X1   g13433(.A(new_n13269_), .B(\a[11] ), .Y(new_n13498_));
  XOR2X1   g13434(.A(new_n13498_), .B(new_n13497_), .Y(new_n13499_));
  NAND2X1  g13435(.A(new_n13499_), .B(new_n13496_), .Y(new_n13500_));
  XOR2X1   g13436(.A(new_n13499_), .B(new_n13495_), .Y(new_n13501_));
  NOR2X1   g13437(.A(new_n13266_), .B(new_n2911_), .Y(new_n13502_));
  XOR2X1   g13438(.A(new_n13502_), .B(new_n13265_), .Y(new_n13503_));
  OAI22X1  g13439(.A0(new_n12168_), .A1(new_n4634_), .B0(new_n12329_), .B1(new_n4869_), .Y(new_n13504_));
  AOI21X1  g13440(.A0(new_n12158_), .A1(new_n5097_), .B0(new_n13504_), .Y(new_n13505_));
  OAI21X1  g13441(.A0(new_n12368_), .A1(new_n4868_), .B0(new_n13505_), .Y(new_n13506_));
  XOR2X1   g13442(.A(new_n13506_), .B(new_n2995_), .Y(new_n13507_));
  NOR2X1   g13443(.A(new_n13507_), .B(new_n13503_), .Y(new_n13508_));
  OAI22X1  g13444(.A0(new_n12176_), .A1(new_n4869_), .B0(new_n12170_), .B1(new_n5096_), .Y(new_n13509_));
  AOI21X1  g13445(.A0(new_n12337_), .A1(new_n4637_), .B0(new_n13509_), .Y(new_n13510_));
  XOR2X1   g13446(.A(new_n13510_), .B(\a[8] ), .Y(new_n13511_));
  AOI21X1  g13447(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n4630_), .Y(new_n13512_));
  OAI22X1  g13448(.A0(new_n12176_), .A1(new_n4634_), .B0(new_n12170_), .B1(new_n4869_), .Y(new_n13513_));
  AOI21X1  g13449(.A0(new_n12165_), .A1(new_n5097_), .B0(new_n13513_), .Y(new_n13514_));
  OAI21X1  g13450(.A0(new_n12344_), .A1(new_n4868_), .B0(new_n13514_), .Y(new_n13515_));
  NOR4X1   g13451(.A(new_n13515_), .B(new_n13512_), .C(new_n13511_), .D(new_n2995_), .Y(new_n13516_));
  NAND2X1  g13452(.A(new_n13516_), .B(new_n13266_), .Y(new_n13517_));
  INVX1    g13453(.A(new_n13516_), .Y(new_n13518_));
  XOR2X1   g13454(.A(new_n13518_), .B(new_n13266_), .Y(new_n13519_));
  AOI22X1  g13455(.A0(new_n12331_), .A1(new_n4635_), .B0(new_n12165_), .B1(new_n4870_), .Y(new_n13520_));
  OAI21X1  g13456(.A0(new_n12329_), .A1(new_n5096_), .B0(new_n13520_), .Y(new_n13521_));
  AOI21X1  g13457(.A0(new_n12328_), .A1(new_n4637_), .B0(new_n13521_), .Y(new_n13522_));
  XOR2X1   g13458(.A(new_n13522_), .B(\a[8] ), .Y(new_n13523_));
  OAI21X1  g13459(.A0(new_n13523_), .A1(new_n13519_), .B0(new_n13517_), .Y(new_n13524_));
  XOR2X1   g13460(.A(new_n13507_), .B(new_n13503_), .Y(new_n13525_));
  AOI21X1  g13461(.A0(new_n13525_), .A1(new_n13524_), .B0(new_n13508_), .Y(new_n13526_));
  OAI21X1  g13462(.A0(new_n13526_), .A1(new_n13501_), .B0(new_n13500_), .Y(new_n13527_));
  XOR2X1   g13463(.A(new_n13490_), .B(new_n13486_), .Y(new_n13528_));
  AOI21X1  g13464(.A0(new_n13528_), .A1(new_n13527_), .B0(new_n13491_), .Y(new_n13529_));
  OR2X1    g13465(.A(new_n13529_), .B(new_n13484_), .Y(new_n13530_));
  XOR2X1   g13466(.A(new_n13475_), .B(new_n13470_), .Y(new_n13531_));
  AOI21X1  g13467(.A0(new_n13530_), .A1(new_n13483_), .B0(new_n13531_), .Y(new_n13532_));
  NOR2X1   g13468(.A(new_n13532_), .B(new_n13476_), .Y(new_n13533_));
  XOR2X1   g13469(.A(new_n13468_), .B(new_n13463_), .Y(new_n13534_));
  OAI21X1  g13470(.A0(new_n13534_), .A1(new_n13533_), .B0(new_n13469_), .Y(new_n13535_));
  XOR2X1   g13471(.A(new_n13461_), .B(new_n13457_), .Y(new_n13536_));
  AOI21X1  g13472(.A0(new_n13536_), .A1(new_n13535_), .B0(new_n13462_), .Y(new_n13537_));
  OR2X1    g13473(.A(new_n13537_), .B(new_n13455_), .Y(new_n13538_));
  AND2X1   g13474(.A(new_n13538_), .B(new_n13453_), .Y(new_n13539_));
  OR2X1    g13475(.A(new_n13539_), .B(new_n13445_), .Y(new_n13540_));
  AND2X1   g13476(.A(new_n13540_), .B(new_n13443_), .Y(new_n13541_));
  NOR2X1   g13477(.A(new_n13541_), .B(new_n13436_), .Y(new_n13542_));
  AOI21X1  g13478(.A0(new_n13435_), .A1(new_n13434_), .B0(new_n13542_), .Y(new_n13543_));
  XOR2X1   g13479(.A(new_n13428_), .B(new_n13423_), .Y(new_n13544_));
  OR2X1    g13480(.A(new_n13544_), .B(new_n13543_), .Y(new_n13545_));
  XOR2X1   g13481(.A(new_n13421_), .B(new_n2995_), .Y(new_n13546_));
  XOR2X1   g13482(.A(new_n13546_), .B(new_n13418_), .Y(new_n13547_));
  AOI21X1  g13483(.A0(new_n13545_), .A1(new_n13429_), .B0(new_n13547_), .Y(new_n13548_));
  AOI21X1  g13484(.A0(new_n13422_), .A1(new_n13418_), .B0(new_n13548_), .Y(new_n13549_));
  INVX1    g13485(.A(new_n13549_), .Y(new_n13550_));
  XOR2X1   g13486(.A(new_n13416_), .B(new_n13412_), .Y(new_n13551_));
  AOI21X1  g13487(.A0(new_n13551_), .A1(new_n13550_), .B0(new_n13417_), .Y(new_n13552_));
  OR2X1    g13488(.A(new_n13552_), .B(new_n13410_), .Y(new_n13553_));
  AOI21X1  g13489(.A0(new_n13553_), .A1(new_n13408_), .B0(new_n13401_), .Y(new_n13554_));
  NOR2X1   g13490(.A(new_n13554_), .B(new_n13399_), .Y(new_n13555_));
  NOR2X1   g13491(.A(new_n13555_), .B(new_n13392_), .Y(new_n13556_));
  AOI21X1  g13492(.A0(new_n13391_), .A1(new_n13390_), .B0(new_n13556_), .Y(new_n13557_));
  XOR2X1   g13493(.A(new_n13383_), .B(new_n13379_), .Y(new_n13558_));
  OAI21X1  g13494(.A0(new_n13558_), .A1(new_n13557_), .B0(new_n13385_), .Y(new_n13559_));
  XOR2X1   g13495(.A(new_n13376_), .B(new_n2995_), .Y(new_n13560_));
  XOR2X1   g13496(.A(new_n13560_), .B(new_n13373_), .Y(new_n13561_));
  INVX1    g13497(.A(new_n13561_), .Y(new_n13562_));
  AOI21X1  g13498(.A0(new_n13562_), .A1(new_n13559_), .B0(new_n13378_), .Y(new_n13563_));
  INVX1    g13499(.A(new_n13563_), .Y(new_n13564_));
  XOR2X1   g13500(.A(new_n13370_), .B(new_n13365_), .Y(new_n13565_));
  AOI21X1  g13501(.A0(new_n13565_), .A1(new_n13564_), .B0(new_n13371_), .Y(new_n13566_));
  OR2X1    g13502(.A(new_n13566_), .B(new_n13363_), .Y(new_n13567_));
  AOI21X1  g13503(.A0(new_n13567_), .A1(new_n13361_), .B0(new_n13354_), .Y(new_n13568_));
  AOI21X1  g13504(.A0(new_n13353_), .A1(new_n13352_), .B0(new_n13568_), .Y(new_n13569_));
  XOR2X1   g13505(.A(new_n13347_), .B(new_n13339_), .Y(new_n13570_));
  OR2X1    g13506(.A(new_n13570_), .B(new_n13569_), .Y(new_n13571_));
  OAI21X1  g13507(.A0(new_n13347_), .A1(new_n13340_), .B0(new_n13571_), .Y(new_n13572_));
  XOR2X1   g13508(.A(new_n13336_), .B(new_n2995_), .Y(new_n13573_));
  XOR2X1   g13509(.A(new_n13573_), .B(new_n13328_), .Y(new_n13574_));
  INVX1    g13510(.A(new_n13574_), .Y(new_n13575_));
  AOI21X1  g13511(.A0(new_n13575_), .A1(new_n13572_), .B0(new_n13338_), .Y(new_n13576_));
  XOR2X1   g13512(.A(new_n13327_), .B(new_n13318_), .Y(new_n13577_));
  OR2X1    g13513(.A(new_n13577_), .B(new_n13576_), .Y(new_n13578_));
  OAI21X1  g13514(.A0(new_n13327_), .A1(new_n13319_), .B0(new_n13578_), .Y(new_n13579_));
  AOI22X1  g13515(.A0(new_n12088_), .A1(new_n4078_), .B0(new_n12085_), .B1(new_n4247_), .Y(new_n13580_));
  OAI21X1  g13516(.A0(new_n13321_), .A1(new_n4427_), .B0(new_n13580_), .Y(new_n13581_));
  AOI21X1  g13517(.A0(new_n13344_), .A1(new_n4080_), .B0(new_n13581_), .Y(new_n13582_));
  XOR2X1   g13518(.A(new_n13582_), .B(\a[11] ), .Y(new_n13583_));
  XOR2X1   g13519(.A(new_n13095_), .B(\a[14] ), .Y(new_n13584_));
  AND2X1   g13520(.A(new_n13584_), .B(new_n13089_), .Y(new_n13585_));
  INVX1    g13521(.A(new_n13585_), .Y(new_n13586_));
  OAI21X1  g13522(.A0(new_n13025_), .A1(new_n12849_), .B0(new_n13098_), .Y(new_n13587_));
  AND2X1   g13523(.A(new_n13587_), .B(new_n13586_), .Y(new_n13588_));
  AOI22X1  g13524(.A0(new_n12102_), .A1(new_n3232_), .B0(new_n12099_), .B1(new_n3390_), .Y(new_n13589_));
  OAI21X1  g13525(.A0(new_n12839_), .A1(new_n3545_), .B0(new_n13589_), .Y(new_n13590_));
  AOI21X1  g13526(.A0(new_n12855_), .A1(new_n3234_), .B0(new_n13590_), .Y(new_n13591_));
  XOR2X1   g13527(.A(new_n13591_), .B(\a[17] ), .Y(new_n13592_));
  INVX1    g13528(.A(new_n13077_), .Y(new_n13593_));
  NOR2X1   g13529(.A(new_n13081_), .B(new_n13593_), .Y(new_n13594_));
  INVX1    g13530(.A(new_n13594_), .Y(new_n13595_));
  OAI21X1  g13531(.A0(new_n13082_), .A1(new_n13033_), .B0(new_n13595_), .Y(new_n13596_));
  AOI22X1  g13532(.A0(new_n12133_), .A1(new_n2657_), .B0(new_n12720_), .B1(new_n2696_), .Y(new_n13597_));
  OAI21X1  g13533(.A0(new_n12113_), .A1(new_n2753_), .B0(new_n13597_), .Y(new_n13598_));
  AOI21X1  g13534(.A0(new_n12719_), .A1(new_n2658_), .B0(new_n13598_), .Y(new_n13599_));
  XOR2X1   g13535(.A(new_n13599_), .B(\a[23] ), .Y(new_n13600_));
  INVX1    g13536(.A(new_n13042_), .Y(new_n13601_));
  INVX1    g13537(.A(new_n13066_), .Y(new_n13602_));
  NOR2X1   g13538(.A(new_n13070_), .B(new_n13602_), .Y(new_n13603_));
  INVX1    g13539(.A(new_n13603_), .Y(new_n13604_));
  OAI21X1  g13540(.A0(new_n13071_), .A1(new_n13601_), .B0(new_n13604_), .Y(new_n13605_));
  INVX1    g13541(.A(new_n13605_), .Y(new_n13606_));
  AOI22X1  g13542(.A0(new_n12155_), .A1(new_n2185_), .B0(new_n12151_), .B1(new_n2095_), .Y(new_n13607_));
  OAI21X1  g13543(.A0(new_n12186_), .A1(new_n2140_), .B0(new_n13607_), .Y(new_n13608_));
  AOI21X1  g13544(.A0(new_n12430_), .A1(new_n2062_), .B0(new_n13608_), .Y(new_n13609_));
  XOR2X1   g13545(.A(new_n13609_), .B(\a[29] ), .Y(new_n13610_));
  NOR2X1   g13546(.A(new_n13060_), .B(new_n13056_), .Y(new_n13611_));
  XOR2X1   g13547(.A(new_n13060_), .B(new_n13056_), .Y(new_n13612_));
  AOI21X1  g13548(.A0(new_n13612_), .A1(new_n13049_), .B0(new_n13611_), .Y(new_n13613_));
  NOR3X1   g13549(.A(new_n497_), .B(new_n455_), .C(new_n1284_), .Y(new_n13614_));
  NOR3X1   g13550(.A(new_n249_), .B(new_n124_), .C(new_n114_), .Y(new_n13615_));
  NOR4X1   g13551(.A(new_n547_), .B(new_n419_), .C(new_n998_), .D(new_n149_), .Y(new_n13616_));
  NAND3X1  g13552(.A(new_n13616_), .B(new_n13615_), .C(new_n13614_), .Y(new_n13617_));
  OR4X1    g13553(.A(new_n668_), .B(new_n1316_), .C(new_n395_), .D(new_n247_), .Y(new_n13618_));
  NOR4X1   g13554(.A(new_n13618_), .B(new_n13617_), .C(new_n236_), .D(new_n186_), .Y(new_n13619_));
  NAND3X1  g13555(.A(new_n13619_), .B(new_n12029_), .C(new_n8673_), .Y(new_n13620_));
  AOI22X1  g13556(.A0(new_n12165_), .A1(new_n1890_), .B0(new_n12162_), .B1(new_n1884_), .Y(new_n13621_));
  OAI21X1  g13557(.A0(new_n12396_), .A1(new_n3498_), .B0(new_n13621_), .Y(new_n13622_));
  AOI21X1  g13558(.A0(new_n12395_), .A1(new_n407_), .B0(new_n13622_), .Y(new_n13623_));
  XOR2X1   g13559(.A(new_n13623_), .B(new_n13620_), .Y(new_n13624_));
  INVX1    g13560(.A(new_n13624_), .Y(new_n13625_));
  XOR2X1   g13561(.A(new_n13625_), .B(new_n13613_), .Y(new_n13626_));
  XOR2X1   g13562(.A(new_n13626_), .B(new_n13610_), .Y(new_n13627_));
  INVX1    g13563(.A(new_n13627_), .Y(new_n13628_));
  NOR2X1   g13564(.A(new_n13062_), .B(new_n13046_), .Y(new_n13629_));
  AOI21X1  g13565(.A0(new_n13065_), .A1(new_n13063_), .B0(new_n13629_), .Y(new_n13630_));
  XOR2X1   g13566(.A(new_n13630_), .B(new_n13628_), .Y(new_n13631_));
  AOI22X1  g13567(.A0(new_n12144_), .A1(new_n2424_), .B0(new_n12141_), .B1(new_n2418_), .Y(new_n13632_));
  OAI21X1  g13568(.A0(new_n12314_), .A1(new_n2626_), .B0(new_n13632_), .Y(new_n13633_));
  AOI21X1  g13569(.A0(new_n12313_), .A1(new_n2301_), .B0(new_n13633_), .Y(new_n13634_));
  XOR2X1   g13570(.A(new_n13634_), .B(\a[26] ), .Y(new_n13635_));
  XOR2X1   g13571(.A(new_n13635_), .B(new_n13631_), .Y(new_n13636_));
  XOR2X1   g13572(.A(new_n13636_), .B(new_n13606_), .Y(new_n13637_));
  XOR2X1   g13573(.A(new_n13637_), .B(new_n13600_), .Y(new_n13638_));
  OR2X1    g13574(.A(new_n13072_), .B(new_n13037_), .Y(new_n13639_));
  OR2X1    g13575(.A(new_n13076_), .B(new_n13074_), .Y(new_n13640_));
  AND2X1   g13576(.A(new_n13640_), .B(new_n13639_), .Y(new_n13641_));
  XOR2X1   g13577(.A(new_n13641_), .B(new_n13638_), .Y(new_n13642_));
  OAI22X1  g13578(.A0(new_n12111_), .A1(new_n3250_), .B0(new_n12109_), .B1(new_n3144_), .Y(new_n13643_));
  AOI21X1  g13579(.A0(new_n12104_), .A1(new_n3146_), .B0(new_n13643_), .Y(new_n13644_));
  OAI21X1  g13580(.A0(new_n12693_), .A1(new_n3098_), .B0(new_n13644_), .Y(new_n13645_));
  XOR2X1   g13581(.A(new_n13645_), .B(new_n1920_), .Y(new_n13646_));
  XOR2X1   g13582(.A(new_n13646_), .B(new_n13642_), .Y(new_n13647_));
  XOR2X1   g13583(.A(new_n13647_), .B(new_n13596_), .Y(new_n13648_));
  XOR2X1   g13584(.A(new_n13648_), .B(new_n13592_), .Y(new_n13649_));
  OR2X1    g13585(.A(new_n13084_), .B(new_n13030_), .Y(new_n13650_));
  OAI21X1  g13586(.A0(new_n13088_), .A1(new_n13086_), .B0(new_n13650_), .Y(new_n13651_));
  XOR2X1   g13587(.A(new_n13651_), .B(new_n13649_), .Y(new_n13652_));
  OAI22X1  g13588(.A0(new_n13090_), .A1(new_n3627_), .B0(new_n13366_), .B1(new_n3907_), .Y(new_n13653_));
  AOI21X1  g13589(.A0(new_n12090_), .A1(new_n3984_), .B0(new_n13653_), .Y(new_n13654_));
  OAI21X1  g13590(.A0(new_n13116_), .A1(new_n3906_), .B0(new_n13654_), .Y(new_n13655_));
  XOR2X1   g13591(.A(new_n13655_), .B(new_n2529_), .Y(new_n13656_));
  XOR2X1   g13592(.A(new_n13656_), .B(new_n13652_), .Y(new_n13657_));
  INVX1    g13593(.A(new_n13657_), .Y(new_n13658_));
  XOR2X1   g13594(.A(new_n13658_), .B(new_n13588_), .Y(new_n13659_));
  XOR2X1   g13595(.A(new_n13659_), .B(new_n13583_), .Y(new_n13660_));
  INVX1    g13596(.A(new_n13660_), .Y(new_n13661_));
  NOR2X1   g13597(.A(new_n13099_), .B(new_n12302_), .Y(new_n13662_));
  AOI21X1  g13598(.A0(new_n13317_), .A1(new_n13100_), .B0(new_n13662_), .Y(new_n13663_));
  XOR2X1   g13599(.A(new_n13663_), .B(new_n13661_), .Y(new_n13664_));
  INVX1    g13600(.A(new_n12079_), .Y(new_n13665_));
  OAI22X1  g13601(.A0(new_n13320_), .A1(new_n4634_), .B0(new_n13665_), .B1(new_n4869_), .Y(new_n13666_));
  AOI21X1  g13602(.A0(new_n12076_), .A1(new_n5097_), .B0(new_n13666_), .Y(new_n13667_));
  NOR2X1   g13603(.A(new_n12079_), .B(new_n12076_), .Y(new_n13668_));
  OAI21X1  g13604(.A0(new_n13668_), .A1(new_n12080_), .B0(new_n12237_), .Y(new_n13669_));
  NOR3X1   g13605(.A(new_n13668_), .B(new_n12237_), .C(new_n12080_), .Y(new_n13670_));
  INVX1    g13606(.A(new_n13670_), .Y(new_n13671_));
  AND2X1   g13607(.A(new_n13671_), .B(new_n13669_), .Y(new_n13672_));
  OAI21X1  g13608(.A0(new_n13672_), .A1(new_n4868_), .B0(new_n13667_), .Y(new_n13673_));
  XOR2X1   g13609(.A(new_n13673_), .B(new_n2995_), .Y(new_n13674_));
  XOR2X1   g13610(.A(new_n13674_), .B(new_n13664_), .Y(new_n13675_));
  XOR2X1   g13611(.A(new_n13675_), .B(new_n13579_), .Y(new_n13676_));
  XOR2X1   g13612(.A(new_n13676_), .B(new_n12296_), .Y(new_n13677_));
  XOR2X1   g13613(.A(new_n12242_), .B(new_n12241_), .Y(new_n13678_));
  INVX1    g13614(.A(new_n12074_), .Y(new_n13679_));
  AOI22X1  g13615(.A0(new_n12076_), .A1(new_n5373_), .B0(new_n12018_), .B1(new_n5659_), .Y(new_n13680_));
  OAI21X1  g13616(.A0(new_n13679_), .A1(new_n5959_), .B0(new_n13680_), .Y(new_n13681_));
  AOI21X1  g13617(.A0(new_n13678_), .A1(new_n67_), .B0(new_n13681_), .Y(new_n13682_));
  XOR2X1   g13618(.A(new_n13682_), .B(\a[5] ), .Y(new_n13683_));
  INVX1    g13619(.A(new_n13577_), .Y(new_n13684_));
  XOR2X1   g13620(.A(new_n13684_), .B(new_n13576_), .Y(new_n13685_));
  NOR2X1   g13621(.A(new_n13685_), .B(new_n13683_), .Y(new_n13686_));
  XOR2X1   g13622(.A(new_n13685_), .B(new_n13683_), .Y(new_n13687_));
  XOR2X1   g13623(.A(new_n12076_), .B(new_n12018_), .Y(new_n13688_));
  OR2X1    g13624(.A(new_n13688_), .B(new_n12239_), .Y(new_n13689_));
  OAI21X1  g13625(.A0(new_n12241_), .A1(new_n12240_), .B0(new_n13689_), .Y(new_n13690_));
  INVX1    g13626(.A(new_n12018_), .Y(new_n13691_));
  AOI22X1  g13627(.A0(new_n12079_), .A1(new_n5373_), .B0(new_n12076_), .B1(new_n5659_), .Y(new_n13692_));
  OAI21X1  g13628(.A0(new_n13691_), .A1(new_n5959_), .B0(new_n13692_), .Y(new_n13693_));
  AOI21X1  g13629(.A0(new_n13690_), .A1(new_n67_), .B0(new_n13693_), .Y(new_n13694_));
  XOR2X1   g13630(.A(new_n13694_), .B(\a[5] ), .Y(new_n13695_));
  XOR2X1   g13631(.A(new_n13574_), .B(new_n13572_), .Y(new_n13696_));
  XOR2X1   g13632(.A(new_n13696_), .B(new_n13695_), .Y(new_n13697_));
  INVX1    g13633(.A(new_n13697_), .Y(new_n13698_));
  INVX1    g13634(.A(new_n13672_), .Y(new_n13699_));
  INVX1    g13635(.A(new_n12076_), .Y(new_n13700_));
  AOI22X1  g13636(.A0(new_n12081_), .A1(new_n5373_), .B0(new_n12079_), .B1(new_n5659_), .Y(new_n13701_));
  OAI21X1  g13637(.A0(new_n13700_), .A1(new_n5959_), .B0(new_n13701_), .Y(new_n13702_));
  AOI21X1  g13638(.A0(new_n13699_), .A1(new_n67_), .B0(new_n13702_), .Y(new_n13703_));
  XOR2X1   g13639(.A(new_n13703_), .B(\a[5] ), .Y(new_n13704_));
  INVX1    g13640(.A(new_n13570_), .Y(new_n13705_));
  XOR2X1   g13641(.A(new_n13705_), .B(new_n13569_), .Y(new_n13706_));
  NOR2X1   g13642(.A(new_n13706_), .B(new_n13704_), .Y(new_n13707_));
  XOR2X1   g13643(.A(new_n13706_), .B(new_n13704_), .Y(new_n13708_));
  INVX1    g13644(.A(new_n13354_), .Y(new_n13709_));
  AND2X1   g13645(.A(new_n13567_), .B(new_n13361_), .Y(new_n13710_));
  XOR2X1   g13646(.A(new_n13710_), .B(new_n13709_), .Y(new_n13711_));
  OAI22X1  g13647(.A0(new_n13321_), .A1(new_n5372_), .B0(new_n13320_), .B1(new_n5658_), .Y(new_n13712_));
  AOI21X1  g13648(.A0(new_n12079_), .A1(new_n5960_), .B0(new_n13712_), .Y(new_n13713_));
  OAI21X1  g13649(.A0(new_n13325_), .A1(new_n5657_), .B0(new_n13713_), .Y(new_n13714_));
  XOR2X1   g13650(.A(new_n13714_), .B(new_n3289_), .Y(new_n13715_));
  XOR2X1   g13651(.A(new_n13566_), .B(new_n13363_), .Y(new_n13716_));
  OAI22X1  g13652(.A0(new_n12298_), .A1(new_n5372_), .B0(new_n13321_), .B1(new_n5658_), .Y(new_n13717_));
  AOI21X1  g13653(.A0(new_n12081_), .A1(new_n5960_), .B0(new_n13717_), .Y(new_n13718_));
  OAI21X1  g13654(.A0(new_n13335_), .A1(new_n5657_), .B0(new_n13718_), .Y(new_n13719_));
  XOR2X1   g13655(.A(new_n13719_), .B(\a[5] ), .Y(new_n13720_));
  AND2X1   g13656(.A(new_n13720_), .B(new_n13716_), .Y(new_n13721_));
  AOI22X1  g13657(.A0(new_n12088_), .A1(new_n5373_), .B0(new_n12085_), .B1(new_n5659_), .Y(new_n13722_));
  OAI21X1  g13658(.A0(new_n13321_), .A1(new_n5959_), .B0(new_n13722_), .Y(new_n13723_));
  AOI21X1  g13659(.A0(new_n13344_), .A1(new_n67_), .B0(new_n13723_), .Y(new_n13724_));
  XOR2X1   g13660(.A(new_n13724_), .B(\a[5] ), .Y(new_n13725_));
  XOR2X1   g13661(.A(new_n13565_), .B(new_n13563_), .Y(new_n13726_));
  INVX1    g13662(.A(new_n13725_), .Y(new_n13727_));
  XOR2X1   g13663(.A(new_n13726_), .B(new_n13727_), .Y(new_n13728_));
  AOI22X1  g13664(.A0(new_n12090_), .A1(new_n5373_), .B0(new_n12088_), .B1(new_n5659_), .Y(new_n13729_));
  OAI21X1  g13665(.A0(new_n12298_), .A1(new_n5959_), .B0(new_n13729_), .Y(new_n13730_));
  AOI21X1  g13666(.A0(new_n12297_), .A1(new_n67_), .B0(new_n13730_), .Y(new_n13731_));
  XOR2X1   g13667(.A(new_n13731_), .B(\a[5] ), .Y(new_n13732_));
  XOR2X1   g13668(.A(new_n13561_), .B(new_n13559_), .Y(new_n13733_));
  NOR2X1   g13669(.A(new_n13733_), .B(new_n13732_), .Y(new_n13734_));
  XOR2X1   g13670(.A(new_n13733_), .B(new_n13732_), .Y(new_n13735_));
  AOI22X1  g13671(.A0(new_n12093_), .A1(new_n5373_), .B0(new_n12090_), .B1(new_n5659_), .Y(new_n13736_));
  OAI21X1  g13672(.A0(new_n13104_), .A1(new_n5959_), .B0(new_n13736_), .Y(new_n13737_));
  AOI21X1  g13673(.A0(new_n13103_), .A1(new_n67_), .B0(new_n13737_), .Y(new_n13738_));
  XOR2X1   g13674(.A(new_n13738_), .B(\a[5] ), .Y(new_n13739_));
  INVX1    g13675(.A(new_n13558_), .Y(new_n13740_));
  XOR2X1   g13676(.A(new_n13740_), .B(new_n13557_), .Y(new_n13741_));
  OR2X1    g13677(.A(new_n13741_), .B(new_n13739_), .Y(new_n13742_));
  XOR2X1   g13678(.A(new_n13741_), .B(new_n13739_), .Y(new_n13743_));
  INVX1    g13679(.A(new_n13743_), .Y(new_n13744_));
  XOR2X1   g13680(.A(new_n13555_), .B(new_n13392_), .Y(new_n13745_));
  OAI22X1  g13681(.A0(new_n13090_), .A1(new_n5372_), .B0(new_n13366_), .B1(new_n5658_), .Y(new_n13746_));
  AOI21X1  g13682(.A0(new_n12090_), .A1(new_n5960_), .B0(new_n13746_), .Y(new_n13747_));
  OAI21X1  g13683(.A0(new_n13116_), .A1(new_n5657_), .B0(new_n13747_), .Y(new_n13748_));
  XOR2X1   g13684(.A(new_n13748_), .B(new_n3289_), .Y(new_n13749_));
  INVX1    g13685(.A(new_n13749_), .Y(new_n13750_));
  AND2X1   g13686(.A(new_n13750_), .B(new_n13745_), .Y(new_n13751_));
  AND2X1   g13687(.A(new_n13553_), .B(new_n13408_), .Y(new_n13752_));
  XOR2X1   g13688(.A(new_n13752_), .B(new_n13401_), .Y(new_n13753_));
  INVX1    g13689(.A(new_n13753_), .Y(new_n13754_));
  OAI22X1  g13690(.A0(new_n12839_), .A1(new_n5372_), .B0(new_n13090_), .B1(new_n5658_), .Y(new_n13755_));
  AOI21X1  g13691(.A0(new_n12093_), .A1(new_n5960_), .B0(new_n13755_), .Y(new_n13756_));
  OAI21X1  g13692(.A0(new_n13094_), .A1(new_n5657_), .B0(new_n13756_), .Y(new_n13757_));
  XOR2X1   g13693(.A(new_n13757_), .B(new_n3289_), .Y(new_n13758_));
  OR2X1    g13694(.A(new_n13758_), .B(new_n13754_), .Y(new_n13759_));
  XOR2X1   g13695(.A(new_n13552_), .B(new_n13410_), .Y(new_n13760_));
  OAI22X1  g13696(.A0(new_n12840_), .A1(new_n5372_), .B0(new_n12839_), .B1(new_n5658_), .Y(new_n13761_));
  AOI21X1  g13697(.A0(new_n12095_), .A1(new_n5960_), .B0(new_n13761_), .Y(new_n13762_));
  OAI21X1  g13698(.A0(new_n12846_), .A1(new_n5657_), .B0(new_n13762_), .Y(new_n13763_));
  XOR2X1   g13699(.A(new_n13763_), .B(\a[5] ), .Y(new_n13764_));
  AND2X1   g13700(.A(new_n13764_), .B(new_n13760_), .Y(new_n13765_));
  AOI22X1  g13701(.A0(new_n12102_), .A1(new_n5373_), .B0(new_n12099_), .B1(new_n5659_), .Y(new_n13766_));
  OAI21X1  g13702(.A0(new_n12839_), .A1(new_n5959_), .B0(new_n13766_), .Y(new_n13767_));
  AOI21X1  g13703(.A0(new_n12855_), .A1(new_n67_), .B0(new_n13767_), .Y(new_n13768_));
  XOR2X1   g13704(.A(new_n13768_), .B(\a[5] ), .Y(new_n13769_));
  XOR2X1   g13705(.A(new_n13551_), .B(new_n13549_), .Y(new_n13770_));
  INVX1    g13706(.A(new_n13769_), .Y(new_n13771_));
  XOR2X1   g13707(.A(new_n13770_), .B(new_n13771_), .Y(new_n13772_));
  AOI22X1  g13708(.A0(new_n12104_), .A1(new_n5373_), .B0(new_n12102_), .B1(new_n5659_), .Y(new_n13773_));
  OAI21X1  g13709(.A0(new_n12840_), .A1(new_n5959_), .B0(new_n13773_), .Y(new_n13774_));
  AOI21X1  g13710(.A0(new_n12859_), .A1(new_n67_), .B0(new_n13774_), .Y(new_n13775_));
  XOR2X1   g13711(.A(new_n13775_), .B(\a[5] ), .Y(new_n13776_));
  INVX1    g13712(.A(new_n13776_), .Y(new_n13777_));
  AND2X1   g13713(.A(new_n13545_), .B(new_n13429_), .Y(new_n13778_));
  XOR2X1   g13714(.A(new_n13547_), .B(new_n13778_), .Y(new_n13779_));
  AND2X1   g13715(.A(new_n13779_), .B(new_n13777_), .Y(new_n13780_));
  XOR2X1   g13716(.A(new_n13779_), .B(new_n13776_), .Y(new_n13781_));
  INVX1    g13717(.A(new_n13781_), .Y(new_n13782_));
  AOI22X1  g13718(.A0(new_n12107_), .A1(new_n5373_), .B0(new_n12104_), .B1(new_n5659_), .Y(new_n13783_));
  OAI21X1  g13719(.A0(new_n12306_), .A1(new_n5959_), .B0(new_n13783_), .Y(new_n13784_));
  AOI21X1  g13720(.A0(new_n12305_), .A1(new_n67_), .B0(new_n13784_), .Y(new_n13785_));
  XOR2X1   g13721(.A(new_n13785_), .B(\a[5] ), .Y(new_n13786_));
  INVX1    g13722(.A(new_n13544_), .Y(new_n13787_));
  XOR2X1   g13723(.A(new_n13787_), .B(new_n13543_), .Y(new_n13788_));
  OR2X1    g13724(.A(new_n13788_), .B(new_n13786_), .Y(new_n13789_));
  XOR2X1   g13725(.A(new_n13788_), .B(new_n13786_), .Y(new_n13790_));
  INVX1    g13726(.A(new_n13790_), .Y(new_n13791_));
  XOR2X1   g13727(.A(new_n13541_), .B(new_n13436_), .Y(new_n13792_));
  INVX1    g13728(.A(new_n13792_), .Y(new_n13793_));
  OAI22X1  g13729(.A0(new_n12111_), .A1(new_n5372_), .B0(new_n12109_), .B1(new_n5658_), .Y(new_n13794_));
  AOI21X1  g13730(.A0(new_n12104_), .A1(new_n5960_), .B0(new_n13794_), .Y(new_n13795_));
  OAI21X1  g13731(.A0(new_n12693_), .A1(new_n5657_), .B0(new_n13795_), .Y(new_n13796_));
  XOR2X1   g13732(.A(new_n13796_), .B(new_n3289_), .Y(new_n13797_));
  NOR2X1   g13733(.A(new_n13797_), .B(new_n13793_), .Y(new_n13798_));
  XOR2X1   g13734(.A(new_n13539_), .B(new_n13445_), .Y(new_n13799_));
  INVX1    g13735(.A(new_n13799_), .Y(new_n13800_));
  OAI22X1  g13736(.A0(new_n12113_), .A1(new_n5372_), .B0(new_n12111_), .B1(new_n5658_), .Y(new_n13801_));
  AOI21X1  g13737(.A0(new_n12107_), .A1(new_n5960_), .B0(new_n13801_), .Y(new_n13802_));
  OAI21X1  g13738(.A0(new_n12708_), .A1(new_n5657_), .B0(new_n13802_), .Y(new_n13803_));
  XOR2X1   g13739(.A(new_n13803_), .B(new_n3289_), .Y(new_n13804_));
  XOR2X1   g13740(.A(new_n13537_), .B(new_n13455_), .Y(new_n13805_));
  INVX1    g13741(.A(new_n13805_), .Y(new_n13806_));
  OAI22X1  g13742(.A0(new_n12117_), .A1(new_n5372_), .B0(new_n12113_), .B1(new_n5658_), .Y(new_n13807_));
  AOI21X1  g13743(.A0(new_n12208_), .A1(new_n5960_), .B0(new_n13807_), .Y(new_n13808_));
  OAI21X1  g13744(.A0(new_n12685_), .A1(new_n5657_), .B0(new_n13808_), .Y(new_n13809_));
  XOR2X1   g13745(.A(new_n13809_), .B(new_n3289_), .Y(new_n13810_));
  OR2X1    g13746(.A(new_n13810_), .B(new_n13806_), .Y(new_n13811_));
  AOI22X1  g13747(.A0(new_n12133_), .A1(new_n5373_), .B0(new_n12720_), .B1(new_n5659_), .Y(new_n13812_));
  OAI21X1  g13748(.A0(new_n12113_), .A1(new_n5959_), .B0(new_n13812_), .Y(new_n13813_));
  AOI21X1  g13749(.A0(new_n12719_), .A1(new_n67_), .B0(new_n13813_), .Y(new_n13814_));
  XOR2X1   g13750(.A(new_n13814_), .B(\a[5] ), .Y(new_n13815_));
  INVX1    g13751(.A(new_n13815_), .Y(new_n13816_));
  XOR2X1   g13752(.A(new_n13536_), .B(new_n13535_), .Y(new_n13817_));
  NAND2X1  g13753(.A(new_n13817_), .B(new_n13816_), .Y(new_n13818_));
  XOR2X1   g13754(.A(new_n13817_), .B(new_n13815_), .Y(new_n13819_));
  AOI22X1  g13755(.A0(new_n12138_), .A1(new_n5373_), .B0(new_n12133_), .B1(new_n5659_), .Y(new_n13820_));
  OAI21X1  g13756(.A0(new_n12117_), .A1(new_n5959_), .B0(new_n13820_), .Y(new_n13821_));
  AOI21X1  g13757(.A0(new_n12526_), .A1(new_n67_), .B0(new_n13821_), .Y(new_n13822_));
  XOR2X1   g13758(.A(new_n13822_), .B(\a[5] ), .Y(new_n13823_));
  INVX1    g13759(.A(new_n13534_), .Y(new_n13824_));
  XOR2X1   g13760(.A(new_n13824_), .B(new_n13533_), .Y(new_n13825_));
  NOR2X1   g13761(.A(new_n13825_), .B(new_n13823_), .Y(new_n13826_));
  XOR2X1   g13762(.A(new_n13825_), .B(new_n13823_), .Y(new_n13827_));
  INVX1    g13763(.A(new_n13827_), .Y(new_n13828_));
  AOI22X1  g13764(.A0(new_n12141_), .A1(new_n5373_), .B0(new_n12138_), .B1(new_n5659_), .Y(new_n13829_));
  OAI21X1  g13765(.A0(new_n12134_), .A1(new_n5959_), .B0(new_n13829_), .Y(new_n13830_));
  AOI21X1  g13766(.A0(new_n12536_), .A1(new_n67_), .B0(new_n13830_), .Y(new_n13831_));
  XOR2X1   g13767(.A(new_n13831_), .B(new_n3289_), .Y(new_n13832_));
  AND2X1   g13768(.A(new_n13530_), .B(new_n13483_), .Y(new_n13833_));
  XOR2X1   g13769(.A(new_n13531_), .B(new_n13833_), .Y(new_n13834_));
  INVX1    g13770(.A(new_n13834_), .Y(new_n13835_));
  XOR2X1   g13771(.A(new_n13835_), .B(new_n13832_), .Y(new_n13836_));
  INVX1    g13772(.A(new_n13484_), .Y(new_n13837_));
  XOR2X1   g13773(.A(new_n13529_), .B(new_n13837_), .Y(new_n13838_));
  AOI22X1  g13774(.A0(new_n12144_), .A1(new_n5373_), .B0(new_n12141_), .B1(new_n5659_), .Y(new_n13839_));
  OAI21X1  g13775(.A0(new_n12314_), .A1(new_n5959_), .B0(new_n13839_), .Y(new_n13840_));
  AOI21X1  g13776(.A0(new_n12313_), .A1(new_n67_), .B0(new_n13840_), .Y(new_n13841_));
  XOR2X1   g13777(.A(new_n13841_), .B(\a[5] ), .Y(new_n13842_));
  NOR2X1   g13778(.A(new_n13842_), .B(new_n13838_), .Y(new_n13843_));
  XOR2X1   g13779(.A(new_n13528_), .B(new_n13527_), .Y(new_n13844_));
  NAND2X1  g13780(.A(new_n12141_), .B(new_n5960_), .Y(new_n13845_));
  AOI22X1  g13781(.A0(new_n12148_), .A1(new_n5373_), .B0(new_n12144_), .B1(new_n5659_), .Y(new_n13846_));
  AND2X1   g13782(.A(new_n13846_), .B(new_n13845_), .Y(new_n13847_));
  OAI21X1  g13783(.A0(new_n12444_), .A1(new_n5657_), .B0(new_n13847_), .Y(new_n13848_));
  XOR2X1   g13784(.A(new_n13848_), .B(new_n3289_), .Y(new_n13849_));
  INVX1    g13785(.A(new_n13849_), .Y(new_n13850_));
  NAND2X1  g13786(.A(new_n13850_), .B(new_n13844_), .Y(new_n13851_));
  XOR2X1   g13787(.A(new_n13526_), .B(new_n13501_), .Y(new_n13852_));
  INVX1    g13788(.A(new_n13852_), .Y(new_n13853_));
  OAI22X1  g13789(.A0(new_n12322_), .A1(new_n5372_), .B0(new_n12186_), .B1(new_n5658_), .Y(new_n13854_));
  AOI21X1  g13790(.A0(new_n12144_), .A1(new_n5960_), .B0(new_n13854_), .Y(new_n13855_));
  OAI21X1  g13791(.A0(new_n12453_), .A1(new_n5657_), .B0(new_n13855_), .Y(new_n13856_));
  XOR2X1   g13792(.A(new_n13856_), .B(new_n3289_), .Y(new_n13857_));
  NOR2X1   g13793(.A(new_n13857_), .B(new_n13853_), .Y(new_n13858_));
  AOI22X1  g13794(.A0(new_n12155_), .A1(new_n5373_), .B0(new_n12151_), .B1(new_n5659_), .Y(new_n13859_));
  OAI21X1  g13795(.A0(new_n12186_), .A1(new_n5959_), .B0(new_n13859_), .Y(new_n13860_));
  AOI21X1  g13796(.A0(new_n12430_), .A1(new_n67_), .B0(new_n13860_), .Y(new_n13861_));
  XOR2X1   g13797(.A(new_n13861_), .B(\a[5] ), .Y(new_n13862_));
  INVX1    g13798(.A(new_n13862_), .Y(new_n13863_));
  XOR2X1   g13799(.A(new_n13525_), .B(new_n13524_), .Y(new_n13864_));
  NAND2X1  g13800(.A(new_n13864_), .B(new_n13863_), .Y(new_n13865_));
  XOR2X1   g13801(.A(new_n13864_), .B(new_n13862_), .Y(new_n13866_));
  XOR2X1   g13802(.A(new_n13522_), .B(new_n2995_), .Y(new_n13867_));
  XOR2X1   g13803(.A(new_n13867_), .B(new_n13519_), .Y(new_n13868_));
  AOI22X1  g13804(.A0(new_n12158_), .A1(new_n5373_), .B0(new_n12155_), .B1(new_n5659_), .Y(new_n13869_));
  OAI21X1  g13805(.A0(new_n12322_), .A1(new_n5959_), .B0(new_n13869_), .Y(new_n13870_));
  AOI21X1  g13806(.A0(new_n12321_), .A1(new_n67_), .B0(new_n13870_), .Y(new_n13871_));
  XOR2X1   g13807(.A(new_n13871_), .B(\a[5] ), .Y(new_n13872_));
  NOR2X1   g13808(.A(new_n13872_), .B(new_n13868_), .Y(new_n13873_));
  AOI22X1  g13809(.A0(new_n12162_), .A1(new_n5373_), .B0(new_n12158_), .B1(new_n5659_), .Y(new_n13874_));
  OAI21X1  g13810(.A0(new_n12353_), .A1(new_n5959_), .B0(new_n13874_), .Y(new_n13875_));
  AOI21X1  g13811(.A0(new_n12352_), .A1(new_n67_), .B0(new_n13875_), .Y(new_n13876_));
  XOR2X1   g13812(.A(new_n13876_), .B(\a[5] ), .Y(new_n13877_));
  INVX1    g13813(.A(new_n13877_), .Y(new_n13878_));
  NOR3X1   g13814(.A(new_n13512_), .B(new_n13511_), .C(new_n2995_), .Y(new_n13879_));
  XOR2X1   g13815(.A(new_n13515_), .B(\a[8] ), .Y(new_n13880_));
  XOR2X1   g13816(.A(new_n13880_), .B(new_n13879_), .Y(new_n13881_));
  NAND2X1  g13817(.A(new_n13881_), .B(new_n13878_), .Y(new_n13882_));
  XOR2X1   g13818(.A(new_n13881_), .B(new_n13877_), .Y(new_n13883_));
  NOR2X1   g13819(.A(new_n13512_), .B(new_n2995_), .Y(new_n13884_));
  XOR2X1   g13820(.A(new_n13884_), .B(new_n13511_), .Y(new_n13885_));
  OAI22X1  g13821(.A0(new_n12168_), .A1(new_n5372_), .B0(new_n12329_), .B1(new_n5658_), .Y(new_n13886_));
  AOI21X1  g13822(.A0(new_n12158_), .A1(new_n5960_), .B0(new_n13886_), .Y(new_n13887_));
  OAI21X1  g13823(.A0(new_n12368_), .A1(new_n5657_), .B0(new_n13887_), .Y(new_n13888_));
  XOR2X1   g13824(.A(new_n13888_), .B(new_n3289_), .Y(new_n13889_));
  NOR2X1   g13825(.A(new_n13889_), .B(new_n13885_), .Y(new_n13890_));
  OAI22X1  g13826(.A0(new_n12176_), .A1(new_n5658_), .B0(new_n12170_), .B1(new_n5959_), .Y(new_n13891_));
  AOI21X1  g13827(.A0(new_n12337_), .A1(new_n67_), .B0(new_n13891_), .Y(new_n13892_));
  XOR2X1   g13828(.A(new_n13892_), .B(\a[5] ), .Y(new_n13893_));
  AOI21X1  g13829(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n5369_), .Y(new_n13894_));
  OAI22X1  g13830(.A0(new_n12176_), .A1(new_n5372_), .B0(new_n12170_), .B1(new_n5658_), .Y(new_n13895_));
  AOI21X1  g13831(.A0(new_n12165_), .A1(new_n5960_), .B0(new_n13895_), .Y(new_n13896_));
  OAI21X1  g13832(.A0(new_n12344_), .A1(new_n5657_), .B0(new_n13896_), .Y(new_n13897_));
  NOR4X1   g13833(.A(new_n13897_), .B(new_n13894_), .C(new_n13893_), .D(new_n3289_), .Y(new_n13898_));
  AND2X1   g13834(.A(new_n13898_), .B(new_n13512_), .Y(new_n13899_));
  INVX1    g13835(.A(new_n13899_), .Y(new_n13900_));
  INVX1    g13836(.A(new_n13898_), .Y(new_n13901_));
  XOR2X1   g13837(.A(new_n13901_), .B(new_n13512_), .Y(new_n13902_));
  AOI22X1  g13838(.A0(new_n12331_), .A1(new_n5373_), .B0(new_n12165_), .B1(new_n5659_), .Y(new_n13903_));
  OAI21X1  g13839(.A0(new_n12329_), .A1(new_n5959_), .B0(new_n13903_), .Y(new_n13904_));
  AOI21X1  g13840(.A0(new_n12328_), .A1(new_n67_), .B0(new_n13904_), .Y(new_n13905_));
  XOR2X1   g13841(.A(new_n13905_), .B(\a[5] ), .Y(new_n13906_));
  OR2X1    g13842(.A(new_n13906_), .B(new_n13902_), .Y(new_n13907_));
  AND2X1   g13843(.A(new_n13907_), .B(new_n13900_), .Y(new_n13908_));
  INVX1    g13844(.A(new_n13908_), .Y(new_n13909_));
  XOR2X1   g13845(.A(new_n13889_), .B(new_n13885_), .Y(new_n13910_));
  AOI21X1  g13846(.A0(new_n13910_), .A1(new_n13909_), .B0(new_n13890_), .Y(new_n13911_));
  OAI21X1  g13847(.A0(new_n13911_), .A1(new_n13883_), .B0(new_n13882_), .Y(new_n13912_));
  XOR2X1   g13848(.A(new_n13872_), .B(new_n13868_), .Y(new_n13913_));
  AOI21X1  g13849(.A0(new_n13913_), .A1(new_n13912_), .B0(new_n13873_), .Y(new_n13914_));
  OAI21X1  g13850(.A0(new_n13914_), .A1(new_n13866_), .B0(new_n13865_), .Y(new_n13915_));
  XOR2X1   g13851(.A(new_n13857_), .B(new_n13852_), .Y(new_n13916_));
  INVX1    g13852(.A(new_n13916_), .Y(new_n13917_));
  AOI21X1  g13853(.A0(new_n13917_), .A1(new_n13915_), .B0(new_n13858_), .Y(new_n13918_));
  XOR2X1   g13854(.A(new_n13849_), .B(new_n13844_), .Y(new_n13919_));
  OR2X1    g13855(.A(new_n13919_), .B(new_n13918_), .Y(new_n13920_));
  NAND2X1  g13856(.A(new_n13920_), .B(new_n13851_), .Y(new_n13921_));
  XOR2X1   g13857(.A(new_n13842_), .B(new_n13838_), .Y(new_n13922_));
  AOI21X1  g13858(.A0(new_n13922_), .A1(new_n13921_), .B0(new_n13843_), .Y(new_n13923_));
  NOR2X1   g13859(.A(new_n13923_), .B(new_n13836_), .Y(new_n13924_));
  AOI21X1  g13860(.A0(new_n13834_), .A1(new_n13832_), .B0(new_n13924_), .Y(new_n13925_));
  NOR2X1   g13861(.A(new_n13925_), .B(new_n13828_), .Y(new_n13926_));
  NOR2X1   g13862(.A(new_n13926_), .B(new_n13826_), .Y(new_n13927_));
  OAI21X1  g13863(.A0(new_n13927_), .A1(new_n13819_), .B0(new_n13818_), .Y(new_n13928_));
  INVX1    g13864(.A(new_n13928_), .Y(new_n13929_));
  XOR2X1   g13865(.A(new_n13810_), .B(new_n13805_), .Y(new_n13930_));
  OAI21X1  g13866(.A0(new_n13930_), .A1(new_n13929_), .B0(new_n13811_), .Y(new_n13931_));
  INVX1    g13867(.A(new_n13931_), .Y(new_n13932_));
  XOR2X1   g13868(.A(new_n13804_), .B(new_n13799_), .Y(new_n13933_));
  OR2X1    g13869(.A(new_n13933_), .B(new_n13932_), .Y(new_n13934_));
  OAI21X1  g13870(.A0(new_n13804_), .A1(new_n13800_), .B0(new_n13934_), .Y(new_n13935_));
  XOR2X1   g13871(.A(new_n13797_), .B(new_n13793_), .Y(new_n13936_));
  AOI21X1  g13872(.A0(new_n13936_), .A1(new_n13935_), .B0(new_n13798_), .Y(new_n13937_));
  OAI21X1  g13873(.A0(new_n13937_), .A1(new_n13791_), .B0(new_n13789_), .Y(new_n13938_));
  AOI21X1  g13874(.A0(new_n13938_), .A1(new_n13782_), .B0(new_n13780_), .Y(new_n13939_));
  OR2X1    g13875(.A(new_n13939_), .B(new_n13772_), .Y(new_n13940_));
  OAI21X1  g13876(.A0(new_n13770_), .A1(new_n13769_), .B0(new_n13940_), .Y(new_n13941_));
  XOR2X1   g13877(.A(new_n13763_), .B(new_n3289_), .Y(new_n13942_));
  XOR2X1   g13878(.A(new_n13942_), .B(new_n13760_), .Y(new_n13943_));
  INVX1    g13879(.A(new_n13943_), .Y(new_n13944_));
  AOI21X1  g13880(.A0(new_n13944_), .A1(new_n13941_), .B0(new_n13765_), .Y(new_n13945_));
  XOR2X1   g13881(.A(new_n13758_), .B(new_n13753_), .Y(new_n13946_));
  OAI21X1  g13882(.A0(new_n13946_), .A1(new_n13945_), .B0(new_n13759_), .Y(new_n13947_));
  XOR2X1   g13883(.A(new_n13750_), .B(new_n13745_), .Y(new_n13948_));
  AOI21X1  g13884(.A0(new_n13948_), .A1(new_n13947_), .B0(new_n13751_), .Y(new_n13949_));
  OAI21X1  g13885(.A0(new_n13949_), .A1(new_n13744_), .B0(new_n13742_), .Y(new_n13950_));
  AOI21X1  g13886(.A0(new_n13950_), .A1(new_n13735_), .B0(new_n13734_), .Y(new_n13951_));
  OR2X1    g13887(.A(new_n13951_), .B(new_n13728_), .Y(new_n13952_));
  OAI21X1  g13888(.A0(new_n13726_), .A1(new_n13725_), .B0(new_n13952_), .Y(new_n13953_));
  XOR2X1   g13889(.A(new_n13719_), .B(new_n3289_), .Y(new_n13954_));
  XOR2X1   g13890(.A(new_n13954_), .B(new_n13716_), .Y(new_n13955_));
  INVX1    g13891(.A(new_n13955_), .Y(new_n13956_));
  AOI21X1  g13892(.A0(new_n13956_), .A1(new_n13953_), .B0(new_n13721_), .Y(new_n13957_));
  INVX1    g13893(.A(new_n13957_), .Y(new_n13958_));
  XOR2X1   g13894(.A(new_n13715_), .B(new_n13711_), .Y(new_n13959_));
  NAND2X1  g13895(.A(new_n13959_), .B(new_n13958_), .Y(new_n13960_));
  OAI21X1  g13896(.A0(new_n13715_), .A1(new_n13711_), .B0(new_n13960_), .Y(new_n13961_));
  AOI21X1  g13897(.A0(new_n13961_), .A1(new_n13708_), .B0(new_n13707_), .Y(new_n13962_));
  OR2X1    g13898(.A(new_n13962_), .B(new_n13698_), .Y(new_n13963_));
  OAI21X1  g13899(.A0(new_n13696_), .A1(new_n13695_), .B0(new_n13963_), .Y(new_n13964_));
  AOI21X1  g13900(.A0(new_n13964_), .A1(new_n13687_), .B0(new_n13686_), .Y(new_n13965_));
  XOR2X1   g13901(.A(new_n13965_), .B(new_n13677_), .Y(new_n13966_));
  NOR2X1   g13902(.A(new_n12275_), .B(new_n12273_), .Y(new_n13967_));
  INVX1    g13903(.A(new_n13967_), .Y(new_n13968_));
  INVX1    g13904(.A(new_n12276_), .Y(new_n13969_));
  OAI21X1  g13905(.A0(new_n12280_), .A1(new_n13969_), .B0(new_n13968_), .Y(new_n13970_));
  AND2X1   g13906(.A(new_n12268_), .B(new_n12258_), .Y(new_n13971_));
  INVX1    g13907(.A(new_n13971_), .Y(new_n13972_));
  INVX1    g13908(.A(new_n12269_), .Y(new_n13973_));
  OAI21X1  g13909(.A0(new_n12272_), .A1(new_n13973_), .B0(new_n13972_), .Y(new_n13974_));
  INVX1    g13910(.A(new_n13974_), .Y(new_n13975_));
  NOR2X1   g13911(.A(new_n12266_), .B(new_n12035_), .Y(new_n13976_));
  AOI21X1  g13912(.A0(new_n12267_), .A1(new_n12261_), .B0(new_n13976_), .Y(new_n13977_));
  OR2X1    g13913(.A(new_n1306_), .B(new_n766_), .Y(new_n13978_));
  OR4X1    g13914(.A(new_n365_), .B(new_n691_), .C(new_n137_), .D(new_n981_), .Y(new_n13979_));
  OR4X1    g13915(.A(new_n13979_), .B(new_n13978_), .C(new_n3794_), .D(new_n2302_), .Y(new_n13980_));
  OR4X1    g13916(.A(new_n1780_), .B(new_n1225_), .C(new_n1114_), .D(new_n777_), .Y(new_n13981_));
  OR4X1    g13917(.A(new_n13981_), .B(new_n510_), .C(new_n299_), .D(new_n149_), .Y(new_n13982_));
  NOR4X1   g13918(.A(new_n13982_), .B(new_n13980_), .C(new_n7101_), .D(new_n2281_), .Y(new_n13983_));
  NAND3X1  g13919(.A(new_n13983_), .B(new_n2121_), .C(new_n2107_), .Y(new_n13984_));
  INVX1    g13920(.A(new_n13984_), .Y(new_n13985_));
  XOR2X1   g13921(.A(new_n13985_), .B(new_n13977_), .Y(new_n13986_));
  AOI22X1  g13922(.A0(new_n7529_), .A1(new_n1884_), .B0(new_n7522_), .B1(new_n1890_), .Y(new_n13987_));
  OAI21X1  g13923(.A0(new_n7581_), .A1(new_n3498_), .B0(new_n13987_), .Y(new_n13988_));
  AOI21X1  g13924(.A0(new_n7565_), .A1(new_n407_), .B0(new_n13988_), .Y(new_n13989_));
  XOR2X1   g13925(.A(new_n13989_), .B(new_n13986_), .Y(new_n13990_));
  XOR2X1   g13926(.A(new_n13990_), .B(new_n13975_), .Y(new_n13991_));
  OAI22X1  g13927(.A0(new_n7602_), .A1(new_n2431_), .B0(new_n7623_), .B1(new_n2186_), .Y(new_n13992_));
  AOI21X1  g13928(.A0(new_n7590_), .A1(new_n2139_), .B0(new_n13992_), .Y(new_n13993_));
  OAI21X1  g13929(.A0(new_n11583_), .A1(new_n2063_), .B0(new_n13993_), .Y(new_n13994_));
  XOR2X1   g13930(.A(new_n13994_), .B(new_n74_), .Y(new_n13995_));
  XOR2X1   g13931(.A(new_n13995_), .B(new_n13991_), .Y(new_n13996_));
  AND2X1   g13932(.A(new_n13996_), .B(new_n13970_), .Y(new_n13997_));
  INVX1    g13933(.A(new_n13997_), .Y(new_n13998_));
  XOR2X1   g13934(.A(new_n13996_), .B(new_n13970_), .Y(new_n13999_));
  INVX1    g13935(.A(new_n13999_), .Y(new_n14000_));
  AOI22X1  g13936(.A0(new_n7657_), .A1(new_n2424_), .B0(new_n7341_), .B1(new_n2423_), .Y(new_n14001_));
  OAI21X1  g13937(.A0(new_n7644_), .A1(new_n2419_), .B0(new_n14001_), .Y(new_n14002_));
  AOI21X1  g13938(.A0(new_n7656_), .A1(new_n2301_), .B0(new_n14002_), .Y(new_n14003_));
  XOR2X1   g13939(.A(new_n14003_), .B(\a[26] ), .Y(new_n14004_));
  OAI21X1  g13940(.A0(new_n14004_), .A1(new_n14000_), .B0(new_n13998_), .Y(new_n14005_));
  AOI22X1  g13941(.A0(new_n7558_), .A1(new_n1884_), .B0(new_n7529_), .B1(new_n1890_), .Y(new_n14006_));
  OAI21X1  g13942(.A0(new_n7623_), .A1(new_n3498_), .B0(new_n14006_), .Y(new_n14007_));
  AOI21X1  g13943(.A0(new_n7622_), .A1(new_n407_), .B0(new_n14007_), .Y(new_n14008_));
  NOR3X1   g13944(.A(new_n382_), .B(new_n301_), .C(new_n200_), .Y(new_n14009_));
  NOR4X1   g13945(.A(new_n510_), .B(new_n396_), .C(new_n356_), .D(new_n197_), .Y(new_n14010_));
  NOR3X1   g13946(.A(new_n1478_), .B(new_n431_), .C(new_n111_), .Y(new_n14011_));
  NAND4X1  g13947(.A(new_n14011_), .B(new_n14010_), .C(new_n14009_), .D(new_n538_), .Y(new_n14012_));
  OR4X1    g13948(.A(new_n14012_), .B(new_n7101_), .C(new_n2373_), .D(new_n1273_), .Y(new_n14013_));
  NOR3X1   g13949(.A(new_n14013_), .B(new_n2273_), .C(new_n2264_), .Y(new_n14014_));
  AND2X1   g13950(.A(new_n14014_), .B(new_n13984_), .Y(new_n14015_));
  NOR2X1   g13951(.A(new_n14014_), .B(new_n13984_), .Y(new_n14016_));
  NOR3X1   g13952(.A(new_n14016_), .B(new_n14015_), .C(new_n14008_), .Y(new_n14017_));
  NOR2X1   g13953(.A(new_n14017_), .B(new_n14016_), .Y(new_n14018_));
  INVX1    g13954(.A(new_n14018_), .Y(new_n14019_));
  OAI22X1  g13955(.A0(new_n14019_), .A1(new_n14015_), .B0(new_n14017_), .B1(new_n14008_), .Y(new_n14020_));
  INVX1    g13956(.A(new_n14020_), .Y(new_n14021_));
  OR2X1    g13957(.A(new_n13984_), .B(new_n13977_), .Y(new_n14022_));
  OR2X1    g13958(.A(new_n13989_), .B(new_n13986_), .Y(new_n14023_));
  AND2X1   g13959(.A(new_n14023_), .B(new_n14022_), .Y(new_n14024_));
  XOR2X1   g13960(.A(new_n14024_), .B(new_n14021_), .Y(new_n14025_));
  NAND2X1  g13961(.A(new_n13990_), .B(new_n13974_), .Y(new_n14026_));
  OR2X1    g13962(.A(new_n13995_), .B(new_n13991_), .Y(new_n14027_));
  AND2X1   g13963(.A(new_n14027_), .B(new_n14026_), .Y(new_n14028_));
  XOR2X1   g13964(.A(new_n14028_), .B(new_n14025_), .Y(new_n14029_));
  AOI21X1  g13965(.A0(new_n2300_), .A1(new_n2422_), .B0(new_n2418_), .Y(new_n14030_));
  OAI22X1  g13966(.A0(new_n14030_), .A1(new_n8172_), .B0(new_n7644_), .B1(new_n2666_), .Y(new_n14031_));
  AOI21X1  g13967(.A0(new_n7807_), .A1(new_n2301_), .B0(new_n14031_), .Y(new_n14032_));
  XOR2X1   g13968(.A(new_n14032_), .B(\a[26] ), .Y(new_n14033_));
  AOI22X1  g13969(.A0(new_n7590_), .A1(new_n2095_), .B0(new_n7578_), .B1(new_n2185_), .Y(new_n14034_));
  OAI21X1  g13970(.A0(new_n7642_), .A1(new_n2140_), .B0(new_n14034_), .Y(new_n14035_));
  AOI21X1  g13971(.A0(new_n7712_), .A1(new_n2062_), .B0(new_n14035_), .Y(new_n14036_));
  XOR2X1   g13972(.A(new_n14036_), .B(new_n74_), .Y(new_n14037_));
  XOR2X1   g13973(.A(new_n14037_), .B(new_n14033_), .Y(new_n14038_));
  XOR2X1   g13974(.A(new_n14038_), .B(new_n14029_), .Y(new_n14039_));
  AND2X1   g13975(.A(new_n14039_), .B(new_n14005_), .Y(new_n14040_));
  INVX1    g13976(.A(new_n14040_), .Y(new_n14041_));
  XOR2X1   g13977(.A(new_n14004_), .B(new_n13999_), .Y(new_n14042_));
  NOR2X1   g13978(.A(new_n12255_), .B(new_n12251_), .Y(new_n14043_));
  INVX1    g13979(.A(new_n12281_), .Y(new_n14044_));
  AOI21X1  g13980(.A0(new_n14044_), .A1(new_n12256_), .B0(new_n14043_), .Y(new_n14045_));
  NOR2X1   g13981(.A(new_n14045_), .B(new_n14042_), .Y(new_n14046_));
  XOR2X1   g13982(.A(new_n14045_), .B(new_n14042_), .Y(new_n14047_));
  NOR2X1   g13983(.A(new_n12282_), .B(new_n12248_), .Y(new_n14048_));
  INVX1    g13984(.A(new_n14048_), .Y(new_n14049_));
  OAI21X1  g13985(.A0(new_n12284_), .A1(new_n12245_), .B0(new_n14049_), .Y(new_n14050_));
  AOI21X1  g13986(.A0(new_n14050_), .A1(new_n14047_), .B0(new_n14046_), .Y(new_n14051_));
  XOR2X1   g13987(.A(new_n14039_), .B(new_n14005_), .Y(new_n14052_));
  INVX1    g13988(.A(new_n14052_), .Y(new_n14053_));
  OAI21X1  g13989(.A0(new_n14053_), .A1(new_n14051_), .B0(new_n14041_), .Y(new_n14054_));
  OR4X1    g13990(.A(new_n2424_), .B(new_n2423_), .C(new_n2418_), .D(new_n2301_), .Y(new_n14055_));
  AND2X1   g13991(.A(new_n14055_), .B(new_n7341_), .Y(new_n14056_));
  XOR2X1   g13992(.A(new_n14056_), .B(new_n89_), .Y(new_n14057_));
  NOR4X1   g13993(.A(new_n2403_), .B(new_n2402_), .C(new_n2376_), .D(new_n510_), .Y(new_n14058_));
  INVX1    g13994(.A(new_n14058_), .Y(new_n14059_));
  OR4X1    g13995(.A(new_n460_), .B(new_n420_), .C(new_n260_), .D(new_n197_), .Y(new_n14060_));
  NOR4X1   g13996(.A(new_n14060_), .B(new_n14059_), .C(new_n2370_), .D(new_n2360_), .Y(new_n14061_));
  XOR2X1   g13997(.A(new_n14061_), .B(new_n13985_), .Y(new_n14062_));
  XOR2X1   g13998(.A(new_n14062_), .B(new_n14057_), .Y(new_n14063_));
  XOR2X1   g13999(.A(new_n14063_), .B(new_n14019_), .Y(new_n14064_));
  AOI22X1  g14000(.A0(new_n7571_), .A1(new_n1884_), .B0(new_n7558_), .B1(new_n1890_), .Y(new_n14065_));
  OAI21X1  g14001(.A0(new_n7602_), .A1(new_n3498_), .B0(new_n14065_), .Y(new_n14066_));
  AOI21X1  g14002(.A0(new_n7601_), .A1(new_n407_), .B0(new_n14066_), .Y(new_n14067_));
  XOR2X1   g14003(.A(new_n14067_), .B(new_n14064_), .Y(new_n14068_));
  AOI22X1  g14004(.A0(new_n7643_), .A1(new_n2139_), .B0(new_n7590_), .B1(new_n2185_), .Y(new_n14069_));
  OAI21X1  g14005(.A0(new_n7642_), .A1(new_n2431_), .B0(new_n14069_), .Y(new_n14070_));
  AOI21X1  g14006(.A0(new_n7718_), .A1(new_n2062_), .B0(new_n14070_), .Y(new_n14071_));
  XOR2X1   g14007(.A(new_n14071_), .B(\a[29] ), .Y(new_n14072_));
  XOR2X1   g14008(.A(new_n14072_), .B(new_n14068_), .Y(new_n14073_));
  INVX1    g14009(.A(new_n14073_), .Y(new_n14074_));
  NOR2X1   g14010(.A(new_n14024_), .B(new_n14021_), .Y(new_n14075_));
  INVX1    g14011(.A(new_n14028_), .Y(new_n14076_));
  AOI21X1  g14012(.A0(new_n14076_), .A1(new_n14025_), .B0(new_n14075_), .Y(new_n14077_));
  XOR2X1   g14013(.A(new_n14077_), .B(new_n14074_), .Y(new_n14078_));
  INVX1    g14014(.A(new_n14078_), .Y(new_n14079_));
  INVX1    g14015(.A(new_n14033_), .Y(new_n14080_));
  NOR2X1   g14016(.A(new_n14038_), .B(new_n14029_), .Y(new_n14081_));
  AOI21X1  g14017(.A0(new_n14037_), .A1(new_n14080_), .B0(new_n14081_), .Y(new_n14082_));
  XOR2X1   g14018(.A(new_n14082_), .B(new_n14079_), .Y(new_n14083_));
  XOR2X1   g14019(.A(new_n14083_), .B(new_n14054_), .Y(new_n14084_));
  XOR2X1   g14020(.A(new_n14050_), .B(new_n14047_), .Y(new_n14085_));
  INVX1    g14021(.A(new_n14085_), .Y(new_n14086_));
  XOR2X1   g14022(.A(new_n14053_), .B(new_n14051_), .Y(new_n14087_));
  INVX1    g14023(.A(new_n14087_), .Y(new_n14088_));
  OAI22X1  g14024(.A0(new_n14088_), .A1(new_n6307_), .B0(new_n14086_), .B1(new_n6325_), .Y(new_n14089_));
  AOI21X1  g14025(.A0(new_n14084_), .A1(new_n6308_), .B0(new_n14089_), .Y(new_n14090_));
  AND2X1   g14026(.A(new_n14087_), .B(new_n14085_), .Y(new_n14091_));
  INVX1    g14027(.A(new_n14091_), .Y(new_n14092_));
  AND2X1   g14028(.A(new_n14085_), .B(new_n12285_), .Y(new_n14093_));
  NOR2X1   g14029(.A(new_n14085_), .B(new_n12285_), .Y(new_n14094_));
  INVX1    g14030(.A(new_n14094_), .Y(new_n14095_));
  AOI21X1  g14031(.A0(new_n14095_), .A1(new_n12290_), .B0(new_n14093_), .Y(new_n14096_));
  NOR2X1   g14032(.A(new_n14087_), .B(new_n14085_), .Y(new_n14097_));
  OAI21X1  g14033(.A0(new_n14097_), .A1(new_n14096_), .B0(new_n14092_), .Y(new_n14098_));
  INVX1    g14034(.A(new_n14098_), .Y(new_n14099_));
  NOR2X1   g14035(.A(new_n14087_), .B(new_n14084_), .Y(new_n14100_));
  XOR2X1   g14036(.A(new_n14087_), .B(new_n14084_), .Y(new_n14101_));
  AND2X1   g14037(.A(new_n14087_), .B(new_n14084_), .Y(new_n14102_));
  INVX1    g14038(.A(new_n14100_), .Y(new_n14103_));
  AOI21X1  g14039(.A0(new_n14103_), .A1(new_n14098_), .B0(new_n14102_), .Y(new_n14104_));
  INVX1    g14040(.A(new_n14104_), .Y(new_n14105_));
  OAI22X1  g14041(.A0(new_n14105_), .A1(new_n14100_), .B0(new_n14101_), .B1(new_n14099_), .Y(new_n14106_));
  INVX1    g14042(.A(new_n14106_), .Y(new_n14107_));
  OAI21X1  g14043(.A0(new_n14107_), .A1(new_n6298_), .B0(new_n14090_), .Y(new_n14108_));
  XOR2X1   g14044(.A(new_n14108_), .B(new_n3431_), .Y(new_n14109_));
  OR2X1    g14045(.A(new_n14109_), .B(new_n13966_), .Y(new_n14110_));
  XOR2X1   g14046(.A(new_n13959_), .B(new_n13958_), .Y(new_n14111_));
  XOR2X1   g14047(.A(new_n13948_), .B(new_n13947_), .Y(new_n14112_));
  INVX1    g14048(.A(new_n13936_), .Y(new_n14113_));
  XOR2X1   g14049(.A(new_n14113_), .B(new_n13935_), .Y(new_n14114_));
  XOR2X1   g14050(.A(new_n13922_), .B(new_n13921_), .Y(new_n14115_));
  XOR2X1   g14051(.A(new_n13910_), .B(new_n13909_), .Y(new_n14116_));
  INVX1    g14052(.A(new_n14116_), .Y(new_n14117_));
  NOR2X1   g14053(.A(new_n13894_), .B(new_n3289_), .Y(new_n14118_));
  INVX1    g14054(.A(new_n14118_), .Y(new_n14119_));
  NOR2X1   g14055(.A(new_n14119_), .B(new_n13893_), .Y(new_n14120_));
  XOR2X1   g14056(.A(new_n13897_), .B(new_n3289_), .Y(new_n14121_));
  XOR2X1   g14057(.A(new_n14121_), .B(new_n14120_), .Y(new_n14122_));
  INVX1    g14058(.A(new_n14122_), .Y(new_n14123_));
  OAI22X1  g14059(.A0(new_n12176_), .A1(new_n6325_), .B0(new_n12170_), .B1(new_n6307_), .Y(new_n14124_));
  AOI21X1  g14060(.A0(new_n12165_), .A1(new_n6308_), .B0(new_n14124_), .Y(new_n14125_));
  NOR2X1   g14061(.A(new_n14125_), .B(new_n3431_), .Y(new_n14126_));
  NOR2X1   g14062(.A(new_n12344_), .B(new_n6351_), .Y(new_n14127_));
  AND2X1   g14063(.A(new_n12337_), .B(new_n6350_), .Y(new_n14128_));
  NOR2X1   g14064(.A(new_n12170_), .B(new_n6362_), .Y(new_n14129_));
  AOI21X1  g14065(.A0(new_n12175_), .A1(new_n12171_), .B0(new_n6361_), .Y(new_n14130_));
  OAI21X1  g14066(.A0(new_n12176_), .A1(new_n6357_), .B0(\a[2] ), .Y(new_n14131_));
  OR4X1    g14067(.A(new_n14131_), .B(new_n14130_), .C(new_n14129_), .D(new_n14128_), .Y(new_n14132_));
  NOR3X1   g14068(.A(new_n14132_), .B(new_n14127_), .C(new_n14126_), .Y(new_n14133_));
  AND2X1   g14069(.A(new_n14133_), .B(new_n13894_), .Y(new_n14134_));
  NOR2X1   g14070(.A(new_n14133_), .B(new_n13894_), .Y(new_n14135_));
  AND2X1   g14071(.A(new_n12328_), .B(new_n5972_), .Y(new_n14136_));
  AOI22X1  g14072(.A0(new_n12331_), .A1(new_n5970_), .B0(new_n12165_), .B1(new_n6300_), .Y(new_n14137_));
  OAI21X1  g14073(.A0(new_n12329_), .A1(new_n6309_), .B0(new_n14137_), .Y(new_n14138_));
  OAI21X1  g14074(.A0(new_n14138_), .A1(new_n14136_), .B0(new_n3431_), .Y(new_n14139_));
  NAND2X1  g14075(.A(new_n12328_), .B(new_n5972_), .Y(new_n14140_));
  INVX1    g14076(.A(new_n14138_), .Y(new_n14141_));
  NAND3X1  g14077(.A(new_n14141_), .B(new_n14140_), .C(\a[2] ), .Y(new_n14142_));
  AOI21X1  g14078(.A0(new_n14142_), .A1(new_n14139_), .B0(new_n14135_), .Y(new_n14143_));
  OAI22X1  g14079(.A0(new_n12168_), .A1(new_n6325_), .B0(new_n12329_), .B1(new_n6307_), .Y(new_n14144_));
  AOI21X1  g14080(.A0(new_n12158_), .A1(new_n6308_), .B0(new_n14144_), .Y(new_n14145_));
  NAND2X1  g14081(.A(new_n14145_), .B(new_n6298_), .Y(new_n14146_));
  NAND2X1  g14082(.A(new_n14145_), .B(new_n12368_), .Y(new_n14147_));
  AOI21X1  g14083(.A0(new_n14147_), .A1(new_n14146_), .B0(new_n3431_), .Y(new_n14148_));
  AND2X1   g14084(.A(new_n14145_), .B(new_n6298_), .Y(new_n14149_));
  AND2X1   g14085(.A(new_n14145_), .B(new_n12368_), .Y(new_n14150_));
  NOR3X1   g14086(.A(new_n14150_), .B(new_n14149_), .C(\a[2] ), .Y(new_n14151_));
  NOR4X1   g14087(.A(new_n14151_), .B(new_n14148_), .C(new_n14143_), .D(new_n14134_), .Y(new_n14152_));
  XOR2X1   g14088(.A(new_n14119_), .B(new_n13893_), .Y(new_n14153_));
  INVX1    g14089(.A(new_n14153_), .Y(new_n14154_));
  OAI22X1  g14090(.A0(new_n14151_), .A1(new_n14148_), .B0(new_n14143_), .B1(new_n14134_), .Y(new_n14155_));
  OAI21X1  g14091(.A0(new_n14154_), .A1(new_n14152_), .B0(new_n14155_), .Y(new_n14156_));
  NAND2X1  g14092(.A(new_n14156_), .B(new_n14123_), .Y(new_n14157_));
  AOI22X1  g14093(.A0(new_n12162_), .A1(new_n5970_), .B0(new_n12158_), .B1(new_n6300_), .Y(new_n14158_));
  OAI21X1  g14094(.A0(new_n12353_), .A1(new_n6309_), .B0(new_n14158_), .Y(new_n14159_));
  AOI21X1  g14095(.A0(new_n12352_), .A1(new_n5972_), .B0(new_n14159_), .Y(new_n14160_));
  XOR2X1   g14096(.A(new_n14160_), .B(new_n3431_), .Y(new_n14161_));
  OAI21X1  g14097(.A0(new_n14156_), .A1(new_n14123_), .B0(new_n14161_), .Y(new_n14162_));
  OAI22X1  g14098(.A0(new_n12396_), .A1(new_n6325_), .B0(new_n12353_), .B1(new_n6307_), .Y(new_n14163_));
  AOI21X1  g14099(.A0(new_n12151_), .A1(new_n6308_), .B0(new_n14163_), .Y(new_n14164_));
  OAI21X1  g14100(.A0(new_n12320_), .A1(new_n6298_), .B0(new_n14164_), .Y(new_n14165_));
  XOR2X1   g14101(.A(new_n14165_), .B(new_n3431_), .Y(new_n14166_));
  AOI21X1  g14102(.A0(new_n14162_), .A1(new_n14157_), .B0(new_n14166_), .Y(new_n14167_));
  NAND3X1  g14103(.A(new_n14166_), .B(new_n14162_), .C(new_n14157_), .Y(new_n14168_));
  XOR2X1   g14104(.A(new_n13906_), .B(new_n13902_), .Y(new_n14169_));
  AOI21X1  g14105(.A0(new_n14169_), .A1(new_n14168_), .B0(new_n14167_), .Y(new_n14170_));
  NOR2X1   g14106(.A(new_n14170_), .B(new_n14117_), .Y(new_n14171_));
  AOI22X1  g14107(.A0(new_n12155_), .A1(new_n5970_), .B0(new_n12151_), .B1(new_n6300_), .Y(new_n14172_));
  OAI21X1  g14108(.A0(new_n12186_), .A1(new_n6309_), .B0(new_n14172_), .Y(new_n14173_));
  AOI21X1  g14109(.A0(new_n12430_), .A1(new_n5972_), .B0(new_n14173_), .Y(new_n14174_));
  XOR2X1   g14110(.A(new_n14174_), .B(\a[2] ), .Y(new_n14175_));
  AOI21X1  g14111(.A0(new_n14170_), .A1(new_n14117_), .B0(new_n14175_), .Y(new_n14176_));
  OAI22X1  g14112(.A0(new_n12322_), .A1(new_n6325_), .B0(new_n12186_), .B1(new_n6307_), .Y(new_n14177_));
  AOI21X1  g14113(.A0(new_n12144_), .A1(new_n6308_), .B0(new_n14177_), .Y(new_n14178_));
  OAI21X1  g14114(.A0(new_n12453_), .A1(new_n6298_), .B0(new_n14178_), .Y(new_n14179_));
  XOR2X1   g14115(.A(new_n14179_), .B(\a[2] ), .Y(new_n14180_));
  NOR3X1   g14116(.A(new_n14180_), .B(new_n14176_), .C(new_n14171_), .Y(new_n14181_));
  XOR2X1   g14117(.A(new_n13911_), .B(new_n13883_), .Y(new_n14182_));
  INVX1    g14118(.A(new_n14182_), .Y(new_n14183_));
  OAI21X1  g14119(.A0(new_n14176_), .A1(new_n14171_), .B0(new_n14180_), .Y(new_n14184_));
  OAI21X1  g14120(.A0(new_n14183_), .A1(new_n14181_), .B0(new_n14184_), .Y(new_n14185_));
  OAI22X1  g14121(.A0(new_n12186_), .A1(new_n6325_), .B0(new_n12192_), .B1(new_n6307_), .Y(new_n14186_));
  AOI21X1  g14122(.A0(new_n12141_), .A1(new_n6308_), .B0(new_n14186_), .Y(new_n14187_));
  OAI21X1  g14123(.A0(new_n12444_), .A1(new_n6298_), .B0(new_n14187_), .Y(new_n14188_));
  XOR2X1   g14124(.A(new_n14188_), .B(\a[2] ), .Y(new_n14189_));
  XOR2X1   g14125(.A(new_n13913_), .B(new_n13912_), .Y(new_n14190_));
  OAI21X1  g14126(.A0(new_n14189_), .A1(new_n14185_), .B0(new_n14190_), .Y(new_n14191_));
  NAND2X1  g14127(.A(new_n14189_), .B(new_n14185_), .Y(new_n14192_));
  INVX1    g14128(.A(new_n12313_), .Y(new_n14193_));
  INVX1    g14129(.A(new_n12141_), .Y(new_n14194_));
  OAI22X1  g14130(.A0(new_n12192_), .A1(new_n6325_), .B0(new_n14194_), .B1(new_n6307_), .Y(new_n14195_));
  AOI21X1  g14131(.A0(new_n12138_), .A1(new_n6308_), .B0(new_n14195_), .Y(new_n14196_));
  OAI21X1  g14132(.A0(new_n14193_), .A1(new_n6298_), .B0(new_n14196_), .Y(new_n14197_));
  XOR2X1   g14133(.A(new_n14197_), .B(new_n3431_), .Y(new_n14198_));
  NAND3X1  g14134(.A(new_n14198_), .B(new_n14192_), .C(new_n14191_), .Y(new_n14199_));
  XOR2X1   g14135(.A(new_n13914_), .B(new_n13866_), .Y(new_n14200_));
  AOI21X1  g14136(.A0(new_n14192_), .A1(new_n14191_), .B0(new_n14198_), .Y(new_n14201_));
  AOI21X1  g14137(.A0(new_n14200_), .A1(new_n14199_), .B0(new_n14201_), .Y(new_n14202_));
  XOR2X1   g14138(.A(new_n13917_), .B(new_n13915_), .Y(new_n14203_));
  INVX1    g14139(.A(new_n14203_), .Y(new_n14204_));
  NOR2X1   g14140(.A(new_n14204_), .B(new_n14202_), .Y(new_n14205_));
  AOI22X1  g14141(.A0(new_n12141_), .A1(new_n5970_), .B0(new_n12138_), .B1(new_n6300_), .Y(new_n14206_));
  OAI21X1  g14142(.A0(new_n12134_), .A1(new_n6309_), .B0(new_n14206_), .Y(new_n14207_));
  AOI21X1  g14143(.A0(new_n12536_), .A1(new_n5972_), .B0(new_n14207_), .Y(new_n14208_));
  XOR2X1   g14144(.A(new_n14208_), .B(\a[2] ), .Y(new_n14209_));
  AOI21X1  g14145(.A0(new_n14204_), .A1(new_n14202_), .B0(new_n14209_), .Y(new_n14210_));
  NAND2X1  g14146(.A(new_n13849_), .B(new_n13844_), .Y(new_n14211_));
  OR2X1    g14147(.A(new_n13849_), .B(new_n13844_), .Y(new_n14212_));
  NAND3X1  g14148(.A(new_n14212_), .B(new_n14211_), .C(new_n13918_), .Y(new_n14213_));
  AND2X1   g14149(.A(new_n14213_), .B(new_n13920_), .Y(new_n14214_));
  OAI21X1  g14150(.A0(new_n14210_), .A1(new_n14205_), .B0(new_n14214_), .Y(new_n14215_));
  NOR3X1   g14151(.A(new_n14214_), .B(new_n14210_), .C(new_n14205_), .Y(new_n14216_));
  AOI22X1  g14152(.A0(new_n12138_), .A1(new_n5970_), .B0(new_n12133_), .B1(new_n6300_), .Y(new_n14217_));
  OAI21X1  g14153(.A0(new_n12117_), .A1(new_n6309_), .B0(new_n14217_), .Y(new_n14218_));
  AOI21X1  g14154(.A0(new_n12526_), .A1(new_n5972_), .B0(new_n14218_), .Y(new_n14219_));
  XOR2X1   g14155(.A(new_n14219_), .B(\a[2] ), .Y(new_n14220_));
  OAI21X1  g14156(.A0(new_n14220_), .A1(new_n14216_), .B0(new_n14215_), .Y(new_n14221_));
  NAND2X1  g14157(.A(new_n14221_), .B(new_n14115_), .Y(new_n14222_));
  AOI22X1  g14158(.A0(new_n12133_), .A1(new_n5970_), .B0(new_n12720_), .B1(new_n6300_), .Y(new_n14223_));
  OAI21X1  g14159(.A0(new_n12113_), .A1(new_n6309_), .B0(new_n14223_), .Y(new_n14224_));
  AOI21X1  g14160(.A0(new_n12719_), .A1(new_n5972_), .B0(new_n14224_), .Y(new_n14225_));
  XOR2X1   g14161(.A(new_n14225_), .B(new_n3431_), .Y(new_n14226_));
  OAI21X1  g14162(.A0(new_n14221_), .A1(new_n14115_), .B0(new_n14226_), .Y(new_n14227_));
  OAI22X1  g14163(.A0(new_n12117_), .A1(new_n6325_), .B0(new_n12113_), .B1(new_n6307_), .Y(new_n14228_));
  AOI21X1  g14164(.A0(new_n12208_), .A1(new_n6308_), .B0(new_n14228_), .Y(new_n14229_));
  OAI21X1  g14165(.A0(new_n12685_), .A1(new_n6298_), .B0(new_n14229_), .Y(new_n14230_));
  XOR2X1   g14166(.A(new_n14230_), .B(new_n3431_), .Y(new_n14231_));
  NAND3X1  g14167(.A(new_n14231_), .B(new_n14227_), .C(new_n14222_), .Y(new_n14232_));
  XOR2X1   g14168(.A(new_n13923_), .B(new_n13836_), .Y(new_n14233_));
  AOI21X1  g14169(.A0(new_n14227_), .A1(new_n14222_), .B0(new_n14231_), .Y(new_n14234_));
  AOI21X1  g14170(.A0(new_n14233_), .A1(new_n14232_), .B0(new_n14234_), .Y(new_n14235_));
  OAI22X1  g14171(.A0(new_n12113_), .A1(new_n6325_), .B0(new_n12111_), .B1(new_n6307_), .Y(new_n14236_));
  AOI21X1  g14172(.A0(new_n12107_), .A1(new_n6308_), .B0(new_n14236_), .Y(new_n14237_));
  OAI21X1  g14173(.A0(new_n12708_), .A1(new_n6298_), .B0(new_n14237_), .Y(new_n14238_));
  XOR2X1   g14174(.A(new_n14238_), .B(new_n3431_), .Y(new_n14239_));
  XOR2X1   g14175(.A(new_n13925_), .B(new_n13828_), .Y(new_n14240_));
  INVX1    g14176(.A(new_n14240_), .Y(new_n14241_));
  AOI21X1  g14177(.A0(new_n14239_), .A1(new_n14235_), .B0(new_n14241_), .Y(new_n14242_));
  NOR2X1   g14178(.A(new_n14239_), .B(new_n14235_), .Y(new_n14243_));
  OAI22X1  g14179(.A0(new_n12111_), .A1(new_n6325_), .B0(new_n12109_), .B1(new_n6307_), .Y(new_n14244_));
  AOI21X1  g14180(.A0(new_n12104_), .A1(new_n6308_), .B0(new_n14244_), .Y(new_n14245_));
  OAI21X1  g14181(.A0(new_n12693_), .A1(new_n6298_), .B0(new_n14245_), .Y(new_n14246_));
  XOR2X1   g14182(.A(new_n14246_), .B(new_n3431_), .Y(new_n14247_));
  INVX1    g14183(.A(new_n14247_), .Y(new_n14248_));
  NOR3X1   g14184(.A(new_n14248_), .B(new_n14243_), .C(new_n14242_), .Y(new_n14249_));
  XOR2X1   g14185(.A(new_n13927_), .B(new_n13819_), .Y(new_n14250_));
  INVX1    g14186(.A(new_n14250_), .Y(new_n14251_));
  OAI21X1  g14187(.A0(new_n14243_), .A1(new_n14242_), .B0(new_n14248_), .Y(new_n14252_));
  OAI21X1  g14188(.A0(new_n14251_), .A1(new_n14249_), .B0(new_n14252_), .Y(new_n14253_));
  XOR2X1   g14189(.A(new_n13930_), .B(new_n13929_), .Y(new_n14254_));
  NAND2X1  g14190(.A(new_n14254_), .B(new_n14253_), .Y(new_n14255_));
  AOI22X1  g14191(.A0(new_n12107_), .A1(new_n5970_), .B0(new_n12104_), .B1(new_n6300_), .Y(new_n14256_));
  OAI21X1  g14192(.A0(new_n12306_), .A1(new_n6309_), .B0(new_n14256_), .Y(new_n14257_));
  AOI21X1  g14193(.A0(new_n12305_), .A1(new_n5972_), .B0(new_n14257_), .Y(new_n14258_));
  XOR2X1   g14194(.A(new_n14258_), .B(\a[2] ), .Y(new_n14259_));
  INVX1    g14195(.A(new_n14259_), .Y(new_n14260_));
  OAI21X1  g14196(.A0(new_n14254_), .A1(new_n14253_), .B0(new_n14260_), .Y(new_n14261_));
  XOR2X1   g14197(.A(new_n13933_), .B(new_n13931_), .Y(new_n14262_));
  AOI21X1  g14198(.A0(new_n14261_), .A1(new_n14255_), .B0(new_n14262_), .Y(new_n14263_));
  NAND3X1  g14199(.A(new_n14262_), .B(new_n14261_), .C(new_n14255_), .Y(new_n14264_));
  AOI22X1  g14200(.A0(new_n12104_), .A1(new_n5970_), .B0(new_n12102_), .B1(new_n6300_), .Y(new_n14265_));
  OAI21X1  g14201(.A0(new_n12840_), .A1(new_n6309_), .B0(new_n14265_), .Y(new_n14266_));
  AOI21X1  g14202(.A0(new_n12859_), .A1(new_n5972_), .B0(new_n14266_), .Y(new_n14267_));
  XOR2X1   g14203(.A(new_n14267_), .B(\a[2] ), .Y(new_n14268_));
  INVX1    g14204(.A(new_n14268_), .Y(new_n14269_));
  AOI21X1  g14205(.A0(new_n14269_), .A1(new_n14264_), .B0(new_n14263_), .Y(new_n14270_));
  NOR2X1   g14206(.A(new_n14270_), .B(new_n14114_), .Y(new_n14271_));
  AOI22X1  g14207(.A0(new_n12102_), .A1(new_n5970_), .B0(new_n12099_), .B1(new_n6300_), .Y(new_n14272_));
  OAI21X1  g14208(.A0(new_n12839_), .A1(new_n6309_), .B0(new_n14272_), .Y(new_n14273_));
  AOI21X1  g14209(.A0(new_n12855_), .A1(new_n5972_), .B0(new_n14273_), .Y(new_n14274_));
  XOR2X1   g14210(.A(new_n14274_), .B(\a[2] ), .Y(new_n14275_));
  AOI21X1  g14211(.A0(new_n14270_), .A1(new_n14114_), .B0(new_n14275_), .Y(new_n14276_));
  OAI22X1  g14212(.A0(new_n12840_), .A1(new_n6325_), .B0(new_n12839_), .B1(new_n6307_), .Y(new_n14277_));
  AOI21X1  g14213(.A0(new_n12095_), .A1(new_n6308_), .B0(new_n14277_), .Y(new_n14278_));
  OAI21X1  g14214(.A0(new_n12846_), .A1(new_n6298_), .B0(new_n14278_), .Y(new_n14279_));
  XOR2X1   g14215(.A(new_n14279_), .B(new_n3431_), .Y(new_n14280_));
  INVX1    g14216(.A(new_n14280_), .Y(new_n14281_));
  NOR3X1   g14217(.A(new_n14281_), .B(new_n14276_), .C(new_n14271_), .Y(new_n14282_));
  XOR2X1   g14218(.A(new_n13937_), .B(new_n13791_), .Y(new_n14283_));
  INVX1    g14219(.A(new_n14283_), .Y(new_n14284_));
  OAI21X1  g14220(.A0(new_n14276_), .A1(new_n14271_), .B0(new_n14281_), .Y(new_n14285_));
  OAI21X1  g14221(.A0(new_n14284_), .A1(new_n14282_), .B0(new_n14285_), .Y(new_n14286_));
  OAI22X1  g14222(.A0(new_n12839_), .A1(new_n6325_), .B0(new_n13090_), .B1(new_n6307_), .Y(new_n14287_));
  AOI21X1  g14223(.A0(new_n12093_), .A1(new_n6308_), .B0(new_n14287_), .Y(new_n14288_));
  OAI21X1  g14224(.A0(new_n13094_), .A1(new_n6298_), .B0(new_n14288_), .Y(new_n14289_));
  XOR2X1   g14225(.A(new_n14289_), .B(new_n3431_), .Y(new_n14290_));
  INVX1    g14226(.A(new_n14290_), .Y(new_n14291_));
  XOR2X1   g14227(.A(new_n13938_), .B(new_n13782_), .Y(new_n14292_));
  OAI21X1  g14228(.A0(new_n14291_), .A1(new_n14286_), .B0(new_n14292_), .Y(new_n14293_));
  NAND2X1  g14229(.A(new_n14291_), .B(new_n14286_), .Y(new_n14294_));
  OAI22X1  g14230(.A0(new_n13090_), .A1(new_n6325_), .B0(new_n13366_), .B1(new_n6307_), .Y(new_n14295_));
  AOI21X1  g14231(.A0(new_n12090_), .A1(new_n6308_), .B0(new_n14295_), .Y(new_n14296_));
  OAI21X1  g14232(.A0(new_n13116_), .A1(new_n6298_), .B0(new_n14296_), .Y(new_n14297_));
  XOR2X1   g14233(.A(new_n14297_), .B(new_n3431_), .Y(new_n14298_));
  NAND3X1  g14234(.A(new_n14298_), .B(new_n14294_), .C(new_n14293_), .Y(new_n14299_));
  XOR2X1   g14235(.A(new_n13939_), .B(new_n13772_), .Y(new_n14300_));
  AOI21X1  g14236(.A0(new_n14294_), .A1(new_n14293_), .B0(new_n14298_), .Y(new_n14301_));
  AOI21X1  g14237(.A0(new_n14300_), .A1(new_n14299_), .B0(new_n14301_), .Y(new_n14302_));
  XOR2X1   g14238(.A(new_n13944_), .B(new_n13941_), .Y(new_n14303_));
  INVX1    g14239(.A(new_n14303_), .Y(new_n14304_));
  NOR2X1   g14240(.A(new_n14304_), .B(new_n14302_), .Y(new_n14305_));
  AOI22X1  g14241(.A0(new_n12093_), .A1(new_n5970_), .B0(new_n12090_), .B1(new_n6300_), .Y(new_n14306_));
  OAI21X1  g14242(.A0(new_n13104_), .A1(new_n6309_), .B0(new_n14306_), .Y(new_n14307_));
  AOI21X1  g14243(.A0(new_n13103_), .A1(new_n5972_), .B0(new_n14307_), .Y(new_n14308_));
  XOR2X1   g14244(.A(new_n14308_), .B(\a[2] ), .Y(new_n14309_));
  AOI21X1  g14245(.A0(new_n14304_), .A1(new_n14302_), .B0(new_n14309_), .Y(new_n14310_));
  XOR2X1   g14246(.A(new_n13946_), .B(new_n13945_), .Y(new_n14311_));
  OAI21X1  g14247(.A0(new_n14310_), .A1(new_n14305_), .B0(new_n14311_), .Y(new_n14312_));
  NOR3X1   g14248(.A(new_n14311_), .B(new_n14310_), .C(new_n14305_), .Y(new_n14313_));
  AOI22X1  g14249(.A0(new_n12090_), .A1(new_n5970_), .B0(new_n12088_), .B1(new_n6300_), .Y(new_n14314_));
  OAI21X1  g14250(.A0(new_n12298_), .A1(new_n6309_), .B0(new_n14314_), .Y(new_n14315_));
  AOI21X1  g14251(.A0(new_n12297_), .A1(new_n5972_), .B0(new_n14315_), .Y(new_n14316_));
  XOR2X1   g14252(.A(new_n14316_), .B(\a[2] ), .Y(new_n14317_));
  OAI21X1  g14253(.A0(new_n14317_), .A1(new_n14313_), .B0(new_n14312_), .Y(new_n14318_));
  NAND2X1  g14254(.A(new_n14318_), .B(new_n14112_), .Y(new_n14319_));
  AOI22X1  g14255(.A0(new_n12088_), .A1(new_n5970_), .B0(new_n12085_), .B1(new_n6300_), .Y(new_n14320_));
  OAI21X1  g14256(.A0(new_n13321_), .A1(new_n6309_), .B0(new_n14320_), .Y(new_n14321_));
  AOI21X1  g14257(.A0(new_n13344_), .A1(new_n5972_), .B0(new_n14321_), .Y(new_n14322_));
  XOR2X1   g14258(.A(new_n14322_), .B(\a[2] ), .Y(new_n14323_));
  INVX1    g14259(.A(new_n14323_), .Y(new_n14324_));
  OAI21X1  g14260(.A0(new_n14318_), .A1(new_n14112_), .B0(new_n14324_), .Y(new_n14325_));
  OAI22X1  g14261(.A0(new_n12298_), .A1(new_n6325_), .B0(new_n13321_), .B1(new_n6307_), .Y(new_n14326_));
  AOI21X1  g14262(.A0(new_n12081_), .A1(new_n6308_), .B0(new_n14326_), .Y(new_n14327_));
  OAI21X1  g14263(.A0(new_n13335_), .A1(new_n6298_), .B0(new_n14327_), .Y(new_n14328_));
  XOR2X1   g14264(.A(new_n14328_), .B(new_n3431_), .Y(new_n14329_));
  NAND3X1  g14265(.A(new_n14329_), .B(new_n14325_), .C(new_n14319_), .Y(new_n14330_));
  XOR2X1   g14266(.A(new_n13949_), .B(new_n13743_), .Y(new_n14331_));
  INVX1    g14267(.A(new_n14331_), .Y(new_n14332_));
  AOI21X1  g14268(.A0(new_n14325_), .A1(new_n14319_), .B0(new_n14329_), .Y(new_n14333_));
  AOI21X1  g14269(.A0(new_n14332_), .A1(new_n14330_), .B0(new_n14333_), .Y(new_n14334_));
  OAI22X1  g14270(.A0(new_n13321_), .A1(new_n6325_), .B0(new_n13320_), .B1(new_n6307_), .Y(new_n14335_));
  AOI21X1  g14271(.A0(new_n12079_), .A1(new_n6308_), .B0(new_n14335_), .Y(new_n14336_));
  OAI21X1  g14272(.A0(new_n13325_), .A1(new_n6298_), .B0(new_n14336_), .Y(new_n14337_));
  XOR2X1   g14273(.A(new_n14337_), .B(new_n3431_), .Y(new_n14338_));
  XOR2X1   g14274(.A(new_n13950_), .B(new_n13735_), .Y(new_n14339_));
  INVX1    g14275(.A(new_n14339_), .Y(new_n14340_));
  AOI21X1  g14276(.A0(new_n14338_), .A1(new_n14334_), .B0(new_n14340_), .Y(new_n14341_));
  NOR2X1   g14277(.A(new_n14338_), .B(new_n14334_), .Y(new_n14342_));
  OAI22X1  g14278(.A0(new_n13320_), .A1(new_n6325_), .B0(new_n13665_), .B1(new_n6307_), .Y(new_n14343_));
  AOI21X1  g14279(.A0(new_n12076_), .A1(new_n6308_), .B0(new_n14343_), .Y(new_n14344_));
  OAI21X1  g14280(.A0(new_n13672_), .A1(new_n6298_), .B0(new_n14344_), .Y(new_n14345_));
  XOR2X1   g14281(.A(new_n14345_), .B(new_n3431_), .Y(new_n14346_));
  INVX1    g14282(.A(new_n14346_), .Y(new_n14347_));
  NOR3X1   g14283(.A(new_n14347_), .B(new_n14342_), .C(new_n14341_), .Y(new_n14348_));
  XOR2X1   g14284(.A(new_n13951_), .B(new_n13728_), .Y(new_n14349_));
  INVX1    g14285(.A(new_n14349_), .Y(new_n14350_));
  OAI21X1  g14286(.A0(new_n14342_), .A1(new_n14341_), .B0(new_n14347_), .Y(new_n14351_));
  OAI21X1  g14287(.A0(new_n14350_), .A1(new_n14348_), .B0(new_n14351_), .Y(new_n14352_));
  XOR2X1   g14288(.A(new_n13956_), .B(new_n13953_), .Y(new_n14353_));
  AND2X1   g14289(.A(new_n14353_), .B(new_n14352_), .Y(new_n14354_));
  AND2X1   g14290(.A(new_n14318_), .B(new_n14112_), .Y(new_n14355_));
  INVX1    g14291(.A(new_n14112_), .Y(new_n14356_));
  OR2X1    g14292(.A(new_n14304_), .B(new_n14302_), .Y(new_n14357_));
  OR2X1    g14293(.A(new_n14270_), .B(new_n14114_), .Y(new_n14358_));
  XOR2X1   g14294(.A(new_n13936_), .B(new_n13935_), .Y(new_n14359_));
  AND2X1   g14295(.A(new_n14254_), .B(new_n14253_), .Y(new_n14360_));
  AND2X1   g14296(.A(new_n14221_), .B(new_n14115_), .Y(new_n14361_));
  INVX1    g14297(.A(new_n14115_), .Y(new_n14362_));
  OR2X1    g14298(.A(new_n14204_), .B(new_n14202_), .Y(new_n14363_));
  OR2X1    g14299(.A(new_n14170_), .B(new_n14117_), .Y(new_n14364_));
  AND2X1   g14300(.A(new_n14156_), .B(new_n14123_), .Y(new_n14365_));
  OR4X1    g14301(.A(new_n14151_), .B(new_n14148_), .C(new_n14143_), .D(new_n14134_), .Y(new_n14366_));
  INVX1    g14302(.A(new_n14134_), .Y(new_n14367_));
  AOI21X1  g14303(.A0(new_n14141_), .A1(new_n14140_), .B0(\a[2] ), .Y(new_n14368_));
  NOR3X1   g14304(.A(new_n14138_), .B(new_n14136_), .C(new_n3431_), .Y(new_n14369_));
  OAI22X1  g14305(.A0(new_n14369_), .A1(new_n14368_), .B0(new_n14133_), .B1(new_n13894_), .Y(new_n14370_));
  OAI21X1  g14306(.A0(new_n14150_), .A1(new_n14149_), .B0(\a[2] ), .Y(new_n14371_));
  NAND3X1  g14307(.A(new_n14147_), .B(new_n14146_), .C(new_n3431_), .Y(new_n14372_));
  AOI22X1  g14308(.A0(new_n14372_), .A1(new_n14371_), .B0(new_n14370_), .B1(new_n14367_), .Y(new_n14373_));
  AOI21X1  g14309(.A0(new_n14153_), .A1(new_n14366_), .B0(new_n14373_), .Y(new_n14374_));
  XOR2X1   g14310(.A(new_n14160_), .B(\a[2] ), .Y(new_n14375_));
  AOI21X1  g14311(.A0(new_n14374_), .A1(new_n14122_), .B0(new_n14375_), .Y(new_n14376_));
  XOR2X1   g14312(.A(new_n14165_), .B(\a[2] ), .Y(new_n14377_));
  OAI21X1  g14313(.A0(new_n14376_), .A1(new_n14365_), .B0(new_n14377_), .Y(new_n14378_));
  NOR3X1   g14314(.A(new_n14377_), .B(new_n14376_), .C(new_n14365_), .Y(new_n14379_));
  INVX1    g14315(.A(new_n14169_), .Y(new_n14380_));
  OAI21X1  g14316(.A0(new_n14380_), .A1(new_n14379_), .B0(new_n14378_), .Y(new_n14381_));
  XOR2X1   g14317(.A(new_n14174_), .B(new_n3431_), .Y(new_n14382_));
  OAI21X1  g14318(.A0(new_n14381_), .A1(new_n14116_), .B0(new_n14382_), .Y(new_n14383_));
  XOR2X1   g14319(.A(new_n14179_), .B(new_n3431_), .Y(new_n14384_));
  NAND3X1  g14320(.A(new_n14384_), .B(new_n14383_), .C(new_n14364_), .Y(new_n14385_));
  AOI21X1  g14321(.A0(new_n14383_), .A1(new_n14364_), .B0(new_n14384_), .Y(new_n14386_));
  AOI21X1  g14322(.A0(new_n14182_), .A1(new_n14385_), .B0(new_n14386_), .Y(new_n14387_));
  XOR2X1   g14323(.A(new_n14188_), .B(new_n3431_), .Y(new_n14388_));
  INVX1    g14324(.A(new_n14190_), .Y(new_n14389_));
  AOI21X1  g14325(.A0(new_n14388_), .A1(new_n14387_), .B0(new_n14389_), .Y(new_n14390_));
  AND2X1   g14326(.A(new_n14189_), .B(new_n14185_), .Y(new_n14391_));
  XOR2X1   g14327(.A(new_n14197_), .B(\a[2] ), .Y(new_n14392_));
  NOR3X1   g14328(.A(new_n14392_), .B(new_n14391_), .C(new_n14390_), .Y(new_n14393_));
  INVX1    g14329(.A(new_n14200_), .Y(new_n14394_));
  OAI21X1  g14330(.A0(new_n14391_), .A1(new_n14390_), .B0(new_n14392_), .Y(new_n14395_));
  OAI21X1  g14331(.A0(new_n14394_), .A1(new_n14393_), .B0(new_n14395_), .Y(new_n14396_));
  INVX1    g14332(.A(new_n14209_), .Y(new_n14397_));
  OAI21X1  g14333(.A0(new_n14203_), .A1(new_n14396_), .B0(new_n14397_), .Y(new_n14398_));
  INVX1    g14334(.A(new_n14214_), .Y(new_n14399_));
  AOI21X1  g14335(.A0(new_n14398_), .A1(new_n14363_), .B0(new_n14399_), .Y(new_n14400_));
  NAND3X1  g14336(.A(new_n14399_), .B(new_n14398_), .C(new_n14363_), .Y(new_n14401_));
  INVX1    g14337(.A(new_n14220_), .Y(new_n14402_));
  AOI21X1  g14338(.A0(new_n14402_), .A1(new_n14401_), .B0(new_n14400_), .Y(new_n14403_));
  XOR2X1   g14339(.A(new_n14225_), .B(\a[2] ), .Y(new_n14404_));
  AOI21X1  g14340(.A0(new_n14403_), .A1(new_n14362_), .B0(new_n14404_), .Y(new_n14405_));
  XOR2X1   g14341(.A(new_n14230_), .B(\a[2] ), .Y(new_n14406_));
  NOR3X1   g14342(.A(new_n14406_), .B(new_n14405_), .C(new_n14361_), .Y(new_n14407_));
  INVX1    g14343(.A(new_n14233_), .Y(new_n14408_));
  OAI21X1  g14344(.A0(new_n14405_), .A1(new_n14361_), .B0(new_n14406_), .Y(new_n14409_));
  OAI21X1  g14345(.A0(new_n14408_), .A1(new_n14407_), .B0(new_n14409_), .Y(new_n14410_));
  INVX1    g14346(.A(new_n14239_), .Y(new_n14411_));
  OAI21X1  g14347(.A0(new_n14411_), .A1(new_n14410_), .B0(new_n14240_), .Y(new_n14412_));
  OR2X1    g14348(.A(new_n14239_), .B(new_n14235_), .Y(new_n14413_));
  NAND3X1  g14349(.A(new_n14247_), .B(new_n14413_), .C(new_n14412_), .Y(new_n14414_));
  AOI21X1  g14350(.A0(new_n14413_), .A1(new_n14412_), .B0(new_n14247_), .Y(new_n14415_));
  AOI21X1  g14351(.A0(new_n14250_), .A1(new_n14414_), .B0(new_n14415_), .Y(new_n14416_));
  INVX1    g14352(.A(new_n14254_), .Y(new_n14417_));
  AOI21X1  g14353(.A0(new_n14417_), .A1(new_n14416_), .B0(new_n14259_), .Y(new_n14418_));
  INVX1    g14354(.A(new_n14262_), .Y(new_n14419_));
  OAI21X1  g14355(.A0(new_n14418_), .A1(new_n14360_), .B0(new_n14419_), .Y(new_n14420_));
  NOR3X1   g14356(.A(new_n14419_), .B(new_n14418_), .C(new_n14360_), .Y(new_n14421_));
  OAI21X1  g14357(.A0(new_n14268_), .A1(new_n14421_), .B0(new_n14420_), .Y(new_n14422_));
  INVX1    g14358(.A(new_n14275_), .Y(new_n14423_));
  OAI21X1  g14359(.A0(new_n14422_), .A1(new_n14359_), .B0(new_n14423_), .Y(new_n14424_));
  NAND3X1  g14360(.A(new_n14280_), .B(new_n14424_), .C(new_n14358_), .Y(new_n14425_));
  AOI21X1  g14361(.A0(new_n14424_), .A1(new_n14358_), .B0(new_n14280_), .Y(new_n14426_));
  AOI21X1  g14362(.A0(new_n14283_), .A1(new_n14425_), .B0(new_n14426_), .Y(new_n14427_));
  INVX1    g14363(.A(new_n14292_), .Y(new_n14428_));
  AOI21X1  g14364(.A0(new_n14290_), .A1(new_n14427_), .B0(new_n14428_), .Y(new_n14429_));
  AND2X1   g14365(.A(new_n14291_), .B(new_n14286_), .Y(new_n14430_));
  INVX1    g14366(.A(new_n14298_), .Y(new_n14431_));
  NOR3X1   g14367(.A(new_n14431_), .B(new_n14430_), .C(new_n14429_), .Y(new_n14432_));
  INVX1    g14368(.A(new_n14300_), .Y(new_n14433_));
  OAI21X1  g14369(.A0(new_n14430_), .A1(new_n14429_), .B0(new_n14431_), .Y(new_n14434_));
  OAI21X1  g14370(.A0(new_n14433_), .A1(new_n14432_), .B0(new_n14434_), .Y(new_n14435_));
  INVX1    g14371(.A(new_n14309_), .Y(new_n14436_));
  OAI21X1  g14372(.A0(new_n14303_), .A1(new_n14435_), .B0(new_n14436_), .Y(new_n14437_));
  INVX1    g14373(.A(new_n14311_), .Y(new_n14438_));
  AOI21X1  g14374(.A0(new_n14437_), .A1(new_n14357_), .B0(new_n14438_), .Y(new_n14439_));
  NAND3X1  g14375(.A(new_n14438_), .B(new_n14437_), .C(new_n14357_), .Y(new_n14440_));
  INVX1    g14376(.A(new_n14317_), .Y(new_n14441_));
  AOI21X1  g14377(.A0(new_n14441_), .A1(new_n14440_), .B0(new_n14439_), .Y(new_n14442_));
  AOI21X1  g14378(.A0(new_n14442_), .A1(new_n14356_), .B0(new_n14323_), .Y(new_n14443_));
  INVX1    g14379(.A(new_n14329_), .Y(new_n14444_));
  NOR3X1   g14380(.A(new_n14444_), .B(new_n14443_), .C(new_n14355_), .Y(new_n14445_));
  OAI21X1  g14381(.A0(new_n14443_), .A1(new_n14355_), .B0(new_n14444_), .Y(new_n14446_));
  OAI21X1  g14382(.A0(new_n14331_), .A1(new_n14445_), .B0(new_n14446_), .Y(new_n14447_));
  INVX1    g14383(.A(new_n14338_), .Y(new_n14448_));
  OAI21X1  g14384(.A0(new_n14448_), .A1(new_n14447_), .B0(new_n14339_), .Y(new_n14449_));
  OR2X1    g14385(.A(new_n14338_), .B(new_n14334_), .Y(new_n14450_));
  NAND3X1  g14386(.A(new_n14346_), .B(new_n14450_), .C(new_n14449_), .Y(new_n14451_));
  AOI21X1  g14387(.A0(new_n14450_), .A1(new_n14449_), .B0(new_n14346_), .Y(new_n14452_));
  AOI21X1  g14388(.A0(new_n14349_), .A1(new_n14451_), .B0(new_n14452_), .Y(new_n14453_));
  INVX1    g14389(.A(new_n14353_), .Y(new_n14454_));
  AOI22X1  g14390(.A0(new_n12079_), .A1(new_n5970_), .B0(new_n12076_), .B1(new_n6300_), .Y(new_n14455_));
  OAI21X1  g14391(.A0(new_n13691_), .A1(new_n6309_), .B0(new_n14455_), .Y(new_n14456_));
  AOI21X1  g14392(.A0(new_n13690_), .A1(new_n5972_), .B0(new_n14456_), .Y(new_n14457_));
  XOR2X1   g14393(.A(new_n14457_), .B(\a[2] ), .Y(new_n14458_));
  AOI21X1  g14394(.A0(new_n14454_), .A1(new_n14453_), .B0(new_n14458_), .Y(new_n14459_));
  OAI21X1  g14395(.A0(new_n14459_), .A1(new_n14354_), .B0(new_n14111_), .Y(new_n14460_));
  NOR3X1   g14396(.A(new_n14459_), .B(new_n14354_), .C(new_n14111_), .Y(new_n14461_));
  AOI22X1  g14397(.A0(new_n12076_), .A1(new_n5970_), .B0(new_n12018_), .B1(new_n6300_), .Y(new_n14462_));
  OAI21X1  g14398(.A0(new_n13679_), .A1(new_n6309_), .B0(new_n14462_), .Y(new_n14463_));
  AOI21X1  g14399(.A0(new_n13678_), .A1(new_n5972_), .B0(new_n14463_), .Y(new_n14464_));
  XOR2X1   g14400(.A(new_n14464_), .B(\a[2] ), .Y(new_n14465_));
  OAI21X1  g14401(.A0(new_n14465_), .A1(new_n14461_), .B0(new_n14460_), .Y(new_n14466_));
  INVX1    g14402(.A(new_n12291_), .Y(new_n14467_));
  OAI22X1  g14403(.A0(new_n13679_), .A1(new_n6307_), .B0(new_n13691_), .B1(new_n6325_), .Y(new_n14468_));
  AOI21X1  g14404(.A0(new_n12285_), .A1(new_n6308_), .B0(new_n14468_), .Y(new_n14469_));
  OAI21X1  g14405(.A0(new_n14467_), .A1(new_n6298_), .B0(new_n14469_), .Y(new_n14470_));
  XOR2X1   g14406(.A(new_n14470_), .B(new_n3431_), .Y(new_n14471_));
  INVX1    g14407(.A(new_n14471_), .Y(new_n14472_));
  XOR2X1   g14408(.A(new_n13961_), .B(new_n13708_), .Y(new_n14473_));
  OAI21X1  g14409(.A0(new_n14472_), .A1(new_n14466_), .B0(new_n14473_), .Y(new_n14474_));
  NAND2X1  g14410(.A(new_n14472_), .B(new_n14466_), .Y(new_n14475_));
  OAI22X1  g14411(.A0(new_n12292_), .A1(new_n6307_), .B0(new_n13679_), .B1(new_n6325_), .Y(new_n14476_));
  AOI21X1  g14412(.A0(new_n14085_), .A1(new_n6308_), .B0(new_n14476_), .Y(new_n14477_));
  INVX1    g14413(.A(new_n14096_), .Y(new_n14478_));
  OAI21X1  g14414(.A0(new_n14094_), .A1(new_n14093_), .B0(new_n12290_), .Y(new_n14479_));
  OAI21X1  g14415(.A0(new_n14478_), .A1(new_n14094_), .B0(new_n14479_), .Y(new_n14480_));
  INVX1    g14416(.A(new_n14480_), .Y(new_n14481_));
  OAI21X1  g14417(.A0(new_n14481_), .A1(new_n6298_), .B0(new_n14477_), .Y(new_n14482_));
  XOR2X1   g14418(.A(new_n14482_), .B(new_n3431_), .Y(new_n14483_));
  NAND3X1  g14419(.A(new_n14483_), .B(new_n14475_), .C(new_n14474_), .Y(new_n14484_));
  XOR2X1   g14420(.A(new_n13962_), .B(new_n13698_), .Y(new_n14485_));
  AOI21X1  g14421(.A0(new_n14475_), .A1(new_n14474_), .B0(new_n14483_), .Y(new_n14486_));
  AOI21X1  g14422(.A0(new_n14485_), .A1(new_n14484_), .B0(new_n14486_), .Y(new_n14487_));
  OAI22X1  g14423(.A0(new_n14086_), .A1(new_n6307_), .B0(new_n12292_), .B1(new_n6325_), .Y(new_n14488_));
  AOI21X1  g14424(.A0(new_n14087_), .A1(new_n6308_), .B0(new_n14488_), .Y(new_n14489_));
  XOR2X1   g14425(.A(new_n14087_), .B(new_n14085_), .Y(new_n14490_));
  OAI22X1  g14426(.A0(new_n14098_), .A1(new_n14097_), .B0(new_n14490_), .B1(new_n14096_), .Y(new_n14491_));
  INVX1    g14427(.A(new_n14491_), .Y(new_n14492_));
  OAI21X1  g14428(.A0(new_n14492_), .A1(new_n6298_), .B0(new_n14489_), .Y(new_n14493_));
  XOR2X1   g14429(.A(new_n14493_), .B(new_n3431_), .Y(new_n14494_));
  INVX1    g14430(.A(new_n13687_), .Y(new_n14495_));
  XOR2X1   g14431(.A(new_n13964_), .B(new_n14495_), .Y(new_n14496_));
  AOI21X1  g14432(.A0(new_n14494_), .A1(new_n14487_), .B0(new_n14496_), .Y(new_n14497_));
  NOR2X1   g14433(.A(new_n14494_), .B(new_n14487_), .Y(new_n14498_));
  XOR2X1   g14434(.A(new_n14109_), .B(new_n13966_), .Y(new_n14499_));
  OAI21X1  g14435(.A0(new_n14498_), .A1(new_n14497_), .B0(new_n14499_), .Y(new_n14500_));
  NAND2X1  g14436(.A(new_n14500_), .B(new_n14110_), .Y(new_n14501_));
  AOI22X1  g14437(.A0(new_n12285_), .A1(new_n5659_), .B0(new_n12074_), .B1(new_n5373_), .Y(new_n14502_));
  OAI21X1  g14438(.A0(new_n14086_), .A1(new_n5959_), .B0(new_n14502_), .Y(new_n14503_));
  AOI21X1  g14439(.A0(new_n14480_), .A1(new_n67_), .B0(new_n14503_), .Y(new_n14504_));
  XOR2X1   g14440(.A(new_n14504_), .B(\a[5] ), .Y(new_n14505_));
  XOR2X1   g14441(.A(new_n13673_), .B(\a[8] ), .Y(new_n14506_));
  AND2X1   g14442(.A(new_n14506_), .B(new_n13664_), .Y(new_n14507_));
  INVX1    g14443(.A(new_n13675_), .Y(new_n14508_));
  AOI21X1  g14444(.A0(new_n14508_), .A1(new_n13579_), .B0(new_n14507_), .Y(new_n14509_));
  INVX1    g14445(.A(new_n13335_), .Y(new_n14510_));
  AOI22X1  g14446(.A0(new_n12085_), .A1(new_n4078_), .B0(new_n12083_), .B1(new_n4247_), .Y(new_n14511_));
  OAI21X1  g14447(.A0(new_n13320_), .A1(new_n4427_), .B0(new_n14511_), .Y(new_n14512_));
  AOI21X1  g14448(.A0(new_n14510_), .A1(new_n4080_), .B0(new_n14512_), .Y(new_n14513_));
  XOR2X1   g14449(.A(new_n14513_), .B(\a[11] ), .Y(new_n14514_));
  XOR2X1   g14450(.A(new_n13655_), .B(\a[14] ), .Y(new_n14515_));
  AND2X1   g14451(.A(new_n14515_), .B(new_n13652_), .Y(new_n14516_));
  AOI21X1  g14452(.A0(new_n13587_), .A1(new_n13586_), .B0(new_n13657_), .Y(new_n14517_));
  NOR2X1   g14453(.A(new_n14517_), .B(new_n14516_), .Y(new_n14518_));
  INVX1    g14454(.A(new_n12846_), .Y(new_n14519_));
  AOI22X1  g14455(.A0(new_n12099_), .A1(new_n3232_), .B0(new_n12097_), .B1(new_n3390_), .Y(new_n14520_));
  OAI21X1  g14456(.A0(new_n13090_), .A1(new_n3545_), .B0(new_n14520_), .Y(new_n14521_));
  AOI21X1  g14457(.A0(new_n14519_), .A1(new_n3234_), .B0(new_n14521_), .Y(new_n14522_));
  XOR2X1   g14458(.A(new_n14522_), .B(\a[17] ), .Y(new_n14523_));
  INVX1    g14459(.A(new_n13596_), .Y(new_n14524_));
  AND2X1   g14460(.A(new_n13641_), .B(new_n13638_), .Y(new_n14525_));
  NOR2X1   g14461(.A(new_n13641_), .B(new_n13638_), .Y(new_n14526_));
  NOR3X1   g14462(.A(new_n13646_), .B(new_n14526_), .C(new_n14525_), .Y(new_n14527_));
  INVX1    g14463(.A(new_n14527_), .Y(new_n14528_));
  OAI21X1  g14464(.A0(new_n13647_), .A1(new_n14524_), .B0(new_n14528_), .Y(new_n14529_));
  NOR2X1   g14465(.A(new_n12685_), .B(new_n2692_), .Y(new_n14530_));
  AOI22X1  g14466(.A0(new_n12720_), .A1(new_n2657_), .B0(new_n12516_), .B1(new_n2696_), .Y(new_n14531_));
  OAI21X1  g14467(.A0(new_n12111_), .A1(new_n2753_), .B0(new_n14531_), .Y(new_n14532_));
  NOR2X1   g14468(.A(new_n14532_), .B(new_n14530_), .Y(new_n14533_));
  XOR2X1   g14469(.A(new_n14533_), .B(\a[23] ), .Y(new_n14534_));
  XOR2X1   g14470(.A(new_n13634_), .B(new_n89_), .Y(new_n14535_));
  AND2X1   g14471(.A(new_n14535_), .B(new_n13631_), .Y(new_n14536_));
  INVX1    g14472(.A(new_n14536_), .Y(new_n14537_));
  OAI21X1  g14473(.A0(new_n13636_), .A1(new_n13606_), .B0(new_n14537_), .Y(new_n14538_));
  INVX1    g14474(.A(new_n14538_), .Y(new_n14539_));
  INVX1    g14475(.A(new_n12453_), .Y(new_n14540_));
  AOI22X1  g14476(.A0(new_n12151_), .A1(new_n2185_), .B0(new_n12148_), .B1(new_n2095_), .Y(new_n14541_));
  OAI21X1  g14477(.A0(new_n12192_), .A1(new_n2140_), .B0(new_n14541_), .Y(new_n14542_));
  AOI21X1  g14478(.A0(new_n14540_), .A1(new_n2062_), .B0(new_n14542_), .Y(new_n14543_));
  XOR2X1   g14479(.A(new_n14543_), .B(\a[29] ), .Y(new_n14544_));
  INVX1    g14480(.A(new_n13620_), .Y(new_n14545_));
  NOR2X1   g14481(.A(new_n13623_), .B(new_n14545_), .Y(new_n14546_));
  INVX1    g14482(.A(new_n14546_), .Y(new_n14547_));
  OAI21X1  g14483(.A0(new_n13624_), .A1(new_n13613_), .B0(new_n14547_), .Y(new_n14548_));
  NOR2X1   g14484(.A(new_n489_), .B(new_n465_), .Y(new_n14549_));
  NOR3X1   g14485(.A(new_n835_), .B(new_n843_), .C(new_n981_), .Y(new_n14550_));
  NAND3X1  g14486(.A(new_n14550_), .B(new_n14549_), .C(new_n2801_), .Y(new_n14551_));
  OR4X1    g14487(.A(new_n1082_), .B(new_n232_), .C(new_n226_), .D(new_n522_), .Y(new_n14552_));
  OR4X1    g14488(.A(new_n14552_), .B(new_n1342_), .C(new_n1057_), .D(new_n154_), .Y(new_n14553_));
  NOR4X1   g14489(.A(new_n14553_), .B(new_n14551_), .C(new_n7375_), .D(new_n1976_), .Y(new_n14554_));
  NAND3X1  g14490(.A(new_n14554_), .B(new_n7434_), .C(new_n2546_), .Y(new_n14555_));
  AOI22X1  g14491(.A0(new_n12162_), .A1(new_n1890_), .B0(new_n12158_), .B1(new_n1884_), .Y(new_n14556_));
  OAI21X1  g14492(.A0(new_n12353_), .A1(new_n3498_), .B0(new_n14556_), .Y(new_n14557_));
  AOI21X1  g14493(.A0(new_n12352_), .A1(new_n407_), .B0(new_n14557_), .Y(new_n14558_));
  XOR2X1   g14494(.A(new_n14558_), .B(new_n14555_), .Y(new_n14559_));
  XOR2X1   g14495(.A(new_n14559_), .B(new_n14548_), .Y(new_n14560_));
  XOR2X1   g14496(.A(new_n14560_), .B(new_n14544_), .Y(new_n14561_));
  INVX1    g14497(.A(new_n14561_), .Y(new_n14562_));
  OR2X1    g14498(.A(new_n13626_), .B(new_n13610_), .Y(new_n14563_));
  OR2X1    g14499(.A(new_n13630_), .B(new_n13628_), .Y(new_n14564_));
  AND2X1   g14500(.A(new_n14564_), .B(new_n14563_), .Y(new_n14565_));
  XOR2X1   g14501(.A(new_n14565_), .B(new_n14562_), .Y(new_n14566_));
  INVX1    g14502(.A(new_n12536_), .Y(new_n14567_));
  OAI22X1  g14503(.A0(new_n14194_), .A1(new_n2666_), .B0(new_n12314_), .B1(new_n2419_), .Y(new_n14568_));
  AOI21X1  g14504(.A0(new_n12133_), .A1(new_n2423_), .B0(new_n14568_), .Y(new_n14569_));
  OAI21X1  g14505(.A0(new_n14567_), .A1(new_n2665_), .B0(new_n14569_), .Y(new_n14570_));
  XOR2X1   g14506(.A(new_n14570_), .B(new_n89_), .Y(new_n14571_));
  XOR2X1   g14507(.A(new_n14571_), .B(new_n14566_), .Y(new_n14572_));
  XOR2X1   g14508(.A(new_n14572_), .B(new_n14539_), .Y(new_n14573_));
  XOR2X1   g14509(.A(new_n14573_), .B(new_n14534_), .Y(new_n14574_));
  INVX1    g14510(.A(new_n13600_), .Y(new_n14575_));
  AOI21X1  g14511(.A0(new_n13637_), .A1(new_n14575_), .B0(new_n14526_), .Y(new_n14576_));
  XOR2X1   g14512(.A(new_n14576_), .B(new_n14574_), .Y(new_n14577_));
  INVX1    g14513(.A(new_n12305_), .Y(new_n14578_));
  OAI22X1  g14514(.A0(new_n12109_), .A1(new_n3250_), .B0(new_n12695_), .B1(new_n3144_), .Y(new_n14579_));
  AOI21X1  g14515(.A0(new_n12102_), .A1(new_n3146_), .B0(new_n14579_), .Y(new_n14580_));
  OAI21X1  g14516(.A0(new_n14578_), .A1(new_n3098_), .B0(new_n14580_), .Y(new_n14581_));
  XOR2X1   g14517(.A(new_n14581_), .B(new_n1920_), .Y(new_n14582_));
  XOR2X1   g14518(.A(new_n14582_), .B(new_n14577_), .Y(new_n14583_));
  XOR2X1   g14519(.A(new_n14583_), .B(new_n14529_), .Y(new_n14584_));
  XOR2X1   g14520(.A(new_n14584_), .B(new_n14523_), .Y(new_n14585_));
  INVX1    g14521(.A(new_n14585_), .Y(new_n14586_));
  NOR2X1   g14522(.A(new_n13648_), .B(new_n13592_), .Y(new_n14587_));
  AOI21X1  g14523(.A0(new_n13651_), .A1(new_n13649_), .B0(new_n14587_), .Y(new_n14588_));
  XOR2X1   g14524(.A(new_n14588_), .B(new_n14586_), .Y(new_n14589_));
  INVX1    g14525(.A(new_n13103_), .Y(new_n14590_));
  OAI22X1  g14526(.A0(new_n13366_), .A1(new_n3627_), .B0(new_n13118_), .B1(new_n3907_), .Y(new_n14591_));
  AOI21X1  g14527(.A0(new_n12088_), .A1(new_n3984_), .B0(new_n14591_), .Y(new_n14592_));
  OAI21X1  g14528(.A0(new_n14590_), .A1(new_n3906_), .B0(new_n14592_), .Y(new_n14593_));
  XOR2X1   g14529(.A(new_n14593_), .B(new_n2529_), .Y(new_n14594_));
  XOR2X1   g14530(.A(new_n14594_), .B(new_n14589_), .Y(new_n14595_));
  INVX1    g14531(.A(new_n14595_), .Y(new_n14596_));
  XOR2X1   g14532(.A(new_n14596_), .B(new_n14518_), .Y(new_n14597_));
  XOR2X1   g14533(.A(new_n14597_), .B(new_n14514_), .Y(new_n14598_));
  INVX1    g14534(.A(new_n14598_), .Y(new_n14599_));
  NOR2X1   g14535(.A(new_n13659_), .B(new_n13583_), .Y(new_n14600_));
  INVX1    g14536(.A(new_n13663_), .Y(new_n14601_));
  AOI21X1  g14537(.A0(new_n14601_), .A1(new_n13660_), .B0(new_n14600_), .Y(new_n14602_));
  XOR2X1   g14538(.A(new_n14602_), .B(new_n14599_), .Y(new_n14603_));
  INVX1    g14539(.A(new_n13690_), .Y(new_n14604_));
  OAI22X1  g14540(.A0(new_n13665_), .A1(new_n4634_), .B0(new_n13700_), .B1(new_n4869_), .Y(new_n14605_));
  AOI21X1  g14541(.A0(new_n12018_), .A1(new_n5097_), .B0(new_n14605_), .Y(new_n14606_));
  OAI21X1  g14542(.A0(new_n14604_), .A1(new_n4868_), .B0(new_n14606_), .Y(new_n14607_));
  XOR2X1   g14543(.A(new_n14607_), .B(new_n2995_), .Y(new_n14608_));
  XOR2X1   g14544(.A(new_n14608_), .B(new_n14603_), .Y(new_n14609_));
  INVX1    g14545(.A(new_n14609_), .Y(new_n14610_));
  XOR2X1   g14546(.A(new_n14610_), .B(new_n14509_), .Y(new_n14611_));
  XOR2X1   g14547(.A(new_n14611_), .B(new_n14505_), .Y(new_n14612_));
  INVX1    g14548(.A(new_n13677_), .Y(new_n14613_));
  OR2X1    g14549(.A(new_n13965_), .B(new_n14613_), .Y(new_n14614_));
  OAI21X1  g14550(.A0(new_n13676_), .A1(new_n12296_), .B0(new_n14614_), .Y(new_n14615_));
  XOR2X1   g14551(.A(new_n14615_), .B(new_n14612_), .Y(new_n14616_));
  NOR2X1   g14552(.A(new_n14082_), .B(new_n14079_), .Y(new_n14617_));
  AOI21X1  g14553(.A0(new_n14083_), .A1(new_n14054_), .B0(new_n14617_), .Y(new_n14618_));
  NOR2X1   g14554(.A(new_n14072_), .B(new_n14068_), .Y(new_n14619_));
  INVX1    g14555(.A(new_n14619_), .Y(new_n14620_));
  OAI21X1  g14556(.A0(new_n14077_), .A1(new_n14074_), .B0(new_n14620_), .Y(new_n14621_));
  AOI22X1  g14557(.A0(new_n7578_), .A1(new_n1884_), .B0(new_n7571_), .B1(new_n1890_), .Y(new_n14622_));
  OAI21X1  g14558(.A0(new_n7594_), .A1(new_n3498_), .B0(new_n14622_), .Y(new_n14623_));
  AOI21X1  g14559(.A0(new_n7593_), .A1(new_n407_), .B0(new_n14623_), .Y(new_n14624_));
  NAND2X1  g14560(.A(new_n14062_), .B(new_n14057_), .Y(new_n14625_));
  OAI21X1  g14561(.A0(new_n14061_), .A1(new_n13985_), .B0(new_n14625_), .Y(new_n14626_));
  NOR4X1   g14562(.A(new_n14059_), .B(new_n2646_), .C(new_n2345_), .D(new_n460_), .Y(new_n14627_));
  XOR2X1   g14563(.A(new_n14627_), .B(new_n14626_), .Y(new_n14628_));
  XOR2X1   g14564(.A(new_n14628_), .B(new_n14624_), .Y(new_n14629_));
  INVX1    g14565(.A(new_n14629_), .Y(new_n14630_));
  INVX1    g14566(.A(new_n14064_), .Y(new_n14631_));
  NOR2X1   g14567(.A(new_n14067_), .B(new_n14631_), .Y(new_n14632_));
  AOI21X1  g14568(.A0(new_n14063_), .A1(new_n14019_), .B0(new_n14632_), .Y(new_n14633_));
  XOR2X1   g14569(.A(new_n14633_), .B(new_n14630_), .Y(new_n14634_));
  OAI22X1  g14570(.A0(new_n7642_), .A1(new_n2186_), .B0(new_n8172_), .B1(new_n2140_), .Y(new_n14635_));
  AOI21X1  g14571(.A0(new_n7643_), .A1(new_n2095_), .B0(new_n14635_), .Y(new_n14636_));
  OAI21X1  g14572(.A0(new_n7655_), .A1(new_n2063_), .B0(new_n14636_), .Y(new_n14637_));
  XOR2X1   g14573(.A(new_n14637_), .B(new_n74_), .Y(new_n14638_));
  XOR2X1   g14574(.A(new_n14638_), .B(new_n14634_), .Y(new_n14639_));
  XOR2X1   g14575(.A(new_n14639_), .B(new_n14621_), .Y(new_n14640_));
  INVX1    g14576(.A(new_n14640_), .Y(new_n14641_));
  XOR2X1   g14577(.A(new_n14641_), .B(new_n14618_), .Y(new_n14642_));
  INVX1    g14578(.A(new_n14084_), .Y(new_n14643_));
  OAI22X1  g14579(.A0(new_n14088_), .A1(new_n6325_), .B0(new_n14643_), .B1(new_n6307_), .Y(new_n14644_));
  AOI21X1  g14580(.A0(new_n14642_), .A1(new_n6308_), .B0(new_n14644_), .Y(new_n14645_));
  NOR2X1   g14581(.A(new_n14642_), .B(new_n14084_), .Y(new_n14646_));
  XOR2X1   g14582(.A(new_n14642_), .B(new_n14084_), .Y(new_n14647_));
  INVX1    g14583(.A(new_n14642_), .Y(new_n14648_));
  NAND2X1  g14584(.A(new_n14647_), .B(new_n14105_), .Y(new_n14649_));
  OAI21X1  g14585(.A0(new_n14648_), .A1(new_n14643_), .B0(new_n14649_), .Y(new_n14650_));
  OAI22X1  g14586(.A0(new_n14650_), .A1(new_n14646_), .B0(new_n14647_), .B1(new_n14104_), .Y(new_n14651_));
  INVX1    g14587(.A(new_n14651_), .Y(new_n14652_));
  OAI21X1  g14588(.A0(new_n14652_), .A1(new_n6298_), .B0(new_n14645_), .Y(new_n14653_));
  XOR2X1   g14589(.A(new_n14653_), .B(new_n3431_), .Y(new_n14654_));
  XOR2X1   g14590(.A(new_n14654_), .B(new_n14616_), .Y(new_n14655_));
  XOR2X1   g14591(.A(new_n14655_), .B(new_n14501_), .Y(new_n14656_));
  NOR2X1   g14592(.A(new_n14498_), .B(new_n14497_), .Y(new_n14657_));
  XOR2X1   g14593(.A(new_n14499_), .B(new_n14657_), .Y(new_n14658_));
  XOR2X1   g14594(.A(new_n14658_), .B(new_n14656_), .Y(\result[0] ));
  NOR2X1   g14595(.A(new_n14658_), .B(new_n14656_), .Y(new_n14660_));
  XOR2X1   g14596(.A(new_n14653_), .B(\a[2] ), .Y(new_n14661_));
  AND2X1   g14597(.A(new_n14661_), .B(new_n14616_), .Y(new_n14662_));
  AOI21X1  g14598(.A0(new_n14500_), .A1(new_n14110_), .B0(new_n14655_), .Y(new_n14663_));
  OR2X1    g14599(.A(new_n14663_), .B(new_n14662_), .Y(new_n14664_));
  AOI22X1  g14600(.A0(new_n14085_), .A1(new_n5659_), .B0(new_n12285_), .B1(new_n5373_), .Y(new_n14665_));
  OAI21X1  g14601(.A0(new_n14088_), .A1(new_n5959_), .B0(new_n14665_), .Y(new_n14666_));
  AOI21X1  g14602(.A0(new_n14491_), .A1(new_n67_), .B0(new_n14666_), .Y(new_n14667_));
  XOR2X1   g14603(.A(new_n14667_), .B(\a[5] ), .Y(new_n14668_));
  INVX1    g14604(.A(new_n14603_), .Y(new_n14669_));
  OR2X1    g14605(.A(new_n14609_), .B(new_n14509_), .Y(new_n14670_));
  OAI21X1  g14606(.A0(new_n14608_), .A1(new_n14669_), .B0(new_n14670_), .Y(new_n14671_));
  INVX1    g14607(.A(new_n13325_), .Y(new_n14672_));
  AOI22X1  g14608(.A0(new_n12083_), .A1(new_n4078_), .B0(new_n12081_), .B1(new_n4247_), .Y(new_n14673_));
  OAI21X1  g14609(.A0(new_n13665_), .A1(new_n4427_), .B0(new_n14673_), .Y(new_n14674_));
  AOI21X1  g14610(.A0(new_n14672_), .A1(new_n4080_), .B0(new_n14674_), .Y(new_n14675_));
  XOR2X1   g14611(.A(new_n14675_), .B(\a[11] ), .Y(new_n14676_));
  XOR2X1   g14612(.A(new_n14593_), .B(\a[14] ), .Y(new_n14677_));
  AND2X1   g14613(.A(new_n14677_), .B(new_n14589_), .Y(new_n14678_));
  INVX1    g14614(.A(new_n14678_), .Y(new_n14679_));
  OAI21X1  g14615(.A0(new_n14517_), .A1(new_n14516_), .B0(new_n14596_), .Y(new_n14680_));
  AND2X1   g14616(.A(new_n14680_), .B(new_n14679_), .Y(new_n14681_));
  AOI22X1  g14617(.A0(new_n12097_), .A1(new_n3232_), .B0(new_n12095_), .B1(new_n3390_), .Y(new_n14682_));
  OAI21X1  g14618(.A0(new_n13366_), .A1(new_n3545_), .B0(new_n14682_), .Y(new_n14683_));
  AOI21X1  g14619(.A0(new_n13093_), .A1(new_n3234_), .B0(new_n14683_), .Y(new_n14684_));
  XOR2X1   g14620(.A(new_n14684_), .B(\a[17] ), .Y(new_n14685_));
  INVX1    g14621(.A(new_n14529_), .Y(new_n14686_));
  AND2X1   g14622(.A(new_n14576_), .B(new_n14574_), .Y(new_n14687_));
  NOR2X1   g14623(.A(new_n14576_), .B(new_n14574_), .Y(new_n14688_));
  NOR3X1   g14624(.A(new_n14582_), .B(new_n14688_), .C(new_n14687_), .Y(new_n14689_));
  INVX1    g14625(.A(new_n14689_), .Y(new_n14690_));
  OAI21X1  g14626(.A0(new_n14583_), .A1(new_n14686_), .B0(new_n14690_), .Y(new_n14691_));
  OAI22X1  g14627(.A0(new_n12113_), .A1(new_n4016_), .B0(new_n12111_), .B1(new_n2743_), .Y(new_n14692_));
  AOI21X1  g14628(.A0(new_n12107_), .A1(new_n2745_), .B0(new_n14692_), .Y(new_n14693_));
  OAI21X1  g14629(.A0(new_n12708_), .A1(new_n2692_), .B0(new_n14693_), .Y(new_n14694_));
  XOR2X1   g14630(.A(new_n14694_), .B(new_n70_), .Y(new_n14695_));
  XOR2X1   g14631(.A(new_n14570_), .B(\a[26] ), .Y(new_n14696_));
  AND2X1   g14632(.A(new_n14696_), .B(new_n14566_), .Y(new_n14697_));
  INVX1    g14633(.A(new_n14697_), .Y(new_n14698_));
  OAI21X1  g14634(.A0(new_n14572_), .A1(new_n14539_), .B0(new_n14698_), .Y(new_n14699_));
  NOR2X1   g14635(.A(new_n14560_), .B(new_n14544_), .Y(new_n14700_));
  OAI21X1  g14636(.A0(new_n13630_), .A1(new_n13628_), .B0(new_n14563_), .Y(new_n14701_));
  AOI21X1  g14637(.A0(new_n14701_), .A1(new_n14561_), .B0(new_n14700_), .Y(new_n14702_));
  INVX1    g14638(.A(new_n14702_), .Y(new_n14703_));
  INVX1    g14639(.A(new_n14548_), .Y(new_n14704_));
  INVX1    g14640(.A(new_n14555_), .Y(new_n14705_));
  NOR2X1   g14641(.A(new_n14558_), .B(new_n14705_), .Y(new_n14706_));
  INVX1    g14642(.A(new_n14706_), .Y(new_n14707_));
  OAI21X1  g14643(.A0(new_n14559_), .A1(new_n14704_), .B0(new_n14707_), .Y(new_n14708_));
  OR4X1    g14644(.A(new_n2089_), .B(new_n1224_), .C(new_n740_), .D(new_n227_), .Y(new_n14709_));
  OR4X1    g14645(.A(new_n220_), .B(new_n648_), .C(new_n746_), .D(new_n1008_), .Y(new_n14710_));
  OR4X1    g14646(.A(new_n14710_), .B(new_n14709_), .C(new_n1136_), .D(new_n1057_), .Y(new_n14711_));
  OR4X1    g14647(.A(new_n848_), .B(new_n510_), .C(new_n819_), .D(new_n400_), .Y(new_n14712_));
  OR4X1    g14648(.A(new_n14712_), .B(new_n2154_), .C(new_n1412_), .D(new_n891_), .Y(new_n14713_));
  OR4X1    g14649(.A(new_n14713_), .B(new_n14711_), .C(new_n3803_), .D(new_n3727_), .Y(new_n14714_));
  NOR4X1   g14650(.A(new_n14714_), .B(new_n7930_), .C(new_n1854_), .D(new_n1611_), .Y(new_n14715_));
  INVX1    g14651(.A(new_n14715_), .Y(new_n14716_));
  AOI22X1  g14652(.A0(new_n12158_), .A1(new_n1890_), .B0(new_n12155_), .B1(new_n1884_), .Y(new_n14717_));
  OAI21X1  g14653(.A0(new_n12322_), .A1(new_n3498_), .B0(new_n14717_), .Y(new_n14718_));
  AOI21X1  g14654(.A0(new_n12321_), .A1(new_n407_), .B0(new_n14718_), .Y(new_n14719_));
  XOR2X1   g14655(.A(new_n14719_), .B(new_n14716_), .Y(new_n14720_));
  XOR2X1   g14656(.A(new_n14720_), .B(new_n14708_), .Y(new_n14721_));
  OAI22X1  g14657(.A0(new_n12186_), .A1(new_n2186_), .B0(new_n12192_), .B1(new_n2431_), .Y(new_n14722_));
  AOI21X1  g14658(.A0(new_n12141_), .A1(new_n2139_), .B0(new_n14722_), .Y(new_n14723_));
  OAI21X1  g14659(.A0(new_n12444_), .A1(new_n2063_), .B0(new_n14723_), .Y(new_n14724_));
  XOR2X1   g14660(.A(new_n14724_), .B(new_n74_), .Y(new_n14725_));
  XOR2X1   g14661(.A(new_n14725_), .B(new_n14721_), .Y(new_n14726_));
  XOR2X1   g14662(.A(new_n14726_), .B(new_n14703_), .Y(new_n14727_));
  AOI22X1  g14663(.A0(new_n12138_), .A1(new_n2424_), .B0(new_n12133_), .B1(new_n2418_), .Y(new_n14728_));
  OAI21X1  g14664(.A0(new_n12117_), .A1(new_n2626_), .B0(new_n14728_), .Y(new_n14729_));
  AOI21X1  g14665(.A0(new_n12526_), .A1(new_n2301_), .B0(new_n14729_), .Y(new_n14730_));
  XOR2X1   g14666(.A(new_n14730_), .B(\a[26] ), .Y(new_n14731_));
  XOR2X1   g14667(.A(new_n14731_), .B(new_n14727_), .Y(new_n14732_));
  XOR2X1   g14668(.A(new_n14732_), .B(new_n14699_), .Y(new_n14733_));
  XOR2X1   g14669(.A(new_n14733_), .B(new_n14695_), .Y(new_n14734_));
  INVX1    g14670(.A(new_n14734_), .Y(new_n14735_));
  INVX1    g14671(.A(new_n14534_), .Y(new_n14736_));
  AOI21X1  g14672(.A0(new_n14573_), .A1(new_n14736_), .B0(new_n14688_), .Y(new_n14737_));
  XOR2X1   g14673(.A(new_n14737_), .B(new_n14735_), .Y(new_n14738_));
  AOI22X1  g14674(.A0(new_n12104_), .A1(new_n2875_), .B0(new_n12102_), .B1(new_n3099_), .Y(new_n14739_));
  OAI21X1  g14675(.A0(new_n12840_), .A1(new_n3152_), .B0(new_n14739_), .Y(new_n14740_));
  AOI21X1  g14676(.A0(new_n12859_), .A1(new_n2876_), .B0(new_n14740_), .Y(new_n14741_));
  XOR2X1   g14677(.A(new_n14741_), .B(\a[20] ), .Y(new_n14742_));
  XOR2X1   g14678(.A(new_n14742_), .B(new_n14738_), .Y(new_n14743_));
  XOR2X1   g14679(.A(new_n14743_), .B(new_n14691_), .Y(new_n14744_));
  XOR2X1   g14680(.A(new_n14744_), .B(new_n14685_), .Y(new_n14745_));
  NOR2X1   g14681(.A(new_n14584_), .B(new_n14523_), .Y(new_n14746_));
  INVX1    g14682(.A(new_n14746_), .Y(new_n14747_));
  OAI21X1  g14683(.A0(new_n14588_), .A1(new_n14586_), .B0(new_n14747_), .Y(new_n14748_));
  XOR2X1   g14684(.A(new_n14748_), .B(new_n14745_), .Y(new_n14749_));
  AOI22X1  g14685(.A0(new_n12090_), .A1(new_n3628_), .B0(new_n12088_), .B1(new_n3908_), .Y(new_n14750_));
  OAI21X1  g14686(.A0(new_n12298_), .A1(new_n3983_), .B0(new_n14750_), .Y(new_n14751_));
  AOI21X1  g14687(.A0(new_n12297_), .A1(new_n3624_), .B0(new_n14751_), .Y(new_n14752_));
  XOR2X1   g14688(.A(new_n14752_), .B(\a[14] ), .Y(new_n14753_));
  XOR2X1   g14689(.A(new_n14753_), .B(new_n14749_), .Y(new_n14754_));
  INVX1    g14690(.A(new_n14754_), .Y(new_n14755_));
  XOR2X1   g14691(.A(new_n14755_), .B(new_n14681_), .Y(new_n14756_));
  XOR2X1   g14692(.A(new_n14756_), .B(new_n14676_), .Y(new_n14757_));
  INVX1    g14693(.A(new_n14757_), .Y(new_n14758_));
  NOR2X1   g14694(.A(new_n14597_), .B(new_n14514_), .Y(new_n14759_));
  INVX1    g14695(.A(new_n14759_), .Y(new_n14760_));
  OR2X1    g14696(.A(new_n14602_), .B(new_n14599_), .Y(new_n14761_));
  AND2X1   g14697(.A(new_n14761_), .B(new_n14760_), .Y(new_n14762_));
  XOR2X1   g14698(.A(new_n14762_), .B(new_n14758_), .Y(new_n14763_));
  AOI22X1  g14699(.A0(new_n12076_), .A1(new_n4635_), .B0(new_n12018_), .B1(new_n4870_), .Y(new_n14764_));
  OAI21X1  g14700(.A0(new_n13679_), .A1(new_n5096_), .B0(new_n14764_), .Y(new_n14765_));
  AOI21X1  g14701(.A0(new_n13678_), .A1(new_n4637_), .B0(new_n14765_), .Y(new_n14766_));
  XOR2X1   g14702(.A(new_n14766_), .B(\a[8] ), .Y(new_n14767_));
  XOR2X1   g14703(.A(new_n14767_), .B(new_n14763_), .Y(new_n14768_));
  XOR2X1   g14704(.A(new_n14768_), .B(new_n14671_), .Y(new_n14769_));
  XOR2X1   g14705(.A(new_n14769_), .B(new_n14668_), .Y(new_n14770_));
  NOR2X1   g14706(.A(new_n14611_), .B(new_n14505_), .Y(new_n14771_));
  AOI21X1  g14707(.A0(new_n14615_), .A1(new_n14612_), .B0(new_n14771_), .Y(new_n14772_));
  XOR2X1   g14708(.A(new_n14772_), .B(new_n14770_), .Y(new_n14773_));
  AND2X1   g14709(.A(new_n14639_), .B(new_n14621_), .Y(new_n14774_));
  INVX1    g14710(.A(new_n14774_), .Y(new_n14775_));
  OAI21X1  g14711(.A0(new_n14641_), .A1(new_n14618_), .B0(new_n14775_), .Y(new_n14776_));
  NOR2X1   g14712(.A(new_n14633_), .B(new_n14629_), .Y(new_n14777_));
  NOR2X1   g14713(.A(new_n14638_), .B(new_n14634_), .Y(new_n14778_));
  NOR2X1   g14714(.A(new_n14778_), .B(new_n14777_), .Y(new_n14779_));
  INVX1    g14715(.A(new_n14627_), .Y(new_n14780_));
  INVX1    g14716(.A(new_n2647_), .Y(new_n14781_));
  NOR2X1   g14717(.A(new_n14781_), .B(new_n2394_), .Y(new_n14782_));
  NOR2X1   g14718(.A(new_n14782_), .B(new_n14780_), .Y(new_n14783_));
  INVX1    g14719(.A(new_n14783_), .Y(new_n14784_));
  INVX1    g14720(.A(new_n14624_), .Y(new_n14785_));
  AND2X1   g14721(.A(new_n14627_), .B(new_n14626_), .Y(new_n14786_));
  AOI21X1  g14722(.A0(new_n14628_), .A1(new_n14785_), .B0(new_n14786_), .Y(new_n14787_));
  XOR2X1   g14723(.A(new_n14782_), .B(new_n14780_), .Y(new_n14788_));
  NOR2X1   g14724(.A(new_n14788_), .B(new_n14787_), .Y(new_n14789_));
  INVX1    g14725(.A(new_n14787_), .Y(new_n14790_));
  NOR3X1   g14726(.A(new_n14627_), .B(new_n14781_), .C(new_n2394_), .Y(new_n14791_));
  AOI21X1  g14727(.A0(new_n14784_), .A1(new_n14790_), .B0(new_n14791_), .Y(new_n14792_));
  AOI21X1  g14728(.A0(new_n14792_), .A1(new_n14784_), .B0(new_n14789_), .Y(new_n14793_));
  OAI21X1  g14729(.A0(new_n2139_), .A1(new_n2095_), .B0(new_n7341_), .Y(new_n14794_));
  OAI21X1  g14730(.A0(new_n7644_), .A1(new_n2186_), .B0(new_n14794_), .Y(new_n14795_));
  AOI21X1  g14731(.A0(new_n7807_), .A1(new_n2062_), .B0(new_n14795_), .Y(new_n14796_));
  XOR2X1   g14732(.A(new_n14796_), .B(\a[29] ), .Y(new_n14797_));
  AOI22X1  g14733(.A0(new_n7590_), .A1(new_n1884_), .B0(new_n7578_), .B1(new_n1890_), .Y(new_n14798_));
  OAI21X1  g14734(.A0(new_n7642_), .A1(new_n3498_), .B0(new_n14798_), .Y(new_n14799_));
  AOI21X1  g14735(.A0(new_n7712_), .A1(new_n407_), .B0(new_n14799_), .Y(new_n14800_));
  XOR2X1   g14736(.A(new_n14800_), .B(new_n14797_), .Y(new_n14801_));
  XOR2X1   g14737(.A(new_n14801_), .B(new_n14793_), .Y(new_n14802_));
  XOR2X1   g14738(.A(new_n14802_), .B(new_n14779_), .Y(new_n14803_));
  XOR2X1   g14739(.A(new_n14803_), .B(new_n14776_), .Y(new_n14804_));
  INVX1    g14740(.A(new_n14804_), .Y(new_n14805_));
  AOI22X1  g14741(.A0(new_n14642_), .A1(new_n6300_), .B0(new_n14084_), .B1(new_n5970_), .Y(new_n14806_));
  OAI21X1  g14742(.A0(new_n14805_), .A1(new_n6309_), .B0(new_n14806_), .Y(new_n14807_));
  XOR2X1   g14743(.A(new_n14804_), .B(new_n14642_), .Y(new_n14808_));
  XOR2X1   g14744(.A(new_n14808_), .B(new_n14650_), .Y(new_n14809_));
  AOI21X1  g14745(.A0(new_n14809_), .A1(new_n5972_), .B0(new_n14807_), .Y(new_n14810_));
  XOR2X1   g14746(.A(new_n14810_), .B(\a[2] ), .Y(new_n14811_));
  XOR2X1   g14747(.A(new_n14811_), .B(new_n14773_), .Y(new_n14812_));
  XOR2X1   g14748(.A(new_n14812_), .B(new_n14664_), .Y(new_n14813_));
  XOR2X1   g14749(.A(new_n14813_), .B(new_n14660_), .Y(\result[1] ));
  AND2X1   g14750(.A(new_n14813_), .B(new_n14660_), .Y(new_n14815_));
  OR2X1    g14751(.A(new_n14811_), .B(new_n14773_), .Y(new_n14816_));
  OAI21X1  g14752(.A0(new_n14663_), .A1(new_n14662_), .B0(new_n14812_), .Y(new_n14817_));
  AND2X1   g14753(.A(new_n14817_), .B(new_n14816_), .Y(new_n14818_));
  AOI22X1  g14754(.A0(new_n14087_), .A1(new_n5659_), .B0(new_n14085_), .B1(new_n5373_), .Y(new_n14819_));
  OAI21X1  g14755(.A0(new_n14643_), .A1(new_n5959_), .B0(new_n14819_), .Y(new_n14820_));
  AOI21X1  g14756(.A0(new_n14106_), .A1(new_n67_), .B0(new_n14820_), .Y(new_n14821_));
  XOR2X1   g14757(.A(new_n14821_), .B(\a[5] ), .Y(new_n14822_));
  XOR2X1   g14758(.A(new_n14766_), .B(new_n2995_), .Y(new_n14823_));
  AND2X1   g14759(.A(new_n14823_), .B(new_n14763_), .Y(new_n14824_));
  INVX1    g14760(.A(new_n14768_), .Y(new_n14825_));
  AOI21X1  g14761(.A0(new_n14825_), .A1(new_n14671_), .B0(new_n14824_), .Y(new_n14826_));
  AOI22X1  g14762(.A0(new_n12081_), .A1(new_n4078_), .B0(new_n12079_), .B1(new_n4247_), .Y(new_n14827_));
  OAI21X1  g14763(.A0(new_n13700_), .A1(new_n4427_), .B0(new_n14827_), .Y(new_n14828_));
  AOI21X1  g14764(.A0(new_n13699_), .A1(new_n4080_), .B0(new_n14828_), .Y(new_n14829_));
  XOR2X1   g14765(.A(new_n14829_), .B(\a[11] ), .Y(new_n14830_));
  XOR2X1   g14766(.A(new_n14752_), .B(new_n2529_), .Y(new_n14831_));
  AND2X1   g14767(.A(new_n14831_), .B(new_n14749_), .Y(new_n14832_));
  AOI21X1  g14768(.A0(new_n14680_), .A1(new_n14679_), .B0(new_n14754_), .Y(new_n14833_));
  NOR2X1   g14769(.A(new_n14833_), .B(new_n14832_), .Y(new_n14834_));
  AOI22X1  g14770(.A0(new_n12095_), .A1(new_n3232_), .B0(new_n12093_), .B1(new_n3390_), .Y(new_n14835_));
  OAI21X1  g14771(.A0(new_n13118_), .A1(new_n3545_), .B0(new_n14835_), .Y(new_n14836_));
  AOI21X1  g14772(.A0(new_n13117_), .A1(new_n3234_), .B0(new_n14836_), .Y(new_n14837_));
  XOR2X1   g14773(.A(new_n14837_), .B(\a[17] ), .Y(new_n14838_));
  INVX1    g14774(.A(new_n14691_), .Y(new_n14839_));
  XOR2X1   g14775(.A(new_n14741_), .B(new_n1920_), .Y(new_n14840_));
  AND2X1   g14776(.A(new_n14840_), .B(new_n14738_), .Y(new_n14841_));
  INVX1    g14777(.A(new_n14841_), .Y(new_n14842_));
  OAI21X1  g14778(.A0(new_n14743_), .A1(new_n14839_), .B0(new_n14842_), .Y(new_n14843_));
  AOI22X1  g14779(.A0(new_n12208_), .A1(new_n2657_), .B0(new_n12107_), .B1(new_n2696_), .Y(new_n14844_));
  OAI21X1  g14780(.A0(new_n12695_), .A1(new_n2753_), .B0(new_n14844_), .Y(new_n14845_));
  AOI21X1  g14781(.A0(new_n12694_), .A1(new_n2658_), .B0(new_n14845_), .Y(new_n14846_));
  XOR2X1   g14782(.A(new_n14846_), .B(\a[23] ), .Y(new_n14847_));
  INVX1    g14783(.A(new_n14847_), .Y(new_n14848_));
  INVX1    g14784(.A(new_n14699_), .Y(new_n14849_));
  INVX1    g14785(.A(new_n14727_), .Y(new_n14850_));
  NOR2X1   g14786(.A(new_n14731_), .B(new_n14850_), .Y(new_n14851_));
  INVX1    g14787(.A(new_n14851_), .Y(new_n14852_));
  OAI21X1  g14788(.A0(new_n14732_), .A1(new_n14849_), .B0(new_n14852_), .Y(new_n14853_));
  NOR2X1   g14789(.A(new_n14725_), .B(new_n14721_), .Y(new_n14854_));
  AOI21X1  g14790(.A0(new_n14726_), .A1(new_n14703_), .B0(new_n14854_), .Y(new_n14855_));
  INVX1    g14791(.A(new_n14855_), .Y(new_n14856_));
  INVX1    g14792(.A(new_n14708_), .Y(new_n14857_));
  NOR2X1   g14793(.A(new_n14719_), .B(new_n14715_), .Y(new_n14858_));
  INVX1    g14794(.A(new_n14858_), .Y(new_n14859_));
  OAI21X1  g14795(.A0(new_n14720_), .A1(new_n14857_), .B0(new_n14859_), .Y(new_n14860_));
  NOR4X1   g14796(.A(new_n1588_), .B(new_n1274_), .C(new_n1156_), .D(new_n1000_), .Y(new_n14861_));
  NOR3X1   g14797(.A(new_n546_), .B(new_n679_), .C(new_n372_), .Y(new_n14862_));
  NOR3X1   g14798(.A(new_n1316_), .B(new_n678_), .C(new_n111_), .Y(new_n14863_));
  NAND3X1  g14799(.A(new_n14863_), .B(new_n14862_), .C(new_n14861_), .Y(new_n14864_));
  OR4X1    g14800(.A(new_n3797_), .B(new_n1304_), .C(new_n887_), .D(new_n104_), .Y(new_n14865_));
  OR4X1    g14801(.A(new_n7939_), .B(new_n2097_), .C(new_n772_), .D(new_n686_), .Y(new_n14866_));
  NOR4X1   g14802(.A(new_n14866_), .B(new_n14865_), .C(new_n14864_), .D(new_n1957_), .Y(new_n14867_));
  NAND3X1  g14803(.A(new_n14867_), .B(new_n1970_), .C(new_n1218_), .Y(new_n14868_));
  AOI22X1  g14804(.A0(new_n12155_), .A1(new_n1890_), .B0(new_n12151_), .B1(new_n1884_), .Y(new_n14869_));
  OAI21X1  g14805(.A0(new_n12186_), .A1(new_n3498_), .B0(new_n14869_), .Y(new_n14870_));
  AOI21X1  g14806(.A0(new_n12430_), .A1(new_n407_), .B0(new_n14870_), .Y(new_n14871_));
  XOR2X1   g14807(.A(new_n14871_), .B(new_n14868_), .Y(new_n14872_));
  XOR2X1   g14808(.A(new_n14872_), .B(new_n14860_), .Y(new_n14873_));
  AOI22X1  g14809(.A0(new_n12144_), .A1(new_n2185_), .B0(new_n12141_), .B1(new_n2095_), .Y(new_n14874_));
  OAI21X1  g14810(.A0(new_n12314_), .A1(new_n2140_), .B0(new_n14874_), .Y(new_n14875_));
  AOI21X1  g14811(.A0(new_n12313_), .A1(new_n2062_), .B0(new_n14875_), .Y(new_n14876_));
  XOR2X1   g14812(.A(new_n14876_), .B(\a[29] ), .Y(new_n14877_));
  XOR2X1   g14813(.A(new_n14877_), .B(new_n14873_), .Y(new_n14878_));
  XOR2X1   g14814(.A(new_n14878_), .B(new_n14856_), .Y(new_n14879_));
  OAI22X1  g14815(.A0(new_n12134_), .A1(new_n2666_), .B0(new_n12117_), .B1(new_n2419_), .Y(new_n14880_));
  AOI21X1  g14816(.A0(new_n12516_), .A1(new_n2423_), .B0(new_n14880_), .Y(new_n14881_));
  OAI21X1  g14817(.A0(new_n12522_), .A1(new_n2665_), .B0(new_n14881_), .Y(new_n14882_));
  XOR2X1   g14818(.A(new_n14882_), .B(new_n89_), .Y(new_n14883_));
  XOR2X1   g14819(.A(new_n14883_), .B(new_n14879_), .Y(new_n14884_));
  XOR2X1   g14820(.A(new_n14884_), .B(new_n14853_), .Y(new_n14885_));
  XOR2X1   g14821(.A(new_n14885_), .B(new_n14848_), .Y(new_n14886_));
  OR2X1    g14822(.A(new_n14733_), .B(new_n14695_), .Y(new_n14887_));
  OR2X1    g14823(.A(new_n14737_), .B(new_n14735_), .Y(new_n14888_));
  AND2X1   g14824(.A(new_n14888_), .B(new_n14887_), .Y(new_n14889_));
  XOR2X1   g14825(.A(new_n14889_), .B(new_n14886_), .Y(new_n14890_));
  OAI22X1  g14826(.A0(new_n12306_), .A1(new_n3250_), .B0(new_n12840_), .B1(new_n3144_), .Y(new_n14891_));
  AOI21X1  g14827(.A0(new_n12097_), .A1(new_n3146_), .B0(new_n14891_), .Y(new_n14892_));
  OAI21X1  g14828(.A0(new_n12856_), .A1(new_n3098_), .B0(new_n14892_), .Y(new_n14893_));
  XOR2X1   g14829(.A(new_n14893_), .B(new_n1920_), .Y(new_n14894_));
  XOR2X1   g14830(.A(new_n14894_), .B(new_n14890_), .Y(new_n14895_));
  XOR2X1   g14831(.A(new_n14895_), .B(new_n14843_), .Y(new_n14896_));
  XOR2X1   g14832(.A(new_n14896_), .B(new_n14838_), .Y(new_n14897_));
  NOR2X1   g14833(.A(new_n14744_), .B(new_n14685_), .Y(new_n14898_));
  AOI21X1  g14834(.A0(new_n14748_), .A1(new_n14745_), .B0(new_n14898_), .Y(new_n14899_));
  INVX1    g14835(.A(new_n14899_), .Y(new_n14900_));
  XOR2X1   g14836(.A(new_n14900_), .B(new_n14897_), .Y(new_n14901_));
  OAI22X1  g14837(.A0(new_n13104_), .A1(new_n3627_), .B0(new_n12298_), .B1(new_n3907_), .Y(new_n14902_));
  AOI21X1  g14838(.A0(new_n12083_), .A1(new_n3984_), .B0(new_n14902_), .Y(new_n14903_));
  OAI21X1  g14839(.A0(new_n13345_), .A1(new_n3906_), .B0(new_n14903_), .Y(new_n14904_));
  XOR2X1   g14840(.A(new_n14904_), .B(new_n2529_), .Y(new_n14905_));
  XOR2X1   g14841(.A(new_n14905_), .B(new_n14901_), .Y(new_n14906_));
  INVX1    g14842(.A(new_n14906_), .Y(new_n14907_));
  XOR2X1   g14843(.A(new_n14907_), .B(new_n14834_), .Y(new_n14908_));
  XOR2X1   g14844(.A(new_n14908_), .B(new_n14830_), .Y(new_n14909_));
  INVX1    g14845(.A(new_n14909_), .Y(new_n14910_));
  NOR2X1   g14846(.A(new_n14756_), .B(new_n14676_), .Y(new_n14911_));
  AOI21X1  g14847(.A0(new_n14761_), .A1(new_n14760_), .B0(new_n14758_), .Y(new_n14912_));
  NOR2X1   g14848(.A(new_n14912_), .B(new_n14911_), .Y(new_n14913_));
  XOR2X1   g14849(.A(new_n14913_), .B(new_n14910_), .Y(new_n14914_));
  OAI22X1  g14850(.A0(new_n13679_), .A1(new_n4869_), .B0(new_n13691_), .B1(new_n4634_), .Y(new_n14915_));
  AOI21X1  g14851(.A0(new_n12285_), .A1(new_n5097_), .B0(new_n14915_), .Y(new_n14916_));
  OAI21X1  g14852(.A0(new_n14467_), .A1(new_n4868_), .B0(new_n14916_), .Y(new_n14917_));
  XOR2X1   g14853(.A(new_n14917_), .B(new_n2995_), .Y(new_n14918_));
  XOR2X1   g14854(.A(new_n14918_), .B(new_n14914_), .Y(new_n14919_));
  INVX1    g14855(.A(new_n14919_), .Y(new_n14920_));
  XOR2X1   g14856(.A(new_n14920_), .B(new_n14826_), .Y(new_n14921_));
  XOR2X1   g14857(.A(new_n14921_), .B(new_n14822_), .Y(new_n14922_));
  INVX1    g14858(.A(new_n14770_), .Y(new_n14923_));
  OR2X1    g14859(.A(new_n14772_), .B(new_n14923_), .Y(new_n14924_));
  OAI21X1  g14860(.A0(new_n14769_), .A1(new_n14668_), .B0(new_n14924_), .Y(new_n14925_));
  XOR2X1   g14861(.A(new_n14925_), .B(new_n14922_), .Y(new_n14926_));
  NOR2X1   g14862(.A(new_n14802_), .B(new_n14779_), .Y(new_n14927_));
  AOI21X1  g14863(.A0(new_n14803_), .A1(new_n14776_), .B0(new_n14927_), .Y(new_n14928_));
  INVX1    g14864(.A(new_n14793_), .Y(new_n14929_));
  NOR2X1   g14865(.A(new_n14800_), .B(new_n14797_), .Y(new_n14930_));
  AOI21X1  g14866(.A0(new_n14801_), .A1(new_n14929_), .B0(new_n14930_), .Y(new_n14931_));
  INVX1    g14867(.A(new_n14931_), .Y(new_n14932_));
  NAND3X1  g14868(.A(new_n2186_), .B(new_n2431_), .C(new_n2061_), .Y(new_n14933_));
  AND2X1   g14869(.A(new_n14933_), .B(new_n7341_), .Y(new_n14934_));
  XOR2X1   g14870(.A(new_n14934_), .B(new_n74_), .Y(new_n14935_));
  INVX1    g14871(.A(new_n14782_), .Y(new_n14936_));
  XOR2X1   g14872(.A(new_n14936_), .B(new_n7094_), .Y(new_n14937_));
  XOR2X1   g14873(.A(new_n14937_), .B(new_n14935_), .Y(new_n14938_));
  AOI22X1  g14874(.A0(new_n7643_), .A1(new_n1889_), .B0(new_n7590_), .B1(new_n1890_), .Y(new_n14939_));
  OAI21X1  g14875(.A0(new_n7642_), .A1(new_n1885_), .B0(new_n14939_), .Y(new_n14940_));
  AOI21X1  g14876(.A0(new_n7718_), .A1(new_n407_), .B0(new_n14940_), .Y(new_n14941_));
  XOR2X1   g14877(.A(new_n14941_), .B(new_n14938_), .Y(new_n14942_));
  XOR2X1   g14878(.A(new_n14942_), .B(new_n14792_), .Y(new_n14943_));
  XOR2X1   g14879(.A(new_n14943_), .B(new_n14932_), .Y(new_n14944_));
  INVX1    g14880(.A(new_n14944_), .Y(new_n14945_));
  XOR2X1   g14881(.A(new_n14945_), .B(new_n14928_), .Y(new_n14946_));
  OAI22X1  g14882(.A0(new_n14805_), .A1(new_n6307_), .B0(new_n14648_), .B1(new_n6325_), .Y(new_n14947_));
  AOI21X1  g14883(.A0(new_n14946_), .A1(new_n6308_), .B0(new_n14947_), .Y(new_n14948_));
  NAND2X1  g14884(.A(new_n14808_), .B(new_n14650_), .Y(new_n14949_));
  OAI21X1  g14885(.A0(new_n14805_), .A1(new_n14648_), .B0(new_n14949_), .Y(new_n14950_));
  XOR2X1   g14886(.A(new_n14946_), .B(new_n14804_), .Y(new_n14951_));
  XOR2X1   g14887(.A(new_n14951_), .B(new_n14950_), .Y(new_n14952_));
  INVX1    g14888(.A(new_n14952_), .Y(new_n14953_));
  OAI21X1  g14889(.A0(new_n14953_), .A1(new_n6298_), .B0(new_n14948_), .Y(new_n14954_));
  XOR2X1   g14890(.A(new_n14954_), .B(new_n3431_), .Y(new_n14955_));
  XOR2X1   g14891(.A(new_n14955_), .B(new_n14926_), .Y(new_n14956_));
  XOR2X1   g14892(.A(new_n14956_), .B(new_n14818_), .Y(new_n14957_));
  XOR2X1   g14893(.A(new_n14957_), .B(new_n14815_), .Y(\result[2] ));
  AND2X1   g14894(.A(new_n14957_), .B(new_n14815_), .Y(new_n14959_));
  XOR2X1   g14895(.A(new_n14954_), .B(\a[2] ), .Y(new_n14960_));
  AND2X1   g14896(.A(new_n14960_), .B(new_n14926_), .Y(new_n14961_));
  AOI21X1  g14897(.A0(new_n14817_), .A1(new_n14816_), .B0(new_n14956_), .Y(new_n14962_));
  OR2X1    g14898(.A(new_n14962_), .B(new_n14961_), .Y(new_n14963_));
  AOI22X1  g14899(.A0(new_n14087_), .A1(new_n5373_), .B0(new_n14084_), .B1(new_n5659_), .Y(new_n14964_));
  OAI21X1  g14900(.A0(new_n14648_), .A1(new_n5959_), .B0(new_n14964_), .Y(new_n14965_));
  AOI21X1  g14901(.A0(new_n14651_), .A1(new_n67_), .B0(new_n14965_), .Y(new_n14966_));
  XOR2X1   g14902(.A(new_n14966_), .B(\a[5] ), .Y(new_n14967_));
  INVX1    g14903(.A(new_n14914_), .Y(new_n14968_));
  OR2X1    g14904(.A(new_n14919_), .B(new_n14826_), .Y(new_n14969_));
  OAI21X1  g14905(.A0(new_n14918_), .A1(new_n14968_), .B0(new_n14969_), .Y(new_n14970_));
  AOI22X1  g14906(.A0(new_n12079_), .A1(new_n4078_), .B0(new_n12076_), .B1(new_n4247_), .Y(new_n14971_));
  OAI21X1  g14907(.A0(new_n13691_), .A1(new_n4427_), .B0(new_n14971_), .Y(new_n14972_));
  AOI21X1  g14908(.A0(new_n13690_), .A1(new_n4080_), .B0(new_n14972_), .Y(new_n14973_));
  XOR2X1   g14909(.A(new_n14973_), .B(\a[11] ), .Y(new_n14974_));
  XOR2X1   g14910(.A(new_n14904_), .B(\a[14] ), .Y(new_n14975_));
  AND2X1   g14911(.A(new_n14975_), .B(new_n14901_), .Y(new_n14976_));
  INVX1    g14912(.A(new_n14976_), .Y(new_n14977_));
  OAI21X1  g14913(.A0(new_n14833_), .A1(new_n14832_), .B0(new_n14907_), .Y(new_n14978_));
  AND2X1   g14914(.A(new_n14978_), .B(new_n14977_), .Y(new_n14979_));
  AOI22X1  g14915(.A0(new_n12093_), .A1(new_n3232_), .B0(new_n12090_), .B1(new_n3390_), .Y(new_n14980_));
  OAI21X1  g14916(.A0(new_n13104_), .A1(new_n3545_), .B0(new_n14980_), .Y(new_n14981_));
  AOI21X1  g14917(.A0(new_n13103_), .A1(new_n3234_), .B0(new_n14981_), .Y(new_n14982_));
  XOR2X1   g14918(.A(new_n14982_), .B(\a[17] ), .Y(new_n14983_));
  INVX1    g14919(.A(new_n14843_), .Y(new_n14984_));
  INVX1    g14920(.A(new_n14894_), .Y(new_n14985_));
  AND2X1   g14921(.A(new_n14985_), .B(new_n14890_), .Y(new_n14986_));
  INVX1    g14922(.A(new_n14986_), .Y(new_n14987_));
  OAI21X1  g14923(.A0(new_n14895_), .A1(new_n14984_), .B0(new_n14987_), .Y(new_n14988_));
  AOI22X1  g14924(.A0(new_n12107_), .A1(new_n2657_), .B0(new_n12104_), .B1(new_n2696_), .Y(new_n14989_));
  OAI21X1  g14925(.A0(new_n12306_), .A1(new_n2753_), .B0(new_n14989_), .Y(new_n14990_));
  AOI21X1  g14926(.A0(new_n12305_), .A1(new_n2658_), .B0(new_n14990_), .Y(new_n14991_));
  XOR2X1   g14927(.A(new_n14991_), .B(\a[23] ), .Y(new_n14992_));
  INVX1    g14928(.A(new_n14992_), .Y(new_n14993_));
  INVX1    g14929(.A(new_n14853_), .Y(new_n14994_));
  XOR2X1   g14930(.A(new_n14882_), .B(\a[26] ), .Y(new_n14995_));
  AND2X1   g14931(.A(new_n14995_), .B(new_n14879_), .Y(new_n14996_));
  INVX1    g14932(.A(new_n14996_), .Y(new_n14997_));
  OAI21X1  g14933(.A0(new_n14884_), .A1(new_n14994_), .B0(new_n14997_), .Y(new_n14998_));
  NOR2X1   g14934(.A(new_n14877_), .B(new_n14873_), .Y(new_n14999_));
  AOI21X1  g14935(.A0(new_n14878_), .A1(new_n14856_), .B0(new_n14999_), .Y(new_n15000_));
  INVX1    g14936(.A(new_n15000_), .Y(new_n15001_));
  INVX1    g14937(.A(new_n14860_), .Y(new_n15002_));
  INVX1    g14938(.A(new_n14868_), .Y(new_n15003_));
  NOR2X1   g14939(.A(new_n14871_), .B(new_n15003_), .Y(new_n15004_));
  INVX1    g14940(.A(new_n15004_), .Y(new_n15005_));
  OAI21X1  g14941(.A0(new_n14872_), .A1(new_n15002_), .B0(new_n15005_), .Y(new_n15006_));
  NOR3X1   g14942(.A(new_n571_), .B(new_n603_), .C(new_n134_), .Y(new_n15007_));
  NOR2X1   g14943(.A(new_n2799_), .B(new_n1267_), .Y(new_n15008_));
  NAND3X1  g14944(.A(new_n15008_), .B(new_n15007_), .C(new_n1281_), .Y(new_n15009_));
  OR4X1    g14945(.A(new_n1647_), .B(new_n432_), .C(new_n412_), .D(new_n100_), .Y(new_n15010_));
  OR4X1    g14946(.A(new_n1588_), .B(new_n959_), .C(new_n474_), .D(new_n291_), .Y(new_n15011_));
  OR4X1    g14947(.A(new_n15011_), .B(new_n15010_), .C(new_n15009_), .D(new_n8568_), .Y(new_n15012_));
  NOR4X1   g14948(.A(new_n15012_), .B(new_n3817_), .C(new_n3799_), .D(new_n1495_), .Y(new_n15013_));
  INVX1    g14949(.A(new_n15013_), .Y(new_n15014_));
  AOI22X1  g14950(.A0(new_n12151_), .A1(new_n1890_), .B0(new_n12148_), .B1(new_n1884_), .Y(new_n15015_));
  OAI21X1  g14951(.A0(new_n12192_), .A1(new_n3498_), .B0(new_n15015_), .Y(new_n15016_));
  AOI21X1  g14952(.A0(new_n14540_), .A1(new_n407_), .B0(new_n15016_), .Y(new_n15017_));
  XOR2X1   g14953(.A(new_n15017_), .B(new_n15014_), .Y(new_n15018_));
  XOR2X1   g14954(.A(new_n15018_), .B(new_n15006_), .Y(new_n15019_));
  OAI22X1  g14955(.A0(new_n14194_), .A1(new_n2186_), .B0(new_n12314_), .B1(new_n2431_), .Y(new_n15020_));
  AOI21X1  g14956(.A0(new_n12133_), .A1(new_n2139_), .B0(new_n15020_), .Y(new_n15021_));
  OAI21X1  g14957(.A0(new_n14567_), .A1(new_n2063_), .B0(new_n15021_), .Y(new_n15022_));
  XOR2X1   g14958(.A(new_n15022_), .B(new_n74_), .Y(new_n15023_));
  XOR2X1   g14959(.A(new_n15023_), .B(new_n15019_), .Y(new_n15024_));
  XOR2X1   g14960(.A(new_n15024_), .B(new_n15001_), .Y(new_n15025_));
  OAI22X1  g14961(.A0(new_n12117_), .A1(new_n2666_), .B0(new_n12113_), .B1(new_n2419_), .Y(new_n15026_));
  AOI21X1  g14962(.A0(new_n12208_), .A1(new_n2423_), .B0(new_n15026_), .Y(new_n15027_));
  OAI21X1  g14963(.A0(new_n12685_), .A1(new_n2665_), .B0(new_n15027_), .Y(new_n15028_));
  XOR2X1   g14964(.A(new_n15028_), .B(new_n89_), .Y(new_n15029_));
  XOR2X1   g14965(.A(new_n15029_), .B(new_n15025_), .Y(new_n15030_));
  XOR2X1   g14966(.A(new_n15030_), .B(new_n14998_), .Y(new_n15031_));
  XOR2X1   g14967(.A(new_n15031_), .B(new_n14993_), .Y(new_n15032_));
  NOR2X1   g14968(.A(new_n14885_), .B(new_n14847_), .Y(new_n15033_));
  AOI21X1  g14969(.A0(new_n14888_), .A1(new_n14887_), .B0(new_n14886_), .Y(new_n15034_));
  NOR2X1   g14970(.A(new_n15034_), .B(new_n15033_), .Y(new_n15035_));
  XOR2X1   g14971(.A(new_n15035_), .B(new_n15032_), .Y(new_n15036_));
  OAI22X1  g14972(.A0(new_n12840_), .A1(new_n3250_), .B0(new_n12839_), .B1(new_n3144_), .Y(new_n15037_));
  AOI21X1  g14973(.A0(new_n12095_), .A1(new_n3146_), .B0(new_n15037_), .Y(new_n15038_));
  OAI21X1  g14974(.A0(new_n12846_), .A1(new_n3098_), .B0(new_n15038_), .Y(new_n15039_));
  XOR2X1   g14975(.A(new_n15039_), .B(new_n1920_), .Y(new_n15040_));
  XOR2X1   g14976(.A(new_n15040_), .B(new_n15036_), .Y(new_n15041_));
  XOR2X1   g14977(.A(new_n15041_), .B(new_n14988_), .Y(new_n15042_));
  XOR2X1   g14978(.A(new_n15042_), .B(new_n14983_), .Y(new_n15043_));
  NOR2X1   g14979(.A(new_n14896_), .B(new_n14838_), .Y(new_n15044_));
  AOI21X1  g14980(.A0(new_n14900_), .A1(new_n14897_), .B0(new_n15044_), .Y(new_n15045_));
  INVX1    g14981(.A(new_n15045_), .Y(new_n15046_));
  XOR2X1   g14982(.A(new_n15046_), .B(new_n15043_), .Y(new_n15047_));
  OAI22X1  g14983(.A0(new_n12298_), .A1(new_n3627_), .B0(new_n13321_), .B1(new_n3907_), .Y(new_n15048_));
  AOI21X1  g14984(.A0(new_n12081_), .A1(new_n3984_), .B0(new_n15048_), .Y(new_n15049_));
  OAI21X1  g14985(.A0(new_n13335_), .A1(new_n3906_), .B0(new_n15049_), .Y(new_n15050_));
  XOR2X1   g14986(.A(new_n15050_), .B(new_n2529_), .Y(new_n15051_));
  XOR2X1   g14987(.A(new_n15051_), .B(new_n15047_), .Y(new_n15052_));
  INVX1    g14988(.A(new_n15052_), .Y(new_n15053_));
  XOR2X1   g14989(.A(new_n15053_), .B(new_n14979_), .Y(new_n15054_));
  XOR2X1   g14990(.A(new_n15054_), .B(new_n14974_), .Y(new_n15055_));
  INVX1    g14991(.A(new_n15055_), .Y(new_n15056_));
  NOR2X1   g14992(.A(new_n14908_), .B(new_n14830_), .Y(new_n15057_));
  INVX1    g14993(.A(new_n15057_), .Y(new_n15058_));
  OAI21X1  g14994(.A0(new_n14912_), .A1(new_n14911_), .B0(new_n14909_), .Y(new_n15059_));
  AND2X1   g14995(.A(new_n15059_), .B(new_n15058_), .Y(new_n15060_));
  XOR2X1   g14996(.A(new_n15060_), .B(new_n15056_), .Y(new_n15061_));
  OAI22X1  g14997(.A0(new_n12292_), .A1(new_n4869_), .B0(new_n13679_), .B1(new_n4634_), .Y(new_n15062_));
  AOI21X1  g14998(.A0(new_n14085_), .A1(new_n5097_), .B0(new_n15062_), .Y(new_n15063_));
  OAI21X1  g14999(.A0(new_n14481_), .A1(new_n4868_), .B0(new_n15063_), .Y(new_n15064_));
  XOR2X1   g15000(.A(new_n15064_), .B(new_n2995_), .Y(new_n15065_));
  XOR2X1   g15001(.A(new_n15065_), .B(new_n15061_), .Y(new_n15066_));
  XOR2X1   g15002(.A(new_n15066_), .B(new_n14970_), .Y(new_n15067_));
  XOR2X1   g15003(.A(new_n15067_), .B(new_n14967_), .Y(new_n15068_));
  NOR2X1   g15004(.A(new_n14921_), .B(new_n14822_), .Y(new_n15069_));
  AOI21X1  g15005(.A0(new_n14925_), .A1(new_n14922_), .B0(new_n15069_), .Y(new_n15070_));
  XOR2X1   g15006(.A(new_n15070_), .B(new_n15068_), .Y(new_n15071_));
  AOI22X1  g15007(.A0(new_n7657_), .A1(new_n1890_), .B0(new_n7341_), .B1(new_n1889_), .Y(new_n15072_));
  OAI21X1  g15008(.A0(new_n7644_), .A1(new_n1885_), .B0(new_n15072_), .Y(new_n15073_));
  AOI21X1  g15009(.A0(new_n7656_), .A1(new_n407_), .B0(new_n15073_), .Y(new_n15074_));
  AND2X1   g15010(.A(new_n14936_), .B(new_n7094_), .Y(new_n15075_));
  AOI21X1  g15011(.A0(new_n14937_), .A1(new_n14935_), .B0(new_n15075_), .Y(new_n15076_));
  XOR2X1   g15012(.A(new_n15076_), .B(new_n2413_), .Y(new_n15077_));
  XOR2X1   g15013(.A(new_n15077_), .B(new_n15074_), .Y(new_n15078_));
  INVX1    g15014(.A(new_n14938_), .Y(new_n15079_));
  OR2X1    g15015(.A(new_n14941_), .B(new_n15079_), .Y(new_n15080_));
  OR2X1    g15016(.A(new_n14942_), .B(new_n14792_), .Y(new_n15081_));
  AND2X1   g15017(.A(new_n15081_), .B(new_n15080_), .Y(new_n15082_));
  XOR2X1   g15018(.A(new_n15082_), .B(new_n15078_), .Y(new_n15083_));
  AND2X1   g15019(.A(new_n14943_), .B(new_n14932_), .Y(new_n15084_));
  INVX1    g15020(.A(new_n15084_), .Y(new_n15085_));
  OAI21X1  g15021(.A0(new_n14945_), .A1(new_n14928_), .B0(new_n15085_), .Y(new_n15086_));
  XOR2X1   g15022(.A(new_n15086_), .B(new_n15083_), .Y(new_n15087_));
  INVX1    g15023(.A(new_n14946_), .Y(new_n15088_));
  OAI22X1  g15024(.A0(new_n15088_), .A1(new_n6307_), .B0(new_n14805_), .B1(new_n6325_), .Y(new_n15089_));
  AOI21X1  g15025(.A0(new_n15087_), .A1(new_n6308_), .B0(new_n15089_), .Y(new_n15090_));
  NAND2X1  g15026(.A(new_n14951_), .B(new_n14950_), .Y(new_n15091_));
  OAI21X1  g15027(.A0(new_n15088_), .A1(new_n14805_), .B0(new_n15091_), .Y(new_n15092_));
  NOR2X1   g15028(.A(new_n15087_), .B(new_n14946_), .Y(new_n15093_));
  INVX1    g15029(.A(new_n15093_), .Y(new_n15094_));
  XOR2X1   g15030(.A(new_n15087_), .B(new_n14946_), .Y(new_n15095_));
  INVX1    g15031(.A(new_n15095_), .Y(new_n15096_));
  AND2X1   g15032(.A(new_n15087_), .B(new_n14946_), .Y(new_n15097_));
  AOI21X1  g15033(.A0(new_n15094_), .A1(new_n15092_), .B0(new_n15097_), .Y(new_n15098_));
  AOI22X1  g15034(.A0(new_n15098_), .A1(new_n15094_), .B0(new_n15096_), .B1(new_n15092_), .Y(new_n15099_));
  OAI21X1  g15035(.A0(new_n15099_), .A1(new_n6298_), .B0(new_n15090_), .Y(new_n15100_));
  XOR2X1   g15036(.A(new_n15100_), .B(new_n3431_), .Y(new_n15101_));
  XOR2X1   g15037(.A(new_n15101_), .B(new_n15071_), .Y(new_n15102_));
  XOR2X1   g15038(.A(new_n15102_), .B(new_n14963_), .Y(new_n15103_));
  XOR2X1   g15039(.A(new_n15103_), .B(new_n14959_), .Y(\result[3] ));
  AND2X1   g15040(.A(new_n15103_), .B(new_n14959_), .Y(new_n15105_));
  OR2X1    g15041(.A(new_n15101_), .B(new_n15071_), .Y(new_n15106_));
  OAI21X1  g15042(.A0(new_n14962_), .A1(new_n14961_), .B0(new_n15102_), .Y(new_n15107_));
  AND2X1   g15043(.A(new_n15107_), .B(new_n15106_), .Y(new_n15108_));
  AOI22X1  g15044(.A0(new_n14642_), .A1(new_n5659_), .B0(new_n14084_), .B1(new_n5373_), .Y(new_n15109_));
  OAI21X1  g15045(.A0(new_n14805_), .A1(new_n5959_), .B0(new_n15109_), .Y(new_n15110_));
  AOI21X1  g15046(.A0(new_n14809_), .A1(new_n67_), .B0(new_n15110_), .Y(new_n15111_));
  XOR2X1   g15047(.A(new_n15111_), .B(\a[5] ), .Y(new_n15112_));
  XOR2X1   g15048(.A(new_n15064_), .B(\a[8] ), .Y(new_n15113_));
  AND2X1   g15049(.A(new_n15113_), .B(new_n15061_), .Y(new_n15114_));
  INVX1    g15050(.A(new_n15066_), .Y(new_n15115_));
  AOI21X1  g15051(.A0(new_n15115_), .A1(new_n14970_), .B0(new_n15114_), .Y(new_n15116_));
  AOI22X1  g15052(.A0(new_n12076_), .A1(new_n4078_), .B0(new_n12018_), .B1(new_n4247_), .Y(new_n15117_));
  OAI21X1  g15053(.A0(new_n13679_), .A1(new_n4427_), .B0(new_n15117_), .Y(new_n15118_));
  AOI21X1  g15054(.A0(new_n13678_), .A1(new_n4080_), .B0(new_n15118_), .Y(new_n15119_));
  XOR2X1   g15055(.A(new_n15119_), .B(\a[11] ), .Y(new_n15120_));
  XOR2X1   g15056(.A(new_n15050_), .B(\a[14] ), .Y(new_n15121_));
  AND2X1   g15057(.A(new_n15121_), .B(new_n15047_), .Y(new_n15122_));
  AOI21X1  g15058(.A0(new_n14978_), .A1(new_n14977_), .B0(new_n15052_), .Y(new_n15123_));
  NOR2X1   g15059(.A(new_n15123_), .B(new_n15122_), .Y(new_n15124_));
  INVX1    g15060(.A(new_n15124_), .Y(new_n15125_));
  AOI22X1  g15061(.A0(new_n12090_), .A1(new_n3232_), .B0(new_n12088_), .B1(new_n3390_), .Y(new_n15126_));
  OAI21X1  g15062(.A0(new_n12298_), .A1(new_n3545_), .B0(new_n15126_), .Y(new_n15127_));
  AOI21X1  g15063(.A0(new_n12297_), .A1(new_n3234_), .B0(new_n15127_), .Y(new_n15128_));
  XOR2X1   g15064(.A(new_n15128_), .B(\a[17] ), .Y(new_n15129_));
  INVX1    g15065(.A(new_n14988_), .Y(new_n15130_));
  INVX1    g15066(.A(new_n15040_), .Y(new_n15131_));
  AND2X1   g15067(.A(new_n15131_), .B(new_n15036_), .Y(new_n15132_));
  INVX1    g15068(.A(new_n15132_), .Y(new_n15133_));
  OAI21X1  g15069(.A0(new_n15041_), .A1(new_n15130_), .B0(new_n15133_), .Y(new_n15134_));
  AOI22X1  g15070(.A0(new_n12104_), .A1(new_n2657_), .B0(new_n12102_), .B1(new_n2696_), .Y(new_n15135_));
  OAI21X1  g15071(.A0(new_n12840_), .A1(new_n2753_), .B0(new_n15135_), .Y(new_n15136_));
  AOI21X1  g15072(.A0(new_n12859_), .A1(new_n2658_), .B0(new_n15136_), .Y(new_n15137_));
  XOR2X1   g15073(.A(new_n15137_), .B(\a[23] ), .Y(new_n15138_));
  INVX1    g15074(.A(new_n14998_), .Y(new_n15139_));
  XOR2X1   g15075(.A(new_n15028_), .B(\a[26] ), .Y(new_n15140_));
  AND2X1   g15076(.A(new_n15140_), .B(new_n15025_), .Y(new_n15141_));
  INVX1    g15077(.A(new_n15141_), .Y(new_n15142_));
  OAI21X1  g15078(.A0(new_n15030_), .A1(new_n15139_), .B0(new_n15142_), .Y(new_n15143_));
  NOR2X1   g15079(.A(new_n15023_), .B(new_n15019_), .Y(new_n15144_));
  AOI21X1  g15080(.A0(new_n15024_), .A1(new_n15001_), .B0(new_n15144_), .Y(new_n15145_));
  INVX1    g15081(.A(new_n15145_), .Y(new_n15146_));
  INVX1    g15082(.A(new_n15006_), .Y(new_n15147_));
  NOR2X1   g15083(.A(new_n15017_), .B(new_n15013_), .Y(new_n15148_));
  INVX1    g15084(.A(new_n15148_), .Y(new_n15149_));
  OAI21X1  g15085(.A0(new_n15018_), .A1(new_n15147_), .B0(new_n15149_), .Y(new_n15150_));
  OR4X1    g15086(.A(new_n1909_), .B(new_n1259_), .C(new_n873_), .D(new_n803_), .Y(new_n15151_));
  OR4X1    g15087(.A(new_n220_), .B(new_n201_), .C(new_n200_), .D(new_n521_), .Y(new_n15152_));
  OR4X1    g15088(.A(new_n15152_), .B(new_n15151_), .C(new_n572_), .D(new_n1978_), .Y(new_n15153_));
  NOR4X1   g15089(.A(new_n2089_), .B(new_n1427_), .C(new_n1224_), .D(new_n1106_), .Y(new_n15154_));
  NOR4X1   g15090(.A(new_n480_), .B(new_n1261_), .C(new_n414_), .D(new_n843_), .Y(new_n15155_));
  NOR4X1   g15091(.A(new_n372_), .B(new_n194_), .C(new_n187_), .D(new_n184_), .Y(new_n15156_));
  NAND3X1  g15092(.A(new_n15156_), .B(new_n15155_), .C(new_n15154_), .Y(new_n15157_));
  NOR2X1   g15093(.A(new_n1244_), .B(new_n814_), .Y(new_n15158_));
  NOR4X1   g15094(.A(new_n946_), .B(new_n679_), .C(new_n681_), .D(new_n111_), .Y(new_n15159_));
  NAND3X1  g15095(.A(new_n15159_), .B(new_n15158_), .C(new_n1050_), .Y(new_n15160_));
  NOR4X1   g15096(.A(new_n15160_), .B(new_n15157_), .C(new_n15153_), .D(new_n1406_), .Y(new_n15161_));
  NAND2X1  g15097(.A(new_n15161_), .B(new_n1946_), .Y(new_n15162_));
  NOR2X1   g15098(.A(new_n15162_), .B(new_n2571_), .Y(new_n15163_));
  INVX1    g15099(.A(new_n15163_), .Y(new_n15164_));
  NOR2X1   g15100(.A(new_n12444_), .B(new_n3178_), .Y(new_n15165_));
  AOI22X1  g15101(.A0(new_n12148_), .A1(new_n1890_), .B0(new_n12144_), .B1(new_n1884_), .Y(new_n15166_));
  OAI21X1  g15102(.A0(new_n14194_), .A1(new_n3498_), .B0(new_n15166_), .Y(new_n15167_));
  NOR2X1   g15103(.A(new_n15167_), .B(new_n15165_), .Y(new_n15168_));
  XOR2X1   g15104(.A(new_n15168_), .B(new_n15164_), .Y(new_n15169_));
  XOR2X1   g15105(.A(new_n15169_), .B(new_n15150_), .Y(new_n15170_));
  AOI22X1  g15106(.A0(new_n12138_), .A1(new_n2185_), .B0(new_n12133_), .B1(new_n2095_), .Y(new_n15171_));
  OAI21X1  g15107(.A0(new_n12117_), .A1(new_n2140_), .B0(new_n15171_), .Y(new_n15172_));
  AOI21X1  g15108(.A0(new_n12526_), .A1(new_n2062_), .B0(new_n15172_), .Y(new_n15173_));
  XOR2X1   g15109(.A(new_n15173_), .B(\a[29] ), .Y(new_n15174_));
  XOR2X1   g15110(.A(new_n15174_), .B(new_n15170_), .Y(new_n15175_));
  XOR2X1   g15111(.A(new_n15175_), .B(new_n15146_), .Y(new_n15176_));
  OAI22X1  g15112(.A0(new_n12113_), .A1(new_n2666_), .B0(new_n12111_), .B1(new_n2419_), .Y(new_n15177_));
  AOI21X1  g15113(.A0(new_n12107_), .A1(new_n2423_), .B0(new_n15177_), .Y(new_n15178_));
  OAI21X1  g15114(.A0(new_n12708_), .A1(new_n2665_), .B0(new_n15178_), .Y(new_n15179_));
  XOR2X1   g15115(.A(new_n15179_), .B(new_n89_), .Y(new_n15180_));
  XOR2X1   g15116(.A(new_n15180_), .B(new_n15176_), .Y(new_n15181_));
  XOR2X1   g15117(.A(new_n15181_), .B(new_n15143_), .Y(new_n15182_));
  XOR2X1   g15118(.A(new_n15182_), .B(new_n15138_), .Y(new_n15183_));
  OR2X1    g15119(.A(new_n15031_), .B(new_n14992_), .Y(new_n15184_));
  OAI21X1  g15120(.A0(new_n15035_), .A1(new_n15032_), .B0(new_n15184_), .Y(new_n15185_));
  XOR2X1   g15121(.A(new_n15185_), .B(new_n15183_), .Y(new_n15186_));
  OAI22X1  g15122(.A0(new_n12839_), .A1(new_n3250_), .B0(new_n13090_), .B1(new_n3144_), .Y(new_n15187_));
  AOI21X1  g15123(.A0(new_n12093_), .A1(new_n3146_), .B0(new_n15187_), .Y(new_n15188_));
  OAI21X1  g15124(.A0(new_n13094_), .A1(new_n3098_), .B0(new_n15188_), .Y(new_n15189_));
  XOR2X1   g15125(.A(new_n15189_), .B(new_n1920_), .Y(new_n15190_));
  XOR2X1   g15126(.A(new_n15190_), .B(new_n15186_), .Y(new_n15191_));
  XOR2X1   g15127(.A(new_n15191_), .B(new_n15134_), .Y(new_n15192_));
  XOR2X1   g15128(.A(new_n15192_), .B(new_n15129_), .Y(new_n15193_));
  NOR2X1   g15129(.A(new_n15042_), .B(new_n14983_), .Y(new_n15194_));
  AOI21X1  g15130(.A0(new_n15046_), .A1(new_n15043_), .B0(new_n15194_), .Y(new_n15195_));
  INVX1    g15131(.A(new_n15195_), .Y(new_n15196_));
  XOR2X1   g15132(.A(new_n15196_), .B(new_n15193_), .Y(new_n15197_));
  OAI22X1  g15133(.A0(new_n13321_), .A1(new_n3627_), .B0(new_n13320_), .B1(new_n3907_), .Y(new_n15198_));
  AOI21X1  g15134(.A0(new_n12079_), .A1(new_n3984_), .B0(new_n15198_), .Y(new_n15199_));
  OAI21X1  g15135(.A0(new_n13325_), .A1(new_n3906_), .B0(new_n15199_), .Y(new_n15200_));
  XOR2X1   g15136(.A(new_n15200_), .B(new_n2529_), .Y(new_n15201_));
  XOR2X1   g15137(.A(new_n15201_), .B(new_n15197_), .Y(new_n15202_));
  XOR2X1   g15138(.A(new_n15202_), .B(new_n15125_), .Y(new_n15203_));
  XOR2X1   g15139(.A(new_n15203_), .B(new_n15120_), .Y(new_n15204_));
  INVX1    g15140(.A(new_n15204_), .Y(new_n15205_));
  NOR2X1   g15141(.A(new_n15054_), .B(new_n14974_), .Y(new_n15206_));
  AOI21X1  g15142(.A0(new_n15059_), .A1(new_n15058_), .B0(new_n15056_), .Y(new_n15207_));
  NOR2X1   g15143(.A(new_n15207_), .B(new_n15206_), .Y(new_n15208_));
  XOR2X1   g15144(.A(new_n15208_), .B(new_n15205_), .Y(new_n15209_));
  OAI22X1  g15145(.A0(new_n14086_), .A1(new_n4869_), .B0(new_n12292_), .B1(new_n4634_), .Y(new_n15210_));
  AOI21X1  g15146(.A0(new_n14087_), .A1(new_n5097_), .B0(new_n15210_), .Y(new_n15211_));
  OAI21X1  g15147(.A0(new_n14492_), .A1(new_n4868_), .B0(new_n15211_), .Y(new_n15212_));
  XOR2X1   g15148(.A(new_n15212_), .B(new_n2995_), .Y(new_n15213_));
  XOR2X1   g15149(.A(new_n15213_), .B(new_n15209_), .Y(new_n15214_));
  INVX1    g15150(.A(new_n15214_), .Y(new_n15215_));
  XOR2X1   g15151(.A(new_n15215_), .B(new_n15116_), .Y(new_n15216_));
  XOR2X1   g15152(.A(new_n15216_), .B(new_n15112_), .Y(new_n15217_));
  NOR2X1   g15153(.A(new_n15067_), .B(new_n14967_), .Y(new_n15218_));
  INVX1    g15154(.A(new_n15218_), .Y(new_n15219_));
  INVX1    g15155(.A(new_n15068_), .Y(new_n15220_));
  OAI21X1  g15156(.A0(new_n15070_), .A1(new_n15220_), .B0(new_n15219_), .Y(new_n15221_));
  XOR2X1   g15157(.A(new_n15221_), .B(new_n15217_), .Y(new_n15222_));
  OAI21X1  g15158(.A0(new_n1889_), .A1(new_n1884_), .B0(new_n7341_), .Y(new_n15223_));
  OAI21X1  g15159(.A0(new_n7644_), .A1(new_n2245_), .B0(new_n15223_), .Y(new_n15224_));
  AOI21X1  g15160(.A0(new_n7807_), .A1(new_n407_), .B0(new_n15224_), .Y(new_n15225_));
  XOR2X1   g15161(.A(new_n15225_), .B(new_n2412_), .Y(new_n15226_));
  INVX1    g15162(.A(new_n15074_), .Y(new_n15227_));
  NOR2X1   g15163(.A(new_n15076_), .B(new_n2413_), .Y(new_n15228_));
  AOI21X1  g15164(.A0(new_n15077_), .A1(new_n15227_), .B0(new_n15228_), .Y(new_n15229_));
  XOR2X1   g15165(.A(new_n15229_), .B(new_n15226_), .Y(new_n15230_));
  INVX1    g15166(.A(new_n15230_), .Y(new_n15231_));
  NOR2X1   g15167(.A(new_n15082_), .B(new_n15078_), .Y(new_n15232_));
  AOI21X1  g15168(.A0(new_n15086_), .A1(new_n15083_), .B0(new_n15232_), .Y(new_n15233_));
  XOR2X1   g15169(.A(new_n15233_), .B(new_n15231_), .Y(new_n15234_));
  INVX1    g15170(.A(new_n15087_), .Y(new_n15235_));
  OAI22X1  g15171(.A0(new_n15235_), .A1(new_n6307_), .B0(new_n15088_), .B1(new_n6325_), .Y(new_n15236_));
  AOI21X1  g15172(.A0(new_n15234_), .A1(new_n6308_), .B0(new_n15236_), .Y(new_n15237_));
  INVX1    g15173(.A(new_n15098_), .Y(new_n15238_));
  XOR2X1   g15174(.A(new_n15234_), .B(new_n15087_), .Y(new_n15239_));
  XOR2X1   g15175(.A(new_n15239_), .B(new_n15238_), .Y(new_n15240_));
  INVX1    g15176(.A(new_n15240_), .Y(new_n15241_));
  OAI21X1  g15177(.A0(new_n15241_), .A1(new_n6298_), .B0(new_n15237_), .Y(new_n15242_));
  XOR2X1   g15178(.A(new_n15242_), .B(new_n3431_), .Y(new_n15243_));
  XOR2X1   g15179(.A(new_n15243_), .B(new_n15222_), .Y(new_n15244_));
  XOR2X1   g15180(.A(new_n15244_), .B(new_n15108_), .Y(new_n15245_));
  XOR2X1   g15181(.A(new_n15245_), .B(new_n15105_), .Y(\result[4] ));
  AND2X1   g15182(.A(new_n15245_), .B(new_n15105_), .Y(new_n15247_));
  XOR2X1   g15183(.A(new_n15242_), .B(\a[2] ), .Y(new_n15248_));
  AND2X1   g15184(.A(new_n15248_), .B(new_n15222_), .Y(new_n15249_));
  AOI21X1  g15185(.A0(new_n15107_), .A1(new_n15106_), .B0(new_n15244_), .Y(new_n15250_));
  OR2X1    g15186(.A(new_n15250_), .B(new_n15249_), .Y(new_n15251_));
  AOI22X1  g15187(.A0(new_n14804_), .A1(new_n5659_), .B0(new_n14642_), .B1(new_n5373_), .Y(new_n15252_));
  OAI21X1  g15188(.A0(new_n15088_), .A1(new_n5959_), .B0(new_n15252_), .Y(new_n15253_));
  AOI21X1  g15189(.A0(new_n14952_), .A1(new_n67_), .B0(new_n15253_), .Y(new_n15254_));
  XOR2X1   g15190(.A(new_n15254_), .B(\a[5] ), .Y(new_n15255_));
  XOR2X1   g15191(.A(new_n15212_), .B(\a[8] ), .Y(new_n15256_));
  AND2X1   g15192(.A(new_n15256_), .B(new_n15209_), .Y(new_n15257_));
  INVX1    g15193(.A(new_n15257_), .Y(new_n15258_));
  OAI21X1  g15194(.A0(new_n15214_), .A1(new_n15116_), .B0(new_n15258_), .Y(new_n15259_));
  AOI22X1  g15195(.A0(new_n12074_), .A1(new_n4247_), .B0(new_n12018_), .B1(new_n4078_), .Y(new_n15260_));
  OAI21X1  g15196(.A0(new_n12292_), .A1(new_n4427_), .B0(new_n15260_), .Y(new_n15261_));
  AOI21X1  g15197(.A0(new_n12291_), .A1(new_n4080_), .B0(new_n15261_), .Y(new_n15262_));
  XOR2X1   g15198(.A(new_n15262_), .B(\a[11] ), .Y(new_n15263_));
  XOR2X1   g15199(.A(new_n15200_), .B(\a[14] ), .Y(new_n15264_));
  NOR2X1   g15200(.A(new_n15202_), .B(new_n15124_), .Y(new_n15265_));
  AOI21X1  g15201(.A0(new_n15264_), .A1(new_n15197_), .B0(new_n15265_), .Y(new_n15266_));
  AOI22X1  g15202(.A0(new_n12088_), .A1(new_n3232_), .B0(new_n12085_), .B1(new_n3390_), .Y(new_n15267_));
  OAI21X1  g15203(.A0(new_n13321_), .A1(new_n3545_), .B0(new_n15267_), .Y(new_n15268_));
  AOI21X1  g15204(.A0(new_n13344_), .A1(new_n3234_), .B0(new_n15268_), .Y(new_n15269_));
  XOR2X1   g15205(.A(new_n15269_), .B(\a[17] ), .Y(new_n15270_));
  INVX1    g15206(.A(new_n15134_), .Y(new_n15271_));
  XOR2X1   g15207(.A(new_n15189_), .B(\a[20] ), .Y(new_n15272_));
  AND2X1   g15208(.A(new_n15272_), .B(new_n15186_), .Y(new_n15273_));
  INVX1    g15209(.A(new_n15273_), .Y(new_n15274_));
  OAI21X1  g15210(.A0(new_n15191_), .A1(new_n15271_), .B0(new_n15274_), .Y(new_n15275_));
  AOI22X1  g15211(.A0(new_n12102_), .A1(new_n2657_), .B0(new_n12099_), .B1(new_n2696_), .Y(new_n15276_));
  OAI21X1  g15212(.A0(new_n12839_), .A1(new_n2753_), .B0(new_n15276_), .Y(new_n15277_));
  AOI21X1  g15213(.A0(new_n12855_), .A1(new_n2658_), .B0(new_n15277_), .Y(new_n15278_));
  XOR2X1   g15214(.A(new_n15278_), .B(\a[23] ), .Y(new_n15279_));
  INVX1    g15215(.A(new_n15143_), .Y(new_n15280_));
  XOR2X1   g15216(.A(new_n15179_), .B(\a[26] ), .Y(new_n15281_));
  AND2X1   g15217(.A(new_n15281_), .B(new_n15176_), .Y(new_n15282_));
  INVX1    g15218(.A(new_n15282_), .Y(new_n15283_));
  OAI21X1  g15219(.A0(new_n15181_), .A1(new_n15280_), .B0(new_n15283_), .Y(new_n15284_));
  INVX1    g15220(.A(new_n15284_), .Y(new_n15285_));
  NOR2X1   g15221(.A(new_n15174_), .B(new_n15170_), .Y(new_n15286_));
  AOI21X1  g15222(.A0(new_n15175_), .A1(new_n15146_), .B0(new_n15286_), .Y(new_n15287_));
  INVX1    g15223(.A(new_n15287_), .Y(new_n15288_));
  INVX1    g15224(.A(new_n15150_), .Y(new_n15289_));
  NOR2X1   g15225(.A(new_n15168_), .B(new_n15163_), .Y(new_n15290_));
  INVX1    g15226(.A(new_n15290_), .Y(new_n15291_));
  OAI21X1  g15227(.A0(new_n15169_), .A1(new_n15289_), .B0(new_n15291_), .Y(new_n15292_));
  OR4X1    g15228(.A(new_n2074_), .B(new_n896_), .C(new_n667_), .D(new_n434_), .Y(new_n15293_));
  OAI22X1  g15229(.A0(new_n143_), .A1(new_n91_), .B0(new_n92_), .B1(new_n79_), .Y(new_n15294_));
  OR4X1    g15230(.A(new_n300_), .B(new_n260_), .C(new_n812_), .D(new_n183_), .Y(new_n15295_));
  OR4X1    g15231(.A(new_n536_), .B(new_n197_), .C(new_n184_), .D(new_n410_), .Y(new_n15296_));
  OR4X1    g15232(.A(new_n15296_), .B(new_n15295_), .C(new_n15294_), .D(new_n1082_), .Y(new_n15297_));
  NOR4X1   g15233(.A(new_n15297_), .B(new_n15293_), .C(new_n6786_), .D(new_n2220_), .Y(new_n15298_));
  NAND3X1  g15234(.A(new_n15298_), .B(new_n8696_), .C(new_n3032_), .Y(new_n15299_));
  AOI22X1  g15235(.A0(new_n12144_), .A1(new_n1890_), .B0(new_n12141_), .B1(new_n1884_), .Y(new_n15300_));
  OAI21X1  g15236(.A0(new_n12314_), .A1(new_n3498_), .B0(new_n15300_), .Y(new_n15301_));
  AOI21X1  g15237(.A0(new_n12313_), .A1(new_n407_), .B0(new_n15301_), .Y(new_n15302_));
  XOR2X1   g15238(.A(new_n15302_), .B(new_n15299_), .Y(new_n15303_));
  XOR2X1   g15239(.A(new_n15303_), .B(new_n15292_), .Y(new_n15304_));
  OAI22X1  g15240(.A0(new_n12134_), .A1(new_n2186_), .B0(new_n12117_), .B1(new_n2431_), .Y(new_n15305_));
  AOI21X1  g15241(.A0(new_n12516_), .A1(new_n2139_), .B0(new_n15305_), .Y(new_n15306_));
  OAI21X1  g15242(.A0(new_n12522_), .A1(new_n2063_), .B0(new_n15306_), .Y(new_n15307_));
  XOR2X1   g15243(.A(new_n15307_), .B(new_n74_), .Y(new_n15308_));
  XOR2X1   g15244(.A(new_n15308_), .B(new_n15304_), .Y(new_n15309_));
  XOR2X1   g15245(.A(new_n15309_), .B(new_n15288_), .Y(new_n15310_));
  OAI22X1  g15246(.A0(new_n12111_), .A1(new_n2666_), .B0(new_n12109_), .B1(new_n2419_), .Y(new_n15311_));
  AOI21X1  g15247(.A0(new_n12104_), .A1(new_n2423_), .B0(new_n15311_), .Y(new_n15312_));
  OAI21X1  g15248(.A0(new_n12693_), .A1(new_n2665_), .B0(new_n15312_), .Y(new_n15313_));
  XOR2X1   g15249(.A(new_n15313_), .B(\a[26] ), .Y(new_n15314_));
  XOR2X1   g15250(.A(new_n15314_), .B(new_n15310_), .Y(new_n15315_));
  XOR2X1   g15251(.A(new_n15315_), .B(new_n15285_), .Y(new_n15316_));
  XOR2X1   g15252(.A(new_n15316_), .B(new_n15279_), .Y(new_n15317_));
  INVX1    g15253(.A(new_n15317_), .Y(new_n15318_));
  NOR2X1   g15254(.A(new_n15182_), .B(new_n15138_), .Y(new_n15319_));
  AOI21X1  g15255(.A0(new_n15185_), .A1(new_n15183_), .B0(new_n15319_), .Y(new_n15320_));
  XOR2X1   g15256(.A(new_n15320_), .B(new_n15318_), .Y(new_n15321_));
  OAI22X1  g15257(.A0(new_n13090_), .A1(new_n3250_), .B0(new_n13366_), .B1(new_n3144_), .Y(new_n15322_));
  AOI21X1  g15258(.A0(new_n12090_), .A1(new_n3146_), .B0(new_n15322_), .Y(new_n15323_));
  OAI21X1  g15259(.A0(new_n13116_), .A1(new_n3098_), .B0(new_n15323_), .Y(new_n15324_));
  XOR2X1   g15260(.A(new_n15324_), .B(new_n1920_), .Y(new_n15325_));
  XOR2X1   g15261(.A(new_n15325_), .B(new_n15321_), .Y(new_n15326_));
  XOR2X1   g15262(.A(new_n15326_), .B(new_n15275_), .Y(new_n15327_));
  XOR2X1   g15263(.A(new_n15327_), .B(new_n15270_), .Y(new_n15328_));
  NOR2X1   g15264(.A(new_n15192_), .B(new_n15129_), .Y(new_n15329_));
  AOI21X1  g15265(.A0(new_n15196_), .A1(new_n15193_), .B0(new_n15329_), .Y(new_n15330_));
  INVX1    g15266(.A(new_n15330_), .Y(new_n15331_));
  XOR2X1   g15267(.A(new_n15331_), .B(new_n15328_), .Y(new_n15332_));
  OAI22X1  g15268(.A0(new_n13320_), .A1(new_n3627_), .B0(new_n13665_), .B1(new_n3907_), .Y(new_n15333_));
  AOI21X1  g15269(.A0(new_n12076_), .A1(new_n3984_), .B0(new_n15333_), .Y(new_n15334_));
  OAI21X1  g15270(.A0(new_n13672_), .A1(new_n3906_), .B0(new_n15334_), .Y(new_n15335_));
  XOR2X1   g15271(.A(new_n15335_), .B(new_n2529_), .Y(new_n15336_));
  XOR2X1   g15272(.A(new_n15336_), .B(new_n15332_), .Y(new_n15337_));
  INVX1    g15273(.A(new_n15337_), .Y(new_n15338_));
  XOR2X1   g15274(.A(new_n15338_), .B(new_n15266_), .Y(new_n15339_));
  XOR2X1   g15275(.A(new_n15339_), .B(new_n15263_), .Y(new_n15340_));
  INVX1    g15276(.A(new_n15340_), .Y(new_n15341_));
  NOR2X1   g15277(.A(new_n15203_), .B(new_n15120_), .Y(new_n15342_));
  NOR2X1   g15278(.A(new_n15208_), .B(new_n15205_), .Y(new_n15343_));
  NOR2X1   g15279(.A(new_n15343_), .B(new_n15342_), .Y(new_n15344_));
  XOR2X1   g15280(.A(new_n15344_), .B(new_n15341_), .Y(new_n15345_));
  OAI22X1  g15281(.A0(new_n14088_), .A1(new_n4869_), .B0(new_n14086_), .B1(new_n4634_), .Y(new_n15346_));
  AOI21X1  g15282(.A0(new_n14084_), .A1(new_n5097_), .B0(new_n15346_), .Y(new_n15347_));
  OAI21X1  g15283(.A0(new_n14107_), .A1(new_n4868_), .B0(new_n15347_), .Y(new_n15348_));
  XOR2X1   g15284(.A(new_n15348_), .B(new_n2995_), .Y(new_n15349_));
  XOR2X1   g15285(.A(new_n15349_), .B(new_n15345_), .Y(new_n15350_));
  XOR2X1   g15286(.A(new_n15350_), .B(new_n15259_), .Y(new_n15351_));
  XOR2X1   g15287(.A(new_n15351_), .B(new_n15255_), .Y(new_n15352_));
  NOR2X1   g15288(.A(new_n15216_), .B(new_n15112_), .Y(new_n15353_));
  AOI21X1  g15289(.A0(new_n15221_), .A1(new_n15217_), .B0(new_n15353_), .Y(new_n15354_));
  XOR2X1   g15290(.A(new_n15354_), .B(new_n15352_), .Y(new_n15355_));
  NOR2X1   g15291(.A(new_n15229_), .B(new_n15226_), .Y(new_n15356_));
  INVX1    g15292(.A(new_n15356_), .Y(new_n15357_));
  OAI21X1  g15293(.A0(new_n15233_), .A1(new_n15231_), .B0(new_n15357_), .Y(new_n15358_));
  AND2X1   g15294(.A(new_n15225_), .B(new_n2412_), .Y(new_n15359_));
  AOI21X1  g15295(.A0(new_n83_), .A1(new_n1888_), .B0(new_n8172_), .Y(new_n15360_));
  XOR2X1   g15296(.A(new_n15360_), .B(new_n15359_), .Y(new_n15361_));
  XOR2X1   g15297(.A(new_n15361_), .B(new_n15358_), .Y(new_n15362_));
  INVX1    g15298(.A(new_n15234_), .Y(new_n15363_));
  OAI22X1  g15299(.A0(new_n15363_), .A1(new_n6307_), .B0(new_n15235_), .B1(new_n6325_), .Y(new_n15364_));
  AOI21X1  g15300(.A0(new_n15362_), .A1(new_n6308_), .B0(new_n15364_), .Y(new_n15365_));
  NAND2X1  g15301(.A(new_n15239_), .B(new_n15238_), .Y(new_n15366_));
  OAI21X1  g15302(.A0(new_n15363_), .A1(new_n15235_), .B0(new_n15366_), .Y(new_n15367_));
  NOR2X1   g15303(.A(new_n15362_), .B(new_n15234_), .Y(new_n15368_));
  INVX1    g15304(.A(new_n15368_), .Y(new_n15369_));
  XOR2X1   g15305(.A(new_n15362_), .B(new_n15234_), .Y(new_n15370_));
  INVX1    g15306(.A(new_n15370_), .Y(new_n15371_));
  AND2X1   g15307(.A(new_n15362_), .B(new_n15234_), .Y(new_n15372_));
  AOI21X1  g15308(.A0(new_n15369_), .A1(new_n15367_), .B0(new_n15372_), .Y(new_n15373_));
  AOI22X1  g15309(.A0(new_n15373_), .A1(new_n15369_), .B0(new_n15371_), .B1(new_n15367_), .Y(new_n15374_));
  OAI21X1  g15310(.A0(new_n15374_), .A1(new_n6298_), .B0(new_n15365_), .Y(new_n15375_));
  XOR2X1   g15311(.A(new_n15375_), .B(new_n3431_), .Y(new_n15376_));
  XOR2X1   g15312(.A(new_n15376_), .B(new_n15355_), .Y(new_n15377_));
  XOR2X1   g15313(.A(new_n15377_), .B(new_n15251_), .Y(new_n15378_));
  XOR2X1   g15314(.A(new_n15378_), .B(new_n15247_), .Y(\result[5] ));
  AND2X1   g15315(.A(new_n15378_), .B(new_n15247_), .Y(new_n15380_));
  INVX1    g15316(.A(new_n15099_), .Y(new_n15381_));
  AOI22X1  g15317(.A0(new_n14946_), .A1(new_n5659_), .B0(new_n14804_), .B1(new_n5373_), .Y(new_n15382_));
  OAI21X1  g15318(.A0(new_n15235_), .A1(new_n5959_), .B0(new_n15382_), .Y(new_n15383_));
  AOI21X1  g15319(.A0(new_n15381_), .A1(new_n67_), .B0(new_n15383_), .Y(new_n15384_));
  XOR2X1   g15320(.A(new_n15384_), .B(\a[5] ), .Y(new_n15385_));
  INVX1    g15321(.A(new_n15259_), .Y(new_n15386_));
  INVX1    g15322(.A(new_n15349_), .Y(new_n15387_));
  NAND2X1  g15323(.A(new_n15387_), .B(new_n15345_), .Y(new_n15388_));
  OAI21X1  g15324(.A0(new_n15350_), .A1(new_n15386_), .B0(new_n15388_), .Y(new_n15389_));
  AOI22X1  g15325(.A0(new_n12285_), .A1(new_n4247_), .B0(new_n12074_), .B1(new_n4078_), .Y(new_n15390_));
  OAI21X1  g15326(.A0(new_n14086_), .A1(new_n4427_), .B0(new_n15390_), .Y(new_n15391_));
  AOI21X1  g15327(.A0(new_n14480_), .A1(new_n4080_), .B0(new_n15391_), .Y(new_n15392_));
  XOR2X1   g15328(.A(new_n15392_), .B(\a[11] ), .Y(new_n15393_));
  INVX1    g15329(.A(new_n15393_), .Y(new_n15394_));
  INVX1    g15330(.A(new_n15336_), .Y(new_n15395_));
  NAND2X1  g15331(.A(new_n15395_), .B(new_n15332_), .Y(new_n15396_));
  OAI21X1  g15332(.A0(new_n15337_), .A1(new_n15266_), .B0(new_n15396_), .Y(new_n15397_));
  AOI22X1  g15333(.A0(new_n12085_), .A1(new_n3232_), .B0(new_n12083_), .B1(new_n3390_), .Y(new_n15398_));
  OAI21X1  g15334(.A0(new_n13320_), .A1(new_n3545_), .B0(new_n15398_), .Y(new_n15399_));
  AOI21X1  g15335(.A0(new_n14510_), .A1(new_n3234_), .B0(new_n15399_), .Y(new_n15400_));
  XOR2X1   g15336(.A(new_n15400_), .B(\a[17] ), .Y(new_n15401_));
  INVX1    g15337(.A(new_n15401_), .Y(new_n15402_));
  INVX1    g15338(.A(new_n15275_), .Y(new_n15403_));
  INVX1    g15339(.A(new_n15325_), .Y(new_n15404_));
  NAND2X1  g15340(.A(new_n15404_), .B(new_n15321_), .Y(new_n15405_));
  OAI21X1  g15341(.A0(new_n15326_), .A1(new_n15403_), .B0(new_n15405_), .Y(new_n15406_));
  AOI22X1  g15342(.A0(new_n12099_), .A1(new_n2657_), .B0(new_n12097_), .B1(new_n2696_), .Y(new_n15407_));
  OAI21X1  g15343(.A0(new_n13090_), .A1(new_n2753_), .B0(new_n15407_), .Y(new_n15408_));
  AOI21X1  g15344(.A0(new_n14519_), .A1(new_n2658_), .B0(new_n15408_), .Y(new_n15409_));
  XOR2X1   g15345(.A(new_n15409_), .B(\a[23] ), .Y(new_n15410_));
  AND2X1   g15346(.A(new_n15314_), .B(new_n15310_), .Y(new_n15411_));
  AND2X1   g15347(.A(new_n15315_), .B(new_n15284_), .Y(new_n15412_));
  OR2X1    g15348(.A(new_n15412_), .B(new_n15411_), .Y(new_n15413_));
  NOR2X1   g15349(.A(new_n15308_), .B(new_n15304_), .Y(new_n15414_));
  AOI21X1  g15350(.A0(new_n15309_), .A1(new_n15288_), .B0(new_n15414_), .Y(new_n15415_));
  INVX1    g15351(.A(new_n15292_), .Y(new_n15416_));
  INVX1    g15352(.A(new_n15299_), .Y(new_n15417_));
  NOR2X1   g15353(.A(new_n15302_), .B(new_n15417_), .Y(new_n15418_));
  INVX1    g15354(.A(new_n15418_), .Y(new_n15419_));
  OAI21X1  g15355(.A0(new_n15303_), .A1(new_n15416_), .B0(new_n15419_), .Y(new_n15420_));
  OR4X1    g15356(.A(new_n7941_), .B(new_n1909_), .C(new_n873_), .D(new_n569_), .Y(new_n15421_));
  OR4X1    g15357(.A(new_n459_), .B(new_n702_), .C(new_n603_), .D(new_n203_), .Y(new_n15422_));
  OR4X1    g15358(.A(new_n1249_), .B(new_n1516_), .C(new_n479_), .D(new_n144_), .Y(new_n15423_));
  OR2X1    g15359(.A(new_n15423_), .B(new_n15422_), .Y(new_n15424_));
  NOR4X1   g15360(.A(new_n530_), .B(new_n1390_), .C(new_n878_), .D(new_n465_), .Y(new_n15425_));
  NOR4X1   g15361(.A(new_n636_), .B(new_n301_), .C(new_n400_), .D(new_n757_), .Y(new_n15426_));
  NOR3X1   g15362(.A(new_n1022_), .B(new_n194_), .C(new_n80_), .Y(new_n15427_));
  NAND3X1  g15363(.A(new_n15427_), .B(new_n15426_), .C(new_n15425_), .Y(new_n15428_));
  OR4X1    g15364(.A(new_n15428_), .B(new_n15424_), .C(new_n15421_), .D(new_n15010_), .Y(new_n15429_));
  NOR4X1   g15365(.A(new_n15429_), .B(new_n8178_), .C(new_n2925_), .D(new_n1611_), .Y(new_n15430_));
  INVX1    g15366(.A(new_n15430_), .Y(new_n15431_));
  AOI22X1  g15367(.A0(new_n12141_), .A1(new_n1890_), .B0(new_n12138_), .B1(new_n1884_), .Y(new_n15432_));
  OAI21X1  g15368(.A0(new_n12134_), .A1(new_n3498_), .B0(new_n15432_), .Y(new_n15433_));
  AOI21X1  g15369(.A0(new_n12536_), .A1(new_n407_), .B0(new_n15433_), .Y(new_n15434_));
  XOR2X1   g15370(.A(new_n15434_), .B(new_n15431_), .Y(new_n15435_));
  XOR2X1   g15371(.A(new_n15435_), .B(new_n15420_), .Y(new_n15436_));
  OAI22X1  g15372(.A0(new_n12117_), .A1(new_n2186_), .B0(new_n12113_), .B1(new_n2431_), .Y(new_n15437_));
  AOI21X1  g15373(.A0(new_n12208_), .A1(new_n2139_), .B0(new_n15437_), .Y(new_n15438_));
  OAI21X1  g15374(.A0(new_n12685_), .A1(new_n2063_), .B0(new_n15438_), .Y(new_n15439_));
  XOR2X1   g15375(.A(new_n15439_), .B(new_n74_), .Y(new_n15440_));
  XOR2X1   g15376(.A(new_n15440_), .B(new_n15436_), .Y(new_n15441_));
  XOR2X1   g15377(.A(new_n15441_), .B(new_n15415_), .Y(new_n15442_));
  OAI22X1  g15378(.A0(new_n12109_), .A1(new_n2666_), .B0(new_n12695_), .B1(new_n2419_), .Y(new_n15443_));
  AOI21X1  g15379(.A0(new_n12102_), .A1(new_n2423_), .B0(new_n15443_), .Y(new_n15444_));
  OAI21X1  g15380(.A0(new_n14578_), .A1(new_n2665_), .B0(new_n15444_), .Y(new_n15445_));
  XOR2X1   g15381(.A(new_n15445_), .B(new_n89_), .Y(new_n15446_));
  XOR2X1   g15382(.A(new_n15446_), .B(new_n15442_), .Y(new_n15447_));
  XOR2X1   g15383(.A(new_n15447_), .B(new_n15413_), .Y(new_n15448_));
  XOR2X1   g15384(.A(new_n15448_), .B(new_n15410_), .Y(new_n15449_));
  INVX1    g15385(.A(new_n15449_), .Y(new_n15450_));
  OR2X1    g15386(.A(new_n15316_), .B(new_n15279_), .Y(new_n15451_));
  OAI21X1  g15387(.A0(new_n15320_), .A1(new_n15318_), .B0(new_n15451_), .Y(new_n15452_));
  XOR2X1   g15388(.A(new_n15452_), .B(new_n15450_), .Y(new_n15453_));
  INVX1    g15389(.A(new_n15453_), .Y(new_n15454_));
  OAI22X1  g15390(.A0(new_n13366_), .A1(new_n3250_), .B0(new_n13118_), .B1(new_n3144_), .Y(new_n15455_));
  AOI21X1  g15391(.A0(new_n12088_), .A1(new_n3146_), .B0(new_n15455_), .Y(new_n15456_));
  OAI21X1  g15392(.A0(new_n14590_), .A1(new_n3098_), .B0(new_n15456_), .Y(new_n15457_));
  XOR2X1   g15393(.A(new_n15457_), .B(new_n1920_), .Y(new_n15458_));
  XOR2X1   g15394(.A(new_n15458_), .B(new_n15454_), .Y(new_n15459_));
  XOR2X1   g15395(.A(new_n15459_), .B(new_n15406_), .Y(new_n15460_));
  XOR2X1   g15396(.A(new_n15460_), .B(new_n15402_), .Y(new_n15461_));
  NOR2X1   g15397(.A(new_n15327_), .B(new_n15270_), .Y(new_n15462_));
  AOI21X1  g15398(.A0(new_n15331_), .A1(new_n15328_), .B0(new_n15462_), .Y(new_n15463_));
  INVX1    g15399(.A(new_n15463_), .Y(new_n15464_));
  XOR2X1   g15400(.A(new_n15464_), .B(new_n15461_), .Y(new_n15465_));
  OAI22X1  g15401(.A0(new_n13665_), .A1(new_n3627_), .B0(new_n13700_), .B1(new_n3907_), .Y(new_n15466_));
  AOI21X1  g15402(.A0(new_n12018_), .A1(new_n3984_), .B0(new_n15466_), .Y(new_n15467_));
  OAI21X1  g15403(.A0(new_n14604_), .A1(new_n3906_), .B0(new_n15467_), .Y(new_n15468_));
  XOR2X1   g15404(.A(new_n15468_), .B(new_n2529_), .Y(new_n15469_));
  INVX1    g15405(.A(new_n15469_), .Y(new_n15470_));
  XOR2X1   g15406(.A(new_n15470_), .B(new_n15465_), .Y(new_n15471_));
  XOR2X1   g15407(.A(new_n15471_), .B(new_n15397_), .Y(new_n15472_));
  XOR2X1   g15408(.A(new_n15472_), .B(new_n15394_), .Y(new_n15473_));
  OR2X1    g15409(.A(new_n15339_), .B(new_n15263_), .Y(new_n15474_));
  OAI21X1  g15410(.A0(new_n15343_), .A1(new_n15342_), .B0(new_n15340_), .Y(new_n15475_));
  AND2X1   g15411(.A(new_n15475_), .B(new_n15474_), .Y(new_n15476_));
  INVX1    g15412(.A(new_n15476_), .Y(new_n15477_));
  XOR2X1   g15413(.A(new_n15477_), .B(new_n15473_), .Y(new_n15478_));
  OAI22X1  g15414(.A0(new_n14088_), .A1(new_n4634_), .B0(new_n14643_), .B1(new_n4869_), .Y(new_n15479_));
  AOI21X1  g15415(.A0(new_n14642_), .A1(new_n5097_), .B0(new_n15479_), .Y(new_n15480_));
  OAI21X1  g15416(.A0(new_n14652_), .A1(new_n4868_), .B0(new_n15480_), .Y(new_n15481_));
  XOR2X1   g15417(.A(new_n15481_), .B(new_n2995_), .Y(new_n15482_));
  INVX1    g15418(.A(new_n15482_), .Y(new_n15483_));
  XOR2X1   g15419(.A(new_n15483_), .B(new_n15478_), .Y(new_n15484_));
  XOR2X1   g15420(.A(new_n15484_), .B(new_n15389_), .Y(new_n15485_));
  XOR2X1   g15421(.A(new_n15485_), .B(new_n15385_), .Y(new_n15486_));
  AOI22X1  g15422(.A0(new_n15362_), .A1(new_n11219_), .B0(new_n15234_), .B1(new_n5970_), .Y(new_n15487_));
  OAI21X1  g15423(.A0(new_n15373_), .A1(new_n6298_), .B0(new_n15487_), .Y(new_n15488_));
  XOR2X1   g15424(.A(new_n15488_), .B(new_n3431_), .Y(new_n15489_));
  XOR2X1   g15425(.A(new_n15489_), .B(new_n15486_), .Y(new_n15490_));
  NOR2X1   g15426(.A(new_n15351_), .B(new_n15255_), .Y(new_n15491_));
  INVX1    g15427(.A(new_n15354_), .Y(new_n15492_));
  AOI21X1  g15428(.A0(new_n15492_), .A1(new_n15352_), .B0(new_n15491_), .Y(new_n15493_));
  XOR2X1   g15429(.A(new_n15493_), .B(new_n15490_), .Y(new_n15494_));
  OR2X1    g15430(.A(new_n15376_), .B(new_n15355_), .Y(new_n15495_));
  OAI21X1  g15431(.A0(new_n15250_), .A1(new_n15249_), .B0(new_n15377_), .Y(new_n15496_));
  AND2X1   g15432(.A(new_n15496_), .B(new_n15495_), .Y(new_n15497_));
  XOR2X1   g15433(.A(new_n15497_), .B(new_n15494_), .Y(new_n15498_));
  XOR2X1   g15434(.A(new_n15498_), .B(new_n15380_), .Y(\result[6] ));
  NAND2X1  g15435(.A(new_n15498_), .B(new_n15380_), .Y(new_n15500_));
  INVX1    g15436(.A(new_n15415_), .Y(new_n15501_));
  NOR2X1   g15437(.A(new_n15440_), .B(new_n15436_), .Y(new_n15502_));
  AOI21X1  g15438(.A0(new_n15441_), .A1(new_n15501_), .B0(new_n15502_), .Y(new_n15503_));
  INVX1    g15439(.A(new_n15503_), .Y(new_n15504_));
  AOI22X1  g15440(.A0(new_n12138_), .A1(new_n1890_), .B0(new_n12133_), .B1(new_n1884_), .Y(new_n15505_));
  OAI21X1  g15441(.A0(new_n12117_), .A1(new_n3498_), .B0(new_n15505_), .Y(new_n15506_));
  AOI21X1  g15442(.A0(new_n12526_), .A1(new_n407_), .B0(new_n15506_), .Y(new_n15507_));
  INVX1    g15443(.A(new_n15507_), .Y(new_n15508_));
  NOR4X1   g15444(.A(new_n3779_), .B(new_n1094_), .C(new_n421_), .D(new_n208_), .Y(new_n15509_));
  NOR4X1   g15445(.A(new_n1599_), .B(new_n1416_), .C(new_n1227_), .D(new_n1205_), .Y(new_n15510_));
  OR4X1    g15446(.A(new_n586_), .B(new_n197_), .C(new_n176_), .D(new_n137_), .Y(new_n15511_));
  NOR4X1   g15447(.A(new_n15511_), .B(new_n1090_), .C(new_n141_), .D(new_n338_), .Y(new_n15512_));
  NAND4X1  g15448(.A(new_n15512_), .B(new_n15510_), .C(new_n15509_), .D(new_n7386_), .Y(new_n15513_));
  INVX1    g15449(.A(new_n260_), .Y(new_n15514_));
  INVX1    g15450(.A(new_n261_), .Y(new_n15515_));
  NAND3X1  g15451(.A(new_n15515_), .B(new_n15514_), .C(new_n1150_), .Y(new_n15516_));
  OR4X1    g15452(.A(new_n2363_), .B(new_n1349_), .C(new_n266_), .D(new_n15516_), .Y(new_n15517_));
  NOR4X1   g15453(.A(new_n15517_), .B(new_n15513_), .C(new_n2264_), .D(new_n1654_), .Y(new_n15518_));
  INVX1    g15454(.A(new_n15518_), .Y(new_n15519_));
  AOI21X1  g15455(.A0(new_n15362_), .A1(new_n8170_), .B0(new_n3431_), .Y(new_n15520_));
  INVX1    g15456(.A(new_n15361_), .Y(new_n15521_));
  XOR2X1   g15457(.A(new_n15521_), .B(new_n15358_), .Y(new_n15522_));
  NOR3X1   g15458(.A(new_n15522_), .B(new_n8169_), .C(\a[2] ), .Y(new_n15523_));
  NOR3X1   g15459(.A(new_n15523_), .B(new_n15520_), .C(new_n15519_), .Y(new_n15524_));
  OAI21X1  g15460(.A0(new_n15522_), .A1(new_n8169_), .B0(\a[2] ), .Y(new_n15525_));
  NAND3X1  g15461(.A(new_n15362_), .B(new_n8170_), .C(new_n3431_), .Y(new_n15526_));
  AOI21X1  g15462(.A0(new_n15526_), .A1(new_n15525_), .B0(new_n15518_), .Y(new_n15527_));
  OAI21X1  g15463(.A0(new_n15527_), .A1(new_n15524_), .B0(new_n15508_), .Y(new_n15528_));
  NAND3X1  g15464(.A(new_n15526_), .B(new_n15525_), .C(new_n15518_), .Y(new_n15529_));
  OAI21X1  g15465(.A0(new_n15523_), .A1(new_n15520_), .B0(new_n15519_), .Y(new_n15530_));
  NAND3X1  g15466(.A(new_n15530_), .B(new_n15529_), .C(new_n15507_), .Y(new_n15531_));
  INVX1    g15467(.A(new_n15420_), .Y(new_n15532_));
  NOR2X1   g15468(.A(new_n15434_), .B(new_n15430_), .Y(new_n15533_));
  INVX1    g15469(.A(new_n15533_), .Y(new_n15534_));
  OAI21X1  g15470(.A0(new_n15435_), .A1(new_n15532_), .B0(new_n15534_), .Y(new_n15535_));
  INVX1    g15471(.A(new_n15535_), .Y(new_n15536_));
  NAND3X1  g15472(.A(new_n15536_), .B(new_n15531_), .C(new_n15528_), .Y(new_n15537_));
  AOI21X1  g15473(.A0(new_n15530_), .A1(new_n15529_), .B0(new_n15507_), .Y(new_n15538_));
  NOR3X1   g15474(.A(new_n15527_), .B(new_n15524_), .C(new_n15508_), .Y(new_n15539_));
  OAI21X1  g15475(.A0(new_n15539_), .A1(new_n15538_), .B0(new_n15535_), .Y(new_n15540_));
  OAI22X1  g15476(.A0(new_n12113_), .A1(new_n2186_), .B0(new_n12111_), .B1(new_n2431_), .Y(new_n15541_));
  AOI21X1  g15477(.A0(new_n12107_), .A1(new_n2139_), .B0(new_n15541_), .Y(new_n15542_));
  OAI21X1  g15478(.A0(new_n12708_), .A1(new_n2063_), .B0(new_n15542_), .Y(new_n15543_));
  XOR2X1   g15479(.A(new_n15543_), .B(new_n74_), .Y(new_n15544_));
  INVX1    g15480(.A(new_n15544_), .Y(new_n15545_));
  NAND3X1  g15481(.A(new_n15545_), .B(new_n15540_), .C(new_n15537_), .Y(new_n15546_));
  NOR3X1   g15482(.A(new_n15535_), .B(new_n15539_), .C(new_n15538_), .Y(new_n15547_));
  AOI21X1  g15483(.A0(new_n15531_), .A1(new_n15528_), .B0(new_n15536_), .Y(new_n15548_));
  OAI21X1  g15484(.A0(new_n15548_), .A1(new_n15547_), .B0(new_n15544_), .Y(new_n15549_));
  NAND3X1  g15485(.A(new_n15549_), .B(new_n15546_), .C(new_n15504_), .Y(new_n15550_));
  NOR3X1   g15486(.A(new_n15544_), .B(new_n15548_), .C(new_n15547_), .Y(new_n15551_));
  AOI21X1  g15487(.A0(new_n15540_), .A1(new_n15537_), .B0(new_n15545_), .Y(new_n15552_));
  OAI21X1  g15488(.A0(new_n15552_), .A1(new_n15551_), .B0(new_n15503_), .Y(new_n15553_));
  AOI22X1  g15489(.A0(new_n12104_), .A1(new_n2424_), .B0(new_n12102_), .B1(new_n2418_), .Y(new_n15554_));
  OAI21X1  g15490(.A0(new_n12840_), .A1(new_n2626_), .B0(new_n15554_), .Y(new_n15555_));
  AOI21X1  g15491(.A0(new_n12859_), .A1(new_n2301_), .B0(new_n15555_), .Y(new_n15556_));
  XOR2X1   g15492(.A(new_n15556_), .B(\a[26] ), .Y(new_n15557_));
  NAND3X1  g15493(.A(new_n15557_), .B(new_n15553_), .C(new_n15550_), .Y(new_n15558_));
  NOR3X1   g15494(.A(new_n15552_), .B(new_n15551_), .C(new_n15503_), .Y(new_n15559_));
  AOI21X1  g15495(.A0(new_n15549_), .A1(new_n15546_), .B0(new_n15504_), .Y(new_n15560_));
  INVX1    g15496(.A(new_n15557_), .Y(new_n15561_));
  OAI21X1  g15497(.A0(new_n15560_), .A1(new_n15559_), .B0(new_n15561_), .Y(new_n15562_));
  NOR2X1   g15498(.A(new_n15446_), .B(new_n15442_), .Y(new_n15563_));
  AOI21X1  g15499(.A0(new_n15447_), .A1(new_n15413_), .B0(new_n15563_), .Y(new_n15564_));
  NAND3X1  g15500(.A(new_n15564_), .B(new_n15562_), .C(new_n15558_), .Y(new_n15565_));
  NOR3X1   g15501(.A(new_n15561_), .B(new_n15560_), .C(new_n15559_), .Y(new_n15566_));
  AOI21X1  g15502(.A0(new_n15553_), .A1(new_n15550_), .B0(new_n15557_), .Y(new_n15567_));
  INVX1    g15503(.A(new_n15564_), .Y(new_n15568_));
  OAI21X1  g15504(.A0(new_n15567_), .A1(new_n15566_), .B0(new_n15568_), .Y(new_n15569_));
  AOI22X1  g15505(.A0(new_n12097_), .A1(new_n2657_), .B0(new_n12095_), .B1(new_n2696_), .Y(new_n15570_));
  OAI21X1  g15506(.A0(new_n13366_), .A1(new_n2753_), .B0(new_n15570_), .Y(new_n15571_));
  AOI21X1  g15507(.A0(new_n13093_), .A1(new_n2658_), .B0(new_n15571_), .Y(new_n15572_));
  XOR2X1   g15508(.A(new_n15572_), .B(\a[23] ), .Y(new_n15573_));
  NAND3X1  g15509(.A(new_n15573_), .B(new_n15569_), .C(new_n15565_), .Y(new_n15574_));
  NOR3X1   g15510(.A(new_n15568_), .B(new_n15567_), .C(new_n15566_), .Y(new_n15575_));
  AOI21X1  g15511(.A0(new_n15562_), .A1(new_n15558_), .B0(new_n15564_), .Y(new_n15576_));
  INVX1    g15512(.A(new_n15573_), .Y(new_n15577_));
  OAI21X1  g15513(.A0(new_n15576_), .A1(new_n15575_), .B0(new_n15577_), .Y(new_n15578_));
  INVX1    g15514(.A(new_n15410_), .Y(new_n15579_));
  AND2X1   g15515(.A(new_n15448_), .B(new_n15579_), .Y(new_n15580_));
  AOI21X1  g15516(.A0(new_n15452_), .A1(new_n15450_), .B0(new_n15580_), .Y(new_n15581_));
  NAND3X1  g15517(.A(new_n15581_), .B(new_n15578_), .C(new_n15574_), .Y(new_n15582_));
  NOR3X1   g15518(.A(new_n15577_), .B(new_n15576_), .C(new_n15575_), .Y(new_n15583_));
  AOI21X1  g15519(.A0(new_n15569_), .A1(new_n15565_), .B0(new_n15573_), .Y(new_n15584_));
  INVX1    g15520(.A(new_n15581_), .Y(new_n15585_));
  OAI21X1  g15521(.A0(new_n15584_), .A1(new_n15583_), .B0(new_n15585_), .Y(new_n15586_));
  AOI22X1  g15522(.A0(new_n12090_), .A1(new_n2875_), .B0(new_n12088_), .B1(new_n3099_), .Y(new_n15587_));
  OAI21X1  g15523(.A0(new_n12298_), .A1(new_n3152_), .B0(new_n15587_), .Y(new_n15588_));
  AOI21X1  g15524(.A0(new_n12297_), .A1(new_n2876_), .B0(new_n15588_), .Y(new_n15589_));
  XOR2X1   g15525(.A(new_n15589_), .B(\a[20] ), .Y(new_n15590_));
  NAND3X1  g15526(.A(new_n15590_), .B(new_n15586_), .C(new_n15582_), .Y(new_n15591_));
  NOR3X1   g15527(.A(new_n15585_), .B(new_n15584_), .C(new_n15583_), .Y(new_n15592_));
  AOI21X1  g15528(.A0(new_n15578_), .A1(new_n15574_), .B0(new_n15581_), .Y(new_n15593_));
  INVX1    g15529(.A(new_n15590_), .Y(new_n15594_));
  OAI21X1  g15530(.A0(new_n15593_), .A1(new_n15592_), .B0(new_n15594_), .Y(new_n15595_));
  NOR2X1   g15531(.A(new_n15458_), .B(new_n15454_), .Y(new_n15596_));
  AOI21X1  g15532(.A0(new_n15459_), .A1(new_n15406_), .B0(new_n15596_), .Y(new_n15597_));
  NAND3X1  g15533(.A(new_n15597_), .B(new_n15595_), .C(new_n15591_), .Y(new_n15598_));
  NOR3X1   g15534(.A(new_n15594_), .B(new_n15593_), .C(new_n15592_), .Y(new_n15599_));
  AOI21X1  g15535(.A0(new_n15586_), .A1(new_n15582_), .B0(new_n15590_), .Y(new_n15600_));
  INVX1    g15536(.A(new_n15597_), .Y(new_n15601_));
  OAI21X1  g15537(.A0(new_n15600_), .A1(new_n15599_), .B0(new_n15601_), .Y(new_n15602_));
  AOI22X1  g15538(.A0(new_n12083_), .A1(new_n3232_), .B0(new_n12081_), .B1(new_n3390_), .Y(new_n15603_));
  OAI21X1  g15539(.A0(new_n13665_), .A1(new_n3545_), .B0(new_n15603_), .Y(new_n15604_));
  AOI21X1  g15540(.A0(new_n14672_), .A1(new_n3234_), .B0(new_n15604_), .Y(new_n15605_));
  XOR2X1   g15541(.A(new_n15605_), .B(\a[17] ), .Y(new_n15606_));
  NAND3X1  g15542(.A(new_n15606_), .B(new_n15602_), .C(new_n15598_), .Y(new_n15607_));
  NOR3X1   g15543(.A(new_n15601_), .B(new_n15600_), .C(new_n15599_), .Y(new_n15608_));
  AOI21X1  g15544(.A0(new_n15595_), .A1(new_n15591_), .B0(new_n15597_), .Y(new_n15609_));
  INVX1    g15545(.A(new_n15606_), .Y(new_n15610_));
  OAI21X1  g15546(.A0(new_n15609_), .A1(new_n15608_), .B0(new_n15610_), .Y(new_n15611_));
  AND2X1   g15547(.A(new_n15460_), .B(new_n15402_), .Y(new_n15612_));
  AOI21X1  g15548(.A0(new_n15464_), .A1(new_n15461_), .B0(new_n15612_), .Y(new_n15613_));
  NAND3X1  g15549(.A(new_n15613_), .B(new_n15611_), .C(new_n15607_), .Y(new_n15614_));
  NOR3X1   g15550(.A(new_n15610_), .B(new_n15609_), .C(new_n15608_), .Y(new_n15615_));
  AOI21X1  g15551(.A0(new_n15602_), .A1(new_n15598_), .B0(new_n15606_), .Y(new_n15616_));
  INVX1    g15552(.A(new_n15613_), .Y(new_n15617_));
  OAI21X1  g15553(.A0(new_n15616_), .A1(new_n15615_), .B0(new_n15617_), .Y(new_n15618_));
  AOI22X1  g15554(.A0(new_n12076_), .A1(new_n3628_), .B0(new_n12018_), .B1(new_n3908_), .Y(new_n15619_));
  OAI21X1  g15555(.A0(new_n13679_), .A1(new_n3983_), .B0(new_n15619_), .Y(new_n15620_));
  AOI21X1  g15556(.A0(new_n13678_), .A1(new_n3624_), .B0(new_n15620_), .Y(new_n15621_));
  XOR2X1   g15557(.A(new_n15621_), .B(\a[14] ), .Y(new_n15622_));
  NAND3X1  g15558(.A(new_n15622_), .B(new_n15618_), .C(new_n15614_), .Y(new_n15623_));
  NOR3X1   g15559(.A(new_n15617_), .B(new_n15616_), .C(new_n15615_), .Y(new_n15624_));
  AOI21X1  g15560(.A0(new_n15611_), .A1(new_n15607_), .B0(new_n15613_), .Y(new_n15625_));
  INVX1    g15561(.A(new_n15622_), .Y(new_n15626_));
  OAI21X1  g15562(.A0(new_n15625_), .A1(new_n15624_), .B0(new_n15626_), .Y(new_n15627_));
  AND2X1   g15563(.A(new_n15470_), .B(new_n15465_), .Y(new_n15628_));
  AOI21X1  g15564(.A0(new_n15471_), .A1(new_n15397_), .B0(new_n15628_), .Y(new_n15629_));
  NAND3X1  g15565(.A(new_n15629_), .B(new_n15627_), .C(new_n15623_), .Y(new_n15630_));
  NOR3X1   g15566(.A(new_n15626_), .B(new_n15625_), .C(new_n15624_), .Y(new_n15631_));
  AOI21X1  g15567(.A0(new_n15618_), .A1(new_n15614_), .B0(new_n15622_), .Y(new_n15632_));
  INVX1    g15568(.A(new_n15629_), .Y(new_n15633_));
  OAI21X1  g15569(.A0(new_n15632_), .A1(new_n15631_), .B0(new_n15633_), .Y(new_n15634_));
  AOI22X1  g15570(.A0(new_n14085_), .A1(new_n4247_), .B0(new_n12285_), .B1(new_n4078_), .Y(new_n15635_));
  OAI21X1  g15571(.A0(new_n14088_), .A1(new_n4427_), .B0(new_n15635_), .Y(new_n15636_));
  AOI21X1  g15572(.A0(new_n14491_), .A1(new_n4080_), .B0(new_n15636_), .Y(new_n15637_));
  XOR2X1   g15573(.A(new_n15637_), .B(\a[11] ), .Y(new_n15638_));
  NAND3X1  g15574(.A(new_n15638_), .B(new_n15634_), .C(new_n15630_), .Y(new_n15639_));
  NOR3X1   g15575(.A(new_n15633_), .B(new_n15632_), .C(new_n15631_), .Y(new_n15640_));
  AOI21X1  g15576(.A0(new_n15627_), .A1(new_n15623_), .B0(new_n15629_), .Y(new_n15641_));
  INVX1    g15577(.A(new_n15638_), .Y(new_n15642_));
  OAI21X1  g15578(.A0(new_n15641_), .A1(new_n15640_), .B0(new_n15642_), .Y(new_n15643_));
  AND2X1   g15579(.A(new_n15472_), .B(new_n15394_), .Y(new_n15644_));
  AOI21X1  g15580(.A0(new_n15477_), .A1(new_n15473_), .B0(new_n15644_), .Y(new_n15645_));
  NAND3X1  g15581(.A(new_n15645_), .B(new_n15643_), .C(new_n15639_), .Y(new_n15646_));
  NOR3X1   g15582(.A(new_n15642_), .B(new_n15641_), .C(new_n15640_), .Y(new_n15647_));
  AOI21X1  g15583(.A0(new_n15634_), .A1(new_n15630_), .B0(new_n15638_), .Y(new_n15648_));
  INVX1    g15584(.A(new_n15645_), .Y(new_n15649_));
  OAI21X1  g15585(.A0(new_n15648_), .A1(new_n15647_), .B0(new_n15649_), .Y(new_n15650_));
  AOI22X1  g15586(.A0(new_n14642_), .A1(new_n4870_), .B0(new_n14084_), .B1(new_n4635_), .Y(new_n15651_));
  OAI21X1  g15587(.A0(new_n14805_), .A1(new_n5096_), .B0(new_n15651_), .Y(new_n15652_));
  AOI21X1  g15588(.A0(new_n14809_), .A1(new_n4637_), .B0(new_n15652_), .Y(new_n15653_));
  XOR2X1   g15589(.A(new_n15653_), .B(\a[8] ), .Y(new_n15654_));
  NAND3X1  g15590(.A(new_n15654_), .B(new_n15650_), .C(new_n15646_), .Y(new_n15655_));
  NOR3X1   g15591(.A(new_n15649_), .B(new_n15648_), .C(new_n15647_), .Y(new_n15656_));
  AOI21X1  g15592(.A0(new_n15643_), .A1(new_n15639_), .B0(new_n15645_), .Y(new_n15657_));
  INVX1    g15593(.A(new_n15654_), .Y(new_n15658_));
  OAI21X1  g15594(.A0(new_n15657_), .A1(new_n15656_), .B0(new_n15658_), .Y(new_n15659_));
  AND2X1   g15595(.A(new_n15483_), .B(new_n15478_), .Y(new_n15660_));
  AOI21X1  g15596(.A0(new_n15484_), .A1(new_n15389_), .B0(new_n15660_), .Y(new_n15661_));
  NAND3X1  g15597(.A(new_n15661_), .B(new_n15659_), .C(new_n15655_), .Y(new_n15662_));
  NOR3X1   g15598(.A(new_n15658_), .B(new_n15657_), .C(new_n15656_), .Y(new_n15663_));
  AOI21X1  g15599(.A0(new_n15650_), .A1(new_n15646_), .B0(new_n15654_), .Y(new_n15664_));
  INVX1    g15600(.A(new_n15661_), .Y(new_n15665_));
  OAI21X1  g15601(.A0(new_n15664_), .A1(new_n15663_), .B0(new_n15665_), .Y(new_n15666_));
  AOI22X1  g15602(.A0(new_n15087_), .A1(new_n5659_), .B0(new_n14946_), .B1(new_n5373_), .Y(new_n15667_));
  OAI21X1  g15603(.A0(new_n15363_), .A1(new_n5959_), .B0(new_n15667_), .Y(new_n15668_));
  AOI21X1  g15604(.A0(new_n15240_), .A1(new_n67_), .B0(new_n15668_), .Y(new_n15669_));
  XOR2X1   g15605(.A(new_n15669_), .B(\a[5] ), .Y(new_n15670_));
  NAND3X1  g15606(.A(new_n15670_), .B(new_n15666_), .C(new_n15662_), .Y(new_n15671_));
  NOR3X1   g15607(.A(new_n15665_), .B(new_n15664_), .C(new_n15663_), .Y(new_n15672_));
  AOI21X1  g15608(.A0(new_n15659_), .A1(new_n15655_), .B0(new_n15661_), .Y(new_n15673_));
  INVX1    g15609(.A(new_n15670_), .Y(new_n15674_));
  OAI21X1  g15610(.A0(new_n15673_), .A1(new_n15672_), .B0(new_n15674_), .Y(new_n15675_));
  XOR2X1   g15611(.A(new_n15384_), .B(new_n3289_), .Y(new_n15676_));
  AND2X1   g15612(.A(new_n15485_), .B(new_n15676_), .Y(new_n15677_));
  NOR2X1   g15613(.A(new_n15489_), .B(new_n15486_), .Y(new_n15678_));
  NOR2X1   g15614(.A(new_n15678_), .B(new_n15677_), .Y(new_n15679_));
  NAND3X1  g15615(.A(new_n15679_), .B(new_n15675_), .C(new_n15671_), .Y(new_n15680_));
  NOR3X1   g15616(.A(new_n15674_), .B(new_n15673_), .C(new_n15672_), .Y(new_n15681_));
  AOI21X1  g15617(.A0(new_n15666_), .A1(new_n15662_), .B0(new_n15670_), .Y(new_n15682_));
  INVX1    g15618(.A(new_n15679_), .Y(new_n15683_));
  OAI21X1  g15619(.A0(new_n15682_), .A1(new_n15681_), .B0(new_n15683_), .Y(new_n15684_));
  AND2X1   g15620(.A(new_n15684_), .B(new_n15680_), .Y(new_n15685_));
  INVX1    g15621(.A(new_n15493_), .Y(new_n15686_));
  AND2X1   g15622(.A(new_n15686_), .B(new_n15490_), .Y(new_n15687_));
  AOI21X1  g15623(.A0(new_n15496_), .A1(new_n15495_), .B0(new_n15494_), .Y(new_n15688_));
  NOR2X1   g15624(.A(new_n15688_), .B(new_n15687_), .Y(new_n15689_));
  XOR2X1   g15625(.A(new_n15689_), .B(new_n15685_), .Y(new_n15690_));
  XOR2X1   g15626(.A(new_n15690_), .B(new_n15500_), .Y(\result[7] ));
  NOR2X1   g15627(.A(new_n15690_), .B(new_n15500_), .Y(new_n15692_));
  OAI21X1  g15628(.A0(new_n15524_), .A1(new_n15507_), .B0(new_n15530_), .Y(new_n15693_));
  AND2X1   g15629(.A(new_n15362_), .B(new_n8170_), .Y(new_n15694_));
  XOR2X1   g15630(.A(new_n15694_), .B(\a[2] ), .Y(new_n15695_));
  NOR2X1   g15631(.A(new_n1030_), .B(new_n1027_), .Y(new_n15696_));
  OR4X1    g15632(.A(new_n634_), .B(new_n540_), .C(new_n158_), .D(new_n100_), .Y(new_n15697_));
  NOR4X1   g15633(.A(new_n15697_), .B(new_n12657_), .C(new_n170_), .D(new_n164_), .Y(new_n15698_));
  OR4X1    g15634(.A(new_n414_), .B(new_n843_), .C(new_n299_), .D(new_n282_), .Y(new_n15699_));
  OR4X1    g15635(.A(new_n830_), .B(new_n607_), .C(new_n3731_), .D(new_n209_), .Y(new_n15700_));
  NOR4X1   g15636(.A(new_n15700_), .B(new_n15699_), .C(new_n1962_), .D(new_n1588_), .Y(new_n15701_));
  OR4X1    g15637(.A(new_n714_), .B(new_n239_), .C(new_n194_), .D(new_n825_), .Y(new_n15702_));
  NOR4X1   g15638(.A(new_n15702_), .B(new_n395_), .C(new_n307_), .D(new_n86_), .Y(new_n15703_));
  NAND4X1  g15639(.A(new_n15703_), .B(new_n15701_), .C(new_n15698_), .D(new_n15696_), .Y(new_n15704_));
  NOR3X1   g15640(.A(new_n15704_), .B(new_n8743_), .C(new_n1454_), .Y(new_n15705_));
  XOR2X1   g15641(.A(new_n15705_), .B(new_n15695_), .Y(new_n15706_));
  AND2X1   g15642(.A(new_n15706_), .B(new_n15693_), .Y(new_n15707_));
  AOI21X1  g15643(.A0(new_n15526_), .A1(new_n15525_), .B0(new_n15705_), .Y(new_n15708_));
  XOR2X1   g15644(.A(new_n15694_), .B(new_n3431_), .Y(new_n15709_));
  AND2X1   g15645(.A(new_n15705_), .B(new_n15709_), .Y(new_n15710_));
  NOR3X1   g15646(.A(new_n15710_), .B(new_n15708_), .C(new_n15693_), .Y(new_n15711_));
  AOI22X1  g15647(.A0(new_n12133_), .A1(new_n1890_), .B0(new_n12720_), .B1(new_n1884_), .Y(new_n15712_));
  OAI21X1  g15648(.A0(new_n12113_), .A1(new_n3498_), .B0(new_n15712_), .Y(new_n15713_));
  AOI21X1  g15649(.A0(new_n12719_), .A1(new_n407_), .B0(new_n15713_), .Y(new_n15714_));
  OAI21X1  g15650(.A0(new_n15711_), .A1(new_n15707_), .B0(new_n15714_), .Y(new_n15715_));
  NAND2X1  g15651(.A(new_n15706_), .B(new_n15693_), .Y(new_n15716_));
  NOR3X1   g15652(.A(new_n15527_), .B(new_n15524_), .C(new_n15507_), .Y(new_n15717_));
  OR4X1    g15653(.A(new_n15710_), .B(new_n15708_), .C(new_n15717_), .D(new_n15527_), .Y(new_n15718_));
  INVX1    g15654(.A(new_n15714_), .Y(new_n15719_));
  NAND3X1  g15655(.A(new_n15719_), .B(new_n15718_), .C(new_n15716_), .Y(new_n15720_));
  AOI21X1  g15656(.A0(new_n15545_), .A1(new_n15537_), .B0(new_n15548_), .Y(new_n15721_));
  NAND3X1  g15657(.A(new_n15721_), .B(new_n15720_), .C(new_n15715_), .Y(new_n15722_));
  AOI21X1  g15658(.A0(new_n15718_), .A1(new_n15716_), .B0(new_n15719_), .Y(new_n15723_));
  NOR3X1   g15659(.A(new_n15714_), .B(new_n15711_), .C(new_n15707_), .Y(new_n15724_));
  OAI21X1  g15660(.A0(new_n15544_), .A1(new_n15547_), .B0(new_n15540_), .Y(new_n15725_));
  OAI21X1  g15661(.A0(new_n15724_), .A1(new_n15723_), .B0(new_n15725_), .Y(new_n15726_));
  AOI22X1  g15662(.A0(new_n12208_), .A1(new_n2185_), .B0(new_n12107_), .B1(new_n2095_), .Y(new_n15727_));
  OAI21X1  g15663(.A0(new_n12695_), .A1(new_n2140_), .B0(new_n15727_), .Y(new_n15728_));
  AOI21X1  g15664(.A0(new_n12694_), .A1(new_n2062_), .B0(new_n15728_), .Y(new_n15729_));
  XOR2X1   g15665(.A(new_n15729_), .B(\a[29] ), .Y(new_n15730_));
  NAND3X1  g15666(.A(new_n15730_), .B(new_n15726_), .C(new_n15722_), .Y(new_n15731_));
  NOR3X1   g15667(.A(new_n15725_), .B(new_n15724_), .C(new_n15723_), .Y(new_n15732_));
  AOI21X1  g15668(.A0(new_n15720_), .A1(new_n15715_), .B0(new_n15721_), .Y(new_n15733_));
  INVX1    g15669(.A(new_n15730_), .Y(new_n15734_));
  OAI21X1  g15670(.A0(new_n15733_), .A1(new_n15732_), .B0(new_n15734_), .Y(new_n15735_));
  AOI22X1  g15671(.A0(new_n12102_), .A1(new_n2424_), .B0(new_n12099_), .B1(new_n2418_), .Y(new_n15736_));
  OAI21X1  g15672(.A0(new_n12839_), .A1(new_n2626_), .B0(new_n15736_), .Y(new_n15737_));
  AOI21X1  g15673(.A0(new_n12855_), .A1(new_n2301_), .B0(new_n15737_), .Y(new_n15738_));
  XOR2X1   g15674(.A(new_n15738_), .B(\a[26] ), .Y(new_n15739_));
  INVX1    g15675(.A(new_n15739_), .Y(new_n15740_));
  AOI21X1  g15676(.A0(new_n15735_), .A1(new_n15731_), .B0(new_n15740_), .Y(new_n15741_));
  NOR3X1   g15677(.A(new_n15734_), .B(new_n15733_), .C(new_n15732_), .Y(new_n15742_));
  AOI21X1  g15678(.A0(new_n15726_), .A1(new_n15722_), .B0(new_n15730_), .Y(new_n15743_));
  NOR3X1   g15679(.A(new_n15739_), .B(new_n15743_), .C(new_n15742_), .Y(new_n15744_));
  OAI21X1  g15680(.A0(new_n15557_), .A1(new_n15560_), .B0(new_n15550_), .Y(new_n15745_));
  NOR3X1   g15681(.A(new_n15745_), .B(new_n15744_), .C(new_n15741_), .Y(new_n15746_));
  OAI21X1  g15682(.A0(new_n15743_), .A1(new_n15742_), .B0(new_n15739_), .Y(new_n15747_));
  NAND3X1  g15683(.A(new_n15740_), .B(new_n15735_), .C(new_n15731_), .Y(new_n15748_));
  AOI21X1  g15684(.A0(new_n15561_), .A1(new_n15553_), .B0(new_n15559_), .Y(new_n15749_));
  AOI21X1  g15685(.A0(new_n15748_), .A1(new_n15747_), .B0(new_n15749_), .Y(new_n15750_));
  AOI22X1  g15686(.A0(new_n12095_), .A1(new_n2657_), .B0(new_n12093_), .B1(new_n2696_), .Y(new_n15751_));
  OAI21X1  g15687(.A0(new_n13118_), .A1(new_n2753_), .B0(new_n15751_), .Y(new_n15752_));
  AOI21X1  g15688(.A0(new_n13117_), .A1(new_n2658_), .B0(new_n15752_), .Y(new_n15753_));
  XOR2X1   g15689(.A(new_n15753_), .B(\a[23] ), .Y(new_n15754_));
  INVX1    g15690(.A(new_n15754_), .Y(new_n15755_));
  NOR3X1   g15691(.A(new_n15755_), .B(new_n15750_), .C(new_n15746_), .Y(new_n15756_));
  NAND3X1  g15692(.A(new_n15749_), .B(new_n15748_), .C(new_n15747_), .Y(new_n15757_));
  OAI21X1  g15693(.A0(new_n15744_), .A1(new_n15741_), .B0(new_n15745_), .Y(new_n15758_));
  AOI21X1  g15694(.A0(new_n15758_), .A1(new_n15757_), .B0(new_n15754_), .Y(new_n15759_));
  OAI21X1  g15695(.A0(new_n15573_), .A1(new_n15575_), .B0(new_n15569_), .Y(new_n15760_));
  NOR3X1   g15696(.A(new_n15760_), .B(new_n15759_), .C(new_n15756_), .Y(new_n15761_));
  NAND3X1  g15697(.A(new_n15754_), .B(new_n15758_), .C(new_n15757_), .Y(new_n15762_));
  OAI21X1  g15698(.A0(new_n15750_), .A1(new_n15746_), .B0(new_n15755_), .Y(new_n15763_));
  AOI21X1  g15699(.A0(new_n15577_), .A1(new_n15565_), .B0(new_n15576_), .Y(new_n15764_));
  AOI21X1  g15700(.A0(new_n15763_), .A1(new_n15762_), .B0(new_n15764_), .Y(new_n15765_));
  AOI22X1  g15701(.A0(new_n12088_), .A1(new_n2875_), .B0(new_n12085_), .B1(new_n3099_), .Y(new_n15766_));
  OAI21X1  g15702(.A0(new_n13321_), .A1(new_n3152_), .B0(new_n15766_), .Y(new_n15767_));
  AOI21X1  g15703(.A0(new_n13344_), .A1(new_n2876_), .B0(new_n15767_), .Y(new_n15768_));
  XOR2X1   g15704(.A(new_n15768_), .B(\a[20] ), .Y(new_n15769_));
  INVX1    g15705(.A(new_n15769_), .Y(new_n15770_));
  NOR3X1   g15706(.A(new_n15770_), .B(new_n15765_), .C(new_n15761_), .Y(new_n15771_));
  NAND3X1  g15707(.A(new_n15764_), .B(new_n15763_), .C(new_n15762_), .Y(new_n15772_));
  OAI21X1  g15708(.A0(new_n15759_), .A1(new_n15756_), .B0(new_n15760_), .Y(new_n15773_));
  AOI21X1  g15709(.A0(new_n15773_), .A1(new_n15772_), .B0(new_n15769_), .Y(new_n15774_));
  OAI21X1  g15710(.A0(new_n15590_), .A1(new_n15592_), .B0(new_n15586_), .Y(new_n15775_));
  NOR3X1   g15711(.A(new_n15775_), .B(new_n15774_), .C(new_n15771_), .Y(new_n15776_));
  NAND3X1  g15712(.A(new_n15769_), .B(new_n15773_), .C(new_n15772_), .Y(new_n15777_));
  OAI21X1  g15713(.A0(new_n15765_), .A1(new_n15761_), .B0(new_n15770_), .Y(new_n15778_));
  AOI21X1  g15714(.A0(new_n15594_), .A1(new_n15582_), .B0(new_n15593_), .Y(new_n15779_));
  AOI21X1  g15715(.A0(new_n15778_), .A1(new_n15777_), .B0(new_n15779_), .Y(new_n15780_));
  AOI22X1  g15716(.A0(new_n12081_), .A1(new_n3232_), .B0(new_n12079_), .B1(new_n3390_), .Y(new_n15781_));
  OAI21X1  g15717(.A0(new_n13700_), .A1(new_n3545_), .B0(new_n15781_), .Y(new_n15782_));
  AOI21X1  g15718(.A0(new_n13699_), .A1(new_n3234_), .B0(new_n15782_), .Y(new_n15783_));
  XOR2X1   g15719(.A(new_n15783_), .B(\a[17] ), .Y(new_n15784_));
  INVX1    g15720(.A(new_n15784_), .Y(new_n15785_));
  NOR3X1   g15721(.A(new_n15785_), .B(new_n15780_), .C(new_n15776_), .Y(new_n15786_));
  NAND3X1  g15722(.A(new_n15779_), .B(new_n15778_), .C(new_n15777_), .Y(new_n15787_));
  OAI21X1  g15723(.A0(new_n15774_), .A1(new_n15771_), .B0(new_n15775_), .Y(new_n15788_));
  AOI21X1  g15724(.A0(new_n15788_), .A1(new_n15787_), .B0(new_n15784_), .Y(new_n15789_));
  OAI21X1  g15725(.A0(new_n15606_), .A1(new_n15608_), .B0(new_n15602_), .Y(new_n15790_));
  NOR3X1   g15726(.A(new_n15790_), .B(new_n15789_), .C(new_n15786_), .Y(new_n15791_));
  NAND3X1  g15727(.A(new_n15784_), .B(new_n15788_), .C(new_n15787_), .Y(new_n15792_));
  OAI21X1  g15728(.A0(new_n15780_), .A1(new_n15776_), .B0(new_n15785_), .Y(new_n15793_));
  AOI21X1  g15729(.A0(new_n15610_), .A1(new_n15598_), .B0(new_n15609_), .Y(new_n15794_));
  AOI21X1  g15730(.A0(new_n15793_), .A1(new_n15792_), .B0(new_n15794_), .Y(new_n15795_));
  AOI22X1  g15731(.A0(new_n12074_), .A1(new_n3908_), .B0(new_n12018_), .B1(new_n3628_), .Y(new_n15796_));
  OAI21X1  g15732(.A0(new_n12292_), .A1(new_n3983_), .B0(new_n15796_), .Y(new_n15797_));
  AOI21X1  g15733(.A0(new_n12291_), .A1(new_n3624_), .B0(new_n15797_), .Y(new_n15798_));
  XOR2X1   g15734(.A(new_n15798_), .B(\a[14] ), .Y(new_n15799_));
  INVX1    g15735(.A(new_n15799_), .Y(new_n15800_));
  NOR3X1   g15736(.A(new_n15800_), .B(new_n15795_), .C(new_n15791_), .Y(new_n15801_));
  NAND3X1  g15737(.A(new_n15794_), .B(new_n15793_), .C(new_n15792_), .Y(new_n15802_));
  OAI21X1  g15738(.A0(new_n15789_), .A1(new_n15786_), .B0(new_n15790_), .Y(new_n15803_));
  AOI21X1  g15739(.A0(new_n15803_), .A1(new_n15802_), .B0(new_n15799_), .Y(new_n15804_));
  OAI21X1  g15740(.A0(new_n15622_), .A1(new_n15624_), .B0(new_n15618_), .Y(new_n15805_));
  NOR3X1   g15741(.A(new_n15805_), .B(new_n15804_), .C(new_n15801_), .Y(new_n15806_));
  NAND3X1  g15742(.A(new_n15799_), .B(new_n15803_), .C(new_n15802_), .Y(new_n15807_));
  OAI21X1  g15743(.A0(new_n15795_), .A1(new_n15791_), .B0(new_n15800_), .Y(new_n15808_));
  AOI21X1  g15744(.A0(new_n15626_), .A1(new_n15614_), .B0(new_n15625_), .Y(new_n15809_));
  AOI21X1  g15745(.A0(new_n15808_), .A1(new_n15807_), .B0(new_n15809_), .Y(new_n15810_));
  AOI22X1  g15746(.A0(new_n14087_), .A1(new_n4247_), .B0(new_n14085_), .B1(new_n4078_), .Y(new_n15811_));
  OAI21X1  g15747(.A0(new_n14643_), .A1(new_n4427_), .B0(new_n15811_), .Y(new_n15812_));
  AOI21X1  g15748(.A0(new_n14106_), .A1(new_n4080_), .B0(new_n15812_), .Y(new_n15813_));
  XOR2X1   g15749(.A(new_n15813_), .B(\a[11] ), .Y(new_n15814_));
  INVX1    g15750(.A(new_n15814_), .Y(new_n15815_));
  NOR3X1   g15751(.A(new_n15815_), .B(new_n15810_), .C(new_n15806_), .Y(new_n15816_));
  NAND3X1  g15752(.A(new_n15809_), .B(new_n15808_), .C(new_n15807_), .Y(new_n15817_));
  OAI21X1  g15753(.A0(new_n15804_), .A1(new_n15801_), .B0(new_n15805_), .Y(new_n15818_));
  AOI21X1  g15754(.A0(new_n15818_), .A1(new_n15817_), .B0(new_n15814_), .Y(new_n15819_));
  OAI21X1  g15755(.A0(new_n15638_), .A1(new_n15640_), .B0(new_n15634_), .Y(new_n15820_));
  NOR3X1   g15756(.A(new_n15820_), .B(new_n15819_), .C(new_n15816_), .Y(new_n15821_));
  NAND3X1  g15757(.A(new_n15814_), .B(new_n15818_), .C(new_n15817_), .Y(new_n15822_));
  OAI21X1  g15758(.A0(new_n15810_), .A1(new_n15806_), .B0(new_n15815_), .Y(new_n15823_));
  AOI21X1  g15759(.A0(new_n15642_), .A1(new_n15630_), .B0(new_n15641_), .Y(new_n15824_));
  AOI21X1  g15760(.A0(new_n15823_), .A1(new_n15822_), .B0(new_n15824_), .Y(new_n15825_));
  AOI22X1  g15761(.A0(new_n14804_), .A1(new_n4870_), .B0(new_n14642_), .B1(new_n4635_), .Y(new_n15826_));
  OAI21X1  g15762(.A0(new_n15088_), .A1(new_n5096_), .B0(new_n15826_), .Y(new_n15827_));
  AOI21X1  g15763(.A0(new_n14952_), .A1(new_n4637_), .B0(new_n15827_), .Y(new_n15828_));
  XOR2X1   g15764(.A(new_n15828_), .B(\a[8] ), .Y(new_n15829_));
  INVX1    g15765(.A(new_n15829_), .Y(new_n15830_));
  NOR3X1   g15766(.A(new_n15830_), .B(new_n15825_), .C(new_n15821_), .Y(new_n15831_));
  NAND3X1  g15767(.A(new_n15824_), .B(new_n15823_), .C(new_n15822_), .Y(new_n15832_));
  OAI21X1  g15768(.A0(new_n15819_), .A1(new_n15816_), .B0(new_n15820_), .Y(new_n15833_));
  AOI21X1  g15769(.A0(new_n15833_), .A1(new_n15832_), .B0(new_n15829_), .Y(new_n15834_));
  OAI21X1  g15770(.A0(new_n15654_), .A1(new_n15656_), .B0(new_n15650_), .Y(new_n15835_));
  NOR3X1   g15771(.A(new_n15835_), .B(new_n15834_), .C(new_n15831_), .Y(new_n15836_));
  NAND3X1  g15772(.A(new_n15829_), .B(new_n15833_), .C(new_n15832_), .Y(new_n15837_));
  OAI21X1  g15773(.A0(new_n15825_), .A1(new_n15821_), .B0(new_n15830_), .Y(new_n15838_));
  AOI21X1  g15774(.A0(new_n15658_), .A1(new_n15646_), .B0(new_n15657_), .Y(new_n15839_));
  AOI21X1  g15775(.A0(new_n15838_), .A1(new_n15837_), .B0(new_n15839_), .Y(new_n15840_));
  INVX1    g15776(.A(new_n15374_), .Y(new_n15841_));
  AOI22X1  g15777(.A0(new_n15234_), .A1(new_n5659_), .B0(new_n15087_), .B1(new_n5373_), .Y(new_n15842_));
  OAI21X1  g15778(.A0(new_n15522_), .A1(new_n5959_), .B0(new_n15842_), .Y(new_n15843_));
  AOI21X1  g15779(.A0(new_n15841_), .A1(new_n67_), .B0(new_n15843_), .Y(new_n15844_));
  XOR2X1   g15780(.A(new_n15844_), .B(\a[5] ), .Y(new_n15845_));
  INVX1    g15781(.A(new_n15845_), .Y(new_n15846_));
  NOR3X1   g15782(.A(new_n15846_), .B(new_n15840_), .C(new_n15836_), .Y(new_n15847_));
  NAND3X1  g15783(.A(new_n15839_), .B(new_n15838_), .C(new_n15837_), .Y(new_n15848_));
  OAI21X1  g15784(.A0(new_n15834_), .A1(new_n15831_), .B0(new_n15835_), .Y(new_n15849_));
  AOI21X1  g15785(.A0(new_n15849_), .A1(new_n15848_), .B0(new_n15845_), .Y(new_n15850_));
  OAI21X1  g15786(.A0(new_n15670_), .A1(new_n15672_), .B0(new_n15666_), .Y(new_n15851_));
  NOR3X1   g15787(.A(new_n15851_), .B(new_n15850_), .C(new_n15847_), .Y(new_n15852_));
  NAND3X1  g15788(.A(new_n15845_), .B(new_n15849_), .C(new_n15848_), .Y(new_n15853_));
  OAI21X1  g15789(.A0(new_n15840_), .A1(new_n15836_), .B0(new_n15846_), .Y(new_n15854_));
  AOI21X1  g15790(.A0(new_n15674_), .A1(new_n15662_), .B0(new_n15673_), .Y(new_n15855_));
  AOI21X1  g15791(.A0(new_n15854_), .A1(new_n15853_), .B0(new_n15855_), .Y(new_n15856_));
  OR2X1    g15792(.A(new_n15856_), .B(new_n15852_), .Y(new_n15857_));
  AOI21X1  g15793(.A0(new_n15675_), .A1(new_n15671_), .B0(new_n15679_), .Y(new_n15858_));
  OR2X1    g15794(.A(new_n15688_), .B(new_n15687_), .Y(new_n15859_));
  AOI21X1  g15795(.A0(new_n15859_), .A1(new_n15680_), .B0(new_n15858_), .Y(new_n15860_));
  XOR2X1   g15796(.A(new_n15860_), .B(new_n15857_), .Y(new_n15861_));
  XOR2X1   g15797(.A(new_n15861_), .B(new_n15692_), .Y(\result[8] ));
  NAND2X1  g15798(.A(new_n15861_), .B(new_n15692_), .Y(new_n15863_));
  NAND3X1  g15799(.A(new_n15705_), .B(new_n15526_), .C(new_n15525_), .Y(new_n15864_));
  AOI21X1  g15800(.A0(new_n15864_), .A1(new_n15693_), .B0(new_n15708_), .Y(new_n15865_));
  OR4X1    g15801(.A(new_n1724_), .B(new_n1600_), .C(new_n959_), .D(new_n904_), .Y(new_n15866_));
  OR4X1    g15802(.A(new_n276_), .B(new_n259_), .C(new_n228_), .D(new_n138_), .Y(new_n15867_));
  OR4X1    g15803(.A(new_n15867_), .B(new_n509_), .C(new_n395_), .D(new_n483_), .Y(new_n15868_));
  OR4X1    g15804(.A(new_n15868_), .B(new_n614_), .C(new_n389_), .D(new_n189_), .Y(new_n15869_));
  OR4X1    g15805(.A(new_n15869_), .B(new_n15866_), .C(new_n8313_), .D(new_n2227_), .Y(new_n15870_));
  NOR3X1   g15806(.A(new_n15870_), .B(new_n1476_), .C(new_n727_), .Y(new_n15871_));
  XOR2X1   g15807(.A(new_n15871_), .B(new_n15709_), .Y(new_n15872_));
  OR2X1    g15808(.A(new_n15872_), .B(new_n15865_), .Y(new_n15873_));
  OR2X1    g15809(.A(new_n15871_), .B(new_n15709_), .Y(new_n15874_));
  NAND3X1  g15810(.A(new_n15871_), .B(new_n15526_), .C(new_n15525_), .Y(new_n15875_));
  NAND3X1  g15811(.A(new_n15875_), .B(new_n15874_), .C(new_n15865_), .Y(new_n15876_));
  NAND2X1  g15812(.A(new_n15876_), .B(new_n15873_), .Y(new_n15877_));
  OR2X1    g15813(.A(new_n12685_), .B(new_n3178_), .Y(new_n15878_));
  OAI22X1  g15814(.A0(new_n12117_), .A1(new_n2245_), .B0(new_n12113_), .B1(new_n1885_), .Y(new_n15879_));
  AOI21X1  g15815(.A0(new_n12208_), .A1(new_n1889_), .B0(new_n15879_), .Y(new_n15880_));
  AND2X1   g15816(.A(new_n15880_), .B(new_n15878_), .Y(new_n15881_));
  XOR2X1   g15817(.A(new_n15881_), .B(new_n15877_), .Y(new_n15882_));
  AOI21X1  g15818(.A0(new_n15718_), .A1(new_n15716_), .B0(new_n15714_), .Y(new_n15883_));
  NOR2X1   g15819(.A(new_n15733_), .B(new_n15883_), .Y(new_n15884_));
  XOR2X1   g15820(.A(new_n15884_), .B(new_n15882_), .Y(new_n15885_));
  AOI22X1  g15821(.A0(new_n12107_), .A1(new_n2185_), .B0(new_n12104_), .B1(new_n2095_), .Y(new_n15886_));
  OAI21X1  g15822(.A0(new_n12306_), .A1(new_n2140_), .B0(new_n15886_), .Y(new_n15887_));
  AOI21X1  g15823(.A0(new_n12305_), .A1(new_n2062_), .B0(new_n15887_), .Y(new_n15888_));
  XOR2X1   g15824(.A(new_n15888_), .B(\a[29] ), .Y(new_n15889_));
  XOR2X1   g15825(.A(new_n15889_), .B(new_n15885_), .Y(new_n15890_));
  AOI22X1  g15826(.A0(new_n12099_), .A1(new_n2424_), .B0(new_n12097_), .B1(new_n2418_), .Y(new_n15891_));
  OAI21X1  g15827(.A0(new_n13090_), .A1(new_n2626_), .B0(new_n15891_), .Y(new_n15892_));
  AOI21X1  g15828(.A0(new_n14519_), .A1(new_n2301_), .B0(new_n15892_), .Y(new_n15893_));
  XOR2X1   g15829(.A(new_n15893_), .B(\a[26] ), .Y(new_n15894_));
  XOR2X1   g15830(.A(new_n15894_), .B(new_n15890_), .Y(new_n15895_));
  NAND3X1  g15831(.A(new_n15734_), .B(new_n15726_), .C(new_n15722_), .Y(new_n15896_));
  OAI21X1  g15832(.A0(new_n15743_), .A1(new_n15742_), .B0(new_n15740_), .Y(new_n15897_));
  AND2X1   g15833(.A(new_n15897_), .B(new_n15896_), .Y(new_n15898_));
  XOR2X1   g15834(.A(new_n15898_), .B(new_n15895_), .Y(new_n15899_));
  AOI22X1  g15835(.A0(new_n12093_), .A1(new_n2657_), .B0(new_n12090_), .B1(new_n2696_), .Y(new_n15900_));
  OAI21X1  g15836(.A0(new_n13104_), .A1(new_n2753_), .B0(new_n15900_), .Y(new_n15901_));
  AOI21X1  g15837(.A0(new_n13103_), .A1(new_n2658_), .B0(new_n15901_), .Y(new_n15902_));
  XOR2X1   g15838(.A(new_n15902_), .B(\a[23] ), .Y(new_n15903_));
  XOR2X1   g15839(.A(new_n15903_), .B(new_n15899_), .Y(new_n15904_));
  AOI21X1  g15840(.A0(new_n15755_), .A1(new_n15757_), .B0(new_n15750_), .Y(new_n15905_));
  XOR2X1   g15841(.A(new_n15905_), .B(new_n15904_), .Y(new_n15906_));
  AOI22X1  g15842(.A0(new_n12085_), .A1(new_n2875_), .B0(new_n12083_), .B1(new_n3099_), .Y(new_n15907_));
  OAI21X1  g15843(.A0(new_n13320_), .A1(new_n3152_), .B0(new_n15907_), .Y(new_n15908_));
  AOI21X1  g15844(.A0(new_n14510_), .A1(new_n2876_), .B0(new_n15908_), .Y(new_n15909_));
  XOR2X1   g15845(.A(new_n15909_), .B(\a[20] ), .Y(new_n15910_));
  XOR2X1   g15846(.A(new_n15910_), .B(new_n15906_), .Y(new_n15911_));
  AOI21X1  g15847(.A0(new_n15770_), .A1(new_n15772_), .B0(new_n15765_), .Y(new_n15912_));
  XOR2X1   g15848(.A(new_n15912_), .B(new_n15911_), .Y(new_n15913_));
  AOI22X1  g15849(.A0(new_n12079_), .A1(new_n3232_), .B0(new_n12076_), .B1(new_n3390_), .Y(new_n15914_));
  OAI21X1  g15850(.A0(new_n13691_), .A1(new_n3545_), .B0(new_n15914_), .Y(new_n15915_));
  AOI21X1  g15851(.A0(new_n13690_), .A1(new_n3234_), .B0(new_n15915_), .Y(new_n15916_));
  XOR2X1   g15852(.A(new_n15916_), .B(\a[17] ), .Y(new_n15917_));
  XOR2X1   g15853(.A(new_n15917_), .B(new_n15913_), .Y(new_n15918_));
  AOI21X1  g15854(.A0(new_n15785_), .A1(new_n15787_), .B0(new_n15780_), .Y(new_n15919_));
  XOR2X1   g15855(.A(new_n15919_), .B(new_n15918_), .Y(new_n15920_));
  AOI22X1  g15856(.A0(new_n12285_), .A1(new_n3908_), .B0(new_n12074_), .B1(new_n3628_), .Y(new_n15921_));
  OAI21X1  g15857(.A0(new_n14086_), .A1(new_n3983_), .B0(new_n15921_), .Y(new_n15922_));
  AOI21X1  g15858(.A0(new_n14480_), .A1(new_n3624_), .B0(new_n15922_), .Y(new_n15923_));
  XOR2X1   g15859(.A(new_n15923_), .B(\a[14] ), .Y(new_n15924_));
  XOR2X1   g15860(.A(new_n15924_), .B(new_n15920_), .Y(new_n15925_));
  AOI21X1  g15861(.A0(new_n15800_), .A1(new_n15802_), .B0(new_n15795_), .Y(new_n15926_));
  XOR2X1   g15862(.A(new_n15926_), .B(new_n15925_), .Y(new_n15927_));
  AOI22X1  g15863(.A0(new_n14087_), .A1(new_n4078_), .B0(new_n14084_), .B1(new_n4247_), .Y(new_n15928_));
  OAI21X1  g15864(.A0(new_n14648_), .A1(new_n4427_), .B0(new_n15928_), .Y(new_n15929_));
  AOI21X1  g15865(.A0(new_n14651_), .A1(new_n4080_), .B0(new_n15929_), .Y(new_n15930_));
  XOR2X1   g15866(.A(new_n15930_), .B(\a[11] ), .Y(new_n15931_));
  XOR2X1   g15867(.A(new_n15931_), .B(new_n15927_), .Y(new_n15932_));
  AOI21X1  g15868(.A0(new_n15815_), .A1(new_n15817_), .B0(new_n15810_), .Y(new_n15933_));
  XOR2X1   g15869(.A(new_n15933_), .B(new_n15932_), .Y(new_n15934_));
  AOI22X1  g15870(.A0(new_n14946_), .A1(new_n4870_), .B0(new_n14804_), .B1(new_n4635_), .Y(new_n15935_));
  OAI21X1  g15871(.A0(new_n15235_), .A1(new_n5096_), .B0(new_n15935_), .Y(new_n15936_));
  AOI21X1  g15872(.A0(new_n15381_), .A1(new_n4637_), .B0(new_n15936_), .Y(new_n15937_));
  XOR2X1   g15873(.A(new_n15937_), .B(\a[8] ), .Y(new_n15938_));
  XOR2X1   g15874(.A(new_n15938_), .B(new_n15934_), .Y(new_n15939_));
  AOI21X1  g15875(.A0(new_n15830_), .A1(new_n15832_), .B0(new_n15825_), .Y(new_n15940_));
  AOI22X1  g15876(.A0(new_n15362_), .A1(new_n10534_), .B0(new_n15234_), .B1(new_n5373_), .Y(new_n15941_));
  OAI21X1  g15877(.A0(new_n15373_), .A1(new_n5657_), .B0(new_n15941_), .Y(new_n15942_));
  XOR2X1   g15878(.A(new_n15942_), .B(new_n3289_), .Y(new_n15943_));
  XOR2X1   g15879(.A(new_n15943_), .B(new_n15940_), .Y(new_n15944_));
  XOR2X1   g15880(.A(new_n15944_), .B(new_n15939_), .Y(new_n15945_));
  AOI21X1  g15881(.A0(new_n15846_), .A1(new_n15848_), .B0(new_n15840_), .Y(new_n15946_));
  XOR2X1   g15882(.A(new_n15946_), .B(new_n15945_), .Y(new_n15947_));
  NAND3X1  g15883(.A(new_n15855_), .B(new_n15854_), .C(new_n15853_), .Y(new_n15948_));
  NOR3X1   g15884(.A(new_n15683_), .B(new_n15682_), .C(new_n15681_), .Y(new_n15949_));
  OAI21X1  g15885(.A0(new_n15689_), .A1(new_n15949_), .B0(new_n15684_), .Y(new_n15950_));
  AOI21X1  g15886(.A0(new_n15950_), .A1(new_n15948_), .B0(new_n15856_), .Y(new_n15951_));
  XOR2X1   g15887(.A(new_n15951_), .B(new_n15947_), .Y(new_n15952_));
  INVX1    g15888(.A(new_n15952_), .Y(new_n15953_));
  XOR2X1   g15889(.A(new_n15953_), .B(new_n15863_), .Y(\result[9] ));
  NOR2X1   g15890(.A(new_n15953_), .B(new_n15863_), .Y(new_n15955_));
  AND2X1   g15891(.A(new_n15876_), .B(new_n15873_), .Y(new_n15956_));
  XOR2X1   g15892(.A(new_n15881_), .B(new_n15956_), .Y(new_n15957_));
  XOR2X1   g15893(.A(new_n15884_), .B(new_n15957_), .Y(new_n15958_));
  XOR2X1   g15894(.A(new_n15889_), .B(new_n15958_), .Y(new_n15959_));
  XOR2X1   g15895(.A(new_n15894_), .B(new_n15959_), .Y(new_n15960_));
  XOR2X1   g15896(.A(new_n15898_), .B(new_n15960_), .Y(new_n15961_));
  XOR2X1   g15897(.A(new_n15903_), .B(new_n15961_), .Y(new_n15962_));
  XOR2X1   g15898(.A(new_n15905_), .B(new_n15962_), .Y(new_n15963_));
  XOR2X1   g15899(.A(new_n15910_), .B(new_n15963_), .Y(new_n15964_));
  XOR2X1   g15900(.A(new_n15912_), .B(new_n15964_), .Y(new_n15965_));
  XOR2X1   g15901(.A(new_n15917_), .B(new_n15965_), .Y(new_n15966_));
  XOR2X1   g15902(.A(new_n15919_), .B(new_n15966_), .Y(new_n15967_));
  XOR2X1   g15903(.A(new_n15924_), .B(new_n15967_), .Y(new_n15968_));
  XOR2X1   g15904(.A(new_n15926_), .B(new_n15968_), .Y(new_n15969_));
  XOR2X1   g15905(.A(new_n15931_), .B(new_n15969_), .Y(new_n15970_));
  XOR2X1   g15906(.A(new_n15933_), .B(new_n15970_), .Y(new_n15971_));
  XOR2X1   g15907(.A(new_n15938_), .B(new_n15971_), .Y(new_n15972_));
  XOR2X1   g15908(.A(new_n15944_), .B(new_n15972_), .Y(new_n15973_));
  OR2X1    g15909(.A(new_n15946_), .B(new_n15973_), .Y(new_n15974_));
  OAI21X1  g15910(.A0(new_n15951_), .A1(new_n15947_), .B0(new_n15974_), .Y(new_n15975_));
  NAND2X1  g15911(.A(new_n15944_), .B(new_n15939_), .Y(new_n15976_));
  OAI21X1  g15912(.A0(new_n15943_), .A1(new_n15940_), .B0(new_n15976_), .Y(new_n15977_));
  OR2X1    g15913(.A(new_n15881_), .B(new_n15956_), .Y(new_n15978_));
  OAI21X1  g15914(.A0(new_n15884_), .A1(new_n15882_), .B0(new_n15978_), .Y(new_n15979_));
  INVX1    g15915(.A(new_n15875_), .Y(new_n15980_));
  OAI21X1  g15916(.A0(new_n15980_), .A1(new_n15865_), .B0(new_n15874_), .Y(new_n15981_));
  NOR4X1   g15917(.A(new_n740_), .B(new_n396_), .C(new_n276_), .D(new_n193_), .Y(new_n15982_));
  NOR4X1   g15918(.A(new_n1608_), .B(new_n935_), .C(new_n1183_), .D(new_n572_), .Y(new_n15983_));
  OR4X1    g15919(.A(new_n2580_), .B(new_n3434_), .C(new_n2302_), .D(new_n1646_), .Y(new_n15984_));
  NOR4X1   g15920(.A(new_n15984_), .B(new_n7457_), .C(new_n1105_), .D(new_n561_), .Y(new_n15985_));
  NAND3X1  g15921(.A(new_n15985_), .B(new_n15983_), .C(new_n15982_), .Y(new_n15986_));
  NOR4X1   g15922(.A(new_n15986_), .B(new_n12405_), .C(new_n1918_), .D(new_n1310_), .Y(new_n15987_));
  XOR2X1   g15923(.A(new_n15987_), .B(new_n15709_), .Y(new_n15988_));
  AND2X1   g15924(.A(new_n15362_), .B(new_n8194_), .Y(new_n15989_));
  XOR2X1   g15925(.A(new_n15989_), .B(new_n3289_), .Y(new_n15990_));
  XOR2X1   g15926(.A(new_n15990_), .B(new_n15988_), .Y(new_n15991_));
  XOR2X1   g15927(.A(new_n15991_), .B(new_n15981_), .Y(new_n15992_));
  OR2X1    g15928(.A(new_n12708_), .B(new_n3178_), .Y(new_n15993_));
  OAI22X1  g15929(.A0(new_n12113_), .A1(new_n2245_), .B0(new_n12111_), .B1(new_n1885_), .Y(new_n15994_));
  AOI21X1  g15930(.A0(new_n12107_), .A1(new_n1889_), .B0(new_n15994_), .Y(new_n15995_));
  AND2X1   g15931(.A(new_n15995_), .B(new_n15993_), .Y(new_n15996_));
  XOR2X1   g15932(.A(new_n15996_), .B(new_n15992_), .Y(new_n15997_));
  XOR2X1   g15933(.A(new_n15997_), .B(new_n15979_), .Y(new_n15998_));
  AOI22X1  g15934(.A0(new_n12104_), .A1(new_n2185_), .B0(new_n12102_), .B1(new_n2095_), .Y(new_n15999_));
  OAI21X1  g15935(.A0(new_n12840_), .A1(new_n2140_), .B0(new_n15999_), .Y(new_n16000_));
  AOI21X1  g15936(.A0(new_n12859_), .A1(new_n2062_), .B0(new_n16000_), .Y(new_n16001_));
  XOR2X1   g15937(.A(new_n16001_), .B(\a[29] ), .Y(new_n16002_));
  XOR2X1   g15938(.A(new_n16002_), .B(new_n15998_), .Y(new_n16003_));
  AOI22X1  g15939(.A0(new_n12097_), .A1(new_n2424_), .B0(new_n12095_), .B1(new_n2418_), .Y(new_n16004_));
  OAI21X1  g15940(.A0(new_n13366_), .A1(new_n2626_), .B0(new_n16004_), .Y(new_n16005_));
  AOI21X1  g15941(.A0(new_n13093_), .A1(new_n2301_), .B0(new_n16005_), .Y(new_n16006_));
  XOR2X1   g15942(.A(new_n16006_), .B(\a[26] ), .Y(new_n16007_));
  XOR2X1   g15943(.A(new_n16007_), .B(new_n16003_), .Y(new_n16008_));
  OR2X1    g15944(.A(new_n15889_), .B(new_n15958_), .Y(new_n16009_));
  OR2X1    g15945(.A(new_n15894_), .B(new_n15890_), .Y(new_n16010_));
  AND2X1   g15946(.A(new_n16010_), .B(new_n16009_), .Y(new_n16011_));
  XOR2X1   g15947(.A(new_n16011_), .B(new_n16008_), .Y(new_n16012_));
  AOI22X1  g15948(.A0(new_n12090_), .A1(new_n2657_), .B0(new_n12088_), .B1(new_n2696_), .Y(new_n16013_));
  OAI21X1  g15949(.A0(new_n12298_), .A1(new_n2753_), .B0(new_n16013_), .Y(new_n16014_));
  AOI21X1  g15950(.A0(new_n12297_), .A1(new_n2658_), .B0(new_n16014_), .Y(new_n16015_));
  XOR2X1   g15951(.A(new_n16015_), .B(\a[23] ), .Y(new_n16016_));
  XOR2X1   g15952(.A(new_n16016_), .B(new_n16012_), .Y(new_n16017_));
  OR2X1    g15953(.A(new_n15898_), .B(new_n15960_), .Y(new_n16018_));
  OAI21X1  g15954(.A0(new_n15903_), .A1(new_n15899_), .B0(new_n16018_), .Y(new_n16019_));
  XOR2X1   g15955(.A(new_n16019_), .B(new_n16017_), .Y(new_n16020_));
  AOI22X1  g15956(.A0(new_n12083_), .A1(new_n2875_), .B0(new_n12081_), .B1(new_n3099_), .Y(new_n16021_));
  OAI21X1  g15957(.A0(new_n13665_), .A1(new_n3152_), .B0(new_n16021_), .Y(new_n16022_));
  AOI21X1  g15958(.A0(new_n14672_), .A1(new_n2876_), .B0(new_n16022_), .Y(new_n16023_));
  XOR2X1   g15959(.A(new_n16023_), .B(\a[20] ), .Y(new_n16024_));
  XOR2X1   g15960(.A(new_n16024_), .B(new_n16020_), .Y(new_n16025_));
  OR2X1    g15961(.A(new_n15905_), .B(new_n15962_), .Y(new_n16026_));
  OAI21X1  g15962(.A0(new_n15910_), .A1(new_n15906_), .B0(new_n16026_), .Y(new_n16027_));
  XOR2X1   g15963(.A(new_n16027_), .B(new_n16025_), .Y(new_n16028_));
  AOI22X1  g15964(.A0(new_n12076_), .A1(new_n3232_), .B0(new_n12018_), .B1(new_n3390_), .Y(new_n16029_));
  OAI21X1  g15965(.A0(new_n13679_), .A1(new_n3545_), .B0(new_n16029_), .Y(new_n16030_));
  AOI21X1  g15966(.A0(new_n13678_), .A1(new_n3234_), .B0(new_n16030_), .Y(new_n16031_));
  XOR2X1   g15967(.A(new_n16031_), .B(\a[17] ), .Y(new_n16032_));
  INVX1    g15968(.A(new_n16032_), .Y(new_n16033_));
  XOR2X1   g15969(.A(new_n16033_), .B(new_n16028_), .Y(new_n16034_));
  NOR2X1   g15970(.A(new_n15912_), .B(new_n15964_), .Y(new_n16035_));
  XOR2X1   g15971(.A(new_n15916_), .B(new_n2445_), .Y(new_n16036_));
  AOI21X1  g15972(.A0(new_n16036_), .A1(new_n15965_), .B0(new_n16035_), .Y(new_n16037_));
  XOR2X1   g15973(.A(new_n16037_), .B(new_n16034_), .Y(new_n16038_));
  OR2X1    g15974(.A(new_n15919_), .B(new_n15966_), .Y(new_n16039_));
  OAI21X1  g15975(.A0(new_n15924_), .A1(new_n15920_), .B0(new_n16039_), .Y(new_n16040_));
  AOI22X1  g15976(.A0(new_n14085_), .A1(new_n3908_), .B0(new_n12285_), .B1(new_n3628_), .Y(new_n16041_));
  OAI21X1  g15977(.A0(new_n14088_), .A1(new_n3983_), .B0(new_n16041_), .Y(new_n16042_));
  AOI21X1  g15978(.A0(new_n14491_), .A1(new_n3624_), .B0(new_n16042_), .Y(new_n16043_));
  XOR2X1   g15979(.A(new_n16043_), .B(\a[14] ), .Y(new_n16044_));
  INVX1    g15980(.A(new_n16044_), .Y(new_n16045_));
  XOR2X1   g15981(.A(new_n16045_), .B(new_n16040_), .Y(new_n16046_));
  XOR2X1   g15982(.A(new_n16046_), .B(new_n16038_), .Y(new_n16047_));
  AOI22X1  g15983(.A0(new_n14642_), .A1(new_n4247_), .B0(new_n14084_), .B1(new_n4078_), .Y(new_n16048_));
  OAI21X1  g15984(.A0(new_n14805_), .A1(new_n4427_), .B0(new_n16048_), .Y(new_n16049_));
  AOI21X1  g15985(.A0(new_n14809_), .A1(new_n4080_), .B0(new_n16049_), .Y(new_n16050_));
  XOR2X1   g15986(.A(new_n16050_), .B(\a[11] ), .Y(new_n16051_));
  INVX1    g15987(.A(new_n16051_), .Y(new_n16052_));
  XOR2X1   g15988(.A(new_n16052_), .B(new_n16047_), .Y(new_n16053_));
  OR2X1    g15989(.A(new_n15926_), .B(new_n15968_), .Y(new_n16054_));
  OAI21X1  g15990(.A0(new_n15931_), .A1(new_n15927_), .B0(new_n16054_), .Y(new_n16055_));
  XOR2X1   g15991(.A(new_n16055_), .B(new_n16053_), .Y(new_n16056_));
  OR2X1    g15992(.A(new_n15933_), .B(new_n15970_), .Y(new_n16057_));
  OAI21X1  g15993(.A0(new_n15938_), .A1(new_n15934_), .B0(new_n16057_), .Y(new_n16058_));
  AOI22X1  g15994(.A0(new_n15087_), .A1(new_n4870_), .B0(new_n14946_), .B1(new_n4635_), .Y(new_n16059_));
  OAI21X1  g15995(.A0(new_n15363_), .A1(new_n5096_), .B0(new_n16059_), .Y(new_n16060_));
  AOI21X1  g15996(.A0(new_n15240_), .A1(new_n4637_), .B0(new_n16060_), .Y(new_n16061_));
  XOR2X1   g15997(.A(new_n16061_), .B(new_n2995_), .Y(new_n16062_));
  XOR2X1   g15998(.A(new_n16062_), .B(new_n16058_), .Y(new_n16063_));
  XOR2X1   g15999(.A(new_n16063_), .B(new_n16056_), .Y(new_n16064_));
  XOR2X1   g16000(.A(new_n16064_), .B(new_n15977_), .Y(new_n16065_));
  XOR2X1   g16001(.A(new_n16065_), .B(new_n15975_), .Y(new_n16066_));
  XOR2X1   g16002(.A(new_n16066_), .B(new_n15955_), .Y(\result[10] ));
  NAND4X1  g16003(.A(new_n16066_), .B(new_n15952_), .C(new_n15861_), .D(new_n15692_), .Y(new_n16068_));
  AND2X1   g16004(.A(new_n15997_), .B(new_n15979_), .Y(new_n16069_));
  INVX1    g16005(.A(new_n16002_), .Y(new_n16070_));
  AOI21X1  g16006(.A0(new_n16070_), .A1(new_n15998_), .B0(new_n16069_), .Y(new_n16071_));
  AOI22X1  g16007(.A0(new_n12208_), .A1(new_n1890_), .B0(new_n12107_), .B1(new_n1884_), .Y(new_n16072_));
  OAI21X1  g16008(.A0(new_n12695_), .A1(new_n3498_), .B0(new_n16072_), .Y(new_n16073_));
  AOI21X1  g16009(.A0(new_n12694_), .A1(new_n407_), .B0(new_n16073_), .Y(new_n16074_));
  OR4X1    g16010(.A(new_n3445_), .B(new_n1062_), .C(new_n1021_), .D(new_n947_), .Y(new_n16075_));
  OR4X1    g16011(.A(new_n1261_), .B(new_n273_), .C(new_n399_), .D(new_n100_), .Y(new_n16076_));
  OR4X1    g16012(.A(new_n16076_), .B(new_n980_), .C(new_n830_), .D(new_n629_), .Y(new_n16077_));
  OR4X1    g16013(.A(new_n16077_), .B(new_n16075_), .C(new_n3784_), .D(new_n2165_), .Y(new_n16078_));
  OR4X1    g16014(.A(new_n3283_), .B(new_n1850_), .C(new_n1269_), .D(new_n1136_), .Y(new_n16079_));
  OR4X1    g16015(.A(new_n16079_), .B(new_n3808_), .C(new_n665_), .D(new_n663_), .Y(new_n16080_));
  OR4X1    g16016(.A(new_n414_), .B(new_n393_), .C(new_n259_), .D(new_n1008_), .Y(new_n16081_));
  OR4X1    g16017(.A(new_n1732_), .B(new_n1082_), .C(new_n504_), .D(new_n579_), .Y(new_n16082_));
  OR4X1    g16018(.A(new_n16082_), .B(new_n16081_), .C(new_n857_), .D(new_n311_), .Y(new_n16083_));
  OR4X1    g16019(.A(new_n16083_), .B(new_n1117_), .C(new_n1115_), .D(new_n1114_), .Y(new_n16084_));
  NOR4X1   g16020(.A(new_n16084_), .B(new_n16080_), .C(new_n16078_), .D(new_n564_), .Y(new_n16085_));
  INVX1    g16021(.A(new_n15988_), .Y(new_n16086_));
  NOR3X1   g16022(.A(new_n15987_), .B(new_n15523_), .C(new_n15520_), .Y(new_n16087_));
  AOI21X1  g16023(.A0(new_n15990_), .A1(new_n16086_), .B0(new_n16087_), .Y(new_n16088_));
  XOR2X1   g16024(.A(new_n16088_), .B(new_n16085_), .Y(new_n16089_));
  XOR2X1   g16025(.A(new_n16089_), .B(new_n16074_), .Y(new_n16090_));
  NOR2X1   g16026(.A(new_n15996_), .B(new_n15992_), .Y(new_n16091_));
  INVX1    g16027(.A(new_n15991_), .Y(new_n16092_));
  AND2X1   g16028(.A(new_n16092_), .B(new_n15981_), .Y(new_n16093_));
  NOR2X1   g16029(.A(new_n16093_), .B(new_n16091_), .Y(new_n16094_));
  XOR2X1   g16030(.A(new_n16094_), .B(new_n16090_), .Y(new_n16095_));
  OAI22X1  g16031(.A0(new_n12306_), .A1(new_n2186_), .B0(new_n12840_), .B1(new_n2431_), .Y(new_n16096_));
  AOI21X1  g16032(.A0(new_n12097_), .A1(new_n2139_), .B0(new_n16096_), .Y(new_n16097_));
  OAI21X1  g16033(.A0(new_n12856_), .A1(new_n2063_), .B0(new_n16097_), .Y(new_n16098_));
  XOR2X1   g16034(.A(new_n16098_), .B(new_n74_), .Y(new_n16099_));
  XOR2X1   g16035(.A(new_n16099_), .B(new_n16095_), .Y(new_n16100_));
  XOR2X1   g16036(.A(new_n16100_), .B(new_n16071_), .Y(new_n16101_));
  AOI22X1  g16037(.A0(new_n12095_), .A1(new_n2424_), .B0(new_n12093_), .B1(new_n2418_), .Y(new_n16102_));
  OAI21X1  g16038(.A0(new_n13118_), .A1(new_n2626_), .B0(new_n16102_), .Y(new_n16103_));
  AOI21X1  g16039(.A0(new_n13117_), .A1(new_n2301_), .B0(new_n16103_), .Y(new_n16104_));
  XOR2X1   g16040(.A(new_n16104_), .B(\a[26] ), .Y(new_n16105_));
  INVX1    g16041(.A(new_n16105_), .Y(new_n16106_));
  XOR2X1   g16042(.A(new_n16106_), .B(new_n16101_), .Y(new_n16107_));
  NOR2X1   g16043(.A(new_n16007_), .B(new_n16003_), .Y(new_n16108_));
  OAI21X1  g16044(.A0(new_n15894_), .A1(new_n15890_), .B0(new_n16009_), .Y(new_n16109_));
  AOI21X1  g16045(.A0(new_n16109_), .A1(new_n16008_), .B0(new_n16108_), .Y(new_n16110_));
  XOR2X1   g16046(.A(new_n16110_), .B(new_n16107_), .Y(new_n16111_));
  AOI22X1  g16047(.A0(new_n12088_), .A1(new_n2657_), .B0(new_n12085_), .B1(new_n2696_), .Y(new_n16112_));
  OAI21X1  g16048(.A0(new_n13321_), .A1(new_n2753_), .B0(new_n16112_), .Y(new_n16113_));
  AOI21X1  g16049(.A0(new_n13344_), .A1(new_n2658_), .B0(new_n16113_), .Y(new_n16114_));
  XOR2X1   g16050(.A(new_n16114_), .B(\a[23] ), .Y(new_n16115_));
  XOR2X1   g16051(.A(new_n16115_), .B(new_n16111_), .Y(new_n16116_));
  NOR2X1   g16052(.A(new_n16016_), .B(new_n16012_), .Y(new_n16117_));
  AOI21X1  g16053(.A0(new_n16019_), .A1(new_n16017_), .B0(new_n16117_), .Y(new_n16118_));
  XOR2X1   g16054(.A(new_n16118_), .B(new_n16116_), .Y(new_n16119_));
  AOI22X1  g16055(.A0(new_n12081_), .A1(new_n2875_), .B0(new_n12079_), .B1(new_n3099_), .Y(new_n16120_));
  OAI21X1  g16056(.A0(new_n13700_), .A1(new_n3152_), .B0(new_n16120_), .Y(new_n16121_));
  AOI21X1  g16057(.A0(new_n13699_), .A1(new_n2876_), .B0(new_n16121_), .Y(new_n16122_));
  XOR2X1   g16058(.A(new_n16122_), .B(\a[20] ), .Y(new_n16123_));
  XOR2X1   g16059(.A(new_n16123_), .B(new_n16119_), .Y(new_n16124_));
  INVX1    g16060(.A(new_n16024_), .Y(new_n16125_));
  XOR2X1   g16061(.A(new_n16125_), .B(new_n16020_), .Y(new_n16126_));
  AND2X1   g16062(.A(new_n16027_), .B(new_n16126_), .Y(new_n16127_));
  AOI21X1  g16063(.A0(new_n16125_), .A1(new_n16020_), .B0(new_n16127_), .Y(new_n16128_));
  XOR2X1   g16064(.A(new_n16128_), .B(new_n16124_), .Y(new_n16129_));
  AOI22X1  g16065(.A0(new_n12074_), .A1(new_n3390_), .B0(new_n12018_), .B1(new_n3232_), .Y(new_n16130_));
  OAI21X1  g16066(.A0(new_n12292_), .A1(new_n3545_), .B0(new_n16130_), .Y(new_n16131_));
  AOI21X1  g16067(.A0(new_n12291_), .A1(new_n3234_), .B0(new_n16131_), .Y(new_n16132_));
  XOR2X1   g16068(.A(new_n16132_), .B(\a[17] ), .Y(new_n16133_));
  XOR2X1   g16069(.A(new_n16133_), .B(new_n16129_), .Y(new_n16134_));
  NOR2X1   g16070(.A(new_n16032_), .B(new_n16028_), .Y(new_n16135_));
  NOR2X1   g16071(.A(new_n16037_), .B(new_n16034_), .Y(new_n16136_));
  NOR2X1   g16072(.A(new_n16136_), .B(new_n16135_), .Y(new_n16137_));
  XOR2X1   g16073(.A(new_n16137_), .B(new_n16134_), .Y(new_n16138_));
  AOI22X1  g16074(.A0(new_n14087_), .A1(new_n3908_), .B0(new_n14085_), .B1(new_n3628_), .Y(new_n16139_));
  OAI21X1  g16075(.A0(new_n14643_), .A1(new_n3983_), .B0(new_n16139_), .Y(new_n16140_));
  AOI21X1  g16076(.A0(new_n14106_), .A1(new_n3624_), .B0(new_n16140_), .Y(new_n16141_));
  XOR2X1   g16077(.A(new_n16141_), .B(\a[14] ), .Y(new_n16142_));
  XOR2X1   g16078(.A(new_n16142_), .B(new_n16138_), .Y(new_n16143_));
  AND2X1   g16079(.A(new_n16045_), .B(new_n16040_), .Y(new_n16144_));
  AOI21X1  g16080(.A0(new_n16046_), .A1(new_n16038_), .B0(new_n16144_), .Y(new_n16145_));
  XOR2X1   g16081(.A(new_n16145_), .B(new_n16143_), .Y(new_n16146_));
  AOI22X1  g16082(.A0(new_n14804_), .A1(new_n4247_), .B0(new_n14642_), .B1(new_n4078_), .Y(new_n16147_));
  OAI21X1  g16083(.A0(new_n15088_), .A1(new_n4427_), .B0(new_n16147_), .Y(new_n16148_));
  AOI21X1  g16084(.A0(new_n14952_), .A1(new_n4080_), .B0(new_n16148_), .Y(new_n16149_));
  XOR2X1   g16085(.A(new_n16149_), .B(\a[11] ), .Y(new_n16150_));
  XOR2X1   g16086(.A(new_n16150_), .B(new_n16146_), .Y(new_n16151_));
  AND2X1   g16087(.A(new_n16052_), .B(new_n16047_), .Y(new_n16152_));
  AOI21X1  g16088(.A0(new_n16055_), .A1(new_n16053_), .B0(new_n16152_), .Y(new_n16153_));
  XOR2X1   g16089(.A(new_n16153_), .B(new_n16151_), .Y(new_n16154_));
  AOI22X1  g16090(.A0(new_n15234_), .A1(new_n4870_), .B0(new_n15087_), .B1(new_n4635_), .Y(new_n16155_));
  OAI21X1  g16091(.A0(new_n15522_), .A1(new_n5096_), .B0(new_n16155_), .Y(new_n16156_));
  AOI21X1  g16092(.A0(new_n15841_), .A1(new_n4637_), .B0(new_n16156_), .Y(new_n16157_));
  XOR2X1   g16093(.A(new_n16157_), .B(\a[8] ), .Y(new_n16158_));
  XOR2X1   g16094(.A(new_n16158_), .B(new_n16154_), .Y(new_n16159_));
  AND2X1   g16095(.A(new_n16062_), .B(new_n16058_), .Y(new_n16160_));
  AOI21X1  g16096(.A0(new_n16063_), .A1(new_n16056_), .B0(new_n16160_), .Y(new_n16161_));
  XOR2X1   g16097(.A(new_n16161_), .B(new_n16159_), .Y(new_n16162_));
  AND2X1   g16098(.A(new_n16064_), .B(new_n15977_), .Y(new_n16163_));
  AOI21X1  g16099(.A0(new_n16065_), .A1(new_n15975_), .B0(new_n16163_), .Y(new_n16164_));
  XOR2X1   g16100(.A(new_n16164_), .B(new_n16162_), .Y(new_n16165_));
  XOR2X1   g16101(.A(new_n16165_), .B(new_n16068_), .Y(\result[11] ));
  NOR2X1   g16102(.A(new_n16165_), .B(new_n16068_), .Y(new_n16167_));
  INVX1    g16103(.A(new_n16085_), .Y(new_n16168_));
  NOR2X1   g16104(.A(new_n16088_), .B(new_n16168_), .Y(new_n16169_));
  NOR2X1   g16105(.A(new_n16089_), .B(new_n16074_), .Y(new_n16170_));
  OR2X1    g16106(.A(new_n16170_), .B(new_n16169_), .Y(new_n16171_));
  NAND3X1  g16107(.A(new_n8566_), .B(new_n1940_), .C(new_n2161_), .Y(new_n16172_));
  OR4X1    g16108(.A(new_n247_), .B(new_n757_), .C(new_n825_), .D(new_n111_), .Y(new_n16173_));
  OR4X1    g16109(.A(new_n16173_), .B(new_n16172_), .C(new_n7022_), .D(new_n216_), .Y(new_n16174_));
  OR4X1    g16110(.A(new_n786_), .B(new_n301_), .C(new_n1613_), .D(new_n200_), .Y(new_n16175_));
  OR4X1    g16111(.A(new_n16175_), .B(new_n16174_), .C(new_n1590_), .D(new_n824_), .Y(new_n16176_));
  OAI22X1  g16112(.A0(new_n152_), .A1(new_n108_), .B0(new_n129_), .B1(new_n115_), .Y(new_n16177_));
  OR2X1    g16113(.A(new_n16177_), .B(new_n642_), .Y(new_n16178_));
  OR4X1    g16114(.A(new_n414_), .B(new_n483_), .C(new_n175_), .D(new_n664_), .Y(new_n16179_));
  OR4X1    g16115(.A(new_n16179_), .B(new_n16178_), .C(new_n616_), .D(new_n390_), .Y(new_n16180_));
  NOR3X1   g16116(.A(new_n2640_), .B(new_n459_), .C(new_n429_), .Y(new_n16181_));
  NOR4X1   g16117(.A(new_n348_), .B(new_n219_), .C(new_n141_), .D(new_n116_), .Y(new_n16182_));
  NOR4X1   g16118(.A(new_n3713_), .B(new_n497_), .C(new_n255_), .D(new_n254_), .Y(new_n16183_));
  NAND3X1  g16119(.A(new_n16183_), .B(new_n16182_), .C(new_n16181_), .Y(new_n16184_));
  OR4X1    g16120(.A(new_n16184_), .B(new_n16180_), .C(new_n6772_), .D(new_n1897_), .Y(new_n16185_));
  OR4X1    g16121(.A(new_n16185_), .B(new_n16176_), .C(new_n7449_), .D(new_n2947_), .Y(new_n16186_));
  XOR2X1   g16122(.A(new_n16186_), .B(new_n16085_), .Y(new_n16187_));
  INVX1    g16123(.A(new_n16187_), .Y(new_n16188_));
  NOR2X1   g16124(.A(new_n16186_), .B(new_n16085_), .Y(new_n16189_));
  AND2X1   g16125(.A(new_n16186_), .B(new_n16085_), .Y(new_n16190_));
  NOR4X1   g16126(.A(new_n16190_), .B(new_n16189_), .C(new_n16170_), .D(new_n16169_), .Y(new_n16191_));
  AOI21X1  g16127(.A0(new_n16188_), .A1(new_n16171_), .B0(new_n16191_), .Y(new_n16192_));
  AOI22X1  g16128(.A0(new_n12107_), .A1(new_n1890_), .B0(new_n12104_), .B1(new_n1884_), .Y(new_n16193_));
  OAI21X1  g16129(.A0(new_n12306_), .A1(new_n3498_), .B0(new_n16193_), .Y(new_n16194_));
  AOI21X1  g16130(.A0(new_n12305_), .A1(new_n407_), .B0(new_n16194_), .Y(new_n16195_));
  XOR2X1   g16131(.A(new_n16195_), .B(new_n16192_), .Y(new_n16196_));
  OAI21X1  g16132(.A0(new_n16093_), .A1(new_n16091_), .B0(new_n16090_), .Y(new_n16197_));
  OAI21X1  g16133(.A0(new_n16099_), .A1(new_n16095_), .B0(new_n16197_), .Y(new_n16198_));
  XOR2X1   g16134(.A(new_n16198_), .B(new_n16196_), .Y(new_n16199_));
  AOI22X1  g16135(.A0(new_n12099_), .A1(new_n2185_), .B0(new_n12097_), .B1(new_n2095_), .Y(new_n16200_));
  OAI21X1  g16136(.A0(new_n13090_), .A1(new_n2140_), .B0(new_n16200_), .Y(new_n16201_));
  AOI21X1  g16137(.A0(new_n14519_), .A1(new_n2062_), .B0(new_n16201_), .Y(new_n16202_));
  XOR2X1   g16138(.A(new_n16202_), .B(\a[29] ), .Y(new_n16203_));
  XOR2X1   g16139(.A(new_n16203_), .B(new_n16199_), .Y(new_n16204_));
  AOI22X1  g16140(.A0(new_n12093_), .A1(new_n2424_), .B0(new_n12090_), .B1(new_n2418_), .Y(new_n16205_));
  OAI21X1  g16141(.A0(new_n13104_), .A1(new_n2626_), .B0(new_n16205_), .Y(new_n16206_));
  AOI21X1  g16142(.A0(new_n13103_), .A1(new_n2301_), .B0(new_n16206_), .Y(new_n16207_));
  XOR2X1   g16143(.A(new_n16207_), .B(\a[26] ), .Y(new_n16208_));
  INVX1    g16144(.A(new_n16208_), .Y(new_n16209_));
  XOR2X1   g16145(.A(new_n16209_), .B(new_n16204_), .Y(new_n16210_));
  AND2X1   g16146(.A(new_n16070_), .B(new_n15998_), .Y(new_n16211_));
  OAI21X1  g16147(.A0(new_n16211_), .A1(new_n16069_), .B0(new_n16100_), .Y(new_n16212_));
  OR2X1    g16148(.A(new_n16105_), .B(new_n16101_), .Y(new_n16213_));
  AND2X1   g16149(.A(new_n16213_), .B(new_n16212_), .Y(new_n16214_));
  XOR2X1   g16150(.A(new_n16214_), .B(new_n16210_), .Y(new_n16215_));
  AOI22X1  g16151(.A0(new_n12085_), .A1(new_n2657_), .B0(new_n12083_), .B1(new_n2696_), .Y(new_n16216_));
  OAI21X1  g16152(.A0(new_n13320_), .A1(new_n2753_), .B0(new_n16216_), .Y(new_n16217_));
  AOI21X1  g16153(.A0(new_n14510_), .A1(new_n2658_), .B0(new_n16217_), .Y(new_n16218_));
  XOR2X1   g16154(.A(new_n16218_), .B(\a[23] ), .Y(new_n16219_));
  XOR2X1   g16155(.A(new_n16219_), .B(new_n16215_), .Y(new_n16220_));
  NOR2X1   g16156(.A(new_n16110_), .B(new_n16107_), .Y(new_n16221_));
  INVX1    g16157(.A(new_n16115_), .Y(new_n16222_));
  AOI21X1  g16158(.A0(new_n16222_), .A1(new_n16111_), .B0(new_n16221_), .Y(new_n16223_));
  XOR2X1   g16159(.A(new_n16223_), .B(new_n16220_), .Y(new_n16224_));
  AOI22X1  g16160(.A0(new_n12079_), .A1(new_n2875_), .B0(new_n12076_), .B1(new_n3099_), .Y(new_n16225_));
  OAI21X1  g16161(.A0(new_n13691_), .A1(new_n3152_), .B0(new_n16225_), .Y(new_n16226_));
  AOI21X1  g16162(.A0(new_n13690_), .A1(new_n2876_), .B0(new_n16226_), .Y(new_n16227_));
  XOR2X1   g16163(.A(new_n16227_), .B(\a[20] ), .Y(new_n16228_));
  XOR2X1   g16164(.A(new_n16228_), .B(new_n16224_), .Y(new_n16229_));
  NOR2X1   g16165(.A(new_n16118_), .B(new_n16116_), .Y(new_n16230_));
  INVX1    g16166(.A(new_n16123_), .Y(new_n16231_));
  AOI21X1  g16167(.A0(new_n16231_), .A1(new_n16119_), .B0(new_n16230_), .Y(new_n16232_));
  XOR2X1   g16168(.A(new_n16232_), .B(new_n16229_), .Y(new_n16233_));
  AOI22X1  g16169(.A0(new_n12285_), .A1(new_n3390_), .B0(new_n12074_), .B1(new_n3232_), .Y(new_n16234_));
  OAI21X1  g16170(.A0(new_n14086_), .A1(new_n3545_), .B0(new_n16234_), .Y(new_n16235_));
  AOI21X1  g16171(.A0(new_n14480_), .A1(new_n3234_), .B0(new_n16235_), .Y(new_n16236_));
  XOR2X1   g16172(.A(new_n16236_), .B(\a[17] ), .Y(new_n16237_));
  XOR2X1   g16173(.A(new_n16237_), .B(new_n16233_), .Y(new_n16238_));
  NOR2X1   g16174(.A(new_n16128_), .B(new_n16124_), .Y(new_n16239_));
  INVX1    g16175(.A(new_n16133_), .Y(new_n16240_));
  AOI21X1  g16176(.A0(new_n16240_), .A1(new_n16129_), .B0(new_n16239_), .Y(new_n16241_));
  XOR2X1   g16177(.A(new_n16241_), .B(new_n16238_), .Y(new_n16242_));
  AOI22X1  g16178(.A0(new_n14087_), .A1(new_n3628_), .B0(new_n14084_), .B1(new_n3908_), .Y(new_n16243_));
  OAI21X1  g16179(.A0(new_n14648_), .A1(new_n3983_), .B0(new_n16243_), .Y(new_n16244_));
  AOI21X1  g16180(.A0(new_n14651_), .A1(new_n3624_), .B0(new_n16244_), .Y(new_n16245_));
  XOR2X1   g16181(.A(new_n16245_), .B(\a[14] ), .Y(new_n16246_));
  XOR2X1   g16182(.A(new_n16246_), .B(new_n16242_), .Y(new_n16247_));
  NOR2X1   g16183(.A(new_n16137_), .B(new_n16134_), .Y(new_n16248_));
  INVX1    g16184(.A(new_n16142_), .Y(new_n16249_));
  AOI21X1  g16185(.A0(new_n16249_), .A1(new_n16138_), .B0(new_n16248_), .Y(new_n16250_));
  XOR2X1   g16186(.A(new_n16250_), .B(new_n16247_), .Y(new_n16251_));
  AOI22X1  g16187(.A0(new_n14946_), .A1(new_n4247_), .B0(new_n14804_), .B1(new_n4078_), .Y(new_n16252_));
  OAI21X1  g16188(.A0(new_n15235_), .A1(new_n4427_), .B0(new_n16252_), .Y(new_n16253_));
  AOI21X1  g16189(.A0(new_n15381_), .A1(new_n4080_), .B0(new_n16253_), .Y(new_n16254_));
  XOR2X1   g16190(.A(new_n16254_), .B(\a[11] ), .Y(new_n16255_));
  XOR2X1   g16191(.A(new_n16255_), .B(new_n16251_), .Y(new_n16256_));
  NOR2X1   g16192(.A(new_n16145_), .B(new_n16143_), .Y(new_n16257_));
  INVX1    g16193(.A(new_n16150_), .Y(new_n16258_));
  AOI21X1  g16194(.A0(new_n16258_), .A1(new_n16146_), .B0(new_n16257_), .Y(new_n16259_));
  AOI22X1  g16195(.A0(new_n15362_), .A1(new_n9681_), .B0(new_n15234_), .B1(new_n4635_), .Y(new_n16260_));
  OAI21X1  g16196(.A0(new_n15373_), .A1(new_n4868_), .B0(new_n16260_), .Y(new_n16261_));
  XOR2X1   g16197(.A(new_n16261_), .B(new_n2995_), .Y(new_n16262_));
  XOR2X1   g16198(.A(new_n16262_), .B(new_n16259_), .Y(new_n16263_));
  XOR2X1   g16199(.A(new_n16263_), .B(new_n16256_), .Y(new_n16264_));
  NOR2X1   g16200(.A(new_n16153_), .B(new_n16151_), .Y(new_n16265_));
  INVX1    g16201(.A(new_n16158_), .Y(new_n16266_));
  AOI21X1  g16202(.A0(new_n16266_), .A1(new_n16154_), .B0(new_n16265_), .Y(new_n16267_));
  XOR2X1   g16203(.A(new_n16267_), .B(new_n16264_), .Y(new_n16268_));
  OR2X1    g16204(.A(new_n16161_), .B(new_n16159_), .Y(new_n16269_));
  XOR2X1   g16205(.A(new_n16266_), .B(new_n16154_), .Y(new_n16270_));
  XOR2X1   g16206(.A(new_n16161_), .B(new_n16270_), .Y(new_n16271_));
  OAI21X1  g16207(.A0(new_n16164_), .A1(new_n16271_), .B0(new_n16269_), .Y(new_n16272_));
  XOR2X1   g16208(.A(new_n16272_), .B(new_n16268_), .Y(new_n16273_));
  XOR2X1   g16209(.A(new_n16273_), .B(new_n16167_), .Y(\result[12] ));
  AND2X1   g16210(.A(new_n16273_), .B(new_n16167_), .Y(new_n16275_));
  NOR2X1   g16211(.A(new_n16267_), .B(new_n16264_), .Y(new_n16276_));
  AOI21X1  g16212(.A0(new_n16272_), .A1(new_n16268_), .B0(new_n16276_), .Y(new_n16277_));
  OR2X1    g16213(.A(new_n16262_), .B(new_n16259_), .Y(new_n16278_));
  INVX1    g16214(.A(new_n16256_), .Y(new_n16279_));
  NAND2X1  g16215(.A(new_n16263_), .B(new_n16279_), .Y(new_n16280_));
  AND2X1   g16216(.A(new_n16280_), .B(new_n16278_), .Y(new_n16281_));
  AND2X1   g16217(.A(new_n16187_), .B(new_n16171_), .Y(new_n16282_));
  OR2X1    g16218(.A(new_n16282_), .B(new_n16190_), .Y(new_n16283_));
  AND2X1   g16219(.A(new_n15362_), .B(new_n7946_), .Y(new_n16284_));
  XOR2X1   g16220(.A(new_n16284_), .B(new_n2995_), .Y(new_n16285_));
  NAND3X1  g16221(.A(new_n2166_), .B(new_n1110_), .C(new_n476_), .Y(new_n16286_));
  OAI22X1  g16222(.A0(new_n102_), .A1(new_n72_), .B0(new_n81_), .B1(new_n69_), .Y(new_n16287_));
  OR4X1    g16223(.A(new_n16287_), .B(new_n1183_), .C(new_n511_), .D(new_n432_), .Y(new_n16288_));
  OR4X1    g16224(.A(new_n16288_), .B(new_n1639_), .C(new_n1478_), .D(new_n1224_), .Y(new_n16289_));
  OR4X1    g16225(.A(new_n16289_), .B(new_n16286_), .C(new_n7432_), .D(new_n1396_), .Y(new_n16290_));
  NOR3X1   g16226(.A(new_n16290_), .B(new_n1866_), .C(new_n1716_), .Y(new_n16291_));
  XOR2X1   g16227(.A(new_n16291_), .B(new_n16085_), .Y(new_n16292_));
  XOR2X1   g16228(.A(new_n16292_), .B(new_n16285_), .Y(new_n16293_));
  XOR2X1   g16229(.A(new_n16293_), .B(new_n16283_), .Y(new_n16294_));
  AOI22X1  g16230(.A0(new_n12104_), .A1(new_n1890_), .B0(new_n12102_), .B1(new_n1884_), .Y(new_n16295_));
  OAI21X1  g16231(.A0(new_n12840_), .A1(new_n3498_), .B0(new_n16295_), .Y(new_n16296_));
  AOI21X1  g16232(.A0(new_n12859_), .A1(new_n407_), .B0(new_n16296_), .Y(new_n16297_));
  XOR2X1   g16233(.A(new_n16297_), .B(new_n16294_), .Y(new_n16298_));
  AOI22X1  g16234(.A0(new_n12097_), .A1(new_n2185_), .B0(new_n12095_), .B1(new_n2095_), .Y(new_n16299_));
  OAI21X1  g16235(.A0(new_n13366_), .A1(new_n2140_), .B0(new_n16299_), .Y(new_n16300_));
  AOI21X1  g16236(.A0(new_n13093_), .A1(new_n2062_), .B0(new_n16300_), .Y(new_n16301_));
  XOR2X1   g16237(.A(new_n16301_), .B(\a[29] ), .Y(new_n16302_));
  XOR2X1   g16238(.A(new_n16302_), .B(new_n16298_), .Y(new_n16303_));
  NOR2X1   g16239(.A(new_n16195_), .B(new_n16192_), .Y(new_n16304_));
  AOI21X1  g16240(.A0(new_n16198_), .A1(new_n16196_), .B0(new_n16304_), .Y(new_n16305_));
  XOR2X1   g16241(.A(new_n16305_), .B(new_n16303_), .Y(new_n16306_));
  AOI22X1  g16242(.A0(new_n12090_), .A1(new_n2424_), .B0(new_n12088_), .B1(new_n2418_), .Y(new_n16307_));
  OAI21X1  g16243(.A0(new_n12298_), .A1(new_n2626_), .B0(new_n16307_), .Y(new_n16308_));
  AOI21X1  g16244(.A0(new_n12297_), .A1(new_n2301_), .B0(new_n16308_), .Y(new_n16309_));
  XOR2X1   g16245(.A(new_n16309_), .B(\a[26] ), .Y(new_n16310_));
  XOR2X1   g16246(.A(new_n16310_), .B(new_n16306_), .Y(new_n16311_));
  INVX1    g16247(.A(new_n16203_), .Y(new_n16312_));
  NOR2X1   g16248(.A(new_n16208_), .B(new_n16204_), .Y(new_n16313_));
  AOI21X1  g16249(.A0(new_n16312_), .A1(new_n16199_), .B0(new_n16313_), .Y(new_n16314_));
  XOR2X1   g16250(.A(new_n16314_), .B(new_n16311_), .Y(new_n16315_));
  AOI22X1  g16251(.A0(new_n12083_), .A1(new_n2657_), .B0(new_n12081_), .B1(new_n2696_), .Y(new_n16316_));
  OAI21X1  g16252(.A0(new_n13665_), .A1(new_n2753_), .B0(new_n16316_), .Y(new_n16317_));
  AOI21X1  g16253(.A0(new_n14672_), .A1(new_n2658_), .B0(new_n16317_), .Y(new_n16318_));
  XOR2X1   g16254(.A(new_n16318_), .B(\a[23] ), .Y(new_n16319_));
  XOR2X1   g16255(.A(new_n16319_), .B(new_n16315_), .Y(new_n16320_));
  NOR2X1   g16256(.A(new_n16214_), .B(new_n16210_), .Y(new_n16321_));
  INVX1    g16257(.A(new_n16219_), .Y(new_n16322_));
  AOI21X1  g16258(.A0(new_n16322_), .A1(new_n16215_), .B0(new_n16321_), .Y(new_n16323_));
  XOR2X1   g16259(.A(new_n16323_), .B(new_n16320_), .Y(new_n16324_));
  AOI22X1  g16260(.A0(new_n12076_), .A1(new_n2875_), .B0(new_n12018_), .B1(new_n3099_), .Y(new_n16325_));
  OAI21X1  g16261(.A0(new_n13679_), .A1(new_n3152_), .B0(new_n16325_), .Y(new_n16326_));
  AOI21X1  g16262(.A0(new_n13678_), .A1(new_n2876_), .B0(new_n16326_), .Y(new_n16327_));
  XOR2X1   g16263(.A(new_n16327_), .B(\a[20] ), .Y(new_n16328_));
  XOR2X1   g16264(.A(new_n16328_), .B(new_n16324_), .Y(new_n16329_));
  NOR2X1   g16265(.A(new_n16223_), .B(new_n16220_), .Y(new_n16330_));
  INVX1    g16266(.A(new_n16228_), .Y(new_n16331_));
  AOI21X1  g16267(.A0(new_n16331_), .A1(new_n16224_), .B0(new_n16330_), .Y(new_n16332_));
  XOR2X1   g16268(.A(new_n16332_), .B(new_n16329_), .Y(new_n16333_));
  INVX1    g16269(.A(new_n16333_), .Y(new_n16334_));
  OR2X1    g16270(.A(new_n16232_), .B(new_n16229_), .Y(new_n16335_));
  INVX1    g16271(.A(new_n16233_), .Y(new_n16336_));
  OAI21X1  g16272(.A0(new_n16237_), .A1(new_n16336_), .B0(new_n16335_), .Y(new_n16337_));
  AOI22X1  g16273(.A0(new_n14085_), .A1(new_n3390_), .B0(new_n12285_), .B1(new_n3232_), .Y(new_n16338_));
  OAI21X1  g16274(.A0(new_n14088_), .A1(new_n3545_), .B0(new_n16338_), .Y(new_n16339_));
  AOI21X1  g16275(.A0(new_n14491_), .A1(new_n3234_), .B0(new_n16339_), .Y(new_n16340_));
  XOR2X1   g16276(.A(new_n16340_), .B(\a[17] ), .Y(new_n16341_));
  XOR2X1   g16277(.A(new_n16341_), .B(new_n16337_), .Y(new_n16342_));
  XOR2X1   g16278(.A(new_n16342_), .B(new_n16334_), .Y(new_n16343_));
  AOI22X1  g16279(.A0(new_n14642_), .A1(new_n3908_), .B0(new_n14084_), .B1(new_n3628_), .Y(new_n16344_));
  OAI21X1  g16280(.A0(new_n14805_), .A1(new_n3983_), .B0(new_n16344_), .Y(new_n16345_));
  AOI21X1  g16281(.A0(new_n14809_), .A1(new_n3624_), .B0(new_n16345_), .Y(new_n16346_));
  XOR2X1   g16282(.A(new_n16346_), .B(\a[14] ), .Y(new_n16347_));
  XOR2X1   g16283(.A(new_n16347_), .B(new_n16343_), .Y(new_n16348_));
  OR2X1    g16284(.A(new_n16241_), .B(new_n16238_), .Y(new_n16349_));
  INVX1    g16285(.A(new_n16242_), .Y(new_n16350_));
  OAI21X1  g16286(.A0(new_n16246_), .A1(new_n16350_), .B0(new_n16349_), .Y(new_n16351_));
  INVX1    g16287(.A(new_n16351_), .Y(new_n16352_));
  XOR2X1   g16288(.A(new_n16352_), .B(new_n16348_), .Y(new_n16353_));
  AND2X1   g16289(.A(new_n16250_), .B(new_n16247_), .Y(new_n16354_));
  OR2X1    g16290(.A(new_n16250_), .B(new_n16247_), .Y(new_n16355_));
  OAI21X1  g16291(.A0(new_n16255_), .A1(new_n16354_), .B0(new_n16355_), .Y(new_n16356_));
  AOI22X1  g16292(.A0(new_n15087_), .A1(new_n4247_), .B0(new_n14946_), .B1(new_n4078_), .Y(new_n16357_));
  OAI21X1  g16293(.A0(new_n15363_), .A1(new_n4427_), .B0(new_n16357_), .Y(new_n16358_));
  AOI21X1  g16294(.A0(new_n15240_), .A1(new_n4080_), .B0(new_n16358_), .Y(new_n16359_));
  XOR2X1   g16295(.A(new_n16359_), .B(\a[11] ), .Y(new_n16360_));
  XOR2X1   g16296(.A(new_n16360_), .B(new_n16356_), .Y(new_n16361_));
  XOR2X1   g16297(.A(new_n16361_), .B(new_n16353_), .Y(new_n16362_));
  XOR2X1   g16298(.A(new_n16362_), .B(new_n16281_), .Y(new_n16363_));
  XOR2X1   g16299(.A(new_n16363_), .B(new_n16277_), .Y(new_n16364_));
  XOR2X1   g16300(.A(new_n16364_), .B(new_n16275_), .Y(\result[13] ));
  AND2X1   g16301(.A(new_n16364_), .B(new_n16275_), .Y(new_n16366_));
  OR2X1    g16302(.A(new_n16302_), .B(new_n16298_), .Y(new_n16367_));
  INVX1    g16303(.A(new_n16303_), .Y(new_n16368_));
  OAI21X1  g16304(.A0(new_n16305_), .A1(new_n16368_), .B0(new_n16367_), .Y(new_n16369_));
  AOI22X1  g16305(.A0(new_n12102_), .A1(new_n1890_), .B0(new_n12099_), .B1(new_n1884_), .Y(new_n16370_));
  OAI21X1  g16306(.A0(new_n12839_), .A1(new_n3498_), .B0(new_n16370_), .Y(new_n16371_));
  AOI21X1  g16307(.A0(new_n12855_), .A1(new_n407_), .B0(new_n16371_), .Y(new_n16372_));
  NAND2X1  g16308(.A(new_n16292_), .B(new_n16285_), .Y(new_n16373_));
  OAI21X1  g16309(.A0(new_n16291_), .A1(new_n16085_), .B0(new_n16373_), .Y(new_n16374_));
  OR4X1    g16310(.A(new_n1153_), .B(new_n546_), .C(new_n579_), .D(new_n395_), .Y(new_n16375_));
  OR4X1    g16311(.A(new_n350_), .B(new_n850_), .C(new_n183_), .D(new_n175_), .Y(new_n16376_));
  OR4X1    g16312(.A(new_n16376_), .B(new_n2806_), .C(new_n2794_), .D(new_n887_), .Y(new_n16377_));
  OR4X1    g16313(.A(new_n16377_), .B(new_n16375_), .C(new_n8642_), .D(new_n7137_), .Y(new_n16378_));
  OR4X1    g16314(.A(new_n16378_), .B(new_n7856_), .C(new_n2091_), .D(new_n946_), .Y(new_n16379_));
  NOR2X1   g16315(.A(new_n16379_), .B(new_n1264_), .Y(new_n16380_));
  XOR2X1   g16316(.A(new_n16380_), .B(new_n16374_), .Y(new_n16381_));
  XOR2X1   g16317(.A(new_n16381_), .B(new_n16372_), .Y(new_n16382_));
  INVX1    g16318(.A(new_n16382_), .Y(new_n16383_));
  AND2X1   g16319(.A(new_n16293_), .B(new_n16283_), .Y(new_n16384_));
  INVX1    g16320(.A(new_n16297_), .Y(new_n16385_));
  AOI21X1  g16321(.A0(new_n16385_), .A1(new_n16294_), .B0(new_n16384_), .Y(new_n16386_));
  XOR2X1   g16322(.A(new_n16386_), .B(new_n16383_), .Y(new_n16387_));
  OAI22X1  g16323(.A0(new_n13090_), .A1(new_n2186_), .B0(new_n13366_), .B1(new_n2431_), .Y(new_n16388_));
  AOI21X1  g16324(.A0(new_n12090_), .A1(new_n2139_), .B0(new_n16388_), .Y(new_n16389_));
  OAI21X1  g16325(.A0(new_n13116_), .A1(new_n2063_), .B0(new_n16389_), .Y(new_n16390_));
  XOR2X1   g16326(.A(new_n16390_), .B(new_n74_), .Y(new_n16391_));
  XOR2X1   g16327(.A(new_n16391_), .B(new_n16387_), .Y(new_n16392_));
  XOR2X1   g16328(.A(new_n16392_), .B(new_n16369_), .Y(new_n16393_));
  AOI22X1  g16329(.A0(new_n12088_), .A1(new_n2424_), .B0(new_n12085_), .B1(new_n2418_), .Y(new_n16394_));
  OAI21X1  g16330(.A0(new_n13321_), .A1(new_n2626_), .B0(new_n16394_), .Y(new_n16395_));
  AOI21X1  g16331(.A0(new_n13344_), .A1(new_n2301_), .B0(new_n16395_), .Y(new_n16396_));
  XOR2X1   g16332(.A(new_n16396_), .B(\a[26] ), .Y(new_n16397_));
  XOR2X1   g16333(.A(new_n16397_), .B(new_n16393_), .Y(new_n16398_));
  OR2X1    g16334(.A(new_n16310_), .B(new_n16306_), .Y(new_n16399_));
  INVX1    g16335(.A(new_n16311_), .Y(new_n16400_));
  OAI21X1  g16336(.A0(new_n16314_), .A1(new_n16400_), .B0(new_n16399_), .Y(new_n16401_));
  XOR2X1   g16337(.A(new_n16401_), .B(new_n16398_), .Y(new_n16402_));
  AOI22X1  g16338(.A0(new_n12081_), .A1(new_n2657_), .B0(new_n12079_), .B1(new_n2696_), .Y(new_n16403_));
  OAI21X1  g16339(.A0(new_n13700_), .A1(new_n2753_), .B0(new_n16403_), .Y(new_n16404_));
  AOI21X1  g16340(.A0(new_n13699_), .A1(new_n2658_), .B0(new_n16404_), .Y(new_n16405_));
  XOR2X1   g16341(.A(new_n16405_), .B(new_n70_), .Y(new_n16406_));
  XOR2X1   g16342(.A(new_n16406_), .B(new_n16402_), .Y(new_n16407_));
  OR2X1    g16343(.A(new_n16319_), .B(new_n16315_), .Y(new_n16408_));
  INVX1    g16344(.A(new_n16320_), .Y(new_n16409_));
  OAI21X1  g16345(.A0(new_n16323_), .A1(new_n16409_), .B0(new_n16408_), .Y(new_n16410_));
  XOR2X1   g16346(.A(new_n16410_), .B(new_n16407_), .Y(new_n16411_));
  AOI22X1  g16347(.A0(new_n12074_), .A1(new_n3099_), .B0(new_n12018_), .B1(new_n2875_), .Y(new_n16412_));
  OAI21X1  g16348(.A0(new_n12292_), .A1(new_n3152_), .B0(new_n16412_), .Y(new_n16413_));
  AOI21X1  g16349(.A0(new_n12291_), .A1(new_n2876_), .B0(new_n16413_), .Y(new_n16414_));
  XOR2X1   g16350(.A(new_n16414_), .B(new_n1920_), .Y(new_n16415_));
  XOR2X1   g16351(.A(new_n16415_), .B(new_n16411_), .Y(new_n16416_));
  OR2X1    g16352(.A(new_n16328_), .B(new_n16324_), .Y(new_n16417_));
  INVX1    g16353(.A(new_n16329_), .Y(new_n16418_));
  OAI21X1  g16354(.A0(new_n16332_), .A1(new_n16418_), .B0(new_n16417_), .Y(new_n16419_));
  XOR2X1   g16355(.A(new_n16419_), .B(new_n16416_), .Y(new_n16420_));
  AOI22X1  g16356(.A0(new_n14087_), .A1(new_n3390_), .B0(new_n14085_), .B1(new_n3232_), .Y(new_n16421_));
  OAI21X1  g16357(.A0(new_n14643_), .A1(new_n3545_), .B0(new_n16421_), .Y(new_n16422_));
  AOI21X1  g16358(.A0(new_n14106_), .A1(new_n3234_), .B0(new_n16422_), .Y(new_n16423_));
  XOR2X1   g16359(.A(new_n16423_), .B(\a[17] ), .Y(new_n16424_));
  XOR2X1   g16360(.A(new_n16424_), .B(new_n16420_), .Y(new_n16425_));
  OR2X1    g16361(.A(new_n16237_), .B(new_n16336_), .Y(new_n16426_));
  AOI21X1  g16362(.A0(new_n16426_), .A1(new_n16335_), .B0(new_n16341_), .Y(new_n16427_));
  NOR2X1   g16363(.A(new_n16342_), .B(new_n16333_), .Y(new_n16428_));
  NOR2X1   g16364(.A(new_n16428_), .B(new_n16427_), .Y(new_n16429_));
  XOR2X1   g16365(.A(new_n16429_), .B(new_n16425_), .Y(new_n16430_));
  AOI22X1  g16366(.A0(new_n14804_), .A1(new_n3908_), .B0(new_n14642_), .B1(new_n3628_), .Y(new_n16431_));
  OAI21X1  g16367(.A0(new_n15088_), .A1(new_n3983_), .B0(new_n16431_), .Y(new_n16432_));
  AOI21X1  g16368(.A0(new_n14952_), .A1(new_n3624_), .B0(new_n16432_), .Y(new_n16433_));
  XOR2X1   g16369(.A(new_n16433_), .B(\a[14] ), .Y(new_n16434_));
  INVX1    g16370(.A(new_n16434_), .Y(new_n16435_));
  XOR2X1   g16371(.A(new_n16435_), .B(new_n16430_), .Y(new_n16436_));
  NOR2X1   g16372(.A(new_n16347_), .B(new_n16343_), .Y(new_n16437_));
  AOI21X1  g16373(.A0(new_n16351_), .A1(new_n16348_), .B0(new_n16437_), .Y(new_n16438_));
  XOR2X1   g16374(.A(new_n16438_), .B(new_n16436_), .Y(new_n16439_));
  AOI22X1  g16375(.A0(new_n15234_), .A1(new_n4247_), .B0(new_n15087_), .B1(new_n4078_), .Y(new_n16440_));
  OAI21X1  g16376(.A0(new_n15522_), .A1(new_n4427_), .B0(new_n16440_), .Y(new_n16441_));
  AOI21X1  g16377(.A0(new_n15841_), .A1(new_n4080_), .B0(new_n16441_), .Y(new_n16442_));
  XOR2X1   g16378(.A(new_n16442_), .B(\a[11] ), .Y(new_n16443_));
  INVX1    g16379(.A(new_n16443_), .Y(new_n16444_));
  XOR2X1   g16380(.A(new_n16444_), .B(new_n16439_), .Y(new_n16445_));
  INVX1    g16381(.A(new_n16360_), .Y(new_n16446_));
  NOR2X1   g16382(.A(new_n16361_), .B(new_n16353_), .Y(new_n16447_));
  AOI21X1  g16383(.A0(new_n16446_), .A1(new_n16356_), .B0(new_n16447_), .Y(new_n16448_));
  XOR2X1   g16384(.A(new_n16448_), .B(new_n16445_), .Y(new_n16449_));
  AND2X1   g16385(.A(new_n16267_), .B(new_n16264_), .Y(new_n16450_));
  OR2X1    g16386(.A(new_n16267_), .B(new_n16264_), .Y(new_n16451_));
  NOR2X1   g16387(.A(new_n16161_), .B(new_n16159_), .Y(new_n16452_));
  NOR2X1   g16388(.A(new_n15946_), .B(new_n15973_), .Y(new_n16453_));
  XOR2X1   g16389(.A(new_n15946_), .B(new_n15973_), .Y(new_n16454_));
  OAI21X1  g16390(.A0(new_n15850_), .A1(new_n15847_), .B0(new_n15851_), .Y(new_n16455_));
  OAI21X1  g16391(.A0(new_n15860_), .A1(new_n15852_), .B0(new_n16455_), .Y(new_n16456_));
  AOI21X1  g16392(.A0(new_n16456_), .A1(new_n16454_), .B0(new_n16453_), .Y(new_n16457_));
  NAND2X1  g16393(.A(new_n16064_), .B(new_n15977_), .Y(new_n16458_));
  NOR2X1   g16394(.A(new_n16064_), .B(new_n15977_), .Y(new_n16459_));
  OAI21X1  g16395(.A0(new_n16459_), .A1(new_n16457_), .B0(new_n16458_), .Y(new_n16460_));
  AOI21X1  g16396(.A0(new_n16460_), .A1(new_n16162_), .B0(new_n16452_), .Y(new_n16461_));
  OAI21X1  g16397(.A0(new_n16461_), .A1(new_n16450_), .B0(new_n16451_), .Y(new_n16462_));
  NAND2X1  g16398(.A(new_n16280_), .B(new_n16278_), .Y(new_n16463_));
  AND2X1   g16399(.A(new_n16362_), .B(new_n16463_), .Y(new_n16464_));
  XOR2X1   g16400(.A(new_n16362_), .B(new_n16463_), .Y(new_n16465_));
  AOI21X1  g16401(.A0(new_n16465_), .A1(new_n16462_), .B0(new_n16464_), .Y(new_n16466_));
  XOR2X1   g16402(.A(new_n16466_), .B(new_n16449_), .Y(new_n16467_));
  XOR2X1   g16403(.A(new_n16467_), .B(new_n16366_), .Y(\result[14] ));
  OR2X1    g16404(.A(new_n16386_), .B(new_n16382_), .Y(new_n16469_));
  OAI21X1  g16405(.A0(new_n16391_), .A1(new_n16387_), .B0(new_n16469_), .Y(new_n16470_));
  OAI22X1  g16406(.A0(new_n152_), .A1(new_n129_), .B0(new_n119_), .B1(new_n92_), .Y(new_n16471_));
  NAND3X1  g16407(.A(new_n2282_), .B(new_n1071_), .C(new_n971_), .Y(new_n16472_));
  OR4X1    g16408(.A(new_n16472_), .B(new_n1775_), .C(new_n16471_), .D(new_n515_), .Y(new_n16473_));
  OR4X1    g16409(.A(new_n1725_), .B(new_n1701_), .C(new_n1402_), .D(new_n1018_), .Y(new_n16474_));
  OR4X1    g16410(.A(new_n723_), .B(new_n293_), .C(new_n239_), .D(new_n220_), .Y(new_n16475_));
  OR4X1    g16411(.A(new_n16475_), .B(new_n16474_), .C(new_n1005_), .D(new_n1461_), .Y(new_n16476_));
  OR4X1    g16412(.A(new_n16476_), .B(new_n16473_), .C(new_n8327_), .D(new_n7438_), .Y(new_n16477_));
  NOR4X1   g16413(.A(new_n16477_), .B(new_n16380_), .C(new_n16078_), .D(new_n3033_), .Y(new_n16478_));
  INVX1    g16414(.A(new_n16372_), .Y(new_n16479_));
  AND2X1   g16415(.A(new_n16380_), .B(new_n16374_), .Y(new_n16480_));
  AOI21X1  g16416(.A0(new_n16381_), .A1(new_n16479_), .B0(new_n16480_), .Y(new_n16481_));
  NOR3X1   g16417(.A(new_n16477_), .B(new_n16078_), .C(new_n3033_), .Y(new_n16482_));
  NOR3X1   g16418(.A(new_n16482_), .B(new_n16379_), .C(new_n1264_), .Y(new_n16483_));
  NOR3X1   g16419(.A(new_n16483_), .B(new_n16478_), .C(new_n16481_), .Y(new_n16484_));
  OR2X1    g16420(.A(new_n16484_), .B(new_n16481_), .Y(new_n16485_));
  NOR2X1   g16421(.A(new_n16484_), .B(new_n16483_), .Y(new_n16486_));
  INVX1    g16422(.A(new_n16486_), .Y(new_n16487_));
  OAI21X1  g16423(.A0(new_n16487_), .A1(new_n16478_), .B0(new_n16485_), .Y(new_n16488_));
  AOI22X1  g16424(.A0(new_n12099_), .A1(new_n1890_), .B0(new_n12097_), .B1(new_n1884_), .Y(new_n16489_));
  OAI21X1  g16425(.A0(new_n13090_), .A1(new_n3498_), .B0(new_n16489_), .Y(new_n16490_));
  AOI21X1  g16426(.A0(new_n14519_), .A1(new_n407_), .B0(new_n16490_), .Y(new_n16491_));
  XOR2X1   g16427(.A(new_n16491_), .B(new_n16488_), .Y(new_n16492_));
  OAI22X1  g16428(.A0(new_n13366_), .A1(new_n2186_), .B0(new_n13118_), .B1(new_n2431_), .Y(new_n16493_));
  AOI21X1  g16429(.A0(new_n12088_), .A1(new_n2139_), .B0(new_n16493_), .Y(new_n16494_));
  OAI21X1  g16430(.A0(new_n14590_), .A1(new_n2063_), .B0(new_n16494_), .Y(new_n16495_));
  XOR2X1   g16431(.A(new_n16495_), .B(new_n74_), .Y(new_n16496_));
  XOR2X1   g16432(.A(new_n16496_), .B(new_n16492_), .Y(new_n16497_));
  XOR2X1   g16433(.A(new_n16497_), .B(new_n16470_), .Y(new_n16498_));
  AOI22X1  g16434(.A0(new_n12085_), .A1(new_n2424_), .B0(new_n12083_), .B1(new_n2418_), .Y(new_n16499_));
  OAI21X1  g16435(.A0(new_n13320_), .A1(new_n2626_), .B0(new_n16499_), .Y(new_n16500_));
  AOI21X1  g16436(.A0(new_n14510_), .A1(new_n2301_), .B0(new_n16500_), .Y(new_n16501_));
  XOR2X1   g16437(.A(new_n16501_), .B(\a[26] ), .Y(new_n16502_));
  XOR2X1   g16438(.A(new_n16502_), .B(new_n16498_), .Y(new_n16503_));
  AND2X1   g16439(.A(new_n16392_), .B(new_n16369_), .Y(new_n16504_));
  INVX1    g16440(.A(new_n16397_), .Y(new_n16505_));
  AOI21X1  g16441(.A0(new_n16505_), .A1(new_n16393_), .B0(new_n16504_), .Y(new_n16506_));
  XOR2X1   g16442(.A(new_n16506_), .B(new_n16503_), .Y(new_n16507_));
  AOI22X1  g16443(.A0(new_n12079_), .A1(new_n2657_), .B0(new_n12076_), .B1(new_n2696_), .Y(new_n16508_));
  OAI21X1  g16444(.A0(new_n13691_), .A1(new_n2753_), .B0(new_n16508_), .Y(new_n16509_));
  AOI21X1  g16445(.A0(new_n13690_), .A1(new_n2658_), .B0(new_n16509_), .Y(new_n16510_));
  XOR2X1   g16446(.A(new_n16510_), .B(\a[23] ), .Y(new_n16511_));
  XOR2X1   g16447(.A(new_n16511_), .B(new_n16507_), .Y(new_n16512_));
  OR2X1    g16448(.A(new_n16314_), .B(new_n16400_), .Y(new_n16513_));
  NAND3X1  g16449(.A(new_n16398_), .B(new_n16513_), .C(new_n16399_), .Y(new_n16514_));
  AOI21X1  g16450(.A0(new_n16513_), .A1(new_n16399_), .B0(new_n16398_), .Y(new_n16515_));
  AOI21X1  g16451(.A0(new_n16406_), .A1(new_n16514_), .B0(new_n16515_), .Y(new_n16516_));
  XOR2X1   g16452(.A(new_n16516_), .B(new_n16512_), .Y(new_n16517_));
  AOI22X1  g16453(.A0(new_n12285_), .A1(new_n3099_), .B0(new_n12074_), .B1(new_n2875_), .Y(new_n16518_));
  OAI21X1  g16454(.A0(new_n14086_), .A1(new_n3152_), .B0(new_n16518_), .Y(new_n16519_));
  AOI21X1  g16455(.A0(new_n14480_), .A1(new_n2876_), .B0(new_n16519_), .Y(new_n16520_));
  XOR2X1   g16456(.A(new_n16520_), .B(\a[20] ), .Y(new_n16521_));
  XOR2X1   g16457(.A(new_n16521_), .B(new_n16517_), .Y(new_n16522_));
  OR2X1    g16458(.A(new_n16323_), .B(new_n16409_), .Y(new_n16523_));
  NAND3X1  g16459(.A(new_n16407_), .B(new_n16523_), .C(new_n16408_), .Y(new_n16524_));
  AOI21X1  g16460(.A0(new_n16523_), .A1(new_n16408_), .B0(new_n16407_), .Y(new_n16525_));
  AOI21X1  g16461(.A0(new_n16415_), .A1(new_n16524_), .B0(new_n16525_), .Y(new_n16526_));
  XOR2X1   g16462(.A(new_n16526_), .B(new_n16522_), .Y(new_n16527_));
  AOI22X1  g16463(.A0(new_n14087_), .A1(new_n3232_), .B0(new_n14084_), .B1(new_n3390_), .Y(new_n16528_));
  OAI21X1  g16464(.A0(new_n14648_), .A1(new_n3545_), .B0(new_n16528_), .Y(new_n16529_));
  AOI21X1  g16465(.A0(new_n14651_), .A1(new_n3234_), .B0(new_n16529_), .Y(new_n16530_));
  XOR2X1   g16466(.A(new_n16530_), .B(\a[17] ), .Y(new_n16531_));
  XOR2X1   g16467(.A(new_n16531_), .B(new_n16527_), .Y(new_n16532_));
  INVX1    g16468(.A(new_n16532_), .Y(new_n16533_));
  OR2X1    g16469(.A(new_n16332_), .B(new_n16418_), .Y(new_n16534_));
  AOI21X1  g16470(.A0(new_n16534_), .A1(new_n16417_), .B0(new_n16416_), .Y(new_n16535_));
  NOR2X1   g16471(.A(new_n16424_), .B(new_n16420_), .Y(new_n16536_));
  NOR2X1   g16472(.A(new_n16536_), .B(new_n16535_), .Y(new_n16537_));
  XOR2X1   g16473(.A(new_n16537_), .B(new_n16533_), .Y(new_n16538_));
  AOI22X1  g16474(.A0(new_n14946_), .A1(new_n3908_), .B0(new_n14804_), .B1(new_n3628_), .Y(new_n16539_));
  OAI21X1  g16475(.A0(new_n15235_), .A1(new_n3983_), .B0(new_n16539_), .Y(new_n16540_));
  AOI21X1  g16476(.A0(new_n15381_), .A1(new_n3624_), .B0(new_n16540_), .Y(new_n16541_));
  XOR2X1   g16477(.A(new_n16541_), .B(\a[14] ), .Y(new_n16542_));
  XOR2X1   g16478(.A(new_n16542_), .B(new_n16538_), .Y(new_n16543_));
  OAI21X1  g16479(.A0(new_n16428_), .A1(new_n16427_), .B0(new_n16425_), .Y(new_n16544_));
  OAI21X1  g16480(.A0(new_n16434_), .A1(new_n16430_), .B0(new_n16544_), .Y(new_n16545_));
  AOI22X1  g16481(.A0(new_n15362_), .A1(new_n9026_), .B0(new_n15234_), .B1(new_n4078_), .Y(new_n16546_));
  OAI21X1  g16482(.A0(new_n15373_), .A1(new_n4245_), .B0(new_n16546_), .Y(new_n16547_));
  XOR2X1   g16483(.A(new_n16547_), .B(new_n2911_), .Y(new_n16548_));
  XOR2X1   g16484(.A(new_n16548_), .B(new_n16545_), .Y(new_n16549_));
  XOR2X1   g16485(.A(new_n16549_), .B(new_n16543_), .Y(new_n16550_));
  NOR2X1   g16486(.A(new_n16438_), .B(new_n16436_), .Y(new_n16551_));
  AOI21X1  g16487(.A0(new_n16444_), .A1(new_n16439_), .B0(new_n16551_), .Y(new_n16552_));
  XOR2X1   g16488(.A(new_n16552_), .B(new_n16550_), .Y(new_n16553_));
  INVX1    g16489(.A(new_n16553_), .Y(new_n16554_));
  XOR2X1   g16490(.A(new_n16443_), .B(new_n16439_), .Y(new_n16555_));
  NOR2X1   g16491(.A(new_n16448_), .B(new_n16555_), .Y(new_n16556_));
  XOR2X1   g16492(.A(new_n16448_), .B(new_n16555_), .Y(new_n16557_));
  NAND2X1  g16493(.A(new_n16362_), .B(new_n16463_), .Y(new_n16558_));
  OAI21X1  g16494(.A0(new_n16363_), .A1(new_n16277_), .B0(new_n16558_), .Y(new_n16559_));
  AOI21X1  g16495(.A0(new_n16559_), .A1(new_n16557_), .B0(new_n16556_), .Y(new_n16560_));
  XOR2X1   g16496(.A(new_n16560_), .B(new_n16554_), .Y(new_n16561_));
  AND2X1   g16497(.A(new_n16467_), .B(new_n16366_), .Y(new_n16562_));
  XOR2X1   g16498(.A(new_n16562_), .B(new_n16561_), .Y(\result[15] ));
  AND2X1   g16499(.A(new_n16562_), .B(new_n16561_), .Y(new_n16564_));
  NOR2X1   g16500(.A(new_n16552_), .B(new_n16550_), .Y(new_n16565_));
  INVX1    g16501(.A(new_n16565_), .Y(new_n16566_));
  OAI21X1  g16502(.A0(new_n16560_), .A1(new_n16554_), .B0(new_n16566_), .Y(new_n16567_));
  INVX1    g16503(.A(new_n16545_), .Y(new_n16568_));
  INVX1    g16504(.A(new_n16549_), .Y(new_n16569_));
  NAND2X1  g16505(.A(new_n16569_), .B(new_n16543_), .Y(new_n16570_));
  OAI21X1  g16506(.A0(new_n16548_), .A1(new_n16568_), .B0(new_n16570_), .Y(new_n16571_));
  OR2X1    g16507(.A(new_n16487_), .B(new_n16478_), .Y(new_n16572_));
  AOI21X1  g16508(.A0(new_n16572_), .A1(new_n16485_), .B0(new_n16491_), .Y(new_n16573_));
  NOR2X1   g16509(.A(new_n16496_), .B(new_n16492_), .Y(new_n16574_));
  NOR2X1   g16510(.A(new_n16574_), .B(new_n16573_), .Y(new_n16575_));
  AND2X1   g16511(.A(new_n15362_), .B(new_n7865_), .Y(new_n16576_));
  XOR2X1   g16512(.A(new_n16576_), .B(new_n2911_), .Y(new_n16577_));
  INVX1    g16513(.A(new_n1103_), .Y(new_n16578_));
  NOR4X1   g16514(.A(new_n1133_), .B(new_n640_), .C(new_n488_), .D(new_n992_), .Y(new_n16579_));
  NOR4X1   g16515(.A(new_n183_), .B(new_n158_), .C(new_n116_), .D(new_n585_), .Y(new_n16580_));
  NAND3X1  g16516(.A(new_n16580_), .B(new_n16579_), .C(new_n2916_), .Y(new_n16581_));
  OR4X1    g16517(.A(new_n2302_), .B(new_n1210_), .C(new_n429_), .D(new_n194_), .Y(new_n16582_));
  OR4X1    g16518(.A(new_n16582_), .B(new_n1351_), .C(new_n432_), .D(new_n390_), .Y(new_n16583_));
  OR4X1    g16519(.A(new_n16583_), .B(new_n16581_), .C(new_n2930_), .D(new_n1073_), .Y(new_n16584_));
  NOR3X1   g16520(.A(new_n16584_), .B(new_n2148_), .C(new_n16578_), .Y(new_n16585_));
  XOR2X1   g16521(.A(new_n16585_), .B(new_n16380_), .Y(new_n16586_));
  XOR2X1   g16522(.A(new_n16586_), .B(new_n16577_), .Y(new_n16587_));
  AOI22X1  g16523(.A0(new_n12097_), .A1(new_n1890_), .B0(new_n12095_), .B1(new_n1884_), .Y(new_n16588_));
  OAI21X1  g16524(.A0(new_n13366_), .A1(new_n3498_), .B0(new_n16588_), .Y(new_n16589_));
  AOI21X1  g16525(.A0(new_n13093_), .A1(new_n407_), .B0(new_n16589_), .Y(new_n16590_));
  XOR2X1   g16526(.A(new_n16590_), .B(new_n16587_), .Y(new_n16591_));
  XOR2X1   g16527(.A(new_n16591_), .B(new_n16487_), .Y(new_n16592_));
  XOR2X1   g16528(.A(new_n16592_), .B(new_n16575_), .Y(new_n16593_));
  AOI22X1  g16529(.A0(new_n12090_), .A1(new_n2185_), .B0(new_n12088_), .B1(new_n2095_), .Y(new_n16594_));
  OAI21X1  g16530(.A0(new_n12298_), .A1(new_n2140_), .B0(new_n16594_), .Y(new_n16595_));
  AOI21X1  g16531(.A0(new_n12297_), .A1(new_n2062_), .B0(new_n16595_), .Y(new_n16596_));
  XOR2X1   g16532(.A(new_n16596_), .B(\a[29] ), .Y(new_n16597_));
  XOR2X1   g16533(.A(new_n16597_), .B(new_n16593_), .Y(new_n16598_));
  AOI22X1  g16534(.A0(new_n12083_), .A1(new_n2424_), .B0(new_n12081_), .B1(new_n2418_), .Y(new_n16599_));
  OAI21X1  g16535(.A0(new_n13665_), .A1(new_n2626_), .B0(new_n16599_), .Y(new_n16600_));
  AOI21X1  g16536(.A0(new_n14672_), .A1(new_n2301_), .B0(new_n16600_), .Y(new_n16601_));
  XOR2X1   g16537(.A(new_n16601_), .B(\a[26] ), .Y(new_n16602_));
  XOR2X1   g16538(.A(new_n16602_), .B(new_n16598_), .Y(new_n16603_));
  NAND2X1  g16539(.A(new_n16497_), .B(new_n16470_), .Y(new_n16604_));
  INVX1    g16540(.A(new_n16498_), .Y(new_n16605_));
  OAI21X1  g16541(.A0(new_n16502_), .A1(new_n16605_), .B0(new_n16604_), .Y(new_n16606_));
  XOR2X1   g16542(.A(new_n16606_), .B(new_n16603_), .Y(new_n16607_));
  AOI22X1  g16543(.A0(new_n12076_), .A1(new_n2657_), .B0(new_n12018_), .B1(new_n2696_), .Y(new_n16608_));
  OAI21X1  g16544(.A0(new_n13679_), .A1(new_n2753_), .B0(new_n16608_), .Y(new_n16609_));
  AOI21X1  g16545(.A0(new_n13678_), .A1(new_n2658_), .B0(new_n16609_), .Y(new_n16610_));
  XOR2X1   g16546(.A(new_n16610_), .B(\a[23] ), .Y(new_n16611_));
  XOR2X1   g16547(.A(new_n16611_), .B(new_n16607_), .Y(new_n16612_));
  NOR2X1   g16548(.A(new_n16506_), .B(new_n16503_), .Y(new_n16613_));
  INVX1    g16549(.A(new_n16511_), .Y(new_n16614_));
  AOI21X1  g16550(.A0(new_n16614_), .A1(new_n16507_), .B0(new_n16613_), .Y(new_n16615_));
  XOR2X1   g16551(.A(new_n16615_), .B(new_n16612_), .Y(new_n16616_));
  INVX1    g16552(.A(new_n16616_), .Y(new_n16617_));
  INVX1    g16553(.A(new_n16517_), .Y(new_n16618_));
  OR2X1    g16554(.A(new_n16521_), .B(new_n16618_), .Y(new_n16619_));
  OAI21X1  g16555(.A0(new_n16516_), .A1(new_n16512_), .B0(new_n16619_), .Y(new_n16620_));
  AOI22X1  g16556(.A0(new_n14085_), .A1(new_n3099_), .B0(new_n12285_), .B1(new_n2875_), .Y(new_n16621_));
  OAI21X1  g16557(.A0(new_n14088_), .A1(new_n3152_), .B0(new_n16621_), .Y(new_n16622_));
  AOI21X1  g16558(.A0(new_n14491_), .A1(new_n2876_), .B0(new_n16622_), .Y(new_n16623_));
  XOR2X1   g16559(.A(new_n16623_), .B(\a[20] ), .Y(new_n16624_));
  XOR2X1   g16560(.A(new_n16624_), .B(new_n16620_), .Y(new_n16625_));
  XOR2X1   g16561(.A(new_n16625_), .B(new_n16617_), .Y(new_n16626_));
  AOI22X1  g16562(.A0(new_n14642_), .A1(new_n3390_), .B0(new_n14084_), .B1(new_n3232_), .Y(new_n16627_));
  OAI21X1  g16563(.A0(new_n14805_), .A1(new_n3545_), .B0(new_n16627_), .Y(new_n16628_));
  AOI21X1  g16564(.A0(new_n14809_), .A1(new_n3234_), .B0(new_n16628_), .Y(new_n16629_));
  XOR2X1   g16565(.A(new_n16629_), .B(\a[17] ), .Y(new_n16630_));
  XOR2X1   g16566(.A(new_n16630_), .B(new_n16626_), .Y(new_n16631_));
  INVX1    g16567(.A(new_n16631_), .Y(new_n16632_));
  NOR2X1   g16568(.A(new_n16526_), .B(new_n16522_), .Y(new_n16633_));
  INVX1    g16569(.A(new_n16531_), .Y(new_n16634_));
  AOI21X1  g16570(.A0(new_n16634_), .A1(new_n16527_), .B0(new_n16633_), .Y(new_n16635_));
  XOR2X1   g16571(.A(new_n16635_), .B(new_n16632_), .Y(new_n16636_));
  NOR2X1   g16572(.A(new_n16537_), .B(new_n16532_), .Y(new_n16637_));
  INVX1    g16573(.A(new_n16637_), .Y(new_n16638_));
  OR2X1    g16574(.A(new_n16542_), .B(new_n16538_), .Y(new_n16639_));
  NAND2X1  g16575(.A(new_n16639_), .B(new_n16638_), .Y(new_n16640_));
  AOI22X1  g16576(.A0(new_n15087_), .A1(new_n3908_), .B0(new_n14946_), .B1(new_n3628_), .Y(new_n16641_));
  OAI21X1  g16577(.A0(new_n15363_), .A1(new_n3983_), .B0(new_n16641_), .Y(new_n16642_));
  AOI21X1  g16578(.A0(new_n15240_), .A1(new_n3624_), .B0(new_n16642_), .Y(new_n16643_));
  XOR2X1   g16579(.A(new_n16643_), .B(\a[14] ), .Y(new_n16644_));
  XOR2X1   g16580(.A(new_n16644_), .B(new_n16640_), .Y(new_n16645_));
  XOR2X1   g16581(.A(new_n16645_), .B(new_n16636_), .Y(new_n16646_));
  XOR2X1   g16582(.A(new_n16646_), .B(new_n16571_), .Y(new_n16647_));
  XOR2X1   g16583(.A(new_n16647_), .B(new_n16567_), .Y(new_n16648_));
  XOR2X1   g16584(.A(new_n16648_), .B(new_n16564_), .Y(\result[16] ));
  AND2X1   g16585(.A(new_n16648_), .B(new_n16564_), .Y(new_n16650_));
  INVX1    g16586(.A(new_n16593_), .Y(new_n16651_));
  OR2X1    g16587(.A(new_n16597_), .B(new_n16651_), .Y(new_n16652_));
  OAI21X1  g16588(.A0(new_n16592_), .A1(new_n16575_), .B0(new_n16652_), .Y(new_n16653_));
  AOI22X1  g16589(.A0(new_n12095_), .A1(new_n1890_), .B0(new_n12093_), .B1(new_n1884_), .Y(new_n16654_));
  OAI21X1  g16590(.A0(new_n13118_), .A1(new_n3498_), .B0(new_n16654_), .Y(new_n16655_));
  AOI21X1  g16591(.A0(new_n13117_), .A1(new_n407_), .B0(new_n16655_), .Y(new_n16656_));
  NAND2X1  g16592(.A(new_n16586_), .B(new_n16577_), .Y(new_n16657_));
  OAI21X1  g16593(.A0(new_n16585_), .A1(new_n16380_), .B0(new_n16657_), .Y(new_n16658_));
  OR4X1    g16594(.A(new_n840_), .B(new_n252_), .C(new_n234_), .D(new_n536_), .Y(new_n16659_));
  OR4X1    g16595(.A(new_n16659_), .B(new_n396_), .C(new_n678_), .D(new_n1087_), .Y(new_n16660_));
  OR4X1    g16596(.A(new_n1447_), .B(new_n1100_), .C(new_n728_), .D(new_n306_), .Y(new_n16661_));
  OR4X1    g16597(.A(new_n16661_), .B(new_n16660_), .C(new_n1921_), .D(new_n1163_), .Y(new_n16662_));
  OR2X1    g16598(.A(new_n15424_), .B(new_n15157_), .Y(new_n16663_));
  NOR4X1   g16599(.A(new_n16663_), .B(new_n16662_), .C(new_n8329_), .D(new_n7350_), .Y(new_n16664_));
  XOR2X1   g16600(.A(new_n16664_), .B(new_n16658_), .Y(new_n16665_));
  XOR2X1   g16601(.A(new_n16665_), .B(new_n16656_), .Y(new_n16666_));
  INVX1    g16602(.A(new_n16666_), .Y(new_n16667_));
  INVX1    g16603(.A(new_n16587_), .Y(new_n16668_));
  NOR2X1   g16604(.A(new_n16590_), .B(new_n16668_), .Y(new_n16669_));
  NOR2X1   g16605(.A(new_n16591_), .B(new_n16486_), .Y(new_n16670_));
  NOR2X1   g16606(.A(new_n16670_), .B(new_n16669_), .Y(new_n16671_));
  XOR2X1   g16607(.A(new_n16671_), .B(new_n16667_), .Y(new_n16672_));
  OAI22X1  g16608(.A0(new_n13104_), .A1(new_n2186_), .B0(new_n12298_), .B1(new_n2431_), .Y(new_n16673_));
  AOI21X1  g16609(.A0(new_n12083_), .A1(new_n2139_), .B0(new_n16673_), .Y(new_n16674_));
  OAI21X1  g16610(.A0(new_n13345_), .A1(new_n2063_), .B0(new_n16674_), .Y(new_n16675_));
  XOR2X1   g16611(.A(new_n16675_), .B(new_n74_), .Y(new_n16676_));
  XOR2X1   g16612(.A(new_n16676_), .B(new_n16672_), .Y(new_n16677_));
  XOR2X1   g16613(.A(new_n16677_), .B(new_n16653_), .Y(new_n16678_));
  AOI22X1  g16614(.A0(new_n12081_), .A1(new_n2424_), .B0(new_n12079_), .B1(new_n2418_), .Y(new_n16679_));
  OAI21X1  g16615(.A0(new_n13700_), .A1(new_n2626_), .B0(new_n16679_), .Y(new_n16680_));
  AOI21X1  g16616(.A0(new_n13699_), .A1(new_n2301_), .B0(new_n16680_), .Y(new_n16681_));
  XOR2X1   g16617(.A(new_n16681_), .B(\a[26] ), .Y(new_n16682_));
  XOR2X1   g16618(.A(new_n16682_), .B(new_n16678_), .Y(new_n16683_));
  NOR2X1   g16619(.A(new_n16602_), .B(new_n16598_), .Y(new_n16684_));
  AOI21X1  g16620(.A0(new_n16606_), .A1(new_n16603_), .B0(new_n16684_), .Y(new_n16685_));
  XOR2X1   g16621(.A(new_n16685_), .B(new_n16683_), .Y(new_n16686_));
  AOI22X1  g16622(.A0(new_n12074_), .A1(new_n2696_), .B0(new_n12018_), .B1(new_n2657_), .Y(new_n16687_));
  OAI21X1  g16623(.A0(new_n12292_), .A1(new_n2753_), .B0(new_n16687_), .Y(new_n16688_));
  AOI21X1  g16624(.A0(new_n12291_), .A1(new_n2658_), .B0(new_n16688_), .Y(new_n16689_));
  XOR2X1   g16625(.A(new_n16689_), .B(\a[23] ), .Y(new_n16690_));
  XOR2X1   g16626(.A(new_n16690_), .B(new_n16686_), .Y(new_n16691_));
  INVX1    g16627(.A(new_n16611_), .Y(new_n16692_));
  NOR2X1   g16628(.A(new_n16615_), .B(new_n16612_), .Y(new_n16693_));
  AOI21X1  g16629(.A0(new_n16692_), .A1(new_n16607_), .B0(new_n16693_), .Y(new_n16694_));
  XOR2X1   g16630(.A(new_n16694_), .B(new_n16691_), .Y(new_n16695_));
  AOI22X1  g16631(.A0(new_n14087_), .A1(new_n3099_), .B0(new_n14085_), .B1(new_n2875_), .Y(new_n16696_));
  OAI21X1  g16632(.A0(new_n14643_), .A1(new_n3152_), .B0(new_n16696_), .Y(new_n16697_));
  AOI21X1  g16633(.A0(new_n14106_), .A1(new_n2876_), .B0(new_n16697_), .Y(new_n16698_));
  XOR2X1   g16634(.A(new_n16698_), .B(\a[20] ), .Y(new_n16699_));
  XOR2X1   g16635(.A(new_n16699_), .B(new_n16695_), .Y(new_n16700_));
  INVX1    g16636(.A(new_n16624_), .Y(new_n16701_));
  NOR2X1   g16637(.A(new_n16625_), .B(new_n16617_), .Y(new_n16702_));
  AOI21X1  g16638(.A0(new_n16701_), .A1(new_n16620_), .B0(new_n16702_), .Y(new_n16703_));
  XOR2X1   g16639(.A(new_n16703_), .B(new_n16700_), .Y(new_n16704_));
  AOI22X1  g16640(.A0(new_n14804_), .A1(new_n3390_), .B0(new_n14642_), .B1(new_n3232_), .Y(new_n16705_));
  OAI21X1  g16641(.A0(new_n15088_), .A1(new_n3545_), .B0(new_n16705_), .Y(new_n16706_));
  AOI21X1  g16642(.A0(new_n14952_), .A1(new_n3234_), .B0(new_n16706_), .Y(new_n16707_));
  XOR2X1   g16643(.A(new_n16707_), .B(\a[17] ), .Y(new_n16708_));
  XOR2X1   g16644(.A(new_n16708_), .B(new_n16704_), .Y(new_n16709_));
  INVX1    g16645(.A(new_n16630_), .Y(new_n16710_));
  NOR2X1   g16646(.A(new_n16635_), .B(new_n16631_), .Y(new_n16711_));
  AOI21X1  g16647(.A0(new_n16710_), .A1(new_n16626_), .B0(new_n16711_), .Y(new_n16712_));
  XOR2X1   g16648(.A(new_n16712_), .B(new_n16709_), .Y(new_n16713_));
  AOI22X1  g16649(.A0(new_n15234_), .A1(new_n3908_), .B0(new_n15087_), .B1(new_n3628_), .Y(new_n16714_));
  OAI21X1  g16650(.A0(new_n15522_), .A1(new_n3983_), .B0(new_n16714_), .Y(new_n16715_));
  AOI21X1  g16651(.A0(new_n15841_), .A1(new_n3624_), .B0(new_n16715_), .Y(new_n16716_));
  XOR2X1   g16652(.A(new_n16716_), .B(\a[14] ), .Y(new_n16717_));
  INVX1    g16653(.A(new_n16717_), .Y(new_n16718_));
  XOR2X1   g16654(.A(new_n16718_), .B(new_n16713_), .Y(new_n16719_));
  AOI21X1  g16655(.A0(new_n16639_), .A1(new_n16638_), .B0(new_n16644_), .Y(new_n16720_));
  NOR2X1   g16656(.A(new_n16645_), .B(new_n16636_), .Y(new_n16721_));
  NOR2X1   g16657(.A(new_n16721_), .B(new_n16720_), .Y(new_n16722_));
  XOR2X1   g16658(.A(new_n16722_), .B(new_n16719_), .Y(new_n16723_));
  AND2X1   g16659(.A(new_n16646_), .B(new_n16571_), .Y(new_n16724_));
  AOI21X1  g16660(.A0(new_n16647_), .A1(new_n16567_), .B0(new_n16724_), .Y(new_n16725_));
  XOR2X1   g16661(.A(new_n16725_), .B(new_n16723_), .Y(new_n16726_));
  XOR2X1   g16662(.A(new_n16726_), .B(new_n16650_), .Y(\result[17] ));
  AND2X1   g16663(.A(new_n16726_), .B(new_n16650_), .Y(new_n16728_));
  AOI22X1  g16664(.A0(new_n12093_), .A1(new_n1890_), .B0(new_n12090_), .B1(new_n1884_), .Y(new_n16729_));
  OAI21X1  g16665(.A0(new_n13104_), .A1(new_n3498_), .B0(new_n16729_), .Y(new_n16730_));
  AOI21X1  g16666(.A0(new_n13103_), .A1(new_n407_), .B0(new_n16730_), .Y(new_n16731_));
  INVX1    g16667(.A(new_n1477_), .Y(new_n16732_));
  OR2X1    g16668(.A(new_n7017_), .B(new_n7016_), .Y(new_n16733_));
  NOR3X1   g16669(.A(new_n3457_), .B(new_n1756_), .C(new_n669_), .Y(new_n16734_));
  NOR4X1   g16670(.A(new_n596_), .B(new_n1044_), .C(new_n579_), .D(new_n273_), .Y(new_n16735_));
  NOR4X1   g16671(.A(new_n247_), .B(new_n1087_), .C(new_n155_), .D(new_n1046_), .Y(new_n16736_));
  NAND3X1  g16672(.A(new_n16736_), .B(new_n16735_), .C(new_n16734_), .Y(new_n16737_));
  OR4X1    g16673(.A(new_n16737_), .B(new_n16733_), .C(new_n1629_), .D(new_n16732_), .Y(new_n16738_));
  OR4X1    g16674(.A(new_n16738_), .B(new_n7136_), .C(new_n2113_), .D(new_n402_), .Y(new_n16739_));
  NOR3X1   g16675(.A(new_n16739_), .B(new_n16664_), .C(new_n1937_), .Y(new_n16740_));
  OAI21X1  g16676(.A0(new_n16739_), .A1(new_n1937_), .B0(new_n16664_), .Y(new_n16741_));
  INVX1    g16677(.A(new_n16741_), .Y(new_n16742_));
  NOR3X1   g16678(.A(new_n16742_), .B(new_n16740_), .C(new_n16731_), .Y(new_n16743_));
  NOR2X1   g16679(.A(new_n16743_), .B(new_n16742_), .Y(new_n16744_));
  INVX1    g16680(.A(new_n16744_), .Y(new_n16745_));
  OAI22X1  g16681(.A0(new_n16745_), .A1(new_n16740_), .B0(new_n16743_), .B1(new_n16731_), .Y(new_n16746_));
  INVX1    g16682(.A(new_n16746_), .Y(new_n16747_));
  INVX1    g16683(.A(new_n16656_), .Y(new_n16748_));
  AND2X1   g16684(.A(new_n16664_), .B(new_n16658_), .Y(new_n16749_));
  AOI21X1  g16685(.A0(new_n16665_), .A1(new_n16748_), .B0(new_n16749_), .Y(new_n16750_));
  XOR2X1   g16686(.A(new_n16750_), .B(new_n16747_), .Y(new_n16751_));
  OAI21X1  g16687(.A0(new_n16670_), .A1(new_n16669_), .B0(new_n16667_), .Y(new_n16752_));
  OAI21X1  g16688(.A0(new_n16676_), .A1(new_n16672_), .B0(new_n16752_), .Y(new_n16753_));
  XOR2X1   g16689(.A(new_n16753_), .B(new_n16751_), .Y(new_n16754_));
  AOI22X1  g16690(.A0(new_n12085_), .A1(new_n2185_), .B0(new_n12083_), .B1(new_n2095_), .Y(new_n16755_));
  OAI21X1  g16691(.A0(new_n13320_), .A1(new_n2140_), .B0(new_n16755_), .Y(new_n16756_));
  AOI21X1  g16692(.A0(new_n14510_), .A1(new_n2062_), .B0(new_n16756_), .Y(new_n16757_));
  XOR2X1   g16693(.A(new_n16757_), .B(\a[29] ), .Y(new_n16758_));
  XOR2X1   g16694(.A(new_n16758_), .B(new_n16754_), .Y(new_n16759_));
  AOI22X1  g16695(.A0(new_n12079_), .A1(new_n2424_), .B0(new_n12076_), .B1(new_n2418_), .Y(new_n16760_));
  OAI21X1  g16696(.A0(new_n13691_), .A1(new_n2626_), .B0(new_n16760_), .Y(new_n16761_));
  AOI21X1  g16697(.A0(new_n13690_), .A1(new_n2301_), .B0(new_n16761_), .Y(new_n16762_));
  XOR2X1   g16698(.A(new_n16762_), .B(\a[26] ), .Y(new_n16763_));
  XOR2X1   g16699(.A(new_n16763_), .B(new_n16759_), .Y(new_n16764_));
  INVX1    g16700(.A(new_n16764_), .Y(new_n16765_));
  AND2X1   g16701(.A(new_n16677_), .B(new_n16653_), .Y(new_n16766_));
  INVX1    g16702(.A(new_n16682_), .Y(new_n16767_));
  AOI21X1  g16703(.A0(new_n16767_), .A1(new_n16678_), .B0(new_n16766_), .Y(new_n16768_));
  XOR2X1   g16704(.A(new_n16768_), .B(new_n16765_), .Y(new_n16769_));
  AOI22X1  g16705(.A0(new_n12285_), .A1(new_n2696_), .B0(new_n12074_), .B1(new_n2657_), .Y(new_n16770_));
  OAI21X1  g16706(.A0(new_n14086_), .A1(new_n2753_), .B0(new_n16770_), .Y(new_n16771_));
  AOI21X1  g16707(.A0(new_n14480_), .A1(new_n2658_), .B0(new_n16771_), .Y(new_n16772_));
  XOR2X1   g16708(.A(new_n16772_), .B(\a[23] ), .Y(new_n16773_));
  XOR2X1   g16709(.A(new_n16773_), .B(new_n16769_), .Y(new_n16774_));
  NOR2X1   g16710(.A(new_n16685_), .B(new_n16683_), .Y(new_n16775_));
  INVX1    g16711(.A(new_n16690_), .Y(new_n16776_));
  AOI21X1  g16712(.A0(new_n16776_), .A1(new_n16686_), .B0(new_n16775_), .Y(new_n16777_));
  XOR2X1   g16713(.A(new_n16777_), .B(new_n16774_), .Y(new_n16778_));
  AOI22X1  g16714(.A0(new_n14087_), .A1(new_n2875_), .B0(new_n14084_), .B1(new_n3099_), .Y(new_n16779_));
  OAI21X1  g16715(.A0(new_n14648_), .A1(new_n3152_), .B0(new_n16779_), .Y(new_n16780_));
  AOI21X1  g16716(.A0(new_n14651_), .A1(new_n2876_), .B0(new_n16780_), .Y(new_n16781_));
  XOR2X1   g16717(.A(new_n16781_), .B(\a[20] ), .Y(new_n16782_));
  XOR2X1   g16718(.A(new_n16782_), .B(new_n16778_), .Y(new_n16783_));
  NOR2X1   g16719(.A(new_n16694_), .B(new_n16691_), .Y(new_n16784_));
  INVX1    g16720(.A(new_n16699_), .Y(new_n16785_));
  AOI21X1  g16721(.A0(new_n16785_), .A1(new_n16695_), .B0(new_n16784_), .Y(new_n16786_));
  XOR2X1   g16722(.A(new_n16786_), .B(new_n16783_), .Y(new_n16787_));
  AOI22X1  g16723(.A0(new_n14946_), .A1(new_n3390_), .B0(new_n14804_), .B1(new_n3232_), .Y(new_n16788_));
  OAI21X1  g16724(.A0(new_n15235_), .A1(new_n3545_), .B0(new_n16788_), .Y(new_n16789_));
  AOI21X1  g16725(.A0(new_n15381_), .A1(new_n3234_), .B0(new_n16789_), .Y(new_n16790_));
  XOR2X1   g16726(.A(new_n16790_), .B(\a[17] ), .Y(new_n16791_));
  XOR2X1   g16727(.A(new_n16791_), .B(new_n16787_), .Y(new_n16792_));
  NOR2X1   g16728(.A(new_n16703_), .B(new_n16700_), .Y(new_n16793_));
  INVX1    g16729(.A(new_n16708_), .Y(new_n16794_));
  AOI21X1  g16730(.A0(new_n16794_), .A1(new_n16704_), .B0(new_n16793_), .Y(new_n16795_));
  AOI22X1  g16731(.A0(new_n15362_), .A1(new_n8502_), .B0(new_n15234_), .B1(new_n3628_), .Y(new_n16796_));
  OAI21X1  g16732(.A0(new_n15373_), .A1(new_n3906_), .B0(new_n16796_), .Y(new_n16797_));
  XOR2X1   g16733(.A(new_n16797_), .B(new_n2529_), .Y(new_n16798_));
  XOR2X1   g16734(.A(new_n16798_), .B(new_n16795_), .Y(new_n16799_));
  XOR2X1   g16735(.A(new_n16799_), .B(new_n16792_), .Y(new_n16800_));
  NOR2X1   g16736(.A(new_n16712_), .B(new_n16709_), .Y(new_n16801_));
  AOI21X1  g16737(.A0(new_n16718_), .A1(new_n16713_), .B0(new_n16801_), .Y(new_n16802_));
  XOR2X1   g16738(.A(new_n16802_), .B(new_n16800_), .Y(new_n16803_));
  XOR2X1   g16739(.A(new_n16717_), .B(new_n16713_), .Y(new_n16804_));
  OR2X1    g16740(.A(new_n16722_), .B(new_n16804_), .Y(new_n16805_));
  OAI21X1  g16741(.A0(new_n16725_), .A1(new_n16723_), .B0(new_n16805_), .Y(new_n16806_));
  XOR2X1   g16742(.A(new_n16806_), .B(new_n16803_), .Y(new_n16807_));
  XOR2X1   g16743(.A(new_n16807_), .B(new_n16728_), .Y(\result[18] ));
  AND2X1   g16744(.A(new_n16807_), .B(new_n16728_), .Y(new_n16809_));
  NOR2X1   g16745(.A(new_n16802_), .B(new_n16800_), .Y(new_n16810_));
  AOI21X1  g16746(.A0(new_n16806_), .A1(new_n16803_), .B0(new_n16810_), .Y(new_n16811_));
  INVX1    g16747(.A(new_n16792_), .Y(new_n16812_));
  NOR2X1   g16748(.A(new_n16798_), .B(new_n16795_), .Y(new_n16813_));
  AOI21X1  g16749(.A0(new_n16799_), .A1(new_n16812_), .B0(new_n16813_), .Y(new_n16814_));
  INVX1    g16750(.A(new_n16814_), .Y(new_n16815_));
  AND2X1   g16751(.A(new_n15362_), .B(new_n7464_), .Y(new_n16816_));
  XOR2X1   g16752(.A(new_n16816_), .B(new_n2529_), .Y(new_n16817_));
  OR4X1    g16753(.A(new_n1916_), .B(new_n1664_), .C(new_n1663_), .D(new_n1500_), .Y(new_n16818_));
  NAND3X1  g16754(.A(new_n1468_), .B(new_n749_), .C(new_n364_), .Y(new_n16819_));
  OR4X1    g16755(.A(new_n16819_), .B(new_n7899_), .C(new_n7345_), .D(new_n945_), .Y(new_n16820_));
  OR4X1    g16756(.A(new_n16820_), .B(new_n16818_), .C(new_n3791_), .D(new_n894_), .Y(new_n16821_));
  NOR4X1   g16757(.A(new_n16821_), .B(new_n7749_), .C(new_n1014_), .D(new_n997_), .Y(new_n16822_));
  XOR2X1   g16758(.A(new_n16822_), .B(new_n16664_), .Y(new_n16823_));
  XOR2X1   g16759(.A(new_n16823_), .B(new_n16817_), .Y(new_n16824_));
  XOR2X1   g16760(.A(new_n16824_), .B(new_n16745_), .Y(new_n16825_));
  AOI22X1  g16761(.A0(new_n12090_), .A1(new_n1890_), .B0(new_n12088_), .B1(new_n1884_), .Y(new_n16826_));
  OAI21X1  g16762(.A0(new_n12298_), .A1(new_n3498_), .B0(new_n16826_), .Y(new_n16827_));
  AOI21X1  g16763(.A0(new_n12297_), .A1(new_n407_), .B0(new_n16827_), .Y(new_n16828_));
  XOR2X1   g16764(.A(new_n16828_), .B(new_n16825_), .Y(new_n16829_));
  AOI22X1  g16765(.A0(new_n12083_), .A1(new_n2185_), .B0(new_n12081_), .B1(new_n2095_), .Y(new_n16830_));
  OAI21X1  g16766(.A0(new_n13665_), .A1(new_n2140_), .B0(new_n16830_), .Y(new_n16831_));
  AOI21X1  g16767(.A0(new_n14672_), .A1(new_n2062_), .B0(new_n16831_), .Y(new_n16832_));
  XOR2X1   g16768(.A(new_n16832_), .B(\a[29] ), .Y(new_n16833_));
  XOR2X1   g16769(.A(new_n16833_), .B(new_n16829_), .Y(new_n16834_));
  INVX1    g16770(.A(new_n16834_), .Y(new_n16835_));
  NOR2X1   g16771(.A(new_n16750_), .B(new_n16747_), .Y(new_n16836_));
  AOI21X1  g16772(.A0(new_n16753_), .A1(new_n16751_), .B0(new_n16836_), .Y(new_n16837_));
  XOR2X1   g16773(.A(new_n16837_), .B(new_n16835_), .Y(new_n16838_));
  AOI22X1  g16774(.A0(new_n12076_), .A1(new_n2424_), .B0(new_n12018_), .B1(new_n2418_), .Y(new_n16839_));
  OAI21X1  g16775(.A0(new_n13679_), .A1(new_n2626_), .B0(new_n16839_), .Y(new_n16840_));
  AOI21X1  g16776(.A0(new_n13678_), .A1(new_n2301_), .B0(new_n16840_), .Y(new_n16841_));
  XOR2X1   g16777(.A(new_n16841_), .B(\a[26] ), .Y(new_n16842_));
  XOR2X1   g16778(.A(new_n16842_), .B(new_n16838_), .Y(new_n16843_));
  INVX1    g16779(.A(new_n16758_), .Y(new_n16844_));
  NOR2X1   g16780(.A(new_n16763_), .B(new_n16759_), .Y(new_n16845_));
  AOI21X1  g16781(.A0(new_n16844_), .A1(new_n16754_), .B0(new_n16845_), .Y(new_n16846_));
  XOR2X1   g16782(.A(new_n16846_), .B(new_n16843_), .Y(new_n16847_));
  INVX1    g16783(.A(new_n16847_), .Y(new_n16848_));
  NOR2X1   g16784(.A(new_n16768_), .B(new_n16765_), .Y(new_n16849_));
  INVX1    g16785(.A(new_n16849_), .Y(new_n16850_));
  INVX1    g16786(.A(new_n16769_), .Y(new_n16851_));
  OAI21X1  g16787(.A0(new_n16773_), .A1(new_n16851_), .B0(new_n16850_), .Y(new_n16852_));
  AOI22X1  g16788(.A0(new_n14085_), .A1(new_n2696_), .B0(new_n12285_), .B1(new_n2657_), .Y(new_n16853_));
  OAI21X1  g16789(.A0(new_n14088_), .A1(new_n2753_), .B0(new_n16853_), .Y(new_n16854_));
  AOI21X1  g16790(.A0(new_n14491_), .A1(new_n2658_), .B0(new_n16854_), .Y(new_n16855_));
  XOR2X1   g16791(.A(new_n16855_), .B(\a[23] ), .Y(new_n16856_));
  XOR2X1   g16792(.A(new_n16856_), .B(new_n16852_), .Y(new_n16857_));
  XOR2X1   g16793(.A(new_n16857_), .B(new_n16848_), .Y(new_n16858_));
  AOI22X1  g16794(.A0(new_n14642_), .A1(new_n3099_), .B0(new_n14084_), .B1(new_n2875_), .Y(new_n16859_));
  OAI21X1  g16795(.A0(new_n14805_), .A1(new_n3152_), .B0(new_n16859_), .Y(new_n16860_));
  AOI21X1  g16796(.A0(new_n14809_), .A1(new_n2876_), .B0(new_n16860_), .Y(new_n16861_));
  XOR2X1   g16797(.A(new_n16861_), .B(\a[20] ), .Y(new_n16862_));
  XOR2X1   g16798(.A(new_n16862_), .B(new_n16858_), .Y(new_n16863_));
  INVX1    g16799(.A(new_n16863_), .Y(new_n16864_));
  NOR2X1   g16800(.A(new_n16777_), .B(new_n16774_), .Y(new_n16865_));
  INVX1    g16801(.A(new_n16782_), .Y(new_n16866_));
  AOI21X1  g16802(.A0(new_n16866_), .A1(new_n16778_), .B0(new_n16865_), .Y(new_n16867_));
  XOR2X1   g16803(.A(new_n16867_), .B(new_n16864_), .Y(new_n16868_));
  NOR2X1   g16804(.A(new_n16786_), .B(new_n16783_), .Y(new_n16869_));
  INVX1    g16805(.A(new_n16869_), .Y(new_n16870_));
  INVX1    g16806(.A(new_n16787_), .Y(new_n16871_));
  OAI21X1  g16807(.A0(new_n16791_), .A1(new_n16871_), .B0(new_n16870_), .Y(new_n16872_));
  AOI22X1  g16808(.A0(new_n15087_), .A1(new_n3390_), .B0(new_n14946_), .B1(new_n3232_), .Y(new_n16873_));
  OAI21X1  g16809(.A0(new_n15363_), .A1(new_n3545_), .B0(new_n16873_), .Y(new_n16874_));
  AOI21X1  g16810(.A0(new_n15240_), .A1(new_n3234_), .B0(new_n16874_), .Y(new_n16875_));
  XOR2X1   g16811(.A(new_n16875_), .B(\a[17] ), .Y(new_n16876_));
  XOR2X1   g16812(.A(new_n16876_), .B(new_n16872_), .Y(new_n16877_));
  XOR2X1   g16813(.A(new_n16877_), .B(new_n16868_), .Y(new_n16878_));
  XOR2X1   g16814(.A(new_n16878_), .B(new_n16815_), .Y(new_n16879_));
  INVX1    g16815(.A(new_n16879_), .Y(new_n16880_));
  XOR2X1   g16816(.A(new_n16880_), .B(new_n16811_), .Y(new_n16881_));
  XOR2X1   g16817(.A(new_n16881_), .B(new_n16809_), .Y(\result[19] ));
  AND2X1   g16818(.A(new_n16881_), .B(new_n16809_), .Y(new_n16883_));
  NOR2X1   g16819(.A(new_n16833_), .B(new_n16829_), .Y(new_n16884_));
  INVX1    g16820(.A(new_n16884_), .Y(new_n16885_));
  OAI21X1  g16821(.A0(new_n16837_), .A1(new_n16835_), .B0(new_n16885_), .Y(new_n16886_));
  AOI22X1  g16822(.A0(new_n12088_), .A1(new_n1890_), .B0(new_n12085_), .B1(new_n1884_), .Y(new_n16887_));
  OAI21X1  g16823(.A0(new_n13321_), .A1(new_n3498_), .B0(new_n16887_), .Y(new_n16888_));
  AOI21X1  g16824(.A0(new_n13344_), .A1(new_n407_), .B0(new_n16888_), .Y(new_n16889_));
  NAND2X1  g16825(.A(new_n16823_), .B(new_n16817_), .Y(new_n16890_));
  OAI21X1  g16826(.A0(new_n16822_), .A1(new_n16664_), .B0(new_n16890_), .Y(new_n16891_));
  OAI22X1  g16827(.A0(new_n129_), .A1(new_n75_), .B0(new_n117_), .B1(new_n81_), .Y(new_n16892_));
  OR4X1    g16828(.A(new_n537_), .B(new_n272_), .C(new_n170_), .D(new_n93_), .Y(new_n16893_));
  OR4X1    g16829(.A(new_n421_), .B(new_n264_), .C(new_n193_), .D(new_n410_), .Y(new_n16894_));
  OR4X1    g16830(.A(new_n16894_), .B(new_n16893_), .C(new_n16892_), .D(new_n603_), .Y(new_n16895_));
  OR4X1    g16831(.A(new_n2119_), .B(new_n1547_), .C(new_n1540_), .D(new_n602_), .Y(new_n16896_));
  OR4X1    g16832(.A(new_n16896_), .B(new_n16895_), .C(new_n7919_), .D(new_n3318_), .Y(new_n16897_));
  NOR3X1   g16833(.A(new_n16897_), .B(new_n2933_), .C(new_n1716_), .Y(new_n16898_));
  XOR2X1   g16834(.A(new_n16898_), .B(new_n16891_), .Y(new_n16899_));
  XOR2X1   g16835(.A(new_n16899_), .B(new_n16889_), .Y(new_n16900_));
  INVX1    g16836(.A(new_n16900_), .Y(new_n16901_));
  INVX1    g16837(.A(new_n16825_), .Y(new_n16902_));
  NOR2X1   g16838(.A(new_n16828_), .B(new_n16902_), .Y(new_n16903_));
  AOI21X1  g16839(.A0(new_n16824_), .A1(new_n16745_), .B0(new_n16903_), .Y(new_n16904_));
  XOR2X1   g16840(.A(new_n16904_), .B(new_n16901_), .Y(new_n16905_));
  OAI22X1  g16841(.A0(new_n13320_), .A1(new_n2186_), .B0(new_n13665_), .B1(new_n2431_), .Y(new_n16906_));
  AOI21X1  g16842(.A0(new_n12076_), .A1(new_n2139_), .B0(new_n16906_), .Y(new_n16907_));
  OAI21X1  g16843(.A0(new_n13672_), .A1(new_n2063_), .B0(new_n16907_), .Y(new_n16908_));
  XOR2X1   g16844(.A(new_n16908_), .B(new_n74_), .Y(new_n16909_));
  XOR2X1   g16845(.A(new_n16909_), .B(new_n16905_), .Y(new_n16910_));
  XOR2X1   g16846(.A(new_n16910_), .B(new_n16886_), .Y(new_n16911_));
  AOI22X1  g16847(.A0(new_n12074_), .A1(new_n2418_), .B0(new_n12018_), .B1(new_n2424_), .Y(new_n16912_));
  OAI21X1  g16848(.A0(new_n12292_), .A1(new_n2626_), .B0(new_n16912_), .Y(new_n16913_));
  AOI21X1  g16849(.A0(new_n12291_), .A1(new_n2301_), .B0(new_n16913_), .Y(new_n16914_));
  XOR2X1   g16850(.A(new_n16914_), .B(\a[26] ), .Y(new_n16915_));
  XOR2X1   g16851(.A(new_n16915_), .B(new_n16911_), .Y(new_n16916_));
  INVX1    g16852(.A(new_n16842_), .Y(new_n16917_));
  NOR2X1   g16853(.A(new_n16846_), .B(new_n16843_), .Y(new_n16918_));
  AOI21X1  g16854(.A0(new_n16917_), .A1(new_n16838_), .B0(new_n16918_), .Y(new_n16919_));
  XOR2X1   g16855(.A(new_n16919_), .B(new_n16916_), .Y(new_n16920_));
  AOI22X1  g16856(.A0(new_n14087_), .A1(new_n2696_), .B0(new_n14085_), .B1(new_n2657_), .Y(new_n16921_));
  OAI21X1  g16857(.A0(new_n14643_), .A1(new_n2753_), .B0(new_n16921_), .Y(new_n16922_));
  AOI21X1  g16858(.A0(new_n14106_), .A1(new_n2658_), .B0(new_n16922_), .Y(new_n16923_));
  XOR2X1   g16859(.A(new_n16923_), .B(\a[23] ), .Y(new_n16924_));
  XOR2X1   g16860(.A(new_n16924_), .B(new_n16920_), .Y(new_n16925_));
  INVX1    g16861(.A(new_n16856_), .Y(new_n16926_));
  NOR2X1   g16862(.A(new_n16857_), .B(new_n16848_), .Y(new_n16927_));
  AOI21X1  g16863(.A0(new_n16926_), .A1(new_n16852_), .B0(new_n16927_), .Y(new_n16928_));
  XOR2X1   g16864(.A(new_n16928_), .B(new_n16925_), .Y(new_n16929_));
  AOI22X1  g16865(.A0(new_n14804_), .A1(new_n3099_), .B0(new_n14642_), .B1(new_n2875_), .Y(new_n16930_));
  OAI21X1  g16866(.A0(new_n15088_), .A1(new_n3152_), .B0(new_n16930_), .Y(new_n16931_));
  AOI21X1  g16867(.A0(new_n14952_), .A1(new_n2876_), .B0(new_n16931_), .Y(new_n16932_));
  XOR2X1   g16868(.A(new_n16932_), .B(\a[20] ), .Y(new_n16933_));
  XOR2X1   g16869(.A(new_n16933_), .B(new_n16929_), .Y(new_n16934_));
  INVX1    g16870(.A(new_n16862_), .Y(new_n16935_));
  NOR2X1   g16871(.A(new_n16867_), .B(new_n16863_), .Y(new_n16936_));
  AOI21X1  g16872(.A0(new_n16935_), .A1(new_n16858_), .B0(new_n16936_), .Y(new_n16937_));
  XOR2X1   g16873(.A(new_n16937_), .B(new_n16934_), .Y(new_n16938_));
  AOI22X1  g16874(.A0(new_n15234_), .A1(new_n3390_), .B0(new_n15087_), .B1(new_n3232_), .Y(new_n16939_));
  OAI21X1  g16875(.A0(new_n15522_), .A1(new_n3545_), .B0(new_n16939_), .Y(new_n16940_));
  AOI21X1  g16876(.A0(new_n15841_), .A1(new_n3234_), .B0(new_n16940_), .Y(new_n16941_));
  XOR2X1   g16877(.A(new_n16941_), .B(\a[17] ), .Y(new_n16942_));
  XOR2X1   g16878(.A(new_n16942_), .B(new_n16938_), .Y(new_n16943_));
  INVX1    g16879(.A(new_n16876_), .Y(new_n16944_));
  NOR2X1   g16880(.A(new_n16877_), .B(new_n16868_), .Y(new_n16945_));
  AOI21X1  g16881(.A0(new_n16944_), .A1(new_n16872_), .B0(new_n16945_), .Y(new_n16946_));
  XOR2X1   g16882(.A(new_n16946_), .B(new_n16943_), .Y(new_n16947_));
  INVX1    g16883(.A(new_n16947_), .Y(new_n16948_));
  INVX1    g16884(.A(new_n16810_), .Y(new_n16949_));
  INVX1    g16885(.A(new_n16803_), .Y(new_n16950_));
  NOR2X1   g16886(.A(new_n16722_), .B(new_n16804_), .Y(new_n16951_));
  XOR2X1   g16887(.A(new_n16722_), .B(new_n16804_), .Y(new_n16952_));
  OR2X1    g16888(.A(new_n16448_), .B(new_n16555_), .Y(new_n16953_));
  OAI21X1  g16889(.A0(new_n16466_), .A1(new_n16449_), .B0(new_n16953_), .Y(new_n16954_));
  AOI21X1  g16890(.A0(new_n16954_), .A1(new_n16553_), .B0(new_n16565_), .Y(new_n16955_));
  NAND2X1  g16891(.A(new_n16646_), .B(new_n16571_), .Y(new_n16956_));
  NOR2X1   g16892(.A(new_n16646_), .B(new_n16571_), .Y(new_n16957_));
  OAI21X1  g16893(.A0(new_n16957_), .A1(new_n16955_), .B0(new_n16956_), .Y(new_n16958_));
  AOI21X1  g16894(.A0(new_n16958_), .A1(new_n16952_), .B0(new_n16951_), .Y(new_n16959_));
  OAI21X1  g16895(.A0(new_n16959_), .A1(new_n16950_), .B0(new_n16949_), .Y(new_n16960_));
  AND2X1   g16896(.A(new_n16878_), .B(new_n16815_), .Y(new_n16961_));
  AOI21X1  g16897(.A0(new_n16879_), .A1(new_n16960_), .B0(new_n16961_), .Y(new_n16962_));
  XOR2X1   g16898(.A(new_n16962_), .B(new_n16948_), .Y(new_n16963_));
  XOR2X1   g16899(.A(new_n16963_), .B(new_n16883_), .Y(\result[20] ));
  NOR2X1   g16900(.A(new_n16904_), .B(new_n16900_), .Y(new_n16965_));
  NOR2X1   g16901(.A(new_n16909_), .B(new_n16905_), .Y(new_n16966_));
  NOR2X1   g16902(.A(new_n16966_), .B(new_n16965_), .Y(new_n16967_));
  INVX1    g16903(.A(new_n16967_), .Y(new_n16968_));
  OR2X1    g16904(.A(new_n3017_), .B(new_n2586_), .Y(new_n16969_));
  INVX1    g16905(.A(new_n1632_), .Y(new_n16970_));
  OAI22X1  g16906(.A0(new_n152_), .A1(new_n129_), .B0(new_n99_), .B1(new_n75_), .Y(new_n16971_));
  OR4X1    g16907(.A(new_n468_), .B(new_n819_), .C(new_n183_), .D(new_n1284_), .Y(new_n16972_));
  OR4X1    g16908(.A(new_n1028_), .B(new_n286_), .C(new_n142_), .D(new_n884_), .Y(new_n16973_));
  OR4X1    g16909(.A(new_n16973_), .B(new_n16972_), .C(new_n16971_), .D(new_n450_), .Y(new_n16974_));
  OR4X1    g16910(.A(new_n1850_), .B(new_n1417_), .C(new_n1336_), .D(new_n1100_), .Y(new_n16975_));
  OR4X1    g16911(.A(new_n16975_), .B(new_n16974_), .C(new_n2259_), .D(new_n16970_), .Y(new_n16976_));
  NOR4X1   g16912(.A(new_n16976_), .B(new_n7196_), .C(new_n16969_), .D(new_n942_), .Y(new_n16977_));
  NOR4X1   g16913(.A(new_n16977_), .B(new_n16897_), .C(new_n2933_), .D(new_n1716_), .Y(new_n16978_));
  INVX1    g16914(.A(new_n16889_), .Y(new_n16979_));
  AND2X1   g16915(.A(new_n16898_), .B(new_n16891_), .Y(new_n16980_));
  AOI21X1  g16916(.A0(new_n16899_), .A1(new_n16979_), .B0(new_n16980_), .Y(new_n16981_));
  OR2X1    g16917(.A(new_n16969_), .B(new_n942_), .Y(new_n16982_));
  NOR4X1   g16918(.A(new_n16982_), .B(new_n16976_), .C(new_n16898_), .D(new_n7196_), .Y(new_n16983_));
  NOR3X1   g16919(.A(new_n16983_), .B(new_n16978_), .C(new_n16981_), .Y(new_n16984_));
  OR2X1    g16920(.A(new_n16984_), .B(new_n16981_), .Y(new_n16985_));
  NOR2X1   g16921(.A(new_n16984_), .B(new_n16983_), .Y(new_n16986_));
  INVX1    g16922(.A(new_n16986_), .Y(new_n16987_));
  OAI21X1  g16923(.A0(new_n16987_), .A1(new_n16978_), .B0(new_n16985_), .Y(new_n16988_));
  AOI22X1  g16924(.A0(new_n12085_), .A1(new_n1890_), .B0(new_n12083_), .B1(new_n1884_), .Y(new_n16989_));
  OAI21X1  g16925(.A0(new_n13320_), .A1(new_n3498_), .B0(new_n16989_), .Y(new_n16990_));
  AOI21X1  g16926(.A0(new_n14510_), .A1(new_n407_), .B0(new_n16990_), .Y(new_n16991_));
  XOR2X1   g16927(.A(new_n16991_), .B(new_n16988_), .Y(new_n16992_));
  OAI22X1  g16928(.A0(new_n13665_), .A1(new_n2186_), .B0(new_n13700_), .B1(new_n2431_), .Y(new_n16993_));
  AOI21X1  g16929(.A0(new_n12018_), .A1(new_n2139_), .B0(new_n16993_), .Y(new_n16994_));
  OAI21X1  g16930(.A0(new_n14604_), .A1(new_n2063_), .B0(new_n16994_), .Y(new_n16995_));
  XOR2X1   g16931(.A(new_n16995_), .B(new_n74_), .Y(new_n16996_));
  XOR2X1   g16932(.A(new_n16996_), .B(new_n16992_), .Y(new_n16997_));
  XOR2X1   g16933(.A(new_n16997_), .B(new_n16968_), .Y(new_n16998_));
  AOI22X1  g16934(.A0(new_n12285_), .A1(new_n2418_), .B0(new_n12074_), .B1(new_n2424_), .Y(new_n16999_));
  OAI21X1  g16935(.A0(new_n14086_), .A1(new_n2626_), .B0(new_n16999_), .Y(new_n17000_));
  AOI21X1  g16936(.A0(new_n14480_), .A1(new_n2301_), .B0(new_n17000_), .Y(new_n17001_));
  XOR2X1   g16937(.A(new_n17001_), .B(\a[26] ), .Y(new_n17002_));
  XOR2X1   g16938(.A(new_n17002_), .B(new_n16998_), .Y(new_n17003_));
  AND2X1   g16939(.A(new_n16910_), .B(new_n16886_), .Y(new_n17004_));
  INVX1    g16940(.A(new_n16915_), .Y(new_n17005_));
  AOI21X1  g16941(.A0(new_n17005_), .A1(new_n16911_), .B0(new_n17004_), .Y(new_n17006_));
  XOR2X1   g16942(.A(new_n17006_), .B(new_n17003_), .Y(new_n17007_));
  AOI22X1  g16943(.A0(new_n14087_), .A1(new_n2657_), .B0(new_n14084_), .B1(new_n2696_), .Y(new_n17008_));
  OAI21X1  g16944(.A0(new_n14648_), .A1(new_n2753_), .B0(new_n17008_), .Y(new_n17009_));
  AOI21X1  g16945(.A0(new_n14651_), .A1(new_n2658_), .B0(new_n17009_), .Y(new_n17010_));
  XOR2X1   g16946(.A(new_n17010_), .B(\a[23] ), .Y(new_n17011_));
  XOR2X1   g16947(.A(new_n17011_), .B(new_n17007_), .Y(new_n17012_));
  NOR2X1   g16948(.A(new_n16919_), .B(new_n16916_), .Y(new_n17013_));
  INVX1    g16949(.A(new_n16924_), .Y(new_n17014_));
  AOI21X1  g16950(.A0(new_n17014_), .A1(new_n16920_), .B0(new_n17013_), .Y(new_n17015_));
  XOR2X1   g16951(.A(new_n17015_), .B(new_n17012_), .Y(new_n17016_));
  AOI22X1  g16952(.A0(new_n14946_), .A1(new_n3099_), .B0(new_n14804_), .B1(new_n2875_), .Y(new_n17017_));
  OAI21X1  g16953(.A0(new_n15235_), .A1(new_n3152_), .B0(new_n17017_), .Y(new_n17018_));
  AOI21X1  g16954(.A0(new_n15381_), .A1(new_n2876_), .B0(new_n17018_), .Y(new_n17019_));
  XOR2X1   g16955(.A(new_n17019_), .B(\a[20] ), .Y(new_n17020_));
  XOR2X1   g16956(.A(new_n17020_), .B(new_n17016_), .Y(new_n17021_));
  NOR2X1   g16957(.A(new_n16928_), .B(new_n16925_), .Y(new_n17022_));
  INVX1    g16958(.A(new_n16933_), .Y(new_n17023_));
  AOI21X1  g16959(.A0(new_n17023_), .A1(new_n16929_), .B0(new_n17022_), .Y(new_n17024_));
  AOI22X1  g16960(.A0(new_n15362_), .A1(new_n8123_), .B0(new_n15234_), .B1(new_n3232_), .Y(new_n17025_));
  OAI21X1  g16961(.A0(new_n15373_), .A1(new_n3388_), .B0(new_n17025_), .Y(new_n17026_));
  XOR2X1   g16962(.A(new_n17026_), .B(new_n2445_), .Y(new_n17027_));
  XOR2X1   g16963(.A(new_n17027_), .B(new_n17024_), .Y(new_n17028_));
  XOR2X1   g16964(.A(new_n17028_), .B(new_n17021_), .Y(new_n17029_));
  NOR2X1   g16965(.A(new_n16937_), .B(new_n16934_), .Y(new_n17030_));
  INVX1    g16966(.A(new_n16942_), .Y(new_n17031_));
  AOI21X1  g16967(.A0(new_n17031_), .A1(new_n16938_), .B0(new_n17030_), .Y(new_n17032_));
  XOR2X1   g16968(.A(new_n17032_), .B(new_n17029_), .Y(new_n17033_));
  INVX1    g16969(.A(new_n17033_), .Y(new_n17034_));
  NOR2X1   g16970(.A(new_n16946_), .B(new_n16943_), .Y(new_n17035_));
  INVX1    g16971(.A(new_n16961_), .Y(new_n17036_));
  OAI21X1  g16972(.A0(new_n16880_), .A1(new_n16811_), .B0(new_n17036_), .Y(new_n17037_));
  AOI21X1  g16973(.A0(new_n17037_), .A1(new_n16947_), .B0(new_n17035_), .Y(new_n17038_));
  XOR2X1   g16974(.A(new_n17038_), .B(new_n17034_), .Y(new_n17039_));
  AND2X1   g16975(.A(new_n16963_), .B(new_n16883_), .Y(new_n17040_));
  XOR2X1   g16976(.A(new_n17040_), .B(new_n17039_), .Y(\result[21] ));
  AND2X1   g16977(.A(new_n17040_), .B(new_n17039_), .Y(new_n17042_));
  NOR2X1   g16978(.A(new_n17032_), .B(new_n17029_), .Y(new_n17043_));
  INVX1    g16979(.A(new_n17043_), .Y(new_n17044_));
  OAI21X1  g16980(.A0(new_n17038_), .A1(new_n17034_), .B0(new_n17044_), .Y(new_n17045_));
  INVX1    g16981(.A(new_n17021_), .Y(new_n17046_));
  NOR2X1   g16982(.A(new_n17027_), .B(new_n17024_), .Y(new_n17047_));
  AOI21X1  g16983(.A0(new_n17028_), .A1(new_n17046_), .B0(new_n17047_), .Y(new_n17048_));
  INVX1    g16984(.A(new_n17048_), .Y(new_n17049_));
  NOR2X1   g16985(.A(new_n17006_), .B(new_n17003_), .Y(new_n17050_));
  INVX1    g16986(.A(new_n17050_), .Y(new_n17051_));
  INVX1    g16987(.A(new_n17007_), .Y(new_n17052_));
  OAI21X1  g16988(.A0(new_n17011_), .A1(new_n17052_), .B0(new_n17051_), .Y(new_n17053_));
  INVX1    g16989(.A(new_n17053_), .Y(new_n17054_));
  AND2X1   g16990(.A(new_n16997_), .B(new_n16968_), .Y(new_n17055_));
  INVX1    g16991(.A(new_n17002_), .Y(new_n17056_));
  AOI21X1  g16992(.A0(new_n17056_), .A1(new_n16998_), .B0(new_n17055_), .Y(new_n17057_));
  AOI22X1  g16993(.A0(new_n14085_), .A1(new_n2418_), .B0(new_n12285_), .B1(new_n2424_), .Y(new_n17058_));
  OAI21X1  g16994(.A0(new_n14088_), .A1(new_n2626_), .B0(new_n17058_), .Y(new_n17059_));
  AOI21X1  g16995(.A0(new_n14491_), .A1(new_n2301_), .B0(new_n17059_), .Y(new_n17060_));
  XOR2X1   g16996(.A(new_n17060_), .B(\a[26] ), .Y(new_n17061_));
  XOR2X1   g16997(.A(new_n17061_), .B(new_n17057_), .Y(new_n17062_));
  OR2X1    g16998(.A(new_n16987_), .B(new_n16978_), .Y(new_n17063_));
  AOI21X1  g16999(.A0(new_n17063_), .A1(new_n16985_), .B0(new_n16991_), .Y(new_n17064_));
  NOR2X1   g17000(.A(new_n16996_), .B(new_n16992_), .Y(new_n17065_));
  NOR2X1   g17001(.A(new_n17065_), .B(new_n17064_), .Y(new_n17066_));
  AND2X1   g17002(.A(new_n15362_), .B(new_n7394_), .Y(new_n17067_));
  XOR2X1   g17003(.A(new_n17067_), .B(new_n2445_), .Y(new_n17068_));
  OR4X1    g17004(.A(new_n497_), .B(new_n496_), .C(new_n399_), .D(new_n142_), .Y(new_n17069_));
  NOR4X1   g17005(.A(new_n17069_), .B(new_n612_), .C(new_n819_), .D(new_n139_), .Y(new_n17070_));
  NAND3X1  g17006(.A(new_n17070_), .B(new_n13051_), .C(new_n948_), .Y(new_n17071_));
  OR4X1    g17007(.A(new_n17071_), .B(new_n1722_), .C(new_n828_), .D(new_n205_), .Y(new_n17072_));
  NOR4X1   g17008(.A(new_n17072_), .B(new_n2804_), .C(new_n2026_), .D(new_n534_), .Y(new_n17073_));
  XOR2X1   g17009(.A(new_n17073_), .B(new_n16977_), .Y(new_n17074_));
  XOR2X1   g17010(.A(new_n17074_), .B(new_n17068_), .Y(new_n17075_));
  AOI22X1  g17011(.A0(new_n12083_), .A1(new_n1890_), .B0(new_n12081_), .B1(new_n1884_), .Y(new_n17076_));
  OAI21X1  g17012(.A0(new_n13665_), .A1(new_n3498_), .B0(new_n17076_), .Y(new_n17077_));
  AOI21X1  g17013(.A0(new_n14672_), .A1(new_n407_), .B0(new_n17077_), .Y(new_n17078_));
  XOR2X1   g17014(.A(new_n17078_), .B(new_n17075_), .Y(new_n17079_));
  XOR2X1   g17015(.A(new_n17079_), .B(new_n16987_), .Y(new_n17080_));
  XOR2X1   g17016(.A(new_n17080_), .B(new_n17066_), .Y(new_n17081_));
  AOI22X1  g17017(.A0(new_n12076_), .A1(new_n2185_), .B0(new_n12018_), .B1(new_n2095_), .Y(new_n17082_));
  OAI21X1  g17018(.A0(new_n13679_), .A1(new_n2140_), .B0(new_n17082_), .Y(new_n17083_));
  AOI21X1  g17019(.A0(new_n13678_), .A1(new_n2062_), .B0(new_n17083_), .Y(new_n17084_));
  XOR2X1   g17020(.A(new_n17084_), .B(\a[29] ), .Y(new_n17085_));
  XOR2X1   g17021(.A(new_n17085_), .B(new_n17081_), .Y(new_n17086_));
  XOR2X1   g17022(.A(new_n17086_), .B(new_n17062_), .Y(new_n17087_));
  AOI22X1  g17023(.A0(new_n14642_), .A1(new_n2696_), .B0(new_n14084_), .B1(new_n2657_), .Y(new_n17088_));
  OAI21X1  g17024(.A0(new_n14805_), .A1(new_n2753_), .B0(new_n17088_), .Y(new_n17089_));
  AOI21X1  g17025(.A0(new_n14809_), .A1(new_n2658_), .B0(new_n17089_), .Y(new_n17090_));
  XOR2X1   g17026(.A(new_n17090_), .B(\a[23] ), .Y(new_n17091_));
  XOR2X1   g17027(.A(new_n17091_), .B(new_n17087_), .Y(new_n17092_));
  XOR2X1   g17028(.A(new_n17092_), .B(new_n17054_), .Y(new_n17093_));
  NOR2X1   g17029(.A(new_n17015_), .B(new_n17012_), .Y(new_n17094_));
  INVX1    g17030(.A(new_n17094_), .Y(new_n17095_));
  INVX1    g17031(.A(new_n17016_), .Y(new_n17096_));
  OAI21X1  g17032(.A0(new_n17020_), .A1(new_n17096_), .B0(new_n17095_), .Y(new_n17097_));
  AOI22X1  g17033(.A0(new_n15087_), .A1(new_n3099_), .B0(new_n14946_), .B1(new_n2875_), .Y(new_n17098_));
  OAI21X1  g17034(.A0(new_n15363_), .A1(new_n3152_), .B0(new_n17098_), .Y(new_n17099_));
  AOI21X1  g17035(.A0(new_n15240_), .A1(new_n2876_), .B0(new_n17099_), .Y(new_n17100_));
  XOR2X1   g17036(.A(new_n17100_), .B(\a[20] ), .Y(new_n17101_));
  XOR2X1   g17037(.A(new_n17101_), .B(new_n17097_), .Y(new_n17102_));
  XOR2X1   g17038(.A(new_n17102_), .B(new_n17093_), .Y(new_n17103_));
  XOR2X1   g17039(.A(new_n17103_), .B(new_n17049_), .Y(new_n17104_));
  XOR2X1   g17040(.A(new_n17104_), .B(new_n17045_), .Y(new_n17105_));
  XOR2X1   g17041(.A(new_n17105_), .B(new_n17042_), .Y(\result[22] ));
  AND2X1   g17042(.A(new_n17105_), .B(new_n17042_), .Y(new_n17107_));
  NOR2X1   g17043(.A(new_n17080_), .B(new_n17066_), .Y(new_n17108_));
  INVX1    g17044(.A(new_n17108_), .Y(new_n17109_));
  INVX1    g17045(.A(new_n17081_), .Y(new_n17110_));
  OAI21X1  g17046(.A0(new_n17085_), .A1(new_n17110_), .B0(new_n17109_), .Y(new_n17111_));
  AOI21X1  g17047(.A0(new_n13671_), .A1(new_n13669_), .B0(new_n3178_), .Y(new_n17112_));
  AOI22X1  g17048(.A0(new_n12081_), .A1(new_n1890_), .B0(new_n12079_), .B1(new_n1884_), .Y(new_n17113_));
  OAI21X1  g17049(.A0(new_n13700_), .A1(new_n3498_), .B0(new_n17113_), .Y(new_n17114_));
  NOR2X1   g17050(.A(new_n17114_), .B(new_n17112_), .Y(new_n17115_));
  NAND2X1  g17051(.A(new_n17074_), .B(new_n17068_), .Y(new_n17116_));
  OAI21X1  g17052(.A0(new_n17073_), .A1(new_n16977_), .B0(new_n17116_), .Y(new_n17117_));
  OR4X1    g17053(.A(new_n740_), .B(new_n418_), .C(new_n319_), .D(new_n137_), .Y(new_n17118_));
  OR4X1    g17054(.A(new_n354_), .B(new_n220_), .C(new_n149_), .D(new_n103_), .Y(new_n17119_));
  OR4X1    g17055(.A(new_n17119_), .B(new_n17118_), .C(new_n7063_), .D(new_n1697_), .Y(new_n17120_));
  OR4X1    g17056(.A(new_n17120_), .B(new_n2451_), .C(new_n653_), .D(new_n561_), .Y(new_n17121_));
  OR2X1    g17057(.A(new_n2147_), .B(new_n1668_), .Y(new_n17122_));
  NOR4X1   g17058(.A(new_n17122_), .B(new_n17121_), .C(new_n16176_), .D(new_n3695_), .Y(new_n17123_));
  XOR2X1   g17059(.A(new_n17123_), .B(new_n17117_), .Y(new_n17124_));
  XOR2X1   g17060(.A(new_n17124_), .B(new_n17115_), .Y(new_n17125_));
  INVX1    g17061(.A(new_n17125_), .Y(new_n17126_));
  INVX1    g17062(.A(new_n17075_), .Y(new_n17127_));
  NOR2X1   g17063(.A(new_n17078_), .B(new_n17127_), .Y(new_n17128_));
  NOR2X1   g17064(.A(new_n17079_), .B(new_n16986_), .Y(new_n17129_));
  NOR2X1   g17065(.A(new_n17129_), .B(new_n17128_), .Y(new_n17130_));
  XOR2X1   g17066(.A(new_n17130_), .B(new_n17126_), .Y(new_n17131_));
  OAI22X1  g17067(.A0(new_n13679_), .A1(new_n2431_), .B0(new_n13691_), .B1(new_n2186_), .Y(new_n17132_));
  AOI21X1  g17068(.A0(new_n12285_), .A1(new_n2139_), .B0(new_n17132_), .Y(new_n17133_));
  OAI21X1  g17069(.A0(new_n14467_), .A1(new_n2063_), .B0(new_n17133_), .Y(new_n17134_));
  XOR2X1   g17070(.A(new_n17134_), .B(new_n74_), .Y(new_n17135_));
  XOR2X1   g17071(.A(new_n17135_), .B(new_n17131_), .Y(new_n17136_));
  XOR2X1   g17072(.A(new_n17136_), .B(new_n17111_), .Y(new_n17137_));
  AOI22X1  g17073(.A0(new_n14087_), .A1(new_n2418_), .B0(new_n14085_), .B1(new_n2424_), .Y(new_n17138_));
  OAI21X1  g17074(.A0(new_n14643_), .A1(new_n2626_), .B0(new_n17138_), .Y(new_n17139_));
  AOI21X1  g17075(.A0(new_n14106_), .A1(new_n2301_), .B0(new_n17139_), .Y(new_n17140_));
  XOR2X1   g17076(.A(new_n17140_), .B(\a[26] ), .Y(new_n17141_));
  XOR2X1   g17077(.A(new_n17141_), .B(new_n17137_), .Y(new_n17142_));
  NOR2X1   g17078(.A(new_n17061_), .B(new_n17057_), .Y(new_n17143_));
  INVX1    g17079(.A(new_n17086_), .Y(new_n17144_));
  AOI21X1  g17080(.A0(new_n17144_), .A1(new_n17062_), .B0(new_n17143_), .Y(new_n17145_));
  XOR2X1   g17081(.A(new_n17145_), .B(new_n17142_), .Y(new_n17146_));
  AOI22X1  g17082(.A0(new_n14804_), .A1(new_n2696_), .B0(new_n14642_), .B1(new_n2657_), .Y(new_n17147_));
  OAI21X1  g17083(.A0(new_n15088_), .A1(new_n2753_), .B0(new_n17147_), .Y(new_n17148_));
  AOI21X1  g17084(.A0(new_n14952_), .A1(new_n2658_), .B0(new_n17148_), .Y(new_n17149_));
  XOR2X1   g17085(.A(new_n17149_), .B(\a[23] ), .Y(new_n17150_));
  XOR2X1   g17086(.A(new_n17150_), .B(new_n17146_), .Y(new_n17151_));
  NOR2X1   g17087(.A(new_n17091_), .B(new_n17087_), .Y(new_n17152_));
  AOI21X1  g17088(.A0(new_n17092_), .A1(new_n17053_), .B0(new_n17152_), .Y(new_n17153_));
  XOR2X1   g17089(.A(new_n17153_), .B(new_n17151_), .Y(new_n17154_));
  AOI22X1  g17090(.A0(new_n15234_), .A1(new_n3099_), .B0(new_n15087_), .B1(new_n2875_), .Y(new_n17155_));
  OAI21X1  g17091(.A0(new_n15522_), .A1(new_n3152_), .B0(new_n17155_), .Y(new_n17156_));
  AOI21X1  g17092(.A0(new_n15841_), .A1(new_n2876_), .B0(new_n17156_), .Y(new_n17157_));
  XOR2X1   g17093(.A(new_n17157_), .B(\a[20] ), .Y(new_n17158_));
  XOR2X1   g17094(.A(new_n17158_), .B(new_n17154_), .Y(new_n17159_));
  INVX1    g17095(.A(new_n17101_), .Y(new_n17160_));
  NOR2X1   g17096(.A(new_n17102_), .B(new_n17093_), .Y(new_n17161_));
  AOI21X1  g17097(.A0(new_n17160_), .A1(new_n17097_), .B0(new_n17161_), .Y(new_n17162_));
  XOR2X1   g17098(.A(new_n17162_), .B(new_n17159_), .Y(new_n17163_));
  INVX1    g17099(.A(new_n17163_), .Y(new_n17164_));
  AND2X1   g17100(.A(new_n17103_), .B(new_n17049_), .Y(new_n17165_));
  AOI21X1  g17101(.A0(new_n17104_), .A1(new_n17045_), .B0(new_n17165_), .Y(new_n17166_));
  XOR2X1   g17102(.A(new_n17166_), .B(new_n17164_), .Y(new_n17167_));
  XOR2X1   g17103(.A(new_n17167_), .B(new_n17107_), .Y(\result[23] ));
  AND2X1   g17104(.A(new_n17167_), .B(new_n17107_), .Y(new_n17169_));
  AOI22X1  g17105(.A0(new_n12079_), .A1(new_n1890_), .B0(new_n12076_), .B1(new_n1884_), .Y(new_n17170_));
  OAI21X1  g17106(.A0(new_n13691_), .A1(new_n3498_), .B0(new_n17170_), .Y(new_n17171_));
  AOI21X1  g17107(.A0(new_n13690_), .A1(new_n407_), .B0(new_n17171_), .Y(new_n17172_));
  INVX1    g17108(.A(new_n17123_), .Y(new_n17173_));
  OR4X1    g17109(.A(new_n1701_), .B(new_n998_), .C(new_n478_), .D(new_n254_), .Y(new_n17174_));
  OR4X1    g17110(.A(new_n869_), .B(new_n681_), .C(new_n226_), .D(new_n431_), .Y(new_n17175_));
  NOR4X1   g17111(.A(new_n17175_), .B(new_n17174_), .C(new_n16972_), .D(new_n15516_), .Y(new_n17176_));
  NAND3X1  g17112(.A(new_n17176_), .B(new_n15703_), .C(new_n2022_), .Y(new_n17177_));
  NOR4X1   g17113(.A(new_n17177_), .B(new_n3717_), .C(new_n2583_), .D(new_n564_), .Y(new_n17178_));
  AND2X1   g17114(.A(new_n17178_), .B(new_n17173_), .Y(new_n17179_));
  NOR2X1   g17115(.A(new_n17178_), .B(new_n17173_), .Y(new_n17180_));
  NOR3X1   g17116(.A(new_n17180_), .B(new_n17179_), .C(new_n17172_), .Y(new_n17181_));
  NOR2X1   g17117(.A(new_n17181_), .B(new_n17180_), .Y(new_n17182_));
  INVX1    g17118(.A(new_n17182_), .Y(new_n17183_));
  OAI22X1  g17119(.A0(new_n17183_), .A1(new_n17179_), .B0(new_n17181_), .B1(new_n17172_), .Y(new_n17184_));
  INVX1    g17120(.A(new_n17184_), .Y(new_n17185_));
  INVX1    g17121(.A(new_n17115_), .Y(new_n17186_));
  AND2X1   g17122(.A(new_n17123_), .B(new_n17117_), .Y(new_n17187_));
  AOI21X1  g17123(.A0(new_n17124_), .A1(new_n17186_), .B0(new_n17187_), .Y(new_n17188_));
  XOR2X1   g17124(.A(new_n17188_), .B(new_n17185_), .Y(new_n17189_));
  OAI21X1  g17125(.A0(new_n17129_), .A1(new_n17128_), .B0(new_n17126_), .Y(new_n17190_));
  OAI21X1  g17126(.A0(new_n17135_), .A1(new_n17131_), .B0(new_n17190_), .Y(new_n17191_));
  XOR2X1   g17127(.A(new_n17191_), .B(new_n17189_), .Y(new_n17192_));
  AOI22X1  g17128(.A0(new_n12285_), .A1(new_n2095_), .B0(new_n12074_), .B1(new_n2185_), .Y(new_n17193_));
  OAI21X1  g17129(.A0(new_n14086_), .A1(new_n2140_), .B0(new_n17193_), .Y(new_n17194_));
  AOI21X1  g17130(.A0(new_n14480_), .A1(new_n2062_), .B0(new_n17194_), .Y(new_n17195_));
  XOR2X1   g17131(.A(new_n17195_), .B(\a[29] ), .Y(new_n17196_));
  XOR2X1   g17132(.A(new_n17196_), .B(new_n17192_), .Y(new_n17197_));
  AOI22X1  g17133(.A0(new_n14087_), .A1(new_n2424_), .B0(new_n14084_), .B1(new_n2418_), .Y(new_n17198_));
  OAI21X1  g17134(.A0(new_n14648_), .A1(new_n2626_), .B0(new_n17198_), .Y(new_n17199_));
  AOI21X1  g17135(.A0(new_n14651_), .A1(new_n2301_), .B0(new_n17199_), .Y(new_n17200_));
  XOR2X1   g17136(.A(new_n17200_), .B(\a[26] ), .Y(new_n17201_));
  XOR2X1   g17137(.A(new_n17201_), .B(new_n17197_), .Y(new_n17202_));
  INVX1    g17138(.A(new_n17202_), .Y(new_n17203_));
  AND2X1   g17139(.A(new_n17136_), .B(new_n17111_), .Y(new_n17204_));
  INVX1    g17140(.A(new_n17141_), .Y(new_n17205_));
  AOI21X1  g17141(.A0(new_n17205_), .A1(new_n17137_), .B0(new_n17204_), .Y(new_n17206_));
  XOR2X1   g17142(.A(new_n17206_), .B(new_n17203_), .Y(new_n17207_));
  AOI22X1  g17143(.A0(new_n14946_), .A1(new_n2696_), .B0(new_n14804_), .B1(new_n2657_), .Y(new_n17208_));
  OAI21X1  g17144(.A0(new_n15235_), .A1(new_n2753_), .B0(new_n17208_), .Y(new_n17209_));
  AOI21X1  g17145(.A0(new_n15381_), .A1(new_n2658_), .B0(new_n17209_), .Y(new_n17210_));
  XOR2X1   g17146(.A(new_n17210_), .B(\a[23] ), .Y(new_n17211_));
  XOR2X1   g17147(.A(new_n17211_), .B(new_n17207_), .Y(new_n17212_));
  NOR2X1   g17148(.A(new_n17145_), .B(new_n17142_), .Y(new_n17213_));
  INVX1    g17149(.A(new_n17150_), .Y(new_n17214_));
  AOI21X1  g17150(.A0(new_n17214_), .A1(new_n17146_), .B0(new_n17213_), .Y(new_n17215_));
  AOI22X1  g17151(.A0(new_n15362_), .A1(new_n7805_), .B0(new_n15234_), .B1(new_n2875_), .Y(new_n17216_));
  OAI21X1  g17152(.A0(new_n15373_), .A1(new_n3098_), .B0(new_n17216_), .Y(new_n17217_));
  XOR2X1   g17153(.A(new_n17217_), .B(new_n1920_), .Y(new_n17218_));
  XOR2X1   g17154(.A(new_n17218_), .B(new_n17215_), .Y(new_n17219_));
  XOR2X1   g17155(.A(new_n17219_), .B(new_n17212_), .Y(new_n17220_));
  NOR2X1   g17156(.A(new_n17153_), .B(new_n17151_), .Y(new_n17221_));
  INVX1    g17157(.A(new_n17158_), .Y(new_n17222_));
  AOI21X1  g17158(.A0(new_n17222_), .A1(new_n17154_), .B0(new_n17221_), .Y(new_n17223_));
  XOR2X1   g17159(.A(new_n17223_), .B(new_n17220_), .Y(new_n17224_));
  NOR2X1   g17160(.A(new_n17162_), .B(new_n17159_), .Y(new_n17225_));
  INVX1    g17161(.A(new_n17225_), .Y(new_n17226_));
  OAI21X1  g17162(.A0(new_n17166_), .A1(new_n17164_), .B0(new_n17226_), .Y(new_n17227_));
  XOR2X1   g17163(.A(new_n17227_), .B(new_n17224_), .Y(new_n17228_));
  XOR2X1   g17164(.A(new_n17228_), .B(new_n17169_), .Y(\result[24] ));
  AND2X1   g17165(.A(new_n17228_), .B(new_n17169_), .Y(new_n17230_));
  NOR2X1   g17166(.A(new_n17223_), .B(new_n17220_), .Y(new_n17231_));
  INVX1    g17167(.A(new_n17231_), .Y(new_n17232_));
  INVX1    g17168(.A(new_n17224_), .Y(new_n17233_));
  INVX1    g17169(.A(new_n17035_), .Y(new_n17234_));
  OAI21X1  g17170(.A0(new_n16962_), .A1(new_n16948_), .B0(new_n17234_), .Y(new_n17235_));
  AOI21X1  g17171(.A0(new_n17235_), .A1(new_n17033_), .B0(new_n17043_), .Y(new_n17236_));
  INVX1    g17172(.A(new_n17165_), .Y(new_n17237_));
  INVX1    g17173(.A(new_n17104_), .Y(new_n17238_));
  OAI21X1  g17174(.A0(new_n17238_), .A1(new_n17236_), .B0(new_n17237_), .Y(new_n17239_));
  AOI21X1  g17175(.A0(new_n17239_), .A1(new_n17163_), .B0(new_n17225_), .Y(new_n17240_));
  OAI21X1  g17176(.A0(new_n17240_), .A1(new_n17233_), .B0(new_n17232_), .Y(new_n17241_));
  INVX1    g17177(.A(new_n17212_), .Y(new_n17242_));
  NOR2X1   g17178(.A(new_n17218_), .B(new_n17215_), .Y(new_n17243_));
  AOI21X1  g17179(.A0(new_n17219_), .A1(new_n17242_), .B0(new_n17243_), .Y(new_n17244_));
  INVX1    g17180(.A(new_n17244_), .Y(new_n17245_));
  AND2X1   g17181(.A(new_n15362_), .B(new_n7342_), .Y(new_n17246_));
  XOR2X1   g17182(.A(new_n17246_), .B(new_n1920_), .Y(new_n17247_));
  OR4X1    g17183(.A(new_n1227_), .B(new_n666_), .C(new_n299_), .D(new_n118_), .Y(new_n17248_));
  OR4X1    g17184(.A(new_n596_), .B(new_n523_), .C(new_n383_), .D(new_n365_), .Y(new_n17249_));
  OR4X1    g17185(.A(new_n17249_), .B(new_n334_), .C(new_n321_), .D(new_n426_), .Y(new_n17250_));
  OR4X1    g17186(.A(new_n17250_), .B(new_n17248_), .C(new_n8179_), .D(new_n16970_), .Y(new_n17251_));
  OR4X1    g17187(.A(new_n8695_), .B(new_n2134_), .C(new_n1764_), .D(new_n802_), .Y(new_n17252_));
  NOR4X1   g17188(.A(new_n17252_), .B(new_n17251_), .C(new_n2539_), .D(new_n880_), .Y(new_n17253_));
  XOR2X1   g17189(.A(new_n17253_), .B(new_n17123_), .Y(new_n17254_));
  XOR2X1   g17190(.A(new_n17254_), .B(new_n17247_), .Y(new_n17255_));
  XOR2X1   g17191(.A(new_n17255_), .B(new_n17183_), .Y(new_n17256_));
  AOI22X1  g17192(.A0(new_n12076_), .A1(new_n1890_), .B0(new_n12018_), .B1(new_n1884_), .Y(new_n17257_));
  OAI21X1  g17193(.A0(new_n13679_), .A1(new_n3498_), .B0(new_n17257_), .Y(new_n17258_));
  AOI21X1  g17194(.A0(new_n13678_), .A1(new_n407_), .B0(new_n17258_), .Y(new_n17259_));
  XOR2X1   g17195(.A(new_n17259_), .B(new_n17256_), .Y(new_n17260_));
  NOR2X1   g17196(.A(new_n17188_), .B(new_n17185_), .Y(new_n17261_));
  AOI21X1  g17197(.A0(new_n17191_), .A1(new_n17189_), .B0(new_n17261_), .Y(new_n17262_));
  XOR2X1   g17198(.A(new_n17262_), .B(new_n17260_), .Y(new_n17263_));
  AOI22X1  g17199(.A0(new_n14085_), .A1(new_n2095_), .B0(new_n12285_), .B1(new_n2185_), .Y(new_n17264_));
  OAI21X1  g17200(.A0(new_n14088_), .A1(new_n2140_), .B0(new_n17264_), .Y(new_n17265_));
  AOI21X1  g17201(.A0(new_n14491_), .A1(new_n2062_), .B0(new_n17265_), .Y(new_n17266_));
  XOR2X1   g17202(.A(new_n17266_), .B(\a[29] ), .Y(new_n17267_));
  XOR2X1   g17203(.A(new_n17267_), .B(new_n17263_), .Y(new_n17268_));
  AOI22X1  g17204(.A0(new_n14642_), .A1(new_n2418_), .B0(new_n14084_), .B1(new_n2424_), .Y(new_n17269_));
  OAI21X1  g17205(.A0(new_n14805_), .A1(new_n2626_), .B0(new_n17269_), .Y(new_n17270_));
  AOI21X1  g17206(.A0(new_n14809_), .A1(new_n2301_), .B0(new_n17270_), .Y(new_n17271_));
  XOR2X1   g17207(.A(new_n17271_), .B(\a[26] ), .Y(new_n17272_));
  XOR2X1   g17208(.A(new_n17272_), .B(new_n17268_), .Y(new_n17273_));
  INVX1    g17209(.A(new_n17196_), .Y(new_n17274_));
  NOR2X1   g17210(.A(new_n17201_), .B(new_n17197_), .Y(new_n17275_));
  AOI21X1  g17211(.A0(new_n17274_), .A1(new_n17192_), .B0(new_n17275_), .Y(new_n17276_));
  XOR2X1   g17212(.A(new_n17276_), .B(new_n17273_), .Y(new_n17277_));
  NOR2X1   g17213(.A(new_n17206_), .B(new_n17203_), .Y(new_n17278_));
  INVX1    g17214(.A(new_n17278_), .Y(new_n17279_));
  INVX1    g17215(.A(new_n17207_), .Y(new_n17280_));
  OAI21X1  g17216(.A0(new_n17211_), .A1(new_n17280_), .B0(new_n17279_), .Y(new_n17281_));
  AOI22X1  g17217(.A0(new_n15087_), .A1(new_n2696_), .B0(new_n14946_), .B1(new_n2657_), .Y(new_n17282_));
  OAI21X1  g17218(.A0(new_n15363_), .A1(new_n2753_), .B0(new_n17282_), .Y(new_n17283_));
  AOI21X1  g17219(.A0(new_n15240_), .A1(new_n2658_), .B0(new_n17283_), .Y(new_n17284_));
  XOR2X1   g17220(.A(new_n17284_), .B(\a[23] ), .Y(new_n17285_));
  XOR2X1   g17221(.A(new_n17285_), .B(new_n17281_), .Y(new_n17286_));
  XOR2X1   g17222(.A(new_n17286_), .B(new_n17277_), .Y(new_n17287_));
  XOR2X1   g17223(.A(new_n17287_), .B(new_n17245_), .Y(new_n17288_));
  XOR2X1   g17224(.A(new_n17288_), .B(new_n17241_), .Y(new_n17289_));
  XOR2X1   g17225(.A(new_n17289_), .B(new_n17230_), .Y(\result[25] ));
  AND2X1   g17226(.A(new_n17289_), .B(new_n17230_), .Y(new_n17291_));
  NOR2X1   g17227(.A(new_n17262_), .B(new_n17260_), .Y(new_n17292_));
  INVX1    g17228(.A(new_n17292_), .Y(new_n17293_));
  INVX1    g17229(.A(new_n17263_), .Y(new_n17294_));
  OAI21X1  g17230(.A0(new_n17267_), .A1(new_n17294_), .B0(new_n17293_), .Y(new_n17295_));
  AOI22X1  g17231(.A0(new_n12074_), .A1(new_n1884_), .B0(new_n12018_), .B1(new_n1890_), .Y(new_n17296_));
  OAI21X1  g17232(.A0(new_n12292_), .A1(new_n3498_), .B0(new_n17296_), .Y(new_n17297_));
  AOI21X1  g17233(.A0(new_n12291_), .A1(new_n407_), .B0(new_n17297_), .Y(new_n17298_));
  NAND2X1  g17234(.A(new_n17254_), .B(new_n17247_), .Y(new_n17299_));
  OAI21X1  g17235(.A0(new_n17253_), .A1(new_n17123_), .B0(new_n17299_), .Y(new_n17300_));
  NOR2X1   g17236(.A(new_n565_), .B(new_n681_), .Y(new_n17301_));
  NOR4X1   g17237(.A(new_n293_), .B(new_n292_), .C(new_n291_), .D(new_n1008_), .Y(new_n17302_));
  NAND4X1  g17238(.A(new_n17302_), .B(new_n17301_), .C(new_n855_), .D(new_n345_), .Y(new_n17303_));
  OR4X1    g17239(.A(new_n2795_), .B(new_n1277_), .C(new_n1222_), .D(new_n1191_), .Y(new_n17304_));
  OR4X1    g17240(.A(new_n17304_), .B(new_n17303_), .C(new_n8739_), .D(new_n1908_), .Y(new_n17305_));
  NOR4X1   g17241(.A(new_n17305_), .B(new_n7926_), .C(new_n2026_), .D(new_n1243_), .Y(new_n17306_));
  XOR2X1   g17242(.A(new_n17306_), .B(new_n17300_), .Y(new_n17307_));
  XOR2X1   g17243(.A(new_n17307_), .B(new_n17298_), .Y(new_n17308_));
  INVX1    g17244(.A(new_n17308_), .Y(new_n17309_));
  INVX1    g17245(.A(new_n17256_), .Y(new_n17310_));
  NOR2X1   g17246(.A(new_n17259_), .B(new_n17310_), .Y(new_n17311_));
  AOI21X1  g17247(.A0(new_n17255_), .A1(new_n17183_), .B0(new_n17311_), .Y(new_n17312_));
  XOR2X1   g17248(.A(new_n17312_), .B(new_n17309_), .Y(new_n17313_));
  OAI22X1  g17249(.A0(new_n14088_), .A1(new_n2431_), .B0(new_n14086_), .B1(new_n2186_), .Y(new_n17314_));
  AOI21X1  g17250(.A0(new_n14084_), .A1(new_n2139_), .B0(new_n17314_), .Y(new_n17315_));
  OAI21X1  g17251(.A0(new_n14107_), .A1(new_n2063_), .B0(new_n17315_), .Y(new_n17316_));
  XOR2X1   g17252(.A(new_n17316_), .B(new_n74_), .Y(new_n17317_));
  XOR2X1   g17253(.A(new_n17317_), .B(new_n17313_), .Y(new_n17318_));
  XOR2X1   g17254(.A(new_n17318_), .B(new_n17295_), .Y(new_n17319_));
  AOI22X1  g17255(.A0(new_n14804_), .A1(new_n2418_), .B0(new_n14642_), .B1(new_n2424_), .Y(new_n17320_));
  OAI21X1  g17256(.A0(new_n15088_), .A1(new_n2626_), .B0(new_n17320_), .Y(new_n17321_));
  AOI21X1  g17257(.A0(new_n14952_), .A1(new_n2301_), .B0(new_n17321_), .Y(new_n17322_));
  XOR2X1   g17258(.A(new_n17322_), .B(\a[26] ), .Y(new_n17323_));
  XOR2X1   g17259(.A(new_n17323_), .B(new_n17319_), .Y(new_n17324_));
  OR2X1    g17260(.A(new_n17272_), .B(new_n17268_), .Y(new_n17325_));
  AND2X1   g17261(.A(new_n17274_), .B(new_n17192_), .Y(new_n17326_));
  OAI21X1  g17262(.A0(new_n17275_), .A1(new_n17326_), .B0(new_n17273_), .Y(new_n17327_));
  AND2X1   g17263(.A(new_n17327_), .B(new_n17325_), .Y(new_n17328_));
  XOR2X1   g17264(.A(new_n17328_), .B(new_n17324_), .Y(new_n17329_));
  AOI22X1  g17265(.A0(new_n15234_), .A1(new_n2696_), .B0(new_n15087_), .B1(new_n2657_), .Y(new_n17330_));
  OAI21X1  g17266(.A0(new_n15522_), .A1(new_n2753_), .B0(new_n17330_), .Y(new_n17331_));
  AOI21X1  g17267(.A0(new_n15841_), .A1(new_n2658_), .B0(new_n17331_), .Y(new_n17332_));
  XOR2X1   g17268(.A(new_n17332_), .B(\a[23] ), .Y(new_n17333_));
  XOR2X1   g17269(.A(new_n17333_), .B(new_n17329_), .Y(new_n17334_));
  INVX1    g17270(.A(new_n17285_), .Y(new_n17335_));
  NOR2X1   g17271(.A(new_n17286_), .B(new_n17277_), .Y(new_n17336_));
  AOI21X1  g17272(.A0(new_n17335_), .A1(new_n17281_), .B0(new_n17336_), .Y(new_n17337_));
  XOR2X1   g17273(.A(new_n17337_), .B(new_n17334_), .Y(new_n17338_));
  AOI21X1  g17274(.A0(new_n17227_), .A1(new_n17224_), .B0(new_n17231_), .Y(new_n17339_));
  AND2X1   g17275(.A(new_n17287_), .B(new_n17245_), .Y(new_n17340_));
  INVX1    g17276(.A(new_n17340_), .Y(new_n17341_));
  INVX1    g17277(.A(new_n17288_), .Y(new_n17342_));
  OAI21X1  g17278(.A0(new_n17342_), .A1(new_n17339_), .B0(new_n17341_), .Y(new_n17343_));
  XOR2X1   g17279(.A(new_n17343_), .B(new_n17338_), .Y(new_n17344_));
  XOR2X1   g17280(.A(new_n17344_), .B(new_n17291_), .Y(\result[26] ));
  INVX1    g17281(.A(new_n17298_), .Y(new_n17346_));
  AND2X1   g17282(.A(new_n17306_), .B(new_n17300_), .Y(new_n17347_));
  AOI21X1  g17283(.A0(new_n17307_), .A1(new_n17346_), .B0(new_n17347_), .Y(new_n17348_));
  OR4X1    g17284(.A(new_n7179_), .B(new_n1701_), .C(new_n7923_), .D(new_n714_), .Y(new_n17349_));
  OR4X1    g17285(.A(new_n724_), .B(new_n1166_), .C(new_n370_), .D(new_n327_), .Y(new_n17350_));
  OR4X1    g17286(.A(new_n17350_), .B(new_n513_), .C(new_n292_), .D(new_n291_), .Y(new_n17351_));
  OR4X1    g17287(.A(new_n17351_), .B(new_n17349_), .C(new_n8653_), .D(new_n7065_), .Y(new_n17352_));
  OR2X1    g17288(.A(new_n16180_), .B(new_n13980_), .Y(new_n17353_));
  NOR4X1   g17289(.A(new_n17353_), .B(new_n17352_), .C(new_n12415_), .D(new_n2509_), .Y(new_n17354_));
  XOR2X1   g17290(.A(new_n17354_), .B(new_n17306_), .Y(new_n17355_));
  NOR2X1   g17291(.A(new_n17355_), .B(new_n17348_), .Y(new_n17356_));
  OR2X1    g17292(.A(new_n17356_), .B(new_n17348_), .Y(new_n17357_));
  INVX1    g17293(.A(new_n17306_), .Y(new_n17358_));
  AND2X1   g17294(.A(new_n17354_), .B(new_n17358_), .Y(new_n17359_));
  NOR2X1   g17295(.A(new_n17356_), .B(new_n17359_), .Y(new_n17360_));
  OAI21X1  g17296(.A0(new_n17354_), .A1(new_n17358_), .B0(new_n17360_), .Y(new_n17361_));
  AND2X1   g17297(.A(new_n17361_), .B(new_n17357_), .Y(new_n17362_));
  AOI22X1  g17298(.A0(new_n12285_), .A1(new_n1884_), .B0(new_n12074_), .B1(new_n1890_), .Y(new_n17363_));
  OAI21X1  g17299(.A0(new_n14086_), .A1(new_n3498_), .B0(new_n17363_), .Y(new_n17364_));
  AOI21X1  g17300(.A0(new_n14480_), .A1(new_n407_), .B0(new_n17364_), .Y(new_n17365_));
  XOR2X1   g17301(.A(new_n17365_), .B(new_n17362_), .Y(new_n17366_));
  OR2X1    g17302(.A(new_n17312_), .B(new_n17308_), .Y(new_n17367_));
  OAI21X1  g17303(.A0(new_n17317_), .A1(new_n17313_), .B0(new_n17367_), .Y(new_n17368_));
  XOR2X1   g17304(.A(new_n17368_), .B(new_n17366_), .Y(new_n17369_));
  AOI22X1  g17305(.A0(new_n14087_), .A1(new_n2185_), .B0(new_n14084_), .B1(new_n2095_), .Y(new_n17370_));
  OAI21X1  g17306(.A0(new_n14648_), .A1(new_n2140_), .B0(new_n17370_), .Y(new_n17371_));
  AOI21X1  g17307(.A0(new_n14651_), .A1(new_n2062_), .B0(new_n17371_), .Y(new_n17372_));
  XOR2X1   g17308(.A(new_n17372_), .B(\a[29] ), .Y(new_n17373_));
  XOR2X1   g17309(.A(new_n17373_), .B(new_n17369_), .Y(new_n17374_));
  AOI22X1  g17310(.A0(new_n14946_), .A1(new_n2418_), .B0(new_n14804_), .B1(new_n2424_), .Y(new_n17375_));
  OAI21X1  g17311(.A0(new_n15235_), .A1(new_n2626_), .B0(new_n17375_), .Y(new_n17376_));
  AOI21X1  g17312(.A0(new_n15381_), .A1(new_n2301_), .B0(new_n17376_), .Y(new_n17377_));
  XOR2X1   g17313(.A(new_n17377_), .B(\a[26] ), .Y(new_n17378_));
  XOR2X1   g17314(.A(new_n17378_), .B(new_n17374_), .Y(new_n17379_));
  AND2X1   g17315(.A(new_n17318_), .B(new_n17295_), .Y(new_n17380_));
  INVX1    g17316(.A(new_n17323_), .Y(new_n17381_));
  AOI21X1  g17317(.A0(new_n17381_), .A1(new_n17319_), .B0(new_n17380_), .Y(new_n17382_));
  AOI22X1  g17318(.A0(new_n15362_), .A1(new_n12061_), .B0(new_n15234_), .B1(new_n2657_), .Y(new_n17383_));
  OAI21X1  g17319(.A0(new_n15373_), .A1(new_n2692_), .B0(new_n17383_), .Y(new_n17384_));
  XOR2X1   g17320(.A(new_n17384_), .B(new_n70_), .Y(new_n17385_));
  XOR2X1   g17321(.A(new_n17385_), .B(new_n17382_), .Y(new_n17386_));
  XOR2X1   g17322(.A(new_n17386_), .B(new_n17379_), .Y(new_n17387_));
  INVX1    g17323(.A(new_n17387_), .Y(new_n17388_));
  NOR2X1   g17324(.A(new_n17328_), .B(new_n17324_), .Y(new_n17389_));
  INVX1    g17325(.A(new_n17333_), .Y(new_n17390_));
  AOI21X1  g17326(.A0(new_n17390_), .A1(new_n17329_), .B0(new_n17389_), .Y(new_n17391_));
  XOR2X1   g17327(.A(new_n17391_), .B(new_n17388_), .Y(new_n17392_));
  INVX1    g17328(.A(new_n17392_), .Y(new_n17393_));
  NOR2X1   g17329(.A(new_n17337_), .B(new_n17334_), .Y(new_n17394_));
  AOI21X1  g17330(.A0(new_n17343_), .A1(new_n17338_), .B0(new_n17394_), .Y(new_n17395_));
  XOR2X1   g17331(.A(new_n17395_), .B(new_n17393_), .Y(new_n17396_));
  AND2X1   g17332(.A(new_n17344_), .B(new_n17291_), .Y(new_n17397_));
  XOR2X1   g17333(.A(new_n17397_), .B(new_n17396_), .Y(\result[27] ));
  AND2X1   g17334(.A(new_n17397_), .B(new_n17396_), .Y(new_n17399_));
  NOR2X1   g17335(.A(new_n17391_), .B(new_n17388_), .Y(new_n17400_));
  INVX1    g17336(.A(new_n17400_), .Y(new_n17401_));
  OAI21X1  g17337(.A0(new_n17395_), .A1(new_n17393_), .B0(new_n17401_), .Y(new_n17402_));
  NOR2X1   g17338(.A(new_n17385_), .B(new_n17382_), .Y(new_n17403_));
  AOI21X1  g17339(.A0(new_n17386_), .A1(new_n17379_), .B0(new_n17403_), .Y(new_n17404_));
  INVX1    g17340(.A(new_n17373_), .Y(new_n17405_));
  NOR2X1   g17341(.A(new_n17378_), .B(new_n17374_), .Y(new_n17406_));
  AOI21X1  g17342(.A0(new_n17405_), .A1(new_n17369_), .B0(new_n17406_), .Y(new_n17407_));
  AOI22X1  g17343(.A0(new_n15087_), .A1(new_n2418_), .B0(new_n14946_), .B1(new_n2424_), .Y(new_n17408_));
  OAI21X1  g17344(.A0(new_n15363_), .A1(new_n2626_), .B0(new_n17408_), .Y(new_n17409_));
  AOI21X1  g17345(.A0(new_n15240_), .A1(new_n2301_), .B0(new_n17409_), .Y(new_n17410_));
  XOR2X1   g17346(.A(new_n17410_), .B(\a[26] ), .Y(new_n17411_));
  XOR2X1   g17347(.A(new_n17411_), .B(new_n17407_), .Y(new_n17412_));
  AND2X1   g17348(.A(new_n15362_), .B(new_n12259_), .Y(new_n17413_));
  XOR2X1   g17349(.A(new_n17413_), .B(new_n70_), .Y(new_n17414_));
  INVX1    g17350(.A(new_n2400_), .Y(new_n17415_));
  NOR4X1   g17351(.A(new_n632_), .B(new_n259_), .C(new_n199_), .D(new_n124_), .Y(new_n17416_));
  NOR3X1   g17352(.A(new_n427_), .B(new_n479_), .C(new_n746_), .Y(new_n17417_));
  NAND3X1  g17353(.A(new_n17417_), .B(new_n17416_), .C(new_n1164_), .Y(new_n17418_));
  OR4X1    g17354(.A(new_n2805_), .B(new_n921_), .C(new_n823_), .D(new_n514_), .Y(new_n17419_));
  OR4X1    g17355(.A(new_n17419_), .B(new_n17418_), .C(new_n17415_), .D(new_n2357_), .Y(new_n17420_));
  NOR2X1   g17356(.A(new_n17420_), .B(new_n7147_), .Y(new_n17421_));
  XOR2X1   g17357(.A(new_n17421_), .B(new_n17354_), .Y(new_n17422_));
  XOR2X1   g17358(.A(new_n17422_), .B(new_n17414_), .Y(new_n17423_));
  XOR2X1   g17359(.A(new_n17423_), .B(new_n17360_), .Y(new_n17424_));
  AOI22X1  g17360(.A0(new_n14085_), .A1(new_n1884_), .B0(new_n12285_), .B1(new_n1890_), .Y(new_n17425_));
  OAI21X1  g17361(.A0(new_n14088_), .A1(new_n3498_), .B0(new_n17425_), .Y(new_n17426_));
  AOI21X1  g17362(.A0(new_n14491_), .A1(new_n407_), .B0(new_n17426_), .Y(new_n17427_));
  XOR2X1   g17363(.A(new_n17427_), .B(new_n17424_), .Y(new_n17428_));
  INVX1    g17364(.A(new_n17428_), .Y(new_n17429_));
  AOI21X1  g17365(.A0(new_n17361_), .A1(new_n17357_), .B0(new_n17365_), .Y(new_n17430_));
  AOI21X1  g17366(.A0(new_n17368_), .A1(new_n17366_), .B0(new_n17430_), .Y(new_n17431_));
  XOR2X1   g17367(.A(new_n17431_), .B(new_n17429_), .Y(new_n17432_));
  AOI22X1  g17368(.A0(new_n14642_), .A1(new_n2095_), .B0(new_n14084_), .B1(new_n2185_), .Y(new_n17433_));
  OAI21X1  g17369(.A0(new_n14805_), .A1(new_n2140_), .B0(new_n17433_), .Y(new_n17434_));
  AOI21X1  g17370(.A0(new_n14809_), .A1(new_n2062_), .B0(new_n17434_), .Y(new_n17435_));
  XOR2X1   g17371(.A(new_n17435_), .B(\a[29] ), .Y(new_n17436_));
  XOR2X1   g17372(.A(new_n17436_), .B(new_n17432_), .Y(new_n17437_));
  XOR2X1   g17373(.A(new_n17437_), .B(new_n17412_), .Y(new_n17438_));
  XOR2X1   g17374(.A(new_n17438_), .B(new_n17404_), .Y(new_n17439_));
  XOR2X1   g17375(.A(new_n17439_), .B(new_n17402_), .Y(new_n17440_));
  XOR2X1   g17376(.A(new_n17440_), .B(new_n17399_), .Y(\result[28] ));
  AND2X1   g17377(.A(new_n17440_), .B(new_n17399_), .Y(new_n17442_));
  NOR2X1   g17378(.A(new_n17431_), .B(new_n17429_), .Y(new_n17443_));
  INVX1    g17379(.A(new_n17436_), .Y(new_n17444_));
  AOI21X1  g17380(.A0(new_n17444_), .A1(new_n17432_), .B0(new_n17443_), .Y(new_n17445_));
  AOI22X1  g17381(.A0(new_n14087_), .A1(new_n1884_), .B0(new_n14085_), .B1(new_n1890_), .Y(new_n17446_));
  OAI21X1  g17382(.A0(new_n14643_), .A1(new_n3498_), .B0(new_n17446_), .Y(new_n17447_));
  AOI21X1  g17383(.A0(new_n14106_), .A1(new_n407_), .B0(new_n17447_), .Y(new_n17448_));
  NAND2X1  g17384(.A(new_n17422_), .B(new_n17414_), .Y(new_n17449_));
  OAI21X1  g17385(.A0(new_n17421_), .A1(new_n17354_), .B0(new_n17449_), .Y(new_n17450_));
  NOR3X1   g17386(.A(new_n945_), .B(new_n229_), .C(new_n194_), .Y(new_n17451_));
  NOR4X1   g17387(.A(new_n1105_), .B(new_n463_), .C(new_n335_), .D(new_n272_), .Y(new_n17452_));
  NOR3X1   g17388(.A(new_n1975_), .B(new_n383_), .C(new_n565_), .Y(new_n17453_));
  NAND3X1  g17389(.A(new_n17453_), .B(new_n17452_), .C(new_n17451_), .Y(new_n17454_));
  OR4X1    g17390(.A(new_n3741_), .B(new_n1320_), .C(new_n1275_), .D(new_n1142_), .Y(new_n17455_));
  NOR4X1   g17391(.A(new_n17455_), .B(new_n17454_), .C(new_n2352_), .D(new_n2331_), .Y(new_n17456_));
  NAND3X1  g17392(.A(new_n17456_), .B(new_n14058_), .C(new_n8638_), .Y(new_n17457_));
  INVX1    g17393(.A(new_n17457_), .Y(new_n17458_));
  XOR2X1   g17394(.A(new_n17458_), .B(new_n17450_), .Y(new_n17459_));
  XOR2X1   g17395(.A(new_n17459_), .B(new_n17448_), .Y(new_n17460_));
  INVX1    g17396(.A(new_n17460_), .Y(new_n17461_));
  OAI21X1  g17397(.A0(new_n17356_), .A1(new_n17359_), .B0(new_n17423_), .Y(new_n17462_));
  OAI21X1  g17398(.A0(new_n17427_), .A1(new_n17424_), .B0(new_n17462_), .Y(new_n17463_));
  XOR2X1   g17399(.A(new_n17463_), .B(new_n17461_), .Y(new_n17464_));
  INVX1    g17400(.A(new_n17464_), .Y(new_n17465_));
  OAI22X1  g17401(.A0(new_n14805_), .A1(new_n2431_), .B0(new_n14648_), .B1(new_n2186_), .Y(new_n17466_));
  AOI21X1  g17402(.A0(new_n14946_), .A1(new_n2139_), .B0(new_n17466_), .Y(new_n17467_));
  OAI21X1  g17403(.A0(new_n14953_), .A1(new_n2063_), .B0(new_n17467_), .Y(new_n17468_));
  XOR2X1   g17404(.A(new_n17468_), .B(new_n74_), .Y(new_n17469_));
  XOR2X1   g17405(.A(new_n17469_), .B(new_n17465_), .Y(new_n17470_));
  XOR2X1   g17406(.A(new_n17470_), .B(new_n17445_), .Y(new_n17471_));
  AOI22X1  g17407(.A0(new_n15234_), .A1(new_n2418_), .B0(new_n15087_), .B1(new_n2424_), .Y(new_n17472_));
  OAI21X1  g17408(.A0(new_n15522_), .A1(new_n2626_), .B0(new_n17472_), .Y(new_n17473_));
  AOI21X1  g17409(.A0(new_n15841_), .A1(new_n2301_), .B0(new_n17473_), .Y(new_n17474_));
  XOR2X1   g17410(.A(new_n17474_), .B(\a[26] ), .Y(new_n17475_));
  XOR2X1   g17411(.A(new_n17475_), .B(new_n17471_), .Y(new_n17476_));
  NOR2X1   g17412(.A(new_n17411_), .B(new_n17407_), .Y(new_n17477_));
  INVX1    g17413(.A(new_n17437_), .Y(new_n17478_));
  AOI21X1  g17414(.A0(new_n17478_), .A1(new_n17412_), .B0(new_n17477_), .Y(new_n17479_));
  XOR2X1   g17415(.A(new_n17479_), .B(new_n17476_), .Y(new_n17480_));
  NOR2X1   g17416(.A(new_n17438_), .B(new_n17404_), .Y(new_n17481_));
  AOI21X1  g17417(.A0(new_n17439_), .A1(new_n17402_), .B0(new_n17481_), .Y(new_n17482_));
  XOR2X1   g17418(.A(new_n17482_), .B(new_n17480_), .Y(new_n17483_));
  XOR2X1   g17419(.A(new_n17483_), .B(new_n17442_), .Y(\result[29] ));
  AND2X1   g17420(.A(new_n17483_), .B(new_n17442_), .Y(new_n17485_));
  INVX1    g17421(.A(new_n17476_), .Y(new_n17486_));
  NOR2X1   g17422(.A(new_n17479_), .B(new_n17486_), .Y(new_n17487_));
  INVX1    g17423(.A(new_n17487_), .Y(new_n17488_));
  OAI21X1  g17424(.A0(new_n17482_), .A1(new_n17480_), .B0(new_n17488_), .Y(new_n17489_));
  INVX1    g17425(.A(new_n17470_), .Y(new_n17490_));
  OR2X1    g17426(.A(new_n17490_), .B(new_n17445_), .Y(new_n17491_));
  OAI21X1  g17427(.A0(new_n17475_), .A1(new_n17471_), .B0(new_n17491_), .Y(new_n17492_));
  INVX1    g17428(.A(new_n17448_), .Y(new_n17493_));
  AND2X1   g17429(.A(new_n17458_), .B(new_n17450_), .Y(new_n17494_));
  AOI21X1  g17430(.A0(new_n17459_), .A1(new_n17493_), .B0(new_n17494_), .Y(new_n17495_));
  INVX1    g17431(.A(new_n17495_), .Y(new_n17496_));
  OR4X1    g17432(.A(new_n7103_), .B(new_n2392_), .C(new_n2363_), .D(new_n199_), .Y(new_n17497_));
  NAND3X1  g17433(.A(new_n2412_), .B(new_n2348_), .C(new_n1511_), .Y(new_n17498_));
  NOR3X1   g17434(.A(new_n17498_), .B(new_n17497_), .C(new_n14059_), .Y(new_n17499_));
  XOR2X1   g17435(.A(new_n17499_), .B(new_n17458_), .Y(new_n17500_));
  OR2X1    g17436(.A(new_n17499_), .B(new_n17457_), .Y(new_n17501_));
  OAI21X1  g17437(.A0(new_n17500_), .A1(new_n17495_), .B0(new_n17501_), .Y(new_n17502_));
  AOI21X1  g17438(.A0(new_n17499_), .A1(new_n17457_), .B0(new_n17502_), .Y(new_n17503_));
  AOI21X1  g17439(.A0(new_n17500_), .A1(new_n17496_), .B0(new_n17503_), .Y(new_n17504_));
  AOI22X1  g17440(.A0(new_n14087_), .A1(new_n1890_), .B0(new_n14084_), .B1(new_n1884_), .Y(new_n17505_));
  OAI21X1  g17441(.A0(new_n14648_), .A1(new_n3498_), .B0(new_n17505_), .Y(new_n17506_));
  AOI21X1  g17442(.A0(new_n14651_), .A1(new_n407_), .B0(new_n17506_), .Y(new_n17507_));
  XOR2X1   g17443(.A(new_n17507_), .B(new_n17504_), .Y(new_n17508_));
  AND2X1   g17444(.A(new_n17463_), .B(new_n17461_), .Y(new_n17509_));
  INVX1    g17445(.A(new_n17509_), .Y(new_n17510_));
  OAI21X1  g17446(.A0(new_n17469_), .A1(new_n17465_), .B0(new_n17510_), .Y(new_n17511_));
  INVX1    g17447(.A(new_n17511_), .Y(new_n17512_));
  XOR2X1   g17448(.A(new_n17512_), .B(new_n17508_), .Y(new_n17513_));
  NOR2X1   g17449(.A(new_n15373_), .B(new_n2665_), .Y(new_n17514_));
  OAI22X1  g17450(.A0(new_n15522_), .A1(new_n14030_), .B0(new_n15363_), .B1(new_n2666_), .Y(new_n17515_));
  NOR2X1   g17451(.A(new_n17515_), .B(new_n17514_), .Y(new_n17516_));
  XOR2X1   g17452(.A(new_n17516_), .B(\a[26] ), .Y(new_n17517_));
  AOI22X1  g17453(.A0(new_n14946_), .A1(new_n2095_), .B0(new_n14804_), .B1(new_n2185_), .Y(new_n17518_));
  OAI21X1  g17454(.A0(new_n15235_), .A1(new_n2140_), .B0(new_n17518_), .Y(new_n17519_));
  AOI21X1  g17455(.A0(new_n15381_), .A1(new_n2062_), .B0(new_n17519_), .Y(new_n17520_));
  XOR2X1   g17456(.A(new_n17520_), .B(\a[29] ), .Y(new_n17521_));
  INVX1    g17457(.A(new_n17521_), .Y(new_n17522_));
  XOR2X1   g17458(.A(new_n17522_), .B(new_n17517_), .Y(new_n17523_));
  XOR2X1   g17459(.A(new_n17523_), .B(new_n17513_), .Y(new_n17524_));
  XOR2X1   g17460(.A(new_n17524_), .B(new_n17492_), .Y(new_n17525_));
  XOR2X1   g17461(.A(new_n17525_), .B(new_n17489_), .Y(new_n17526_));
  XOR2X1   g17462(.A(new_n17526_), .B(new_n17485_), .Y(\result[30] ));
  NAND2X1  g17463(.A(new_n17526_), .B(new_n17485_), .Y(new_n17528_));
  AND2X1   g17464(.A(new_n17524_), .B(new_n17492_), .Y(new_n17529_));
  AOI21X1  g17465(.A0(new_n17525_), .A1(new_n17489_), .B0(new_n17529_), .Y(new_n17530_));
  OAI22X1  g17466(.A0(new_n15235_), .A1(new_n2431_), .B0(new_n15088_), .B1(new_n2186_), .Y(new_n17531_));
  AOI21X1  g17467(.A0(new_n15234_), .A1(new_n2139_), .B0(new_n17531_), .Y(new_n17532_));
  OAI21X1  g17468(.A0(new_n15241_), .A1(new_n2063_), .B0(new_n17532_), .Y(new_n17533_));
  NOR2X1   g17469(.A(new_n17507_), .B(new_n17504_), .Y(new_n17534_));
  AOI21X1  g17470(.A0(new_n17511_), .A1(new_n17508_), .B0(new_n17534_), .Y(new_n17535_));
  XOR2X1   g17471(.A(new_n17535_), .B(new_n74_), .Y(new_n17536_));
  XOR2X1   g17472(.A(new_n17536_), .B(new_n17533_), .Y(new_n17537_));
  AOI22X1  g17473(.A0(new_n14642_), .A1(new_n1884_), .B0(new_n14084_), .B1(new_n1890_), .Y(new_n17538_));
  OAI21X1  g17474(.A0(new_n14805_), .A1(new_n3498_), .B0(new_n17538_), .Y(new_n17539_));
  AOI21X1  g17475(.A0(new_n14809_), .A1(new_n407_), .B0(new_n17539_), .Y(new_n17540_));
  XOR2X1   g17476(.A(new_n17540_), .B(new_n17502_), .Y(new_n17541_));
  XOR2X1   g17477(.A(new_n17541_), .B(new_n17537_), .Y(new_n17542_));
  OR2X1    g17478(.A(new_n17521_), .B(new_n17517_), .Y(new_n17543_));
  OAI21X1  g17479(.A0(new_n17523_), .A1(new_n17513_), .B0(new_n17543_), .Y(new_n17544_));
  NOR3X1   g17480(.A(new_n2646_), .B(new_n2405_), .C(new_n197_), .Y(new_n17545_));
  XOR2X1   g17481(.A(new_n17545_), .B(new_n89_), .Y(new_n17546_));
  AND2X1   g17482(.A(new_n15362_), .B(new_n14055_), .Y(new_n17547_));
  XOR2X1   g17483(.A(new_n17547_), .B(new_n17457_), .Y(new_n17548_));
  XOR2X1   g17484(.A(new_n17548_), .B(new_n17546_), .Y(new_n17549_));
  XOR2X1   g17485(.A(new_n17549_), .B(new_n17544_), .Y(new_n17550_));
  XOR2X1   g17486(.A(new_n17550_), .B(new_n17542_), .Y(new_n17551_));
  XOR2X1   g17487(.A(new_n17551_), .B(new_n17530_), .Y(new_n17552_));
  XOR2X1   g17488(.A(new_n17552_), .B(new_n17528_), .Y(\result[31] ));
endmodule


