// Benchmark "c432.blif" written by ABC on Sun Apr 15 22:34:58 2018

module c432.blif ( 
    G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat, G27gat,
    G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat, G56gat,
    G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat, G86gat,
    G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat, G112gat,
    G115gat,
    G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat  );
  input  G1gat, G4gat, G8gat, G11gat, G14gat, G17gat, G21gat, G24gat,
    G27gat, G30gat, G34gat, G37gat, G40gat, G43gat, G47gat, G50gat, G53gat,
    G56gat, G60gat, G63gat, G66gat, G69gat, G73gat, G76gat, G79gat, G82gat,
    G86gat, G89gat, G92gat, G95gat, G99gat, G102gat, G105gat, G108gat,
    G112gat, G115gat;
  output G223gat, G329gat, G370gat, G421gat, G430gat, G431gat, G432gat;
  wire n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n71, n72,
    n73, n74, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n103,
    n104, n105, n109, n110, n111, n112, n113, n117, n118, n119, n123, n124,
    n125, n126, n129, n130, n131, n132, n135, n136, n137, n138, n139, n142,
    n143, n144, n145, n148, n149, n150, n151, n152, n153, n154, n158, n159,
    n160, n162, n163, n164, n165, n167, n168, n169, n170, n171, n172, n173,
    n175, n176, n177, n179, n180, n181, n182, n185, n186, n189, n190, n191,
    n194, n195, n198, n199, n200, n201, n202, n203, n204, n206, n207, n208,
    n209, n210, n213, n214, n215, n216, n217, n218, n219, n222, n223, n224,
    n225, n226, n229, n230, n231, n232, n233, n234, n237, n238, n239, n240,
    n243, n244, n245, n246, n247, n250, n251, n252, n253, n256, n257, n258,
    n259, n260, n261, n262, n264, n265, n268, n269, n272, n273, n274, n275,
    n278, n279, n282, n283, n284, n287, n288, n289, n292, n293, n294, n295,
    n298, n299, n300, n303, n304, n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
    n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378, n379, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416;
  "!a"     g000(.a(G108gat), .O(n43));
  "(a+b)'" g001(.a(n43), .b(G102gat), .O(n44));
  "!a"     g002(.a(G89gat), .O(n45));
  "(ab)'"  g003(.a(G95gat), .b(n45), .O(n46));
  "!a"     g004(.a(G76gat), .O(n47));
  "(ab)'"  g005(.a(G82gat), .b(n47), .O(n48));
  "(ab)'"  g006(.a(n48), .b(n46), .O(n49));
  "(a+b)'" g007(.a(n49), .b(n44), .O(n50));
  "!a"     g008(.a(G1gat), .O(n51));
  "(ab)'"  g009(.a(G4gat), .b(n51), .O(n52));
  "!a"     g010(.a(G11gat), .O(n53));
  "(ab)'"  g011(.a(G17gat), .b(n53), .O(n54));
  "(ab)'"  g012(.a(n54), .b(n52), .O(n55));
  "!a"     g013(.a(G43gat), .O(n56));
  "(a+b)'" g014(.a(n56), .b(G37gat), .O(n57));
  "!a"     g015(.a(G30gat), .O(n58));
  "(a+b)'" g016(.a(n58), .b(G24gat), .O(n59));
  "(a+b)'" g017(.a(n59), .b(n57), .O(n60));
  "!a"     g018(.a(G69gat), .O(n61));
  "(a+b)'" g019(.a(n61), .b(G63gat), .O(n62));
  "!a"     g020(.a(G56gat), .O(n63));
  "(a+b)'" g021(.a(n63), .b(G50gat), .O(n64));
  "(a+b)'" g022(.a(n64), .b(n62), .O(n65));
  "(ab)'"  g023(.a(n65), .b(n60), .O(n66));
  "(a+b)'" g024(.a(n66), .b(n55), .O(n67));
  "(ab)'"  g025(.a(n67), .b(n50), .O(G223gat));
  "!a"     g026(.a(G95gat), .O(n70));
  "(a+b)'" g027(.a(n70), .b(G89gat), .O(n71));
  "!a"     g028(.a(G82gat), .O(n72));
  "(a+b)'" g029(.a(n72), .b(G76gat), .O(n73));
  "(a+b)'" g030(.a(n73), .b(n71), .O(n74));
  "(a+b)'" g031(.a(n44), .b(n99), .O(n76));
  "(a+b)'" g032(.a(G112gat), .b(n43), .O(n77));
  "!a"     g033(.a(n77), .O(n78));
  "(a+b)'" g034(.a(n78), .b(n76), .O(n79));
  "!a"     g035(.a(n44), .O(n80));
  "(ab)'"  g036(.a(n74), .b(n80), .O(n81));
  "!a"     g037(.a(G4gat), .O(n82));
  "(a+b)'" g038(.a(n82), .b(G1gat), .O(n83));
  "!a"     g039(.a(G17gat), .O(n84));
  "(a+b)'" g040(.a(n84), .b(G11gat), .O(n85));
  "(a+b)'" g041(.a(n85), .b(n83), .O(n86));
  "!a"     g042(.a(G37gat), .O(n87));
  "(ab)'"  g043(.a(G43gat), .b(n87), .O(n88));
  "!a"     g044(.a(G24gat), .O(n89));
  "(ab)'"  g045(.a(G30gat), .b(n89), .O(n90));
  "(ab)'"  g046(.a(n90), .b(n88), .O(n91));
  "!a"     g047(.a(G63gat), .O(n92));
  "(ab)'"  g048(.a(G69gat), .b(n92), .O(n93));
  "!a"     g049(.a(G50gat), .O(n94));
  "(ab)'"  g050(.a(G56gat), .b(n94), .O(n95));
  "(ab)'"  g051(.a(n95), .b(n93), .O(n96));
  "(a+b)'" g052(.a(n96), .b(n91), .O(n97));
  "(ab)'"  g053(.a(n97), .b(n86), .O(n98));
  "(a+b)'" g054(.a(n98), .b(n81), .O(n99));
  "(ab)'"  g055(.a(n99), .b(n46), .O(n100));
  "(ab)'"  g056(.a(n46), .b(n100), .O(n103));
  "(a+b)'" g057(.a(G99gat), .b(n70), .O(n104));
  "(ab)'"  g058(.a(n104), .b(n103), .O(n105));
  "(ab)'"  g059(.a(n48), .b(n100), .O(n109));
  "(a+b)'" g060(.a(G86gat), .b(n72), .O(n110));
  "(ab)'"  g061(.a(n110), .b(n109), .O(n111));
  "(ab)'"  g062(.a(n111), .b(n105), .O(n112));
  "(a+b)'" g063(.a(n112), .b(n79), .O(n113));
  "(ab)'"  g064(.a(n52), .b(n100), .O(n117));
  "(a+b)'" g065(.a(G8gat), .b(n82), .O(n118));
  "(ab)'"  g066(.a(n118), .b(n117), .O(n119));
  "(ab)'"  g067(.a(n54), .b(n100), .O(n123));
  "(a+b)'" g068(.a(G21gat), .b(n84), .O(n124));
  "(ab)'"  g069(.a(n124), .b(n123), .O(n125));
  "(ab)'"  g070(.a(n125), .b(n119), .O(n126));
  "(a+b)'" g071(.a(n57), .b(n99), .O(n129));
  "(a+b)'" g072(.a(G47gat), .b(n56), .O(n130));
  "!a"     g073(.a(n130), .O(n131));
  "(a+b)'" g074(.a(n131), .b(n129), .O(n132));
  "(a+b)'" g075(.a(n59), .b(n99), .O(n135));
  "(a+b)'" g076(.a(G34gat), .b(n58), .O(n136));
  "!a"     g077(.a(n136), .O(n137));
  "(a+b)'" g078(.a(n137), .b(n135), .O(n138));
  "(a+b)'" g079(.a(n138), .b(n132), .O(n139));
  "(a+b)'" g080(.a(n62), .b(n99), .O(n142));
  "(a+b)'" g081(.a(G73gat), .b(n61), .O(n143));
  "!a"     g082(.a(n143), .O(n144));
  "(a+b)'" g083(.a(n144), .b(n142), .O(n145));
  "(a+b)'" g084(.a(n64), .b(n99), .O(n148));
  "(a+b)'" g085(.a(G60gat), .b(n63), .O(n149));
  "!a"     g086(.a(n149), .O(n150));
  "(a+b)'" g087(.a(n150), .b(n148), .O(n151));
  "(a+b)'" g088(.a(n151), .b(n145), .O(n152));
  "(ab)'"  g089(.a(n152), .b(n139), .O(n153));
  "(a+b)'" g090(.a(n153), .b(n126), .O(n154));
  "(ab)'"  g091(.a(n154), .b(n113), .O(G329gat));
  "(a+b)'" g092(.a(n71), .b(n99), .O(n158));
  "!a"     g093(.a(n104), .O(n159));
  "(a+b)'" g094(.a(n159), .b(n158), .O(n160));
  "(a+b)'" g095(.a(n73), .b(n99), .O(n162));
  "!a"     g096(.a(n110), .O(n163));
  "(a+b)'" g097(.a(n163), .b(n162), .O(n164));
  "(a+b)'" g098(.a(n164), .b(n160), .O(n165));
  "(a+b)'" g099(.a(n79), .b(n203), .O(n167));
  "!a"     g100(.a(n76), .O(n168));
  "(a+b)'" g101(.a(G115gat), .b(n43), .O(n169));
  "(ab)'"  g102(.a(n169), .b(n168), .O(n170));
  "(a+b)'" g103(.a(n170), .b(n167), .O(n171));
  "!a"     g104(.a(n79), .O(n172));
  "(ab)'"  g105(.a(n165), .b(n172), .O(n173));
  "(a+b)'" g106(.a(n83), .b(n99), .O(n175));
  "!a"     g107(.a(n118), .O(n176));
  "(a+b)'" g108(.a(n176), .b(n175), .O(n177));
  "(a+b)'" g109(.a(n85), .b(n99), .O(n179));
  "!a"     g110(.a(n124), .O(n180));
  "(a+b)'" g111(.a(n180), .b(n179), .O(n181));
  "(a+b)'" g112(.a(n181), .b(n177), .O(n182));
  "(ab)'"  g113(.a(n88), .b(n100), .O(n185));
  "(ab)'"  g114(.a(n130), .b(n185), .O(n186));
  "(ab)'"  g115(.a(n90), .b(n100), .O(n189));
  "(ab)'"  g116(.a(n136), .b(n189), .O(n190));
  "(ab)'"  g117(.a(n190), .b(n186), .O(n191));
  "(ab)'"  g118(.a(n93), .b(n100), .O(n194));
  "(ab)'"  g119(.a(n143), .b(n194), .O(n195));
  "(ab)'"  g120(.a(n95), .b(n100), .O(n198));
  "(ab)'"  g121(.a(n149), .b(n198), .O(n199));
  "(ab)'"  g122(.a(n199), .b(n195), .O(n200));
  "(a+b)'" g123(.a(n200), .b(n191), .O(n201));
  "(ab)'"  g124(.a(n201), .b(n182), .O(n202));
  "(a+b)'" g125(.a(n202), .b(n173), .O(n203));
  "(ab)'"  g126(.a(n203), .b(n105), .O(n204));
  "(ab)'"  g127(.a(n105), .b(n204), .O(n206));
  "(a+b)'" g128(.a(G105gat), .b(n70), .O(n207));
  "(ab)'"  g129(.a(n207), .b(n103), .O(n208));
  "!a"     g130(.a(n208), .O(n209));
  "(ab)'"  g131(.a(n209), .b(n206), .O(n210));
  "(ab)'"  g132(.a(n111), .b(n204), .O(n213));
  "(a+b)'" g133(.a(G92gat), .b(n72), .O(n214));
  "(ab)'"  g134(.a(n214), .b(n109), .O(n215));
  "!a"     g135(.a(n215), .O(n216));
  "(ab)'"  g136(.a(n216), .b(n213), .O(n217));
  "(ab)'"  g137(.a(n217), .b(n210), .O(n218));
  "(a+b)'" g138(.a(n218), .b(n171), .O(n219));
  "(ab)'"  g139(.a(n119), .b(n204), .O(n222));
  "(a+b)'" g140(.a(G14gat), .b(n82), .O(n223));
  "(ab)'"  g141(.a(n223), .b(n117), .O(n224));
  "!a"     g142(.a(n224), .O(n225));
  "(ab)'"  g143(.a(n225), .b(n222), .O(n226));
  "(ab)'"  g144(.a(n125), .b(n204), .O(n229));
  "(a+b)'" g145(.a(G27gat), .b(n84), .O(n230));
  "(ab)'"  g146(.a(n230), .b(n123), .O(n231));
  "!a"     g147(.a(n231), .O(n232));
  "(ab)'"  g148(.a(n232), .b(n229), .O(n233));
  "(ab)'"  g149(.a(n233), .b(n226), .O(n234));
  "(a+b)'" g150(.a(n132), .b(n203), .O(n237));
  "(a+b)'" g151(.a(G53gat), .b(n56), .O(n238));
  "(ab)'"  g152(.a(n238), .b(n185), .O(n239));
  "(a+b)'" g153(.a(n239), .b(n237), .O(n240));
  "(a+b)'" g154(.a(n138), .b(n203), .O(n243));
  "(a+b)'" g155(.a(G40gat), .b(n58), .O(n244));
  "(ab)'"  g156(.a(n244), .b(n189), .O(n245));
  "(a+b)'" g157(.a(n245), .b(n243), .O(n246));
  "(a+b)'" g158(.a(n246), .b(n240), .O(n247));
  "(a+b)'" g159(.a(n145), .b(n203), .O(n250));
  "(a+b)'" g160(.a(G79gat), .b(n61), .O(n251));
  "(ab)'"  g161(.a(n251), .b(n194), .O(n252));
  "(a+b)'" g162(.a(n252), .b(n250), .O(n253));
  "(a+b)'" g163(.a(n151), .b(n203), .O(n256));
  "(a+b)'" g164(.a(G66gat), .b(n63), .O(n257));
  "(ab)'"  g165(.a(n257), .b(n198), .O(n258));
  "(a+b)'" g166(.a(n258), .b(n256), .O(n259));
  "(a+b)'" g167(.a(n259), .b(n253), .O(n260));
  "(ab)'"  g168(.a(n260), .b(n247), .O(n261));
  "(a+b)'" g169(.a(n261), .b(n234), .O(n262));
  "(ab)'"  g170(.a(n262), .b(n219), .O(G370gat));
  "!a"     g171(.a(G14gat), .O(n264));
  "!a"     g172(.a(n171), .O(n265));
  "(a+b)'" g173(.a(n160), .b(n203), .O(n268));
  "(a+b)'" g174(.a(n208), .b(n268), .O(n269));
  "(a+b)'" g175(.a(n164), .b(n203), .O(n272));
  "(a+b)'" g176(.a(n215), .b(n272), .O(n273));
  "(a+b)'" g177(.a(n273), .b(n269), .O(n274));
  "(ab)'"  g178(.a(n274), .b(n265), .O(n275));
  "(a+b)'" g179(.a(n177), .b(n203), .O(n278));
  "(a+b)'" g180(.a(n224), .b(n278), .O(n279));
  "(a+b)'" g181(.a(n181), .b(n203), .O(n282));
  "(a+b)'" g182(.a(n231), .b(n282), .O(n283));
  "(a+b)'" g183(.a(n283), .b(n279), .O(n284));
  "(ab)'"  g184(.a(n186), .b(n204), .O(n287));
  "!a"     g185(.a(n239), .O(n288));
  "(ab)'"  g186(.a(n288), .b(n287), .O(n289));
  "(ab)'"  g187(.a(n190), .b(n204), .O(n292));
  "!a"     g188(.a(n245), .O(n293));
  "(ab)'"  g189(.a(n293), .b(n292), .O(n294));
  "(ab)'"  g190(.a(n294), .b(n289), .O(n295));
  "(ab)'"  g191(.a(n195), .b(n204), .O(n298));
  "!a"     g192(.a(n252), .O(n299));
  "(ab)'"  g193(.a(n299), .b(n298), .O(n300));
  "(ab)'"  g194(.a(n199), .b(n204), .O(n303));
  "!a"     g195(.a(n258), .O(n304));
  "(ab)'"  g196(.a(n304), .b(n303), .O(n305));
  "(ab)'"  g197(.a(n305), .b(n300), .O(n306));
  "(a+b)'" g198(.a(n306), .b(n295), .O(n307));
  "(ab)'"  g199(.a(n307), .b(n284), .O(n308));
  "(a+b)'" g200(.a(n308), .b(n275), .O(n309));
  "(a+b)'" g201(.a(n309), .b(n264), .O(n310));
  "(ab)'"  g202(.a(G329gat), .b(G8gat), .O(n311));
  "(a+b)'" g203(.a(n99), .b(n51), .O(n312));
  "(a+b)'" g204(.a(n312), .b(n82), .O(n313));
  "(ab)'"  g205(.a(n313), .b(n311), .O(n314));
  "(a+b)'" g206(.a(n314), .b(n310), .O(n315));
  "!a"     g207(.a(G66gat), .O(n316));
  "(a+b)'" g208(.a(n309), .b(n316), .O(n317));
  "(ab)'"  g209(.a(G329gat), .b(G60gat), .O(n318));
  "(a+b)'" g210(.a(n99), .b(n94), .O(n319));
  "(a+b)'" g211(.a(n319), .b(n63), .O(n320));
  "(ab)'"  g212(.a(n320), .b(n318), .O(n321));
  "(a+b)'" g213(.a(n321), .b(n317), .O(n322));
  "!a"     g214(.a(G53gat), .O(n323));
  "(a+b)'" g215(.a(n309), .b(n323), .O(n324));
  "(ab)'"  g216(.a(G329gat), .b(G47gat), .O(n325));
  "(a+b)'" g217(.a(n99), .b(n87), .O(n326));
  "(a+b)'" g218(.a(n326), .b(n56), .O(n327));
  "(ab)'"  g219(.a(n327), .b(n325), .O(n328));
  "(a+b)'" g220(.a(n328), .b(n324), .O(n329));
  "(a+b)'" g221(.a(n329), .b(n322), .O(n330));
  "!a"     g222(.a(G92gat), .O(n331));
  "(a+b)'" g223(.a(n309), .b(n331), .O(n332));
  "(ab)'"  g224(.a(G329gat), .b(G86gat), .O(n333));
  "(a+b)'" g225(.a(n99), .b(n47), .O(n334));
  "(a+b)'" g226(.a(n334), .b(n72), .O(n335));
  "(ab)'"  g227(.a(n335), .b(n333), .O(n336));
  "(a+b)'" g228(.a(n336), .b(n332), .O(n337));
  "!a"     g229(.a(G79gat), .O(n338));
  "(a+b)'" g230(.a(n309), .b(n338), .O(n339));
  "(ab)'"  g231(.a(G329gat), .b(G73gat), .O(n340));
  "(a+b)'" g232(.a(n99), .b(n92), .O(n341));
  "(a+b)'" g233(.a(n341), .b(n61), .O(n342));
  "(ab)'"  g234(.a(n342), .b(n340), .O(n343));
  "(a+b)'" g235(.a(n343), .b(n339), .O(n344));
  "(a+b)'" g236(.a(n344), .b(n337), .O(n345));
  "(ab)'"  g237(.a(n345), .b(n330), .O(n346));
  "!a"     g238(.a(G27gat), .O(n347));
  "(a+b)'" g239(.a(n309), .b(n347), .O(n348));
  "(ab)'"  g240(.a(G329gat), .b(G21gat), .O(n349));
  "(a+b)'" g241(.a(n99), .b(n53), .O(n350));
  "(a+b)'" g242(.a(n350), .b(n84), .O(n351));
  "(ab)'"  g243(.a(n351), .b(n349), .O(n352));
  "(a+b)'" g244(.a(n352), .b(n348), .O(n353));
  "!a"     g245(.a(G40gat), .O(n354));
  "(a+b)'" g246(.a(n309), .b(n354), .O(n355));
  "(ab)'"  g247(.a(G329gat), .b(G34gat), .O(n356));
  "(a+b)'" g248(.a(n99), .b(n89), .O(n357));
  "(a+b)'" g249(.a(n357), .b(n58), .O(n358));
  "(ab)'"  g250(.a(n358), .b(n356), .O(n359));
  "(a+b)'" g251(.a(n359), .b(n355), .O(n360));
  "(a+b)'" g252(.a(n360), .b(n353), .O(n361));
  "!a"     g253(.a(G115gat), .O(n362));
  "(a+b)'" g254(.a(n309), .b(n362), .O(n363));
  "(ab)'"  g255(.a(G329gat), .b(G112gat), .O(n364));
  "!a"     g256(.a(G102gat), .O(n365));
  "(a+b)'" g257(.a(n99), .b(n365), .O(n366));
  "(a+b)'" g258(.a(n366), .b(n43), .O(n367));
  "(ab)'"  g259(.a(n367), .b(n364), .O(n368));
  "(a+b)'" g260(.a(n368), .b(n363), .O(n369));
  "!a"     g261(.a(G105gat), .O(n370));
  "(a+b)'" g262(.a(n309), .b(n370), .O(n371));
  "(ab)'"  g263(.a(G329gat), .b(G99gat), .O(n372));
  "(a+b)'" g264(.a(n99), .b(n45), .O(n373));
  "(a+b)'" g265(.a(n373), .b(n70), .O(n374));
  "(ab)'"  g266(.a(n374), .b(n372), .O(n375));
  "(a+b)'" g267(.a(n375), .b(n371), .O(n376));
  "(a+b)'" g268(.a(n376), .b(n369), .O(n377));
  "(ab)'"  g269(.a(n377), .b(n361), .O(n378));
  "(a+b)'" g270(.a(n378), .b(n346), .O(n379));
  "(a+b)'" g271(.a(n379), .b(n315), .O(G421gat));
  "(ab)'"  g272(.a(G370gat), .b(G40gat), .O(n381));
  "!a"     g273(.a(n359), .O(n382));
  "(ab)'"  g274(.a(n382), .b(n381), .O(n383));
  "(ab)'"  g275(.a(n383), .b(n329), .O(n384));
  "(ab)'"  g276(.a(G370gat), .b(G27gat), .O(n385));
  "!a"     g277(.a(n352), .O(n386));
  "(ab)'"  g278(.a(n386), .b(n385), .O(n387));
  "(ab)'"  g279(.a(n383), .b(n387), .O(n388));
  "(a+b)'" g280(.a(n388), .b(n322), .O(n389));
  "(ab)'"  g281(.a(n389), .b(n384), .O(G430gat));
  "(a+b)'" g282(.a(n360), .b(n329), .O(n391));
  "(ab)'"  g283(.a(G370gat), .b(G79gat), .O(n392));
  "!a"     g284(.a(n343), .O(n393));
  "(ab)'"  g285(.a(n393), .b(n392), .O(n394));
  "(a+b)'" g286(.a(n394), .b(n322), .O(n395));
  "(ab)'"  g287(.a(n395), .b(n391), .O(n396));
  "(ab)'"  g288(.a(G370gat), .b(G66gat), .O(n397));
  "!a"     g289(.a(n321), .O(n398));
  "(ab)'"  g290(.a(n398), .b(n397), .O(n399));
  "(ab)'"  g291(.a(n337), .b(n399), .O(n400));
  "(a+b)'" g292(.a(n400), .b(n329), .O(n401));
  "(a+b)'" g293(.a(n401), .b(n388), .O(n402));
  "(ab)'"  g294(.a(n402), .b(n396), .O(G431gat));
  "(ab)'"  g295(.a(G370gat), .b(G105gat), .O(n404));
  "!a"     g296(.a(n375), .O(n405));
  "(ab)'"  g297(.a(n405), .b(n404), .O(n406));
  "(a+b)'" g298(.a(n406), .b(n337), .O(n407));
  "(ab)'"  g299(.a(n407), .b(n391), .O(n408));
  "(ab)'"  g300(.a(G370gat), .b(G53gat), .O(n409));
  "!a"     g301(.a(n328), .O(n410));
  "(ab)'"  g302(.a(n410), .b(n409), .O(n411));
  "(ab)'"  g303(.a(n383), .b(n411), .O(n412));
  "(ab)'"  g304(.a(n344), .b(n399), .O(n413));
  "(a+b)'" g305(.a(n413), .b(n412), .O(n414));
  "(ab)'"  g306(.a(n384), .b(n387), .O(n415));
  "(a+b)'" g307(.a(n415), .b(n414), .O(n416));
  "(ab)'"  g308(.a(n416), .b(n408), .O(G432gat));
endmodule


